
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module cr_kme_tlv_parser ( stitcher_rd, parser_kimreader_valid, 
	.parser_kimreader_data( {\parser_kimreader_data.sot [0], 
	\parser_kimreader_data.eoi [0], \parser_kimreader_data.eot [0], 
	\parser_kimreader_data.id [3], \parser_kimreader_data.id [2], 
	\parser_kimreader_data.id [1], \parser_kimreader_data.id [0], 
	\parser_kimreader_data.tdata [63], \parser_kimreader_data.tdata [62], 
	\parser_kimreader_data.tdata [61], \parser_kimreader_data.tdata [60], 
	\parser_kimreader_data.tdata [59], \parser_kimreader_data.tdata [58], 
	\parser_kimreader_data.tdata [57], \parser_kimreader_data.tdata [56], 
	\parser_kimreader_data.tdata [55], \parser_kimreader_data.tdata [54], 
	\parser_kimreader_data.tdata [53], \parser_kimreader_data.tdata [52], 
	\parser_kimreader_data.tdata [51], \parser_kimreader_data.tdata [50], 
	\parser_kimreader_data.tdata [49], \parser_kimreader_data.tdata [48], 
	\parser_kimreader_data.tdata [47], \parser_kimreader_data.tdata [46], 
	\parser_kimreader_data.tdata [45], \parser_kimreader_data.tdata [44], 
	\parser_kimreader_data.tdata [43], \parser_kimreader_data.tdata [42], 
	\parser_kimreader_data.tdata [41], \parser_kimreader_data.tdata [40], 
	\parser_kimreader_data.tdata [39], \parser_kimreader_data.tdata [38], 
	\parser_kimreader_data.tdata [37], \parser_kimreader_data.tdata [36], 
	\parser_kimreader_data.tdata [35], \parser_kimreader_data.tdata [34], 
	\parser_kimreader_data.tdata [33], \parser_kimreader_data.tdata [32], 
	\parser_kimreader_data.tdata [31], \parser_kimreader_data.tdata [30], 
	\parser_kimreader_data.tdata [29], \parser_kimreader_data.tdata [28], 
	\parser_kimreader_data.tdata [27], \parser_kimreader_data.tdata [26], 
	\parser_kimreader_data.tdata [25], \parser_kimreader_data.tdata [24], 
	\parser_kimreader_data.tdata [23], \parser_kimreader_data.tdata [22], 
	\parser_kimreader_data.tdata [21], \parser_kimreader_data.tdata [20], 
	\parser_kimreader_data.tdata [19], \parser_kimreader_data.tdata [18], 
	\parser_kimreader_data.tdata [17], \parser_kimreader_data.tdata [16], 
	\parser_kimreader_data.tdata [15], \parser_kimreader_data.tdata [14], 
	\parser_kimreader_data.tdata [13], \parser_kimreader_data.tdata [12], 
	\parser_kimreader_data.tdata [11], \parser_kimreader_data.tdata [10], 
	\parser_kimreader_data.tdata [9], \parser_kimreader_data.tdata [8], 
	\parser_kimreader_data.tdata [7], \parser_kimreader_data.tdata [6], 
	\parser_kimreader_data.tdata [5], \parser_kimreader_data.tdata [4], 
	\parser_kimreader_data.tdata [3], \parser_kimreader_data.tdata [2], 
	\parser_kimreader_data.tdata [1], \parser_kimreader_data.tdata [0]} ), 
	tlv_parser_idle, tlv_parser_int_tlv_start_pulse, clk, rst_n, 
	disable_debug_cmd_q, always_validate_kim_ref, .stitcher_out( {
	\stitcher_out.tvalid , \stitcher_out.tlast , \stitcher_out.tid [0], 
	\stitcher_out.tstrb [7], \stitcher_out.tstrb [6], 
	\stitcher_out.tstrb [5], \stitcher_out.tstrb [4], 
	\stitcher_out.tstrb [3], \stitcher_out.tstrb [2], 
	\stitcher_out.tstrb [1], \stitcher_out.tstrb [0], 
	\stitcher_out.tuser [7], \stitcher_out.tuser [6], 
	\stitcher_out.tuser [5], \stitcher_out.tuser [4], 
	\stitcher_out.tuser [3], \stitcher_out.tuser [2], 
	\stitcher_out.tuser [1], \stitcher_out.tuser [0], 
	\stitcher_out.tdata [63], \stitcher_out.tdata [62], 
	\stitcher_out.tdata [61], \stitcher_out.tdata [60], 
	\stitcher_out.tdata [59], \stitcher_out.tdata [58], 
	\stitcher_out.tdata [57], \stitcher_out.tdata [56], 
	\stitcher_out.tdata [55], \stitcher_out.tdata [54], 
	\stitcher_out.tdata [53], \stitcher_out.tdata [52], 
	\stitcher_out.tdata [51], \stitcher_out.tdata [50], 
	\stitcher_out.tdata [49], \stitcher_out.tdata [48], 
	\stitcher_out.tdata [47], \stitcher_out.tdata [46], 
	\stitcher_out.tdata [45], \stitcher_out.tdata [44], 
	\stitcher_out.tdata [43], \stitcher_out.tdata [42], 
	\stitcher_out.tdata [41], \stitcher_out.tdata [40], 
	\stitcher_out.tdata [39], \stitcher_out.tdata [38], 
	\stitcher_out.tdata [37], \stitcher_out.tdata [36], 
	\stitcher_out.tdata [35], \stitcher_out.tdata [34], 
	\stitcher_out.tdata [33], \stitcher_out.tdata [32], 
	\stitcher_out.tdata [31], \stitcher_out.tdata [30], 
	\stitcher_out.tdata [29], \stitcher_out.tdata [28], 
	\stitcher_out.tdata [27], \stitcher_out.tdata [26], 
	\stitcher_out.tdata [25], \stitcher_out.tdata [24], 
	\stitcher_out.tdata [23], \stitcher_out.tdata [22], 
	\stitcher_out.tdata [21], \stitcher_out.tdata [20], 
	\stitcher_out.tdata [19], \stitcher_out.tdata [18], 
	\stitcher_out.tdata [17], \stitcher_out.tdata [16], 
	\stitcher_out.tdata [15], \stitcher_out.tdata [14], 
	\stitcher_out.tdata [13], \stitcher_out.tdata [12], 
	\stitcher_out.tdata [11], \stitcher_out.tdata [10], 
	\stitcher_out.tdata [9], \stitcher_out.tdata [8], 
	\stitcher_out.tdata [7], \stitcher_out.tdata [6], 
	\stitcher_out.tdata [5], \stitcher_out.tdata [4], 
	\stitcher_out.tdata [3], \stitcher_out.tdata [2], 
	\stitcher_out.tdata [1], \stitcher_out.tdata [0]} ), stitcher_empty, 
	kimreader_parser_ack);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output stitcher_rd;
output parser_kimreader_valid;
output [0:0] \parser_kimreader_data.sot ;
output [0:0] \parser_kimreader_data.eoi ;
output [0:0] \parser_kimreader_data.eot ;
output [3:0] \parser_kimreader_data.id ;
output [63:0] \parser_kimreader_data.tdata ;
wire [70:0] parser_kimreader_data;
output tlv_parser_idle;
output tlv_parser_int_tlv_start_pulse;
input clk;
input rst_n;
input disable_debug_cmd_q;
input always_validate_kim_ref;
input \stitcher_out.tvalid ;
input \stitcher_out.tlast ;
input [0:0] \stitcher_out.tid ;
input [7:0] \stitcher_out.tstrb ;
input [7:0] \stitcher_out.tuser ;
input [63:0] \stitcher_out.tdata ;
wire [82:0] stitcher_out;
input stitcher_empty;
input kimreader_parser_ack;
wire fifo_in_stall;
wire stitcher_sot;
wire stitcher_eot;
wire _zy_simnet_stitcher_rd_0_w$;
wire [0:70] _zy_simnet_parser_kimreader_data_1_w$;
wire [0:70] _zy_simnet_parser_kimreader_data_2_w$;
wire _zy_simnet_dio_3;
wire _zy_simnet_dio_4;
wire [0:70] _zy_simnet_fifo_in_5_w$;
wire _zy_simnet_fifo_in_valid_6_w$;
wire _zy_simnet_cio_7;
wire _zy_sva_key_type0_line4_1_reset_or;
wire _zy_sva_key_type0_line5a_2_reset_or;
wire _zy_sva_key_type0_line5b_3_reset_or;
wire _zy_sva_key_type1_line7a_4_reset_or;
wire _zy_sva_key_type1_line7b_5_reset_or;
wire _zy_sva_key_type1_line8a_6_reset_or;
wire _zy_sva_key_type1_line8b_7_reset_or;
wire _zy_sva_key_type1_line9_8_reset_or;
wire _zy_sva_key_type1_line10_9_reset_or;
wire _zy_sva_key_type1_line11a_10_reset_or;
wire _zy_sva_key_type1_line11b_11_reset_or;
wire _zy_sva_key_type1_line11c_12_reset_or;
wire _zy_sva_key_type1_line11d_13_reset_or;
wire _zy_sva_key_type1_line12a_14_reset_or;
wire _zy_sva_key_type1_line12b_15_reset_or;
wire _zy_sva_key_type9_line14_16_reset_or;
wire _zy_sva_key_type9_line15_17_reset_or;
wire _zy_sva_key_type9_line16a_18_reset_or;
wire _zy_sva_key_type9_line16b_19_reset_or;
wire _zy_sva_key_type9_line17a_20_reset_or;
wire _zy_sva_key_type9_line17b_21_reset_or;
wire _zy_sva_key_type9_line18a_22_reset_or;
wire _zy_sva_key_type9_line18b_23_reset_or;
wire _zy_sva_key_type9_line19a_24_reset_or;
wire _zy_sva_key_type9_line19b_25_reset_or;
wire _zy_sva_key_type9_line19c_26_reset_or;
wire _zy_sva_key_type9_line19d_27_reset_or;
wire _zy_sva_guid_miss_aux_cmd_0_28_reset_or;
wire _zy_sva_guid_miss_aux_cmd_1_29_reset_or;
wire _zy_sva_guid_miss_aux_cmd_2_30_reset_or;
wire _zy_sva_guid_miss_aux_cmd_3_31_reset_or;
wire _zy_sva_guid_miss_aux_cmd_iv_0_32_reset_or;
wire _zy_sva_guid_miss_aux_cmd_iv_1_33_reset_or;
wire _zy_sva_guid_miss_aux_cmd_iv_2_34_reset_or;
wire _zy_sva_guid_miss_aux_cmd_iv_3_35_reset_or;
wire _zy_sva_iv_miss_aux_cmd_0_36_reset_or;
wire _zy_sva_iv_miss_aux_cmd_1_37_reset_or;
wire _zy_sva_iv_miss_aux_cmd_guid_38_reset_or;
wire _zy_sva_brcm_aux_cmd_39_reset_or;
wire _zy_sva_brcm_aux_cmd_iv_40_reset_or;
wire _zy_sva_brcm_aux_cmd_guid_41_reset_or;
wire _zy_sva_brcm_aux_cmd_guid_iv_42_reset_or;
wire _zy_sva_brcm_key_type_43_reset_or;
wire _zy_sva_brcm_aux_cmd_44_reset_or;
wire _zy_sva_brcm_aux_cmd_iv_45_reset_or;
wire _zy_sva_brcm_aux_cmd_guid_46_reset_or;
wire _zy_sva_brcm_aux_cmd_guid_iv_47_reset_or;
wire _zy_sva_brcm_key_type_48_reset_or;
wire _zy_sva_brcm_aux_cmd_49_reset_or;
wire _zy_sva_brcm_aux_cmd_iv_50_reset_or;
wire _zy_sva_brcm_aux_cmd_guid_51_reset_or;
wire _zy_sva_brcm_aux_cmd_guid_iv_52_reset_or;
wire _zy_sva_brcm_key_type_53_reset_or;
wire _zy_sva_brcm_aux_cmd_54_reset_or;
wire _zy_sva_brcm_aux_cmd_iv_55_reset_or;
wire _zy_sva_brcm_aux_cmd_guid_56_reset_or;
wire _zy_sva_brcm_aux_cmd_guid_iv_57_reset_or;
wire _zy_sva_brcm_key_type_58_reset_or;
wire _zy_sva_brcm_aux_cmd_59_reset_or;
wire _zy_sva_brcm_aux_cmd_iv_60_reset_or;
wire _zy_sva_brcm_aux_cmd_guid_61_reset_or;
wire _zy_sva_brcm_aux_cmd_guid_iv_62_reset_or;
wire _zy_sva_brcm_key_type_63_reset_or;
wire _zy_sva_brcm_aux_cmd_64_reset_or;
wire _zy_sva_brcm_aux_cmd_iv_65_reset_or;
wire _zy_sva_brcm_aux_cmd_guid_66_reset_or;
wire _zy_sva_brcm_aux_cmd_guid_iv_67_reset_or;
wire _zy_sva_brcm_key_type_68_reset_or;
wire _zy_sva_brcm_aux_cmd_69_reset_or;
wire _zy_sva_brcm_aux_cmd_iv_70_reset_or;
wire _zy_sva_brcm_aux_cmd_guid_71_reset_or;
wire _zy_sva_brcm_aux_cmd_guid_iv_72_reset_or;
wire _zy_sva_brcm_key_type_73_reset_or;
wire _zy_sva_brcm_aux_cmd_74_reset_or;
wire _zy_sva_brcm_aux_cmd_iv_75_reset_or;
wire _zy_sva_brcm_aux_cmd_guid_76_reset_or;
wire _zy_sva_brcm_aux_cmd_guid_iv_77_reset_or;
wire _zy_sva_brcm_key_type_78_reset_or;
wire _zy_sva_brcm_aux_cmd_79_reset_or;
wire _zy_sva_brcm_aux_cmd_iv_80_reset_or;
wire _zy_sva_brcm_aux_cmd_guid_81_reset_or;
wire _zy_sva_brcm_aux_cmd_guid_iv_82_reset_or;
wire _zy_sva_brcm_key_type_83_reset_or;
wire _zy_sva_brcm_aux_cmd_84_reset_or;
wire _zy_sva_brcm_aux_cmd_iv_85_reset_or;
wire _zy_sva_brcm_aux_cmd_guid_86_reset_or;
wire _zy_sva_brcm_aux_cmd_guid_iv_87_reset_or;
wire _zy_sva_brcm_key_type_88_reset_or;
wire _zy_sva_brcm_aux_cmd_89_reset_or;
wire _zy_sva_brcm_aux_cmd_iv_90_reset_or;
wire _zy_sva_brcm_aux_cmd_guid_91_reset_or;
wire _zy_sva_brcm_aux_cmd_guid_iv_92_reset_or;
wire _zy_sva_brcm_key_type_93_reset_or;
wire _zy_sva_brcm_aux_cmd_94_reset_or;
wire _zy_sva_brcm_aux_cmd_iv_95_reset_or;
wire _zy_sva_brcm_aux_cmd_guid_96_reset_or;
wire _zy_sva_brcm_aux_cmd_guid_iv_97_reset_or;
wire _zy_sva_brcm_key_type_98_reset_or;
wire _zy_sva_brcm_aux_cmd_99_reset_or;
wire _zy_sva_brcm_aux_cmd_iv_100_reset_or;
wire _zy_sva_brcm_aux_cmd_guid_101_reset_or;
wire _zy_sva_brcm_aux_cmd_guid_iv_102_reset_or;
wire _zy_sva_brcm_key_type_103_reset_or;
wire _zy_sva_brcm_aux_cmd_104_reset_or;
wire _zy_sva_brcm_aux_cmd_iv_105_reset_or;
wire _zy_sva_brcm_aux_cmd_guid_106_reset_or;
wire _zy_sva_brcm_aux_cmd_guid_iv_107_reset_or;
wire _zy_sva_brcm_key_type_108_reset_or;
wire _zy_sva_brcm_kdf_ops_109_reset_or;
wire _zy_sva_brcm_kdf_ops_110_reset_or;
wire _zy_sva_brcm_kdf_ops_111_reset_or;
wire _zy_sva_brcm_kdf_ops_112_reset_or;
wire _zy_sva_brcm_kdf_ops_113_reset_or;
wire _zy_sva_brcm_kdf_ops_114_reset_or;
wire _zy_sva_brcm_kdf_ops_115_reset_or;
wire _zy_sva_brcm_kdf_ops_116_reset_or;
wire _zy_sva_brcm_kdf_ops_117_reset_or;
wire _zy_sva_brcm_kdf_ops_118_reset_or;
wire _zy_sva_brcm_kdf_ops_119_reset_or;
wire _zy_sva_brcm_kdf_ops_120_reset_or;
wire _zy_sva_brcm_kdf_ops_121_reset_or;
wire _zy_sva_brcm_kdf_ops_122_reset_or;
wire _zy_sva_brcm_kdf_ops_123_reset_or;
wire _zy_sva_brcm_kdf_ops_124_reset_or;
wire _zy_sva_null_gcm_125_reset_or;
wire _zy_sva_sha_gcm_126_reset_or;
wire _zy_sva_null_xts_127_reset_or;
wire _zy_sva_sha_xts_128_reset_or;
wire _zy_sva_null_null_129_reset_or;
wire _zy_sva_sha_null_130_reset_or;
wire _zy_sva_hmac_gcm_131_reset_or;
wire _zy_sva_hmac_xts_132_reset_or;
wire _zy_sva_hmac_null_133_reset_or;
wire _zy_sva_null_gcm_134_reset_or;
wire _zy_sva_sha_gcm_135_reset_or;
wire _zy_sva_null_xts_136_reset_or;
wire _zy_sva_sha_xts_137_reset_or;
wire _zy_sva_null_null_138_reset_or;
wire _zy_sva_sha_null_139_reset_or;
wire _zy_sva_hmac_gcm_140_reset_or;
wire _zy_sva_hmac_xts_141_reset_or;
wire _zy_sva_hmac_null_142_reset_or;
wire _zy_sva_null_gcm_143_reset_or;
wire _zy_sva_sha_gcm_144_reset_or;
wire _zy_sva_null_xts_145_reset_or;
wire _zy_sva_sha_xts_146_reset_or;
wire _zy_sva_null_null_147_reset_or;
wire _zy_sva_sha_null_148_reset_or;
wire _zy_sva_hmac_gcm_149_reset_or;
wire _zy_sva_hmac_xts_150_reset_or;
wire _zy_sva_hmac_null_151_reset_or;
wire _zy_sva_null_gcm_152_reset_or;
wire _zy_sva_sha_gcm_153_reset_or;
wire _zy_sva_null_xts_154_reset_or;
wire _zy_sva_sha_xts_155_reset_or;
wire _zy_sva_null_null_156_reset_or;
wire _zy_sva_sha_null_157_reset_or;
wire _zy_sva_hmac_gcm_158_reset_or;
wire _zy_sva_hmac_xts_159_reset_or;
wire _zy_sva_hmac_null_160_reset_or;
wire _zy_sva_null_gcm_161_reset_or;
wire _zy_sva_sha_gcm_162_reset_or;
wire _zy_sva_null_xts_163_reset_or;
wire _zy_sva_sha_xts_164_reset_or;
wire _zy_sva_null_null_165_reset_or;
wire _zy_sva_sha_null_166_reset_or;
wire _zy_sva_hmac_gcm_167_reset_or;
wire _zy_sva_hmac_xts_168_reset_or;
wire _zy_sva_hmac_null_169_reset_or;
wire _zy_sva_null_gcm_170_reset_or;
wire _zy_sva_sha_gcm_171_reset_or;
wire _zy_sva_null_xts_172_reset_or;
wire _zy_sva_sha_xts_173_reset_or;
wire _zy_sva_null_null_174_reset_or;
wire _zy_sva_sha_null_175_reset_or;
wire _zy_sva_hmac_gcm_176_reset_or;
wire _zy_sva_hmac_xts_177_reset_or;
wire _zy_sva_hmac_null_178_reset_or;
wire _zy_sva_b0_t;
wire _zy_sva_b1_t;
wire _zy_sva_b2_t;
wire _zy_sva_b3_t;
wire _zy_sva_b4_t;
wire _zy_sva_b5_t;
wire _zy_sva_b6_t;
wire _zy_sva_b7_t;
wire _zy_sva_b8_t;
wire _zy_sva_b9_t;
wire _zy_sva_b10_t;
wire _zy_sva_b11_t;
wire _zy_sva_b12_t;
wire _zy_sva_b13_t;
wire _zy_sva_b14_t;
wire _zy_sva_b15_t;
wire _zy_sva_b16_t;
wire _zy_sva_b17_t;
wire _zy_sva_b18_t;
wire _zy_sva_b19_t;
wire _zy_sva_b20_t;
wire _zy_sva_b21_t;
wire _zy_sva_b22_t;
wire _zy_sva_b23_t;
wire _zy_sva_b24_t;
wire _zy_sva_b25_t;
wire _zy_sva_b26_t;
wire _zy_sva_b27_t;
wire _zy_sva_b28_t;
wire _zy_sva_b29_t;
wire _zy_sva_b30_t;
wire _zy_sva_b31_t;
wire _zy_sva_b32_t;
wire _zy_sva_b33_t;
wire _zy_sva_b34_t;
wire _zy_sva_b35_t;
wire _zy_sva_b36_t;
wire _zy_sva_b37_t;
wire _zy_sva_b38_t;
wire _zy_sva_b39_t;
wire _zy_sva_b40_t;
wire _zy_sva_b41_t;
wire _zy_sva_b42_t;
wire _zy_sva_b43_t;
wire _zy_sva_b44_t;
wire _zy_sva_b45_t;
wire _zy_sva_b46_t;
wire _zy_sva_b47_t;
wire _zy_sva_b48_t;
wire _zy_sva_b49_t;
wire _zy_sva_b50_t;
wire _zy_sva_b51_t;
wire _zy_sva_b52_t;
wire _zy_sva_b53_t;
wire _zy_sva_b54_t;
wire _zy_sva_b55_t;
wire _zy_sva_b56_t;
wire _zy_sva_b57_t;
wire _zy_sva_b58_t;
wire _zy_sva_b59_t;
wire _zy_sva_b60_t;
wire _zy_sva_b61_t;
wire _zy_sva_b62_t;
wire _zy_sva_b63_t;
wire _zy_sva_b64_t;
wire _zy_sva_b65_t;
wire _zy_sva_b66_t;
wire _zy_sva_b67_t;
wire _zy_sva_b68_t;
wire _zy_sva_b69_t;
wire _zy_sva_b70_t;
wire _zy_sva_b71_t;
wire _zy_sva_b72_t;
wire _zy_sva_b73_t;
wire _zy_sva_b74_t;
wire _zy_sva_b75_t;
wire _zy_sva_b76_t;
wire _zy_sva_b77_t;
wire _zy_sva_b78_t;
wire _zy_sva_b79_t;
wire _zy_sva_b80_t;
wire _zy_sva_b81_t;
wire _zy_sva_b82_t;
wire _zy_sva_b83_t;
wire _zy_sva_b84_t;
wire _zy_sva_b85_t;
wire _zy_sva_b86_t;
wire _zy_sva_b87_t;
wire _zy_sva_b88_t;
wire _zy_sva_b89_t;
wire _zy_sva_b90_t;
wire _zy_sva_b91_t;
wire _zy_sva_b92_t;
wire _zy_sva_b93_t;
wire _zy_sva_b94_t;
wire _zy_sva_b95_t;
wire _zy_sva_b96_t;
wire _zy_sva_b97_t;
wire _zy_sva_b98_t;
wire _zy_sva_b99_t;
wire _zy_sva_b100_t;
wire _zy_sva_b101_t;
wire _zy_sva_b102_t;
wire _zy_sva_b103_t;
wire _zy_sva_b104_t;
wire _zy_sva_b105_t;
wire _zy_sva_b106_t;
wire _zy_sva_b107_t;
wire _zy_sva_b108_t;
wire _zy_sva_b109_t;
wire _zy_sva_b110_t;
wire _zy_sva_b111_t;
wire _zy_sva_b112_t;
wire _zy_sva_b113_t;
wire _zy_sva_b114_t;
wire _zy_sva_b115_t;
wire _zy_sva_b116_t;
wire _zy_sva_b117_t;
wire _zy_sva_b118_t;
wire _zy_sva_b119_t;
wire _zy_sva_b120_t;
wire _zy_sva_b121_t;
wire _zy_sva_b122_t;
wire _zy_sva_b123_t;
wire _zy_sva_b124_t;
wire _zy_sva_b125_t;
wire _zy_sva_b126_t;
wire _zy_sva_b127_t;
wire _zy_sva_b128_t;
wire _zy_sva_b129_t;
wire _zy_sva_b130_t;
wire _zy_sva_b131_t;
wire _zy_sva_b132_t;
wire _zy_sva_b133_t;
wire _zy_sva_b134_t;
wire _zy_sva_b135_t;
wire _zy_sva_b136_t;
wire _zy_sva_b137_t;
wire _zy_sva_b138_t;
wire _zy_sva_b139_t;
wire _zy_sva_b140_t;
wire _zy_sva_b141_t;
wire _zy_sva_b142_t;
wire _zy_sva_b143_t;
wire _zy_sva_b144_t;
wire _zy_sva_b145_t;
wire _zy_sva_b146_t;
wire _zy_sva_b147_t;
wire _zy_sva_b148_t;
wire _zy_sva_b149_t;
wire _zy_sva_b150_t;
wire _zy_sva_b151_t;
wire _zy_sva_b152_t;
wire _zy_sva_b153_t;
wire _zy_sva_b154_t;
wire _zy_sva_b155_t;
wire _zy_sva_b156_t;
wire _zy_sva_b157_t;
wire _zy_sva_b158_t;
wire _zy_sva_b159_t;
wire _zy_sva_b160_t;
wire _zy_sva_b161_t;
wire _zy_sva_b162_t;
wire _zy_sva_b163_t;
wire _zy_sva_b164_t;
wire _zy_sva_b165_t;
wire _zy_sva_b166_t;
wire _zy_sva_b167_t;
wire _zy_sva_b168_t;
wire _zy_sva_b169_t;
wire _zy_sva_b170_t;
wire _zy_sva_b171_t;
wire _zy_sva_b172_t;
wire _zy_sva_b173_t;
wire _zy_sva_b174_t;
wire _zy_sva_b175_t;
wire _zy_sva_b176_t;
wire _zy_sva_b177_t;
wire [70:0] fifo_in;
wire fifo_in_valid;
wire key_blob_region;
wire [5:0] int_tlv_counter;
wire [4:0] tlv_counter;
wire [63:0] tlv_word0;
wire [63:0] tlv_word1;
wire [63:0] tlv_word2;
wire [3:0] nxt_fifo_in_id;
wire [63:0] frame_word;
wire [63:0] kme_internal_word0;
wire [63:0] nxt_kme_internal_word0;
wire [63:0] kme_internal_dek_kim_word;
wire [63:0] nxt_kme_internal_dek_kim_word;
wire [63:0] kme_internal_dak_kim_word;
wire [63:0] nxt_kme_internal_dak_kim_word;
wire [7:0] tlv_type;
wire [7:0] nxt_tlv_type;
wire [5:0] aux_key_type;
wire [5:0] nxt_aux_key_type;
wire [1:0] aux_iv_op;
wire [1:0] nxt_aux_iv_op;
wire [3:0] aux_cipher_op;
wire [3:0] nxt_aux_cipher_op;
wire [3:0] aux_auth_op;
wire [3:0] nxt_aux_auth_op;
wire [3:0] aux_raw_auth_op;
wire [3:0] nxt_aux_raw_auth_op;
wire [31:0] debug_cmd;
wire [31:0] nxt_debug_cmd;
wire [31:0] aux_key_header;
wire [31:0] nxt_aux_key_header;
wire [6:0] skip;
wire [6:0] nxt_skip;
wire [63:0] guid0;
wire [63:0] nxt_guid0;
wire [63:0] guid1;
wire [63:0] nxt_guid1;
wire [63:0] guid2;
wire [63:0] nxt_guid2;
wire [63:0] guid3;
wire [63:0] nxt_guid3;
wire [63:0] iv0;
wire [63:0] nxt_iv0;
wire [63:0] iv1;
wire [63:0] nxt_iv1;
wire [31:0] buffer;
wire [31:0] nxt_buffer;
`_2_ wire [0:0] _zy_sva_key_type0_line4_1_ccheck;
`_2_ wire [0:0] _zy_sva_key_type0_line4_1_cpass;
`_2_ wire _zy_sva_b0;
`_2_ wire [0:0] _zy_sva_key_type0_line5a_2_ccheck;
`_2_ wire [0:0] _zy_sva_key_type0_line5a_2_cpass;
`_2_ wire _zy_sva_b1;
`_2_ wire [0:0] _zy_sva_key_type0_line5b_3_ccheck;
`_2_ wire [0:0] _zy_sva_key_type0_line5b_3_cpass;
`_2_ wire _zy_sva_b2;
`_2_ wire [0:0] _zy_sva_key_type1_line7a_4_ccheck;
`_2_ wire [0:0] _zy_sva_key_type1_line7a_4_cpass;
`_2_ wire _zy_sva_b3;
`_2_ wire [0:0] _zy_sva_key_type1_line7b_5_ccheck;
`_2_ wire [0:0] _zy_sva_key_type1_line7b_5_cpass;
`_2_ wire _zy_sva_b4;
`_2_ wire [0:0] _zy_sva_key_type1_line8a_6_ccheck;
`_2_ wire [0:0] _zy_sva_key_type1_line8a_6_cpass;
`_2_ wire _zy_sva_b5;
`_2_ wire [0:0] _zy_sva_key_type1_line8b_7_ccheck;
`_2_ wire [0:0] _zy_sva_key_type1_line8b_7_cpass;
`_2_ wire _zy_sva_b6;
`_2_ wire [0:0] _zy_sva_key_type1_line9_8_ccheck;
`_2_ wire [0:0] _zy_sva_key_type1_line9_8_cpass;
`_2_ wire _zy_sva_b7;
`_2_ wire [0:0] _zy_sva_key_type1_line10_9_ccheck;
`_2_ wire [0:0] _zy_sva_key_type1_line10_9_cpass;
`_2_ wire _zy_sva_b8;
`_2_ wire [0:0] _zy_sva_key_type1_line11a_10_ccheck;
`_2_ wire [0:0] _zy_sva_key_type1_line11a_10_cpass;
`_2_ wire _zy_sva_b9;
`_2_ wire [0:0] _zy_sva_key_type1_line11b_11_ccheck;
`_2_ wire [0:0] _zy_sva_key_type1_line11b_11_cpass;
`_2_ wire _zy_sva_b10;
`_2_ wire [0:0] _zy_sva_key_type1_line11c_12_ccheck;
`_2_ wire [0:0] _zy_sva_key_type1_line11c_12_cpass;
`_2_ wire _zy_sva_b11;
`_2_ wire [0:0] _zy_sva_key_type1_line11d_13_ccheck;
`_2_ wire [0:0] _zy_sva_key_type1_line11d_13_cpass;
`_2_ wire _zy_sva_b12;
`_2_ wire [0:0] _zy_sva_key_type1_line12a_14_ccheck;
`_2_ wire [0:0] _zy_sva_key_type1_line12a_14_cpass;
`_2_ wire _zy_sva_b13;
`_2_ wire [0:0] _zy_sva_key_type1_line12b_15_ccheck;
`_2_ wire [0:0] _zy_sva_key_type1_line12b_15_cpass;
`_2_ wire _zy_sva_b14;
`_2_ wire [0:0] _zy_sva_key_type9_line14_16_ccheck;
`_2_ wire [0:0] _zy_sva_key_type9_line14_16_cpass;
`_2_ wire _zy_sva_b15;
`_2_ wire [0:0] _zy_sva_key_type9_line15_17_ccheck;
`_2_ wire [0:0] _zy_sva_key_type9_line15_17_cpass;
`_2_ wire _zy_sva_b16;
`_2_ wire [0:0] _zy_sva_key_type9_line16a_18_ccheck;
`_2_ wire [0:0] _zy_sva_key_type9_line16a_18_cpass;
`_2_ wire _zy_sva_b17;
`_2_ wire [0:0] _zy_sva_key_type9_line16b_19_ccheck;
`_2_ wire [0:0] _zy_sva_key_type9_line16b_19_cpass;
`_2_ wire _zy_sva_b18;
`_2_ wire [0:0] _zy_sva_key_type9_line17a_20_ccheck;
`_2_ wire [0:0] _zy_sva_key_type9_line17a_20_cpass;
`_2_ wire _zy_sva_b19;
`_2_ wire [0:0] _zy_sva_key_type9_line17b_21_ccheck;
`_2_ wire [0:0] _zy_sva_key_type9_line17b_21_cpass;
`_2_ wire _zy_sva_b20;
`_2_ wire [0:0] _zy_sva_key_type9_line18a_22_ccheck;
`_2_ wire [0:0] _zy_sva_key_type9_line18a_22_cpass;
`_2_ wire _zy_sva_b21;
`_2_ wire [0:0] _zy_sva_key_type9_line18b_23_ccheck;
`_2_ wire [0:0] _zy_sva_key_type9_line18b_23_cpass;
`_2_ wire _zy_sva_b22;
`_2_ wire [0:0] _zy_sva_key_type9_line19a_24_ccheck;
`_2_ wire [0:0] _zy_sva_key_type9_line19a_24_cpass;
`_2_ wire _zy_sva_b23;
`_2_ wire [0:0] _zy_sva_key_type9_line19b_25_ccheck;
`_2_ wire [0:0] _zy_sva_key_type9_line19b_25_cpass;
`_2_ wire _zy_sva_b24;
`_2_ wire [0:0] _zy_sva_key_type9_line19c_26_ccheck;
`_2_ wire [0:0] _zy_sva_key_type9_line19c_26_cpass;
`_2_ wire _zy_sva_b25;
`_2_ wire [0:0] _zy_sva_key_type9_line19d_27_ccheck;
`_2_ wire [0:0] _zy_sva_key_type9_line19d_27_cpass;
`_2_ wire _zy_sva_b26;
`_2_ wire [0:0] _zy_sva_guid_miss_aux_cmd_0_28_ccheck;
`_2_ wire [0:0] _zy_sva_guid_miss_aux_cmd_0_28_cpass;
`_2_ wire _zy_sva_b27;
`_2_ wire [0:0] _zy_sva_guid_miss_aux_cmd_1_29_ccheck;
`_2_ wire [0:0] _zy_sva_guid_miss_aux_cmd_1_29_cpass;
`_2_ wire _zy_sva_b28;
`_2_ wire [0:0] _zy_sva_guid_miss_aux_cmd_2_30_ccheck;
`_2_ wire [0:0] _zy_sva_guid_miss_aux_cmd_2_30_cpass;
`_2_ wire _zy_sva_b29;
`_2_ wire [0:0] _zy_sva_guid_miss_aux_cmd_3_31_ccheck;
`_2_ wire [0:0] _zy_sva_guid_miss_aux_cmd_3_31_cpass;
`_2_ wire _zy_sva_b30;
`_2_ wire [0:0] _zy_sva_guid_miss_aux_cmd_iv_0_32_ccheck;
`_2_ wire [0:0] _zy_sva_guid_miss_aux_cmd_iv_0_32_cpass;
`_2_ wire _zy_sva_b31;
`_2_ wire [0:0] _zy_sva_guid_miss_aux_cmd_iv_1_33_ccheck;
`_2_ wire [0:0] _zy_sva_guid_miss_aux_cmd_iv_1_33_cpass;
`_2_ wire _zy_sva_b32;
`_2_ wire [0:0] _zy_sva_guid_miss_aux_cmd_iv_2_34_ccheck;
`_2_ wire [0:0] _zy_sva_guid_miss_aux_cmd_iv_2_34_cpass;
`_2_ wire _zy_sva_b33;
`_2_ wire [0:0] _zy_sva_guid_miss_aux_cmd_iv_3_35_ccheck;
`_2_ wire [0:0] _zy_sva_guid_miss_aux_cmd_iv_3_35_cpass;
`_2_ wire _zy_sva_b34;
`_2_ wire [0:0] _zy_sva_iv_miss_aux_cmd_0_36_ccheck;
`_2_ wire [0:0] _zy_sva_iv_miss_aux_cmd_0_36_cpass;
`_2_ wire _zy_sva_b35;
`_2_ wire [0:0] _zy_sva_iv_miss_aux_cmd_1_37_ccheck;
`_2_ wire [0:0] _zy_sva_iv_miss_aux_cmd_1_37_cpass;
`_2_ wire _zy_sva_b36;
`_2_ wire [0:0] _zy_sva_iv_miss_aux_cmd_guid_38_ccheck;
`_2_ wire [0:0] _zy_sva_iv_miss_aux_cmd_guid_38_cpass;
`_2_ wire _zy_sva_b37;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_39_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_39_cpass;
`_2_ wire _zy_sva_b38;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_iv_40_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_iv_40_cpass;
`_2_ wire _zy_sva_b39;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_41_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_41_cpass;
`_2_ wire _zy_sva_b40;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_iv_42_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_iv_42_cpass;
`_2_ wire _zy_sva_b41;
`_2_ wire [0:0] _zy_sva_brcm_key_type_43_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_key_type_43_cpass;
`_2_ wire _zy_sva_b42;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_44_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_44_cpass;
`_2_ wire _zy_sva_b43;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_iv_45_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_iv_45_cpass;
`_2_ wire _zy_sva_b44;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_46_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_46_cpass;
`_2_ wire _zy_sva_b45;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_iv_47_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_iv_47_cpass;
`_2_ wire _zy_sva_b46;
`_2_ wire [0:0] _zy_sva_brcm_key_type_48_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_key_type_48_cpass;
`_2_ wire _zy_sva_b47;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_49_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_49_cpass;
`_2_ wire _zy_sva_b48;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_iv_50_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_iv_50_cpass;
`_2_ wire _zy_sva_b49;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_51_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_51_cpass;
`_2_ wire _zy_sva_b50;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_iv_52_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_iv_52_cpass;
`_2_ wire _zy_sva_b51;
`_2_ wire [0:0] _zy_sva_brcm_key_type_53_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_key_type_53_cpass;
`_2_ wire _zy_sva_b52;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_54_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_54_cpass;
`_2_ wire _zy_sva_b53;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_iv_55_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_iv_55_cpass;
`_2_ wire _zy_sva_b54;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_56_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_56_cpass;
`_2_ wire _zy_sva_b55;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_iv_57_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_iv_57_cpass;
`_2_ wire _zy_sva_b56;
`_2_ wire [0:0] _zy_sva_brcm_key_type_58_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_key_type_58_cpass;
`_2_ wire _zy_sva_b57;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_59_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_59_cpass;
`_2_ wire _zy_sva_b58;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_iv_60_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_iv_60_cpass;
`_2_ wire _zy_sva_b59;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_61_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_61_cpass;
`_2_ wire _zy_sva_b60;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_iv_62_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_iv_62_cpass;
`_2_ wire _zy_sva_b61;
`_2_ wire [0:0] _zy_sva_brcm_key_type_63_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_key_type_63_cpass;
`_2_ wire _zy_sva_b62;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_64_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_64_cpass;
`_2_ wire _zy_sva_b63;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_iv_65_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_iv_65_cpass;
`_2_ wire _zy_sva_b64;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_66_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_66_cpass;
`_2_ wire _zy_sva_b65;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_iv_67_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_iv_67_cpass;
`_2_ wire _zy_sva_b66;
`_2_ wire [0:0] _zy_sva_brcm_key_type_68_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_key_type_68_cpass;
`_2_ wire _zy_sva_b67;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_69_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_69_cpass;
`_2_ wire _zy_sva_b68;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_iv_70_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_iv_70_cpass;
`_2_ wire _zy_sva_b69;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_71_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_71_cpass;
`_2_ wire _zy_sva_b70;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_iv_72_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_iv_72_cpass;
`_2_ wire _zy_sva_b71;
`_2_ wire [0:0] _zy_sva_brcm_key_type_73_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_key_type_73_cpass;
`_2_ wire _zy_sva_b72;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_74_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_74_cpass;
`_2_ wire _zy_sva_b73;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_iv_75_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_iv_75_cpass;
`_2_ wire _zy_sva_b74;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_76_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_76_cpass;
`_2_ wire _zy_sva_b75;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_iv_77_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_iv_77_cpass;
`_2_ wire _zy_sva_b76;
`_2_ wire [0:0] _zy_sva_brcm_key_type_78_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_key_type_78_cpass;
`_2_ wire _zy_sva_b77;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_79_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_79_cpass;
`_2_ wire _zy_sva_b78;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_iv_80_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_iv_80_cpass;
`_2_ wire _zy_sva_b79;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_81_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_81_cpass;
`_2_ wire _zy_sva_b80;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_iv_82_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_iv_82_cpass;
`_2_ wire _zy_sva_b81;
`_2_ wire [0:0] _zy_sva_brcm_key_type_83_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_key_type_83_cpass;
`_2_ wire _zy_sva_b82;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_84_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_84_cpass;
`_2_ wire _zy_sva_b83;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_iv_85_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_iv_85_cpass;
`_2_ wire _zy_sva_b84;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_86_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_86_cpass;
`_2_ wire _zy_sva_b85;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_iv_87_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_iv_87_cpass;
`_2_ wire _zy_sva_b86;
`_2_ wire [0:0] _zy_sva_brcm_key_type_88_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_key_type_88_cpass;
`_2_ wire _zy_sva_b87;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_89_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_89_cpass;
`_2_ wire _zy_sva_b88;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_iv_90_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_iv_90_cpass;
`_2_ wire _zy_sva_b89;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_91_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_91_cpass;
`_2_ wire _zy_sva_b90;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_iv_92_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_iv_92_cpass;
`_2_ wire _zy_sva_b91;
`_2_ wire [0:0] _zy_sva_brcm_key_type_93_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_key_type_93_cpass;
`_2_ wire _zy_sva_b92;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_94_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_94_cpass;
`_2_ wire _zy_sva_b93;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_iv_95_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_iv_95_cpass;
`_2_ wire _zy_sva_b94;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_96_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_96_cpass;
`_2_ wire _zy_sva_b95;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_iv_97_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_iv_97_cpass;
`_2_ wire _zy_sva_b96;
`_2_ wire [0:0] _zy_sva_brcm_key_type_98_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_key_type_98_cpass;
`_2_ wire _zy_sva_b97;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_99_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_99_cpass;
`_2_ wire _zy_sva_b98;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_iv_100_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_iv_100_cpass;
`_2_ wire _zy_sva_b99;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_101_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_101_cpass;
`_2_ wire _zy_sva_b100;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_iv_102_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_iv_102_cpass;
`_2_ wire _zy_sva_b101;
`_2_ wire [0:0] _zy_sva_brcm_key_type_103_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_key_type_103_cpass;
`_2_ wire _zy_sva_b102;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_104_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_104_cpass;
`_2_ wire _zy_sva_b103;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_iv_105_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_iv_105_cpass;
`_2_ wire _zy_sva_b104;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_106_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_106_cpass;
`_2_ wire _zy_sva_b105;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_iv_107_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_aux_cmd_guid_iv_107_cpass;
`_2_ wire _zy_sva_b106;
`_2_ wire [0:0] _zy_sva_brcm_key_type_108_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_key_type_108_cpass;
`_2_ wire _zy_sva_b107;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_109_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_109_cpass;
`_2_ wire _zy_sva_b108;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_110_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_110_cpass;
`_2_ wire _zy_sva_b109;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_111_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_111_cpass;
`_2_ wire _zy_sva_b110;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_112_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_112_cpass;
`_2_ wire _zy_sva_b111;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_113_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_113_cpass;
`_2_ wire _zy_sva_b112;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_114_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_114_cpass;
`_2_ wire _zy_sva_b113;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_115_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_115_cpass;
`_2_ wire _zy_sva_b114;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_116_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_116_cpass;
`_2_ wire _zy_sva_b115;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_117_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_117_cpass;
`_2_ wire _zy_sva_b116;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_118_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_118_cpass;
`_2_ wire _zy_sva_b117;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_119_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_119_cpass;
`_2_ wire _zy_sva_b118;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_120_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_120_cpass;
`_2_ wire _zy_sva_b119;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_121_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_121_cpass;
`_2_ wire _zy_sva_b120;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_122_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_122_cpass;
`_2_ wire _zy_sva_b121;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_123_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_123_cpass;
`_2_ wire _zy_sva_b122;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_124_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_ops_124_cpass;
`_2_ wire _zy_sva_b123;
`_2_ wire [0:0] _zy_sva_null_gcm_125_ccheck;
`_2_ wire [0:0] _zy_sva_null_gcm_125_cpass;
`_2_ wire _zy_sva_b124;
`_2_ wire [0:0] _zy_sva_sha_gcm_126_ccheck;
`_2_ wire [0:0] _zy_sva_sha_gcm_126_cpass;
`_2_ wire _zy_sva_b125;
`_2_ wire [0:0] _zy_sva_null_xts_127_ccheck;
`_2_ wire [0:0] _zy_sva_null_xts_127_cpass;
`_2_ wire _zy_sva_b126;
`_2_ wire [0:0] _zy_sva_sha_xts_128_ccheck;
`_2_ wire [0:0] _zy_sva_sha_xts_128_cpass;
`_2_ wire _zy_sva_b127;
`_2_ wire [0:0] _zy_sva_null_null_129_ccheck;
`_2_ wire [0:0] _zy_sva_null_null_129_cpass;
`_2_ wire _zy_sva_b128;
`_2_ wire [0:0] _zy_sva_sha_null_130_ccheck;
`_2_ wire [0:0] _zy_sva_sha_null_130_cpass;
`_2_ wire _zy_sva_b129;
`_2_ wire [0:0] _zy_sva_hmac_gcm_131_ccheck;
`_2_ wire [0:0] _zy_sva_hmac_gcm_131_cpass;
`_2_ wire _zy_sva_b130;
`_2_ wire [0:0] _zy_sva_hmac_xts_132_ccheck;
`_2_ wire [0:0] _zy_sva_hmac_xts_132_cpass;
`_2_ wire _zy_sva_b131;
`_2_ wire [0:0] _zy_sva_hmac_null_133_ccheck;
`_2_ wire [0:0] _zy_sva_hmac_null_133_cpass;
`_2_ wire _zy_sva_b132;
`_2_ wire [0:0] _zy_sva_null_gcm_134_ccheck;
`_2_ wire [0:0] _zy_sva_null_gcm_134_cpass;
`_2_ wire _zy_sva_b133;
`_2_ wire [0:0] _zy_sva_sha_gcm_135_ccheck;
`_2_ wire [0:0] _zy_sva_sha_gcm_135_cpass;
`_2_ wire _zy_sva_b134;
`_2_ wire [0:0] _zy_sva_null_xts_136_ccheck;
`_2_ wire [0:0] _zy_sva_null_xts_136_cpass;
`_2_ wire _zy_sva_b135;
`_2_ wire [0:0] _zy_sva_sha_xts_137_ccheck;
`_2_ wire [0:0] _zy_sva_sha_xts_137_cpass;
`_2_ wire _zy_sva_b136;
`_2_ wire [0:0] _zy_sva_null_null_138_ccheck;
`_2_ wire [0:0] _zy_sva_null_null_138_cpass;
`_2_ wire _zy_sva_b137;
`_2_ wire [0:0] _zy_sva_sha_null_139_ccheck;
`_2_ wire [0:0] _zy_sva_sha_null_139_cpass;
`_2_ wire _zy_sva_b138;
`_2_ wire [0:0] _zy_sva_hmac_gcm_140_ccheck;
`_2_ wire [0:0] _zy_sva_hmac_gcm_140_cpass;
`_2_ wire _zy_sva_b139;
`_2_ wire [0:0] _zy_sva_hmac_xts_141_ccheck;
`_2_ wire [0:0] _zy_sva_hmac_xts_141_cpass;
`_2_ wire _zy_sva_b140;
`_2_ wire [0:0] _zy_sva_hmac_null_142_ccheck;
`_2_ wire [0:0] _zy_sva_hmac_null_142_cpass;
`_2_ wire _zy_sva_b141;
`_2_ wire [0:0] _zy_sva_null_gcm_143_ccheck;
`_2_ wire [0:0] _zy_sva_null_gcm_143_cpass;
`_2_ wire _zy_sva_b142;
`_2_ wire [0:0] _zy_sva_sha_gcm_144_ccheck;
`_2_ wire [0:0] _zy_sva_sha_gcm_144_cpass;
`_2_ wire _zy_sva_b143;
`_2_ wire [0:0] _zy_sva_null_xts_145_ccheck;
`_2_ wire [0:0] _zy_sva_null_xts_145_cpass;
`_2_ wire _zy_sva_b144;
`_2_ wire [0:0] _zy_sva_sha_xts_146_ccheck;
`_2_ wire [0:0] _zy_sva_sha_xts_146_cpass;
`_2_ wire _zy_sva_b145;
`_2_ wire [0:0] _zy_sva_null_null_147_ccheck;
`_2_ wire [0:0] _zy_sva_null_null_147_cpass;
`_2_ wire _zy_sva_b146;
`_2_ wire [0:0] _zy_sva_sha_null_148_ccheck;
`_2_ wire [0:0] _zy_sva_sha_null_148_cpass;
`_2_ wire _zy_sva_b147;
`_2_ wire [0:0] _zy_sva_hmac_gcm_149_ccheck;
`_2_ wire [0:0] _zy_sva_hmac_gcm_149_cpass;
`_2_ wire _zy_sva_b148;
`_2_ wire [0:0] _zy_sva_hmac_xts_150_ccheck;
`_2_ wire [0:0] _zy_sva_hmac_xts_150_cpass;
`_2_ wire _zy_sva_b149;
`_2_ wire [0:0] _zy_sva_hmac_null_151_ccheck;
`_2_ wire [0:0] _zy_sva_hmac_null_151_cpass;
`_2_ wire _zy_sva_b150;
`_2_ wire [0:0] _zy_sva_null_gcm_152_ccheck;
`_2_ wire [0:0] _zy_sva_null_gcm_152_cpass;
`_2_ wire _zy_sva_b151;
`_2_ wire [0:0] _zy_sva_sha_gcm_153_ccheck;
`_2_ wire [0:0] _zy_sva_sha_gcm_153_cpass;
`_2_ wire _zy_sva_b152;
`_2_ wire [0:0] _zy_sva_null_xts_154_ccheck;
`_2_ wire [0:0] _zy_sva_null_xts_154_cpass;
`_2_ wire _zy_sva_b153;
`_2_ wire [0:0] _zy_sva_sha_xts_155_ccheck;
`_2_ wire [0:0] _zy_sva_sha_xts_155_cpass;
`_2_ wire _zy_sva_b154;
`_2_ wire [0:0] _zy_sva_null_null_156_ccheck;
`_2_ wire [0:0] _zy_sva_null_null_156_cpass;
`_2_ wire _zy_sva_b155;
`_2_ wire [0:0] _zy_sva_sha_null_157_ccheck;
`_2_ wire [0:0] _zy_sva_sha_null_157_cpass;
`_2_ wire _zy_sva_b156;
`_2_ wire [0:0] _zy_sva_hmac_gcm_158_ccheck;
`_2_ wire [0:0] _zy_sva_hmac_gcm_158_cpass;
`_2_ wire _zy_sva_b157;
`_2_ wire [0:0] _zy_sva_hmac_xts_159_ccheck;
`_2_ wire [0:0] _zy_sva_hmac_xts_159_cpass;
`_2_ wire _zy_sva_b158;
`_2_ wire [0:0] _zy_sva_hmac_null_160_ccheck;
`_2_ wire [0:0] _zy_sva_hmac_null_160_cpass;
`_2_ wire _zy_sva_b159;
`_2_ wire [0:0] _zy_sva_null_gcm_161_ccheck;
`_2_ wire [0:0] _zy_sva_null_gcm_161_cpass;
`_2_ wire _zy_sva_b160;
`_2_ wire [0:0] _zy_sva_sha_gcm_162_ccheck;
`_2_ wire [0:0] _zy_sva_sha_gcm_162_cpass;
`_2_ wire _zy_sva_b161;
`_2_ wire [0:0] _zy_sva_null_xts_163_ccheck;
`_2_ wire [0:0] _zy_sva_null_xts_163_cpass;
`_2_ wire _zy_sva_b162;
`_2_ wire [0:0] _zy_sva_sha_xts_164_ccheck;
`_2_ wire [0:0] _zy_sva_sha_xts_164_cpass;
`_2_ wire _zy_sva_b163;
`_2_ wire [0:0] _zy_sva_null_null_165_ccheck;
`_2_ wire [0:0] _zy_sva_null_null_165_cpass;
`_2_ wire _zy_sva_b164;
`_2_ wire [0:0] _zy_sva_sha_null_166_ccheck;
`_2_ wire [0:0] _zy_sva_sha_null_166_cpass;
`_2_ wire _zy_sva_b165;
`_2_ wire [0:0] _zy_sva_hmac_gcm_167_ccheck;
`_2_ wire [0:0] _zy_sva_hmac_gcm_167_cpass;
`_2_ wire _zy_sva_b166;
`_2_ wire [0:0] _zy_sva_hmac_xts_168_ccheck;
`_2_ wire [0:0] _zy_sva_hmac_xts_168_cpass;
`_2_ wire _zy_sva_b167;
`_2_ wire [0:0] _zy_sva_hmac_null_169_ccheck;
`_2_ wire [0:0] _zy_sva_hmac_null_169_cpass;
`_2_ wire _zy_sva_b168;
`_2_ wire [0:0] _zy_sva_null_gcm_170_ccheck;
`_2_ wire [0:0] _zy_sva_null_gcm_170_cpass;
`_2_ wire _zy_sva_b169;
`_2_ wire [0:0] _zy_sva_sha_gcm_171_ccheck;
`_2_ wire [0:0] _zy_sva_sha_gcm_171_cpass;
`_2_ wire _zy_sva_b170;
`_2_ wire [0:0] _zy_sva_null_xts_172_ccheck;
`_2_ wire [0:0] _zy_sva_null_xts_172_cpass;
`_2_ wire _zy_sva_b171;
`_2_ wire [0:0] _zy_sva_sha_xts_173_ccheck;
`_2_ wire [0:0] _zy_sva_sha_xts_173_cpass;
`_2_ wire _zy_sva_b172;
`_2_ wire [0:0] _zy_sva_null_null_174_ccheck;
`_2_ wire [0:0] _zy_sva_null_null_174_cpass;
`_2_ wire _zy_sva_b173;
`_2_ wire [0:0] _zy_sva_sha_null_175_ccheck;
`_2_ wire [0:0] _zy_sva_sha_null_175_cpass;
`_2_ wire _zy_sva_b174;
`_2_ wire [0:0] _zy_sva_hmac_gcm_176_ccheck;
`_2_ wire [0:0] _zy_sva_hmac_gcm_176_cpass;
`_2_ wire _zy_sva_b175;
`_2_ wire [0:0] _zy_sva_hmac_xts_177_ccheck;
`_2_ wire [0:0] _zy_sva_hmac_xts_177_cpass;
`_2_ wire _zy_sva_b176;
`_2_ wire [0:0] _zy_sva_hmac_null_178_ccheck;
`_2_ wire [0:0] _zy_sva_hmac_null_178_cpass;
`_2_ wire _zy_sva_b177;
wire [63:0] _zyL234_tfiRv52;
wire _zyL252_tfiRv53;
wire _zyL253_tfiRv54;
wire _zyL254_tfiRv55;
wire _zyL255_tfiRv56;
wire [63:0] _zyL288_tfiRv57;
wire [63:0] _zyL293_tfiRv58;
wire [63:0] _zyL301_tfiRv59;
wire [63:0] _zyL306_tfiRv60;
wire [63:0] _zyL313_tfiRv61;
wire [63:0] _zyL321_tfiRv62;
wire [63:0] _zyL327_tfiRv63;
wire [63:0] _zyL337_tfiRv64;
wire [63:0] _zyL346_tfiRv65;
wire [63:0] _zyL354_tfiRv66;
wire [63:0] _zyL359_tfiRv67;
wire [63:0] _zyL368_tfiRv68;
wire [63:0] _zyL373_tfiRv69;
wire [63:0] _zyL382_tfiRv70;
wire [63:0] _zyL390_tfiRv71;
wire [63:0] _zyL395_tfiRv72;
wire [63:0] _zyL410_tfiRv73;
wire _zyL485_tfiRv74;
wire _zyL486_tfiRv75;
wire _zyL489_tfiRv76;
wire _zyL489_tfiRv77;
wire _zyL492_tfiRv78;
wire [63:0] _zyL526_tfiRv79;
wire [63:0] _zyL527_tfiRv80;
wire [63:0] _zyL541_tfiRv81;
wire [63:0] _zyL542_tfiRv82;
wire [63:0] _zyL555_tfiRv83;
wire [63:0] _zyL556_tfiRv84;
wire [63:0] _zyL569_tfiRv85;
wire [63:0] _zyL570_tfiRv86;
supply1 n47;
supply0 n1735;
wire [0:0] \fifo_in.sot ;
wire [0:0] \fifo_in.eoi ;
wire [0:0] \fifo_in.eot ;
wire [3:0] \fifo_in.id ;
wire [63:0] \fifo_in.tdata ;
wire [1:0] \tlv_word0.tlv_bip2 ;
wire \tlv_word0.no_data ;
wire \tlv_word0.aux_frmd_crc ;
wire [3:0] \tlv_word0.frame_size ;
wire \tlv_word0.vf_valid ;
wire [0:0] \tlv_word0.trace ;
wire [10:0] \tlv_word0.unused ;
wire [10:0] \tlv_word0.tlv_frame_num ;
wire [3:0] \tlv_word0.resv0 ;
wire [3:0] \tlv_word0.tlv_eng_id ;
wire [7:0] \tlv_word0.tlv_seq_num ;
wire [7:0] \tlv_word0.tlv_len ;
wire [7:0] \tlv_word0.tlv_type ;
wire [3:0] \tlv_word1.pf_number ;
wire [11:0] \tlv_word1.vf_number ;
wire [15:0] \tlv_word1.scheduler_handle ;
wire [31:0] \tlv_word1.src_data_len ;
wire \tlv_word2.rsvd2 ;
wire [5:0] \tlv_word2.key_type ;
wire [1:0] \tlv_word2.rsvd1 ;
wire [0:0] \tlv_word2.cipher_pad ;
wire [1:0] \tlv_word2.iv_op ;
wire [7:0] \tlv_word2.aad_len ;
wire [3:0] \tlv_word2.cipher_op ;
wire [3:0] \tlv_word2.auth_op ;
wire [3:0] \tlv_word2.raw_auth_op ;
wire [7:0] \tlv_word2.rsvd0 ;
wire [1:0] \tlv_word2.chu_comp_thrsh ;
wire [0:0] \tlv_word2.xp10_crc_mode ;
wire [5:0] \tlv_word2.xp10_user_prefix_size ;
wire [1:0] \tlv_word2.xp10_prefix_mode ;
wire [1:0] \tlv_word2.lz77_max_symb_len ;
wire [0:0] \tlv_word2.lz77_min_match_len ;
wire [1:0] \tlv_word2.lz77_dly_match_win ;
wire [3:0] \tlv_word2.lz77_win_size ;
wire [3:0] \tlv_word2.comp_mode ;
wire [0:0] \frame_word.debug.tlvp_corrupt ;
wire [1:0] \frame_word.debug.cmd_mode ;
wire [4:0] \frame_word.debug.module_id ;
wire [0:0] \frame_word.debug.cmd_type ;
wire [4:0] \frame_word.debug.tlv_num ;
wire [9:0] \frame_word.debug.byte_num ;
wire [7:0] \frame_word.debug.byte_msk ;
wire \frame_word.trace ;
wire \frame_word.dst_guid_present ;
wire [6:0] \frame_word.frmd_out_type ;
wire [1:0] \frame_word.md_op ;
wire [1:0] \frame_word.md_type ;
wire [6:0] \frame_word.frmd_in_type ;
wire [5:0] \frame_word.frmd_in_aux ;
wire [0:0] \frame_word.frmd_crc_in ;
wire [0:0] \frame_word.src_guid_present ;
wire [3:0] \frame_word.compound_cmd_frm_size ;
wire [1:0] \kme_internal_word0.tlv_bip2 ;
wire [12:0] \kme_internal_word0.resv0 ;
wire [0:0] \kme_internal_word0.kdf_dek_iter ;
wire [0:0] \kme_internal_word0.keyless_algos ;
wire [0:0] \kme_internal_word0.needs_dek ;
wire [0:0] \kme_internal_word0.needs_dak ;
wire [5:0] \kme_internal_word0.key_type ;
wire [10:0] \kme_internal_word0.tlv_frame_num ;
wire [3:0] \kme_internal_word0.tlv_eng_id ;
wire [7:0] \kme_internal_word0.tlv_seq_num ;
wire [7:0] \kme_internal_word0.tlv_len ;
wire [7:0] \kme_internal_word0.tlv_type ;
wire [1:0] \nxt_kme_internal_word0.tlv_bip2 ;
wire [12:0] \nxt_kme_internal_word0.resv0 ;
wire [0:0] \nxt_kme_internal_word0.kdf_dek_iter ;
wire [0:0] \nxt_kme_internal_word0.keyless_algos ;
wire [0:0] \nxt_kme_internal_word0.needs_dek ;
wire [0:0] \nxt_kme_internal_word0.needs_dak ;
wire [5:0] \nxt_kme_internal_word0.key_type ;
wire [10:0] \nxt_kme_internal_word0.tlv_frame_num ;
wire [3:0] \nxt_kme_internal_word0.tlv_eng_id ;
wire [7:0] \nxt_kme_internal_word0.tlv_seq_num ;
wire [7:0] \nxt_kme_internal_word0.tlv_len ;
wire [7:0] \nxt_kme_internal_word0.tlv_type ;
wire [0:0] \kme_internal_dek_kim_word.dek_kim_entry.valid ;
wire [2:0] \kme_internal_dek_kim_word.dek_kim_entry.label_index ;
wire [1:0] \kme_internal_dek_kim_word.dek_kim_entry.ckv_length ;
wire [14:0] \kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer ;
wire [3:0] \kme_internal_dek_kim_word.dek_kim_entry.pf_num ;
wire [11:0] \kme_internal_dek_kim_word.dek_kim_entry.vf_num ;
wire [0:0] \kme_internal_dek_kim_word.dek_kim_entry.vf_valid ;
wire [5:0] \kme_internal_dek_kim_word.unused ;
wire [0:0] \kme_internal_dek_kim_word.missing_iv ;
wire [0:0] \kme_internal_dek_kim_word.missing_guid ;
wire [0:0] \kme_internal_dek_kim_word.validate_dek ;
wire [0:0] \kme_internal_dek_kim_word.vf_valid ;
wire [3:0] \kme_internal_dek_kim_word.pf_num ;
wire [11:0] \kme_internal_dek_kim_word.vf_num ;
wire [0:0] \nxt_kme_internal_dek_kim_word.dek_kim_entry.valid ;
wire [2:0] \nxt_kme_internal_dek_kim_word.dek_kim_entry.label_index ;
wire [1:0] \nxt_kme_internal_dek_kim_word.dek_kim_entry.ckv_length ;
wire [14:0] \nxt_kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer ;
wire [3:0] \nxt_kme_internal_dek_kim_word.dek_kim_entry.pf_num ;
wire [11:0] \nxt_kme_internal_dek_kim_word.dek_kim_entry.vf_num ;
wire [0:0] \nxt_kme_internal_dek_kim_word.dek_kim_entry.vf_valid ;
wire [5:0] \nxt_kme_internal_dek_kim_word.unused ;
wire [0:0] \nxt_kme_internal_dek_kim_word.missing_iv ;
wire [0:0] \nxt_kme_internal_dek_kim_word.missing_guid ;
wire [0:0] \nxt_kme_internal_dek_kim_word.validate_dek ;
wire [0:0] \nxt_kme_internal_dek_kim_word.vf_valid ;
wire [3:0] \nxt_kme_internal_dek_kim_word.pf_num ;
wire [11:0] \nxt_kme_internal_dek_kim_word.vf_num ;
wire [0:0] \kme_internal_dak_kim_word.dak_kim_entry.valid ;
wire [2:0] \kme_internal_dak_kim_word.dak_kim_entry.label_index ;
wire [1:0] \kme_internal_dak_kim_word.dak_kim_entry.ckv_length ;
wire [14:0] \kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer ;
wire [3:0] \kme_internal_dak_kim_word.dak_kim_entry.pf_num ;
wire [11:0] \kme_internal_dak_kim_word.dak_kim_entry.vf_num ;
wire [0:0] \kme_internal_dak_kim_word.dak_kim_entry.vf_valid ;
wire [7:0] \kme_internal_dak_kim_word.unused ;
wire [0:0] \kme_internal_dak_kim_word.validate_dak ;
wire [0:0] \kme_internal_dak_kim_word.vf_valid ;
wire [3:0] \kme_internal_dak_kim_word.pf_num ;
wire [11:0] \kme_internal_dak_kim_word.vf_num ;
wire [0:0] \nxt_kme_internal_dak_kim_word.dak_kim_entry.valid ;
wire [2:0] \nxt_kme_internal_dak_kim_word.dak_kim_entry.label_index ;
wire [1:0] \nxt_kme_internal_dak_kim_word.dak_kim_entry.ckv_length ;
wire [14:0] \nxt_kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer ;
wire [3:0] \nxt_kme_internal_dak_kim_word.dak_kim_entry.pf_num ;
wire [11:0] \nxt_kme_internal_dak_kim_word.dak_kim_entry.vf_num ;
wire [0:0] \nxt_kme_internal_dak_kim_word.dak_kim_entry.vf_valid ;
wire [7:0] \nxt_kme_internal_dak_kim_word.unused ;
wire [0:0] \nxt_kme_internal_dak_kim_word.validate_dak ;
wire [0:0] \nxt_kme_internal_dak_kim_word.vf_valid ;
wire [3:0] \nxt_kme_internal_dak_kim_word.pf_num ;
wire [11:0] \nxt_kme_internal_dak_kim_word.vf_num ;
wire [0:0] \debug_cmd.tlvp_corrupt ;
wire [1:0] \debug_cmd.cmd_mode ;
wire [4:0] \debug_cmd.module_id ;
wire [0:0] \debug_cmd.cmd_type ;
wire [4:0] \debug_cmd.tlv_num ;
wire [9:0] \debug_cmd.byte_num ;
wire [7:0] \debug_cmd.byte_msk ;
wire [0:0] \nxt_debug_cmd.tlvp_corrupt ;
wire [1:0] \nxt_debug_cmd.cmd_mode ;
wire [4:0] \nxt_debug_cmd.module_id ;
wire [0:0] \nxt_debug_cmd.cmd_type ;
wire [4:0] \nxt_debug_cmd.tlv_num ;
wire [9:0] \nxt_debug_cmd.byte_num ;
wire [7:0] \nxt_debug_cmd.byte_msk ;
wire [0:0] \aux_key_header.dak_key_op ;
wire [13:0] \aux_key_header.dak_key_ref ;
wire [1:0] \aux_key_header.kdf_mode ;
wire [0:0] \aux_key_header.dek_key_op ;
wire [13:0] \aux_key_header.dek_key_ref ;
wire [0:0] \nxt_aux_key_header.dak_key_op ;
wire [13:0] \nxt_aux_key_header.dak_key_ref ;
wire [1:0] \nxt_aux_key_header.kdf_mode ;
wire [0:0] \nxt_aux_key_header.dek_key_op ;
wire [13:0] \nxt_aux_key_header.dek_key_ref ;
wire [0:0] \skip.start ;
wire [0:0] \skip.partial ;
wire [0:0] \skip.endian_swap ;
wire [3:0] \skip.till ;
wire [0:0] \nxt_skip.start ;
wire [0:0] \nxt_skip.partial ;
wire [0:0] \nxt_skip.endian_swap ;
wire [3:0] \nxt_skip.till ;
tran (parser_kimreader_data[70], \parser_kimreader_data.sot [0]);
tran (parser_kimreader_data[69], \parser_kimreader_data.eoi [0]);
tran (parser_kimreader_data[68], \parser_kimreader_data.eot [0]);
tran (parser_kimreader_data[67], \parser_kimreader_data.id [3]);
tran (parser_kimreader_data[66], \parser_kimreader_data.id [2]);
tran (parser_kimreader_data[65], \parser_kimreader_data.id [1]);
tran (parser_kimreader_data[64], \parser_kimreader_data.id [0]);
tran (parser_kimreader_data[63], \parser_kimreader_data.tdata [63]);
tran (parser_kimreader_data[62], \parser_kimreader_data.tdata [62]);
tran (parser_kimreader_data[61], \parser_kimreader_data.tdata [61]);
tran (parser_kimreader_data[60], \parser_kimreader_data.tdata [60]);
tran (parser_kimreader_data[59], \parser_kimreader_data.tdata [59]);
tran (parser_kimreader_data[58], \parser_kimreader_data.tdata [58]);
tran (parser_kimreader_data[57], \parser_kimreader_data.tdata [57]);
tran (parser_kimreader_data[56], \parser_kimreader_data.tdata [56]);
tran (parser_kimreader_data[55], \parser_kimreader_data.tdata [55]);
tran (parser_kimreader_data[54], \parser_kimreader_data.tdata [54]);
tran (parser_kimreader_data[53], \parser_kimreader_data.tdata [53]);
tran (parser_kimreader_data[52], \parser_kimreader_data.tdata [52]);
tran (parser_kimreader_data[51], \parser_kimreader_data.tdata [51]);
tran (parser_kimreader_data[50], \parser_kimreader_data.tdata [50]);
tran (parser_kimreader_data[49], \parser_kimreader_data.tdata [49]);
tran (parser_kimreader_data[48], \parser_kimreader_data.tdata [48]);
tran (parser_kimreader_data[47], \parser_kimreader_data.tdata [47]);
tran (parser_kimreader_data[46], \parser_kimreader_data.tdata [46]);
tran (parser_kimreader_data[45], \parser_kimreader_data.tdata [45]);
tran (parser_kimreader_data[44], \parser_kimreader_data.tdata [44]);
tran (parser_kimreader_data[43], \parser_kimreader_data.tdata [43]);
tran (parser_kimreader_data[42], \parser_kimreader_data.tdata [42]);
tran (parser_kimreader_data[41], \parser_kimreader_data.tdata [41]);
tran (parser_kimreader_data[40], \parser_kimreader_data.tdata [40]);
tran (parser_kimreader_data[39], \parser_kimreader_data.tdata [39]);
tran (parser_kimreader_data[38], \parser_kimreader_data.tdata [38]);
tran (parser_kimreader_data[37], \parser_kimreader_data.tdata [37]);
tran (parser_kimreader_data[36], \parser_kimreader_data.tdata [36]);
tran (parser_kimreader_data[35], \parser_kimreader_data.tdata [35]);
tran (parser_kimreader_data[34], \parser_kimreader_data.tdata [34]);
tran (parser_kimreader_data[33], \parser_kimreader_data.tdata [33]);
tran (parser_kimreader_data[32], \parser_kimreader_data.tdata [32]);
tran (parser_kimreader_data[31], \parser_kimreader_data.tdata [31]);
tran (parser_kimreader_data[30], \parser_kimreader_data.tdata [30]);
tran (parser_kimreader_data[29], \parser_kimreader_data.tdata [29]);
tran (parser_kimreader_data[28], \parser_kimreader_data.tdata [28]);
tran (parser_kimreader_data[27], \parser_kimreader_data.tdata [27]);
tran (parser_kimreader_data[26], \parser_kimreader_data.tdata [26]);
tran (parser_kimreader_data[25], \parser_kimreader_data.tdata [25]);
tran (parser_kimreader_data[24], \parser_kimreader_data.tdata [24]);
tran (parser_kimreader_data[23], \parser_kimreader_data.tdata [23]);
tran (parser_kimreader_data[22], \parser_kimreader_data.tdata [22]);
tran (parser_kimreader_data[21], \parser_kimreader_data.tdata [21]);
tran (parser_kimreader_data[20], \parser_kimreader_data.tdata [20]);
tran (parser_kimreader_data[19], \parser_kimreader_data.tdata [19]);
tran (parser_kimreader_data[18], \parser_kimreader_data.tdata [18]);
tran (parser_kimreader_data[17], \parser_kimreader_data.tdata [17]);
tran (parser_kimreader_data[16], \parser_kimreader_data.tdata [16]);
tran (parser_kimreader_data[15], \parser_kimreader_data.tdata [15]);
tran (parser_kimreader_data[14], \parser_kimreader_data.tdata [14]);
tran (parser_kimreader_data[13], \parser_kimreader_data.tdata [13]);
tran (parser_kimreader_data[12], \parser_kimreader_data.tdata [12]);
tran (parser_kimreader_data[11], \parser_kimreader_data.tdata [11]);
tran (parser_kimreader_data[10], \parser_kimreader_data.tdata [10]);
tran (parser_kimreader_data[9], \parser_kimreader_data.tdata [9]);
tran (parser_kimreader_data[8], \parser_kimreader_data.tdata [8]);
tran (parser_kimreader_data[7], \parser_kimreader_data.tdata [7]);
tran (parser_kimreader_data[6], \parser_kimreader_data.tdata [6]);
tran (parser_kimreader_data[5], \parser_kimreader_data.tdata [5]);
tran (parser_kimreader_data[4], \parser_kimreader_data.tdata [4]);
tran (parser_kimreader_data[3], \parser_kimreader_data.tdata [3]);
tran (parser_kimreader_data[2], \parser_kimreader_data.tdata [2]);
tran (parser_kimreader_data[1], \parser_kimreader_data.tdata [1]);
tran (parser_kimreader_data[0], \parser_kimreader_data.tdata [0]);
tran (stitcher_out[82], \stitcher_out.tvalid );
tran (stitcher_out[81], \stitcher_out.tlast );
tran (stitcher_out[80], \stitcher_out.tid [0]);
tran (stitcher_out[79], \stitcher_out.tstrb [7]);
tran (stitcher_out[78], \stitcher_out.tstrb [6]);
tran (stitcher_out[77], \stitcher_out.tstrb [5]);
tran (stitcher_out[76], \stitcher_out.tstrb [4]);
tran (stitcher_out[75], \stitcher_out.tstrb [3]);
tran (stitcher_out[74], \stitcher_out.tstrb [2]);
tran (stitcher_out[73], \stitcher_out.tstrb [1]);
tran (stitcher_out[72], \stitcher_out.tstrb [0]);
tran (stitcher_out[71], \stitcher_out.tuser [7]);
tran (stitcher_out[70], \stitcher_out.tuser [6]);
tran (stitcher_out[69], \stitcher_out.tuser [5]);
tran (stitcher_out[68], \stitcher_out.tuser [4]);
tran (stitcher_out[67], \stitcher_out.tuser [3]);
tran (stitcher_out[66], \stitcher_out.tuser [2]);
tran (stitcher_out[65], \stitcher_out.tuser [1]);
tran (stitcher_out[64], \stitcher_out.tuser [0]);
tran (stitcher_out[63], \stitcher_out.tdata [63]);
tran (stitcher_out[62], \stitcher_out.tdata [62]);
tran (stitcher_out[61], \stitcher_out.tdata [61]);
tran (stitcher_out[60], \stitcher_out.tdata [60]);
tran (stitcher_out[59], \stitcher_out.tdata [59]);
tran (stitcher_out[58], \stitcher_out.tdata [58]);
tran (stitcher_out[57], \stitcher_out.tdata [57]);
tran (stitcher_out[56], \stitcher_out.tdata [56]);
tran (stitcher_out[55], \stitcher_out.tdata [55]);
tran (stitcher_out[54], \stitcher_out.tdata [54]);
tran (stitcher_out[53], \stitcher_out.tdata [53]);
tran (stitcher_out[52], \stitcher_out.tdata [52]);
tran (stitcher_out[51], \stitcher_out.tdata [51]);
tran (stitcher_out[50], \stitcher_out.tdata [50]);
tran (stitcher_out[49], \stitcher_out.tdata [49]);
tran (stitcher_out[48], \stitcher_out.tdata [48]);
tran (stitcher_out[47], \stitcher_out.tdata [47]);
tran (stitcher_out[46], \stitcher_out.tdata [46]);
tran (stitcher_out[45], \stitcher_out.tdata [45]);
tran (stitcher_out[44], \stitcher_out.tdata [44]);
tran (stitcher_out[43], \stitcher_out.tdata [43]);
tran (stitcher_out[42], \stitcher_out.tdata [42]);
tran (stitcher_out[41], \stitcher_out.tdata [41]);
tran (stitcher_out[40], \stitcher_out.tdata [40]);
tran (stitcher_out[39], \stitcher_out.tdata [39]);
tran (stitcher_out[38], \stitcher_out.tdata [38]);
tran (stitcher_out[37], \stitcher_out.tdata [37]);
tran (stitcher_out[36], \stitcher_out.tdata [36]);
tran (stitcher_out[35], \stitcher_out.tdata [35]);
tran (stitcher_out[34], \stitcher_out.tdata [34]);
tran (stitcher_out[33], \stitcher_out.tdata [33]);
tran (stitcher_out[32], \stitcher_out.tdata [32]);
tran (stitcher_out[31], \stitcher_out.tdata [31]);
tran (stitcher_out[30], \stitcher_out.tdata [30]);
tran (stitcher_out[29], \stitcher_out.tdata [29]);
tran (stitcher_out[28], \stitcher_out.tdata [28]);
tran (stitcher_out[27], \stitcher_out.tdata [27]);
tran (stitcher_out[26], \stitcher_out.tdata [26]);
tran (stitcher_out[25], \stitcher_out.tdata [25]);
tran (stitcher_out[24], \stitcher_out.tdata [24]);
tran (stitcher_out[23], \stitcher_out.tdata [23]);
tran (stitcher_out[22], \stitcher_out.tdata [22]);
tran (stitcher_out[21], \stitcher_out.tdata [21]);
tran (stitcher_out[20], \stitcher_out.tdata [20]);
tran (stitcher_out[19], \stitcher_out.tdata [19]);
tran (stitcher_out[18], \stitcher_out.tdata [18]);
tran (stitcher_out[17], \stitcher_out.tdata [17]);
tran (stitcher_out[16], \stitcher_out.tdata [16]);
tran (stitcher_out[15], \stitcher_out.tdata [15]);
tran (stitcher_out[14], \stitcher_out.tdata [14]);
tran (stitcher_out[13], \stitcher_out.tdata [13]);
tran (stitcher_out[12], \stitcher_out.tdata [12]);
tran (stitcher_out[11], \stitcher_out.tdata [11]);
tran (stitcher_out[10], \stitcher_out.tdata [10]);
tran (stitcher_out[9], \stitcher_out.tdata [9]);
tran (stitcher_out[8], \stitcher_out.tdata [8]);
tran (stitcher_out[7], \stitcher_out.tdata [7]);
tran (stitcher_out[6], \stitcher_out.tdata [6]);
tran (stitcher_out[5], \stitcher_out.tdata [5]);
tran (stitcher_out[4], \stitcher_out.tdata [4]);
tran (stitcher_out[3], \stitcher_out.tdata [3]);
tran (stitcher_out[2], \stitcher_out.tdata [2]);
tran (stitcher_out[1], \stitcher_out.tdata [1]);
tran (stitcher_out[0], \stitcher_out.tdata [0]);
tran (tlv_word0[63], \tlv_word0.tlv_bip2 [1]);
tran (tlv_word1[63], \tlv_word1.pf_number [3]);
tran (tlv_word2[63], \tlv_word2.rsvd2 );
tran (frame_word[63], \frame_word.debug.tlvp_corrupt [0]);
tran (tlv_word0[62], \tlv_word0.tlv_bip2 [0]);
tran (tlv_word1[62], \tlv_word1.pf_number [2]);
tran (tlv_word2[62], \tlv_word2.key_type [5]);
tran (frame_word[62], \frame_word.debug.cmd_mode [1]);
tran (tlv_word0[61], \tlv_word0.no_data );
tran (tlv_word1[61], \tlv_word1.pf_number [1]);
tran (tlv_word2[61], \tlv_word2.key_type [4]);
tran (frame_word[61], \frame_word.debug.cmd_mode [0]);
tran (tlv_word0[60], \tlv_word0.aux_frmd_crc );
tran (tlv_word1[60], \tlv_word1.pf_number [0]);
tran (tlv_word2[60], \tlv_word2.key_type [3]);
tran (frame_word[60], \frame_word.debug.module_id [4]);
tran (tlv_word0[59], \tlv_word0.frame_size [3]);
tran (tlv_word1[59], \tlv_word1.vf_number [11]);
tran (tlv_word2[59], \tlv_word2.key_type [2]);
tran (frame_word[59], \frame_word.debug.module_id [3]);
tran (tlv_word0[58], \tlv_word0.frame_size [2]);
tran (tlv_word1[58], \tlv_word1.vf_number [10]);
tran (tlv_word2[58], \tlv_word2.key_type [1]);
tran (frame_word[58], \frame_word.debug.module_id [2]);
tran (tlv_word0[57], \tlv_word0.frame_size [1]);
tran (tlv_word1[57], \tlv_word1.vf_number [9]);
tran (tlv_word2[57], \tlv_word2.key_type [0]);
tran (frame_word[57], \frame_word.debug.module_id [1]);
tran (tlv_word0[56], \tlv_word0.frame_size [0]);
tran (tlv_word1[56], \tlv_word1.vf_number [8]);
tran (tlv_word2[56], \tlv_word2.rsvd1 [1]);
tran (frame_word[56], \frame_word.debug.module_id [0]);
tran (tlv_word0[55], \tlv_word0.vf_valid );
tran (tlv_word1[55], \tlv_word1.vf_number [7]);
tran (tlv_word2[55], \tlv_word2.rsvd1 [0]);
tran (frame_word[55], \frame_word.debug.cmd_type [0]);
tran (tlv_word0[54], \tlv_word0.trace [0]);
tran (tlv_word1[54], \tlv_word1.vf_number [6]);
tran (tlv_word2[54], \tlv_word2.cipher_pad [0]);
tran (frame_word[54], \frame_word.debug.tlv_num [4]);
tran (tlv_word0[53], \tlv_word0.unused [10]);
tran (tlv_word1[53], \tlv_word1.vf_number [5]);
tran (tlv_word2[53], \tlv_word2.iv_op [1]);
tran (frame_word[53], \frame_word.debug.tlv_num [3]);
tran (tlv_word0[52], \tlv_word0.unused [9]);
tran (tlv_word1[52], \tlv_word1.vf_number [4]);
tran (tlv_word2[52], \tlv_word2.iv_op [0]);
tran (frame_word[52], \frame_word.debug.tlv_num [2]);
tran (tlv_word0[51], \tlv_word0.unused [8]);
tran (tlv_word1[51], \tlv_word1.vf_number [3]);
tran (tlv_word2[51], \tlv_word2.aad_len [7]);
tran (frame_word[51], \frame_word.debug.tlv_num [1]);
tran (tlv_word0[50], \tlv_word0.unused [7]);
tran (tlv_word1[50], \tlv_word1.vf_number [2]);
tran (tlv_word2[50], \tlv_word2.aad_len [6]);
tran (frame_word[50], \frame_word.debug.tlv_num [0]);
tran (tlv_word0[49], \tlv_word0.unused [6]);
tran (tlv_word1[49], \tlv_word1.vf_number [1]);
tran (tlv_word2[49], \tlv_word2.aad_len [5]);
tran (frame_word[49], \frame_word.debug.byte_num [9]);
tran (tlv_word0[48], \tlv_word0.unused [5]);
tran (tlv_word1[48], \tlv_word1.vf_number [0]);
tran (tlv_word2[48], \tlv_word2.aad_len [4]);
tran (frame_word[48], \frame_word.debug.byte_num [8]);
tran (tlv_word0[47], \tlv_word0.unused [4]);
tran (tlv_word1[47], \tlv_word1.scheduler_handle [15]);
tran (tlv_word2[47], \tlv_word2.aad_len [3]);
tran (frame_word[47], \frame_word.debug.byte_num [7]);
tran (tlv_word0[46], \tlv_word0.unused [3]);
tran (tlv_word1[46], \tlv_word1.scheduler_handle [14]);
tran (tlv_word2[46], \tlv_word2.aad_len [2]);
tran (frame_word[46], \frame_word.debug.byte_num [6]);
tran (tlv_word0[45], \tlv_word0.unused [2]);
tran (tlv_word1[45], \tlv_word1.scheduler_handle [13]);
tran (tlv_word2[45], \tlv_word2.aad_len [1]);
tran (frame_word[45], \frame_word.debug.byte_num [5]);
tran (tlv_word0[44], \tlv_word0.unused [1]);
tran (tlv_word1[44], \tlv_word1.scheduler_handle [12]);
tran (tlv_word2[44], \tlv_word2.aad_len [0]);
tran (frame_word[44], \frame_word.debug.byte_num [4]);
tran (tlv_word0[43], \tlv_word0.unused [0]);
tran (tlv_word1[43], \tlv_word1.scheduler_handle [11]);
tran (tlv_word2[43], \tlv_word2.cipher_op [3]);
tran (frame_word[43], \frame_word.debug.byte_num [3]);
tran (tlv_word0[42], \tlv_word0.tlv_frame_num [10]);
tran (tlv_word1[42], \tlv_word1.scheduler_handle [10]);
tran (tlv_word2[42], \tlv_word2.cipher_op [2]);
tran (frame_word[42], \frame_word.debug.byte_num [2]);
tran (tlv_word0[41], \tlv_word0.tlv_frame_num [9]);
tran (tlv_word1[41], \tlv_word1.scheduler_handle [9]);
tran (tlv_word2[41], \tlv_word2.cipher_op [1]);
tran (frame_word[41], \frame_word.debug.byte_num [1]);
tran (tlv_word0[40], \tlv_word0.tlv_frame_num [8]);
tran (tlv_word1[40], \tlv_word1.scheduler_handle [8]);
tran (tlv_word2[40], \tlv_word2.cipher_op [0]);
tran (frame_word[40], \frame_word.debug.byte_num [0]);
tran (tlv_word0[39], \tlv_word0.tlv_frame_num [7]);
tran (tlv_word1[39], \tlv_word1.scheduler_handle [7]);
tran (tlv_word2[39], \tlv_word2.auth_op [3]);
tran (frame_word[39], \frame_word.debug.byte_msk [7]);
tran (tlv_word0[38], \tlv_word0.tlv_frame_num [6]);
tran (tlv_word1[38], \tlv_word1.scheduler_handle [6]);
tran (tlv_word2[38], \tlv_word2.auth_op [2]);
tran (frame_word[38], \frame_word.debug.byte_msk [6]);
tran (tlv_word0[37], \tlv_word0.tlv_frame_num [5]);
tran (tlv_word1[37], \tlv_word1.scheduler_handle [5]);
tran (tlv_word2[37], \tlv_word2.auth_op [1]);
tran (frame_word[37], \frame_word.debug.byte_msk [5]);
tran (tlv_word0[36], \tlv_word0.tlv_frame_num [4]);
tran (tlv_word1[36], \tlv_word1.scheduler_handle [4]);
tran (tlv_word2[36], \tlv_word2.auth_op [0]);
tran (frame_word[36], \frame_word.debug.byte_msk [4]);
tran (tlv_word0[35], \tlv_word0.tlv_frame_num [3]);
tran (tlv_word1[35], \tlv_word1.scheduler_handle [3]);
tran (tlv_word2[35], \tlv_word2.raw_auth_op [3]);
tran (frame_word[35], \frame_word.debug.byte_msk [3]);
tran (tlv_word0[34], \tlv_word0.tlv_frame_num [2]);
tran (tlv_word1[34], \tlv_word1.scheduler_handle [2]);
tran (tlv_word2[34], \tlv_word2.raw_auth_op [2]);
tran (frame_word[34], \frame_word.debug.byte_msk [2]);
tran (tlv_word0[33], \tlv_word0.tlv_frame_num [1]);
tran (tlv_word1[33], \tlv_word1.scheduler_handle [1]);
tran (tlv_word2[33], \tlv_word2.raw_auth_op [1]);
tran (frame_word[33], \frame_word.debug.byte_msk [1]);
tran (tlv_word0[32], \tlv_word0.tlv_frame_num [0]);
tran (tlv_word1[32], \tlv_word1.scheduler_handle [0]);
tran (tlv_word2[32], \tlv_word2.raw_auth_op [0]);
tran (frame_word[32], \frame_word.debug.byte_msk [0]);
tran (tlv_word0[31], \tlv_word0.resv0 [3]);
tran (tlv_word1[31], \tlv_word1.src_data_len [31]);
tran (tlv_word2[31], \tlv_word2.rsvd0 [7]);
tran (frame_word[31], \frame_word.trace );
tran (tlv_word0[30], \tlv_word0.resv0 [2]);
tran (tlv_word1[30], \tlv_word1.src_data_len [30]);
tran (tlv_word2[30], \tlv_word2.rsvd0 [6]);
tran (frame_word[30], \frame_word.dst_guid_present );
tran (tlv_word0[29], \tlv_word0.resv0 [1]);
tran (tlv_word1[29], \tlv_word1.src_data_len [29]);
tran (tlv_word2[29], \tlv_word2.rsvd0 [5]);
tran (frame_word[29], \frame_word.frmd_out_type [6]);
tran (tlv_word0[28], \tlv_word0.resv0 [0]);
tran (tlv_word1[28], \tlv_word1.src_data_len [28]);
tran (tlv_word2[28], \tlv_word2.rsvd0 [4]);
tran (frame_word[28], \frame_word.frmd_out_type [5]);
tran (tlv_word0[27], \tlv_word0.tlv_eng_id [3]);
tran (tlv_word1[27], \tlv_word1.src_data_len [27]);
tran (tlv_word2[27], \tlv_word2.rsvd0 [3]);
tran (frame_word[27], \frame_word.frmd_out_type [4]);
tran (tlv_word0[26], \tlv_word0.tlv_eng_id [2]);
tran (tlv_word1[26], \tlv_word1.src_data_len [26]);
tran (tlv_word2[26], \tlv_word2.rsvd0 [2]);
tran (frame_word[26], \frame_word.frmd_out_type [3]);
tran (tlv_word0[25], \tlv_word0.tlv_eng_id [1]);
tran (tlv_word1[25], \tlv_word1.src_data_len [25]);
tran (tlv_word2[25], \tlv_word2.rsvd0 [1]);
tran (frame_word[25], \frame_word.frmd_out_type [2]);
tran (tlv_word0[24], \tlv_word0.tlv_eng_id [0]);
tran (tlv_word1[24], \tlv_word1.src_data_len [24]);
tran (tlv_word2[24], \tlv_word2.rsvd0 [0]);
tran (frame_word[24], \frame_word.frmd_out_type [1]);
tran (tlv_word0[23], \tlv_word0.tlv_seq_num [7]);
tran (tlv_word1[23], \tlv_word1.src_data_len [23]);
tran (tlv_word2[23], \tlv_word2.chu_comp_thrsh [1]);
tran (frame_word[23], \frame_word.frmd_out_type [0]);
tran (tlv_word0[22], \tlv_word0.tlv_seq_num [6]);
tran (tlv_word1[22], \tlv_word1.src_data_len [22]);
tran (tlv_word2[22], \tlv_word2.chu_comp_thrsh [0]);
tran (frame_word[22], \frame_word.md_op [1]);
tran (tlv_word0[21], \tlv_word0.tlv_seq_num [5]);
tran (tlv_word1[21], \tlv_word1.src_data_len [21]);
tran (tlv_word2[21], \tlv_word2.xp10_crc_mode [0]);
tran (frame_word[21], \frame_word.md_op [0]);
tran (tlv_word0[20], \tlv_word0.tlv_seq_num [4]);
tran (tlv_word1[20], \tlv_word1.src_data_len [20]);
tran (tlv_word2[20], \tlv_word2.xp10_user_prefix_size [5]);
tran (frame_word[20], \frame_word.md_type [1]);
tran (tlv_word0[19], \tlv_word0.tlv_seq_num [3]);
tran (tlv_word1[19], \tlv_word1.src_data_len [19]);
tran (tlv_word2[19], \tlv_word2.xp10_user_prefix_size [4]);
tran (frame_word[19], \frame_word.md_type [0]);
tran (tlv_word0[18], \tlv_word0.tlv_seq_num [2]);
tran (tlv_word1[18], \tlv_word1.src_data_len [18]);
tran (tlv_word2[18], \tlv_word2.xp10_user_prefix_size [3]);
tran (frame_word[18], \frame_word.frmd_in_type [6]);
tran (tlv_word0[17], \tlv_word0.tlv_seq_num [1]);
tran (tlv_word1[17], \tlv_word1.src_data_len [17]);
tran (tlv_word2[17], \tlv_word2.xp10_user_prefix_size [2]);
tran (frame_word[17], \frame_word.frmd_in_type [5]);
tran (tlv_word0[16], \tlv_word0.tlv_seq_num [0]);
tran (tlv_word1[16], \tlv_word1.src_data_len [16]);
tran (tlv_word2[16], \tlv_word2.xp10_user_prefix_size [1]);
tran (frame_word[16], \frame_word.frmd_in_type [4]);
tran (tlv_word0[15], \tlv_word0.tlv_len [7]);
tran (tlv_word1[15], \tlv_word1.src_data_len [15]);
tran (tlv_word2[15], \tlv_word2.xp10_user_prefix_size [0]);
tran (frame_word[15], \frame_word.frmd_in_type [3]);
tran (tlv_word0[14], \tlv_word0.tlv_len [6]);
tran (tlv_word1[14], \tlv_word1.src_data_len [14]);
tran (tlv_word2[14], \tlv_word2.xp10_prefix_mode [1]);
tran (frame_word[14], \frame_word.frmd_in_type [2]);
tran (tlv_word0[13], \tlv_word0.tlv_len [5]);
tran (tlv_word1[13], \tlv_word1.src_data_len [13]);
tran (tlv_word2[13], \tlv_word2.xp10_prefix_mode [0]);
tran (frame_word[13], \frame_word.frmd_in_type [1]);
tran (tlv_word0[12], \tlv_word0.tlv_len [4]);
tran (tlv_word1[12], \tlv_word1.src_data_len [12]);
tran (tlv_word2[12], \tlv_word2.lz77_max_symb_len [1]);
tran (frame_word[12], \frame_word.frmd_in_type [0]);
tran (tlv_word0[11], \tlv_word0.tlv_len [3]);
tran (tlv_word1[11], \tlv_word1.src_data_len [11]);
tran (tlv_word2[11], \tlv_word2.lz77_max_symb_len [0]);
tran (frame_word[11], \frame_word.frmd_in_aux [5]);
tran (tlv_word0[10], \tlv_word0.tlv_len [2]);
tran (tlv_word1[10], \tlv_word1.src_data_len [10]);
tran (tlv_word2[10], \tlv_word2.lz77_min_match_len [0]);
tran (frame_word[10], \frame_word.frmd_in_aux [4]);
tran (tlv_word0[9], \tlv_word0.tlv_len [1]);
tran (tlv_word1[9], \tlv_word1.src_data_len [9]);
tran (tlv_word2[9], \tlv_word2.lz77_dly_match_win [1]);
tran (frame_word[9], \frame_word.frmd_in_aux [3]);
tran (tlv_word0[8], \tlv_word0.tlv_len [0]);
tran (tlv_word1[8], \tlv_word1.src_data_len [8]);
tran (tlv_word2[8], \tlv_word2.lz77_dly_match_win [0]);
tran (frame_word[8], \frame_word.frmd_in_aux [2]);
tran (tlv_word0[7], \tlv_word0.tlv_type [7]);
tran (tlv_word1[7], \tlv_word1.src_data_len [7]);
tran (tlv_word2[7], \tlv_word2.lz77_win_size [3]);
tran (frame_word[7], \frame_word.frmd_in_aux [1]);
tran (tlv_word0[6], \tlv_word0.tlv_type [6]);
tran (tlv_word1[6], \tlv_word1.src_data_len [6]);
tran (tlv_word2[6], \tlv_word2.lz77_win_size [2]);
tran (frame_word[6], \frame_word.frmd_in_aux [0]);
tran (tlv_word0[5], \tlv_word0.tlv_type [5]);
tran (tlv_word1[5], \tlv_word1.src_data_len [5]);
tran (tlv_word2[5], \tlv_word2.lz77_win_size [1]);
tran (frame_word[5], \frame_word.frmd_crc_in [0]);
tran (tlv_word0[4], \tlv_word0.tlv_type [4]);
tran (tlv_word1[4], \tlv_word1.src_data_len [4]);
tran (tlv_word2[4], \tlv_word2.lz77_win_size [0]);
tran (frame_word[4], \frame_word.src_guid_present [0]);
tran (tlv_word0[3], \tlv_word0.tlv_type [3]);
tran (tlv_word1[3], \tlv_word1.src_data_len [3]);
tran (tlv_word2[3], \tlv_word2.comp_mode [3]);
tran (frame_word[3], \frame_word.compound_cmd_frm_size [3]);
tran (tlv_word0[2], \tlv_word0.tlv_type [2]);
tran (tlv_word1[2], \tlv_word1.src_data_len [2]);
tran (tlv_word2[2], \tlv_word2.comp_mode [2]);
tran (frame_word[2], \frame_word.compound_cmd_frm_size [2]);
tran (tlv_word0[1], \tlv_word0.tlv_type [1]);
tran (tlv_word1[1], \tlv_word1.src_data_len [1]);
tran (tlv_word2[1], \tlv_word2.comp_mode [1]);
tran (frame_word[1], \frame_word.compound_cmd_frm_size [1]);
tran (tlv_word0[0], \tlv_word0.tlv_type [0]);
tran (tlv_word1[0], \tlv_word1.src_data_len [0]);
tran (tlv_word2[0], \tlv_word2.comp_mode [0]);
tran (frame_word[0], \frame_word.compound_cmd_frm_size [0]);
tran (skip[4], \skip.endian_swap [0]);
tran (fifo_in[69], \fifo_in.eoi [0]);
tran (fifo_in[70], \fifo_in.sot [0]);
tran (fifo_in[68], \fifo_in.eot [0]);
tran (nxt_skip[0], \nxt_skip.till [0]);
tran (nxt_skip[1], \nxt_skip.till [1]);
tran (nxt_skip[2], \nxt_skip.till [2]);
tran (nxt_skip[3], \nxt_skip.till [3]);
tran (nxt_skip[4], \nxt_skip.endian_swap [0]);
tran (nxt_skip[5], \nxt_skip.partial [0]);
tran (nxt_skip[6], \nxt_skip.start [0]);
tran (nxt_aux_key_header[0], \nxt_aux_key_header.dek_key_ref [0]);
tran (nxt_aux_key_header[1], \nxt_aux_key_header.dek_key_ref [1]);
tran (nxt_aux_key_header[2], \nxt_aux_key_header.dek_key_ref [2]);
tran (nxt_aux_key_header[3], \nxt_aux_key_header.dek_key_ref [3]);
tran (nxt_aux_key_header[4], \nxt_aux_key_header.dek_key_ref [4]);
tran (nxt_aux_key_header[5], \nxt_aux_key_header.dek_key_ref [5]);
tran (nxt_aux_key_header[6], \nxt_aux_key_header.dek_key_ref [6]);
tran (nxt_aux_key_header[7], \nxt_aux_key_header.dek_key_ref [7]);
tran (nxt_aux_key_header[8], \nxt_aux_key_header.dek_key_ref [8]);
tran (nxt_aux_key_header[9], \nxt_aux_key_header.dek_key_ref [9]);
tran (nxt_aux_key_header[10], \nxt_aux_key_header.dek_key_ref [10]);
tran (nxt_aux_key_header[11], \nxt_aux_key_header.dek_key_ref [11]);
tran (nxt_aux_key_header[12], \nxt_aux_key_header.dek_key_ref [12]);
tran (nxt_aux_key_header[13], \nxt_aux_key_header.dek_key_ref [13]);
tran (nxt_aux_key_header[14], \nxt_aux_key_header.dek_key_op [0]);
tran (nxt_aux_key_header[15], \nxt_aux_key_header.kdf_mode [0]);
tran (nxt_aux_key_header[16], \nxt_aux_key_header.kdf_mode [1]);
tran (nxt_aux_key_header[17], \nxt_aux_key_header.dak_key_ref [0]);
tran (nxt_aux_key_header[18], \nxt_aux_key_header.dak_key_ref [1]);
tran (nxt_aux_key_header[19], \nxt_aux_key_header.dak_key_ref [2]);
tran (nxt_aux_key_header[20], \nxt_aux_key_header.dak_key_ref [3]);
tran (nxt_aux_key_header[21], \nxt_aux_key_header.dak_key_ref [4]);
tran (nxt_aux_key_header[22], \nxt_aux_key_header.dak_key_ref [5]);
tran (nxt_aux_key_header[23], \nxt_aux_key_header.dak_key_ref [6]);
tran (nxt_aux_key_header[24], \nxt_aux_key_header.dak_key_ref [7]);
tran (nxt_aux_key_header[25], \nxt_aux_key_header.dak_key_ref [8]);
tran (nxt_aux_key_header[26], \nxt_aux_key_header.dak_key_ref [9]);
tran (nxt_aux_key_header[27], \nxt_aux_key_header.dak_key_ref [10]);
tran (nxt_aux_key_header[28], \nxt_aux_key_header.dak_key_ref [11]);
tran (nxt_aux_key_header[29], \nxt_aux_key_header.dak_key_ref [12]);
tran (nxt_aux_key_header[30], \nxt_aux_key_header.dak_key_ref [13]);
tran (nxt_aux_key_header[31], \nxt_aux_key_header.dak_key_op [0]);
tran (nxt_debug_cmd[0], \nxt_debug_cmd.byte_msk [0]);
tran (nxt_debug_cmd[1], \nxt_debug_cmd.byte_msk [1]);
tran (nxt_debug_cmd[2], \nxt_debug_cmd.byte_msk [2]);
tran (nxt_debug_cmd[3], \nxt_debug_cmd.byte_msk [3]);
tran (nxt_debug_cmd[4], \nxt_debug_cmd.byte_msk [4]);
tran (nxt_debug_cmd[5], \nxt_debug_cmd.byte_msk [5]);
tran (nxt_debug_cmd[6], \nxt_debug_cmd.byte_msk [6]);
tran (nxt_debug_cmd[7], \nxt_debug_cmd.byte_msk [7]);
tran (nxt_debug_cmd[8], \nxt_debug_cmd.byte_num [0]);
tran (nxt_debug_cmd[9], \nxt_debug_cmd.byte_num [1]);
tran (nxt_debug_cmd[10], \nxt_debug_cmd.byte_num [2]);
tran (nxt_debug_cmd[11], \nxt_debug_cmd.byte_num [3]);
tran (nxt_debug_cmd[12], \nxt_debug_cmd.byte_num [4]);
tran (nxt_debug_cmd[13], \nxt_debug_cmd.byte_num [5]);
tran (nxt_debug_cmd[14], \nxt_debug_cmd.byte_num [6]);
tran (nxt_debug_cmd[15], \nxt_debug_cmd.byte_num [7]);
tran (nxt_debug_cmd[16], \nxt_debug_cmd.byte_num [8]);
tran (nxt_debug_cmd[17], \nxt_debug_cmd.byte_num [9]);
tran (nxt_debug_cmd[18], \nxt_debug_cmd.tlv_num [0]);
tran (nxt_debug_cmd[19], \nxt_debug_cmd.tlv_num [1]);
tran (nxt_debug_cmd[20], \nxt_debug_cmd.tlv_num [2]);
tran (nxt_debug_cmd[21], \nxt_debug_cmd.tlv_num [3]);
tran (nxt_debug_cmd[22], \nxt_debug_cmd.tlv_num [4]);
tran (nxt_debug_cmd[23], \nxt_debug_cmd.cmd_type [0]);
tran (nxt_debug_cmd[24], \nxt_debug_cmd.module_id [0]);
tran (nxt_debug_cmd[25], \nxt_debug_cmd.module_id [1]);
tran (nxt_debug_cmd[26], \nxt_debug_cmd.module_id [2]);
tran (nxt_debug_cmd[27], \nxt_debug_cmd.module_id [3]);
tran (nxt_debug_cmd[28], \nxt_debug_cmd.module_id [4]);
tran (nxt_debug_cmd[29], \nxt_debug_cmd.cmd_mode [0]);
tran (nxt_debug_cmd[30], \nxt_debug_cmd.cmd_mode [1]);
tran (nxt_debug_cmd[31], \nxt_debug_cmd.tlvp_corrupt [0]);
tran (nxt_kme_internal_dak_kim_word[0], \nxt_kme_internal_dak_kim_word.vf_num [0]);
tran (nxt_kme_internal_dak_kim_word[1], \nxt_kme_internal_dak_kim_word.vf_num [1]);
tran (nxt_kme_internal_dak_kim_word[2], \nxt_kme_internal_dak_kim_word.vf_num [2]);
tran (nxt_kme_internal_dak_kim_word[3], \nxt_kme_internal_dak_kim_word.vf_num [3]);
tran (nxt_kme_internal_dak_kim_word[4], \nxt_kme_internal_dak_kim_word.vf_num [4]);
tran (nxt_kme_internal_dak_kim_word[5], \nxt_kme_internal_dak_kim_word.vf_num [5]);
tran (nxt_kme_internal_dak_kim_word[6], \nxt_kme_internal_dak_kim_word.vf_num [6]);
tran (nxt_kme_internal_dak_kim_word[7], \nxt_kme_internal_dak_kim_word.vf_num [7]);
tran (nxt_kme_internal_dak_kim_word[8], \nxt_kme_internal_dak_kim_word.vf_num [8]);
tran (nxt_kme_internal_dak_kim_word[9], \nxt_kme_internal_dak_kim_word.vf_num [9]);
tran (nxt_kme_internal_dak_kim_word[10], \nxt_kme_internal_dak_kim_word.vf_num [10]);
tran (nxt_kme_internal_dak_kim_word[11], \nxt_kme_internal_dak_kim_word.vf_num [11]);
tran (nxt_kme_internal_dak_kim_word[12], \nxt_kme_internal_dak_kim_word.pf_num [0]);
tran (nxt_kme_internal_dak_kim_word[13], \nxt_kme_internal_dak_kim_word.pf_num [1]);
tran (nxt_kme_internal_dak_kim_word[14], \nxt_kme_internal_dak_kim_word.pf_num [2]);
tran (nxt_kme_internal_dak_kim_word[15], \nxt_kme_internal_dak_kim_word.pf_num [3]);
tran (nxt_kme_internal_dak_kim_word[16], \nxt_kme_internal_dak_kim_word.vf_valid [0]);
tran (nxt_kme_internal_dak_kim_word[17], \nxt_kme_internal_dak_kim_word.validate_dak [0]);
tran (nxt_kme_internal_dak_kim_word[18], \nxt_kme_internal_dak_kim_word.unused [0]);
tran (nxt_kme_internal_dak_kim_word[19], \nxt_kme_internal_dak_kim_word.unused [1]);
tran (nxt_kme_internal_dak_kim_word[20], \nxt_kme_internal_dak_kim_word.unused [2]);
tran (nxt_kme_internal_dak_kim_word[21], \nxt_kme_internal_dak_kim_word.unused [3]);
tran (nxt_kme_internal_dak_kim_word[22], \nxt_kme_internal_dak_kim_word.unused [4]);
tran (nxt_kme_internal_dak_kim_word[23], \nxt_kme_internal_dak_kim_word.unused [5]);
tran (nxt_kme_internal_dak_kim_word[24], \nxt_kme_internal_dak_kim_word.unused [6]);
tran (nxt_kme_internal_dak_kim_word[25], \nxt_kme_internal_dak_kim_word.unused [7]);
tran (nxt_kme_internal_dak_kim_word[26], \nxt_kme_internal_dak_kim_word.dak_kim_entry.vf_valid [0]);
tran (nxt_kme_internal_dak_kim_word[27], \nxt_kme_internal_dak_kim_word.dak_kim_entry.vf_num [0]);
tran (nxt_kme_internal_dak_kim_word[28], \nxt_kme_internal_dak_kim_word.dak_kim_entry.vf_num [1]);
tran (nxt_kme_internal_dak_kim_word[29], \nxt_kme_internal_dak_kim_word.dak_kim_entry.vf_num [2]);
tran (nxt_kme_internal_dak_kim_word[30], \nxt_kme_internal_dak_kim_word.dak_kim_entry.vf_num [3]);
tran (nxt_kme_internal_dak_kim_word[31], \nxt_kme_internal_dak_kim_word.dak_kim_entry.vf_num [4]);
tran (nxt_kme_internal_dak_kim_word[32], \nxt_kme_internal_dak_kim_word.dak_kim_entry.vf_num [5]);
tran (nxt_kme_internal_dak_kim_word[33], \nxt_kme_internal_dak_kim_word.dak_kim_entry.vf_num [6]);
tran (nxt_kme_internal_dak_kim_word[34], \nxt_kme_internal_dak_kim_word.dak_kim_entry.vf_num [7]);
tran (nxt_kme_internal_dak_kim_word[35], \nxt_kme_internal_dak_kim_word.dak_kim_entry.vf_num [8]);
tran (nxt_kme_internal_dak_kim_word[36], \nxt_kme_internal_dak_kim_word.dak_kim_entry.vf_num [9]);
tran (nxt_kme_internal_dak_kim_word[37], \nxt_kme_internal_dak_kim_word.dak_kim_entry.vf_num [10]);
tran (nxt_kme_internal_dak_kim_word[38], \nxt_kme_internal_dak_kim_word.dak_kim_entry.vf_num [11]);
tran (nxt_kme_internal_dak_kim_word[39], \nxt_kme_internal_dak_kim_word.dak_kim_entry.pf_num [0]);
tran (nxt_kme_internal_dak_kim_word[40], \nxt_kme_internal_dak_kim_word.dak_kim_entry.pf_num [1]);
tran (nxt_kme_internal_dak_kim_word[41], \nxt_kme_internal_dak_kim_word.dak_kim_entry.pf_num [2]);
tran (nxt_kme_internal_dak_kim_word[42], \nxt_kme_internal_dak_kim_word.dak_kim_entry.pf_num [3]);
tran (nxt_kme_internal_dak_kim_word[43], \nxt_kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [0]);
tran (nxt_kme_internal_dak_kim_word[44], \nxt_kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [1]);
tran (nxt_kme_internal_dak_kim_word[45], \nxt_kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [2]);
tran (nxt_kme_internal_dak_kim_word[46], \nxt_kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [3]);
tran (nxt_kme_internal_dak_kim_word[47], \nxt_kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [4]);
tran (nxt_kme_internal_dak_kim_word[48], \nxt_kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [5]);
tran (nxt_kme_internal_dak_kim_word[49], \nxt_kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [6]);
tran (nxt_kme_internal_dak_kim_word[50], \nxt_kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [7]);
tran (nxt_kme_internal_dak_kim_word[51], \nxt_kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [8]);
tran (nxt_kme_internal_dak_kim_word[52], \nxt_kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [9]);
tran (nxt_kme_internal_dak_kim_word[53], \nxt_kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [10]);
tran (nxt_kme_internal_dak_kim_word[54], \nxt_kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [11]);
tran (nxt_kme_internal_dak_kim_word[55], \nxt_kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [12]);
tran (nxt_kme_internal_dak_kim_word[56], \nxt_kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [13]);
tran (nxt_kme_internal_dak_kim_word[57], \nxt_kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [14]);
tran (nxt_kme_internal_dak_kim_word[58], \nxt_kme_internal_dak_kim_word.dak_kim_entry.ckv_length [0]);
tran (nxt_kme_internal_dak_kim_word[59], \nxt_kme_internal_dak_kim_word.dak_kim_entry.ckv_length [1]);
tran (nxt_kme_internal_dak_kim_word[60], \nxt_kme_internal_dak_kim_word.dak_kim_entry.label_index [0]);
tran (nxt_kme_internal_dak_kim_word[61], \nxt_kme_internal_dak_kim_word.dak_kim_entry.label_index [1]);
tran (nxt_kme_internal_dak_kim_word[62], \nxt_kme_internal_dak_kim_word.dak_kim_entry.label_index [2]);
tran (nxt_kme_internal_dak_kim_word[63], \nxt_kme_internal_dak_kim_word.dak_kim_entry.valid [0]);
tran (nxt_kme_internal_dek_kim_word[0], \nxt_kme_internal_dek_kim_word.vf_num [0]);
tran (nxt_kme_internal_dek_kim_word[1], \nxt_kme_internal_dek_kim_word.vf_num [1]);
tran (nxt_kme_internal_dek_kim_word[2], \nxt_kme_internal_dek_kim_word.vf_num [2]);
tran (nxt_kme_internal_dek_kim_word[3], \nxt_kme_internal_dek_kim_word.vf_num [3]);
tran (nxt_kme_internal_dek_kim_word[4], \nxt_kme_internal_dek_kim_word.vf_num [4]);
tran (nxt_kme_internal_dek_kim_word[5], \nxt_kme_internal_dek_kim_word.vf_num [5]);
tran (nxt_kme_internal_dek_kim_word[6], \nxt_kme_internal_dek_kim_word.vf_num [6]);
tran (nxt_kme_internal_dek_kim_word[7], \nxt_kme_internal_dek_kim_word.vf_num [7]);
tran (nxt_kme_internal_dek_kim_word[8], \nxt_kme_internal_dek_kim_word.vf_num [8]);
tran (nxt_kme_internal_dek_kim_word[9], \nxt_kme_internal_dek_kim_word.vf_num [9]);
tran (nxt_kme_internal_dek_kim_word[10], \nxt_kme_internal_dek_kim_word.vf_num [10]);
tran (nxt_kme_internal_dek_kim_word[11], \nxt_kme_internal_dek_kim_word.vf_num [11]);
tran (nxt_kme_internal_dek_kim_word[12], \nxt_kme_internal_dek_kim_word.pf_num [0]);
tran (nxt_kme_internal_dek_kim_word[13], \nxt_kme_internal_dek_kim_word.pf_num [1]);
tran (nxt_kme_internal_dek_kim_word[14], \nxt_kme_internal_dek_kim_word.pf_num [2]);
tran (nxt_kme_internal_dek_kim_word[15], \nxt_kme_internal_dek_kim_word.pf_num [3]);
tran (nxt_kme_internal_dek_kim_word[16], \nxt_kme_internal_dek_kim_word.vf_valid [0]);
tran (nxt_kme_internal_dek_kim_word[17], \nxt_kme_internal_dek_kim_word.validate_dek [0]);
tran (nxt_kme_internal_dek_kim_word[18], \nxt_kme_internal_dek_kim_word.missing_guid [0]);
tran (nxt_kme_internal_dek_kim_word[19], \nxt_kme_internal_dek_kim_word.missing_iv [0]);
tran (nxt_kme_internal_dek_kim_word[20], \nxt_kme_internal_dek_kim_word.unused [0]);
tran (nxt_kme_internal_dek_kim_word[21], \nxt_kme_internal_dek_kim_word.unused [1]);
tran (nxt_kme_internal_dek_kim_word[22], \nxt_kme_internal_dek_kim_word.unused [2]);
tran (nxt_kme_internal_dek_kim_word[23], \nxt_kme_internal_dek_kim_word.unused [3]);
tran (nxt_kme_internal_dek_kim_word[24], \nxt_kme_internal_dek_kim_word.unused [4]);
tran (nxt_kme_internal_dek_kim_word[25], \nxt_kme_internal_dek_kim_word.unused [5]);
tran (nxt_kme_internal_dek_kim_word[26], \nxt_kme_internal_dek_kim_word.dek_kim_entry.vf_valid [0]);
tran (nxt_kme_internal_dek_kim_word[27], \nxt_kme_internal_dek_kim_word.dek_kim_entry.vf_num [0]);
tran (nxt_kme_internal_dek_kim_word[28], \nxt_kme_internal_dek_kim_word.dek_kim_entry.vf_num [1]);
tran (nxt_kme_internal_dek_kim_word[29], \nxt_kme_internal_dek_kim_word.dek_kim_entry.vf_num [2]);
tran (nxt_kme_internal_dek_kim_word[30], \nxt_kme_internal_dek_kim_word.dek_kim_entry.vf_num [3]);
tran (nxt_kme_internal_dek_kim_word[31], \nxt_kme_internal_dek_kim_word.dek_kim_entry.vf_num [4]);
tran (nxt_kme_internal_dek_kim_word[32], \nxt_kme_internal_dek_kim_word.dek_kim_entry.vf_num [5]);
tran (nxt_kme_internal_dek_kim_word[33], \nxt_kme_internal_dek_kim_word.dek_kim_entry.vf_num [6]);
tran (nxt_kme_internal_dek_kim_word[34], \nxt_kme_internal_dek_kim_word.dek_kim_entry.vf_num [7]);
tran (nxt_kme_internal_dek_kim_word[35], \nxt_kme_internal_dek_kim_word.dek_kim_entry.vf_num [8]);
tran (nxt_kme_internal_dek_kim_word[36], \nxt_kme_internal_dek_kim_word.dek_kim_entry.vf_num [9]);
tran (nxt_kme_internal_dek_kim_word[37], \nxt_kme_internal_dek_kim_word.dek_kim_entry.vf_num [10]);
tran (nxt_kme_internal_dek_kim_word[38], \nxt_kme_internal_dek_kim_word.dek_kim_entry.vf_num [11]);
tran (nxt_kme_internal_dek_kim_word[39], \nxt_kme_internal_dek_kim_word.dek_kim_entry.pf_num [0]);
tran (nxt_kme_internal_dek_kim_word[40], \nxt_kme_internal_dek_kim_word.dek_kim_entry.pf_num [1]);
tran (nxt_kme_internal_dek_kim_word[41], \nxt_kme_internal_dek_kim_word.dek_kim_entry.pf_num [2]);
tran (nxt_kme_internal_dek_kim_word[42], \nxt_kme_internal_dek_kim_word.dek_kim_entry.pf_num [3]);
tran (nxt_kme_internal_dek_kim_word[43], \nxt_kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [0]);
tran (nxt_kme_internal_dek_kim_word[44], \nxt_kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [1]);
tran (nxt_kme_internal_dek_kim_word[45], \nxt_kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [2]);
tran (nxt_kme_internal_dek_kim_word[46], \nxt_kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [3]);
tran (nxt_kme_internal_dek_kim_word[47], \nxt_kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [4]);
tran (nxt_kme_internal_dek_kim_word[48], \nxt_kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [5]);
tran (nxt_kme_internal_dek_kim_word[49], \nxt_kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [6]);
tran (nxt_kme_internal_dek_kim_word[50], \nxt_kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [7]);
tran (nxt_kme_internal_dek_kim_word[51], \nxt_kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [8]);
tran (nxt_kme_internal_dek_kim_word[52], \nxt_kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [9]);
tran (nxt_kme_internal_dek_kim_word[53], \nxt_kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [10]);
tran (nxt_kme_internal_dek_kim_word[54], \nxt_kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [11]);
tran (nxt_kme_internal_dek_kim_word[55], \nxt_kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [12]);
tran (nxt_kme_internal_dek_kim_word[56], \nxt_kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [13]);
tran (nxt_kme_internal_dek_kim_word[57], \nxt_kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [14]);
tran (nxt_kme_internal_dek_kim_word[58], \nxt_kme_internal_dek_kim_word.dek_kim_entry.ckv_length [0]);
tran (nxt_kme_internal_dek_kim_word[59], \nxt_kme_internal_dek_kim_word.dek_kim_entry.ckv_length [1]);
tran (nxt_kme_internal_dek_kim_word[60], \nxt_kme_internal_dek_kim_word.dek_kim_entry.label_index [0]);
tran (nxt_kme_internal_dek_kim_word[61], \nxt_kme_internal_dek_kim_word.dek_kim_entry.label_index [1]);
tran (nxt_kme_internal_dek_kim_word[62], \nxt_kme_internal_dek_kim_word.dek_kim_entry.label_index [2]);
tran (nxt_kme_internal_dek_kim_word[63], \nxt_kme_internal_dek_kim_word.dek_kim_entry.valid [0]);
tran (nxt_kme_internal_word0[0], \nxt_kme_internal_word0.tlv_type [0]);
tran (nxt_kme_internal_word0[1], \nxt_kme_internal_word0.tlv_type [1]);
tran (nxt_kme_internal_word0[2], \nxt_kme_internal_word0.tlv_type [2]);
tran (nxt_kme_internal_word0[3], \nxt_kme_internal_word0.tlv_type [3]);
tran (nxt_kme_internal_word0[4], \nxt_kme_internal_word0.tlv_type [4]);
tran (nxt_kme_internal_word0[5], \nxt_kme_internal_word0.tlv_type [5]);
tran (nxt_kme_internal_word0[6], \nxt_kme_internal_word0.tlv_type [6]);
tran (nxt_kme_internal_word0[7], \nxt_kme_internal_word0.tlv_type [7]);
tran (nxt_kme_internal_word0[8], \nxt_kme_internal_word0.tlv_len [0]);
tran (nxt_kme_internal_word0[9], \nxt_kme_internal_word0.tlv_len [1]);
tran (nxt_kme_internal_word0[10], \nxt_kme_internal_word0.tlv_len [2]);
tran (nxt_kme_internal_word0[11], \nxt_kme_internal_word0.tlv_len [3]);
tran (nxt_kme_internal_word0[12], \nxt_kme_internal_word0.tlv_len [4]);
tran (nxt_kme_internal_word0[13], \nxt_kme_internal_word0.tlv_len [5]);
tran (nxt_kme_internal_word0[14], \nxt_kme_internal_word0.tlv_len [6]);
tran (nxt_kme_internal_word0[15], \nxt_kme_internal_word0.tlv_len [7]);
tran (nxt_kme_internal_word0[16], \nxt_kme_internal_word0.tlv_seq_num [0]);
tran (nxt_kme_internal_word0[17], \nxt_kme_internal_word0.tlv_seq_num [1]);
tran (nxt_kme_internal_word0[18], \nxt_kme_internal_word0.tlv_seq_num [2]);
tran (nxt_kme_internal_word0[19], \nxt_kme_internal_word0.tlv_seq_num [3]);
tran (nxt_kme_internal_word0[20], \nxt_kme_internal_word0.tlv_seq_num [4]);
tran (nxt_kme_internal_word0[21], \nxt_kme_internal_word0.tlv_seq_num [5]);
tran (nxt_kme_internal_word0[22], \nxt_kme_internal_word0.tlv_seq_num [6]);
tran (nxt_kme_internal_word0[23], \nxt_kme_internal_word0.tlv_seq_num [7]);
tran (nxt_kme_internal_word0[24], \nxt_kme_internal_word0.tlv_eng_id [0]);
tran (nxt_kme_internal_word0[25], \nxt_kme_internal_word0.tlv_eng_id [1]);
tran (nxt_kme_internal_word0[26], \nxt_kme_internal_word0.tlv_eng_id [2]);
tran (nxt_kme_internal_word0[27], \nxt_kme_internal_word0.tlv_eng_id [3]);
tran (nxt_kme_internal_word0[28], \nxt_kme_internal_word0.tlv_frame_num [0]);
tran (nxt_kme_internal_word0[29], \nxt_kme_internal_word0.tlv_frame_num [1]);
tran (nxt_kme_internal_word0[30], \nxt_kme_internal_word0.tlv_frame_num [2]);
tran (nxt_kme_internal_word0[31], \nxt_kme_internal_word0.tlv_frame_num [3]);
tran (nxt_kme_internal_word0[32], \nxt_kme_internal_word0.tlv_frame_num [4]);
tran (nxt_kme_internal_word0[33], \nxt_kme_internal_word0.tlv_frame_num [5]);
tran (nxt_kme_internal_word0[34], \nxt_kme_internal_word0.tlv_frame_num [6]);
tran (nxt_kme_internal_word0[35], \nxt_kme_internal_word0.tlv_frame_num [7]);
tran (nxt_kme_internal_word0[36], \nxt_kme_internal_word0.tlv_frame_num [8]);
tran (nxt_kme_internal_word0[37], \nxt_kme_internal_word0.tlv_frame_num [9]);
tran (nxt_kme_internal_word0[38], \nxt_kme_internal_word0.tlv_frame_num [10]);
tran (nxt_kme_internal_word0[39], \nxt_kme_internal_word0.key_type [0]);
tran (nxt_kme_internal_word0[40], \nxt_kme_internal_word0.key_type [1]);
tran (nxt_kme_internal_word0[41], \nxt_kme_internal_word0.key_type [2]);
tran (nxt_kme_internal_word0[42], \nxt_kme_internal_word0.key_type [3]);
tran (nxt_kme_internal_word0[43], \nxt_kme_internal_word0.key_type [4]);
tran (nxt_kme_internal_word0[44], \nxt_kme_internal_word0.key_type [5]);
tran (nxt_kme_internal_word0[45], \nxt_kme_internal_word0.needs_dak [0]);
tran (nxt_kme_internal_word0[46], \nxt_kme_internal_word0.needs_dek [0]);
tran (nxt_kme_internal_word0[47], \nxt_kme_internal_word0.keyless_algos [0]);
tran (nxt_kme_internal_word0[48], \nxt_kme_internal_word0.kdf_dek_iter [0]);
tran (nxt_kme_internal_word0[49], \nxt_kme_internal_word0.resv0 [0]);
tran (nxt_kme_internal_word0[50], \nxt_kme_internal_word0.resv0 [1]);
tran (nxt_kme_internal_word0[51], \nxt_kme_internal_word0.resv0 [2]);
tran (nxt_kme_internal_word0[52], \nxt_kme_internal_word0.resv0 [3]);
tran (nxt_kme_internal_word0[53], \nxt_kme_internal_word0.resv0 [4]);
tran (nxt_kme_internal_word0[54], \nxt_kme_internal_word0.resv0 [5]);
tran (nxt_kme_internal_word0[55], \nxt_kme_internal_word0.resv0 [6]);
tran (nxt_kme_internal_word0[56], \nxt_kme_internal_word0.resv0 [7]);
tran (nxt_kme_internal_word0[57], \nxt_kme_internal_word0.resv0 [8]);
tran (nxt_kme_internal_word0[58], \nxt_kme_internal_word0.resv0 [9]);
tran (nxt_kme_internal_word0[59], \nxt_kme_internal_word0.resv0 [10]);
tran (nxt_kme_internal_word0[60], \nxt_kme_internal_word0.resv0 [11]);
tran (nxt_kme_internal_word0[61], \nxt_kme_internal_word0.resv0 [12]);
tran (nxt_kme_internal_word0[62], \nxt_kme_internal_word0.tlv_bip2 [0]);
tran (nxt_kme_internal_word0[63], \nxt_kme_internal_word0.tlv_bip2 [1]);
tran (fifo_in[0], \fifo_in.tdata [0]);
tran (fifo_in[1], \fifo_in.tdata [1]);
tran (fifo_in[2], \fifo_in.tdata [2]);
tran (fifo_in[3], \fifo_in.tdata [3]);
tran (fifo_in[4], \fifo_in.tdata [4]);
tran (fifo_in[5], \fifo_in.tdata [5]);
tran (fifo_in[6], \fifo_in.tdata [6]);
tran (fifo_in[7], \fifo_in.tdata [7]);
tran (fifo_in[8], \fifo_in.tdata [8]);
tran (fifo_in[9], \fifo_in.tdata [9]);
tran (fifo_in[10], \fifo_in.tdata [10]);
tran (fifo_in[11], \fifo_in.tdata [11]);
tran (fifo_in[12], \fifo_in.tdata [12]);
tran (fifo_in[13], \fifo_in.tdata [13]);
tran (fifo_in[14], \fifo_in.tdata [14]);
tran (fifo_in[15], \fifo_in.tdata [15]);
tran (fifo_in[16], \fifo_in.tdata [16]);
tran (fifo_in[17], \fifo_in.tdata [17]);
tran (fifo_in[18], \fifo_in.tdata [18]);
tran (fifo_in[19], \fifo_in.tdata [19]);
tran (fifo_in[20], \fifo_in.tdata [20]);
tran (fifo_in[21], \fifo_in.tdata [21]);
tran (fifo_in[22], \fifo_in.tdata [22]);
tran (fifo_in[23], \fifo_in.tdata [23]);
tran (fifo_in[24], \fifo_in.tdata [24]);
tran (fifo_in[25], \fifo_in.tdata [25]);
tran (fifo_in[26], \fifo_in.tdata [26]);
tran (fifo_in[27], \fifo_in.tdata [27]);
tran (fifo_in[28], \fifo_in.tdata [28]);
tran (fifo_in[29], \fifo_in.tdata [29]);
tran (fifo_in[30], \fifo_in.tdata [30]);
tran (fifo_in[31], \fifo_in.tdata [31]);
tran (fifo_in[32], \fifo_in.tdata [32]);
tran (fifo_in[33], \fifo_in.tdata [33]);
tran (fifo_in[34], \fifo_in.tdata [34]);
tran (fifo_in[35], \fifo_in.tdata [35]);
tran (fifo_in[36], \fifo_in.tdata [36]);
tran (fifo_in[37], \fifo_in.tdata [37]);
tran (fifo_in[38], \fifo_in.tdata [38]);
tran (fifo_in[39], \fifo_in.tdata [39]);
tran (fifo_in[40], \fifo_in.tdata [40]);
tran (fifo_in[41], \fifo_in.tdata [41]);
tran (fifo_in[42], \fifo_in.tdata [42]);
tran (fifo_in[43], \fifo_in.tdata [43]);
tran (fifo_in[44], \fifo_in.tdata [44]);
tran (fifo_in[45], \fifo_in.tdata [45]);
tran (fifo_in[46], \fifo_in.tdata [46]);
tran (fifo_in[47], \fifo_in.tdata [47]);
tran (fifo_in[48], \fifo_in.tdata [48]);
tran (fifo_in[49], \fifo_in.tdata [49]);
tran (fifo_in[50], \fifo_in.tdata [50]);
tran (fifo_in[51], \fifo_in.tdata [51]);
tran (fifo_in[52], \fifo_in.tdata [52]);
tran (fifo_in[53], \fifo_in.tdata [53]);
tran (fifo_in[54], \fifo_in.tdata [54]);
tran (fifo_in[55], \fifo_in.tdata [55]);
tran (fifo_in[56], \fifo_in.tdata [56]);
tran (fifo_in[57], \fifo_in.tdata [57]);
tran (fifo_in[58], \fifo_in.tdata [58]);
tran (fifo_in[59], \fifo_in.tdata [59]);
tran (fifo_in[60], \fifo_in.tdata [60]);
tran (fifo_in[61], \fifo_in.tdata [61]);
tran (fifo_in[62], \fifo_in.tdata [62]);
tran (fifo_in[63], \fifo_in.tdata [63]);
tran (skip[0], \skip.till [0]);
tran (skip[1], \skip.till [1]);
tran (skip[2], \skip.till [2]);
tran (skip[3], \skip.till [3]);
tran (skip[5], \skip.partial [0]);
tran (skip[6], \skip.start [0]);
tran (aux_key_header[0], \aux_key_header.dek_key_ref [0]);
tran (aux_key_header[1], \aux_key_header.dek_key_ref [1]);
tran (aux_key_header[2], \aux_key_header.dek_key_ref [2]);
tran (aux_key_header[3], \aux_key_header.dek_key_ref [3]);
tran (aux_key_header[4], \aux_key_header.dek_key_ref [4]);
tran (aux_key_header[5], \aux_key_header.dek_key_ref [5]);
tran (aux_key_header[6], \aux_key_header.dek_key_ref [6]);
tran (aux_key_header[7], \aux_key_header.dek_key_ref [7]);
tran (aux_key_header[8], \aux_key_header.dek_key_ref [8]);
tran (aux_key_header[9], \aux_key_header.dek_key_ref [9]);
tran (aux_key_header[10], \aux_key_header.dek_key_ref [10]);
tran (aux_key_header[11], \aux_key_header.dek_key_ref [11]);
tran (aux_key_header[12], \aux_key_header.dek_key_ref [12]);
tran (aux_key_header[13], \aux_key_header.dek_key_ref [13]);
tran (aux_key_header[14], \aux_key_header.dek_key_op [0]);
tran (aux_key_header[15], \aux_key_header.kdf_mode [0]);
tran (aux_key_header[16], \aux_key_header.kdf_mode [1]);
tran (aux_key_header[17], \aux_key_header.dak_key_ref [0]);
tran (aux_key_header[18], \aux_key_header.dak_key_ref [1]);
tran (aux_key_header[19], \aux_key_header.dak_key_ref [2]);
tran (aux_key_header[20], \aux_key_header.dak_key_ref [3]);
tran (aux_key_header[21], \aux_key_header.dak_key_ref [4]);
tran (aux_key_header[22], \aux_key_header.dak_key_ref [5]);
tran (aux_key_header[23], \aux_key_header.dak_key_ref [6]);
tran (aux_key_header[24], \aux_key_header.dak_key_ref [7]);
tran (aux_key_header[25], \aux_key_header.dak_key_ref [8]);
tran (aux_key_header[26], \aux_key_header.dak_key_ref [9]);
tran (aux_key_header[27], \aux_key_header.dak_key_ref [10]);
tran (aux_key_header[28], \aux_key_header.dak_key_ref [11]);
tran (aux_key_header[29], \aux_key_header.dak_key_ref [12]);
tran (aux_key_header[30], \aux_key_header.dak_key_ref [13]);
tran (aux_key_header[31], \aux_key_header.dak_key_op [0]);
tran (debug_cmd[0], \debug_cmd.byte_msk [0]);
tran (debug_cmd[1], \debug_cmd.byte_msk [1]);
tran (debug_cmd[2], \debug_cmd.byte_msk [2]);
tran (debug_cmd[3], \debug_cmd.byte_msk [3]);
tran (debug_cmd[4], \debug_cmd.byte_msk [4]);
tran (debug_cmd[5], \debug_cmd.byte_msk [5]);
tran (debug_cmd[6], \debug_cmd.byte_msk [6]);
tran (debug_cmd[7], \debug_cmd.byte_msk [7]);
tran (debug_cmd[8], \debug_cmd.byte_num [0]);
tran (debug_cmd[9], \debug_cmd.byte_num [1]);
tran (debug_cmd[10], \debug_cmd.byte_num [2]);
tran (debug_cmd[11], \debug_cmd.byte_num [3]);
tran (debug_cmd[12], \debug_cmd.byte_num [4]);
tran (debug_cmd[13], \debug_cmd.byte_num [5]);
tran (debug_cmd[14], \debug_cmd.byte_num [6]);
tran (debug_cmd[15], \debug_cmd.byte_num [7]);
tran (debug_cmd[16], \debug_cmd.byte_num [8]);
tran (debug_cmd[17], \debug_cmd.byte_num [9]);
tran (debug_cmd[18], \debug_cmd.tlv_num [0]);
tran (debug_cmd[19], \debug_cmd.tlv_num [1]);
tran (debug_cmd[20], \debug_cmd.tlv_num [2]);
tran (debug_cmd[21], \debug_cmd.tlv_num [3]);
tran (debug_cmd[22], \debug_cmd.tlv_num [4]);
tran (debug_cmd[23], \debug_cmd.cmd_type [0]);
tran (debug_cmd[24], \debug_cmd.module_id [0]);
tran (debug_cmd[25], \debug_cmd.module_id [1]);
tran (debug_cmd[26], \debug_cmd.module_id [2]);
tran (debug_cmd[27], \debug_cmd.module_id [3]);
tran (debug_cmd[28], \debug_cmd.module_id [4]);
tran (debug_cmd[29], \debug_cmd.cmd_mode [0]);
tran (debug_cmd[30], \debug_cmd.cmd_mode [1]);
tran (debug_cmd[31], \debug_cmd.tlvp_corrupt [0]);
tran (kme_internal_dak_kim_word[0], \kme_internal_dak_kim_word.vf_num [0]);
tran (kme_internal_dak_kim_word[1], \kme_internal_dak_kim_word.vf_num [1]);
tran (kme_internal_dak_kim_word[2], \kme_internal_dak_kim_word.vf_num [2]);
tran (kme_internal_dak_kim_word[3], \kme_internal_dak_kim_word.vf_num [3]);
tran (kme_internal_dak_kim_word[4], \kme_internal_dak_kim_word.vf_num [4]);
tran (kme_internal_dak_kim_word[5], \kme_internal_dak_kim_word.vf_num [5]);
tran (kme_internal_dak_kim_word[6], \kme_internal_dak_kim_word.vf_num [6]);
tran (kme_internal_dak_kim_word[7], \kme_internal_dak_kim_word.vf_num [7]);
tran (kme_internal_dak_kim_word[8], \kme_internal_dak_kim_word.vf_num [8]);
tran (kme_internal_dak_kim_word[9], \kme_internal_dak_kim_word.vf_num [9]);
tran (kme_internal_dak_kim_word[10], \kme_internal_dak_kim_word.vf_num [10]);
tran (kme_internal_dak_kim_word[11], \kme_internal_dak_kim_word.vf_num [11]);
tran (kme_internal_dak_kim_word[12], \kme_internal_dak_kim_word.pf_num [0]);
tran (kme_internal_dak_kim_word[13], \kme_internal_dak_kim_word.pf_num [1]);
tran (kme_internal_dak_kim_word[14], \kme_internal_dak_kim_word.pf_num [2]);
tran (kme_internal_dak_kim_word[15], \kme_internal_dak_kim_word.pf_num [3]);
tran (kme_internal_dak_kim_word[16], \kme_internal_dak_kim_word.vf_valid [0]);
tran (kme_internal_dak_kim_word[17], \kme_internal_dak_kim_word.validate_dak [0]);
tran (kme_internal_dak_kim_word[18], \kme_internal_dak_kim_word.unused [0]);
tran (kme_internal_dak_kim_word[19], \kme_internal_dak_kim_word.unused [1]);
tran (kme_internal_dak_kim_word[20], \kme_internal_dak_kim_word.unused [2]);
tran (kme_internal_dak_kim_word[21], \kme_internal_dak_kim_word.unused [3]);
tran (kme_internal_dak_kim_word[22], \kme_internal_dak_kim_word.unused [4]);
tran (kme_internal_dak_kim_word[23], \kme_internal_dak_kim_word.unused [5]);
tran (kme_internal_dak_kim_word[24], \kme_internal_dak_kim_word.unused [6]);
tran (kme_internal_dak_kim_word[25], \kme_internal_dak_kim_word.unused [7]);
tran (kme_internal_dak_kim_word[26], \kme_internal_dak_kim_word.dak_kim_entry.vf_valid [0]);
tran (kme_internal_dak_kim_word[27], \kme_internal_dak_kim_word.dak_kim_entry.vf_num [0]);
tran (kme_internal_dak_kim_word[28], \kme_internal_dak_kim_word.dak_kim_entry.vf_num [1]);
tran (kme_internal_dak_kim_word[29], \kme_internal_dak_kim_word.dak_kim_entry.vf_num [2]);
tran (kme_internal_dak_kim_word[30], \kme_internal_dak_kim_word.dak_kim_entry.vf_num [3]);
tran (kme_internal_dak_kim_word[31], \kme_internal_dak_kim_word.dak_kim_entry.vf_num [4]);
tran (kme_internal_dak_kim_word[32], \kme_internal_dak_kim_word.dak_kim_entry.vf_num [5]);
tran (kme_internal_dak_kim_word[33], \kme_internal_dak_kim_word.dak_kim_entry.vf_num [6]);
tran (kme_internal_dak_kim_word[34], \kme_internal_dak_kim_word.dak_kim_entry.vf_num [7]);
tran (kme_internal_dak_kim_word[35], \kme_internal_dak_kim_word.dak_kim_entry.vf_num [8]);
tran (kme_internal_dak_kim_word[36], \kme_internal_dak_kim_word.dak_kim_entry.vf_num [9]);
tran (kme_internal_dak_kim_word[37], \kme_internal_dak_kim_word.dak_kim_entry.vf_num [10]);
tran (kme_internal_dak_kim_word[38], \kme_internal_dak_kim_word.dak_kim_entry.vf_num [11]);
tran (kme_internal_dak_kim_word[39], \kme_internal_dak_kim_word.dak_kim_entry.pf_num [0]);
tran (kme_internal_dak_kim_word[40], \kme_internal_dak_kim_word.dak_kim_entry.pf_num [1]);
tran (kme_internal_dak_kim_word[41], \kme_internal_dak_kim_word.dak_kim_entry.pf_num [2]);
tran (kme_internal_dak_kim_word[42], \kme_internal_dak_kim_word.dak_kim_entry.pf_num [3]);
tran (kme_internal_dak_kim_word[43], \kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [0]);
tran (kme_internal_dak_kim_word[44], \kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [1]);
tran (kme_internal_dak_kim_word[45], \kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [2]);
tran (kme_internal_dak_kim_word[46], \kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [3]);
tran (kme_internal_dak_kim_word[47], \kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [4]);
tran (kme_internal_dak_kim_word[48], \kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [5]);
tran (kme_internal_dak_kim_word[49], \kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [6]);
tran (kme_internal_dak_kim_word[50], \kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [7]);
tran (kme_internal_dak_kim_word[51], \kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [8]);
tran (kme_internal_dak_kim_word[52], \kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [9]);
tran (kme_internal_dak_kim_word[53], \kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [10]);
tran (kme_internal_dak_kim_word[54], \kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [11]);
tran (kme_internal_dak_kim_word[55], \kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [12]);
tran (kme_internal_dak_kim_word[56], \kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [13]);
tran (kme_internal_dak_kim_word[57], \kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer [14]);
tran (kme_internal_dak_kim_word[58], \kme_internal_dak_kim_word.dak_kim_entry.ckv_length [0]);
tran (kme_internal_dak_kim_word[59], \kme_internal_dak_kim_word.dak_kim_entry.ckv_length [1]);
tran (kme_internal_dak_kim_word[60], \kme_internal_dak_kim_word.dak_kim_entry.label_index [0]);
tran (kme_internal_dak_kim_word[61], \kme_internal_dak_kim_word.dak_kim_entry.label_index [1]);
tran (kme_internal_dak_kim_word[62], \kme_internal_dak_kim_word.dak_kim_entry.label_index [2]);
tran (kme_internal_dak_kim_word[63], \kme_internal_dak_kim_word.dak_kim_entry.valid [0]);
tran (kme_internal_dek_kim_word[0], \kme_internal_dek_kim_word.vf_num [0]);
tran (kme_internal_dek_kim_word[1], \kme_internal_dek_kim_word.vf_num [1]);
tran (kme_internal_dek_kim_word[2], \kme_internal_dek_kim_word.vf_num [2]);
tran (kme_internal_dek_kim_word[3], \kme_internal_dek_kim_word.vf_num [3]);
tran (kme_internal_dek_kim_word[4], \kme_internal_dek_kim_word.vf_num [4]);
tran (kme_internal_dek_kim_word[5], \kme_internal_dek_kim_word.vf_num [5]);
tran (kme_internal_dek_kim_word[6], \kme_internal_dek_kim_word.vf_num [6]);
tran (kme_internal_dek_kim_word[7], \kme_internal_dek_kim_word.vf_num [7]);
tran (kme_internal_dek_kim_word[8], \kme_internal_dek_kim_word.vf_num [8]);
tran (kme_internal_dek_kim_word[9], \kme_internal_dek_kim_word.vf_num [9]);
tran (kme_internal_dek_kim_word[10], \kme_internal_dek_kim_word.vf_num [10]);
tran (kme_internal_dek_kim_word[11], \kme_internal_dek_kim_word.vf_num [11]);
tran (kme_internal_dek_kim_word[12], \kme_internal_dek_kim_word.pf_num [0]);
tran (kme_internal_dek_kim_word[13], \kme_internal_dek_kim_word.pf_num [1]);
tran (kme_internal_dek_kim_word[14], \kme_internal_dek_kim_word.pf_num [2]);
tran (kme_internal_dek_kim_word[15], \kme_internal_dek_kim_word.pf_num [3]);
tran (kme_internal_dek_kim_word[16], \kme_internal_dek_kim_word.vf_valid [0]);
tran (kme_internal_dek_kim_word[17], \kme_internal_dek_kim_word.validate_dek [0]);
tran (kme_internal_dek_kim_word[18], \kme_internal_dek_kim_word.missing_guid [0]);
tran (kme_internal_dek_kim_word[19], \kme_internal_dek_kim_word.missing_iv [0]);
tran (kme_internal_dek_kim_word[20], \kme_internal_dek_kim_word.unused [0]);
tran (kme_internal_dek_kim_word[21], \kme_internal_dek_kim_word.unused [1]);
tran (kme_internal_dek_kim_word[22], \kme_internal_dek_kim_word.unused [2]);
tran (kme_internal_dek_kim_word[23], \kme_internal_dek_kim_word.unused [3]);
tran (kme_internal_dek_kim_word[24], \kme_internal_dek_kim_word.unused [4]);
tran (kme_internal_dek_kim_word[25], \kme_internal_dek_kim_word.unused [5]);
tran (kme_internal_dek_kim_word[26], \kme_internal_dek_kim_word.dek_kim_entry.vf_valid [0]);
tran (kme_internal_dek_kim_word[27], \kme_internal_dek_kim_word.dek_kim_entry.vf_num [0]);
tran (kme_internal_dek_kim_word[28], \kme_internal_dek_kim_word.dek_kim_entry.vf_num [1]);
tran (kme_internal_dek_kim_word[29], \kme_internal_dek_kim_word.dek_kim_entry.vf_num [2]);
tran (kme_internal_dek_kim_word[30], \kme_internal_dek_kim_word.dek_kim_entry.vf_num [3]);
tran (kme_internal_dek_kim_word[31], \kme_internal_dek_kim_word.dek_kim_entry.vf_num [4]);
tran (kme_internal_dek_kim_word[32], \kme_internal_dek_kim_word.dek_kim_entry.vf_num [5]);
tran (kme_internal_dek_kim_word[33], \kme_internal_dek_kim_word.dek_kim_entry.vf_num [6]);
tran (kme_internal_dek_kim_word[34], \kme_internal_dek_kim_word.dek_kim_entry.vf_num [7]);
tran (kme_internal_dek_kim_word[35], \kme_internal_dek_kim_word.dek_kim_entry.vf_num [8]);
tran (kme_internal_dek_kim_word[36], \kme_internal_dek_kim_word.dek_kim_entry.vf_num [9]);
tran (kme_internal_dek_kim_word[37], \kme_internal_dek_kim_word.dek_kim_entry.vf_num [10]);
tran (kme_internal_dek_kim_word[38], \kme_internal_dek_kim_word.dek_kim_entry.vf_num [11]);
tran (kme_internal_dek_kim_word[39], \kme_internal_dek_kim_word.dek_kim_entry.pf_num [0]);
tran (kme_internal_dek_kim_word[40], \kme_internal_dek_kim_word.dek_kim_entry.pf_num [1]);
tran (kme_internal_dek_kim_word[41], \kme_internal_dek_kim_word.dek_kim_entry.pf_num [2]);
tran (kme_internal_dek_kim_word[42], \kme_internal_dek_kim_word.dek_kim_entry.pf_num [3]);
tran (kme_internal_dek_kim_word[43], \kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [0]);
tran (kme_internal_dek_kim_word[44], \kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [1]);
tran (kme_internal_dek_kim_word[45], \kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [2]);
tran (kme_internal_dek_kim_word[46], \kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [3]);
tran (kme_internal_dek_kim_word[47], \kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [4]);
tran (kme_internal_dek_kim_word[48], \kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [5]);
tran (kme_internal_dek_kim_word[49], \kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [6]);
tran (kme_internal_dek_kim_word[50], \kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [7]);
tran (kme_internal_dek_kim_word[51], \kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [8]);
tran (kme_internal_dek_kim_word[52], \kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [9]);
tran (kme_internal_dek_kim_word[53], \kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [10]);
tran (kme_internal_dek_kim_word[54], \kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [11]);
tran (kme_internal_dek_kim_word[55], \kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [12]);
tran (kme_internal_dek_kim_word[56], \kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [13]);
tran (kme_internal_dek_kim_word[57], \kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer [14]);
tran (kme_internal_dek_kim_word[58], \kme_internal_dek_kim_word.dek_kim_entry.ckv_length [0]);
tran (kme_internal_dek_kim_word[59], \kme_internal_dek_kim_word.dek_kim_entry.ckv_length [1]);
tran (kme_internal_dek_kim_word[60], \kme_internal_dek_kim_word.dek_kim_entry.label_index [0]);
tran (kme_internal_dek_kim_word[61], \kme_internal_dek_kim_word.dek_kim_entry.label_index [1]);
tran (kme_internal_dek_kim_word[62], \kme_internal_dek_kim_word.dek_kim_entry.label_index [2]);
tran (kme_internal_dek_kim_word[63], \kme_internal_dek_kim_word.dek_kim_entry.valid [0]);
tran (kme_internal_word0[0], \kme_internal_word0.tlv_type [0]);
tran (kme_internal_word0[1], \kme_internal_word0.tlv_type [1]);
tran (kme_internal_word0[2], \kme_internal_word0.tlv_type [2]);
tran (kme_internal_word0[3], \kme_internal_word0.tlv_type [3]);
tran (kme_internal_word0[4], \kme_internal_word0.tlv_type [4]);
tran (kme_internal_word0[5], \kme_internal_word0.tlv_type [5]);
tran (kme_internal_word0[6], \kme_internal_word0.tlv_type [6]);
tran (kme_internal_word0[7], \kme_internal_word0.tlv_type [7]);
tran (kme_internal_word0[8], \kme_internal_word0.tlv_len [0]);
tran (kme_internal_word0[9], \kme_internal_word0.tlv_len [1]);
tran (kme_internal_word0[10], \kme_internal_word0.tlv_len [2]);
tran (kme_internal_word0[11], \kme_internal_word0.tlv_len [3]);
tran (kme_internal_word0[12], \kme_internal_word0.tlv_len [4]);
tran (kme_internal_word0[13], \kme_internal_word0.tlv_len [5]);
tran (kme_internal_word0[14], \kme_internal_word0.tlv_len [6]);
tran (kme_internal_word0[15], \kme_internal_word0.tlv_len [7]);
tran (kme_internal_word0[16], \kme_internal_word0.tlv_seq_num [0]);
tran (kme_internal_word0[17], \kme_internal_word0.tlv_seq_num [1]);
tran (kme_internal_word0[18], \kme_internal_word0.tlv_seq_num [2]);
tran (kme_internal_word0[19], \kme_internal_word0.tlv_seq_num [3]);
tran (kme_internal_word0[20], \kme_internal_word0.tlv_seq_num [4]);
tran (kme_internal_word0[21], \kme_internal_word0.tlv_seq_num [5]);
tran (kme_internal_word0[22], \kme_internal_word0.tlv_seq_num [6]);
tran (kme_internal_word0[23], \kme_internal_word0.tlv_seq_num [7]);
tran (kme_internal_word0[24], \kme_internal_word0.tlv_eng_id [0]);
tran (kme_internal_word0[25], \kme_internal_word0.tlv_eng_id [1]);
tran (kme_internal_word0[26], \kme_internal_word0.tlv_eng_id [2]);
tran (kme_internal_word0[27], \kme_internal_word0.tlv_eng_id [3]);
tran (kme_internal_word0[28], \kme_internal_word0.tlv_frame_num [0]);
tran (kme_internal_word0[29], \kme_internal_word0.tlv_frame_num [1]);
tran (kme_internal_word0[30], \kme_internal_word0.tlv_frame_num [2]);
tran (kme_internal_word0[31], \kme_internal_word0.tlv_frame_num [3]);
tran (kme_internal_word0[32], \kme_internal_word0.tlv_frame_num [4]);
tran (kme_internal_word0[33], \kme_internal_word0.tlv_frame_num [5]);
tran (kme_internal_word0[34], \kme_internal_word0.tlv_frame_num [6]);
tran (kme_internal_word0[35], \kme_internal_word0.tlv_frame_num [7]);
tran (kme_internal_word0[36], \kme_internal_word0.tlv_frame_num [8]);
tran (kme_internal_word0[37], \kme_internal_word0.tlv_frame_num [9]);
tran (kme_internal_word0[38], \kme_internal_word0.tlv_frame_num [10]);
tran (kme_internal_word0[39], \kme_internal_word0.key_type [0]);
tran (kme_internal_word0[40], \kme_internal_word0.key_type [1]);
tran (kme_internal_word0[41], \kme_internal_word0.key_type [2]);
tran (kme_internal_word0[42], \kme_internal_word0.key_type [3]);
tran (kme_internal_word0[43], \kme_internal_word0.key_type [4]);
tran (kme_internal_word0[44], \kme_internal_word0.key_type [5]);
tran (kme_internal_word0[45], \kme_internal_word0.needs_dak [0]);
tran (kme_internal_word0[46], \kme_internal_word0.needs_dek [0]);
tran (kme_internal_word0[47], \kme_internal_word0.keyless_algos [0]);
tran (kme_internal_word0[48], \kme_internal_word0.kdf_dek_iter [0]);
tran (kme_internal_word0[49], \kme_internal_word0.resv0 [0]);
tran (kme_internal_word0[50], \kme_internal_word0.resv0 [1]);
tran (kme_internal_word0[51], \kme_internal_word0.resv0 [2]);
tran (kme_internal_word0[52], \kme_internal_word0.resv0 [3]);
tran (kme_internal_word0[53], \kme_internal_word0.resv0 [4]);
tran (kme_internal_word0[54], \kme_internal_word0.resv0 [5]);
tran (kme_internal_word0[55], \kme_internal_word0.resv0 [6]);
tran (kme_internal_word0[56], \kme_internal_word0.resv0 [7]);
tran (kme_internal_word0[57], \kme_internal_word0.resv0 [8]);
tran (kme_internal_word0[58], \kme_internal_word0.resv0 [9]);
tran (kme_internal_word0[59], \kme_internal_word0.resv0 [10]);
tran (kme_internal_word0[60], \kme_internal_word0.resv0 [11]);
tran (kme_internal_word0[61], \kme_internal_word0.resv0 [12]);
tran (kme_internal_word0[62], \kme_internal_word0.tlv_bip2 [0]);
tran (kme_internal_word0[63], \kme_internal_word0.tlv_bip2 [1]);
tran (fifo_in[64], \fifo_in.id [0]);
tran (fifo_in[65], \fifo_in.id [1]);
tran (fifo_in[66], \fifo_in.id [2]);
tran (fifo_in[67], \fifo_in.id [3]);
Q_BUF U0 ( .A(n1735), .Z(_zy_simnet_cio_7));
Q_ASSIGN U1 ( .B(stitcher_out[63]), .A(tlv_word0[63]));
Q_ASSIGN U2 ( .B(stitcher_out[63]), .A(tlv_word1[63]));
Q_ASSIGN U3 ( .B(stitcher_out[63]), .A(tlv_word2[63]));
Q_ASSIGN U4 ( .B(stitcher_out[63]), .A(frame_word[63]));
Q_ASSIGN U5 ( .B(stitcher_out[62]), .A(tlv_word0[62]));
Q_ASSIGN U6 ( .B(stitcher_out[62]), .A(tlv_word1[62]));
Q_ASSIGN U7 ( .B(stitcher_out[62]), .A(tlv_word2[62]));
Q_ASSIGN U8 ( .B(stitcher_out[62]), .A(frame_word[62]));
Q_ASSIGN U9 ( .B(stitcher_out[61]), .A(tlv_word0[61]));
Q_ASSIGN U10 ( .B(stitcher_out[61]), .A(tlv_word1[61]));
Q_ASSIGN U11 ( .B(stitcher_out[61]), .A(tlv_word2[61]));
Q_ASSIGN U12 ( .B(stitcher_out[61]), .A(frame_word[61]));
Q_ASSIGN U13 ( .B(stitcher_out[60]), .A(tlv_word0[60]));
Q_ASSIGN U14 ( .B(stitcher_out[60]), .A(tlv_word1[60]));
Q_ASSIGN U15 ( .B(stitcher_out[60]), .A(tlv_word2[60]));
Q_ASSIGN U16 ( .B(stitcher_out[60]), .A(frame_word[60]));
Q_ASSIGN U17 ( .B(stitcher_out[59]), .A(tlv_word0[59]));
Q_ASSIGN U18 ( .B(stitcher_out[59]), .A(tlv_word1[59]));
Q_ASSIGN U19 ( .B(stitcher_out[59]), .A(tlv_word2[59]));
Q_ASSIGN U20 ( .B(stitcher_out[59]), .A(frame_word[59]));
Q_ASSIGN U21 ( .B(stitcher_out[58]), .A(tlv_word0[58]));
Q_ASSIGN U22 ( .B(stitcher_out[58]), .A(tlv_word1[58]));
Q_ASSIGN U23 ( .B(stitcher_out[58]), .A(tlv_word2[58]));
Q_ASSIGN U24 ( .B(stitcher_out[58]), .A(frame_word[58]));
Q_ASSIGN U25 ( .B(stitcher_out[57]), .A(tlv_word0[57]));
Q_ASSIGN U26 ( .B(stitcher_out[57]), .A(tlv_word1[57]));
Q_ASSIGN U27 ( .B(stitcher_out[57]), .A(tlv_word2[57]));
Q_ASSIGN U28 ( .B(stitcher_out[57]), .A(frame_word[57]));
Q_ASSIGN U29 ( .B(stitcher_out[56]), .A(tlv_word0[56]));
Q_ASSIGN U30 ( .B(stitcher_out[56]), .A(tlv_word1[56]));
Q_ASSIGN U31 ( .B(stitcher_out[56]), .A(tlv_word2[56]));
Q_ASSIGN U32 ( .B(stitcher_out[56]), .A(frame_word[56]));
Q_ASSIGN U33 ( .B(stitcher_out[55]), .A(tlv_word0[55]));
Q_ASSIGN U34 ( .B(stitcher_out[55]), .A(tlv_word1[55]));
Q_ASSIGN U35 ( .B(stitcher_out[55]), .A(tlv_word2[55]));
Q_ASSIGN U36 ( .B(stitcher_out[55]), .A(frame_word[55]));
Q_ASSIGN U37 ( .B(stitcher_out[54]), .A(tlv_word0[54]));
Q_ASSIGN U38 ( .B(stitcher_out[54]), .A(tlv_word1[54]));
Q_ASSIGN U39 ( .B(stitcher_out[54]), .A(tlv_word2[54]));
Q_ASSIGN U40 ( .B(stitcher_out[54]), .A(frame_word[54]));
Q_ASSIGN U41 ( .B(stitcher_out[53]), .A(tlv_word0[53]));
Q_ASSIGN U42 ( .B(stitcher_out[53]), .A(tlv_word1[53]));
Q_ASSIGN U43 ( .B(stitcher_out[53]), .A(tlv_word2[53]));
Q_ASSIGN U44 ( .B(stitcher_out[53]), .A(frame_word[53]));
Q_ASSIGN U45 ( .B(stitcher_out[52]), .A(tlv_word0[52]));
Q_ASSIGN U46 ( .B(stitcher_out[52]), .A(tlv_word1[52]));
Q_ASSIGN U47 ( .B(stitcher_out[52]), .A(tlv_word2[52]));
Q_ASSIGN U48 ( .B(stitcher_out[52]), .A(frame_word[52]));
Q_ASSIGN U49 ( .B(stitcher_out[51]), .A(tlv_word0[51]));
Q_ASSIGN U50 ( .B(stitcher_out[51]), .A(tlv_word1[51]));
Q_ASSIGN U51 ( .B(stitcher_out[51]), .A(tlv_word2[51]));
Q_ASSIGN U52 ( .B(stitcher_out[51]), .A(frame_word[51]));
Q_ASSIGN U53 ( .B(stitcher_out[50]), .A(tlv_word0[50]));
Q_ASSIGN U54 ( .B(stitcher_out[50]), .A(tlv_word1[50]));
Q_ASSIGN U55 ( .B(stitcher_out[50]), .A(tlv_word2[50]));
Q_ASSIGN U56 ( .B(stitcher_out[50]), .A(frame_word[50]));
Q_ASSIGN U57 ( .B(stitcher_out[49]), .A(tlv_word0[49]));
Q_ASSIGN U58 ( .B(stitcher_out[49]), .A(tlv_word1[49]));
Q_ASSIGN U59 ( .B(stitcher_out[49]), .A(tlv_word2[49]));
Q_ASSIGN U60 ( .B(stitcher_out[49]), .A(frame_word[49]));
Q_ASSIGN U61 ( .B(stitcher_out[48]), .A(tlv_word0[48]));
Q_ASSIGN U62 ( .B(stitcher_out[48]), .A(tlv_word1[48]));
Q_ASSIGN U63 ( .B(stitcher_out[48]), .A(tlv_word2[48]));
Q_ASSIGN U64 ( .B(stitcher_out[48]), .A(frame_word[48]));
Q_ASSIGN U65 ( .B(stitcher_out[47]), .A(tlv_word0[47]));
Q_ASSIGN U66 ( .B(stitcher_out[47]), .A(tlv_word1[47]));
Q_ASSIGN U67 ( .B(stitcher_out[47]), .A(tlv_word2[47]));
Q_ASSIGN U68 ( .B(stitcher_out[47]), .A(frame_word[47]));
Q_ASSIGN U69 ( .B(stitcher_out[46]), .A(tlv_word0[46]));
Q_ASSIGN U70 ( .B(stitcher_out[46]), .A(tlv_word1[46]));
Q_ASSIGN U71 ( .B(stitcher_out[46]), .A(tlv_word2[46]));
Q_ASSIGN U72 ( .B(stitcher_out[46]), .A(frame_word[46]));
Q_ASSIGN U73 ( .B(stitcher_out[45]), .A(tlv_word0[45]));
Q_ASSIGN U74 ( .B(stitcher_out[45]), .A(tlv_word1[45]));
Q_ASSIGN U75 ( .B(stitcher_out[45]), .A(tlv_word2[45]));
Q_ASSIGN U76 ( .B(stitcher_out[45]), .A(frame_word[45]));
Q_ASSIGN U77 ( .B(stitcher_out[44]), .A(tlv_word0[44]));
Q_ASSIGN U78 ( .B(stitcher_out[44]), .A(tlv_word1[44]));
Q_ASSIGN U79 ( .B(stitcher_out[44]), .A(tlv_word2[44]));
Q_ASSIGN U80 ( .B(stitcher_out[44]), .A(frame_word[44]));
Q_ASSIGN U81 ( .B(stitcher_out[43]), .A(tlv_word0[43]));
Q_ASSIGN U82 ( .B(stitcher_out[43]), .A(tlv_word1[43]));
Q_ASSIGN U83 ( .B(stitcher_out[43]), .A(tlv_word2[43]));
Q_ASSIGN U84 ( .B(stitcher_out[43]), .A(frame_word[43]));
Q_ASSIGN U85 ( .B(stitcher_out[42]), .A(tlv_word0[42]));
Q_ASSIGN U86 ( .B(stitcher_out[42]), .A(tlv_word1[42]));
Q_ASSIGN U87 ( .B(stitcher_out[42]), .A(tlv_word2[42]));
Q_ASSIGN U88 ( .B(stitcher_out[42]), .A(frame_word[42]));
Q_ASSIGN U89 ( .B(stitcher_out[41]), .A(tlv_word0[41]));
Q_ASSIGN U90 ( .B(stitcher_out[41]), .A(tlv_word1[41]));
Q_ASSIGN U91 ( .B(stitcher_out[41]), .A(tlv_word2[41]));
Q_ASSIGN U92 ( .B(stitcher_out[41]), .A(frame_word[41]));
Q_ASSIGN U93 ( .B(stitcher_out[40]), .A(tlv_word0[40]));
Q_ASSIGN U94 ( .B(stitcher_out[40]), .A(tlv_word1[40]));
Q_ASSIGN U95 ( .B(stitcher_out[40]), .A(tlv_word2[40]));
Q_ASSIGN U96 ( .B(stitcher_out[40]), .A(frame_word[40]));
Q_ASSIGN U97 ( .B(stitcher_out[39]), .A(tlv_word0[39]));
Q_ASSIGN U98 ( .B(stitcher_out[39]), .A(tlv_word1[39]));
Q_ASSIGN U99 ( .B(stitcher_out[39]), .A(tlv_word2[39]));
Q_ASSIGN U100 ( .B(stitcher_out[39]), .A(frame_word[39]));
Q_ASSIGN U101 ( .B(stitcher_out[38]), .A(tlv_word0[38]));
Q_ASSIGN U102 ( .B(stitcher_out[38]), .A(tlv_word1[38]));
Q_ASSIGN U103 ( .B(stitcher_out[38]), .A(tlv_word2[38]));
Q_ASSIGN U104 ( .B(stitcher_out[38]), .A(frame_word[38]));
Q_ASSIGN U105 ( .B(stitcher_out[37]), .A(tlv_word0[37]));
Q_ASSIGN U106 ( .B(stitcher_out[37]), .A(tlv_word1[37]));
Q_ASSIGN U107 ( .B(stitcher_out[37]), .A(tlv_word2[37]));
Q_ASSIGN U108 ( .B(stitcher_out[37]), .A(frame_word[37]));
Q_ASSIGN U109 ( .B(stitcher_out[36]), .A(tlv_word0[36]));
Q_ASSIGN U110 ( .B(stitcher_out[36]), .A(tlv_word1[36]));
Q_ASSIGN U111 ( .B(stitcher_out[36]), .A(tlv_word2[36]));
Q_ASSIGN U112 ( .B(stitcher_out[36]), .A(frame_word[36]));
Q_ASSIGN U113 ( .B(stitcher_out[35]), .A(tlv_word0[35]));
Q_ASSIGN U114 ( .B(stitcher_out[35]), .A(tlv_word1[35]));
Q_ASSIGN U115 ( .B(stitcher_out[35]), .A(tlv_word2[35]));
Q_ASSIGN U116 ( .B(stitcher_out[35]), .A(frame_word[35]));
Q_ASSIGN U117 ( .B(stitcher_out[34]), .A(tlv_word0[34]));
Q_ASSIGN U118 ( .B(stitcher_out[34]), .A(tlv_word1[34]));
Q_ASSIGN U119 ( .B(stitcher_out[34]), .A(tlv_word2[34]));
Q_ASSIGN U120 ( .B(stitcher_out[34]), .A(frame_word[34]));
Q_ASSIGN U121 ( .B(stitcher_out[33]), .A(tlv_word0[33]));
Q_ASSIGN U122 ( .B(stitcher_out[33]), .A(tlv_word1[33]));
Q_ASSIGN U123 ( .B(stitcher_out[33]), .A(tlv_word2[33]));
Q_ASSIGN U124 ( .B(stitcher_out[33]), .A(frame_word[33]));
Q_ASSIGN U125 ( .B(stitcher_out[32]), .A(tlv_word0[32]));
Q_ASSIGN U126 ( .B(stitcher_out[32]), .A(tlv_word1[32]));
Q_ASSIGN U127 ( .B(stitcher_out[32]), .A(tlv_word2[32]));
Q_ASSIGN U128 ( .B(stitcher_out[32]), .A(frame_word[32]));
Q_ASSIGN U129 ( .B(stitcher_out[31]), .A(tlv_word0[31]));
Q_ASSIGN U130 ( .B(stitcher_out[31]), .A(tlv_word1[31]));
Q_ASSIGN U131 ( .B(stitcher_out[31]), .A(tlv_word2[31]));
Q_ASSIGN U132 ( .B(stitcher_out[31]), .A(frame_word[31]));
Q_ASSIGN U133 ( .B(stitcher_out[30]), .A(tlv_word0[30]));
Q_ASSIGN U134 ( .B(stitcher_out[30]), .A(tlv_word1[30]));
Q_ASSIGN U135 ( .B(stitcher_out[30]), .A(tlv_word2[30]));
Q_ASSIGN U136 ( .B(stitcher_out[30]), .A(frame_word[30]));
Q_ASSIGN U137 ( .B(stitcher_out[29]), .A(tlv_word0[29]));
Q_ASSIGN U138 ( .B(stitcher_out[29]), .A(tlv_word1[29]));
Q_ASSIGN U139 ( .B(stitcher_out[29]), .A(tlv_word2[29]));
Q_ASSIGN U140 ( .B(stitcher_out[29]), .A(frame_word[29]));
Q_ASSIGN U141 ( .B(stitcher_out[28]), .A(tlv_word0[28]));
Q_ASSIGN U142 ( .B(stitcher_out[28]), .A(tlv_word1[28]));
Q_ASSIGN U143 ( .B(stitcher_out[28]), .A(tlv_word2[28]));
Q_ASSIGN U144 ( .B(stitcher_out[28]), .A(frame_word[28]));
Q_ASSIGN U145 ( .B(stitcher_out[27]), .A(tlv_word0[27]));
Q_ASSIGN U146 ( .B(stitcher_out[27]), .A(tlv_word1[27]));
Q_ASSIGN U147 ( .B(stitcher_out[27]), .A(tlv_word2[27]));
Q_ASSIGN U148 ( .B(stitcher_out[27]), .A(frame_word[27]));
Q_ASSIGN U149 ( .B(stitcher_out[26]), .A(tlv_word0[26]));
Q_ASSIGN U150 ( .B(stitcher_out[26]), .A(tlv_word1[26]));
Q_ASSIGN U151 ( .B(stitcher_out[26]), .A(tlv_word2[26]));
Q_ASSIGN U152 ( .B(stitcher_out[26]), .A(frame_word[26]));
Q_ASSIGN U153 ( .B(stitcher_out[25]), .A(tlv_word0[25]));
Q_ASSIGN U154 ( .B(stitcher_out[25]), .A(tlv_word1[25]));
Q_ASSIGN U155 ( .B(stitcher_out[25]), .A(tlv_word2[25]));
Q_ASSIGN U156 ( .B(stitcher_out[25]), .A(frame_word[25]));
Q_ASSIGN U157 ( .B(stitcher_out[24]), .A(tlv_word0[24]));
Q_ASSIGN U158 ( .B(stitcher_out[24]), .A(tlv_word1[24]));
Q_ASSIGN U159 ( .B(stitcher_out[24]), .A(tlv_word2[24]));
Q_ASSIGN U160 ( .B(stitcher_out[24]), .A(frame_word[24]));
Q_ASSIGN U161 ( .B(stitcher_out[23]), .A(tlv_word0[23]));
Q_ASSIGN U162 ( .B(stitcher_out[23]), .A(tlv_word1[23]));
Q_ASSIGN U163 ( .B(stitcher_out[23]), .A(tlv_word2[23]));
Q_ASSIGN U164 ( .B(stitcher_out[23]), .A(frame_word[23]));
Q_ASSIGN U165 ( .B(stitcher_out[22]), .A(tlv_word0[22]));
Q_ASSIGN U166 ( .B(stitcher_out[22]), .A(tlv_word1[22]));
Q_ASSIGN U167 ( .B(stitcher_out[22]), .A(tlv_word2[22]));
Q_ASSIGN U168 ( .B(stitcher_out[22]), .A(frame_word[22]));
Q_ASSIGN U169 ( .B(stitcher_out[21]), .A(tlv_word0[21]));
Q_ASSIGN U170 ( .B(stitcher_out[21]), .A(tlv_word1[21]));
Q_ASSIGN U171 ( .B(stitcher_out[21]), .A(tlv_word2[21]));
Q_ASSIGN U172 ( .B(stitcher_out[21]), .A(frame_word[21]));
Q_ASSIGN U173 ( .B(stitcher_out[20]), .A(tlv_word0[20]));
Q_ASSIGN U174 ( .B(stitcher_out[20]), .A(tlv_word1[20]));
Q_ASSIGN U175 ( .B(stitcher_out[20]), .A(tlv_word2[20]));
Q_ASSIGN U176 ( .B(stitcher_out[20]), .A(frame_word[20]));
Q_ASSIGN U177 ( .B(stitcher_out[19]), .A(tlv_word0[19]));
Q_ASSIGN U178 ( .B(stitcher_out[19]), .A(tlv_word1[19]));
Q_ASSIGN U179 ( .B(stitcher_out[19]), .A(tlv_word2[19]));
Q_ASSIGN U180 ( .B(stitcher_out[19]), .A(frame_word[19]));
Q_ASSIGN U181 ( .B(stitcher_out[18]), .A(tlv_word0[18]));
Q_ASSIGN U182 ( .B(stitcher_out[18]), .A(tlv_word1[18]));
Q_ASSIGN U183 ( .B(stitcher_out[18]), .A(tlv_word2[18]));
Q_ASSIGN U184 ( .B(stitcher_out[18]), .A(frame_word[18]));
Q_ASSIGN U185 ( .B(stitcher_out[17]), .A(tlv_word0[17]));
Q_ASSIGN U186 ( .B(stitcher_out[17]), .A(tlv_word1[17]));
Q_ASSIGN U187 ( .B(stitcher_out[17]), .A(tlv_word2[17]));
Q_ASSIGN U188 ( .B(stitcher_out[17]), .A(frame_word[17]));
Q_ASSIGN U189 ( .B(stitcher_out[16]), .A(tlv_word0[16]));
Q_ASSIGN U190 ( .B(stitcher_out[16]), .A(tlv_word1[16]));
Q_ASSIGN U191 ( .B(stitcher_out[16]), .A(tlv_word2[16]));
Q_ASSIGN U192 ( .B(stitcher_out[16]), .A(frame_word[16]));
Q_ASSIGN U193 ( .B(stitcher_out[15]), .A(tlv_word0[15]));
Q_ASSIGN U194 ( .B(stitcher_out[15]), .A(tlv_word1[15]));
Q_ASSIGN U195 ( .B(stitcher_out[15]), .A(tlv_word2[15]));
Q_ASSIGN U196 ( .B(stitcher_out[15]), .A(frame_word[15]));
Q_ASSIGN U197 ( .B(stitcher_out[14]), .A(tlv_word0[14]));
Q_ASSIGN U198 ( .B(stitcher_out[14]), .A(tlv_word1[14]));
Q_ASSIGN U199 ( .B(stitcher_out[14]), .A(tlv_word2[14]));
Q_ASSIGN U200 ( .B(stitcher_out[14]), .A(frame_word[14]));
Q_ASSIGN U201 ( .B(stitcher_out[13]), .A(tlv_word0[13]));
Q_ASSIGN U202 ( .B(stitcher_out[13]), .A(tlv_word1[13]));
Q_ASSIGN U203 ( .B(stitcher_out[13]), .A(tlv_word2[13]));
Q_ASSIGN U204 ( .B(stitcher_out[13]), .A(frame_word[13]));
Q_ASSIGN U205 ( .B(stitcher_out[12]), .A(tlv_word0[12]));
Q_ASSIGN U206 ( .B(stitcher_out[12]), .A(tlv_word1[12]));
Q_ASSIGN U207 ( .B(stitcher_out[12]), .A(tlv_word2[12]));
Q_ASSIGN U208 ( .B(stitcher_out[12]), .A(frame_word[12]));
Q_ASSIGN U209 ( .B(stitcher_out[11]), .A(tlv_word0[11]));
Q_ASSIGN U210 ( .B(stitcher_out[11]), .A(tlv_word1[11]));
Q_ASSIGN U211 ( .B(stitcher_out[11]), .A(tlv_word2[11]));
Q_ASSIGN U212 ( .B(stitcher_out[11]), .A(frame_word[11]));
Q_ASSIGN U213 ( .B(stitcher_out[10]), .A(tlv_word0[10]));
Q_ASSIGN U214 ( .B(stitcher_out[10]), .A(tlv_word1[10]));
Q_ASSIGN U215 ( .B(stitcher_out[10]), .A(tlv_word2[10]));
Q_ASSIGN U216 ( .B(stitcher_out[10]), .A(frame_word[10]));
Q_ASSIGN U217 ( .B(stitcher_out[9]), .A(tlv_word0[9]));
Q_ASSIGN U218 ( .B(stitcher_out[9]), .A(tlv_word1[9]));
Q_ASSIGN U219 ( .B(stitcher_out[9]), .A(tlv_word2[9]));
Q_ASSIGN U220 ( .B(stitcher_out[9]), .A(frame_word[9]));
Q_ASSIGN U221 ( .B(stitcher_out[8]), .A(tlv_word0[8]));
Q_ASSIGN U222 ( .B(stitcher_out[8]), .A(tlv_word1[8]));
Q_ASSIGN U223 ( .B(stitcher_out[8]), .A(tlv_word2[8]));
Q_ASSIGN U224 ( .B(stitcher_out[8]), .A(frame_word[8]));
Q_ASSIGN U225 ( .B(stitcher_out[7]), .A(tlv_word0[7]));
Q_ASSIGN U226 ( .B(stitcher_out[7]), .A(tlv_word1[7]));
Q_ASSIGN U227 ( .B(stitcher_out[7]), .A(tlv_word2[7]));
Q_ASSIGN U228 ( .B(stitcher_out[7]), .A(frame_word[7]));
Q_ASSIGN U229 ( .B(stitcher_out[6]), .A(tlv_word0[6]));
Q_ASSIGN U230 ( .B(stitcher_out[6]), .A(tlv_word1[6]));
Q_ASSIGN U231 ( .B(stitcher_out[6]), .A(tlv_word2[6]));
Q_ASSIGN U232 ( .B(stitcher_out[6]), .A(frame_word[6]));
Q_ASSIGN U233 ( .B(stitcher_out[5]), .A(tlv_word0[5]));
Q_ASSIGN U234 ( .B(stitcher_out[5]), .A(tlv_word1[5]));
Q_ASSIGN U235 ( .B(stitcher_out[5]), .A(tlv_word2[5]));
Q_ASSIGN U236 ( .B(stitcher_out[5]), .A(frame_word[5]));
Q_ASSIGN U237 ( .B(stitcher_out[4]), .A(tlv_word0[4]));
Q_ASSIGN U238 ( .B(stitcher_out[4]), .A(tlv_word1[4]));
Q_ASSIGN U239 ( .B(stitcher_out[4]), .A(tlv_word2[4]));
Q_ASSIGN U240 ( .B(stitcher_out[4]), .A(frame_word[4]));
Q_ASSIGN U241 ( .B(stitcher_out[3]), .A(tlv_word0[3]));
Q_ASSIGN U242 ( .B(stitcher_out[3]), .A(tlv_word1[3]));
Q_ASSIGN U243 ( .B(stitcher_out[3]), .A(tlv_word2[3]));
Q_ASSIGN U244 ( .B(stitcher_out[3]), .A(frame_word[3]));
Q_ASSIGN U245 ( .B(stitcher_out[2]), .A(tlv_word0[2]));
Q_ASSIGN U246 ( .B(stitcher_out[2]), .A(tlv_word1[2]));
Q_ASSIGN U247 ( .B(stitcher_out[2]), .A(tlv_word2[2]));
Q_ASSIGN U248 ( .B(stitcher_out[2]), .A(frame_word[2]));
Q_ASSIGN U249 ( .B(stitcher_out[1]), .A(tlv_word0[1]));
Q_ASSIGN U250 ( .B(stitcher_out[1]), .A(tlv_word1[1]));
Q_ASSIGN U251 ( .B(stitcher_out[1]), .A(tlv_word2[1]));
Q_ASSIGN U252 ( .B(stitcher_out[1]), .A(frame_word[1]));
Q_ASSIGN U253 ( .B(stitcher_out[0]), .A(tlv_word0[0]));
Q_ASSIGN U254 ( .B(stitcher_out[0]), .A(tlv_word1[0]));
Q_ASSIGN U255 ( .B(stitcher_out[0]), .A(tlv_word2[0]));
Q_ASSIGN U256 ( .B(stitcher_out[0]), .A(frame_word[0]));
Q_BUF U257 ( .A(_zy_sva_key_type0_line5b_3_reset_or), .Z(_zy_sva_key_type0_line5a_2_reset_or));
Q_BUF U258 ( .A(_zy_sva_key_type1_line7a_4_reset_or), .Z(_zy_sva_key_type0_line5b_3_reset_or));
Q_BUF U259 ( .A(_zy_sva_key_type1_line7b_5_reset_or), .Z(_zy_sva_key_type1_line7a_4_reset_or));
Q_BUF U260 ( .A(_zy_sva_key_type1_line8a_6_reset_or), .Z(_zy_sva_key_type1_line7b_5_reset_or));
Q_BUF U261 ( .A(_zy_sva_key_type1_line8b_7_reset_or), .Z(_zy_sva_key_type1_line8a_6_reset_or));
Q_BUF U262 ( .A(_zy_sva_key_type1_line9_8_reset_or), .Z(_zy_sva_key_type1_line8b_7_reset_or));
Q_BUF U263 ( .A(_zy_sva_key_type1_line10_9_reset_or), .Z(_zy_sva_key_type1_line9_8_reset_or));
Q_BUF U264 ( .A(_zy_sva_key_type1_line11a_10_reset_or), .Z(_zy_sva_key_type1_line10_9_reset_or));
Q_BUF U265 ( .A(_zy_sva_key_type1_line11b_11_reset_or), .Z(_zy_sva_key_type1_line11a_10_reset_or));
Q_BUF U266 ( .A(_zy_sva_key_type1_line11c_12_reset_or), .Z(_zy_sva_key_type1_line11b_11_reset_or));
Q_BUF U267 ( .A(_zy_sva_key_type1_line11d_13_reset_or), .Z(_zy_sva_key_type1_line11c_12_reset_or));
Q_BUF U268 ( .A(_zy_sva_key_type1_line12a_14_reset_or), .Z(_zy_sva_key_type1_line11d_13_reset_or));
Q_BUF U269 ( .A(_zy_sva_key_type1_line12b_15_reset_or), .Z(_zy_sva_key_type1_line12a_14_reset_or));
Q_BUF U270 ( .A(_zy_sva_key_type9_line14_16_reset_or), .Z(_zy_sva_key_type1_line12b_15_reset_or));
Q_BUF U271 ( .A(_zy_sva_key_type9_line15_17_reset_or), .Z(_zy_sva_key_type9_line14_16_reset_or));
Q_BUF U272 ( .A(_zy_sva_key_type9_line16a_18_reset_or), .Z(_zy_sva_key_type9_line15_17_reset_or));
Q_BUF U273 ( .A(_zy_sva_key_type9_line16b_19_reset_or), .Z(_zy_sva_key_type9_line16a_18_reset_or));
Q_BUF U274 ( .A(_zy_sva_key_type9_line17a_20_reset_or), .Z(_zy_sva_key_type9_line16b_19_reset_or));
Q_BUF U275 ( .A(_zy_sva_key_type9_line17b_21_reset_or), .Z(_zy_sva_key_type9_line17a_20_reset_or));
Q_BUF U276 ( .A(_zy_sva_key_type9_line18a_22_reset_or), .Z(_zy_sva_key_type9_line17b_21_reset_or));
Q_BUF U277 ( .A(_zy_sva_key_type9_line18b_23_reset_or), .Z(_zy_sva_key_type9_line18a_22_reset_or));
Q_BUF U278 ( .A(_zy_sva_key_type9_line19a_24_reset_or), .Z(_zy_sva_key_type9_line18b_23_reset_or));
Q_BUF U279 ( .A(_zy_sva_key_type9_line19b_25_reset_or), .Z(_zy_sva_key_type9_line19a_24_reset_or));
Q_BUF U280 ( .A(_zy_sva_key_type9_line19c_26_reset_or), .Z(_zy_sva_key_type9_line19b_25_reset_or));
Q_BUF U281 ( .A(_zy_sva_key_type9_line19d_27_reset_or), .Z(_zy_sva_key_type9_line19c_26_reset_or));
Q_BUF U282 ( .A(_zy_sva_guid_miss_aux_cmd_0_28_reset_or), .Z(_zy_sva_key_type9_line19d_27_reset_or));
Q_BUF U283 ( .A(_zy_sva_guid_miss_aux_cmd_1_29_reset_or), .Z(_zy_sva_guid_miss_aux_cmd_0_28_reset_or));
Q_BUF U284 ( .A(_zy_sva_guid_miss_aux_cmd_2_30_reset_or), .Z(_zy_sva_guid_miss_aux_cmd_1_29_reset_or));
Q_BUF U285 ( .A(_zy_sva_guid_miss_aux_cmd_3_31_reset_or), .Z(_zy_sva_guid_miss_aux_cmd_2_30_reset_or));
Q_BUF U286 ( .A(_zy_sva_guid_miss_aux_cmd_iv_0_32_reset_or), .Z(_zy_sva_guid_miss_aux_cmd_3_31_reset_or));
Q_BUF U287 ( .A(_zy_sva_guid_miss_aux_cmd_iv_1_33_reset_or), .Z(_zy_sva_guid_miss_aux_cmd_iv_0_32_reset_or));
Q_BUF U288 ( .A(_zy_sva_guid_miss_aux_cmd_iv_2_34_reset_or), .Z(_zy_sva_guid_miss_aux_cmd_iv_1_33_reset_or));
Q_BUF U289 ( .A(_zy_sva_guid_miss_aux_cmd_iv_3_35_reset_or), .Z(_zy_sva_guid_miss_aux_cmd_iv_2_34_reset_or));
Q_BUF U290 ( .A(_zy_sva_iv_miss_aux_cmd_0_36_reset_or), .Z(_zy_sva_guid_miss_aux_cmd_iv_3_35_reset_or));
Q_BUF U291 ( .A(_zy_sva_iv_miss_aux_cmd_1_37_reset_or), .Z(_zy_sva_iv_miss_aux_cmd_0_36_reset_or));
Q_BUF U292 ( .A(_zy_sva_iv_miss_aux_cmd_guid_38_reset_or), .Z(_zy_sva_iv_miss_aux_cmd_1_37_reset_or));
Q_BUF U293 ( .A(_zy_sva_brcm_aux_cmd_39_reset_or), .Z(_zy_sva_iv_miss_aux_cmd_guid_38_reset_or));
Q_BUF U294 ( .A(_zy_sva_brcm_aux_cmd_iv_40_reset_or), .Z(_zy_sva_brcm_aux_cmd_39_reset_or));
Q_BUF U295 ( .A(_zy_sva_brcm_aux_cmd_guid_41_reset_or), .Z(_zy_sva_brcm_aux_cmd_iv_40_reset_or));
Q_BUF U296 ( .A(_zy_sva_brcm_aux_cmd_guid_iv_42_reset_or), .Z(_zy_sva_brcm_aux_cmd_guid_41_reset_or));
Q_BUF U297 ( .A(_zy_sva_brcm_key_type_43_reset_or), .Z(_zy_sva_brcm_aux_cmd_guid_iv_42_reset_or));
Q_BUF U298 ( .A(_zy_sva_brcm_aux_cmd_44_reset_or), .Z(_zy_sva_brcm_key_type_43_reset_or));
Q_BUF U299 ( .A(_zy_sva_brcm_aux_cmd_iv_45_reset_or), .Z(_zy_sva_brcm_aux_cmd_44_reset_or));
Q_BUF U300 ( .A(_zy_sva_brcm_aux_cmd_guid_46_reset_or), .Z(_zy_sva_brcm_aux_cmd_iv_45_reset_or));
Q_BUF U301 ( .A(_zy_sva_brcm_aux_cmd_guid_iv_47_reset_or), .Z(_zy_sva_brcm_aux_cmd_guid_46_reset_or));
Q_BUF U302 ( .A(_zy_sva_brcm_key_type_48_reset_or), .Z(_zy_sva_brcm_aux_cmd_guid_iv_47_reset_or));
Q_BUF U303 ( .A(_zy_sva_brcm_aux_cmd_49_reset_or), .Z(_zy_sva_brcm_key_type_48_reset_or));
Q_BUF U304 ( .A(_zy_sva_brcm_aux_cmd_iv_50_reset_or), .Z(_zy_sva_brcm_aux_cmd_49_reset_or));
Q_BUF U305 ( .A(_zy_sva_brcm_aux_cmd_guid_51_reset_or), .Z(_zy_sva_brcm_aux_cmd_iv_50_reset_or));
Q_BUF U306 ( .A(_zy_sva_brcm_aux_cmd_guid_iv_52_reset_or), .Z(_zy_sva_brcm_aux_cmd_guid_51_reset_or));
Q_BUF U307 ( .A(_zy_sva_brcm_key_type_53_reset_or), .Z(_zy_sva_brcm_aux_cmd_guid_iv_52_reset_or));
Q_BUF U308 ( .A(_zy_sva_brcm_aux_cmd_54_reset_or), .Z(_zy_sva_brcm_key_type_53_reset_or));
Q_BUF U309 ( .A(_zy_sva_brcm_aux_cmd_iv_55_reset_or), .Z(_zy_sva_brcm_aux_cmd_54_reset_or));
Q_BUF U310 ( .A(_zy_sva_brcm_aux_cmd_guid_56_reset_or), .Z(_zy_sva_brcm_aux_cmd_iv_55_reset_or));
Q_BUF U311 ( .A(_zy_sva_brcm_aux_cmd_guid_iv_57_reset_or), .Z(_zy_sva_brcm_aux_cmd_guid_56_reset_or));
Q_BUF U312 ( .A(_zy_sva_brcm_key_type_58_reset_or), .Z(_zy_sva_brcm_aux_cmd_guid_iv_57_reset_or));
Q_BUF U313 ( .A(_zy_sva_brcm_aux_cmd_59_reset_or), .Z(_zy_sva_brcm_key_type_58_reset_or));
Q_BUF U314 ( .A(_zy_sva_brcm_aux_cmd_iv_60_reset_or), .Z(_zy_sva_brcm_aux_cmd_59_reset_or));
Q_BUF U315 ( .A(_zy_sva_brcm_aux_cmd_guid_61_reset_or), .Z(_zy_sva_brcm_aux_cmd_iv_60_reset_or));
Q_BUF U316 ( .A(_zy_sva_brcm_aux_cmd_guid_iv_62_reset_or), .Z(_zy_sva_brcm_aux_cmd_guid_61_reset_or));
Q_BUF U317 ( .A(_zy_sva_brcm_key_type_63_reset_or), .Z(_zy_sva_brcm_aux_cmd_guid_iv_62_reset_or));
Q_BUF U318 ( .A(_zy_sva_brcm_aux_cmd_64_reset_or), .Z(_zy_sva_brcm_key_type_63_reset_or));
Q_BUF U319 ( .A(_zy_sva_brcm_aux_cmd_iv_65_reset_or), .Z(_zy_sva_brcm_aux_cmd_64_reset_or));
Q_BUF U320 ( .A(_zy_sva_brcm_aux_cmd_guid_66_reset_or), .Z(_zy_sva_brcm_aux_cmd_iv_65_reset_or));
Q_BUF U321 ( .A(_zy_sva_brcm_aux_cmd_guid_iv_67_reset_or), .Z(_zy_sva_brcm_aux_cmd_guid_66_reset_or));
Q_BUF U322 ( .A(_zy_sva_brcm_key_type_68_reset_or), .Z(_zy_sva_brcm_aux_cmd_guid_iv_67_reset_or));
Q_BUF U323 ( .A(_zy_sva_brcm_aux_cmd_69_reset_or), .Z(_zy_sva_brcm_key_type_68_reset_or));
Q_BUF U324 ( .A(_zy_sva_brcm_aux_cmd_iv_70_reset_or), .Z(_zy_sva_brcm_aux_cmd_69_reset_or));
Q_BUF U325 ( .A(_zy_sva_brcm_aux_cmd_guid_71_reset_or), .Z(_zy_sva_brcm_aux_cmd_iv_70_reset_or));
Q_BUF U326 ( .A(_zy_sva_brcm_aux_cmd_guid_iv_72_reset_or), .Z(_zy_sva_brcm_aux_cmd_guid_71_reset_or));
Q_BUF U327 ( .A(_zy_sva_brcm_key_type_73_reset_or), .Z(_zy_sva_brcm_aux_cmd_guid_iv_72_reset_or));
Q_BUF U328 ( .A(_zy_sva_brcm_aux_cmd_74_reset_or), .Z(_zy_sva_brcm_key_type_73_reset_or));
Q_BUF U329 ( .A(_zy_sva_brcm_aux_cmd_iv_75_reset_or), .Z(_zy_sva_brcm_aux_cmd_74_reset_or));
Q_BUF U330 ( .A(_zy_sva_brcm_aux_cmd_guid_76_reset_or), .Z(_zy_sva_brcm_aux_cmd_iv_75_reset_or));
Q_BUF U331 ( .A(_zy_sva_brcm_aux_cmd_guid_iv_77_reset_or), .Z(_zy_sva_brcm_aux_cmd_guid_76_reset_or));
Q_BUF U332 ( .A(_zy_sva_brcm_key_type_78_reset_or), .Z(_zy_sva_brcm_aux_cmd_guid_iv_77_reset_or));
Q_BUF U333 ( .A(_zy_sva_brcm_aux_cmd_79_reset_or), .Z(_zy_sva_brcm_key_type_78_reset_or));
Q_BUF U334 ( .A(_zy_sva_brcm_aux_cmd_iv_80_reset_or), .Z(_zy_sva_brcm_aux_cmd_79_reset_or));
Q_BUF U335 ( .A(_zy_sva_brcm_aux_cmd_guid_81_reset_or), .Z(_zy_sva_brcm_aux_cmd_iv_80_reset_or));
Q_BUF U336 ( .A(_zy_sva_brcm_aux_cmd_guid_iv_82_reset_or), .Z(_zy_sva_brcm_aux_cmd_guid_81_reset_or));
Q_BUF U337 ( .A(_zy_sva_brcm_key_type_83_reset_or), .Z(_zy_sva_brcm_aux_cmd_guid_iv_82_reset_or));
Q_BUF U338 ( .A(_zy_sva_brcm_aux_cmd_84_reset_or), .Z(_zy_sva_brcm_key_type_83_reset_or));
Q_BUF U339 ( .A(_zy_sva_brcm_aux_cmd_iv_85_reset_or), .Z(_zy_sva_brcm_aux_cmd_84_reset_or));
Q_BUF U340 ( .A(_zy_sva_brcm_aux_cmd_guid_86_reset_or), .Z(_zy_sva_brcm_aux_cmd_iv_85_reset_or));
Q_BUF U341 ( .A(_zy_sva_brcm_aux_cmd_guid_iv_87_reset_or), .Z(_zy_sva_brcm_aux_cmd_guid_86_reset_or));
Q_BUF U342 ( .A(_zy_sva_brcm_key_type_88_reset_or), .Z(_zy_sva_brcm_aux_cmd_guid_iv_87_reset_or));
Q_BUF U343 ( .A(_zy_sva_brcm_aux_cmd_89_reset_or), .Z(_zy_sva_brcm_key_type_88_reset_or));
Q_BUF U344 ( .A(_zy_sva_brcm_aux_cmd_iv_90_reset_or), .Z(_zy_sva_brcm_aux_cmd_89_reset_or));
Q_BUF U345 ( .A(_zy_sva_brcm_aux_cmd_guid_91_reset_or), .Z(_zy_sva_brcm_aux_cmd_iv_90_reset_or));
Q_BUF U346 ( .A(_zy_sva_brcm_aux_cmd_guid_iv_92_reset_or), .Z(_zy_sva_brcm_aux_cmd_guid_91_reset_or));
Q_BUF U347 ( .A(_zy_sva_brcm_key_type_93_reset_or), .Z(_zy_sva_brcm_aux_cmd_guid_iv_92_reset_or));
Q_BUF U348 ( .A(_zy_sva_brcm_aux_cmd_94_reset_or), .Z(_zy_sva_brcm_key_type_93_reset_or));
Q_BUF U349 ( .A(_zy_sva_brcm_aux_cmd_iv_95_reset_or), .Z(_zy_sva_brcm_aux_cmd_94_reset_or));
Q_BUF U350 ( .A(_zy_sva_brcm_aux_cmd_guid_96_reset_or), .Z(_zy_sva_brcm_aux_cmd_iv_95_reset_or));
Q_BUF U351 ( .A(_zy_sva_brcm_aux_cmd_guid_iv_97_reset_or), .Z(_zy_sva_brcm_aux_cmd_guid_96_reset_or));
Q_BUF U352 ( .A(_zy_sva_brcm_key_type_98_reset_or), .Z(_zy_sva_brcm_aux_cmd_guid_iv_97_reset_or));
Q_BUF U353 ( .A(_zy_sva_brcm_aux_cmd_99_reset_or), .Z(_zy_sva_brcm_key_type_98_reset_or));
Q_BUF U354 ( .A(_zy_sva_brcm_aux_cmd_iv_100_reset_or), .Z(_zy_sva_brcm_aux_cmd_99_reset_or));
Q_BUF U355 ( .A(_zy_sva_brcm_aux_cmd_guid_101_reset_or), .Z(_zy_sva_brcm_aux_cmd_iv_100_reset_or));
Q_BUF U356 ( .A(_zy_sva_brcm_aux_cmd_guid_iv_102_reset_or), .Z(_zy_sva_brcm_aux_cmd_guid_101_reset_or));
Q_BUF U357 ( .A(_zy_sva_brcm_key_type_103_reset_or), .Z(_zy_sva_brcm_aux_cmd_guid_iv_102_reset_or));
Q_BUF U358 ( .A(_zy_sva_brcm_aux_cmd_104_reset_or), .Z(_zy_sva_brcm_key_type_103_reset_or));
Q_BUF U359 ( .A(_zy_sva_brcm_aux_cmd_iv_105_reset_or), .Z(_zy_sva_brcm_aux_cmd_104_reset_or));
Q_BUF U360 ( .A(_zy_sva_brcm_aux_cmd_guid_106_reset_or), .Z(_zy_sva_brcm_aux_cmd_iv_105_reset_or));
Q_BUF U361 ( .A(_zy_sva_brcm_aux_cmd_guid_iv_107_reset_or), .Z(_zy_sva_brcm_aux_cmd_guid_106_reset_or));
Q_BUF U362 ( .A(_zy_sva_brcm_key_type_108_reset_or), .Z(_zy_sva_brcm_aux_cmd_guid_iv_107_reset_or));
Q_BUF U363 ( .A(_zy_sva_brcm_kdf_ops_109_reset_or), .Z(_zy_sva_brcm_key_type_108_reset_or));
Q_BUF U364 ( .A(_zy_sva_brcm_kdf_ops_110_reset_or), .Z(_zy_sva_brcm_kdf_ops_109_reset_or));
Q_BUF U365 ( .A(_zy_sva_brcm_kdf_ops_111_reset_or), .Z(_zy_sva_brcm_kdf_ops_110_reset_or));
Q_BUF U366 ( .A(_zy_sva_brcm_kdf_ops_112_reset_or), .Z(_zy_sva_brcm_kdf_ops_111_reset_or));
Q_BUF U367 ( .A(_zy_sva_brcm_kdf_ops_113_reset_or), .Z(_zy_sva_brcm_kdf_ops_112_reset_or));
Q_BUF U368 ( .A(_zy_sva_brcm_kdf_ops_114_reset_or), .Z(_zy_sva_brcm_kdf_ops_113_reset_or));
Q_BUF U369 ( .A(_zy_sva_brcm_kdf_ops_115_reset_or), .Z(_zy_sva_brcm_kdf_ops_114_reset_or));
Q_BUF U370 ( .A(_zy_sva_brcm_kdf_ops_116_reset_or), .Z(_zy_sva_brcm_kdf_ops_115_reset_or));
Q_BUF U371 ( .A(_zy_sva_brcm_kdf_ops_117_reset_or), .Z(_zy_sva_brcm_kdf_ops_116_reset_or));
Q_BUF U372 ( .A(_zy_sva_brcm_kdf_ops_118_reset_or), .Z(_zy_sva_brcm_kdf_ops_117_reset_or));
Q_BUF U373 ( .A(_zy_sva_brcm_kdf_ops_119_reset_or), .Z(_zy_sva_brcm_kdf_ops_118_reset_or));
Q_BUF U374 ( .A(_zy_sva_brcm_kdf_ops_120_reset_or), .Z(_zy_sva_brcm_kdf_ops_119_reset_or));
Q_BUF U375 ( .A(_zy_sva_brcm_kdf_ops_121_reset_or), .Z(_zy_sva_brcm_kdf_ops_120_reset_or));
Q_BUF U376 ( .A(_zy_sva_brcm_kdf_ops_122_reset_or), .Z(_zy_sva_brcm_kdf_ops_121_reset_or));
Q_BUF U377 ( .A(_zy_sva_brcm_kdf_ops_123_reset_or), .Z(_zy_sva_brcm_kdf_ops_122_reset_or));
Q_BUF U378 ( .A(_zy_sva_brcm_kdf_ops_124_reset_or), .Z(_zy_sva_brcm_kdf_ops_123_reset_or));
Q_BUF U379 ( .A(_zy_sva_null_gcm_125_reset_or), .Z(_zy_sva_brcm_kdf_ops_124_reset_or));
Q_BUF U380 ( .A(_zy_sva_sha_gcm_126_reset_or), .Z(_zy_sva_null_gcm_125_reset_or));
Q_BUF U381 ( .A(_zy_sva_null_xts_127_reset_or), .Z(_zy_sva_sha_gcm_126_reset_or));
Q_BUF U382 ( .A(_zy_sva_sha_xts_128_reset_or), .Z(_zy_sva_null_xts_127_reset_or));
Q_BUF U383 ( .A(_zy_sva_null_null_129_reset_or), .Z(_zy_sva_sha_xts_128_reset_or));
Q_BUF U384 ( .A(_zy_sva_sha_null_130_reset_or), .Z(_zy_sva_null_null_129_reset_or));
Q_BUF U385 ( .A(_zy_sva_hmac_gcm_131_reset_or), .Z(_zy_sva_sha_null_130_reset_or));
Q_BUF U386 ( .A(_zy_sva_hmac_xts_132_reset_or), .Z(_zy_sva_hmac_gcm_131_reset_or));
Q_BUF U387 ( .A(_zy_sva_hmac_null_133_reset_or), .Z(_zy_sva_hmac_xts_132_reset_or));
Q_BUF U388 ( .A(_zy_sva_null_gcm_134_reset_or), .Z(_zy_sva_hmac_null_133_reset_or));
Q_BUF U389 ( .A(_zy_sva_sha_gcm_135_reset_or), .Z(_zy_sva_null_gcm_134_reset_or));
Q_BUF U390 ( .A(_zy_sva_null_xts_136_reset_or), .Z(_zy_sva_sha_gcm_135_reset_or));
Q_BUF U391 ( .A(_zy_sva_sha_xts_137_reset_or), .Z(_zy_sva_null_xts_136_reset_or));
Q_BUF U392 ( .A(_zy_sva_null_null_138_reset_or), .Z(_zy_sva_sha_xts_137_reset_or));
Q_BUF U393 ( .A(_zy_sva_sha_null_139_reset_or), .Z(_zy_sva_null_null_138_reset_or));
Q_BUF U394 ( .A(_zy_sva_hmac_gcm_140_reset_or), .Z(_zy_sva_sha_null_139_reset_or));
Q_BUF U395 ( .A(_zy_sva_hmac_xts_141_reset_or), .Z(_zy_sva_hmac_gcm_140_reset_or));
Q_BUF U396 ( .A(_zy_sva_hmac_null_142_reset_or), .Z(_zy_sva_hmac_xts_141_reset_or));
Q_BUF U397 ( .A(_zy_sva_null_gcm_143_reset_or), .Z(_zy_sva_hmac_null_142_reset_or));
Q_BUF U398 ( .A(_zy_sva_sha_gcm_144_reset_or), .Z(_zy_sva_null_gcm_143_reset_or));
Q_BUF U399 ( .A(_zy_sva_null_xts_145_reset_or), .Z(_zy_sva_sha_gcm_144_reset_or));
Q_BUF U400 ( .A(_zy_sva_sha_xts_146_reset_or), .Z(_zy_sva_null_xts_145_reset_or));
Q_BUF U401 ( .A(_zy_sva_null_null_147_reset_or), .Z(_zy_sva_sha_xts_146_reset_or));
Q_BUF U402 ( .A(_zy_sva_sha_null_148_reset_or), .Z(_zy_sva_null_null_147_reset_or));
Q_BUF U403 ( .A(_zy_sva_hmac_gcm_149_reset_or), .Z(_zy_sva_sha_null_148_reset_or));
Q_BUF U404 ( .A(_zy_sva_hmac_xts_150_reset_or), .Z(_zy_sva_hmac_gcm_149_reset_or));
Q_BUF U405 ( .A(_zy_sva_hmac_null_151_reset_or), .Z(_zy_sva_hmac_xts_150_reset_or));
Q_BUF U406 ( .A(_zy_sva_null_gcm_152_reset_or), .Z(_zy_sva_hmac_null_151_reset_or));
Q_BUF U407 ( .A(_zy_sva_sha_gcm_153_reset_or), .Z(_zy_sva_null_gcm_152_reset_or));
Q_BUF U408 ( .A(_zy_sva_null_xts_154_reset_or), .Z(_zy_sva_sha_gcm_153_reset_or));
Q_BUF U409 ( .A(_zy_sva_sha_xts_155_reset_or), .Z(_zy_sva_null_xts_154_reset_or));
Q_BUF U410 ( .A(_zy_sva_null_null_156_reset_or), .Z(_zy_sva_sha_xts_155_reset_or));
Q_BUF U411 ( .A(_zy_sva_sha_null_157_reset_or), .Z(_zy_sva_null_null_156_reset_or));
Q_BUF U412 ( .A(_zy_sva_hmac_gcm_158_reset_or), .Z(_zy_sva_sha_null_157_reset_or));
Q_BUF U413 ( .A(_zy_sva_hmac_xts_159_reset_or), .Z(_zy_sva_hmac_gcm_158_reset_or));
Q_BUF U414 ( .A(_zy_sva_hmac_null_160_reset_or), .Z(_zy_sva_hmac_xts_159_reset_or));
Q_BUF U415 ( .A(_zy_sva_null_gcm_161_reset_or), .Z(_zy_sva_hmac_null_160_reset_or));
Q_BUF U416 ( .A(_zy_sva_sha_gcm_162_reset_or), .Z(_zy_sva_null_gcm_161_reset_or));
Q_BUF U417 ( .A(_zy_sva_null_xts_163_reset_or), .Z(_zy_sva_sha_gcm_162_reset_or));
Q_BUF U418 ( .A(_zy_sva_sha_xts_164_reset_or), .Z(_zy_sva_null_xts_163_reset_or));
Q_BUF U419 ( .A(_zy_sva_null_null_165_reset_or), .Z(_zy_sva_sha_xts_164_reset_or));
Q_BUF U420 ( .A(_zy_sva_sha_null_166_reset_or), .Z(_zy_sva_null_null_165_reset_or));
Q_BUF U421 ( .A(_zy_sva_hmac_gcm_167_reset_or), .Z(_zy_sva_sha_null_166_reset_or));
Q_BUF U422 ( .A(_zy_sva_hmac_xts_168_reset_or), .Z(_zy_sva_hmac_gcm_167_reset_or));
Q_BUF U423 ( .A(_zy_sva_hmac_null_169_reset_or), .Z(_zy_sva_hmac_xts_168_reset_or));
Q_BUF U424 ( .A(_zy_sva_null_gcm_170_reset_or), .Z(_zy_sva_hmac_null_169_reset_or));
Q_BUF U425 ( .A(_zy_sva_sha_gcm_171_reset_or), .Z(_zy_sva_null_gcm_170_reset_or));
Q_BUF U426 ( .A(_zy_sva_null_xts_172_reset_or), .Z(_zy_sva_sha_gcm_171_reset_or));
Q_BUF U427 ( .A(_zy_sva_sha_xts_173_reset_or), .Z(_zy_sva_null_xts_172_reset_or));
Q_BUF U428 ( .A(_zy_sva_null_null_174_reset_or), .Z(_zy_sva_sha_xts_173_reset_or));
Q_BUF U429 ( .A(_zy_sva_sha_null_175_reset_or), .Z(_zy_sva_null_null_174_reset_or));
Q_BUF U430 ( .A(_zy_sva_hmac_gcm_176_reset_or), .Z(_zy_sva_sha_null_175_reset_or));
Q_BUF U431 ( .A(_zy_sva_hmac_xts_177_reset_or), .Z(_zy_sva_hmac_gcm_176_reset_or));
Q_BUF U432 ( .A(_zy_sva_hmac_null_178_reset_or), .Z(_zy_sva_hmac_xts_177_reset_or));
Q_BUF U433 ( .A(_zy_sva_key_type0_line4_1_reset_or), .Z(_zy_sva_hmac_null_178_reset_or));
Q_AN02 U434 ( .A0(n144), .A1(n706), .Z(n1));
Q_AN02 U435 ( .A0(n144), .A1(n3), .Z(n2));
Q_INV U436 ( .A(n528), .Z(n3));
Q_OR02 U437 ( .A0(n5), .A1(int_tlv_counter[5]), .Z(n4));
Q_INV U438 ( .A(n6), .Z(n5));
Q_AN02 U439 ( .A0(int_tlv_counter[4]), .A1(n7), .Z(n6));
Q_INV U440 ( .A(n8), .Z(n7));
Q_OR02 U441 ( .A0(n9), .A1(int_tlv_counter[3]), .Z(n8));
Q_INV U442 ( .A(n10), .Z(n9));
Q_AN02 U443 ( .A0(int_tlv_counter[2]), .A1(int_tlv_counter[1]), .Z(n10));
Q_AN02 U444 ( .A0(int_tlv_counter[4]), .A1(n12), .Z(n11));
Q_AN02 U445 ( .A0(int_tlv_counter[3]), .A1(int_tlv_counter[2]), .Z(n12));
Q_OR02 U446 ( .A0(n14), .A1(int_tlv_counter[5]), .Z(n13));
Q_INV U447 ( .A(n15), .Z(n14));
Q_AN02 U448 ( .A0(int_tlv_counter[4]), .A1(n16), .Z(n15));
Q_INV U449 ( .A(n17), .Z(n16));
Q_OR02 U450 ( .A0(n18), .A1(int_tlv_counter[3]), .Z(n17));
Q_INV U451 ( .A(n19), .Z(n18));
Q_AN02 U452 ( .A0(int_tlv_counter[2]), .A1(n20), .Z(n19));
Q_AN02 U453 ( .A0(int_tlv_counter[1]), .A1(n682), .Z(n20));
Q_AN02 U454 ( .A0(aux_key_type[2]), .A1(n22), .Z(n21));
Q_AN02 U455 ( .A0(aux_key_type[1]), .A1(aux_key_type[0]), .Z(n22));
Q_OR02 U456 ( .A0(n493), .A1(int_tlv_counter[4]), .Z(n23));
Q_OR02 U457 ( .A0(n73), .A1(n64), .Z(n24));
Q_AN02 U458 ( .A0(n139), .A1(n144), .Z(n25));
Q_OR02 U459 ( .A0(n27), .A1(n704), .Z(n26));
Q_OR02 U460 ( .A0(n28), .A1(int_tlv_counter[5]), .Z(n27));
Q_OR02 U461 ( .A0(n29), .A1(int_tlv_counter[4]), .Z(n28));
Q_OR02 U462 ( .A0(n30), .A1(int_tlv_counter[3]), .Z(n29));
Q_OR02 U463 ( .A0(n526), .A1(n2135), .Z(n30));
Q_OR02 U464 ( .A0(n139), .A1(n704), .Z(n31));
Q_INV U465 ( .A(n1708), .Z(n32));
Q_INV U466 ( .A(n2112), .Z(n33));
Q_INV U467 ( .A(n638), .Z(n34));
Q_INV U468 ( .A(n2122), .Z(n35));
Q_INV U469 ( .A(n116), .Z(n36));
Q_INV U470 ( .A(n2030), .Z(n37));
Q_INV U471 ( .A(n2118), .Z(n38));
Q_INV U472 ( .A(n2070), .Z(n39));
Q_INV U473 ( .A(n2055), .Z(n40));
Q_INV U474 ( .A(n2056), .Z(n41));
Q_INV U475 ( .A(n662), .Z(n42));
Q_INV U476 ( .A(n550), .Z(n43));
Q_INV U477 ( .A(n221), .Z(n44));
Q_INV U478 ( .A(n478), .Z(n45));
Q_INV U479 ( .A(n511), .Z(n46));
Q_OR02 U480 ( .A0(int_tlv_counter[3]), .A1(int_tlv_counter[4]), .Z(n92));
Q_MX02 U481 ( .S(int_tlv_counter[1]), .A0(n79), .A1(n92), .Z(n52));
Q_OR02 U482 ( .A0(int_tlv_counter[2]), .A1(n36), .Z(n88));
Q_OR02 U483 ( .A0(n2136), .A1(n88), .Z(n53));
Q_MX02 U484 ( .S(int_tlv_counter[0]), .A0(n53), .A1(n52), .Z(n54));
Q_AN02 U485 ( .A0(n36), .A1(int_tlv_counter[2]), .Z(n56));
Q_AN02 U486 ( .A0(int_tlv_counter[3]), .A1(int_tlv_counter[4]), .Z(n61));
Q_INV U487 ( .A(n76), .Z(n55));
Q_OR03 U488 ( .A0(n56), .A1(n55), .A2(n2136), .Z(n69));
Q_INV U489 ( .A(n61), .Z(n75));
Q_OR02 U490 ( .A0(n75), .A1(int_tlv_counter[1]), .Z(n57));
Q_AN03 U491 ( .A0(n69), .A1(n57), .A2(int_tlv_counter[0]), .Z(n58));
Q_OR02 U492 ( .A0(int_tlv_counter[2]), .A1(n92), .Z(n87));
Q_OR02 U493 ( .A0(int_tlv_counter[1]), .A1(n87), .Z(n65));
Q_NR02 U494 ( .A0(n58), .A1(n98), .Z(n59));
Q_MX02 U495 ( .S(int_tlv_counter[5]), .A0(n59), .A1(n54), .Z(n60));
Q_OR02 U496 ( .A0(n190), .A1(n60), .Z(n48));
Q_INV U497 ( .A(n48), .Z(fifo_in[69]));
Q_MX02 U498 ( .S(int_tlv_counter[1]), .A0(n61), .A1(n95), .Z(n62));
Q_MX02 U499 ( .S(int_tlv_counter[0]), .A0(n65), .A1(n62), .Z(n63));
Q_OR03 U500 ( .A0(n190), .A1(int_tlv_counter[5]), .A2(n63), .Z(n64));
Q_OR02 U501 ( .A0(n682), .A1(n65), .Z(n66));
Q_INV U502 ( .A(n92), .Z(n67));
Q_OR02 U503 ( .A0(n67), .A1(int_tlv_counter[1]), .Z(n68));
Q_AN03 U504 ( .A0(n69), .A1(n68), .A2(int_tlv_counter[0]), .Z(n70));
Q_NR02 U505 ( .A0(n70), .A1(n98), .Z(n71));
Q_MX02 U506 ( .S(int_tlv_counter[5]), .A0(n71), .A1(n66), .Z(n72));
Q_OR02 U507 ( .A0(n190), .A1(n72), .Z(n73));
Q_INV U508 ( .A(n73), .Z(n49));
Q_OR02 U509 ( .A0(n511), .A1(n92), .Z(n74));
Q_ND02 U510 ( .A0(n113), .A1(int_tlv_counter[2]), .Z(n77));
Q_OR02 U511 ( .A0(n75), .A1(int_tlv_counter[2]), .Z(n76));
Q_AN02 U512 ( .A0(n77), .A1(n76), .Z(n78));
Q_ND02 U513 ( .A0(n116), .A1(int_tlv_counter[2]), .Z(n80));
Q_OR02 U514 ( .A0(int_tlv_counter[4]), .A1(int_tlv_counter[2]), .Z(n79));
Q_AN02 U515 ( .A0(n80), .A1(n79), .Z(n81));
Q_MX02 U516 ( .S(int_tlv_counter[1]), .A0(n81), .A1(n78), .Z(n82));
Q_OA21 U517 ( .A0(n82), .A1(n682), .B0(n83), .Z(n84));
Q_INV U518 ( .A(n98), .Z(n83));
Q_MX02 U519 ( .S(int_tlv_counter[5]), .A0(n84), .A1(n74), .Z(n85));
Q_OR02 U520 ( .A0(n190), .A1(n85), .Z(n86));
Q_INV U521 ( .A(n86), .Z(n50));
Q_MX02 U522 ( .S(int_tlv_counter[1]), .A0(n88), .A1(n87), .Z(n89));
Q_OR02 U523 ( .A0(n682), .A1(n89), .Z(n90));
Q_AN02 U524 ( .A0(int_tlv_counter[2]), .A1(int_tlv_counter[4]), .Z(n91));
Q_OR02 U525 ( .A0(n92), .A1(n2135), .Z(n95));
Q_XOR2 U526 ( .A0(int_tlv_counter[3]), .A1(n688), .Z(n93));
Q_OR02 U527 ( .A0(n93), .A1(int_tlv_counter[2]), .Z(n94));
Q_ND02 U528 ( .A0(n95), .A1(n94), .Z(n96));
Q_MX02 U529 ( .S(int_tlv_counter[1]), .A0(n96), .A1(n91), .Z(n97));
Q_AN02 U530 ( .A0(n97), .A1(int_tlv_counter[0]), .Z(n99));
Q_NR02 U531 ( .A0(n65), .A1(int_tlv_counter[0]), .Z(n98));
Q_NR02 U532 ( .A0(n99), .A1(n98), .Z(n100));
Q_MX02 U533 ( .S(int_tlv_counter[5]), .A0(n100), .A1(n90), .Z(n101));
Q_OR02 U534 ( .A0(n190), .A1(n101), .Z(n102));
Q_INV U535 ( .A(n102), .Z(n51));
Q_AO21 U536 ( .A0(n48), .A1(fifo_in[64]), .B0(n108), .Z(nxt_fifo_in_id[0]));
Q_AO21 U537 ( .A0(n48), .A1(fifo_in[65]), .B0(n107), .Z(nxt_fifo_in_id[1]));
Q_AO21 U538 ( .A0(n48), .A1(fifo_in[66]), .B0(n106), .Z(nxt_fifo_in_id[2]));
Q_AO21 U539 ( .A0(n48), .A1(fifo_in[67]), .B0(n104), .Z(nxt_fifo_in_id[3]));
Q_ND02 U540 ( .A0(n86), .A1(n102), .Z(n105));
Q_OR02 U541 ( .A0(n49), .A1(n105), .Z(n103));
Q_XNR2 U542 ( .A0(n64), .A1(n103), .Z(n104));
Q_XNR2 U543 ( .A0(n73), .A1(n105), .Z(n106));
Q_XNR2 U544 ( .A0(n50), .A1(n102), .Z(n107));
Q_MX02 U545 ( .S(n24), .A0(n50), .A1(n51), .Z(n108));
Q_NR02 U546 ( .A0(n190), .A1(n2032), .Z(fifo_in[70]));
Q_AN02 U547 ( .A0(int_tlv_counter[4]), .A1(n697), .Z(n113));
Q_AN03 U548 ( .A0(n706), .A1(n113), .A2(n114), .Z(n111));
Q_AN03 U549 ( .A0(int_tlv_counter[2]), .A1(n2136), .A2(int_tlv_counter[0]), .Z(n114));
Q_AN02 U550 ( .A0(n688), .A1(int_tlv_counter[3]), .Z(n116));
Q_AN03 U551 ( .A0(int_tlv_counter[5]), .A1(n116), .A2(n115), .Z(n120));
Q_AN03 U552 ( .A0(n2135), .A1(int_tlv_counter[1]), .A2(n682), .Z(n115));
Q_OA21 U553 ( .A0(n111), .A1(n120), .B0(fifo_in_valid), .Z(n109));
Q_ND02 U554 ( .A0(n478), .A1(n526), .Z(n118));
Q_AN02 U555 ( .A0(fifo_in_valid), .A1(int_tlv_counter[5]), .Z(n117));
Q_AN03 U556 ( .A0(n117), .A1(n116), .A2(n119), .Z(n110));
Q_AN02 U557 ( .A0(n2135), .A1(n118), .Z(n119));
Q_INV U558 ( .A(n120), .Z(n112));
Q_AN02 U559 ( .A0(n112), .A1(n127), .Z(n121));
Q_AN02 U560 ( .A0(n112), .A1(n129), .Z(n122));
Q_AN02 U561 ( .A0(n112), .A1(n131), .Z(n123));
Q_AN02 U562 ( .A0(n112), .A1(n133), .Z(n124));
Q_AN02 U563 ( .A0(n112), .A1(n134), .Z(n125));
Q_NR02 U564 ( .A0(n120), .A1(int_tlv_counter[0]), .Z(n126));
Q_XOR2 U565 ( .A0(int_tlv_counter[5]), .A1(n128), .Z(n127));
Q_AD01HF U566 ( .A0(int_tlv_counter[4]), .B0(n130), .S(n129), .CO(n128));
Q_AD01HF U567 ( .A0(int_tlv_counter[3]), .B0(n132), .S(n131), .CO(n130));
Q_AD01HF U568 ( .A0(int_tlv_counter[2]), .B0(n46), .S(n133), .CO(n132));
Q_OR02 U569 ( .A0(tlv_counter[0]), .A1(tlv_counter[2]), .Z(n415));
Q_OR02 U570 ( .A0(tlv_counter[3]), .A1(n534), .Z(n466));
Q_OR03 U571 ( .A0(n466), .A1(n415), .A2(tlv_counter[4]), .Z(n618));
Q_OR02 U572 ( .A0(n621), .A1(key_blob_region), .Z(n544));
Q_INV U573 ( .A(stitcher_rd), .Z(n621));
Q_OR02 U574 ( .A0(n544), .A1(n618), .Z(n631));
Q_INV U575 ( .A(n631), .Z(n168));
Q_INV U576 ( .A(n144), .Z(n704));
Q_OR02 U577 ( .A0(n1748), .A1(tlv_counter[2]), .Z(n465));
Q_OA21 U578 ( .A0(tlv_counter[1]), .A1(n465), .B0(tlv_counter[3]), .Z(n540));
Q_MX02 U579 ( .S(tlv_counter[2]), .A0(n2052), .A1(n2034), .Z(n217));
Q_OR02 U580 ( .A0(n444), .A1(tlv_counter[0]), .Z(n532));
Q_AN02 U581 ( .A0(n211), .A1(n532), .Z(n178));
Q_AO21 U582 ( .A0(n178), .A1(tlv_counter[1]), .B0(n218), .Z(n179));
Q_AN02 U583 ( .A0(tlv_counter[2]), .A1(n2042), .Z(n531));
Q_AN03 U584 ( .A0(tlv_counter[0]), .A1(n531), .A2(n534), .Z(n218));
Q_NR02 U585 ( .A0(n179), .A1(tlv_counter[3]), .Z(n180));
Q_OR03 U586 ( .A0(n540), .A1(n180), .A2(tlv_counter[4]), .Z(n181));
Q_OR02 U587 ( .A0(n544), .A1(n181), .Z(n554));
Q_INV U588 ( .A(n181), .Z(n182));
Q_OR02 U589 ( .A0(n182), .A1(key_blob_region), .Z(n183));
Q_AN03 U590 ( .A0(n606), .A1(n183), .A2(stitcher_rd), .Z(n186));
Q_INV U591 ( .A(n186), .Z(n184));
Q_MX02 U592 ( .S(n487), .A0(n184), .A1(n554), .Z(n185));
Q_INV U593 ( .A(n554), .Z(n553));
Q_MX02 U594 ( .S(n732), .A0(n553), .A1(n186), .Z(n187));
Q_INV U595 ( .A(n187), .Z(n188));
Q_MX02 U596 ( .S(aux_key_type[3]), .A0(n188), .A1(n185), .Z(n189));
Q_AN02 U597 ( .A0(n31), .A1(n189), .Z(n190));
Q_INV U598 ( .A(n190), .Z(fifo_in_valid));
Q_OR02 U599 ( .A0(tlv_counter[1]), .A1(n415), .Z(n545));
Q_OR03 U600 ( .A0(tlv_counter[3]), .A1(n1724), .A2(n541), .Z(n191));
Q_OR03 U601 ( .A0(n191), .A1(n545), .A2(n621), .Z(n146));
Q_INV U602 ( .A(n146), .Z(n148));
Q_NR02 U603 ( .A0(n530), .A1(n148), .Z(n192));
Q_AN02 U604 ( .A0(n26), .A1(n146), .Z(n147));
Q_OR02 U605 ( .A0(tlv_counter[2]), .A1(n1722), .Z(n195));
Q_AN02 U606 ( .A0(n195), .A1(tlv_counter[0]), .Z(n193));
Q_OR03 U607 ( .A0(n193), .A1(n203), .A2(tlv_counter[1]), .Z(n194));
Q_OR02 U608 ( .A0(n453), .A1(n195), .Z(n197));
Q_MX02 U609 ( .S(n1724), .A0(n194), .A1(n197), .Z(n196));
Q_OR02 U610 ( .A0(n546), .A1(n196), .Z(n149));
Q_NR02 U611 ( .A0(n546), .A1(n197), .Z(n198));
Q_AN02 U612 ( .A0(tlv_type[0]), .A1(stitcher_out[4]), .Z(n200));
Q_ND02 U613 ( .A0(n136), .A1(n200), .Z(n199));
Q_OR03 U614 ( .A0(n209), .A1(n199), .A2(n546), .Z(n150));
Q_INV U615 ( .A(n200), .Z(n201));
Q_OR03 U616 ( .A0(n1721), .A1(tlv_type[1]), .A2(n201), .Z(n202));
Q_OA21 U617 ( .A0(n208), .A1(n202), .B0(tlv_counter[0]), .Z(n204));
Q_INV U618 ( .A(n532), .Z(n203));
Q_OR03 U619 ( .A0(n204), .A1(n203), .A2(n451), .Z(n205));
Q_OR03 U620 ( .A0(n543), .A1(n415), .A2(n544), .Z(n169));
Q_OR03 U621 ( .A0(n137), .A1(disable_debug_cmd_q), .A2(n465), .Z(n206));
Q_NR03 U622 ( .A0(n450), .A1(n206), .A2(n621), .Z(n207));
Q_OR02 U623 ( .A0(tlv_counter[2]), .A1(n137), .Z(n208));
Q_OR02 U624 ( .A0(n453), .A1(n208), .Z(n209));
Q_OR02 U625 ( .A0(n546), .A1(n209), .Z(n151));
Q_OR02 U626 ( .A0(tlv_counter[1]), .A1(tlv_counter[2]), .Z(n210));
Q_OR02 U627 ( .A0(n1748), .A1(n217), .Z(n211));
Q_AN02 U628 ( .A0(n533), .A1(n415), .Z(n212));
Q_MX02 U629 ( .S(tlv_counter[1]), .A0(n212), .A1(n211), .Z(n213));
Q_INV U630 ( .A(n213), .Z(n214));
Q_MX02 U631 ( .S(tlv_counter[3]), .A0(n214), .A1(n210), .Z(n215));
Q_OR02 U632 ( .A0(tlv_counter[4]), .A1(n215), .Z(n216));
Q_AN03 U633 ( .A0(tlv_counter[0]), .A1(n217), .A2(tlv_counter[1]), .Z(n536));
Q_NR03 U634 ( .A0(n536), .A1(n218), .A2(tlv_counter[3]), .Z(n219));
Q_OR03 U635 ( .A0(n540), .A1(n219), .A2(tlv_counter[4]), .Z(n427));
Q_MX02 U636 ( .S(n2139), .A0(n216), .A1(n427), .Z(n220));
Q_OR02 U637 ( .A0(n544), .A1(n220), .Z(n239));
Q_NR02 U638 ( .A0(n1728), .A1(n2139), .Z(n572));
Q_INV U639 ( .A(n220), .Z(n229));
Q_AN03 U640 ( .A0(n575), .A1(n230), .A2(stitcher_rd), .Z(n244));
Q_INV U641 ( .A(n244), .Z(n242));
Q_OR02 U642 ( .A0(n242), .A1(aux_key_type[1]), .Z(n221));
Q_AN03 U643 ( .A0(n241), .A1(n221), .A2(aux_key_type[2]), .Z(n223));
Q_NR02 U644 ( .A0(n244), .A1(aux_key_type[2]), .Z(n222));
Q_OR02 U645 ( .A0(n223), .A1(n222), .Z(n224));
Q_OR02 U646 ( .A0(n244), .A1(n1960), .Z(n227));
Q_AN02 U647 ( .A0(n244), .A1(aux_key_type[1]), .Z(n225));
Q_OR03 U648 ( .A0(n225), .A1(n437), .A2(aux_key_type[2]), .Z(n226));
Q_ND02 U649 ( .A0(n227), .A1(n226), .Z(n228));
Q_MX02 U650 ( .S(aux_key_type[3]), .A0(n228), .A1(n224), .Z(n266));
Q_OR02 U651 ( .A0(n229), .A1(key_blob_region), .Z(n230));
Q_AN03 U652 ( .A0(n606), .A1(n230), .A2(stitcher_rd), .Z(n436));
Q_INV U653 ( .A(n436), .Z(n254));
Q_OR02 U654 ( .A0(n223), .A1(n255), .Z(n231));
Q_OA21 U655 ( .A0(n231), .A1(n2071), .B0(n257), .Z(n235));
Q_MX02 U656 ( .S(aux_key_type[0]), .A0(n244), .A1(n436), .Z(n246));
Q_AN02 U657 ( .A0(n246), .A1(aux_key_type[1]), .Z(n232));
Q_OR03 U658 ( .A0(n232), .A1(n44), .A2(n1960), .Z(n233));
Q_ND02 U659 ( .A0(n233), .A1(n226), .Z(n234));
Q_AO21 U660 ( .A0(n235), .A1(n682), .B0(n259), .Z(n236));
Q_OA21 U661 ( .A0(n236), .A1(n2136), .B0(n261), .Z(n237));
Q_MX02 U662 ( .S(n23), .A0(n237), .A1(n266), .Z(n238));
Q_OR02 U663 ( .A0(n239), .A1(n1972), .Z(n241));
Q_OR02 U664 ( .A0(n254), .A1(aux_key_type[1]), .Z(n240));
Q_AN03 U665 ( .A0(n241), .A1(n240), .A2(aux_key_type[2]), .Z(n256));
Q_OR02 U666 ( .A0(n256), .A1(n222), .Z(n243));
Q_MX02 U667 ( .S(aux_key_type[0]), .A0(n436), .A1(n244), .Z(n245));
Q_MX02 U668 ( .S(aux_key_type[1]), .A0(n246), .A1(n245), .Z(n247));
Q_OR02 U669 ( .A0(n247), .A1(n1960), .Z(n248));
Q_ND02 U670 ( .A0(n248), .A1(n226), .Z(n249));
Q_MX02 U671 ( .S(aux_key_type[3]), .A0(n249), .A1(n243), .Z(n250));
Q_MX02 U672 ( .S(int_tlv_counter[0]), .A0(n266), .A1(n250), .Z(n251));
Q_OA21 U673 ( .A0(n251), .A1(n2136), .B0(n261), .Z(n252));
Q_AO21 U674 ( .A0(n252), .A1(int_tlv_counter[2]), .B0(n263), .Z(n253));
Q_AN02 U675 ( .A0(n266), .A1(int_tlv_counter[0]), .Z(n259));
Q_NR02 U676 ( .A0(n436), .A1(aux_key_type[2]), .Z(n255));
Q_OR03 U677 ( .A0(n256), .A1(n255), .A2(n2071), .Z(n441));
Q_OR02 U678 ( .A0(n234), .A1(aux_key_type[3]), .Z(n257));
Q_AN02 U679 ( .A0(n441), .A1(n257), .Z(n258));
Q_AO21 U680 ( .A0(n258), .A1(n682), .B0(n259), .Z(n260));
Q_OA21 U681 ( .A0(n260), .A1(n2136), .B0(n261), .Z(n262));
Q_OR02 U682 ( .A0(n266), .A1(int_tlv_counter[1]), .Z(n261));
Q_AO21 U683 ( .A0(n262), .A1(int_tlv_counter[2]), .B0(n263), .Z(n264));
Q_AN02 U684 ( .A0(n266), .A1(n2135), .Z(n263));
Q_MX02 U685 ( .S(int_tlv_counter[3]), .A0(n264), .A1(n253), .Z(n265));
Q_MX03 U686 ( .S0(int_tlv_counter[4]), .S1(int_tlv_counter[5]), .A0(n266), .A1(n265), .A2(n238), .Z(n267));
Q_INV U687 ( .A(n267), .Z(n152));
Q_OR02 U688 ( .A0(n25), .A1(n152), .Z(n268));
Q_AN02 U689 ( .A0(n445), .A1(n419), .Z(n269));
Q_MX02 U690 ( .S(tlv_counter[3]), .A0(n269), .A1(n545), .Z(n270));
Q_OR03 U691 ( .A0(n2139), .A1(tlv_counter[4]), .A2(n270), .Z(n271));
Q_OR02 U692 ( .A0(n544), .A1(n271), .Z(n297));
Q_AO21 U693 ( .A0(n297), .A1(aux_key_type[2]), .B0(n285), .Z(n274));
Q_INV U694 ( .A(n271), .Z(n272));
Q_OR02 U695 ( .A0(n272), .A1(key_blob_region), .Z(n273));
Q_AN03 U696 ( .A0(n606), .A1(n273), .A2(stitcher_rd), .Z(n275));
Q_INV U697 ( .A(n275), .Z(n284));
Q_OA21 U698 ( .A0(n274), .A1(n2071), .B0(n288), .Z(n278));
Q_INV U699 ( .A(n297), .Z(n276));
Q_MX02 U700 ( .S(n21), .A0(n276), .A1(n275), .Z(n277));
Q_INV U701 ( .A(n277), .Z(n287));
Q_AO21 U702 ( .A0(n278), .A1(n682), .B0(n290), .Z(n279));
Q_OA21 U703 ( .A0(n279), .A1(n2136), .B0(n292), .Z(n280));
Q_MX02 U704 ( .S(int_tlv_counter[2]), .A0(n280), .A1(n297), .Z(n281));
Q_OA21 U705 ( .A0(n281), .A1(int_tlv_counter[3]), .B0(n295), .Z(n282));
Q_OR02 U706 ( .A0(n297), .A1(n697), .Z(n295));
Q_AN02 U707 ( .A0(n297), .A1(int_tlv_counter[0]), .Z(n290));
Q_MX02 U708 ( .S(aux_key_type[1]), .A0(n284), .A1(n297), .Z(n283));
Q_AO21 U709 ( .A0(n283), .A1(aux_key_type[2]), .B0(n285), .Z(n286));
Q_NR02 U710 ( .A0(n275), .A1(aux_key_type[2]), .Z(n285));
Q_OA21 U711 ( .A0(n286), .A1(n2071), .B0(n288), .Z(n289));
Q_OR02 U712 ( .A0(n287), .A1(aux_key_type[3]), .Z(n288));
Q_AO21 U713 ( .A0(n289), .A1(n682), .B0(n290), .Z(n291));
Q_OA21 U714 ( .A0(n291), .A1(n2136), .B0(n292), .Z(n293));
Q_OR02 U715 ( .A0(n297), .A1(int_tlv_counter[1]), .Z(n292));
Q_MX02 U716 ( .S(int_tlv_counter[2]), .A0(n297), .A1(n293), .Z(n294));
Q_OA21 U717 ( .A0(n294), .A1(int_tlv_counter[3]), .B0(n295), .Z(n296));
Q_MX04 U718 ( .S0(int_tlv_counter[4]), .S1(int_tlv_counter[5]), .A0(n297), .A1(n296), .A2(n282), .A3(n297), .Z(n298));
Q_INV U719 ( .A(n298), .Z(n153));
Q_OR02 U720 ( .A0(n165), .A1(n153), .Z(n299));
Q_AN03 U721 ( .A0(key_blob_region), .A1(n138), .A2(stitcher_rd), .Z(n548));
Q_INV U722 ( .A(n548), .Z(n506));
Q_AO21 U723 ( .A0(n304), .A1(aux_key_type[3]), .B0(n492), .Z(n302));
Q_AN02 U724 ( .A0(aux_key_type[0]), .A1(n548), .Z(n507));
Q_AN02 U725 ( .A0(aux_key_type[2]), .A1(aux_key_type[1]), .Z(n487));
Q_AN02 U726 ( .A0(n487), .A1(n507), .Z(n300));
Q_OR02 U727 ( .A0(n493), .A1(n526), .Z(n301));
Q_OR03 U728 ( .A0(int_tlv_counter[4]), .A1(n301), .A2(n302), .Z(n303));
Q_OR02 U729 ( .A0(aux_key_type[1]), .A1(n506), .Z(n490));
Q_OA21 U730 ( .A0(n490), .A1(n1960), .B0(n304), .Z(n547));
Q_OR02 U731 ( .A0(n506), .A1(aux_key_type[2]), .Z(n304));
Q_AO21 U732 ( .A0(n547), .A1(aux_key_type[3]), .B0(n492), .Z(n305));
Q_OR03 U733 ( .A0(n688), .A1(n529), .A2(n305), .Z(n306));
Q_MX02 U734 ( .S(int_tlv_counter[5]), .A0(n306), .A1(n303), .Z(n307));
Q_INV U735 ( .A(n307), .Z(n154));
Q_OR02 U736 ( .A0(n165), .A1(n154), .Z(n308));
Q_OR03 U737 ( .A0(key_blob_region), .A1(n1728), .A2(n621), .Z(n322));
Q_INV U738 ( .A(n323), .Z(n309));
Q_OR02 U739 ( .A0(n2098), .A1(n322), .Z(n315));
Q_MX02 U740 ( .S(aux_key_type[1]), .A0(n315), .A1(n322), .Z(n310));
Q_OR02 U741 ( .A0(n1972), .A1(n322), .Z(n317));
Q_MX04 U742 ( .S0(aux_key_type[2]), .S1(aux_key_type[3]), .A0(n317), .A1(n310), .A2(n322), .A3(n309), .Z(n319));
Q_OA21 U743 ( .A0(n1728), .A1(stitcher_eot), .B0(key_blob_region), .Z(n620));
Q_INV U744 ( .A(n368), .Z(n311));
Q_OR03 U745 ( .A0(n620), .A1(n311), .A2(n621), .Z(n313));
Q_OR02 U746 ( .A0(n487), .A1(n313), .Z(n312));
Q_MX02 U747 ( .S(aux_key_type[0]), .A0(n322), .A1(n313), .Z(n314));
Q_MX02 U748 ( .S(aux_key_type[1]), .A0(n315), .A1(n314), .Z(n316));
Q_MX03 U749 ( .S0(aux_key_type[2]), .S1(aux_key_type[3]), .A0(n317), .A1(n316), .A2(n312), .Z(n318));
Q_MX02 U750 ( .S(n13), .A0(n318), .A1(n319), .Z(n155));
Q_OR02 U751 ( .A0(n138), .A1(key_blob_region), .Z(n368));
Q_AN03 U752 ( .A0(n575), .A1(n368), .A2(stitcher_rd), .Z(n373));
Q_INV U753 ( .A(n373), .Z(n339));
Q_OR02 U754 ( .A0(aux_key_type[1]), .A1(n339), .Z(n355));
Q_OR02 U755 ( .A0(n327), .A1(n340), .Z(n320));
Q_AN03 U756 ( .A0(stitcher_rd), .A1(key_blob_region), .A2(n572), .Z(n486));
Q_AN02 U757 ( .A0(n342), .A1(n378), .Z(n380));
Q_AN02 U758 ( .A0(n380), .A1(aux_key_type[1]), .Z(n321));
Q_OA21 U759 ( .A0(n486), .A1(n2098), .B0(n344), .Z(n359));
Q_OR03 U760 ( .A0(n321), .A1(n330), .A2(n1960), .Z(n324));
Q_INV U761 ( .A(n322), .Z(n360));
Q_NR02 U762 ( .A0(n322), .A1(aux_key_type[1]), .Z(n323));
Q_OR03 U763 ( .A0(n474), .A1(n323), .A2(aux_key_type[2]), .Z(n347));
Q_ND02 U764 ( .A0(n324), .A1(n347), .Z(n325));
Q_MX02 U765 ( .S(aux_key_type[3]), .A0(n325), .A1(n320), .Z(n354));
Q_AN02 U766 ( .A0(n355), .A1(aux_key_type[2]), .Z(n327));
Q_AN02 U767 ( .A0(stitcher_rd), .A1(n138), .Z(n372));
Q_INV U768 ( .A(n372), .Z(n337));
Q_NR02 U769 ( .A0(n372), .A1(aux_key_type[2]), .Z(n326));
Q_OR02 U770 ( .A0(n327), .A1(n326), .Z(n328));
Q_OR02 U771 ( .A0(n372), .A1(n2098), .Z(n329));
Q_AN03 U772 ( .A0(n329), .A1(n378), .A2(aux_key_type[1]), .Z(n331));
Q_AN02 U773 ( .A0(n359), .A1(n1972), .Z(n330));
Q_OR03 U774 ( .A0(n331), .A1(n330), .A2(n1960), .Z(n332));
Q_ND02 U775 ( .A0(n332), .A1(n347), .Z(n333));
Q_MX03 U776 ( .S0(aux_key_type[3]), .S1(int_tlv_counter[0]), .A0(n333), .A1(n328), .A2(n354), .Z(n334));
Q_OA21 U777 ( .A0(n334), .A1(n2136), .B0(n352), .Z(n335));
Q_MX02 U778 ( .S(n23), .A0(n335), .A1(n354), .Z(n336));
Q_OR02 U779 ( .A0(aux_key_type[1]), .A1(n337), .Z(n338));
Q_AO21 U780 ( .A0(n338), .A1(aux_key_type[2]), .B0(n340), .Z(n341));
Q_NR02 U781 ( .A0(n373), .A1(aux_key_type[2]), .Z(n340));
Q_OR02 U782 ( .A0(n373), .A1(n2098), .Z(n342));
Q_OA21 U783 ( .A0(n548), .A1(aux_key_type[0]), .B0(n342), .Z(n343));
Q_OA21 U784 ( .A0(n548), .A1(n2098), .B0(n344), .Z(n345));
Q_OR02 U785 ( .A0(n373), .A1(aux_key_type[0]), .Z(n344));
Q_MX02 U786 ( .S(aux_key_type[1]), .A0(n345), .A1(n343), .Z(n346));
Q_OR02 U787 ( .A0(n346), .A1(n1960), .Z(n348));
Q_ND02 U788 ( .A0(n348), .A1(n347), .Z(n349));
Q_MX02 U789 ( .S(aux_key_type[3]), .A0(n349), .A1(n341), .Z(n350));
Q_MX02 U790 ( .S(int_tlv_counter[0]), .A0(n354), .A1(n350), .Z(n351));
Q_OA21 U791 ( .A0(n351), .A1(n2136), .B0(n352), .Z(n353));
Q_OR02 U792 ( .A0(n354), .A1(int_tlv_counter[1]), .Z(n352));
Q_MX03 U793 ( .S0(n11), .S1(int_tlv_counter[5]), .A0(n354), .A1(n353), .A2(n336), .Z(n156));
Q_MX02 U794 ( .S(aux_key_type[1]), .A0(n359), .A1(n373), .Z(n356));
Q_INV U795 ( .A(n356), .Z(n357));
Q_MX02 U796 ( .S(aux_key_type[2]), .A0(n357), .A1(n355), .Z(n358));
Q_MX02 U797 ( .S(aux_key_type[1]), .A0(n360), .A1(n359), .Z(n382));
Q_MX02 U798 ( .S(aux_key_type[2]), .A0(n382), .A1(n380), .Z(n361));
Q_INV U799 ( .A(n361), .Z(n362));
Q_MX02 U800 ( .S(aux_key_type[3]), .A0(n362), .A1(n358), .Z(n386));
Q_ND02 U801 ( .A0(n2139), .A1(n1947), .Z(n363));
Q_AO21 U802 ( .A0(n138), .A1(n363), .B0(n617), .Z(n364));
Q_ND03 U803 ( .A0(n364), .A1(n368), .A2(stitcher_rd), .Z(n365));
Q_OR02 U804 ( .A0(aux_key_type[1]), .A1(n365), .Z(n366));
Q_ND02 U805 ( .A0(n2139), .A1(n1970), .Z(n367));
Q_AO21 U806 ( .A0(n138), .A1(n367), .B0(n617), .Z(n369));
Q_AN03 U807 ( .A0(n369), .A1(n368), .A2(stitcher_rd), .Z(n370));
Q_MX02 U808 ( .S(n1992), .A0(n486), .A1(n548), .Z(n371));
Q_MX02 U809 ( .S(n1992), .A0(n373), .A1(n372), .Z(n377));
Q_MX03 U810 ( .S0(aux_key_type[0]), .S1(aux_key_type[1]), .A0(n377), .A1(n371), .A2(n370), .Z(n374));
Q_INV U811 ( .A(n374), .Z(n375));
Q_MX02 U812 ( .S(aux_key_type[2]), .A0(n375), .A1(n366), .Z(n376));
Q_OA21 U813 ( .A0(n377), .A1(n2098), .B0(n378), .Z(n379));
Q_OR02 U814 ( .A0(n486), .A1(aux_key_type[0]), .Z(n378));
Q_MX02 U815 ( .S(aux_key_type[1]), .A0(n380), .A1(n379), .Z(n381));
Q_MX02 U816 ( .S(aux_key_type[2]), .A0(n382), .A1(n381), .Z(n383));
Q_INV U817 ( .A(n383), .Z(n384));
Q_MX03 U818 ( .S0(aux_key_type[3]), .S1(int_tlv_counter[0]), .A0(n384), .A1(n376), .A2(n386), .Z(n385));
Q_MX02 U819 ( .S(n4), .A0(n385), .A1(n386), .Z(n387));
Q_INV U820 ( .A(n387), .Z(n157));
Q_OR02 U821 ( .A0(n2044), .A1(tlv_type[2]), .Z(n405));
Q_OR02 U822 ( .A0(n1720), .A1(n405), .Z(n459));
Q_OR02 U823 ( .A0(tlv_type[1]), .A1(n459), .Z(n392));
Q_OR02 U824 ( .A0(n465), .A1(n392), .Z(n389));
Q_NR02 U825 ( .A0(n412), .A1(n389), .Z(n388));
Q_AN02 U826 ( .A0(n389), .A1(tlv_counter[1]), .Z(n390));
Q_OR03 U827 ( .A0(n390), .A1(n416), .A2(n546), .Z(n158));
Q_NR02 U828 ( .A0(n461), .A1(n392), .Z(n391));
Q_AN02 U829 ( .A0(tlv_counter[2]), .A1(n392), .Z(n394));
Q_OR02 U830 ( .A0(n543), .A1(n424), .Z(n393));
Q_OR03 U831 ( .A0(n544), .A1(n393), .A2(n394), .Z(n159));
Q_AN02 U832 ( .A0(tlv_counter[2]), .A1(n135), .Z(n399));
Q_ND02 U833 ( .A0(tlv_counter[0]), .A1(n399), .Z(n395));
Q_NR03 U834 ( .A0(n450), .A1(n395), .A2(n621), .Z(n396));
Q_OR02 U835 ( .A0(n399), .A1(n1748), .Z(n397));
Q_ND02 U836 ( .A0(n397), .A1(n532), .Z(n398));
Q_OR02 U837 ( .A0(n451), .A1(n398), .Z(n160));
Q_INV U838 ( .A(n399), .Z(n400));
Q_OR02 U839 ( .A0(tlv_counter[0]), .A1(n400), .Z(n402));
Q_NR03 U840 ( .A0(n411), .A1(n402), .A2(n621), .Z(n401));
Q_AN02 U841 ( .A0(n402), .A1(tlv_counter[1]), .Z(n403));
Q_OR03 U842 ( .A0(n403), .A1(n416), .A2(n546), .Z(n161));
Q_OR02 U843 ( .A0(tlv_type[5]), .A1(n2057), .Z(n404));
Q_OR03 U844 ( .A0(tlv_type[7]), .A1(tlv_type[6]), .A2(n404), .Z(n406));
Q_OR03 U845 ( .A0(n457), .A1(n405), .A2(n406), .Z(n418));
Q_OR02 U846 ( .A0(tlv_type[3]), .A1(n2058), .Z(n407));
Q_OR02 U847 ( .A0(n2059), .A1(n1720), .Z(n408));
Q_OR03 U848 ( .A0(n408), .A1(n407), .A2(n409), .Z(n422));
Q_MX02 U849 ( .S(tlv_counter[2]), .A0(n422), .A1(n418), .Z(n410));
Q_OR02 U850 ( .A0(n1748), .A1(n410), .Z(n414));
Q_OR02 U851 ( .A0(n541), .A1(n466), .Z(n411));
Q_OR02 U852 ( .A0(n621), .A1(n411), .Z(n412));
Q_NR02 U853 ( .A0(n412), .A1(n414), .Z(n413));
Q_AN02 U854 ( .A0(n414), .A1(tlv_counter[1]), .Z(n417));
Q_AN02 U855 ( .A0(n415), .A1(n534), .Z(n416));
Q_OR03 U856 ( .A0(n417), .A1(n416), .A2(n546), .Z(n162));
Q_OA21 U857 ( .A0(n545), .A1(n418), .B0(tlv_counter[3]), .Z(n426));
Q_OR02 U858 ( .A0(tlv_counter[1]), .A1(n532), .Z(n419));
Q_OA21 U859 ( .A0(n419), .A1(n422), .B0(n538), .Z(n420));
Q_NR03 U860 ( .A0(n426), .A1(n420), .A2(n542), .Z(n421));
Q_AN02 U861 ( .A0(tlv_counter[2]), .A1(n422), .Z(n423));
Q_OR02 U862 ( .A0(tlv_counter[1]), .A1(tlv_counter[0]), .Z(n424));
Q_OA21 U863 ( .A0(n424), .A1(n423), .B0(n538), .Z(n425));
Q_OR03 U864 ( .A0(n426), .A1(n425), .A2(n542), .Z(n163));
Q_OR02 U865 ( .A0(n544), .A1(n427), .Z(n591));
Q_INV U866 ( .A(n427), .Z(n573));
Q_AN03 U867 ( .A0(n606), .A1(n574), .A2(stitcher_rd), .Z(n677));
Q_INV U868 ( .A(n677), .Z(n429));
Q_OR02 U869 ( .A0(n429), .A1(aux_key_type[1]), .Z(n428));
Q_AN03 U870 ( .A0(n592), .A1(n428), .A2(aux_key_type[2]), .Z(n576));
Q_NR02 U871 ( .A0(n677), .A1(aux_key_type[2]), .Z(n430));
Q_OR03 U872 ( .A0(n576), .A1(n430), .A2(n2071), .Z(n571));
Q_AO21 U873 ( .A0(n677), .A1(aux_key_type[1]), .B0(n580), .Z(n431));
Q_INV U874 ( .A(n591), .Z(n166));
Q_MX02 U875 ( .S(aux_key_type[2]), .A0(n431), .A1(n677), .Z(n432));
Q_INV U876 ( .A(n432), .Z(n433));
Q_OR02 U877 ( .A0(n433), .A1(aux_key_type[3]), .Z(n434));
Q_ND02 U878 ( .A0(n571), .A1(n434), .Z(n435));
Q_AO21 U879 ( .A0(n436), .A1(aux_key_type[1]), .B0(n437), .Z(n438));
Q_NR02 U880 ( .A0(n239), .A1(aux_key_type[1]), .Z(n437));
Q_MX02 U881 ( .S(aux_key_type[2]), .A0(n438), .A1(n436), .Z(n439));
Q_INV U882 ( .A(n439), .Z(n440));
Q_OA21 U883 ( .A0(n440), .A1(aux_key_type[3]), .B0(n441), .Z(n164));
Q_AN03 U884 ( .A0(tlv_type[0]), .A1(n135), .A2(tlv_counter[2]), .Z(n448));
Q_INV U885 ( .A(n448), .Z(n442));
Q_NR03 U886 ( .A0(n446), .A1(n442), .A2(n544), .Z(n443));
Q_OR03 U887 ( .A0(tlv_type[0]), .A1(n1719), .A2(n444), .Z(n454));
Q_OR02 U888 ( .A0(n534), .A1(tlv_counter[0]), .Z(n445));
Q_OR02 U889 ( .A0(n543), .A1(n445), .Z(n446));
Q_NR03 U890 ( .A0(n446), .A1(n454), .A2(n544), .Z(n447));
Q_ND02 U891 ( .A0(tlv_counter[0]), .A1(n448), .Z(n449));
Q_OR02 U892 ( .A0(n541), .A1(n460), .Z(n450));
Q_OR02 U893 ( .A0(n621), .A1(n450), .Z(n451));
Q_NR02 U894 ( .A0(n451), .A1(n449), .Z(n452));
Q_OR02 U895 ( .A0(tlv_counter[1]), .A1(n1748), .Z(n453));
Q_OR02 U896 ( .A0(n543), .A1(n453), .Z(n455));
Q_NR03 U897 ( .A0(n455), .A1(n454), .A2(n544), .Z(n456));
Q_OR02 U898 ( .A0(tlv_type[1]), .A1(n2059), .Z(n457));
Q_OR02 U899 ( .A0(n457), .A1(n459), .Z(n463));
Q_NR02 U900 ( .A0(n461), .A1(n463), .Z(n458));
Q_OR03 U901 ( .A0(tlv_type[1]), .A1(tlv_type[0]), .A2(n459), .Z(n467));
Q_OR03 U902 ( .A0(n460), .A1(n532), .A2(n542), .Z(n461));
Q_OR02 U903 ( .A0(tlv_counter[3]), .A1(tlv_counter[1]), .Z(n460));
Q_NR02 U904 ( .A0(n461), .A1(n467), .Z(n462));
Q_NR02 U905 ( .A0(n468), .A1(n463), .Z(n464));
Q_OR03 U906 ( .A0(n466), .A1(n465), .A2(n542), .Z(n468));
Q_NR02 U907 ( .A0(n468), .A1(n467), .Z(n469));
Q_INV U908 ( .A(n486), .Z(n501));
Q_OR02 U909 ( .A0(aux_key_type[1]), .A1(n501), .Z(n484));
Q_NR02 U910 ( .A0(n471), .A1(n484), .Z(n470));
Q_ND02 U911 ( .A0(aux_key_type[3]), .A1(aux_key_type[2]), .Z(n471));
Q_OR02 U912 ( .A0(n471), .A1(n490), .Z(n473));
Q_NR03 U913 ( .A0(n514), .A1(n529), .A2(n473), .Z(n472));
Q_AN02 U914 ( .A0(aux_key_type[1]), .A1(n486), .Z(n474));
Q_INV U915 ( .A(n474), .Z(n519));
Q_NR02 U916 ( .A0(n476), .A1(n519), .Z(n475));
Q_AN02 U917 ( .A0(aux_key_type[1]), .A1(n548), .Z(n549));
Q_INV U918 ( .A(n549), .Z(n523));
Q_OR02 U919 ( .A0(n2071), .A1(aux_key_type[2]), .Z(n476));
Q_OR02 U920 ( .A0(n476), .A1(n523), .Z(n483));
Q_OR02 U921 ( .A0(n526), .A1(n483), .Z(n481));
Q_NR02 U922 ( .A0(n495), .A1(n481), .Z(n477));
Q_OR02 U923 ( .A0(int_tlv_counter[1]), .A1(n682), .Z(n478));
Q_OR02 U924 ( .A0(n493), .A1(n478), .Z(n479));
Q_NR03 U925 ( .A0(n494), .A1(n479), .A2(n483), .Z(n480));
Q_NR02 U926 ( .A0(n498), .A1(n481), .Z(n482));
Q_OR02 U927 ( .A0(aux_key_type[2]), .A1(n484), .Z(n485));
Q_AN02 U928 ( .A0(aux_key_type[0]), .A1(n486), .Z(n502));
Q_ND02 U929 ( .A0(n487), .A1(n502), .Z(n488));
Q_MX02 U930 ( .S(aux_key_type[3]), .A0(n488), .A1(n485), .Z(n489));
Q_OR02 U931 ( .A0(aux_key_type[2]), .A1(n490), .Z(n491));
Q_AO21 U932 ( .A0(n491), .A1(aux_key_type[3]), .B0(n492), .Z(n500));
Q_NR02 U933 ( .A0(n300), .A1(aux_key_type[3]), .Z(n492));
Q_OR02 U934 ( .A0(n526), .A1(n500), .Z(n497));
Q_OR02 U935 ( .A0(int_tlv_counter[3]), .A1(int_tlv_counter[2]), .Z(n493));
Q_OR02 U936 ( .A0(n494), .A1(n493), .Z(n495));
Q_OR02 U937 ( .A0(n706), .A1(int_tlv_counter[4]), .Z(n494));
Q_NR02 U938 ( .A0(n495), .A1(n497), .Z(n496));
Q_OR02 U939 ( .A0(n514), .A1(n527), .Z(n498));
Q_NR02 U940 ( .A0(n498), .A1(n497), .Z(n499));
Q_OR02 U941 ( .A0(aux_key_type[0]), .A1(n501), .Z(n517));
Q_INV U942 ( .A(n502), .Z(n503));
Q_MX02 U943 ( .S(aux_key_type[1]), .A0(n503), .A1(n517), .Z(n504));
Q_NR02 U944 ( .A0(n510), .A1(n504), .Z(n505));
Q_OR02 U945 ( .A0(aux_key_type[0]), .A1(n506), .Z(n522));
Q_INV U946 ( .A(n507), .Z(n508));
Q_MX02 U947 ( .S(aux_key_type[1]), .A0(n508), .A1(n522), .Z(n509));
Q_OR02 U948 ( .A0(aux_key_type[3]), .A1(n1960), .Z(n510));
Q_OR02 U949 ( .A0(n510), .A1(n509), .Z(n516));
Q_ND02 U950 ( .A0(int_tlv_counter[1]), .A1(int_tlv_counter[0]), .Z(n511));
Q_OR02 U951 ( .A0(n512), .A1(n511), .Z(n513));
Q_ND02 U952 ( .A0(int_tlv_counter[3]), .A1(int_tlv_counter[2]), .Z(n512));
Q_NR03 U953 ( .A0(n514), .A1(n513), .A2(n516), .Z(n515));
Q_OR02 U954 ( .A0(int_tlv_counter[5]), .A1(n688), .Z(n514));
Q_OR02 U955 ( .A0(aux_key_type[1]), .A1(n517), .Z(n518));
Q_MX02 U956 ( .S(aux_key_type[2]), .A0(n519), .A1(n518), .Z(n520));
Q_NR02 U957 ( .A0(aux_key_type[3]), .A1(n520), .Z(n521));
Q_OA21 U958 ( .A0(aux_key_type[1]), .A1(n522), .B0(aux_key_type[2]), .Z(n524));
Q_NR03 U959 ( .A0(n524), .A1(n43), .A2(aux_key_type[3]), .Z(n525));
Q_OR02 U960 ( .A0(n2136), .A1(int_tlv_counter[0]), .Z(n526));
Q_OR02 U961 ( .A0(int_tlv_counter[3]), .A1(n2135), .Z(n527));
Q_OR02 U962 ( .A0(n527), .A1(n526), .Z(n529));
Q_OR02 U963 ( .A0(int_tlv_counter[5]), .A1(int_tlv_counter[4]), .Z(n528));
Q_OR03 U964 ( .A0(n704), .A1(n528), .A2(n529), .Z(n530));
Q_AN02 U965 ( .A0(n144), .A1(skip[5]), .Z(n165));
Q_OR02 U966 ( .A0(n531), .A1(n1748), .Z(n533));
Q_AN02 U967 ( .A0(n533), .A1(n532), .Z(n535));
Q_AO21 U968 ( .A0(n535), .A1(n534), .B0(n536), .Z(n537));
Q_NR02 U969 ( .A0(n537), .A1(tlv_counter[3]), .Z(n539));
Q_OR03 U970 ( .A0(n540), .A1(n539), .A2(n542), .Z(n167));
Q_OR02 U971 ( .A0(key_blob_region), .A1(tlv_counter[4]), .Z(n541));
Q_OR02 U972 ( .A0(n621), .A1(n541), .Z(n542));
Q_OR02 U973 ( .A0(tlv_counter[4]), .A1(tlv_counter[3]), .Z(n543));
Q_OR02 U974 ( .A0(n544), .A1(n543), .Z(n546));
Q_OR02 U975 ( .A0(n546), .A1(n545), .Z(n170));
Q_OR02 U976 ( .A0(n548), .A1(n1960), .Z(n551));
Q_OR02 U977 ( .A0(n549), .A1(aux_key_type[2]), .Z(n550));
Q_ND02 U978 ( .A0(n551), .A1(n550), .Z(n552));
Q_MX02 U979 ( .S(aux_key_type[3]), .A0(n552), .A1(n547), .Z(n565));
Q_MX02 U980 ( .S(int_tlv_counter[1]), .A0(n553), .A1(n565), .Z(n558));
Q_INV U981 ( .A(n565), .Z(n561));
Q_MX02 U982 ( .S(int_tlv_counter[1]), .A0(n561), .A1(n554), .Z(n560));
Q_INV U983 ( .A(n560), .Z(n555));
Q_MX03 U984 ( .S0(int_tlv_counter[2]), .S1(int_tlv_counter[3]), .A0(n555), .A1(n558), .A2(n565), .Z(n556));
Q_MX02 U985 ( .S(n2), .A0(n565), .A1(n556), .Z(n557));
Q_MX02 U986 ( .S(int_tlv_counter[2]), .A0(n558), .A1(n565), .Z(n559));
Q_MX02 U987 ( .S(int_tlv_counter[2]), .A0(n561), .A1(n560), .Z(n562));
Q_INV U988 ( .A(n562), .Z(n563));
Q_MX03 U989 ( .S0(int_tlv_counter[3]), .S1(int_tlv_counter[4]), .A0(n563), .A1(n559), .A2(n565), .Z(n564));
Q_MX02 U990 ( .S(n1), .A0(n565), .A1(n564), .Z(n566));
Q_INV U991 ( .A(n566), .Z(n171));
Q_OR02 U992 ( .A0(n677), .A1(n2098), .Z(n567));
Q_AN03 U993 ( .A0(n567), .A1(n578), .A2(aux_key_type[1]), .Z(n568));
Q_OR03 U994 ( .A0(n568), .A1(n580), .A2(n1960), .Z(n569));
Q_ND02 U995 ( .A0(n569), .A1(n582), .Z(n570));
Q_OA21 U996 ( .A0(n570), .A1(aux_key_type[3]), .B0(n571), .Z(n612));
Q_OR02 U997 ( .A0(n572), .A1(n617), .Z(n575));
Q_OR02 U998 ( .A0(n573), .A1(key_blob_region), .Z(n574));
Q_AN03 U999 ( .A0(n575), .A1(n574), .A2(stitcher_rd), .Z(n678));
Q_INV U1000 ( .A(n678), .Z(n593));
Q_OR02 U1001 ( .A0(n576), .A1(n594), .Z(n577));
Q_OA21 U1002 ( .A0(n577), .A1(n2071), .B0(n596), .Z(n585));
Q_OR02 U1003 ( .A0(n678), .A1(n2098), .Z(n579));
Q_OR02 U1004 ( .A0(n166), .A1(aux_key_type[0]), .Z(n578));
Q_AN03 U1005 ( .A0(n579), .A1(n578), .A2(aux_key_type[1]), .Z(n581));
Q_NR02 U1006 ( .A0(n591), .A1(aux_key_type[1]), .Z(n580));
Q_OR03 U1007 ( .A0(n581), .A1(n580), .A2(n1960), .Z(n583));
Q_OR02 U1008 ( .A0(n166), .A1(aux_key_type[2]), .Z(n582));
Q_ND02 U1009 ( .A0(n583), .A1(n582), .Z(n584));
Q_AO21 U1010 ( .A0(n585), .A1(n682), .B0(n597), .Z(n586));
Q_OA21 U1011 ( .A0(n586), .A1(n2136), .B0(n599), .Z(n587));
Q_AO21 U1012 ( .A0(n587), .A1(n2135), .B0(n610), .Z(n588));
Q_OA21 U1013 ( .A0(n588), .A1(int_tlv_counter[3]), .B0(n602), .Z(n589));
Q_MX02 U1014 ( .S(int_tlv_counter[4]), .A0(n589), .A1(n612), .Z(n590));
Q_OR02 U1015 ( .A0(n612), .A1(n697), .Z(n602));
Q_AN02 U1016 ( .A0(n612), .A1(int_tlv_counter[0]), .Z(n597));
Q_OR02 U1017 ( .A0(n591), .A1(n1972), .Z(n592));
Q_OA21 U1018 ( .A0(n593), .A1(aux_key_type[1]), .B0(n592), .Z(n676));
Q_AO21 U1019 ( .A0(n676), .A1(aux_key_type[2]), .B0(n594), .Z(n595));
Q_NR02 U1020 ( .A0(n678), .A1(aux_key_type[2]), .Z(n594));
Q_OA21 U1021 ( .A0(n595), .A1(n2071), .B0(n596), .Z(n708));
Q_OR02 U1022 ( .A0(n584), .A1(aux_key_type[3]), .Z(n596));
Q_AO21 U1023 ( .A0(n708), .A1(n682), .B0(n597), .Z(n598));
Q_OA21 U1024 ( .A0(n598), .A1(n2136), .B0(n599), .Z(n600));
Q_OR02 U1025 ( .A0(n612), .A1(int_tlv_counter[1]), .Z(n599));
Q_AO21 U1026 ( .A0(n600), .A1(int_tlv_counter[2]), .B0(n613), .Z(n601));
Q_OA21 U1027 ( .A0(n601), .A1(int_tlv_counter[3]), .B0(n602), .Z(n603));
Q_AN02 U1028 ( .A0(n612), .A1(int_tlv_counter[2]), .Z(n610));
Q_OA21 U1029 ( .A0(n612), .A1(n2136), .B0(n34), .Z(n641));
Q_ND02 U1030 ( .A0(n1728), .A1(key_blob_region), .Z(n606));
Q_INV U1031 ( .A(n618), .Z(n604));
Q_OR02 U1032 ( .A0(n604), .A1(key_blob_region), .Z(n605));
Q_AN03 U1033 ( .A0(n606), .A1(n605), .A2(stitcher_rd), .Z(n608));
Q_INV U1034 ( .A(n608), .Z(n623));
Q_MX02 U1035 ( .S(n22), .A0(n623), .A1(n631), .Z(n607));
Q_MX02 U1036 ( .S(aux_key_type[1]), .A0(n168), .A1(n608), .Z(n609));
Q_INV U1037 ( .A(n609), .Z(n625));
Q_MX03 U1038 ( .S0(aux_key_type[2]), .S1(aux_key_type[3]), .A0(n625), .A1(n607), .A2(n631), .Z(n650));
Q_AO21 U1039 ( .A0(n641), .A1(n2135), .B0(n610), .Z(n611));
Q_AO21 U1040 ( .A0(n641), .A1(int_tlv_counter[2]), .B0(n613), .Z(n614));
Q_AN02 U1041 ( .A0(n612), .A1(n2135), .Z(n613));
Q_MX03 U1042 ( .S0(int_tlv_counter[3]), .S1(int_tlv_counter[4]), .A0(n614), .A1(n611), .A2(n603), .Z(n615));
Q_MX02 U1043 ( .S(int_tlv_counter[5]), .A0(n615), .A1(n590), .Z(n616));
Q_OA21 U1044 ( .A0(n631), .A1(n1960), .B0(n633), .Z(n622));
Q_AN02 U1045 ( .A0(n618), .A1(n617), .Z(n619));
Q_OR03 U1046 ( .A0(n620), .A1(n619), .A2(n621), .Z(n632));
Q_AO21 U1047 ( .A0(n622), .A1(aux_key_type[3]), .B0(n635), .Z(n626));
Q_MX02 U1048 ( .S(n22), .A0(n623), .A1(n632), .Z(n624));
Q_MX02 U1049 ( .S(aux_key_type[2]), .A0(n625), .A1(n624), .Z(n654));
Q_OA21 U1050 ( .A0(n626), .A1(int_tlv_counter[0]), .B0(n636), .Z(n627));
Q_AO21 U1051 ( .A0(n627), .A1(int_tlv_counter[1]), .B0(n638), .Z(n628));
Q_MX02 U1052 ( .S(int_tlv_counter[2]), .A0(n628), .A1(n650), .Z(n629));
Q_AO21 U1053 ( .A0(n629), .A1(n697), .B0(n643), .Z(n630));
Q_MX02 U1054 ( .S(int_tlv_counter[4]), .A0(n630), .A1(n650), .Z(n648));
Q_OR02 U1055 ( .A0(n650), .A1(n682), .Z(n636));
Q_MX02 U1056 ( .S(aux_key_type[1]), .A0(n632), .A1(n631), .Z(n653));
Q_OA21 U1057 ( .A0(n653), .A1(n1960), .B0(n633), .Z(n634));
Q_OR02 U1058 ( .A0(n632), .A1(aux_key_type[2]), .Z(n633));
Q_AO21 U1059 ( .A0(n634), .A1(aux_key_type[3]), .B0(n635), .Z(n661));
Q_AN02 U1060 ( .A0(n654), .A1(n2071), .Z(n635));
Q_OA21 U1061 ( .A0(n661), .A1(int_tlv_counter[0]), .B0(n636), .Z(n637));
Q_AO21 U1062 ( .A0(n637), .A1(int_tlv_counter[1]), .B0(n638), .Z(n639));
Q_AN02 U1063 ( .A0(n650), .A1(n2136), .Z(n638));
Q_MX02 U1064 ( .S(int_tlv_counter[2]), .A0(n650), .A1(n639), .Z(n640));
Q_AO21 U1065 ( .A0(n640), .A1(n697), .B0(n643), .Z(n649));
Q_AN02 U1066 ( .A0(n650), .A1(int_tlv_counter[3]), .Z(n643));
Q_NR02 U1067 ( .A0(n641), .A1(int_tlv_counter[3]), .Z(n642));
Q_OR02 U1068 ( .A0(n643), .A1(n642), .Z(n644));
Q_MX03 U1069 ( .S0(int_tlv_counter[4]), .S1(int_tlv_counter[5]), .A0(n644), .A1(n649), .A2(n648), .Z(n645));
Q_INV U1070 ( .A(n645), .Z(n646));
Q_MX02 U1071 ( .S(skip[5]), .A0(n646), .A1(n616), .Z(n647));
Q_MX03 U1072 ( .S0(int_tlv_counter[4]), .S1(int_tlv_counter[5]), .A0(n650), .A1(n649), .A2(n648), .Z(n651));
Q_INV U1073 ( .A(n651), .Z(n652));
Q_MX02 U1074 ( .S(n144), .A0(n652), .A1(n647), .Z(n172));
Q_MX02 U1075 ( .S(aux_key_type[3]), .A0(n654), .A1(n653), .Z(n655));
Q_AO21 U1076 ( .A0(n655), .A1(int_tlv_counter[0]), .B0(n42), .Z(n656));
Q_OA21 U1077 ( .A0(n656), .A1(int_tlv_counter[1]), .B0(n664), .Z(n657));
Q_AO21 U1078 ( .A0(n657), .A1(n2135), .B0(n666), .Z(n658));
Q_MX02 U1079 ( .S(int_tlv_counter[3]), .A0(n658), .A1(n661), .Z(n659));
Q_AO21 U1080 ( .A0(n659), .A1(n688), .B0(n673), .Z(n660));
Q_AN02 U1081 ( .A0(n661), .A1(int_tlv_counter[4]), .Z(n673));
Q_AN02 U1082 ( .A0(n661), .A1(int_tlv_counter[2]), .Z(n666));
Q_OR02 U1083 ( .A0(n661), .A1(n2136), .Z(n664));
Q_OA21 U1084 ( .A0(n708), .A1(n682), .B0(n662), .Z(n693));
Q_INV U1085 ( .A(n661), .Z(n668));
Q_OR02 U1086 ( .A0(n668), .A1(int_tlv_counter[0]), .Z(n662));
Q_INV U1087 ( .A(n693), .Z(n663));
Q_OA21 U1088 ( .A0(n663), .A1(int_tlv_counter[1]), .B0(n664), .Z(n665));
Q_AO21 U1089 ( .A0(n665), .A1(n2135), .B0(n666), .Z(n667));
Q_NR02 U1090 ( .A0(n661), .A1(int_tlv_counter[1]), .Z(n669));
Q_OR03 U1091 ( .A0(n694), .A1(n669), .A2(int_tlv_counter[2]), .Z(n670));
Q_ND02 U1092 ( .A0(n696), .A1(n670), .Z(n671));
Q_MX02 U1093 ( .S(int_tlv_counter[3]), .A0(n671), .A1(n667), .Z(n672));
Q_AO21 U1094 ( .A0(n672), .A1(n688), .B0(n673), .Z(n674));
Q_MX02 U1095 ( .S(int_tlv_counter[5]), .A0(n674), .A1(n660), .Z(n675));
Q_MX02 U1096 ( .S(aux_key_type[1]), .A0(n678), .A1(n677), .Z(n679));
Q_INV U1097 ( .A(n679), .Z(n680));
Q_MX02 U1098 ( .S(aux_key_type[2]), .A0(n680), .A1(n676), .Z(n681));
Q_MX02 U1099 ( .S(aux_key_type[3]), .A0(n584), .A1(n681), .Z(n683));
Q_MX02 U1100 ( .S(int_tlv_counter[0]), .A0(n708), .A1(n683), .Z(n684));
Q_AO21 U1101 ( .A0(n684), .A1(n2136), .B0(n689), .Z(n685));
Q_OA21 U1102 ( .A0(n685), .A1(int_tlv_counter[2]), .B0(n691), .Z(n686));
Q_MX02 U1103 ( .S(int_tlv_counter[3]), .A0(n686), .A1(n708), .Z(n687));
Q_OA21 U1104 ( .A0(n687), .A1(int_tlv_counter[4]), .B0(n700), .Z(n707));
Q_OR02 U1105 ( .A0(n708), .A1(n688), .Z(n700));
Q_OR02 U1106 ( .A0(n708), .A1(n2135), .Z(n691));
Q_AN02 U1107 ( .A0(n708), .A1(int_tlv_counter[1]), .Z(n689));
Q_AO21 U1108 ( .A0(n693), .A1(n2136), .B0(n689), .Z(n690));
Q_OA21 U1109 ( .A0(n690), .A1(int_tlv_counter[2]), .B0(n691), .Z(n692));
Q_OR02 U1110 ( .A0(n693), .A1(n2135), .Z(n696));
Q_AN02 U1111 ( .A0(n693), .A1(int_tlv_counter[1]), .Z(n694));
Q_AO21 U1112 ( .A0(n708), .A1(n2136), .B0(n694), .Z(n695));
Q_OA21 U1113 ( .A0(n695), .A1(int_tlv_counter[2]), .B0(n696), .Z(n698));
Q_MX02 U1114 ( .S(int_tlv_counter[3]), .A0(n698), .A1(n692), .Z(n699));
Q_OA21 U1115 ( .A0(n699), .A1(int_tlv_counter[4]), .B0(n700), .Z(n701));
Q_MX02 U1116 ( .S(int_tlv_counter[5]), .A0(n701), .A1(n707), .Z(n702));
Q_INV U1117 ( .A(n702), .Z(n703));
Q_MX02 U1118 ( .S(skip[5]), .A0(n703), .A1(n675), .Z(n705));
Q_MX02 U1119 ( .S(int_tlv_counter[5]), .A0(n708), .A1(n707), .Z(n709));
Q_INV U1120 ( .A(n709), .Z(n710));
Q_MX02 U1121 ( .S(n144), .A0(n710), .A1(n705), .Z(n173));
Q_INV U1122 ( .A(n140), .Z(n711));
Q_OR03 U1123 ( .A0(stitcher_out[57]), .A1(n711), .A2(n721), .Z(n712));
Q_AN03 U1124 ( .A0(stitcher_out[57]), .A1(n140), .A2(stitcher_out[58]), .Z(n713));
Q_OA21 U1125 ( .A0(n2026), .A1(n140), .B0(n2023), .Z(n714));
Q_MX02 U1126 ( .S(stitcher_out[59]), .A0(n714), .A1(n713), .Z(n715));
Q_INV U1127 ( .A(n715), .Z(n716));
Q_MX02 U1128 ( .S(stitcher_out[60]), .A0(n716), .A1(n712), .Z(n717));
Q_OR02 U1129 ( .A0(n141), .A1(n717), .Z(n174));
Q_ND02 U1130 ( .A0(stitcher_out[57]), .A1(n145), .Z(n718));
Q_OR02 U1131 ( .A0(stitcher_out[59]), .A1(stitcher_out[58]), .Z(n721));
Q_OR03 U1132 ( .A0(n719), .A1(n721), .A2(n141), .Z(n175));
Q_AN02 U1133 ( .A0(stitcher_out[57]), .A1(n1702), .Z(n720));
Q_MX02 U1134 ( .S(stitcher_out[60]), .A0(n720), .A1(n718), .Z(n719));
Q_OR03 U1135 ( .A0(aux_key_type[0]), .A1(n2122), .A2(n732), .Z(n722));
Q_AN03 U1136 ( .A0(aux_key_type[0]), .A1(n35), .A2(aux_key_type[1]), .Z(n723));
Q_ND02 U1137 ( .A0(aux_key_type[0]), .A1(n2122), .Z(n724));
Q_AN02 U1138 ( .A0(n1972), .A1(n724), .Z(n725));
Q_MX02 U1139 ( .S(aux_key_type[2]), .A0(n725), .A1(n723), .Z(n726));
Q_INV U1140 ( .A(n726), .Z(n727));
Q_MX02 U1141 ( .S(aux_key_type[3]), .A0(n727), .A1(n722), .Z(n728));
Q_OR02 U1142 ( .A0(n143), .A1(n728), .Z(n176));
Q_ND02 U1143 ( .A0(aux_key_type[0]), .A1(n142), .Z(n729));
Q_OR02 U1144 ( .A0(aux_key_type[2]), .A1(aux_key_type[1]), .Z(n732));
Q_OR03 U1145 ( .A0(n730), .A1(n732), .A2(n143), .Z(n177));
Q_NR02 U1146 ( .A0(n2098), .A1(n142), .Z(n731));
Q_MX02 U1147 ( .S(aux_key_type[3]), .A0(n731), .A1(n729), .Z(n730));
Q_LDP0 \_zyL570_tfiRv86_REG[0] ( .G(n443), .D(stitcher_out[56]), .Q(_zyL570_tfiRv86[0]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[1] ( .G(n443), .D(stitcher_out[57]), .Q(_zyL570_tfiRv86[1]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[2] ( .G(n443), .D(stitcher_out[58]), .Q(_zyL570_tfiRv86[2]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[3] ( .G(n443), .D(stitcher_out[59]), .Q(_zyL570_tfiRv86[3]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[4] ( .G(n443), .D(stitcher_out[60]), .Q(_zyL570_tfiRv86[4]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[5] ( .G(n443), .D(stitcher_out[61]), .Q(_zyL570_tfiRv86[5]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[6] ( .G(n443), .D(stitcher_out[62]), .Q(_zyL570_tfiRv86[6]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[7] ( .G(n443), .D(stitcher_out[63]), .Q(_zyL570_tfiRv86[7]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[8] ( .G(n443), .D(stitcher_out[48]), .Q(_zyL570_tfiRv86[8]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[9] ( .G(n443), .D(stitcher_out[49]), .Q(_zyL570_tfiRv86[9]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[10] ( .G(n443), .D(stitcher_out[50]), .Q(_zyL570_tfiRv86[10]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[11] ( .G(n443), .D(stitcher_out[51]), .Q(_zyL570_tfiRv86[11]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[12] ( .G(n443), .D(stitcher_out[52]), .Q(_zyL570_tfiRv86[12]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[13] ( .G(n443), .D(stitcher_out[53]), .Q(_zyL570_tfiRv86[13]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[14] ( .G(n443), .D(stitcher_out[54]), .Q(_zyL570_tfiRv86[14]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[15] ( .G(n443), .D(stitcher_out[55]), .Q(_zyL570_tfiRv86[15]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[16] ( .G(n443), .D(stitcher_out[40]), .Q(_zyL570_tfiRv86[16]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[17] ( .G(n443), .D(stitcher_out[41]), .Q(_zyL570_tfiRv86[17]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[18] ( .G(n443), .D(stitcher_out[42]), .Q(_zyL570_tfiRv86[18]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[19] ( .G(n443), .D(stitcher_out[43]), .Q(_zyL570_tfiRv86[19]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[20] ( .G(n443), .D(stitcher_out[44]), .Q(_zyL570_tfiRv86[20]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[21] ( .G(n443), .D(stitcher_out[45]), .Q(_zyL570_tfiRv86[21]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[22] ( .G(n443), .D(stitcher_out[46]), .Q(_zyL570_tfiRv86[22]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[23] ( .G(n443), .D(stitcher_out[47]), .Q(_zyL570_tfiRv86[23]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[24] ( .G(n443), .D(stitcher_out[32]), .Q(_zyL570_tfiRv86[24]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[25] ( .G(n443), .D(stitcher_out[33]), .Q(_zyL570_tfiRv86[25]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[26] ( .G(n443), .D(stitcher_out[34]), .Q(_zyL570_tfiRv86[26]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[27] ( .G(n443), .D(stitcher_out[35]), .Q(_zyL570_tfiRv86[27]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[28] ( .G(n443), .D(stitcher_out[36]), .Q(_zyL570_tfiRv86[28]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[29] ( .G(n443), .D(stitcher_out[37]), .Q(_zyL570_tfiRv86[29]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[30] ( .G(n443), .D(stitcher_out[38]), .Q(_zyL570_tfiRv86[30]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[31] ( .G(n443), .D(stitcher_out[39]), .Q(_zyL570_tfiRv86[31]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[32] ( .G(n443), .D(stitcher_out[24]), .Q(_zyL570_tfiRv86[32]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[33] ( .G(n443), .D(stitcher_out[25]), .Q(_zyL570_tfiRv86[33]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[34] ( .G(n443), .D(stitcher_out[26]), .Q(_zyL570_tfiRv86[34]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[35] ( .G(n443), .D(stitcher_out[27]), .Q(_zyL570_tfiRv86[35]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[36] ( .G(n443), .D(stitcher_out[28]), .Q(_zyL570_tfiRv86[36]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[37] ( .G(n443), .D(stitcher_out[29]), .Q(_zyL570_tfiRv86[37]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[38] ( .G(n443), .D(stitcher_out[30]), .Q(_zyL570_tfiRv86[38]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[39] ( .G(n443), .D(stitcher_out[31]), .Q(_zyL570_tfiRv86[39]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[40] ( .G(n443), .D(stitcher_out[16]), .Q(_zyL570_tfiRv86[40]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[41] ( .G(n443), .D(stitcher_out[17]), .Q(_zyL570_tfiRv86[41]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[42] ( .G(n443), .D(stitcher_out[18]), .Q(_zyL570_tfiRv86[42]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[43] ( .G(n443), .D(stitcher_out[19]), .Q(_zyL570_tfiRv86[43]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[44] ( .G(n443), .D(stitcher_out[20]), .Q(_zyL570_tfiRv86[44]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[45] ( .G(n443), .D(stitcher_out[21]), .Q(_zyL570_tfiRv86[45]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[46] ( .G(n443), .D(stitcher_out[22]), .Q(_zyL570_tfiRv86[46]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[47] ( .G(n443), .D(stitcher_out[23]), .Q(_zyL570_tfiRv86[47]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[48] ( .G(n443), .D(stitcher_out[8]), .Q(_zyL570_tfiRv86[48]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[49] ( .G(n443), .D(stitcher_out[9]), .Q(_zyL570_tfiRv86[49]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[50] ( .G(n443), .D(stitcher_out[10]), .Q(_zyL570_tfiRv86[50]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[51] ( .G(n443), .D(stitcher_out[11]), .Q(_zyL570_tfiRv86[51]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[52] ( .G(n443), .D(stitcher_out[12]), .Q(_zyL570_tfiRv86[52]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[53] ( .G(n443), .D(stitcher_out[13]), .Q(_zyL570_tfiRv86[53]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[54] ( .G(n443), .D(stitcher_out[14]), .Q(_zyL570_tfiRv86[54]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[55] ( .G(n443), .D(stitcher_out[15]), .Q(_zyL570_tfiRv86[55]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[56] ( .G(n443), .D(stitcher_out[0]), .Q(_zyL570_tfiRv86[56]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[57] ( .G(n443), .D(stitcher_out[1]), .Q(_zyL570_tfiRv86[57]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[58] ( .G(n443), .D(stitcher_out[2]), .Q(_zyL570_tfiRv86[58]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[59] ( .G(n443), .D(stitcher_out[3]), .Q(_zyL570_tfiRv86[59]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[60] ( .G(n443), .D(stitcher_out[4]), .Q(_zyL570_tfiRv86[60]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[61] ( .G(n443), .D(stitcher_out[5]), .Q(_zyL570_tfiRv86[61]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[62] ( .G(n443), .D(stitcher_out[6]), .Q(_zyL570_tfiRv86[62]), .QN( ));
Q_LDP0 \_zyL570_tfiRv86_REG[63] ( .G(n443), .D(stitcher_out[7]), .Q(_zyL570_tfiRv86[63]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[0] ( .G(n447), .D(stitcher_out[56]), .Q(_zyL569_tfiRv85[0]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[1] ( .G(n447), .D(stitcher_out[57]), .Q(_zyL569_tfiRv85[1]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[2] ( .G(n447), .D(stitcher_out[58]), .Q(_zyL569_tfiRv85[2]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[3] ( .G(n447), .D(stitcher_out[59]), .Q(_zyL569_tfiRv85[3]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[4] ( .G(n447), .D(stitcher_out[60]), .Q(_zyL569_tfiRv85[4]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[5] ( .G(n447), .D(stitcher_out[61]), .Q(_zyL569_tfiRv85[5]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[6] ( .G(n447), .D(stitcher_out[62]), .Q(_zyL569_tfiRv85[6]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[7] ( .G(n447), .D(stitcher_out[63]), .Q(_zyL569_tfiRv85[7]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[8] ( .G(n447), .D(stitcher_out[48]), .Q(_zyL569_tfiRv85[8]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[9] ( .G(n447), .D(stitcher_out[49]), .Q(_zyL569_tfiRv85[9]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[10] ( .G(n447), .D(stitcher_out[50]), .Q(_zyL569_tfiRv85[10]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[11] ( .G(n447), .D(stitcher_out[51]), .Q(_zyL569_tfiRv85[11]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[12] ( .G(n447), .D(stitcher_out[52]), .Q(_zyL569_tfiRv85[12]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[13] ( .G(n447), .D(stitcher_out[53]), .Q(_zyL569_tfiRv85[13]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[14] ( .G(n447), .D(stitcher_out[54]), .Q(_zyL569_tfiRv85[14]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[15] ( .G(n447), .D(stitcher_out[55]), .Q(_zyL569_tfiRv85[15]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[16] ( .G(n447), .D(stitcher_out[40]), .Q(_zyL569_tfiRv85[16]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[17] ( .G(n447), .D(stitcher_out[41]), .Q(_zyL569_tfiRv85[17]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[18] ( .G(n447), .D(stitcher_out[42]), .Q(_zyL569_tfiRv85[18]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[19] ( .G(n447), .D(stitcher_out[43]), .Q(_zyL569_tfiRv85[19]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[20] ( .G(n447), .D(stitcher_out[44]), .Q(_zyL569_tfiRv85[20]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[21] ( .G(n447), .D(stitcher_out[45]), .Q(_zyL569_tfiRv85[21]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[22] ( .G(n447), .D(stitcher_out[46]), .Q(_zyL569_tfiRv85[22]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[23] ( .G(n447), .D(stitcher_out[47]), .Q(_zyL569_tfiRv85[23]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[24] ( .G(n447), .D(stitcher_out[32]), .Q(_zyL569_tfiRv85[24]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[25] ( .G(n447), .D(stitcher_out[33]), .Q(_zyL569_tfiRv85[25]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[26] ( .G(n447), .D(stitcher_out[34]), .Q(_zyL569_tfiRv85[26]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[27] ( .G(n447), .D(stitcher_out[35]), .Q(_zyL569_tfiRv85[27]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[28] ( .G(n447), .D(stitcher_out[36]), .Q(_zyL569_tfiRv85[28]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[29] ( .G(n447), .D(stitcher_out[37]), .Q(_zyL569_tfiRv85[29]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[30] ( .G(n447), .D(stitcher_out[38]), .Q(_zyL569_tfiRv85[30]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[31] ( .G(n447), .D(stitcher_out[39]), .Q(_zyL569_tfiRv85[31]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[32] ( .G(n447), .D(stitcher_out[24]), .Q(_zyL569_tfiRv85[32]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[33] ( .G(n447), .D(stitcher_out[25]), .Q(_zyL569_tfiRv85[33]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[34] ( .G(n447), .D(stitcher_out[26]), .Q(_zyL569_tfiRv85[34]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[35] ( .G(n447), .D(stitcher_out[27]), .Q(_zyL569_tfiRv85[35]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[36] ( .G(n447), .D(stitcher_out[28]), .Q(_zyL569_tfiRv85[36]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[37] ( .G(n447), .D(stitcher_out[29]), .Q(_zyL569_tfiRv85[37]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[38] ( .G(n447), .D(stitcher_out[30]), .Q(_zyL569_tfiRv85[38]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[39] ( .G(n447), .D(stitcher_out[31]), .Q(_zyL569_tfiRv85[39]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[40] ( .G(n447), .D(stitcher_out[16]), .Q(_zyL569_tfiRv85[40]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[41] ( .G(n447), .D(stitcher_out[17]), .Q(_zyL569_tfiRv85[41]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[42] ( .G(n447), .D(stitcher_out[18]), .Q(_zyL569_tfiRv85[42]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[43] ( .G(n447), .D(stitcher_out[19]), .Q(_zyL569_tfiRv85[43]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[44] ( .G(n447), .D(stitcher_out[20]), .Q(_zyL569_tfiRv85[44]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[45] ( .G(n447), .D(stitcher_out[21]), .Q(_zyL569_tfiRv85[45]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[46] ( .G(n447), .D(stitcher_out[22]), .Q(_zyL569_tfiRv85[46]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[47] ( .G(n447), .D(stitcher_out[23]), .Q(_zyL569_tfiRv85[47]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[48] ( .G(n447), .D(stitcher_out[8]), .Q(_zyL569_tfiRv85[48]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[49] ( .G(n447), .D(stitcher_out[9]), .Q(_zyL569_tfiRv85[49]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[50] ( .G(n447), .D(stitcher_out[10]), .Q(_zyL569_tfiRv85[50]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[51] ( .G(n447), .D(stitcher_out[11]), .Q(_zyL569_tfiRv85[51]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[52] ( .G(n447), .D(stitcher_out[12]), .Q(_zyL569_tfiRv85[52]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[53] ( .G(n447), .D(stitcher_out[13]), .Q(_zyL569_tfiRv85[53]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[54] ( .G(n447), .D(stitcher_out[14]), .Q(_zyL569_tfiRv85[54]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[55] ( .G(n447), .D(stitcher_out[15]), .Q(_zyL569_tfiRv85[55]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[56] ( .G(n447), .D(stitcher_out[0]), .Q(_zyL569_tfiRv85[56]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[57] ( .G(n447), .D(stitcher_out[1]), .Q(_zyL569_tfiRv85[57]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[58] ( .G(n447), .D(stitcher_out[2]), .Q(_zyL569_tfiRv85[58]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[59] ( .G(n447), .D(stitcher_out[3]), .Q(_zyL569_tfiRv85[59]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[60] ( .G(n447), .D(stitcher_out[4]), .Q(_zyL569_tfiRv85[60]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[61] ( .G(n447), .D(stitcher_out[5]), .Q(_zyL569_tfiRv85[61]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[62] ( .G(n447), .D(stitcher_out[6]), .Q(_zyL569_tfiRv85[62]), .QN( ));
Q_LDP0 \_zyL569_tfiRv85_REG[63] ( .G(n447), .D(stitcher_out[7]), .Q(_zyL569_tfiRv85[63]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[0] ( .G(n452), .D(stitcher_out[56]), .Q(_zyL556_tfiRv84[0]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[1] ( .G(n452), .D(stitcher_out[57]), .Q(_zyL556_tfiRv84[1]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[2] ( .G(n452), .D(stitcher_out[58]), .Q(_zyL556_tfiRv84[2]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[3] ( .G(n452), .D(stitcher_out[59]), .Q(_zyL556_tfiRv84[3]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[4] ( .G(n452), .D(stitcher_out[60]), .Q(_zyL556_tfiRv84[4]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[5] ( .G(n452), .D(stitcher_out[61]), .Q(_zyL556_tfiRv84[5]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[6] ( .G(n452), .D(stitcher_out[62]), .Q(_zyL556_tfiRv84[6]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[7] ( .G(n452), .D(stitcher_out[63]), .Q(_zyL556_tfiRv84[7]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[8] ( .G(n452), .D(stitcher_out[48]), .Q(_zyL556_tfiRv84[8]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[9] ( .G(n452), .D(stitcher_out[49]), .Q(_zyL556_tfiRv84[9]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[10] ( .G(n452), .D(stitcher_out[50]), .Q(_zyL556_tfiRv84[10]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[11] ( .G(n452), .D(stitcher_out[51]), .Q(_zyL556_tfiRv84[11]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[12] ( .G(n452), .D(stitcher_out[52]), .Q(_zyL556_tfiRv84[12]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[13] ( .G(n452), .D(stitcher_out[53]), .Q(_zyL556_tfiRv84[13]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[14] ( .G(n452), .D(stitcher_out[54]), .Q(_zyL556_tfiRv84[14]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[15] ( .G(n452), .D(stitcher_out[55]), .Q(_zyL556_tfiRv84[15]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[16] ( .G(n452), .D(stitcher_out[40]), .Q(_zyL556_tfiRv84[16]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[17] ( .G(n452), .D(stitcher_out[41]), .Q(_zyL556_tfiRv84[17]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[18] ( .G(n452), .D(stitcher_out[42]), .Q(_zyL556_tfiRv84[18]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[19] ( .G(n452), .D(stitcher_out[43]), .Q(_zyL556_tfiRv84[19]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[20] ( .G(n452), .D(stitcher_out[44]), .Q(_zyL556_tfiRv84[20]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[21] ( .G(n452), .D(stitcher_out[45]), .Q(_zyL556_tfiRv84[21]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[22] ( .G(n452), .D(stitcher_out[46]), .Q(_zyL556_tfiRv84[22]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[23] ( .G(n452), .D(stitcher_out[47]), .Q(_zyL556_tfiRv84[23]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[24] ( .G(n452), .D(stitcher_out[32]), .Q(_zyL556_tfiRv84[24]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[25] ( .G(n452), .D(stitcher_out[33]), .Q(_zyL556_tfiRv84[25]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[26] ( .G(n452), .D(stitcher_out[34]), .Q(_zyL556_tfiRv84[26]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[27] ( .G(n452), .D(stitcher_out[35]), .Q(_zyL556_tfiRv84[27]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[28] ( .G(n452), .D(stitcher_out[36]), .Q(_zyL556_tfiRv84[28]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[29] ( .G(n452), .D(stitcher_out[37]), .Q(_zyL556_tfiRv84[29]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[30] ( .G(n452), .D(stitcher_out[38]), .Q(_zyL556_tfiRv84[30]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[31] ( .G(n452), .D(stitcher_out[39]), .Q(_zyL556_tfiRv84[31]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[32] ( .G(n452), .D(stitcher_out[24]), .Q(_zyL556_tfiRv84[32]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[33] ( .G(n452), .D(stitcher_out[25]), .Q(_zyL556_tfiRv84[33]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[34] ( .G(n452), .D(stitcher_out[26]), .Q(_zyL556_tfiRv84[34]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[35] ( .G(n452), .D(stitcher_out[27]), .Q(_zyL556_tfiRv84[35]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[36] ( .G(n452), .D(stitcher_out[28]), .Q(_zyL556_tfiRv84[36]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[37] ( .G(n452), .D(stitcher_out[29]), .Q(_zyL556_tfiRv84[37]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[38] ( .G(n452), .D(stitcher_out[30]), .Q(_zyL556_tfiRv84[38]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[39] ( .G(n452), .D(stitcher_out[31]), .Q(_zyL556_tfiRv84[39]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[40] ( .G(n452), .D(stitcher_out[16]), .Q(_zyL556_tfiRv84[40]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[41] ( .G(n452), .D(stitcher_out[17]), .Q(_zyL556_tfiRv84[41]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[42] ( .G(n452), .D(stitcher_out[18]), .Q(_zyL556_tfiRv84[42]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[43] ( .G(n452), .D(stitcher_out[19]), .Q(_zyL556_tfiRv84[43]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[44] ( .G(n452), .D(stitcher_out[20]), .Q(_zyL556_tfiRv84[44]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[45] ( .G(n452), .D(stitcher_out[21]), .Q(_zyL556_tfiRv84[45]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[46] ( .G(n452), .D(stitcher_out[22]), .Q(_zyL556_tfiRv84[46]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[47] ( .G(n452), .D(stitcher_out[23]), .Q(_zyL556_tfiRv84[47]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[48] ( .G(n452), .D(stitcher_out[8]), .Q(_zyL556_tfiRv84[48]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[49] ( .G(n452), .D(stitcher_out[9]), .Q(_zyL556_tfiRv84[49]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[50] ( .G(n452), .D(stitcher_out[10]), .Q(_zyL556_tfiRv84[50]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[51] ( .G(n452), .D(stitcher_out[11]), .Q(_zyL556_tfiRv84[51]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[52] ( .G(n452), .D(stitcher_out[12]), .Q(_zyL556_tfiRv84[52]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[53] ( .G(n452), .D(stitcher_out[13]), .Q(_zyL556_tfiRv84[53]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[54] ( .G(n452), .D(stitcher_out[14]), .Q(_zyL556_tfiRv84[54]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[55] ( .G(n452), .D(stitcher_out[15]), .Q(_zyL556_tfiRv84[55]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[56] ( .G(n452), .D(stitcher_out[0]), .Q(_zyL556_tfiRv84[56]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[57] ( .G(n452), .D(stitcher_out[1]), .Q(_zyL556_tfiRv84[57]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[58] ( .G(n452), .D(stitcher_out[2]), .Q(_zyL556_tfiRv84[58]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[59] ( .G(n452), .D(stitcher_out[3]), .Q(_zyL556_tfiRv84[59]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[60] ( .G(n452), .D(stitcher_out[4]), .Q(_zyL556_tfiRv84[60]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[61] ( .G(n452), .D(stitcher_out[5]), .Q(_zyL556_tfiRv84[61]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[62] ( .G(n452), .D(stitcher_out[6]), .Q(_zyL556_tfiRv84[62]), .QN( ));
Q_LDP0 \_zyL556_tfiRv84_REG[63] ( .G(n452), .D(stitcher_out[7]), .Q(_zyL556_tfiRv84[63]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[0] ( .G(n456), .D(stitcher_out[56]), .Q(_zyL555_tfiRv83[0]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[1] ( .G(n456), .D(stitcher_out[57]), .Q(_zyL555_tfiRv83[1]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[2] ( .G(n456), .D(stitcher_out[58]), .Q(_zyL555_tfiRv83[2]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[3] ( .G(n456), .D(stitcher_out[59]), .Q(_zyL555_tfiRv83[3]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[4] ( .G(n456), .D(stitcher_out[60]), .Q(_zyL555_tfiRv83[4]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[5] ( .G(n456), .D(stitcher_out[61]), .Q(_zyL555_tfiRv83[5]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[6] ( .G(n456), .D(stitcher_out[62]), .Q(_zyL555_tfiRv83[6]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[7] ( .G(n456), .D(stitcher_out[63]), .Q(_zyL555_tfiRv83[7]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[8] ( .G(n456), .D(stitcher_out[48]), .Q(_zyL555_tfiRv83[8]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[9] ( .G(n456), .D(stitcher_out[49]), .Q(_zyL555_tfiRv83[9]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[10] ( .G(n456), .D(stitcher_out[50]), .Q(_zyL555_tfiRv83[10]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[11] ( .G(n456), .D(stitcher_out[51]), .Q(_zyL555_tfiRv83[11]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[12] ( .G(n456), .D(stitcher_out[52]), .Q(_zyL555_tfiRv83[12]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[13] ( .G(n456), .D(stitcher_out[53]), .Q(_zyL555_tfiRv83[13]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[14] ( .G(n456), .D(stitcher_out[54]), .Q(_zyL555_tfiRv83[14]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[15] ( .G(n456), .D(stitcher_out[55]), .Q(_zyL555_tfiRv83[15]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[16] ( .G(n456), .D(stitcher_out[40]), .Q(_zyL555_tfiRv83[16]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[17] ( .G(n456), .D(stitcher_out[41]), .Q(_zyL555_tfiRv83[17]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[18] ( .G(n456), .D(stitcher_out[42]), .Q(_zyL555_tfiRv83[18]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[19] ( .G(n456), .D(stitcher_out[43]), .Q(_zyL555_tfiRv83[19]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[20] ( .G(n456), .D(stitcher_out[44]), .Q(_zyL555_tfiRv83[20]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[21] ( .G(n456), .D(stitcher_out[45]), .Q(_zyL555_tfiRv83[21]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[22] ( .G(n456), .D(stitcher_out[46]), .Q(_zyL555_tfiRv83[22]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[23] ( .G(n456), .D(stitcher_out[47]), .Q(_zyL555_tfiRv83[23]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[24] ( .G(n456), .D(stitcher_out[32]), .Q(_zyL555_tfiRv83[24]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[25] ( .G(n456), .D(stitcher_out[33]), .Q(_zyL555_tfiRv83[25]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[26] ( .G(n456), .D(stitcher_out[34]), .Q(_zyL555_tfiRv83[26]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[27] ( .G(n456), .D(stitcher_out[35]), .Q(_zyL555_tfiRv83[27]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[28] ( .G(n456), .D(stitcher_out[36]), .Q(_zyL555_tfiRv83[28]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[29] ( .G(n456), .D(stitcher_out[37]), .Q(_zyL555_tfiRv83[29]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[30] ( .G(n456), .D(stitcher_out[38]), .Q(_zyL555_tfiRv83[30]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[31] ( .G(n456), .D(stitcher_out[39]), .Q(_zyL555_tfiRv83[31]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[32] ( .G(n456), .D(stitcher_out[24]), .Q(_zyL555_tfiRv83[32]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[33] ( .G(n456), .D(stitcher_out[25]), .Q(_zyL555_tfiRv83[33]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[34] ( .G(n456), .D(stitcher_out[26]), .Q(_zyL555_tfiRv83[34]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[35] ( .G(n456), .D(stitcher_out[27]), .Q(_zyL555_tfiRv83[35]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[36] ( .G(n456), .D(stitcher_out[28]), .Q(_zyL555_tfiRv83[36]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[37] ( .G(n456), .D(stitcher_out[29]), .Q(_zyL555_tfiRv83[37]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[38] ( .G(n456), .D(stitcher_out[30]), .Q(_zyL555_tfiRv83[38]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[39] ( .G(n456), .D(stitcher_out[31]), .Q(_zyL555_tfiRv83[39]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[40] ( .G(n456), .D(stitcher_out[16]), .Q(_zyL555_tfiRv83[40]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[41] ( .G(n456), .D(stitcher_out[17]), .Q(_zyL555_tfiRv83[41]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[42] ( .G(n456), .D(stitcher_out[18]), .Q(_zyL555_tfiRv83[42]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[43] ( .G(n456), .D(stitcher_out[19]), .Q(_zyL555_tfiRv83[43]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[44] ( .G(n456), .D(stitcher_out[20]), .Q(_zyL555_tfiRv83[44]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[45] ( .G(n456), .D(stitcher_out[21]), .Q(_zyL555_tfiRv83[45]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[46] ( .G(n456), .D(stitcher_out[22]), .Q(_zyL555_tfiRv83[46]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[47] ( .G(n456), .D(stitcher_out[23]), .Q(_zyL555_tfiRv83[47]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[48] ( .G(n456), .D(stitcher_out[8]), .Q(_zyL555_tfiRv83[48]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[49] ( .G(n456), .D(stitcher_out[9]), .Q(_zyL555_tfiRv83[49]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[50] ( .G(n456), .D(stitcher_out[10]), .Q(_zyL555_tfiRv83[50]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[51] ( .G(n456), .D(stitcher_out[11]), .Q(_zyL555_tfiRv83[51]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[52] ( .G(n456), .D(stitcher_out[12]), .Q(_zyL555_tfiRv83[52]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[53] ( .G(n456), .D(stitcher_out[13]), .Q(_zyL555_tfiRv83[53]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[54] ( .G(n456), .D(stitcher_out[14]), .Q(_zyL555_tfiRv83[54]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[55] ( .G(n456), .D(stitcher_out[15]), .Q(_zyL555_tfiRv83[55]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[56] ( .G(n456), .D(stitcher_out[0]), .Q(_zyL555_tfiRv83[56]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[57] ( .G(n456), .D(stitcher_out[1]), .Q(_zyL555_tfiRv83[57]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[58] ( .G(n456), .D(stitcher_out[2]), .Q(_zyL555_tfiRv83[58]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[59] ( .G(n456), .D(stitcher_out[3]), .Q(_zyL555_tfiRv83[59]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[60] ( .G(n456), .D(stitcher_out[4]), .Q(_zyL555_tfiRv83[60]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[61] ( .G(n456), .D(stitcher_out[5]), .Q(_zyL555_tfiRv83[61]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[62] ( .G(n456), .D(stitcher_out[6]), .Q(_zyL555_tfiRv83[62]), .QN( ));
Q_LDP0 \_zyL555_tfiRv83_REG[63] ( .G(n456), .D(stitcher_out[7]), .Q(_zyL555_tfiRv83[63]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[0] ( .G(n458), .D(stitcher_out[56]), .Q(_zyL542_tfiRv82[0]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[1] ( .G(n458), .D(stitcher_out[57]), .Q(_zyL542_tfiRv82[1]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[2] ( .G(n458), .D(stitcher_out[58]), .Q(_zyL542_tfiRv82[2]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[3] ( .G(n458), .D(stitcher_out[59]), .Q(_zyL542_tfiRv82[3]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[4] ( .G(n458), .D(stitcher_out[60]), .Q(_zyL542_tfiRv82[4]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[5] ( .G(n458), .D(stitcher_out[61]), .Q(_zyL542_tfiRv82[5]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[6] ( .G(n458), .D(stitcher_out[62]), .Q(_zyL542_tfiRv82[6]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[7] ( .G(n458), .D(stitcher_out[63]), .Q(_zyL542_tfiRv82[7]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[8] ( .G(n458), .D(stitcher_out[48]), .Q(_zyL542_tfiRv82[8]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[9] ( .G(n458), .D(stitcher_out[49]), .Q(_zyL542_tfiRv82[9]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[10] ( .G(n458), .D(stitcher_out[50]), .Q(_zyL542_tfiRv82[10]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[11] ( .G(n458), .D(stitcher_out[51]), .Q(_zyL542_tfiRv82[11]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[12] ( .G(n458), .D(stitcher_out[52]), .Q(_zyL542_tfiRv82[12]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[13] ( .G(n458), .D(stitcher_out[53]), .Q(_zyL542_tfiRv82[13]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[14] ( .G(n458), .D(stitcher_out[54]), .Q(_zyL542_tfiRv82[14]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[15] ( .G(n458), .D(stitcher_out[55]), .Q(_zyL542_tfiRv82[15]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[16] ( .G(n458), .D(stitcher_out[40]), .Q(_zyL542_tfiRv82[16]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[17] ( .G(n458), .D(stitcher_out[41]), .Q(_zyL542_tfiRv82[17]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[18] ( .G(n458), .D(stitcher_out[42]), .Q(_zyL542_tfiRv82[18]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[19] ( .G(n458), .D(stitcher_out[43]), .Q(_zyL542_tfiRv82[19]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[20] ( .G(n458), .D(stitcher_out[44]), .Q(_zyL542_tfiRv82[20]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[21] ( .G(n458), .D(stitcher_out[45]), .Q(_zyL542_tfiRv82[21]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[22] ( .G(n458), .D(stitcher_out[46]), .Q(_zyL542_tfiRv82[22]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[23] ( .G(n458), .D(stitcher_out[47]), .Q(_zyL542_tfiRv82[23]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[24] ( .G(n458), .D(stitcher_out[32]), .Q(_zyL542_tfiRv82[24]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[25] ( .G(n458), .D(stitcher_out[33]), .Q(_zyL542_tfiRv82[25]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[26] ( .G(n458), .D(stitcher_out[34]), .Q(_zyL542_tfiRv82[26]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[27] ( .G(n458), .D(stitcher_out[35]), .Q(_zyL542_tfiRv82[27]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[28] ( .G(n458), .D(stitcher_out[36]), .Q(_zyL542_tfiRv82[28]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[29] ( .G(n458), .D(stitcher_out[37]), .Q(_zyL542_tfiRv82[29]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[30] ( .G(n458), .D(stitcher_out[38]), .Q(_zyL542_tfiRv82[30]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[31] ( .G(n458), .D(stitcher_out[39]), .Q(_zyL542_tfiRv82[31]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[32] ( .G(n458), .D(stitcher_out[24]), .Q(_zyL542_tfiRv82[32]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[33] ( .G(n458), .D(stitcher_out[25]), .Q(_zyL542_tfiRv82[33]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[34] ( .G(n458), .D(stitcher_out[26]), .Q(_zyL542_tfiRv82[34]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[35] ( .G(n458), .D(stitcher_out[27]), .Q(_zyL542_tfiRv82[35]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[36] ( .G(n458), .D(stitcher_out[28]), .Q(_zyL542_tfiRv82[36]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[37] ( .G(n458), .D(stitcher_out[29]), .Q(_zyL542_tfiRv82[37]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[38] ( .G(n458), .D(stitcher_out[30]), .Q(_zyL542_tfiRv82[38]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[39] ( .G(n458), .D(stitcher_out[31]), .Q(_zyL542_tfiRv82[39]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[40] ( .G(n458), .D(stitcher_out[16]), .Q(_zyL542_tfiRv82[40]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[41] ( .G(n458), .D(stitcher_out[17]), .Q(_zyL542_tfiRv82[41]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[42] ( .G(n458), .D(stitcher_out[18]), .Q(_zyL542_tfiRv82[42]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[43] ( .G(n458), .D(stitcher_out[19]), .Q(_zyL542_tfiRv82[43]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[44] ( .G(n458), .D(stitcher_out[20]), .Q(_zyL542_tfiRv82[44]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[45] ( .G(n458), .D(stitcher_out[21]), .Q(_zyL542_tfiRv82[45]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[46] ( .G(n458), .D(stitcher_out[22]), .Q(_zyL542_tfiRv82[46]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[47] ( .G(n458), .D(stitcher_out[23]), .Q(_zyL542_tfiRv82[47]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[48] ( .G(n458), .D(stitcher_out[8]), .Q(_zyL542_tfiRv82[48]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[49] ( .G(n458), .D(stitcher_out[9]), .Q(_zyL542_tfiRv82[49]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[50] ( .G(n458), .D(stitcher_out[10]), .Q(_zyL542_tfiRv82[50]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[51] ( .G(n458), .D(stitcher_out[11]), .Q(_zyL542_tfiRv82[51]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[52] ( .G(n458), .D(stitcher_out[12]), .Q(_zyL542_tfiRv82[52]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[53] ( .G(n458), .D(stitcher_out[13]), .Q(_zyL542_tfiRv82[53]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[54] ( .G(n458), .D(stitcher_out[14]), .Q(_zyL542_tfiRv82[54]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[55] ( .G(n458), .D(stitcher_out[15]), .Q(_zyL542_tfiRv82[55]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[56] ( .G(n458), .D(stitcher_out[0]), .Q(_zyL542_tfiRv82[56]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[57] ( .G(n458), .D(stitcher_out[1]), .Q(_zyL542_tfiRv82[57]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[58] ( .G(n458), .D(stitcher_out[2]), .Q(_zyL542_tfiRv82[58]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[59] ( .G(n458), .D(stitcher_out[3]), .Q(_zyL542_tfiRv82[59]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[60] ( .G(n458), .D(stitcher_out[4]), .Q(_zyL542_tfiRv82[60]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[61] ( .G(n458), .D(stitcher_out[5]), .Q(_zyL542_tfiRv82[61]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[62] ( .G(n458), .D(stitcher_out[6]), .Q(_zyL542_tfiRv82[62]), .QN( ));
Q_LDP0 \_zyL542_tfiRv82_REG[63] ( .G(n458), .D(stitcher_out[7]), .Q(_zyL542_tfiRv82[63]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[0] ( .G(n462), .D(stitcher_out[56]), .Q(_zyL541_tfiRv81[0]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[1] ( .G(n462), .D(stitcher_out[57]), .Q(_zyL541_tfiRv81[1]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[2] ( .G(n462), .D(stitcher_out[58]), .Q(_zyL541_tfiRv81[2]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[3] ( .G(n462), .D(stitcher_out[59]), .Q(_zyL541_tfiRv81[3]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[4] ( .G(n462), .D(stitcher_out[60]), .Q(_zyL541_tfiRv81[4]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[5] ( .G(n462), .D(stitcher_out[61]), .Q(_zyL541_tfiRv81[5]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[6] ( .G(n462), .D(stitcher_out[62]), .Q(_zyL541_tfiRv81[6]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[7] ( .G(n462), .D(stitcher_out[63]), .Q(_zyL541_tfiRv81[7]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[8] ( .G(n462), .D(stitcher_out[48]), .Q(_zyL541_tfiRv81[8]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[9] ( .G(n462), .D(stitcher_out[49]), .Q(_zyL541_tfiRv81[9]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[10] ( .G(n462), .D(stitcher_out[50]), .Q(_zyL541_tfiRv81[10]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[11] ( .G(n462), .D(stitcher_out[51]), .Q(_zyL541_tfiRv81[11]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[12] ( .G(n462), .D(stitcher_out[52]), .Q(_zyL541_tfiRv81[12]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[13] ( .G(n462), .D(stitcher_out[53]), .Q(_zyL541_tfiRv81[13]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[14] ( .G(n462), .D(stitcher_out[54]), .Q(_zyL541_tfiRv81[14]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[15] ( .G(n462), .D(stitcher_out[55]), .Q(_zyL541_tfiRv81[15]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[16] ( .G(n462), .D(stitcher_out[40]), .Q(_zyL541_tfiRv81[16]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[17] ( .G(n462), .D(stitcher_out[41]), .Q(_zyL541_tfiRv81[17]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[18] ( .G(n462), .D(stitcher_out[42]), .Q(_zyL541_tfiRv81[18]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[19] ( .G(n462), .D(stitcher_out[43]), .Q(_zyL541_tfiRv81[19]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[20] ( .G(n462), .D(stitcher_out[44]), .Q(_zyL541_tfiRv81[20]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[21] ( .G(n462), .D(stitcher_out[45]), .Q(_zyL541_tfiRv81[21]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[22] ( .G(n462), .D(stitcher_out[46]), .Q(_zyL541_tfiRv81[22]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[23] ( .G(n462), .D(stitcher_out[47]), .Q(_zyL541_tfiRv81[23]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[24] ( .G(n462), .D(stitcher_out[32]), .Q(_zyL541_tfiRv81[24]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[25] ( .G(n462), .D(stitcher_out[33]), .Q(_zyL541_tfiRv81[25]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[26] ( .G(n462), .D(stitcher_out[34]), .Q(_zyL541_tfiRv81[26]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[27] ( .G(n462), .D(stitcher_out[35]), .Q(_zyL541_tfiRv81[27]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[28] ( .G(n462), .D(stitcher_out[36]), .Q(_zyL541_tfiRv81[28]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[29] ( .G(n462), .D(stitcher_out[37]), .Q(_zyL541_tfiRv81[29]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[30] ( .G(n462), .D(stitcher_out[38]), .Q(_zyL541_tfiRv81[30]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[31] ( .G(n462), .D(stitcher_out[39]), .Q(_zyL541_tfiRv81[31]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[32] ( .G(n462), .D(stitcher_out[24]), .Q(_zyL541_tfiRv81[32]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[33] ( .G(n462), .D(stitcher_out[25]), .Q(_zyL541_tfiRv81[33]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[34] ( .G(n462), .D(stitcher_out[26]), .Q(_zyL541_tfiRv81[34]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[35] ( .G(n462), .D(stitcher_out[27]), .Q(_zyL541_tfiRv81[35]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[36] ( .G(n462), .D(stitcher_out[28]), .Q(_zyL541_tfiRv81[36]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[37] ( .G(n462), .D(stitcher_out[29]), .Q(_zyL541_tfiRv81[37]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[38] ( .G(n462), .D(stitcher_out[30]), .Q(_zyL541_tfiRv81[38]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[39] ( .G(n462), .D(stitcher_out[31]), .Q(_zyL541_tfiRv81[39]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[40] ( .G(n462), .D(stitcher_out[16]), .Q(_zyL541_tfiRv81[40]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[41] ( .G(n462), .D(stitcher_out[17]), .Q(_zyL541_tfiRv81[41]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[42] ( .G(n462), .D(stitcher_out[18]), .Q(_zyL541_tfiRv81[42]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[43] ( .G(n462), .D(stitcher_out[19]), .Q(_zyL541_tfiRv81[43]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[44] ( .G(n462), .D(stitcher_out[20]), .Q(_zyL541_tfiRv81[44]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[45] ( .G(n462), .D(stitcher_out[21]), .Q(_zyL541_tfiRv81[45]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[46] ( .G(n462), .D(stitcher_out[22]), .Q(_zyL541_tfiRv81[46]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[47] ( .G(n462), .D(stitcher_out[23]), .Q(_zyL541_tfiRv81[47]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[48] ( .G(n462), .D(stitcher_out[8]), .Q(_zyL541_tfiRv81[48]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[49] ( .G(n462), .D(stitcher_out[9]), .Q(_zyL541_tfiRv81[49]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[50] ( .G(n462), .D(stitcher_out[10]), .Q(_zyL541_tfiRv81[50]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[51] ( .G(n462), .D(stitcher_out[11]), .Q(_zyL541_tfiRv81[51]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[52] ( .G(n462), .D(stitcher_out[12]), .Q(_zyL541_tfiRv81[52]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[53] ( .G(n462), .D(stitcher_out[13]), .Q(_zyL541_tfiRv81[53]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[54] ( .G(n462), .D(stitcher_out[14]), .Q(_zyL541_tfiRv81[54]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[55] ( .G(n462), .D(stitcher_out[15]), .Q(_zyL541_tfiRv81[55]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[56] ( .G(n462), .D(stitcher_out[0]), .Q(_zyL541_tfiRv81[56]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[57] ( .G(n462), .D(stitcher_out[1]), .Q(_zyL541_tfiRv81[57]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[58] ( .G(n462), .D(stitcher_out[2]), .Q(_zyL541_tfiRv81[58]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[59] ( .G(n462), .D(stitcher_out[3]), .Q(_zyL541_tfiRv81[59]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[60] ( .G(n462), .D(stitcher_out[4]), .Q(_zyL541_tfiRv81[60]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[61] ( .G(n462), .D(stitcher_out[5]), .Q(_zyL541_tfiRv81[61]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[62] ( .G(n462), .D(stitcher_out[6]), .Q(_zyL541_tfiRv81[62]), .QN( ));
Q_LDP0 \_zyL541_tfiRv81_REG[63] ( .G(n462), .D(stitcher_out[7]), .Q(_zyL541_tfiRv81[63]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[0] ( .G(n464), .D(stitcher_out[56]), .Q(_zyL527_tfiRv80[0]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[1] ( .G(n464), .D(stitcher_out[57]), .Q(_zyL527_tfiRv80[1]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[2] ( .G(n464), .D(stitcher_out[58]), .Q(_zyL527_tfiRv80[2]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[3] ( .G(n464), .D(stitcher_out[59]), .Q(_zyL527_tfiRv80[3]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[4] ( .G(n464), .D(stitcher_out[60]), .Q(_zyL527_tfiRv80[4]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[5] ( .G(n464), .D(stitcher_out[61]), .Q(_zyL527_tfiRv80[5]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[6] ( .G(n464), .D(stitcher_out[62]), .Q(_zyL527_tfiRv80[6]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[7] ( .G(n464), .D(stitcher_out[63]), .Q(_zyL527_tfiRv80[7]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[8] ( .G(n464), .D(stitcher_out[48]), .Q(_zyL527_tfiRv80[8]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[9] ( .G(n464), .D(stitcher_out[49]), .Q(_zyL527_tfiRv80[9]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[10] ( .G(n464), .D(stitcher_out[50]), .Q(_zyL527_tfiRv80[10]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[11] ( .G(n464), .D(stitcher_out[51]), .Q(_zyL527_tfiRv80[11]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[12] ( .G(n464), .D(stitcher_out[52]), .Q(_zyL527_tfiRv80[12]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[13] ( .G(n464), .D(stitcher_out[53]), .Q(_zyL527_tfiRv80[13]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[14] ( .G(n464), .D(stitcher_out[54]), .Q(_zyL527_tfiRv80[14]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[15] ( .G(n464), .D(stitcher_out[55]), .Q(_zyL527_tfiRv80[15]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[16] ( .G(n464), .D(stitcher_out[40]), .Q(_zyL527_tfiRv80[16]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[17] ( .G(n464), .D(stitcher_out[41]), .Q(_zyL527_tfiRv80[17]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[18] ( .G(n464), .D(stitcher_out[42]), .Q(_zyL527_tfiRv80[18]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[19] ( .G(n464), .D(stitcher_out[43]), .Q(_zyL527_tfiRv80[19]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[20] ( .G(n464), .D(stitcher_out[44]), .Q(_zyL527_tfiRv80[20]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[21] ( .G(n464), .D(stitcher_out[45]), .Q(_zyL527_tfiRv80[21]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[22] ( .G(n464), .D(stitcher_out[46]), .Q(_zyL527_tfiRv80[22]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[23] ( .G(n464), .D(stitcher_out[47]), .Q(_zyL527_tfiRv80[23]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[24] ( .G(n464), .D(stitcher_out[32]), .Q(_zyL527_tfiRv80[24]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[25] ( .G(n464), .D(stitcher_out[33]), .Q(_zyL527_tfiRv80[25]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[26] ( .G(n464), .D(stitcher_out[34]), .Q(_zyL527_tfiRv80[26]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[27] ( .G(n464), .D(stitcher_out[35]), .Q(_zyL527_tfiRv80[27]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[28] ( .G(n464), .D(stitcher_out[36]), .Q(_zyL527_tfiRv80[28]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[29] ( .G(n464), .D(stitcher_out[37]), .Q(_zyL527_tfiRv80[29]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[30] ( .G(n464), .D(stitcher_out[38]), .Q(_zyL527_tfiRv80[30]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[31] ( .G(n464), .D(stitcher_out[39]), .Q(_zyL527_tfiRv80[31]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[32] ( .G(n464), .D(stitcher_out[24]), .Q(_zyL527_tfiRv80[32]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[33] ( .G(n464), .D(stitcher_out[25]), .Q(_zyL527_tfiRv80[33]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[34] ( .G(n464), .D(stitcher_out[26]), .Q(_zyL527_tfiRv80[34]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[35] ( .G(n464), .D(stitcher_out[27]), .Q(_zyL527_tfiRv80[35]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[36] ( .G(n464), .D(stitcher_out[28]), .Q(_zyL527_tfiRv80[36]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[37] ( .G(n464), .D(stitcher_out[29]), .Q(_zyL527_tfiRv80[37]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[38] ( .G(n464), .D(stitcher_out[30]), .Q(_zyL527_tfiRv80[38]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[39] ( .G(n464), .D(stitcher_out[31]), .Q(_zyL527_tfiRv80[39]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[40] ( .G(n464), .D(stitcher_out[16]), .Q(_zyL527_tfiRv80[40]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[41] ( .G(n464), .D(stitcher_out[17]), .Q(_zyL527_tfiRv80[41]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[42] ( .G(n464), .D(stitcher_out[18]), .Q(_zyL527_tfiRv80[42]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[43] ( .G(n464), .D(stitcher_out[19]), .Q(_zyL527_tfiRv80[43]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[44] ( .G(n464), .D(stitcher_out[20]), .Q(_zyL527_tfiRv80[44]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[45] ( .G(n464), .D(stitcher_out[21]), .Q(_zyL527_tfiRv80[45]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[46] ( .G(n464), .D(stitcher_out[22]), .Q(_zyL527_tfiRv80[46]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[47] ( .G(n464), .D(stitcher_out[23]), .Q(_zyL527_tfiRv80[47]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[48] ( .G(n464), .D(stitcher_out[8]), .Q(_zyL527_tfiRv80[48]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[49] ( .G(n464), .D(stitcher_out[9]), .Q(_zyL527_tfiRv80[49]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[50] ( .G(n464), .D(stitcher_out[10]), .Q(_zyL527_tfiRv80[50]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[51] ( .G(n464), .D(stitcher_out[11]), .Q(_zyL527_tfiRv80[51]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[52] ( .G(n464), .D(stitcher_out[12]), .Q(_zyL527_tfiRv80[52]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[53] ( .G(n464), .D(stitcher_out[13]), .Q(_zyL527_tfiRv80[53]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[54] ( .G(n464), .D(stitcher_out[14]), .Q(_zyL527_tfiRv80[54]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[55] ( .G(n464), .D(stitcher_out[15]), .Q(_zyL527_tfiRv80[55]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[56] ( .G(n464), .D(stitcher_out[0]), .Q(_zyL527_tfiRv80[56]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[57] ( .G(n464), .D(stitcher_out[1]), .Q(_zyL527_tfiRv80[57]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[58] ( .G(n464), .D(stitcher_out[2]), .Q(_zyL527_tfiRv80[58]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[59] ( .G(n464), .D(stitcher_out[3]), .Q(_zyL527_tfiRv80[59]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[60] ( .G(n464), .D(stitcher_out[4]), .Q(_zyL527_tfiRv80[60]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[61] ( .G(n464), .D(stitcher_out[5]), .Q(_zyL527_tfiRv80[61]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[62] ( .G(n464), .D(stitcher_out[6]), .Q(_zyL527_tfiRv80[62]), .QN( ));
Q_LDP0 \_zyL527_tfiRv80_REG[63] ( .G(n464), .D(stitcher_out[7]), .Q(_zyL527_tfiRv80[63]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[0] ( .G(n469), .D(stitcher_out[56]), .Q(_zyL526_tfiRv79[0]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[1] ( .G(n469), .D(stitcher_out[57]), .Q(_zyL526_tfiRv79[1]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[2] ( .G(n469), .D(stitcher_out[58]), .Q(_zyL526_tfiRv79[2]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[3] ( .G(n469), .D(stitcher_out[59]), .Q(_zyL526_tfiRv79[3]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[4] ( .G(n469), .D(stitcher_out[60]), .Q(_zyL526_tfiRv79[4]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[5] ( .G(n469), .D(stitcher_out[61]), .Q(_zyL526_tfiRv79[5]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[6] ( .G(n469), .D(stitcher_out[62]), .Q(_zyL526_tfiRv79[6]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[7] ( .G(n469), .D(stitcher_out[63]), .Q(_zyL526_tfiRv79[7]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[8] ( .G(n469), .D(stitcher_out[48]), .Q(_zyL526_tfiRv79[8]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[9] ( .G(n469), .D(stitcher_out[49]), .Q(_zyL526_tfiRv79[9]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[10] ( .G(n469), .D(stitcher_out[50]), .Q(_zyL526_tfiRv79[10]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[11] ( .G(n469), .D(stitcher_out[51]), .Q(_zyL526_tfiRv79[11]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[12] ( .G(n469), .D(stitcher_out[52]), .Q(_zyL526_tfiRv79[12]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[13] ( .G(n469), .D(stitcher_out[53]), .Q(_zyL526_tfiRv79[13]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[14] ( .G(n469), .D(stitcher_out[54]), .Q(_zyL526_tfiRv79[14]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[15] ( .G(n469), .D(stitcher_out[55]), .Q(_zyL526_tfiRv79[15]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[16] ( .G(n469), .D(stitcher_out[40]), .Q(_zyL526_tfiRv79[16]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[17] ( .G(n469), .D(stitcher_out[41]), .Q(_zyL526_tfiRv79[17]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[18] ( .G(n469), .D(stitcher_out[42]), .Q(_zyL526_tfiRv79[18]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[19] ( .G(n469), .D(stitcher_out[43]), .Q(_zyL526_tfiRv79[19]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[20] ( .G(n469), .D(stitcher_out[44]), .Q(_zyL526_tfiRv79[20]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[21] ( .G(n469), .D(stitcher_out[45]), .Q(_zyL526_tfiRv79[21]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[22] ( .G(n469), .D(stitcher_out[46]), .Q(_zyL526_tfiRv79[22]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[23] ( .G(n469), .D(stitcher_out[47]), .Q(_zyL526_tfiRv79[23]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[24] ( .G(n469), .D(stitcher_out[32]), .Q(_zyL526_tfiRv79[24]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[25] ( .G(n469), .D(stitcher_out[33]), .Q(_zyL526_tfiRv79[25]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[26] ( .G(n469), .D(stitcher_out[34]), .Q(_zyL526_tfiRv79[26]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[27] ( .G(n469), .D(stitcher_out[35]), .Q(_zyL526_tfiRv79[27]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[28] ( .G(n469), .D(stitcher_out[36]), .Q(_zyL526_tfiRv79[28]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[29] ( .G(n469), .D(stitcher_out[37]), .Q(_zyL526_tfiRv79[29]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[30] ( .G(n469), .D(stitcher_out[38]), .Q(_zyL526_tfiRv79[30]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[31] ( .G(n469), .D(stitcher_out[39]), .Q(_zyL526_tfiRv79[31]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[32] ( .G(n469), .D(stitcher_out[24]), .Q(_zyL526_tfiRv79[32]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[33] ( .G(n469), .D(stitcher_out[25]), .Q(_zyL526_tfiRv79[33]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[34] ( .G(n469), .D(stitcher_out[26]), .Q(_zyL526_tfiRv79[34]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[35] ( .G(n469), .D(stitcher_out[27]), .Q(_zyL526_tfiRv79[35]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[36] ( .G(n469), .D(stitcher_out[28]), .Q(_zyL526_tfiRv79[36]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[37] ( .G(n469), .D(stitcher_out[29]), .Q(_zyL526_tfiRv79[37]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[38] ( .G(n469), .D(stitcher_out[30]), .Q(_zyL526_tfiRv79[38]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[39] ( .G(n469), .D(stitcher_out[31]), .Q(_zyL526_tfiRv79[39]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[40] ( .G(n469), .D(stitcher_out[16]), .Q(_zyL526_tfiRv79[40]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[41] ( .G(n469), .D(stitcher_out[17]), .Q(_zyL526_tfiRv79[41]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[42] ( .G(n469), .D(stitcher_out[18]), .Q(_zyL526_tfiRv79[42]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[43] ( .G(n469), .D(stitcher_out[19]), .Q(_zyL526_tfiRv79[43]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[44] ( .G(n469), .D(stitcher_out[20]), .Q(_zyL526_tfiRv79[44]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[45] ( .G(n469), .D(stitcher_out[21]), .Q(_zyL526_tfiRv79[45]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[46] ( .G(n469), .D(stitcher_out[22]), .Q(_zyL526_tfiRv79[46]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[47] ( .G(n469), .D(stitcher_out[23]), .Q(_zyL526_tfiRv79[47]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[48] ( .G(n469), .D(stitcher_out[8]), .Q(_zyL526_tfiRv79[48]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[49] ( .G(n469), .D(stitcher_out[9]), .Q(_zyL526_tfiRv79[49]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[50] ( .G(n469), .D(stitcher_out[10]), .Q(_zyL526_tfiRv79[50]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[51] ( .G(n469), .D(stitcher_out[11]), .Q(_zyL526_tfiRv79[51]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[52] ( .G(n469), .D(stitcher_out[12]), .Q(_zyL526_tfiRv79[52]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[53] ( .G(n469), .D(stitcher_out[13]), .Q(_zyL526_tfiRv79[53]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[54] ( .G(n469), .D(stitcher_out[14]), .Q(_zyL526_tfiRv79[54]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[55] ( .G(n469), .D(stitcher_out[15]), .Q(_zyL526_tfiRv79[55]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[56] ( .G(n469), .D(stitcher_out[0]), .Q(_zyL526_tfiRv79[56]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[57] ( .G(n469), .D(stitcher_out[1]), .Q(_zyL526_tfiRv79[57]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[58] ( .G(n469), .D(stitcher_out[2]), .Q(_zyL526_tfiRv79[58]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[59] ( .G(n469), .D(stitcher_out[3]), .Q(_zyL526_tfiRv79[59]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[60] ( .G(n469), .D(stitcher_out[4]), .Q(_zyL526_tfiRv79[60]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[61] ( .G(n469), .D(stitcher_out[5]), .Q(_zyL526_tfiRv79[61]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[62] ( .G(n469), .D(stitcher_out[6]), .Q(_zyL526_tfiRv79[62]), .QN( ));
Q_LDP0 \_zyL526_tfiRv79_REG[63] ( .G(n469), .D(stitcher_out[7]), .Q(_zyL526_tfiRv79[63]), .QN( ));
Q_LDN0 _zyL489_tfiRv77_REG  ( .G(n631), .D(n140), .Q(_zyL489_tfiRv77), .QN( ));
Q_LDN0 _zyL489_tfiRv76_REG  ( .G(n631), .D(n145), .Q(_zyL489_tfiRv76), .QN( ));
Q_LDN0 _zyL486_tfiRv75_REG  ( .G(n631), .D(n174), .Q(_zyL486_tfiRv75), .QN( ));
Q_LDN0 _zyL485_tfiRv74_REG  ( .G(n631), .D(n175), .Q(_zyL485_tfiRv74), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[0] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[0]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[1] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[1]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[2] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[2]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[3] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[3]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[4] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[4]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[5] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[5]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[6] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[6]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[7] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[7]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[8] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[8]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[9] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[9]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[10] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[10]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[11] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[11]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[12] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[12]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[13] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[13]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[14] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[14]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[15] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[15]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[16] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[16]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[17] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[17]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[18] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[18]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[19] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[19]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[20] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[20]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[21] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[21]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[22] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[22]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[23] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[23]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[24] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[24]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[25] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[25]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[26] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[26]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[27] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[27]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[28] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[28]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[29] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[29]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[30] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[30]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[31] ( .G(n470), .D(n1735), .Q(_zyL410_tfiRv73[31]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[32] ( .G(n470), .D(stitcher_out[24]), .Q(_zyL410_tfiRv73[32]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[33] ( .G(n470), .D(stitcher_out[25]), .Q(_zyL410_tfiRv73[33]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[34] ( .G(n470), .D(stitcher_out[26]), .Q(_zyL410_tfiRv73[34]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[35] ( .G(n470), .D(stitcher_out[27]), .Q(_zyL410_tfiRv73[35]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[36] ( .G(n470), .D(stitcher_out[28]), .Q(_zyL410_tfiRv73[36]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[37] ( .G(n470), .D(stitcher_out[29]), .Q(_zyL410_tfiRv73[37]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[38] ( .G(n470), .D(stitcher_out[30]), .Q(_zyL410_tfiRv73[38]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[39] ( .G(n470), .D(stitcher_out[31]), .Q(_zyL410_tfiRv73[39]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[40] ( .G(n470), .D(stitcher_out[16]), .Q(_zyL410_tfiRv73[40]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[41] ( .G(n470), .D(stitcher_out[17]), .Q(_zyL410_tfiRv73[41]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[42] ( .G(n470), .D(stitcher_out[18]), .Q(_zyL410_tfiRv73[42]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[43] ( .G(n470), .D(stitcher_out[19]), .Q(_zyL410_tfiRv73[43]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[44] ( .G(n470), .D(stitcher_out[20]), .Q(_zyL410_tfiRv73[44]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[45] ( .G(n470), .D(stitcher_out[21]), .Q(_zyL410_tfiRv73[45]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[46] ( .G(n470), .D(stitcher_out[22]), .Q(_zyL410_tfiRv73[46]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[47] ( .G(n470), .D(stitcher_out[23]), .Q(_zyL410_tfiRv73[47]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[48] ( .G(n470), .D(stitcher_out[8]), .Q(_zyL410_tfiRv73[48]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[49] ( .G(n470), .D(stitcher_out[9]), .Q(_zyL410_tfiRv73[49]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[50] ( .G(n470), .D(stitcher_out[10]), .Q(_zyL410_tfiRv73[50]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[51] ( .G(n470), .D(stitcher_out[11]), .Q(_zyL410_tfiRv73[51]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[52] ( .G(n470), .D(stitcher_out[12]), .Q(_zyL410_tfiRv73[52]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[53] ( .G(n470), .D(stitcher_out[13]), .Q(_zyL410_tfiRv73[53]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[54] ( .G(n470), .D(stitcher_out[14]), .Q(_zyL410_tfiRv73[54]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[55] ( .G(n470), .D(stitcher_out[15]), .Q(_zyL410_tfiRv73[55]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[56] ( .G(n470), .D(stitcher_out[0]), .Q(_zyL410_tfiRv73[56]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[57] ( .G(n470), .D(stitcher_out[1]), .Q(_zyL410_tfiRv73[57]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[58] ( .G(n470), .D(stitcher_out[2]), .Q(_zyL410_tfiRv73[58]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[59] ( .G(n470), .D(stitcher_out[3]), .Q(_zyL410_tfiRv73[59]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[60] ( .G(n470), .D(stitcher_out[4]), .Q(_zyL410_tfiRv73[60]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[61] ( .G(n470), .D(stitcher_out[5]), .Q(_zyL410_tfiRv73[61]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[62] ( .G(n470), .D(stitcher_out[6]), .Q(_zyL410_tfiRv73[62]), .QN( ));
Q_LDP0 \_zyL410_tfiRv73_REG[63] ( .G(n470), .D(stitcher_out[7]), .Q(_zyL410_tfiRv73[63]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[0] ( .G(n472), .D(stitcher_out[24]), .Q(_zyL395_tfiRv72[0]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[1] ( .G(n472), .D(stitcher_out[25]), .Q(_zyL395_tfiRv72[1]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[2] ( .G(n472), .D(stitcher_out[26]), .Q(_zyL395_tfiRv72[2]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[3] ( .G(n472), .D(stitcher_out[27]), .Q(_zyL395_tfiRv72[3]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[4] ( .G(n472), .D(stitcher_out[28]), .Q(_zyL395_tfiRv72[4]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[5] ( .G(n472), .D(stitcher_out[29]), .Q(_zyL395_tfiRv72[5]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[6] ( .G(n472), .D(stitcher_out[30]), .Q(_zyL395_tfiRv72[6]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[7] ( .G(n472), .D(stitcher_out[31]), .Q(_zyL395_tfiRv72[7]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[8] ( .G(n472), .D(stitcher_out[16]), .Q(_zyL395_tfiRv72[8]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[9] ( .G(n472), .D(stitcher_out[17]), .Q(_zyL395_tfiRv72[9]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[10] ( .G(n472), .D(stitcher_out[18]), .Q(_zyL395_tfiRv72[10]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[11] ( .G(n472), .D(stitcher_out[19]), .Q(_zyL395_tfiRv72[11]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[12] ( .G(n472), .D(stitcher_out[20]), .Q(_zyL395_tfiRv72[12]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[13] ( .G(n472), .D(stitcher_out[21]), .Q(_zyL395_tfiRv72[13]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[14] ( .G(n472), .D(stitcher_out[22]), .Q(_zyL395_tfiRv72[14]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[15] ( .G(n472), .D(stitcher_out[23]), .Q(_zyL395_tfiRv72[15]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[16] ( .G(n472), .D(stitcher_out[8]), .Q(_zyL395_tfiRv72[16]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[17] ( .G(n472), .D(stitcher_out[9]), .Q(_zyL395_tfiRv72[17]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[18] ( .G(n472), .D(stitcher_out[10]), .Q(_zyL395_tfiRv72[18]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[19] ( .G(n472), .D(stitcher_out[11]), .Q(_zyL395_tfiRv72[19]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[20] ( .G(n472), .D(stitcher_out[12]), .Q(_zyL395_tfiRv72[20]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[21] ( .G(n472), .D(stitcher_out[13]), .Q(_zyL395_tfiRv72[21]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[22] ( .G(n472), .D(stitcher_out[14]), .Q(_zyL395_tfiRv72[22]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[23] ( .G(n472), .D(stitcher_out[15]), .Q(_zyL395_tfiRv72[23]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[24] ( .G(n472), .D(stitcher_out[0]), .Q(_zyL395_tfiRv72[24]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[25] ( .G(n472), .D(stitcher_out[1]), .Q(_zyL395_tfiRv72[25]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[26] ( .G(n472), .D(stitcher_out[2]), .Q(_zyL395_tfiRv72[26]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[27] ( .G(n472), .D(stitcher_out[3]), .Q(_zyL395_tfiRv72[27]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[28] ( .G(n472), .D(stitcher_out[4]), .Q(_zyL395_tfiRv72[28]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[29] ( .G(n472), .D(stitcher_out[5]), .Q(_zyL395_tfiRv72[29]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[30] ( .G(n472), .D(stitcher_out[6]), .Q(_zyL395_tfiRv72[30]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[31] ( .G(n472), .D(stitcher_out[7]), .Q(_zyL395_tfiRv72[31]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[32] ( .G(n472), .D(buffer[24]), .Q(_zyL395_tfiRv72[32]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[33] ( .G(n472), .D(buffer[25]), .Q(_zyL395_tfiRv72[33]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[34] ( .G(n472), .D(buffer[26]), .Q(_zyL395_tfiRv72[34]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[35] ( .G(n472), .D(buffer[27]), .Q(_zyL395_tfiRv72[35]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[36] ( .G(n472), .D(buffer[28]), .Q(_zyL395_tfiRv72[36]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[37] ( .G(n472), .D(buffer[29]), .Q(_zyL395_tfiRv72[37]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[38] ( .G(n472), .D(buffer[30]), .Q(_zyL395_tfiRv72[38]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[39] ( .G(n472), .D(buffer[31]), .Q(_zyL395_tfiRv72[39]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[40] ( .G(n472), .D(buffer[16]), .Q(_zyL395_tfiRv72[40]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[41] ( .G(n472), .D(buffer[17]), .Q(_zyL395_tfiRv72[41]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[42] ( .G(n472), .D(buffer[18]), .Q(_zyL395_tfiRv72[42]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[43] ( .G(n472), .D(buffer[19]), .Q(_zyL395_tfiRv72[43]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[44] ( .G(n472), .D(buffer[20]), .Q(_zyL395_tfiRv72[44]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[45] ( .G(n472), .D(buffer[21]), .Q(_zyL395_tfiRv72[45]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[46] ( .G(n472), .D(buffer[22]), .Q(_zyL395_tfiRv72[46]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[47] ( .G(n472), .D(buffer[23]), .Q(_zyL395_tfiRv72[47]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[48] ( .G(n472), .D(buffer[8]), .Q(_zyL395_tfiRv72[48]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[49] ( .G(n472), .D(buffer[9]), .Q(_zyL395_tfiRv72[49]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[50] ( .G(n472), .D(buffer[10]), .Q(_zyL395_tfiRv72[50]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[51] ( .G(n472), .D(buffer[11]), .Q(_zyL395_tfiRv72[51]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[52] ( .G(n472), .D(buffer[12]), .Q(_zyL395_tfiRv72[52]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[53] ( .G(n472), .D(buffer[13]), .Q(_zyL395_tfiRv72[53]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[54] ( .G(n472), .D(buffer[14]), .Q(_zyL395_tfiRv72[54]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[55] ( .G(n472), .D(buffer[15]), .Q(_zyL395_tfiRv72[55]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[56] ( .G(n472), .D(buffer[0]), .Q(_zyL395_tfiRv72[56]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[57] ( .G(n472), .D(buffer[1]), .Q(_zyL395_tfiRv72[57]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[58] ( .G(n472), .D(buffer[2]), .Q(_zyL395_tfiRv72[58]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[59] ( .G(n472), .D(buffer[3]), .Q(_zyL395_tfiRv72[59]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[60] ( .G(n472), .D(buffer[4]), .Q(_zyL395_tfiRv72[60]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[61] ( .G(n472), .D(buffer[5]), .Q(_zyL395_tfiRv72[61]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[62] ( .G(n472), .D(buffer[6]), .Q(_zyL395_tfiRv72[62]), .QN( ));
Q_LDP0 \_zyL395_tfiRv72_REG[63] ( .G(n472), .D(buffer[7]), .Q(_zyL395_tfiRv72[63]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[0] ( .G(n473), .D(stitcher_out[56]), .Q(_zyL390_tfiRv71[0]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[1] ( .G(n473), .D(stitcher_out[57]), .Q(_zyL390_tfiRv71[1]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[2] ( .G(n473), .D(stitcher_out[58]), .Q(_zyL390_tfiRv71[2]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[3] ( .G(n473), .D(stitcher_out[59]), .Q(_zyL390_tfiRv71[3]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[4] ( .G(n473), .D(stitcher_out[60]), .Q(_zyL390_tfiRv71[4]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[5] ( .G(n473), .D(stitcher_out[61]), .Q(_zyL390_tfiRv71[5]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[6] ( .G(n473), .D(stitcher_out[62]), .Q(_zyL390_tfiRv71[6]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[7] ( .G(n473), .D(stitcher_out[63]), .Q(_zyL390_tfiRv71[7]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[8] ( .G(n473), .D(stitcher_out[48]), .Q(_zyL390_tfiRv71[8]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[9] ( .G(n473), .D(stitcher_out[49]), .Q(_zyL390_tfiRv71[9]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[10] ( .G(n473), .D(stitcher_out[50]), .Q(_zyL390_tfiRv71[10]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[11] ( .G(n473), .D(stitcher_out[51]), .Q(_zyL390_tfiRv71[11]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[12] ( .G(n473), .D(stitcher_out[52]), .Q(_zyL390_tfiRv71[12]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[13] ( .G(n473), .D(stitcher_out[53]), .Q(_zyL390_tfiRv71[13]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[14] ( .G(n473), .D(stitcher_out[54]), .Q(_zyL390_tfiRv71[14]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[15] ( .G(n473), .D(stitcher_out[55]), .Q(_zyL390_tfiRv71[15]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[16] ( .G(n473), .D(stitcher_out[40]), .Q(_zyL390_tfiRv71[16]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[17] ( .G(n473), .D(stitcher_out[41]), .Q(_zyL390_tfiRv71[17]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[18] ( .G(n473), .D(stitcher_out[42]), .Q(_zyL390_tfiRv71[18]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[19] ( .G(n473), .D(stitcher_out[43]), .Q(_zyL390_tfiRv71[19]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[20] ( .G(n473), .D(stitcher_out[44]), .Q(_zyL390_tfiRv71[20]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[21] ( .G(n473), .D(stitcher_out[45]), .Q(_zyL390_tfiRv71[21]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[22] ( .G(n473), .D(stitcher_out[46]), .Q(_zyL390_tfiRv71[22]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[23] ( .G(n473), .D(stitcher_out[47]), .Q(_zyL390_tfiRv71[23]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[24] ( .G(n473), .D(stitcher_out[32]), .Q(_zyL390_tfiRv71[24]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[25] ( .G(n473), .D(stitcher_out[33]), .Q(_zyL390_tfiRv71[25]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[26] ( .G(n473), .D(stitcher_out[34]), .Q(_zyL390_tfiRv71[26]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[27] ( .G(n473), .D(stitcher_out[35]), .Q(_zyL390_tfiRv71[27]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[28] ( .G(n473), .D(stitcher_out[36]), .Q(_zyL390_tfiRv71[28]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[29] ( .G(n473), .D(stitcher_out[37]), .Q(_zyL390_tfiRv71[29]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[30] ( .G(n473), .D(stitcher_out[38]), .Q(_zyL390_tfiRv71[30]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[31] ( .G(n473), .D(stitcher_out[39]), .Q(_zyL390_tfiRv71[31]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[32] ( .G(n473), .D(stitcher_out[24]), .Q(_zyL390_tfiRv71[32]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[33] ( .G(n473), .D(stitcher_out[25]), .Q(_zyL390_tfiRv71[33]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[34] ( .G(n473), .D(stitcher_out[26]), .Q(_zyL390_tfiRv71[34]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[35] ( .G(n473), .D(stitcher_out[27]), .Q(_zyL390_tfiRv71[35]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[36] ( .G(n473), .D(stitcher_out[28]), .Q(_zyL390_tfiRv71[36]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[37] ( .G(n473), .D(stitcher_out[29]), .Q(_zyL390_tfiRv71[37]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[38] ( .G(n473), .D(stitcher_out[30]), .Q(_zyL390_tfiRv71[38]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[39] ( .G(n473), .D(stitcher_out[31]), .Q(_zyL390_tfiRv71[39]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[40] ( .G(n473), .D(stitcher_out[16]), .Q(_zyL390_tfiRv71[40]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[41] ( .G(n473), .D(stitcher_out[17]), .Q(_zyL390_tfiRv71[41]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[42] ( .G(n473), .D(stitcher_out[18]), .Q(_zyL390_tfiRv71[42]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[43] ( .G(n473), .D(stitcher_out[19]), .Q(_zyL390_tfiRv71[43]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[44] ( .G(n473), .D(stitcher_out[20]), .Q(_zyL390_tfiRv71[44]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[45] ( .G(n473), .D(stitcher_out[21]), .Q(_zyL390_tfiRv71[45]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[46] ( .G(n473), .D(stitcher_out[22]), .Q(_zyL390_tfiRv71[46]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[47] ( .G(n473), .D(stitcher_out[23]), .Q(_zyL390_tfiRv71[47]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[48] ( .G(n473), .D(stitcher_out[8]), .Q(_zyL390_tfiRv71[48]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[49] ( .G(n473), .D(stitcher_out[9]), .Q(_zyL390_tfiRv71[49]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[50] ( .G(n473), .D(stitcher_out[10]), .Q(_zyL390_tfiRv71[50]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[51] ( .G(n473), .D(stitcher_out[11]), .Q(_zyL390_tfiRv71[51]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[52] ( .G(n473), .D(stitcher_out[12]), .Q(_zyL390_tfiRv71[52]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[53] ( .G(n473), .D(stitcher_out[13]), .Q(_zyL390_tfiRv71[53]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[54] ( .G(n473), .D(stitcher_out[14]), .Q(_zyL390_tfiRv71[54]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[55] ( .G(n473), .D(stitcher_out[15]), .Q(_zyL390_tfiRv71[55]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[56] ( .G(n473), .D(stitcher_out[0]), .Q(_zyL390_tfiRv71[56]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[57] ( .G(n473), .D(stitcher_out[1]), .Q(_zyL390_tfiRv71[57]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[58] ( .G(n473), .D(stitcher_out[2]), .Q(_zyL390_tfiRv71[58]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[59] ( .G(n473), .D(stitcher_out[3]), .Q(_zyL390_tfiRv71[59]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[60] ( .G(n473), .D(stitcher_out[4]), .Q(_zyL390_tfiRv71[60]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[61] ( .G(n473), .D(stitcher_out[5]), .Q(_zyL390_tfiRv71[61]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[62] ( .G(n473), .D(stitcher_out[6]), .Q(_zyL390_tfiRv71[62]), .QN( ));
Q_LDN0 \_zyL390_tfiRv71_REG[63] ( .G(n473), .D(stitcher_out[7]), .Q(_zyL390_tfiRv71[63]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[0] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[0]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[1] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[1]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[2] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[2]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[3] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[3]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[4] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[4]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[5] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[5]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[6] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[6]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[7] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[7]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[8] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[8]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[9] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[9]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[10] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[10]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[11] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[11]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[12] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[12]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[13] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[13]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[14] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[14]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[15] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[15]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[16] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[16]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[17] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[17]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[18] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[18]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[19] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[19]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[20] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[20]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[21] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[21]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[22] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[22]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[23] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[23]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[24] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[24]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[25] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[25]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[26] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[26]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[27] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[27]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[28] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[28]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[29] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[29]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[30] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[30]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[31] ( .G(n475), .D(n1735), .Q(_zyL382_tfiRv70[31]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[32] ( .G(n475), .D(stitcher_out[24]), .Q(_zyL382_tfiRv70[32]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[33] ( .G(n475), .D(stitcher_out[25]), .Q(_zyL382_tfiRv70[33]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[34] ( .G(n475), .D(stitcher_out[26]), .Q(_zyL382_tfiRv70[34]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[35] ( .G(n475), .D(stitcher_out[27]), .Q(_zyL382_tfiRv70[35]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[36] ( .G(n475), .D(stitcher_out[28]), .Q(_zyL382_tfiRv70[36]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[37] ( .G(n475), .D(stitcher_out[29]), .Q(_zyL382_tfiRv70[37]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[38] ( .G(n475), .D(stitcher_out[30]), .Q(_zyL382_tfiRv70[38]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[39] ( .G(n475), .D(stitcher_out[31]), .Q(_zyL382_tfiRv70[39]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[40] ( .G(n475), .D(stitcher_out[16]), .Q(_zyL382_tfiRv70[40]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[41] ( .G(n475), .D(stitcher_out[17]), .Q(_zyL382_tfiRv70[41]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[42] ( .G(n475), .D(stitcher_out[18]), .Q(_zyL382_tfiRv70[42]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[43] ( .G(n475), .D(stitcher_out[19]), .Q(_zyL382_tfiRv70[43]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[44] ( .G(n475), .D(stitcher_out[20]), .Q(_zyL382_tfiRv70[44]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[45] ( .G(n475), .D(stitcher_out[21]), .Q(_zyL382_tfiRv70[45]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[46] ( .G(n475), .D(stitcher_out[22]), .Q(_zyL382_tfiRv70[46]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[47] ( .G(n475), .D(stitcher_out[23]), .Q(_zyL382_tfiRv70[47]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[48] ( .G(n475), .D(stitcher_out[8]), .Q(_zyL382_tfiRv70[48]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[49] ( .G(n475), .D(stitcher_out[9]), .Q(_zyL382_tfiRv70[49]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[50] ( .G(n475), .D(stitcher_out[10]), .Q(_zyL382_tfiRv70[50]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[51] ( .G(n475), .D(stitcher_out[11]), .Q(_zyL382_tfiRv70[51]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[52] ( .G(n475), .D(stitcher_out[12]), .Q(_zyL382_tfiRv70[52]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[53] ( .G(n475), .D(stitcher_out[13]), .Q(_zyL382_tfiRv70[53]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[54] ( .G(n475), .D(stitcher_out[14]), .Q(_zyL382_tfiRv70[54]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[55] ( .G(n475), .D(stitcher_out[15]), .Q(_zyL382_tfiRv70[55]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[56] ( .G(n475), .D(stitcher_out[0]), .Q(_zyL382_tfiRv70[56]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[57] ( .G(n475), .D(stitcher_out[1]), .Q(_zyL382_tfiRv70[57]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[58] ( .G(n475), .D(stitcher_out[2]), .Q(_zyL382_tfiRv70[58]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[59] ( .G(n475), .D(stitcher_out[3]), .Q(_zyL382_tfiRv70[59]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[60] ( .G(n475), .D(stitcher_out[4]), .Q(_zyL382_tfiRv70[60]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[61] ( .G(n475), .D(stitcher_out[5]), .Q(_zyL382_tfiRv70[61]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[62] ( .G(n475), .D(stitcher_out[6]), .Q(_zyL382_tfiRv70[62]), .QN( ));
Q_LDP0 \_zyL382_tfiRv70_REG[63] ( .G(n475), .D(stitcher_out[7]), .Q(_zyL382_tfiRv70[63]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[0] ( .G(n477), .D(stitcher_out[24]), .Q(_zyL373_tfiRv69[0]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[1] ( .G(n477), .D(stitcher_out[25]), .Q(_zyL373_tfiRv69[1]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[2] ( .G(n477), .D(stitcher_out[26]), .Q(_zyL373_tfiRv69[2]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[3] ( .G(n477), .D(stitcher_out[27]), .Q(_zyL373_tfiRv69[3]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[4] ( .G(n477), .D(stitcher_out[28]), .Q(_zyL373_tfiRv69[4]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[5] ( .G(n477), .D(stitcher_out[29]), .Q(_zyL373_tfiRv69[5]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[6] ( .G(n477), .D(stitcher_out[30]), .Q(_zyL373_tfiRv69[6]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[7] ( .G(n477), .D(stitcher_out[31]), .Q(_zyL373_tfiRv69[7]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[8] ( .G(n477), .D(stitcher_out[16]), .Q(_zyL373_tfiRv69[8]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[9] ( .G(n477), .D(stitcher_out[17]), .Q(_zyL373_tfiRv69[9]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[10] ( .G(n477), .D(stitcher_out[18]), .Q(_zyL373_tfiRv69[10]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[11] ( .G(n477), .D(stitcher_out[19]), .Q(_zyL373_tfiRv69[11]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[12] ( .G(n477), .D(stitcher_out[20]), .Q(_zyL373_tfiRv69[12]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[13] ( .G(n477), .D(stitcher_out[21]), .Q(_zyL373_tfiRv69[13]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[14] ( .G(n477), .D(stitcher_out[22]), .Q(_zyL373_tfiRv69[14]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[15] ( .G(n477), .D(stitcher_out[23]), .Q(_zyL373_tfiRv69[15]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[16] ( .G(n477), .D(stitcher_out[8]), .Q(_zyL373_tfiRv69[16]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[17] ( .G(n477), .D(stitcher_out[9]), .Q(_zyL373_tfiRv69[17]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[18] ( .G(n477), .D(stitcher_out[10]), .Q(_zyL373_tfiRv69[18]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[19] ( .G(n477), .D(stitcher_out[11]), .Q(_zyL373_tfiRv69[19]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[20] ( .G(n477), .D(stitcher_out[12]), .Q(_zyL373_tfiRv69[20]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[21] ( .G(n477), .D(stitcher_out[13]), .Q(_zyL373_tfiRv69[21]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[22] ( .G(n477), .D(stitcher_out[14]), .Q(_zyL373_tfiRv69[22]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[23] ( .G(n477), .D(stitcher_out[15]), .Q(_zyL373_tfiRv69[23]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[24] ( .G(n477), .D(stitcher_out[0]), .Q(_zyL373_tfiRv69[24]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[25] ( .G(n477), .D(stitcher_out[1]), .Q(_zyL373_tfiRv69[25]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[26] ( .G(n477), .D(stitcher_out[2]), .Q(_zyL373_tfiRv69[26]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[27] ( .G(n477), .D(stitcher_out[3]), .Q(_zyL373_tfiRv69[27]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[28] ( .G(n477), .D(stitcher_out[4]), .Q(_zyL373_tfiRv69[28]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[29] ( .G(n477), .D(stitcher_out[5]), .Q(_zyL373_tfiRv69[29]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[30] ( .G(n477), .D(stitcher_out[6]), .Q(_zyL373_tfiRv69[30]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[31] ( .G(n477), .D(stitcher_out[7]), .Q(_zyL373_tfiRv69[31]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[32] ( .G(n477), .D(buffer[24]), .Q(_zyL373_tfiRv69[32]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[33] ( .G(n477), .D(buffer[25]), .Q(_zyL373_tfiRv69[33]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[34] ( .G(n477), .D(buffer[26]), .Q(_zyL373_tfiRv69[34]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[35] ( .G(n477), .D(buffer[27]), .Q(_zyL373_tfiRv69[35]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[36] ( .G(n477), .D(buffer[28]), .Q(_zyL373_tfiRv69[36]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[37] ( .G(n477), .D(buffer[29]), .Q(_zyL373_tfiRv69[37]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[38] ( .G(n477), .D(buffer[30]), .Q(_zyL373_tfiRv69[38]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[39] ( .G(n477), .D(buffer[31]), .Q(_zyL373_tfiRv69[39]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[40] ( .G(n477), .D(buffer[16]), .Q(_zyL373_tfiRv69[40]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[41] ( .G(n477), .D(buffer[17]), .Q(_zyL373_tfiRv69[41]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[42] ( .G(n477), .D(buffer[18]), .Q(_zyL373_tfiRv69[42]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[43] ( .G(n477), .D(buffer[19]), .Q(_zyL373_tfiRv69[43]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[44] ( .G(n477), .D(buffer[20]), .Q(_zyL373_tfiRv69[44]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[45] ( .G(n477), .D(buffer[21]), .Q(_zyL373_tfiRv69[45]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[46] ( .G(n477), .D(buffer[22]), .Q(_zyL373_tfiRv69[46]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[47] ( .G(n477), .D(buffer[23]), .Q(_zyL373_tfiRv69[47]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[48] ( .G(n477), .D(buffer[8]), .Q(_zyL373_tfiRv69[48]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[49] ( .G(n477), .D(buffer[9]), .Q(_zyL373_tfiRv69[49]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[50] ( .G(n477), .D(buffer[10]), .Q(_zyL373_tfiRv69[50]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[51] ( .G(n477), .D(buffer[11]), .Q(_zyL373_tfiRv69[51]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[52] ( .G(n477), .D(buffer[12]), .Q(_zyL373_tfiRv69[52]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[53] ( .G(n477), .D(buffer[13]), .Q(_zyL373_tfiRv69[53]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[54] ( .G(n477), .D(buffer[14]), .Q(_zyL373_tfiRv69[54]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[55] ( .G(n477), .D(buffer[15]), .Q(_zyL373_tfiRv69[55]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[56] ( .G(n477), .D(buffer[0]), .Q(_zyL373_tfiRv69[56]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[57] ( .G(n477), .D(buffer[1]), .Q(_zyL373_tfiRv69[57]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[58] ( .G(n477), .D(buffer[2]), .Q(_zyL373_tfiRv69[58]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[59] ( .G(n477), .D(buffer[3]), .Q(_zyL373_tfiRv69[59]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[60] ( .G(n477), .D(buffer[4]), .Q(_zyL373_tfiRv69[60]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[61] ( .G(n477), .D(buffer[5]), .Q(_zyL373_tfiRv69[61]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[62] ( .G(n477), .D(buffer[6]), .Q(_zyL373_tfiRv69[62]), .QN( ));
Q_LDP0 \_zyL373_tfiRv69_REG[63] ( .G(n477), .D(buffer[7]), .Q(_zyL373_tfiRv69[63]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[0] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[0]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[1] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[1]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[2] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[2]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[3] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[3]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[4] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[4]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[5] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[5]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[6] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[6]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[7] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[7]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[8] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[8]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[9] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[9]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[10] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[10]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[11] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[11]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[12] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[12]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[13] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[13]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[14] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[14]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[15] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[15]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[16] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[16]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[17] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[17]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[18] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[18]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[19] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[19]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[20] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[20]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[21] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[21]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[22] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[22]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[23] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[23]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[24] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[24]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[25] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[25]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[26] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[26]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[27] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[27]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[28] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[28]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[29] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[29]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[30] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[30]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[31] ( .G(n480), .D(n1735), .Q(_zyL368_tfiRv68[31]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[32] ( .G(n480), .D(stitcher_out[24]), .Q(_zyL368_tfiRv68[32]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[33] ( .G(n480), .D(stitcher_out[25]), .Q(_zyL368_tfiRv68[33]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[34] ( .G(n480), .D(stitcher_out[26]), .Q(_zyL368_tfiRv68[34]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[35] ( .G(n480), .D(stitcher_out[27]), .Q(_zyL368_tfiRv68[35]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[36] ( .G(n480), .D(stitcher_out[28]), .Q(_zyL368_tfiRv68[36]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[37] ( .G(n480), .D(stitcher_out[29]), .Q(_zyL368_tfiRv68[37]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[38] ( .G(n480), .D(stitcher_out[30]), .Q(_zyL368_tfiRv68[38]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[39] ( .G(n480), .D(stitcher_out[31]), .Q(_zyL368_tfiRv68[39]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[40] ( .G(n480), .D(stitcher_out[16]), .Q(_zyL368_tfiRv68[40]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[41] ( .G(n480), .D(stitcher_out[17]), .Q(_zyL368_tfiRv68[41]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[42] ( .G(n480), .D(stitcher_out[18]), .Q(_zyL368_tfiRv68[42]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[43] ( .G(n480), .D(stitcher_out[19]), .Q(_zyL368_tfiRv68[43]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[44] ( .G(n480), .D(stitcher_out[20]), .Q(_zyL368_tfiRv68[44]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[45] ( .G(n480), .D(stitcher_out[21]), .Q(_zyL368_tfiRv68[45]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[46] ( .G(n480), .D(stitcher_out[22]), .Q(_zyL368_tfiRv68[46]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[47] ( .G(n480), .D(stitcher_out[23]), .Q(_zyL368_tfiRv68[47]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[48] ( .G(n480), .D(stitcher_out[8]), .Q(_zyL368_tfiRv68[48]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[49] ( .G(n480), .D(stitcher_out[9]), .Q(_zyL368_tfiRv68[49]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[50] ( .G(n480), .D(stitcher_out[10]), .Q(_zyL368_tfiRv68[50]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[51] ( .G(n480), .D(stitcher_out[11]), .Q(_zyL368_tfiRv68[51]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[52] ( .G(n480), .D(stitcher_out[12]), .Q(_zyL368_tfiRv68[52]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[53] ( .G(n480), .D(stitcher_out[13]), .Q(_zyL368_tfiRv68[53]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[54] ( .G(n480), .D(stitcher_out[14]), .Q(_zyL368_tfiRv68[54]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[55] ( .G(n480), .D(stitcher_out[15]), .Q(_zyL368_tfiRv68[55]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[56] ( .G(n480), .D(stitcher_out[0]), .Q(_zyL368_tfiRv68[56]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[57] ( .G(n480), .D(stitcher_out[1]), .Q(_zyL368_tfiRv68[57]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[58] ( .G(n480), .D(stitcher_out[2]), .Q(_zyL368_tfiRv68[58]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[59] ( .G(n480), .D(stitcher_out[3]), .Q(_zyL368_tfiRv68[59]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[60] ( .G(n480), .D(stitcher_out[4]), .Q(_zyL368_tfiRv68[60]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[61] ( .G(n480), .D(stitcher_out[5]), .Q(_zyL368_tfiRv68[61]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[62] ( .G(n480), .D(stitcher_out[6]), .Q(_zyL368_tfiRv68[62]), .QN( ));
Q_LDP0 \_zyL368_tfiRv68_REG[63] ( .G(n480), .D(stitcher_out[7]), .Q(_zyL368_tfiRv68[63]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[0] ( .G(n482), .D(stitcher_out[24]), .Q(_zyL359_tfiRv67[0]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[1] ( .G(n482), .D(stitcher_out[25]), .Q(_zyL359_tfiRv67[1]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[2] ( .G(n482), .D(stitcher_out[26]), .Q(_zyL359_tfiRv67[2]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[3] ( .G(n482), .D(stitcher_out[27]), .Q(_zyL359_tfiRv67[3]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[4] ( .G(n482), .D(stitcher_out[28]), .Q(_zyL359_tfiRv67[4]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[5] ( .G(n482), .D(stitcher_out[29]), .Q(_zyL359_tfiRv67[5]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[6] ( .G(n482), .D(stitcher_out[30]), .Q(_zyL359_tfiRv67[6]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[7] ( .G(n482), .D(stitcher_out[31]), .Q(_zyL359_tfiRv67[7]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[8] ( .G(n482), .D(stitcher_out[16]), .Q(_zyL359_tfiRv67[8]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[9] ( .G(n482), .D(stitcher_out[17]), .Q(_zyL359_tfiRv67[9]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[10] ( .G(n482), .D(stitcher_out[18]), .Q(_zyL359_tfiRv67[10]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[11] ( .G(n482), .D(stitcher_out[19]), .Q(_zyL359_tfiRv67[11]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[12] ( .G(n482), .D(stitcher_out[20]), .Q(_zyL359_tfiRv67[12]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[13] ( .G(n482), .D(stitcher_out[21]), .Q(_zyL359_tfiRv67[13]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[14] ( .G(n482), .D(stitcher_out[22]), .Q(_zyL359_tfiRv67[14]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[15] ( .G(n482), .D(stitcher_out[23]), .Q(_zyL359_tfiRv67[15]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[16] ( .G(n482), .D(stitcher_out[8]), .Q(_zyL359_tfiRv67[16]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[17] ( .G(n482), .D(stitcher_out[9]), .Q(_zyL359_tfiRv67[17]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[18] ( .G(n482), .D(stitcher_out[10]), .Q(_zyL359_tfiRv67[18]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[19] ( .G(n482), .D(stitcher_out[11]), .Q(_zyL359_tfiRv67[19]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[20] ( .G(n482), .D(stitcher_out[12]), .Q(_zyL359_tfiRv67[20]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[21] ( .G(n482), .D(stitcher_out[13]), .Q(_zyL359_tfiRv67[21]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[22] ( .G(n482), .D(stitcher_out[14]), .Q(_zyL359_tfiRv67[22]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[23] ( .G(n482), .D(stitcher_out[15]), .Q(_zyL359_tfiRv67[23]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[24] ( .G(n482), .D(stitcher_out[0]), .Q(_zyL359_tfiRv67[24]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[25] ( .G(n482), .D(stitcher_out[1]), .Q(_zyL359_tfiRv67[25]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[26] ( .G(n482), .D(stitcher_out[2]), .Q(_zyL359_tfiRv67[26]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[27] ( .G(n482), .D(stitcher_out[3]), .Q(_zyL359_tfiRv67[27]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[28] ( .G(n482), .D(stitcher_out[4]), .Q(_zyL359_tfiRv67[28]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[29] ( .G(n482), .D(stitcher_out[5]), .Q(_zyL359_tfiRv67[29]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[30] ( .G(n482), .D(stitcher_out[6]), .Q(_zyL359_tfiRv67[30]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[31] ( .G(n482), .D(stitcher_out[7]), .Q(_zyL359_tfiRv67[31]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[32] ( .G(n482), .D(buffer[24]), .Q(_zyL359_tfiRv67[32]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[33] ( .G(n482), .D(buffer[25]), .Q(_zyL359_tfiRv67[33]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[34] ( .G(n482), .D(buffer[26]), .Q(_zyL359_tfiRv67[34]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[35] ( .G(n482), .D(buffer[27]), .Q(_zyL359_tfiRv67[35]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[36] ( .G(n482), .D(buffer[28]), .Q(_zyL359_tfiRv67[36]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[37] ( .G(n482), .D(buffer[29]), .Q(_zyL359_tfiRv67[37]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[38] ( .G(n482), .D(buffer[30]), .Q(_zyL359_tfiRv67[38]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[39] ( .G(n482), .D(buffer[31]), .Q(_zyL359_tfiRv67[39]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[40] ( .G(n482), .D(buffer[16]), .Q(_zyL359_tfiRv67[40]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[41] ( .G(n482), .D(buffer[17]), .Q(_zyL359_tfiRv67[41]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[42] ( .G(n482), .D(buffer[18]), .Q(_zyL359_tfiRv67[42]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[43] ( .G(n482), .D(buffer[19]), .Q(_zyL359_tfiRv67[43]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[44] ( .G(n482), .D(buffer[20]), .Q(_zyL359_tfiRv67[44]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[45] ( .G(n482), .D(buffer[21]), .Q(_zyL359_tfiRv67[45]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[46] ( .G(n482), .D(buffer[22]), .Q(_zyL359_tfiRv67[46]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[47] ( .G(n482), .D(buffer[23]), .Q(_zyL359_tfiRv67[47]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[48] ( .G(n482), .D(buffer[8]), .Q(_zyL359_tfiRv67[48]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[49] ( .G(n482), .D(buffer[9]), .Q(_zyL359_tfiRv67[49]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[50] ( .G(n482), .D(buffer[10]), .Q(_zyL359_tfiRv67[50]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[51] ( .G(n482), .D(buffer[11]), .Q(_zyL359_tfiRv67[51]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[52] ( .G(n482), .D(buffer[12]), .Q(_zyL359_tfiRv67[52]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[53] ( .G(n482), .D(buffer[13]), .Q(_zyL359_tfiRv67[53]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[54] ( .G(n482), .D(buffer[14]), .Q(_zyL359_tfiRv67[54]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[55] ( .G(n482), .D(buffer[15]), .Q(_zyL359_tfiRv67[55]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[56] ( .G(n482), .D(buffer[0]), .Q(_zyL359_tfiRv67[56]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[57] ( .G(n482), .D(buffer[1]), .Q(_zyL359_tfiRv67[57]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[58] ( .G(n482), .D(buffer[2]), .Q(_zyL359_tfiRv67[58]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[59] ( .G(n482), .D(buffer[3]), .Q(_zyL359_tfiRv67[59]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[60] ( .G(n482), .D(buffer[4]), .Q(_zyL359_tfiRv67[60]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[61] ( .G(n482), .D(buffer[5]), .Q(_zyL359_tfiRv67[61]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[62] ( .G(n482), .D(buffer[6]), .Q(_zyL359_tfiRv67[62]), .QN( ));
Q_LDP0 \_zyL359_tfiRv67_REG[63] ( .G(n482), .D(buffer[7]), .Q(_zyL359_tfiRv67[63]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[0] ( .G(n483), .D(stitcher_out[56]), .Q(_zyL354_tfiRv66[0]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[1] ( .G(n483), .D(stitcher_out[57]), .Q(_zyL354_tfiRv66[1]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[2] ( .G(n483), .D(stitcher_out[58]), .Q(_zyL354_tfiRv66[2]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[3] ( .G(n483), .D(stitcher_out[59]), .Q(_zyL354_tfiRv66[3]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[4] ( .G(n483), .D(stitcher_out[60]), .Q(_zyL354_tfiRv66[4]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[5] ( .G(n483), .D(stitcher_out[61]), .Q(_zyL354_tfiRv66[5]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[6] ( .G(n483), .D(stitcher_out[62]), .Q(_zyL354_tfiRv66[6]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[7] ( .G(n483), .D(stitcher_out[63]), .Q(_zyL354_tfiRv66[7]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[8] ( .G(n483), .D(stitcher_out[48]), .Q(_zyL354_tfiRv66[8]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[9] ( .G(n483), .D(stitcher_out[49]), .Q(_zyL354_tfiRv66[9]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[10] ( .G(n483), .D(stitcher_out[50]), .Q(_zyL354_tfiRv66[10]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[11] ( .G(n483), .D(stitcher_out[51]), .Q(_zyL354_tfiRv66[11]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[12] ( .G(n483), .D(stitcher_out[52]), .Q(_zyL354_tfiRv66[12]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[13] ( .G(n483), .D(stitcher_out[53]), .Q(_zyL354_tfiRv66[13]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[14] ( .G(n483), .D(stitcher_out[54]), .Q(_zyL354_tfiRv66[14]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[15] ( .G(n483), .D(stitcher_out[55]), .Q(_zyL354_tfiRv66[15]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[16] ( .G(n483), .D(stitcher_out[40]), .Q(_zyL354_tfiRv66[16]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[17] ( .G(n483), .D(stitcher_out[41]), .Q(_zyL354_tfiRv66[17]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[18] ( .G(n483), .D(stitcher_out[42]), .Q(_zyL354_tfiRv66[18]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[19] ( .G(n483), .D(stitcher_out[43]), .Q(_zyL354_tfiRv66[19]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[20] ( .G(n483), .D(stitcher_out[44]), .Q(_zyL354_tfiRv66[20]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[21] ( .G(n483), .D(stitcher_out[45]), .Q(_zyL354_tfiRv66[21]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[22] ( .G(n483), .D(stitcher_out[46]), .Q(_zyL354_tfiRv66[22]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[23] ( .G(n483), .D(stitcher_out[47]), .Q(_zyL354_tfiRv66[23]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[24] ( .G(n483), .D(stitcher_out[32]), .Q(_zyL354_tfiRv66[24]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[25] ( .G(n483), .D(stitcher_out[33]), .Q(_zyL354_tfiRv66[25]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[26] ( .G(n483), .D(stitcher_out[34]), .Q(_zyL354_tfiRv66[26]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[27] ( .G(n483), .D(stitcher_out[35]), .Q(_zyL354_tfiRv66[27]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[28] ( .G(n483), .D(stitcher_out[36]), .Q(_zyL354_tfiRv66[28]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[29] ( .G(n483), .D(stitcher_out[37]), .Q(_zyL354_tfiRv66[29]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[30] ( .G(n483), .D(stitcher_out[38]), .Q(_zyL354_tfiRv66[30]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[31] ( .G(n483), .D(stitcher_out[39]), .Q(_zyL354_tfiRv66[31]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[32] ( .G(n483), .D(stitcher_out[24]), .Q(_zyL354_tfiRv66[32]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[33] ( .G(n483), .D(stitcher_out[25]), .Q(_zyL354_tfiRv66[33]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[34] ( .G(n483), .D(stitcher_out[26]), .Q(_zyL354_tfiRv66[34]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[35] ( .G(n483), .D(stitcher_out[27]), .Q(_zyL354_tfiRv66[35]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[36] ( .G(n483), .D(stitcher_out[28]), .Q(_zyL354_tfiRv66[36]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[37] ( .G(n483), .D(stitcher_out[29]), .Q(_zyL354_tfiRv66[37]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[38] ( .G(n483), .D(stitcher_out[30]), .Q(_zyL354_tfiRv66[38]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[39] ( .G(n483), .D(stitcher_out[31]), .Q(_zyL354_tfiRv66[39]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[40] ( .G(n483), .D(stitcher_out[16]), .Q(_zyL354_tfiRv66[40]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[41] ( .G(n483), .D(stitcher_out[17]), .Q(_zyL354_tfiRv66[41]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[42] ( .G(n483), .D(stitcher_out[18]), .Q(_zyL354_tfiRv66[42]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[43] ( .G(n483), .D(stitcher_out[19]), .Q(_zyL354_tfiRv66[43]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[44] ( .G(n483), .D(stitcher_out[20]), .Q(_zyL354_tfiRv66[44]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[45] ( .G(n483), .D(stitcher_out[21]), .Q(_zyL354_tfiRv66[45]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[46] ( .G(n483), .D(stitcher_out[22]), .Q(_zyL354_tfiRv66[46]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[47] ( .G(n483), .D(stitcher_out[23]), .Q(_zyL354_tfiRv66[47]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[48] ( .G(n483), .D(stitcher_out[8]), .Q(_zyL354_tfiRv66[48]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[49] ( .G(n483), .D(stitcher_out[9]), .Q(_zyL354_tfiRv66[49]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[50] ( .G(n483), .D(stitcher_out[10]), .Q(_zyL354_tfiRv66[50]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[51] ( .G(n483), .D(stitcher_out[11]), .Q(_zyL354_tfiRv66[51]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[52] ( .G(n483), .D(stitcher_out[12]), .Q(_zyL354_tfiRv66[52]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[53] ( .G(n483), .D(stitcher_out[13]), .Q(_zyL354_tfiRv66[53]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[54] ( .G(n483), .D(stitcher_out[14]), .Q(_zyL354_tfiRv66[54]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[55] ( .G(n483), .D(stitcher_out[15]), .Q(_zyL354_tfiRv66[55]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[56] ( .G(n483), .D(stitcher_out[0]), .Q(_zyL354_tfiRv66[56]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[57] ( .G(n483), .D(stitcher_out[1]), .Q(_zyL354_tfiRv66[57]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[58] ( .G(n483), .D(stitcher_out[2]), .Q(_zyL354_tfiRv66[58]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[59] ( .G(n483), .D(stitcher_out[3]), .Q(_zyL354_tfiRv66[59]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[60] ( .G(n483), .D(stitcher_out[4]), .Q(_zyL354_tfiRv66[60]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[61] ( .G(n483), .D(stitcher_out[5]), .Q(_zyL354_tfiRv66[61]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[62] ( .G(n483), .D(stitcher_out[6]), .Q(_zyL354_tfiRv66[62]), .QN( ));
Q_LDN0 \_zyL354_tfiRv66_REG[63] ( .G(n483), .D(stitcher_out[7]), .Q(_zyL354_tfiRv66[63]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[0] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[0]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[1] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[1]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[2] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[2]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[3] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[3]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[4] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[4]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[5] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[5]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[6] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[6]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[7] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[7]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[8] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[8]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[9] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[9]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[10] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[10]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[11] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[11]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[12] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[12]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[13] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[13]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[14] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[14]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[15] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[15]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[16] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[16]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[17] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[17]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[18] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[18]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[19] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[19]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[20] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[20]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[21] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[21]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[22] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[22]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[23] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[23]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[24] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[24]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[25] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[25]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[26] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[26]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[27] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[27]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[28] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[28]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[29] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[29]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[30] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[30]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[31] ( .G(n489), .D(n1735), .Q(_zyL346_tfiRv65[31]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[32] ( .G(n489), .D(stitcher_out[24]), .Q(_zyL346_tfiRv65[32]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[33] ( .G(n489), .D(stitcher_out[25]), .Q(_zyL346_tfiRv65[33]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[34] ( .G(n489), .D(stitcher_out[26]), .Q(_zyL346_tfiRv65[34]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[35] ( .G(n489), .D(stitcher_out[27]), .Q(_zyL346_tfiRv65[35]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[36] ( .G(n489), .D(stitcher_out[28]), .Q(_zyL346_tfiRv65[36]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[37] ( .G(n489), .D(stitcher_out[29]), .Q(_zyL346_tfiRv65[37]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[38] ( .G(n489), .D(stitcher_out[30]), .Q(_zyL346_tfiRv65[38]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[39] ( .G(n489), .D(stitcher_out[31]), .Q(_zyL346_tfiRv65[39]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[40] ( .G(n489), .D(stitcher_out[16]), .Q(_zyL346_tfiRv65[40]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[41] ( .G(n489), .D(stitcher_out[17]), .Q(_zyL346_tfiRv65[41]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[42] ( .G(n489), .D(stitcher_out[18]), .Q(_zyL346_tfiRv65[42]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[43] ( .G(n489), .D(stitcher_out[19]), .Q(_zyL346_tfiRv65[43]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[44] ( .G(n489), .D(stitcher_out[20]), .Q(_zyL346_tfiRv65[44]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[45] ( .G(n489), .D(stitcher_out[21]), .Q(_zyL346_tfiRv65[45]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[46] ( .G(n489), .D(stitcher_out[22]), .Q(_zyL346_tfiRv65[46]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[47] ( .G(n489), .D(stitcher_out[23]), .Q(_zyL346_tfiRv65[47]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[48] ( .G(n489), .D(stitcher_out[8]), .Q(_zyL346_tfiRv65[48]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[49] ( .G(n489), .D(stitcher_out[9]), .Q(_zyL346_tfiRv65[49]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[50] ( .G(n489), .D(stitcher_out[10]), .Q(_zyL346_tfiRv65[50]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[51] ( .G(n489), .D(stitcher_out[11]), .Q(_zyL346_tfiRv65[51]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[52] ( .G(n489), .D(stitcher_out[12]), .Q(_zyL346_tfiRv65[52]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[53] ( .G(n489), .D(stitcher_out[13]), .Q(_zyL346_tfiRv65[53]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[54] ( .G(n489), .D(stitcher_out[14]), .Q(_zyL346_tfiRv65[54]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[55] ( .G(n489), .D(stitcher_out[15]), .Q(_zyL346_tfiRv65[55]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[56] ( .G(n489), .D(stitcher_out[0]), .Q(_zyL346_tfiRv65[56]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[57] ( .G(n489), .D(stitcher_out[1]), .Q(_zyL346_tfiRv65[57]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[58] ( .G(n489), .D(stitcher_out[2]), .Q(_zyL346_tfiRv65[58]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[59] ( .G(n489), .D(stitcher_out[3]), .Q(_zyL346_tfiRv65[59]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[60] ( .G(n489), .D(stitcher_out[4]), .Q(_zyL346_tfiRv65[60]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[61] ( .G(n489), .D(stitcher_out[5]), .Q(_zyL346_tfiRv65[61]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[62] ( .G(n489), .D(stitcher_out[6]), .Q(_zyL346_tfiRv65[62]), .QN( ));
Q_LDN0 \_zyL346_tfiRv65_REG[63] ( .G(n489), .D(stitcher_out[7]), .Q(_zyL346_tfiRv65[63]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[0] ( .G(n496), .D(stitcher_out[24]), .Q(_zyL337_tfiRv64[0]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[1] ( .G(n496), .D(stitcher_out[25]), .Q(_zyL337_tfiRv64[1]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[2] ( .G(n496), .D(stitcher_out[26]), .Q(_zyL337_tfiRv64[2]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[3] ( .G(n496), .D(stitcher_out[27]), .Q(_zyL337_tfiRv64[3]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[4] ( .G(n496), .D(stitcher_out[28]), .Q(_zyL337_tfiRv64[4]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[5] ( .G(n496), .D(stitcher_out[29]), .Q(_zyL337_tfiRv64[5]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[6] ( .G(n496), .D(stitcher_out[30]), .Q(_zyL337_tfiRv64[6]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[7] ( .G(n496), .D(stitcher_out[31]), .Q(_zyL337_tfiRv64[7]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[8] ( .G(n496), .D(stitcher_out[16]), .Q(_zyL337_tfiRv64[8]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[9] ( .G(n496), .D(stitcher_out[17]), .Q(_zyL337_tfiRv64[9]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[10] ( .G(n496), .D(stitcher_out[18]), .Q(_zyL337_tfiRv64[10]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[11] ( .G(n496), .D(stitcher_out[19]), .Q(_zyL337_tfiRv64[11]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[12] ( .G(n496), .D(stitcher_out[20]), .Q(_zyL337_tfiRv64[12]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[13] ( .G(n496), .D(stitcher_out[21]), .Q(_zyL337_tfiRv64[13]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[14] ( .G(n496), .D(stitcher_out[22]), .Q(_zyL337_tfiRv64[14]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[15] ( .G(n496), .D(stitcher_out[23]), .Q(_zyL337_tfiRv64[15]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[16] ( .G(n496), .D(stitcher_out[8]), .Q(_zyL337_tfiRv64[16]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[17] ( .G(n496), .D(stitcher_out[9]), .Q(_zyL337_tfiRv64[17]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[18] ( .G(n496), .D(stitcher_out[10]), .Q(_zyL337_tfiRv64[18]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[19] ( .G(n496), .D(stitcher_out[11]), .Q(_zyL337_tfiRv64[19]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[20] ( .G(n496), .D(stitcher_out[12]), .Q(_zyL337_tfiRv64[20]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[21] ( .G(n496), .D(stitcher_out[13]), .Q(_zyL337_tfiRv64[21]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[22] ( .G(n496), .D(stitcher_out[14]), .Q(_zyL337_tfiRv64[22]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[23] ( .G(n496), .D(stitcher_out[15]), .Q(_zyL337_tfiRv64[23]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[24] ( .G(n496), .D(stitcher_out[0]), .Q(_zyL337_tfiRv64[24]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[25] ( .G(n496), .D(stitcher_out[1]), .Q(_zyL337_tfiRv64[25]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[26] ( .G(n496), .D(stitcher_out[2]), .Q(_zyL337_tfiRv64[26]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[27] ( .G(n496), .D(stitcher_out[3]), .Q(_zyL337_tfiRv64[27]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[28] ( .G(n496), .D(stitcher_out[4]), .Q(_zyL337_tfiRv64[28]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[29] ( .G(n496), .D(stitcher_out[5]), .Q(_zyL337_tfiRv64[29]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[30] ( .G(n496), .D(stitcher_out[6]), .Q(_zyL337_tfiRv64[30]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[31] ( .G(n496), .D(stitcher_out[7]), .Q(_zyL337_tfiRv64[31]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[32] ( .G(n496), .D(buffer[24]), .Q(_zyL337_tfiRv64[32]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[33] ( .G(n496), .D(buffer[25]), .Q(_zyL337_tfiRv64[33]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[34] ( .G(n496), .D(buffer[26]), .Q(_zyL337_tfiRv64[34]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[35] ( .G(n496), .D(buffer[27]), .Q(_zyL337_tfiRv64[35]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[36] ( .G(n496), .D(buffer[28]), .Q(_zyL337_tfiRv64[36]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[37] ( .G(n496), .D(buffer[29]), .Q(_zyL337_tfiRv64[37]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[38] ( .G(n496), .D(buffer[30]), .Q(_zyL337_tfiRv64[38]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[39] ( .G(n496), .D(buffer[31]), .Q(_zyL337_tfiRv64[39]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[40] ( .G(n496), .D(buffer[16]), .Q(_zyL337_tfiRv64[40]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[41] ( .G(n496), .D(buffer[17]), .Q(_zyL337_tfiRv64[41]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[42] ( .G(n496), .D(buffer[18]), .Q(_zyL337_tfiRv64[42]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[43] ( .G(n496), .D(buffer[19]), .Q(_zyL337_tfiRv64[43]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[44] ( .G(n496), .D(buffer[20]), .Q(_zyL337_tfiRv64[44]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[45] ( .G(n496), .D(buffer[21]), .Q(_zyL337_tfiRv64[45]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[46] ( .G(n496), .D(buffer[22]), .Q(_zyL337_tfiRv64[46]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[47] ( .G(n496), .D(buffer[23]), .Q(_zyL337_tfiRv64[47]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[48] ( .G(n496), .D(buffer[8]), .Q(_zyL337_tfiRv64[48]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[49] ( .G(n496), .D(buffer[9]), .Q(_zyL337_tfiRv64[49]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[50] ( .G(n496), .D(buffer[10]), .Q(_zyL337_tfiRv64[50]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[51] ( .G(n496), .D(buffer[11]), .Q(_zyL337_tfiRv64[51]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[52] ( .G(n496), .D(buffer[12]), .Q(_zyL337_tfiRv64[52]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[53] ( .G(n496), .D(buffer[13]), .Q(_zyL337_tfiRv64[53]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[54] ( .G(n496), .D(buffer[14]), .Q(_zyL337_tfiRv64[54]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[55] ( .G(n496), .D(buffer[15]), .Q(_zyL337_tfiRv64[55]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[56] ( .G(n496), .D(buffer[0]), .Q(_zyL337_tfiRv64[56]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[57] ( .G(n496), .D(buffer[1]), .Q(_zyL337_tfiRv64[57]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[58] ( .G(n496), .D(buffer[2]), .Q(_zyL337_tfiRv64[58]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[59] ( .G(n496), .D(buffer[3]), .Q(_zyL337_tfiRv64[59]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[60] ( .G(n496), .D(buffer[4]), .Q(_zyL337_tfiRv64[60]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[61] ( .G(n496), .D(buffer[5]), .Q(_zyL337_tfiRv64[61]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[62] ( .G(n496), .D(buffer[6]), .Q(_zyL337_tfiRv64[62]), .QN( ));
Q_LDP0 \_zyL337_tfiRv64_REG[63] ( .G(n496), .D(buffer[7]), .Q(_zyL337_tfiRv64[63]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[0] ( .G(n499), .D(stitcher_out[24]), .Q(_zyL327_tfiRv63[0]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[1] ( .G(n499), .D(stitcher_out[25]), .Q(_zyL327_tfiRv63[1]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[2] ( .G(n499), .D(stitcher_out[26]), .Q(_zyL327_tfiRv63[2]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[3] ( .G(n499), .D(stitcher_out[27]), .Q(_zyL327_tfiRv63[3]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[4] ( .G(n499), .D(stitcher_out[28]), .Q(_zyL327_tfiRv63[4]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[5] ( .G(n499), .D(stitcher_out[29]), .Q(_zyL327_tfiRv63[5]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[6] ( .G(n499), .D(stitcher_out[30]), .Q(_zyL327_tfiRv63[6]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[7] ( .G(n499), .D(stitcher_out[31]), .Q(_zyL327_tfiRv63[7]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[8] ( .G(n499), .D(stitcher_out[16]), .Q(_zyL327_tfiRv63[8]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[9] ( .G(n499), .D(stitcher_out[17]), .Q(_zyL327_tfiRv63[9]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[10] ( .G(n499), .D(stitcher_out[18]), .Q(_zyL327_tfiRv63[10]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[11] ( .G(n499), .D(stitcher_out[19]), .Q(_zyL327_tfiRv63[11]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[12] ( .G(n499), .D(stitcher_out[20]), .Q(_zyL327_tfiRv63[12]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[13] ( .G(n499), .D(stitcher_out[21]), .Q(_zyL327_tfiRv63[13]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[14] ( .G(n499), .D(stitcher_out[22]), .Q(_zyL327_tfiRv63[14]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[15] ( .G(n499), .D(stitcher_out[23]), .Q(_zyL327_tfiRv63[15]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[16] ( .G(n499), .D(stitcher_out[8]), .Q(_zyL327_tfiRv63[16]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[17] ( .G(n499), .D(stitcher_out[9]), .Q(_zyL327_tfiRv63[17]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[18] ( .G(n499), .D(stitcher_out[10]), .Q(_zyL327_tfiRv63[18]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[19] ( .G(n499), .D(stitcher_out[11]), .Q(_zyL327_tfiRv63[19]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[20] ( .G(n499), .D(stitcher_out[12]), .Q(_zyL327_tfiRv63[20]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[21] ( .G(n499), .D(stitcher_out[13]), .Q(_zyL327_tfiRv63[21]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[22] ( .G(n499), .D(stitcher_out[14]), .Q(_zyL327_tfiRv63[22]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[23] ( .G(n499), .D(stitcher_out[15]), .Q(_zyL327_tfiRv63[23]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[24] ( .G(n499), .D(stitcher_out[0]), .Q(_zyL327_tfiRv63[24]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[25] ( .G(n499), .D(stitcher_out[1]), .Q(_zyL327_tfiRv63[25]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[26] ( .G(n499), .D(stitcher_out[2]), .Q(_zyL327_tfiRv63[26]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[27] ( .G(n499), .D(stitcher_out[3]), .Q(_zyL327_tfiRv63[27]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[28] ( .G(n499), .D(stitcher_out[4]), .Q(_zyL327_tfiRv63[28]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[29] ( .G(n499), .D(stitcher_out[5]), .Q(_zyL327_tfiRv63[29]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[30] ( .G(n499), .D(stitcher_out[6]), .Q(_zyL327_tfiRv63[30]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[31] ( .G(n499), .D(stitcher_out[7]), .Q(_zyL327_tfiRv63[31]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[32] ( .G(n499), .D(buffer[24]), .Q(_zyL327_tfiRv63[32]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[33] ( .G(n499), .D(buffer[25]), .Q(_zyL327_tfiRv63[33]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[34] ( .G(n499), .D(buffer[26]), .Q(_zyL327_tfiRv63[34]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[35] ( .G(n499), .D(buffer[27]), .Q(_zyL327_tfiRv63[35]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[36] ( .G(n499), .D(buffer[28]), .Q(_zyL327_tfiRv63[36]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[37] ( .G(n499), .D(buffer[29]), .Q(_zyL327_tfiRv63[37]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[38] ( .G(n499), .D(buffer[30]), .Q(_zyL327_tfiRv63[38]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[39] ( .G(n499), .D(buffer[31]), .Q(_zyL327_tfiRv63[39]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[40] ( .G(n499), .D(buffer[16]), .Q(_zyL327_tfiRv63[40]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[41] ( .G(n499), .D(buffer[17]), .Q(_zyL327_tfiRv63[41]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[42] ( .G(n499), .D(buffer[18]), .Q(_zyL327_tfiRv63[42]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[43] ( .G(n499), .D(buffer[19]), .Q(_zyL327_tfiRv63[43]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[44] ( .G(n499), .D(buffer[20]), .Q(_zyL327_tfiRv63[44]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[45] ( .G(n499), .D(buffer[21]), .Q(_zyL327_tfiRv63[45]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[46] ( .G(n499), .D(buffer[22]), .Q(_zyL327_tfiRv63[46]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[47] ( .G(n499), .D(buffer[23]), .Q(_zyL327_tfiRv63[47]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[48] ( .G(n499), .D(buffer[8]), .Q(_zyL327_tfiRv63[48]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[49] ( .G(n499), .D(buffer[9]), .Q(_zyL327_tfiRv63[49]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[50] ( .G(n499), .D(buffer[10]), .Q(_zyL327_tfiRv63[50]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[51] ( .G(n499), .D(buffer[11]), .Q(_zyL327_tfiRv63[51]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[52] ( .G(n499), .D(buffer[12]), .Q(_zyL327_tfiRv63[52]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[53] ( .G(n499), .D(buffer[13]), .Q(_zyL327_tfiRv63[53]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[54] ( .G(n499), .D(buffer[14]), .Q(_zyL327_tfiRv63[54]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[55] ( .G(n499), .D(buffer[15]), .Q(_zyL327_tfiRv63[55]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[56] ( .G(n499), .D(buffer[0]), .Q(_zyL327_tfiRv63[56]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[57] ( .G(n499), .D(buffer[1]), .Q(_zyL327_tfiRv63[57]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[58] ( .G(n499), .D(buffer[2]), .Q(_zyL327_tfiRv63[58]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[59] ( .G(n499), .D(buffer[3]), .Q(_zyL327_tfiRv63[59]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[60] ( .G(n499), .D(buffer[4]), .Q(_zyL327_tfiRv63[60]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[61] ( .G(n499), .D(buffer[5]), .Q(_zyL327_tfiRv63[61]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[62] ( .G(n499), .D(buffer[6]), .Q(_zyL327_tfiRv63[62]), .QN( ));
Q_LDP0 \_zyL327_tfiRv63_REG[63] ( .G(n499), .D(buffer[7]), .Q(_zyL327_tfiRv63[63]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[0] ( .G(n500), .D(stitcher_out[56]), .Q(_zyL321_tfiRv62[0]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[1] ( .G(n500), .D(stitcher_out[57]), .Q(_zyL321_tfiRv62[1]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[2] ( .G(n500), .D(stitcher_out[58]), .Q(_zyL321_tfiRv62[2]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[3] ( .G(n500), .D(stitcher_out[59]), .Q(_zyL321_tfiRv62[3]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[4] ( .G(n500), .D(stitcher_out[60]), .Q(_zyL321_tfiRv62[4]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[5] ( .G(n500), .D(stitcher_out[61]), .Q(_zyL321_tfiRv62[5]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[6] ( .G(n500), .D(stitcher_out[62]), .Q(_zyL321_tfiRv62[6]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[7] ( .G(n500), .D(stitcher_out[63]), .Q(_zyL321_tfiRv62[7]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[8] ( .G(n500), .D(stitcher_out[48]), .Q(_zyL321_tfiRv62[8]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[9] ( .G(n500), .D(stitcher_out[49]), .Q(_zyL321_tfiRv62[9]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[10] ( .G(n500), .D(stitcher_out[50]), .Q(_zyL321_tfiRv62[10]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[11] ( .G(n500), .D(stitcher_out[51]), .Q(_zyL321_tfiRv62[11]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[12] ( .G(n500), .D(stitcher_out[52]), .Q(_zyL321_tfiRv62[12]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[13] ( .G(n500), .D(stitcher_out[53]), .Q(_zyL321_tfiRv62[13]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[14] ( .G(n500), .D(stitcher_out[54]), .Q(_zyL321_tfiRv62[14]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[15] ( .G(n500), .D(stitcher_out[55]), .Q(_zyL321_tfiRv62[15]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[16] ( .G(n500), .D(stitcher_out[40]), .Q(_zyL321_tfiRv62[16]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[17] ( .G(n500), .D(stitcher_out[41]), .Q(_zyL321_tfiRv62[17]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[18] ( .G(n500), .D(stitcher_out[42]), .Q(_zyL321_tfiRv62[18]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[19] ( .G(n500), .D(stitcher_out[43]), .Q(_zyL321_tfiRv62[19]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[20] ( .G(n500), .D(stitcher_out[44]), .Q(_zyL321_tfiRv62[20]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[21] ( .G(n500), .D(stitcher_out[45]), .Q(_zyL321_tfiRv62[21]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[22] ( .G(n500), .D(stitcher_out[46]), .Q(_zyL321_tfiRv62[22]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[23] ( .G(n500), .D(stitcher_out[47]), .Q(_zyL321_tfiRv62[23]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[24] ( .G(n500), .D(stitcher_out[32]), .Q(_zyL321_tfiRv62[24]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[25] ( .G(n500), .D(stitcher_out[33]), .Q(_zyL321_tfiRv62[25]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[26] ( .G(n500), .D(stitcher_out[34]), .Q(_zyL321_tfiRv62[26]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[27] ( .G(n500), .D(stitcher_out[35]), .Q(_zyL321_tfiRv62[27]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[28] ( .G(n500), .D(stitcher_out[36]), .Q(_zyL321_tfiRv62[28]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[29] ( .G(n500), .D(stitcher_out[37]), .Q(_zyL321_tfiRv62[29]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[30] ( .G(n500), .D(stitcher_out[38]), .Q(_zyL321_tfiRv62[30]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[31] ( .G(n500), .D(stitcher_out[39]), .Q(_zyL321_tfiRv62[31]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[32] ( .G(n500), .D(stitcher_out[24]), .Q(_zyL321_tfiRv62[32]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[33] ( .G(n500), .D(stitcher_out[25]), .Q(_zyL321_tfiRv62[33]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[34] ( .G(n500), .D(stitcher_out[26]), .Q(_zyL321_tfiRv62[34]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[35] ( .G(n500), .D(stitcher_out[27]), .Q(_zyL321_tfiRv62[35]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[36] ( .G(n500), .D(stitcher_out[28]), .Q(_zyL321_tfiRv62[36]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[37] ( .G(n500), .D(stitcher_out[29]), .Q(_zyL321_tfiRv62[37]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[38] ( .G(n500), .D(stitcher_out[30]), .Q(_zyL321_tfiRv62[38]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[39] ( .G(n500), .D(stitcher_out[31]), .Q(_zyL321_tfiRv62[39]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[40] ( .G(n500), .D(stitcher_out[16]), .Q(_zyL321_tfiRv62[40]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[41] ( .G(n500), .D(stitcher_out[17]), .Q(_zyL321_tfiRv62[41]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[42] ( .G(n500), .D(stitcher_out[18]), .Q(_zyL321_tfiRv62[42]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[43] ( .G(n500), .D(stitcher_out[19]), .Q(_zyL321_tfiRv62[43]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[44] ( .G(n500), .D(stitcher_out[20]), .Q(_zyL321_tfiRv62[44]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[45] ( .G(n500), .D(stitcher_out[21]), .Q(_zyL321_tfiRv62[45]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[46] ( .G(n500), .D(stitcher_out[22]), .Q(_zyL321_tfiRv62[46]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[47] ( .G(n500), .D(stitcher_out[23]), .Q(_zyL321_tfiRv62[47]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[48] ( .G(n500), .D(stitcher_out[8]), .Q(_zyL321_tfiRv62[48]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[49] ( .G(n500), .D(stitcher_out[9]), .Q(_zyL321_tfiRv62[49]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[50] ( .G(n500), .D(stitcher_out[10]), .Q(_zyL321_tfiRv62[50]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[51] ( .G(n500), .D(stitcher_out[11]), .Q(_zyL321_tfiRv62[51]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[52] ( .G(n500), .D(stitcher_out[12]), .Q(_zyL321_tfiRv62[52]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[53] ( .G(n500), .D(stitcher_out[13]), .Q(_zyL321_tfiRv62[53]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[54] ( .G(n500), .D(stitcher_out[14]), .Q(_zyL321_tfiRv62[54]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[55] ( .G(n500), .D(stitcher_out[15]), .Q(_zyL321_tfiRv62[55]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[56] ( .G(n500), .D(stitcher_out[0]), .Q(_zyL321_tfiRv62[56]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[57] ( .G(n500), .D(stitcher_out[1]), .Q(_zyL321_tfiRv62[57]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[58] ( .G(n500), .D(stitcher_out[2]), .Q(_zyL321_tfiRv62[58]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[59] ( .G(n500), .D(stitcher_out[3]), .Q(_zyL321_tfiRv62[59]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[60] ( .G(n500), .D(stitcher_out[4]), .Q(_zyL321_tfiRv62[60]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[61] ( .G(n500), .D(stitcher_out[5]), .Q(_zyL321_tfiRv62[61]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[62] ( .G(n500), .D(stitcher_out[6]), .Q(_zyL321_tfiRv62[62]), .QN( ));
Q_LDN0 \_zyL321_tfiRv62_REG[63] ( .G(n500), .D(stitcher_out[7]), .Q(_zyL321_tfiRv62[63]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[0] ( .G(n505), .D(stitcher_out[24]), .Q(_zyL313_tfiRv61[0]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[1] ( .G(n505), .D(stitcher_out[25]), .Q(_zyL313_tfiRv61[1]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[2] ( .G(n505), .D(stitcher_out[26]), .Q(_zyL313_tfiRv61[2]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[3] ( .G(n505), .D(stitcher_out[27]), .Q(_zyL313_tfiRv61[3]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[4] ( .G(n505), .D(stitcher_out[28]), .Q(_zyL313_tfiRv61[4]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[5] ( .G(n505), .D(stitcher_out[29]), .Q(_zyL313_tfiRv61[5]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[6] ( .G(n505), .D(stitcher_out[30]), .Q(_zyL313_tfiRv61[6]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[7] ( .G(n505), .D(stitcher_out[31]), .Q(_zyL313_tfiRv61[7]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[8] ( .G(n505), .D(stitcher_out[16]), .Q(_zyL313_tfiRv61[8]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[9] ( .G(n505), .D(stitcher_out[17]), .Q(_zyL313_tfiRv61[9]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[10] ( .G(n505), .D(stitcher_out[18]), .Q(_zyL313_tfiRv61[10]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[11] ( .G(n505), .D(stitcher_out[19]), .Q(_zyL313_tfiRv61[11]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[12] ( .G(n505), .D(stitcher_out[20]), .Q(_zyL313_tfiRv61[12]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[13] ( .G(n505), .D(stitcher_out[21]), .Q(_zyL313_tfiRv61[13]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[14] ( .G(n505), .D(stitcher_out[22]), .Q(_zyL313_tfiRv61[14]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[15] ( .G(n505), .D(stitcher_out[23]), .Q(_zyL313_tfiRv61[15]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[16] ( .G(n505), .D(stitcher_out[8]), .Q(_zyL313_tfiRv61[16]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[17] ( .G(n505), .D(stitcher_out[9]), .Q(_zyL313_tfiRv61[17]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[18] ( .G(n505), .D(stitcher_out[10]), .Q(_zyL313_tfiRv61[18]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[19] ( .G(n505), .D(stitcher_out[11]), .Q(_zyL313_tfiRv61[19]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[20] ( .G(n505), .D(stitcher_out[12]), .Q(_zyL313_tfiRv61[20]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[21] ( .G(n505), .D(stitcher_out[13]), .Q(_zyL313_tfiRv61[21]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[22] ( .G(n505), .D(stitcher_out[14]), .Q(_zyL313_tfiRv61[22]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[23] ( .G(n505), .D(stitcher_out[15]), .Q(_zyL313_tfiRv61[23]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[24] ( .G(n505), .D(stitcher_out[0]), .Q(_zyL313_tfiRv61[24]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[25] ( .G(n505), .D(stitcher_out[1]), .Q(_zyL313_tfiRv61[25]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[26] ( .G(n505), .D(stitcher_out[2]), .Q(_zyL313_tfiRv61[26]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[27] ( .G(n505), .D(stitcher_out[3]), .Q(_zyL313_tfiRv61[27]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[28] ( .G(n505), .D(stitcher_out[4]), .Q(_zyL313_tfiRv61[28]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[29] ( .G(n505), .D(stitcher_out[5]), .Q(_zyL313_tfiRv61[29]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[30] ( .G(n505), .D(stitcher_out[6]), .Q(_zyL313_tfiRv61[30]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[31] ( .G(n505), .D(stitcher_out[7]), .Q(_zyL313_tfiRv61[31]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[32] ( .G(n505), .D(buffer[24]), .Q(_zyL313_tfiRv61[32]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[33] ( .G(n505), .D(buffer[25]), .Q(_zyL313_tfiRv61[33]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[34] ( .G(n505), .D(buffer[26]), .Q(_zyL313_tfiRv61[34]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[35] ( .G(n505), .D(buffer[27]), .Q(_zyL313_tfiRv61[35]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[36] ( .G(n505), .D(buffer[28]), .Q(_zyL313_tfiRv61[36]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[37] ( .G(n505), .D(buffer[29]), .Q(_zyL313_tfiRv61[37]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[38] ( .G(n505), .D(buffer[30]), .Q(_zyL313_tfiRv61[38]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[39] ( .G(n505), .D(buffer[31]), .Q(_zyL313_tfiRv61[39]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[40] ( .G(n505), .D(buffer[16]), .Q(_zyL313_tfiRv61[40]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[41] ( .G(n505), .D(buffer[17]), .Q(_zyL313_tfiRv61[41]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[42] ( .G(n505), .D(buffer[18]), .Q(_zyL313_tfiRv61[42]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[43] ( .G(n505), .D(buffer[19]), .Q(_zyL313_tfiRv61[43]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[44] ( .G(n505), .D(buffer[20]), .Q(_zyL313_tfiRv61[44]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[45] ( .G(n505), .D(buffer[21]), .Q(_zyL313_tfiRv61[45]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[46] ( .G(n505), .D(buffer[22]), .Q(_zyL313_tfiRv61[46]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[47] ( .G(n505), .D(buffer[23]), .Q(_zyL313_tfiRv61[47]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[48] ( .G(n505), .D(buffer[8]), .Q(_zyL313_tfiRv61[48]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[49] ( .G(n505), .D(buffer[9]), .Q(_zyL313_tfiRv61[49]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[50] ( .G(n505), .D(buffer[10]), .Q(_zyL313_tfiRv61[50]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[51] ( .G(n505), .D(buffer[11]), .Q(_zyL313_tfiRv61[51]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[52] ( .G(n505), .D(buffer[12]), .Q(_zyL313_tfiRv61[52]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[53] ( .G(n505), .D(buffer[13]), .Q(_zyL313_tfiRv61[53]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[54] ( .G(n505), .D(buffer[14]), .Q(_zyL313_tfiRv61[54]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[55] ( .G(n505), .D(buffer[15]), .Q(_zyL313_tfiRv61[55]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[56] ( .G(n505), .D(buffer[0]), .Q(_zyL313_tfiRv61[56]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[57] ( .G(n505), .D(buffer[1]), .Q(_zyL313_tfiRv61[57]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[58] ( .G(n505), .D(buffer[2]), .Q(_zyL313_tfiRv61[58]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[59] ( .G(n505), .D(buffer[3]), .Q(_zyL313_tfiRv61[59]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[60] ( .G(n505), .D(buffer[4]), .Q(_zyL313_tfiRv61[60]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[61] ( .G(n505), .D(buffer[5]), .Q(_zyL313_tfiRv61[61]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[62] ( .G(n505), .D(buffer[6]), .Q(_zyL313_tfiRv61[62]), .QN( ));
Q_LDP0 \_zyL313_tfiRv61_REG[63] ( .G(n505), .D(buffer[7]), .Q(_zyL313_tfiRv61[63]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[0] ( .G(n515), .D(stitcher_out[24]), .Q(_zyL306_tfiRv60[0]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[1] ( .G(n515), .D(stitcher_out[25]), .Q(_zyL306_tfiRv60[1]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[2] ( .G(n515), .D(stitcher_out[26]), .Q(_zyL306_tfiRv60[2]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[3] ( .G(n515), .D(stitcher_out[27]), .Q(_zyL306_tfiRv60[3]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[4] ( .G(n515), .D(stitcher_out[28]), .Q(_zyL306_tfiRv60[4]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[5] ( .G(n515), .D(stitcher_out[29]), .Q(_zyL306_tfiRv60[5]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[6] ( .G(n515), .D(stitcher_out[30]), .Q(_zyL306_tfiRv60[6]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[7] ( .G(n515), .D(stitcher_out[31]), .Q(_zyL306_tfiRv60[7]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[8] ( .G(n515), .D(stitcher_out[16]), .Q(_zyL306_tfiRv60[8]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[9] ( .G(n515), .D(stitcher_out[17]), .Q(_zyL306_tfiRv60[9]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[10] ( .G(n515), .D(stitcher_out[18]), .Q(_zyL306_tfiRv60[10]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[11] ( .G(n515), .D(stitcher_out[19]), .Q(_zyL306_tfiRv60[11]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[12] ( .G(n515), .D(stitcher_out[20]), .Q(_zyL306_tfiRv60[12]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[13] ( .G(n515), .D(stitcher_out[21]), .Q(_zyL306_tfiRv60[13]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[14] ( .G(n515), .D(stitcher_out[22]), .Q(_zyL306_tfiRv60[14]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[15] ( .G(n515), .D(stitcher_out[23]), .Q(_zyL306_tfiRv60[15]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[16] ( .G(n515), .D(stitcher_out[8]), .Q(_zyL306_tfiRv60[16]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[17] ( .G(n515), .D(stitcher_out[9]), .Q(_zyL306_tfiRv60[17]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[18] ( .G(n515), .D(stitcher_out[10]), .Q(_zyL306_tfiRv60[18]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[19] ( .G(n515), .D(stitcher_out[11]), .Q(_zyL306_tfiRv60[19]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[20] ( .G(n515), .D(stitcher_out[12]), .Q(_zyL306_tfiRv60[20]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[21] ( .G(n515), .D(stitcher_out[13]), .Q(_zyL306_tfiRv60[21]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[22] ( .G(n515), .D(stitcher_out[14]), .Q(_zyL306_tfiRv60[22]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[23] ( .G(n515), .D(stitcher_out[15]), .Q(_zyL306_tfiRv60[23]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[24] ( .G(n515), .D(stitcher_out[0]), .Q(_zyL306_tfiRv60[24]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[25] ( .G(n515), .D(stitcher_out[1]), .Q(_zyL306_tfiRv60[25]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[26] ( .G(n515), .D(stitcher_out[2]), .Q(_zyL306_tfiRv60[26]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[27] ( .G(n515), .D(stitcher_out[3]), .Q(_zyL306_tfiRv60[27]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[28] ( .G(n515), .D(stitcher_out[4]), .Q(_zyL306_tfiRv60[28]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[29] ( .G(n515), .D(stitcher_out[5]), .Q(_zyL306_tfiRv60[29]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[30] ( .G(n515), .D(stitcher_out[6]), .Q(_zyL306_tfiRv60[30]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[31] ( .G(n515), .D(stitcher_out[7]), .Q(_zyL306_tfiRv60[31]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[32] ( .G(n515), .D(buffer[24]), .Q(_zyL306_tfiRv60[32]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[33] ( .G(n515), .D(buffer[25]), .Q(_zyL306_tfiRv60[33]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[34] ( .G(n515), .D(buffer[26]), .Q(_zyL306_tfiRv60[34]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[35] ( .G(n515), .D(buffer[27]), .Q(_zyL306_tfiRv60[35]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[36] ( .G(n515), .D(buffer[28]), .Q(_zyL306_tfiRv60[36]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[37] ( .G(n515), .D(buffer[29]), .Q(_zyL306_tfiRv60[37]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[38] ( .G(n515), .D(buffer[30]), .Q(_zyL306_tfiRv60[38]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[39] ( .G(n515), .D(buffer[31]), .Q(_zyL306_tfiRv60[39]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[40] ( .G(n515), .D(buffer[16]), .Q(_zyL306_tfiRv60[40]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[41] ( .G(n515), .D(buffer[17]), .Q(_zyL306_tfiRv60[41]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[42] ( .G(n515), .D(buffer[18]), .Q(_zyL306_tfiRv60[42]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[43] ( .G(n515), .D(buffer[19]), .Q(_zyL306_tfiRv60[43]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[44] ( .G(n515), .D(buffer[20]), .Q(_zyL306_tfiRv60[44]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[45] ( .G(n515), .D(buffer[21]), .Q(_zyL306_tfiRv60[45]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[46] ( .G(n515), .D(buffer[22]), .Q(_zyL306_tfiRv60[46]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[47] ( .G(n515), .D(buffer[23]), .Q(_zyL306_tfiRv60[47]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[48] ( .G(n515), .D(buffer[8]), .Q(_zyL306_tfiRv60[48]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[49] ( .G(n515), .D(buffer[9]), .Q(_zyL306_tfiRv60[49]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[50] ( .G(n515), .D(buffer[10]), .Q(_zyL306_tfiRv60[50]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[51] ( .G(n515), .D(buffer[11]), .Q(_zyL306_tfiRv60[51]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[52] ( .G(n515), .D(buffer[12]), .Q(_zyL306_tfiRv60[52]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[53] ( .G(n515), .D(buffer[13]), .Q(_zyL306_tfiRv60[53]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[54] ( .G(n515), .D(buffer[14]), .Q(_zyL306_tfiRv60[54]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[55] ( .G(n515), .D(buffer[15]), .Q(_zyL306_tfiRv60[55]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[56] ( .G(n515), .D(buffer[0]), .Q(_zyL306_tfiRv60[56]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[57] ( .G(n515), .D(buffer[1]), .Q(_zyL306_tfiRv60[57]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[58] ( .G(n515), .D(buffer[2]), .Q(_zyL306_tfiRv60[58]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[59] ( .G(n515), .D(buffer[3]), .Q(_zyL306_tfiRv60[59]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[60] ( .G(n515), .D(buffer[4]), .Q(_zyL306_tfiRv60[60]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[61] ( .G(n515), .D(buffer[5]), .Q(_zyL306_tfiRv60[61]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[62] ( .G(n515), .D(buffer[6]), .Q(_zyL306_tfiRv60[62]), .QN( ));
Q_LDP0 \_zyL306_tfiRv60_REG[63] ( .G(n515), .D(buffer[7]), .Q(_zyL306_tfiRv60[63]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[0] ( .G(n516), .D(stitcher_out[24]), .Q(_zyL301_tfiRv59[0]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[1] ( .G(n516), .D(stitcher_out[25]), .Q(_zyL301_tfiRv59[1]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[2] ( .G(n516), .D(stitcher_out[26]), .Q(_zyL301_tfiRv59[2]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[3] ( .G(n516), .D(stitcher_out[27]), .Q(_zyL301_tfiRv59[3]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[4] ( .G(n516), .D(stitcher_out[28]), .Q(_zyL301_tfiRv59[4]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[5] ( .G(n516), .D(stitcher_out[29]), .Q(_zyL301_tfiRv59[5]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[6] ( .G(n516), .D(stitcher_out[30]), .Q(_zyL301_tfiRv59[6]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[7] ( .G(n516), .D(stitcher_out[31]), .Q(_zyL301_tfiRv59[7]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[8] ( .G(n516), .D(stitcher_out[16]), .Q(_zyL301_tfiRv59[8]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[9] ( .G(n516), .D(stitcher_out[17]), .Q(_zyL301_tfiRv59[9]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[10] ( .G(n516), .D(stitcher_out[18]), .Q(_zyL301_tfiRv59[10]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[11] ( .G(n516), .D(stitcher_out[19]), .Q(_zyL301_tfiRv59[11]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[12] ( .G(n516), .D(stitcher_out[20]), .Q(_zyL301_tfiRv59[12]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[13] ( .G(n516), .D(stitcher_out[21]), .Q(_zyL301_tfiRv59[13]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[14] ( .G(n516), .D(stitcher_out[22]), .Q(_zyL301_tfiRv59[14]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[15] ( .G(n516), .D(stitcher_out[23]), .Q(_zyL301_tfiRv59[15]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[16] ( .G(n516), .D(stitcher_out[8]), .Q(_zyL301_tfiRv59[16]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[17] ( .G(n516), .D(stitcher_out[9]), .Q(_zyL301_tfiRv59[17]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[18] ( .G(n516), .D(stitcher_out[10]), .Q(_zyL301_tfiRv59[18]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[19] ( .G(n516), .D(stitcher_out[11]), .Q(_zyL301_tfiRv59[19]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[20] ( .G(n516), .D(stitcher_out[12]), .Q(_zyL301_tfiRv59[20]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[21] ( .G(n516), .D(stitcher_out[13]), .Q(_zyL301_tfiRv59[21]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[22] ( .G(n516), .D(stitcher_out[14]), .Q(_zyL301_tfiRv59[22]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[23] ( .G(n516), .D(stitcher_out[15]), .Q(_zyL301_tfiRv59[23]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[24] ( .G(n516), .D(stitcher_out[0]), .Q(_zyL301_tfiRv59[24]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[25] ( .G(n516), .D(stitcher_out[1]), .Q(_zyL301_tfiRv59[25]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[26] ( .G(n516), .D(stitcher_out[2]), .Q(_zyL301_tfiRv59[26]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[27] ( .G(n516), .D(stitcher_out[3]), .Q(_zyL301_tfiRv59[27]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[28] ( .G(n516), .D(stitcher_out[4]), .Q(_zyL301_tfiRv59[28]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[29] ( .G(n516), .D(stitcher_out[5]), .Q(_zyL301_tfiRv59[29]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[30] ( .G(n516), .D(stitcher_out[6]), .Q(_zyL301_tfiRv59[30]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[31] ( .G(n516), .D(stitcher_out[7]), .Q(_zyL301_tfiRv59[31]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[32] ( .G(n516), .D(buffer[24]), .Q(_zyL301_tfiRv59[32]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[33] ( .G(n516), .D(buffer[25]), .Q(_zyL301_tfiRv59[33]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[34] ( .G(n516), .D(buffer[26]), .Q(_zyL301_tfiRv59[34]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[35] ( .G(n516), .D(buffer[27]), .Q(_zyL301_tfiRv59[35]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[36] ( .G(n516), .D(buffer[28]), .Q(_zyL301_tfiRv59[36]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[37] ( .G(n516), .D(buffer[29]), .Q(_zyL301_tfiRv59[37]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[38] ( .G(n516), .D(buffer[30]), .Q(_zyL301_tfiRv59[38]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[39] ( .G(n516), .D(buffer[31]), .Q(_zyL301_tfiRv59[39]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[40] ( .G(n516), .D(buffer[16]), .Q(_zyL301_tfiRv59[40]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[41] ( .G(n516), .D(buffer[17]), .Q(_zyL301_tfiRv59[41]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[42] ( .G(n516), .D(buffer[18]), .Q(_zyL301_tfiRv59[42]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[43] ( .G(n516), .D(buffer[19]), .Q(_zyL301_tfiRv59[43]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[44] ( .G(n516), .D(buffer[20]), .Q(_zyL301_tfiRv59[44]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[45] ( .G(n516), .D(buffer[21]), .Q(_zyL301_tfiRv59[45]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[46] ( .G(n516), .D(buffer[22]), .Q(_zyL301_tfiRv59[46]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[47] ( .G(n516), .D(buffer[23]), .Q(_zyL301_tfiRv59[47]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[48] ( .G(n516), .D(buffer[8]), .Q(_zyL301_tfiRv59[48]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[49] ( .G(n516), .D(buffer[9]), .Q(_zyL301_tfiRv59[49]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[50] ( .G(n516), .D(buffer[10]), .Q(_zyL301_tfiRv59[50]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[51] ( .G(n516), .D(buffer[11]), .Q(_zyL301_tfiRv59[51]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[52] ( .G(n516), .D(buffer[12]), .Q(_zyL301_tfiRv59[52]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[53] ( .G(n516), .D(buffer[13]), .Q(_zyL301_tfiRv59[53]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[54] ( .G(n516), .D(buffer[14]), .Q(_zyL301_tfiRv59[54]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[55] ( .G(n516), .D(buffer[15]), .Q(_zyL301_tfiRv59[55]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[56] ( .G(n516), .D(buffer[0]), .Q(_zyL301_tfiRv59[56]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[57] ( .G(n516), .D(buffer[1]), .Q(_zyL301_tfiRv59[57]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[58] ( .G(n516), .D(buffer[2]), .Q(_zyL301_tfiRv59[58]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[59] ( .G(n516), .D(buffer[3]), .Q(_zyL301_tfiRv59[59]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[60] ( .G(n516), .D(buffer[4]), .Q(_zyL301_tfiRv59[60]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[61] ( .G(n516), .D(buffer[5]), .Q(_zyL301_tfiRv59[61]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[62] ( .G(n516), .D(buffer[6]), .Q(_zyL301_tfiRv59[62]), .QN( ));
Q_LDN0 \_zyL301_tfiRv59_REG[63] ( .G(n516), .D(buffer[7]), .Q(_zyL301_tfiRv59[63]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[0] ( .G(n521), .D(stitcher_out[24]), .Q(_zyL293_tfiRv58[0]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[1] ( .G(n521), .D(stitcher_out[25]), .Q(_zyL293_tfiRv58[1]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[2] ( .G(n521), .D(stitcher_out[26]), .Q(_zyL293_tfiRv58[2]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[3] ( .G(n521), .D(stitcher_out[27]), .Q(_zyL293_tfiRv58[3]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[4] ( .G(n521), .D(stitcher_out[28]), .Q(_zyL293_tfiRv58[4]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[5] ( .G(n521), .D(stitcher_out[29]), .Q(_zyL293_tfiRv58[5]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[6] ( .G(n521), .D(stitcher_out[30]), .Q(_zyL293_tfiRv58[6]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[7] ( .G(n521), .D(stitcher_out[31]), .Q(_zyL293_tfiRv58[7]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[8] ( .G(n521), .D(stitcher_out[16]), .Q(_zyL293_tfiRv58[8]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[9] ( .G(n521), .D(stitcher_out[17]), .Q(_zyL293_tfiRv58[9]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[10] ( .G(n521), .D(stitcher_out[18]), .Q(_zyL293_tfiRv58[10]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[11] ( .G(n521), .D(stitcher_out[19]), .Q(_zyL293_tfiRv58[11]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[12] ( .G(n521), .D(stitcher_out[20]), .Q(_zyL293_tfiRv58[12]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[13] ( .G(n521), .D(stitcher_out[21]), .Q(_zyL293_tfiRv58[13]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[14] ( .G(n521), .D(stitcher_out[22]), .Q(_zyL293_tfiRv58[14]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[15] ( .G(n521), .D(stitcher_out[23]), .Q(_zyL293_tfiRv58[15]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[16] ( .G(n521), .D(stitcher_out[8]), .Q(_zyL293_tfiRv58[16]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[17] ( .G(n521), .D(stitcher_out[9]), .Q(_zyL293_tfiRv58[17]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[18] ( .G(n521), .D(stitcher_out[10]), .Q(_zyL293_tfiRv58[18]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[19] ( .G(n521), .D(stitcher_out[11]), .Q(_zyL293_tfiRv58[19]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[20] ( .G(n521), .D(stitcher_out[12]), .Q(_zyL293_tfiRv58[20]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[21] ( .G(n521), .D(stitcher_out[13]), .Q(_zyL293_tfiRv58[21]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[22] ( .G(n521), .D(stitcher_out[14]), .Q(_zyL293_tfiRv58[22]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[23] ( .G(n521), .D(stitcher_out[15]), .Q(_zyL293_tfiRv58[23]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[24] ( .G(n521), .D(stitcher_out[0]), .Q(_zyL293_tfiRv58[24]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[25] ( .G(n521), .D(stitcher_out[1]), .Q(_zyL293_tfiRv58[25]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[26] ( .G(n521), .D(stitcher_out[2]), .Q(_zyL293_tfiRv58[26]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[27] ( .G(n521), .D(stitcher_out[3]), .Q(_zyL293_tfiRv58[27]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[28] ( .G(n521), .D(stitcher_out[4]), .Q(_zyL293_tfiRv58[28]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[29] ( .G(n521), .D(stitcher_out[5]), .Q(_zyL293_tfiRv58[29]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[30] ( .G(n521), .D(stitcher_out[6]), .Q(_zyL293_tfiRv58[30]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[31] ( .G(n521), .D(stitcher_out[7]), .Q(_zyL293_tfiRv58[31]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[32] ( .G(n521), .D(buffer[24]), .Q(_zyL293_tfiRv58[32]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[33] ( .G(n521), .D(buffer[25]), .Q(_zyL293_tfiRv58[33]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[34] ( .G(n521), .D(buffer[26]), .Q(_zyL293_tfiRv58[34]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[35] ( .G(n521), .D(buffer[27]), .Q(_zyL293_tfiRv58[35]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[36] ( .G(n521), .D(buffer[28]), .Q(_zyL293_tfiRv58[36]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[37] ( .G(n521), .D(buffer[29]), .Q(_zyL293_tfiRv58[37]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[38] ( .G(n521), .D(buffer[30]), .Q(_zyL293_tfiRv58[38]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[39] ( .G(n521), .D(buffer[31]), .Q(_zyL293_tfiRv58[39]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[40] ( .G(n521), .D(buffer[16]), .Q(_zyL293_tfiRv58[40]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[41] ( .G(n521), .D(buffer[17]), .Q(_zyL293_tfiRv58[41]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[42] ( .G(n521), .D(buffer[18]), .Q(_zyL293_tfiRv58[42]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[43] ( .G(n521), .D(buffer[19]), .Q(_zyL293_tfiRv58[43]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[44] ( .G(n521), .D(buffer[20]), .Q(_zyL293_tfiRv58[44]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[45] ( .G(n521), .D(buffer[21]), .Q(_zyL293_tfiRv58[45]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[46] ( .G(n521), .D(buffer[22]), .Q(_zyL293_tfiRv58[46]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[47] ( .G(n521), .D(buffer[23]), .Q(_zyL293_tfiRv58[47]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[48] ( .G(n521), .D(buffer[8]), .Q(_zyL293_tfiRv58[48]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[49] ( .G(n521), .D(buffer[9]), .Q(_zyL293_tfiRv58[49]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[50] ( .G(n521), .D(buffer[10]), .Q(_zyL293_tfiRv58[50]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[51] ( .G(n521), .D(buffer[11]), .Q(_zyL293_tfiRv58[51]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[52] ( .G(n521), .D(buffer[12]), .Q(_zyL293_tfiRv58[52]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[53] ( .G(n521), .D(buffer[13]), .Q(_zyL293_tfiRv58[53]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[54] ( .G(n521), .D(buffer[14]), .Q(_zyL293_tfiRv58[54]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[55] ( .G(n521), .D(buffer[15]), .Q(_zyL293_tfiRv58[55]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[56] ( .G(n521), .D(buffer[0]), .Q(_zyL293_tfiRv58[56]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[57] ( .G(n521), .D(buffer[1]), .Q(_zyL293_tfiRv58[57]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[58] ( .G(n521), .D(buffer[2]), .Q(_zyL293_tfiRv58[58]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[59] ( .G(n521), .D(buffer[3]), .Q(_zyL293_tfiRv58[59]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[60] ( .G(n521), .D(buffer[4]), .Q(_zyL293_tfiRv58[60]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[61] ( .G(n521), .D(buffer[5]), .Q(_zyL293_tfiRv58[61]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[62] ( .G(n521), .D(buffer[6]), .Q(_zyL293_tfiRv58[62]), .QN( ));
Q_LDP0 \_zyL293_tfiRv58_REG[63] ( .G(n521), .D(buffer[7]), .Q(_zyL293_tfiRv58[63]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[0] ( .G(n525), .D(stitcher_out[24]), .Q(_zyL288_tfiRv57[0]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[1] ( .G(n525), .D(stitcher_out[25]), .Q(_zyL288_tfiRv57[1]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[2] ( .G(n525), .D(stitcher_out[26]), .Q(_zyL288_tfiRv57[2]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[3] ( .G(n525), .D(stitcher_out[27]), .Q(_zyL288_tfiRv57[3]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[4] ( .G(n525), .D(stitcher_out[28]), .Q(_zyL288_tfiRv57[4]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[5] ( .G(n525), .D(stitcher_out[29]), .Q(_zyL288_tfiRv57[5]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[6] ( .G(n525), .D(stitcher_out[30]), .Q(_zyL288_tfiRv57[6]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[7] ( .G(n525), .D(stitcher_out[31]), .Q(_zyL288_tfiRv57[7]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[8] ( .G(n525), .D(stitcher_out[16]), .Q(_zyL288_tfiRv57[8]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[9] ( .G(n525), .D(stitcher_out[17]), .Q(_zyL288_tfiRv57[9]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[10] ( .G(n525), .D(stitcher_out[18]), .Q(_zyL288_tfiRv57[10]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[11] ( .G(n525), .D(stitcher_out[19]), .Q(_zyL288_tfiRv57[11]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[12] ( .G(n525), .D(stitcher_out[20]), .Q(_zyL288_tfiRv57[12]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[13] ( .G(n525), .D(stitcher_out[21]), .Q(_zyL288_tfiRv57[13]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[14] ( .G(n525), .D(stitcher_out[22]), .Q(_zyL288_tfiRv57[14]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[15] ( .G(n525), .D(stitcher_out[23]), .Q(_zyL288_tfiRv57[15]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[16] ( .G(n525), .D(stitcher_out[8]), .Q(_zyL288_tfiRv57[16]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[17] ( .G(n525), .D(stitcher_out[9]), .Q(_zyL288_tfiRv57[17]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[18] ( .G(n525), .D(stitcher_out[10]), .Q(_zyL288_tfiRv57[18]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[19] ( .G(n525), .D(stitcher_out[11]), .Q(_zyL288_tfiRv57[19]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[20] ( .G(n525), .D(stitcher_out[12]), .Q(_zyL288_tfiRv57[20]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[21] ( .G(n525), .D(stitcher_out[13]), .Q(_zyL288_tfiRv57[21]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[22] ( .G(n525), .D(stitcher_out[14]), .Q(_zyL288_tfiRv57[22]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[23] ( .G(n525), .D(stitcher_out[15]), .Q(_zyL288_tfiRv57[23]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[24] ( .G(n525), .D(stitcher_out[0]), .Q(_zyL288_tfiRv57[24]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[25] ( .G(n525), .D(stitcher_out[1]), .Q(_zyL288_tfiRv57[25]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[26] ( .G(n525), .D(stitcher_out[2]), .Q(_zyL288_tfiRv57[26]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[27] ( .G(n525), .D(stitcher_out[3]), .Q(_zyL288_tfiRv57[27]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[28] ( .G(n525), .D(stitcher_out[4]), .Q(_zyL288_tfiRv57[28]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[29] ( .G(n525), .D(stitcher_out[5]), .Q(_zyL288_tfiRv57[29]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[30] ( .G(n525), .D(stitcher_out[6]), .Q(_zyL288_tfiRv57[30]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[31] ( .G(n525), .D(stitcher_out[7]), .Q(_zyL288_tfiRv57[31]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[32] ( .G(n525), .D(buffer[24]), .Q(_zyL288_tfiRv57[32]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[33] ( .G(n525), .D(buffer[25]), .Q(_zyL288_tfiRv57[33]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[34] ( .G(n525), .D(buffer[26]), .Q(_zyL288_tfiRv57[34]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[35] ( .G(n525), .D(buffer[27]), .Q(_zyL288_tfiRv57[35]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[36] ( .G(n525), .D(buffer[28]), .Q(_zyL288_tfiRv57[36]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[37] ( .G(n525), .D(buffer[29]), .Q(_zyL288_tfiRv57[37]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[38] ( .G(n525), .D(buffer[30]), .Q(_zyL288_tfiRv57[38]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[39] ( .G(n525), .D(buffer[31]), .Q(_zyL288_tfiRv57[39]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[40] ( .G(n525), .D(buffer[16]), .Q(_zyL288_tfiRv57[40]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[41] ( .G(n525), .D(buffer[17]), .Q(_zyL288_tfiRv57[41]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[42] ( .G(n525), .D(buffer[18]), .Q(_zyL288_tfiRv57[42]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[43] ( .G(n525), .D(buffer[19]), .Q(_zyL288_tfiRv57[43]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[44] ( .G(n525), .D(buffer[20]), .Q(_zyL288_tfiRv57[44]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[45] ( .G(n525), .D(buffer[21]), .Q(_zyL288_tfiRv57[45]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[46] ( .G(n525), .D(buffer[22]), .Q(_zyL288_tfiRv57[46]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[47] ( .G(n525), .D(buffer[23]), .Q(_zyL288_tfiRv57[47]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[48] ( .G(n525), .D(buffer[8]), .Q(_zyL288_tfiRv57[48]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[49] ( .G(n525), .D(buffer[9]), .Q(_zyL288_tfiRv57[49]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[50] ( .G(n525), .D(buffer[10]), .Q(_zyL288_tfiRv57[50]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[51] ( .G(n525), .D(buffer[11]), .Q(_zyL288_tfiRv57[51]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[52] ( .G(n525), .D(buffer[12]), .Q(_zyL288_tfiRv57[52]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[53] ( .G(n525), .D(buffer[13]), .Q(_zyL288_tfiRv57[53]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[54] ( .G(n525), .D(buffer[14]), .Q(_zyL288_tfiRv57[54]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[55] ( .G(n525), .D(buffer[15]), .Q(_zyL288_tfiRv57[55]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[56] ( .G(n525), .D(buffer[0]), .Q(_zyL288_tfiRv57[56]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[57] ( .G(n525), .D(buffer[1]), .Q(_zyL288_tfiRv57[57]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[58] ( .G(n525), .D(buffer[2]), .Q(_zyL288_tfiRv57[58]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[59] ( .G(n525), .D(buffer[3]), .Q(_zyL288_tfiRv57[59]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[60] ( .G(n525), .D(buffer[4]), .Q(_zyL288_tfiRv57[60]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[61] ( .G(n525), .D(buffer[5]), .Q(_zyL288_tfiRv57[61]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[62] ( .G(n525), .D(buffer[6]), .Q(_zyL288_tfiRv57[62]), .QN( ));
Q_LDP0 \_zyL288_tfiRv57_REG[63] ( .G(n525), .D(buffer[7]), .Q(_zyL288_tfiRv57[63]), .QN( ));
Q_LDN0 _zyL255_tfiRv56_REG  ( .G(n530), .D(n176), .Q(_zyL255_tfiRv56), .QN( ));
Q_LDN0 _zyL254_tfiRv55_REG  ( .G(n530), .D(n1710), .Q(_zyL254_tfiRv55), .QN( ));
Q_LDN0 _zyL253_tfiRv54_REG  ( .G(n530), .D(n1712), .Q(_zyL253_tfiRv54), .QN( ));
Q_LDN0 _zyL252_tfiRv53_REG  ( .G(n530), .D(n177), .Q(_zyL252_tfiRv53), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[0] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[0]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[1] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[1]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[2] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[2]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[3] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[3]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[4] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[4]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[5] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[5]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[6] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[6]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[7] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[7]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[8] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[8]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[9] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[9]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[10] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[10]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[11] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[11]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[12] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[12]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[13] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[13]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[14] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[14]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[15] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[15]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[16] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[16]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[17] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[17]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[18] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[18]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[19] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[19]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[20] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[20]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[21] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[21]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[22] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[22]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[23] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[23]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[24] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[24]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[25] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[25]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[26] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[26]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[27] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[27]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[28] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[28]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[29] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[29]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[30] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[30]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[31] ( .G(n165), .D(n1735), .Q(_zyL234_tfiRv52[31]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[32] ( .G(n165), .D(buffer[24]), .Q(_zyL234_tfiRv52[32]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[33] ( .G(n165), .D(buffer[25]), .Q(_zyL234_tfiRv52[33]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[34] ( .G(n165), .D(buffer[26]), .Q(_zyL234_tfiRv52[34]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[35] ( .G(n165), .D(buffer[27]), .Q(_zyL234_tfiRv52[35]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[36] ( .G(n165), .D(buffer[28]), .Q(_zyL234_tfiRv52[36]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[37] ( .G(n165), .D(buffer[29]), .Q(_zyL234_tfiRv52[37]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[38] ( .G(n165), .D(buffer[30]), .Q(_zyL234_tfiRv52[38]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[39] ( .G(n165), .D(buffer[31]), .Q(_zyL234_tfiRv52[39]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[40] ( .G(n165), .D(buffer[16]), .Q(_zyL234_tfiRv52[40]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[41] ( .G(n165), .D(buffer[17]), .Q(_zyL234_tfiRv52[41]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[42] ( .G(n165), .D(buffer[18]), .Q(_zyL234_tfiRv52[42]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[43] ( .G(n165), .D(buffer[19]), .Q(_zyL234_tfiRv52[43]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[44] ( .G(n165), .D(buffer[20]), .Q(_zyL234_tfiRv52[44]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[45] ( .G(n165), .D(buffer[21]), .Q(_zyL234_tfiRv52[45]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[46] ( .G(n165), .D(buffer[22]), .Q(_zyL234_tfiRv52[46]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[47] ( .G(n165), .D(buffer[23]), .Q(_zyL234_tfiRv52[47]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[48] ( .G(n165), .D(buffer[8]), .Q(_zyL234_tfiRv52[48]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[49] ( .G(n165), .D(buffer[9]), .Q(_zyL234_tfiRv52[49]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[50] ( .G(n165), .D(buffer[10]), .Q(_zyL234_tfiRv52[50]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[51] ( .G(n165), .D(buffer[11]), .Q(_zyL234_tfiRv52[51]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[52] ( .G(n165), .D(buffer[12]), .Q(_zyL234_tfiRv52[52]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[53] ( .G(n165), .D(buffer[13]), .Q(_zyL234_tfiRv52[53]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[54] ( .G(n165), .D(buffer[14]), .Q(_zyL234_tfiRv52[54]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[55] ( .G(n165), .D(buffer[15]), .Q(_zyL234_tfiRv52[55]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[56] ( .G(n165), .D(buffer[0]), .Q(_zyL234_tfiRv52[56]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[57] ( .G(n165), .D(buffer[1]), .Q(_zyL234_tfiRv52[57]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[58] ( .G(n165), .D(buffer[2]), .Q(_zyL234_tfiRv52[58]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[59] ( .G(n165), .D(buffer[3]), .Q(_zyL234_tfiRv52[59]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[60] ( .G(n165), .D(buffer[4]), .Q(_zyL234_tfiRv52[60]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[61] ( .G(n165), .D(buffer[5]), .Q(_zyL234_tfiRv52[61]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[62] ( .G(n165), .D(buffer[6]), .Q(_zyL234_tfiRv52[62]), .QN( ));
Q_LDP0 \_zyL234_tfiRv52_REG[63] ( .G(n165), .D(buffer[7]), .Q(_zyL234_tfiRv52[63]), .QN( ));
Q_MX02 U2820 ( .S(n192), .A0(n733), .A1(n177), .Z(nxt_kme_internal_dek_kim_word[17]));
Q_AN02 U2821 ( .A0(n147), .A1(kme_internal_dek_kim_word[17]), .Z(n733));
Q_MX02 U2822 ( .S(n192), .A0(n734), .A1(n176), .Z(nxt_kme_internal_dak_kim_word[17]));
Q_AN02 U2823 ( .A0(n147), .A1(kme_internal_dak_kim_word[17]), .Z(n734));
Q_MX02 U2824 ( .S(n631), .A0(n174), .A1(n735), .Z(nxt_kme_internal_word0[45]));
Q_AN02 U2825 ( .A0(n169), .A1(kme_internal_word0[45]), .Z(n735));
Q_MX02 U2826 ( .S(n631), .A0(n175), .A1(n736), .Z(nxt_kme_internal_word0[46]));
Q_AN02 U2827 ( .A0(n169), .A1(kme_internal_word0[46]), .Z(n736));
Q_MX03 U2828 ( .S0(n566), .S1(n557), .A0(n742), .A1(n741), .A2(n737), .Z(fifo_in[63]));
Q_MX03 U2829 ( .S0(n172), .S1(n171), .A0(n738), .A1(n739), .A2(n740), .Z(n737));
Q_AN02 U2830 ( .A0(n173), .A1(debug_cmd[31]), .Z(n738));
Q_MX02 U2831 ( .S(n173), .A0(kme_internal_word0[63]), .A1(n1664), .Z(n739));
Q_MX04 U2832 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[63]), .A1(kme_internal_dek_kim_word[63]), .A2(iv1[63]), .A3(iv0[63]), .Z(n740));
Q_MX04 U2833 ( .S0(n173), .S1(n172), .A0(guid3[63]), .A1(guid2[63]), .A2(guid1[63]), .A3(guid0[63]), .Z(n741));
Q_MX02 U2834 ( .S(n172), .A0(stitcher_out[7]), .A1(buffer[7]), .Z(n742));
Q_MX03 U2835 ( .S0(n566), .S1(n557), .A0(n748), .A1(n747), .A2(n743), .Z(fifo_in[62]));
Q_MX03 U2836 ( .S0(n172), .S1(n171), .A0(n744), .A1(n745), .A2(n746), .Z(n743));
Q_AN02 U2837 ( .A0(n173), .A1(debug_cmd[30]), .Z(n744));
Q_MX02 U2838 ( .S(n173), .A0(kme_internal_word0[62]), .A1(n1665), .Z(n745));
Q_MX04 U2839 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[62]), .A1(kme_internal_dek_kim_word[62]), .A2(iv1[62]), .A3(iv0[62]), .Z(n746));
Q_MX04 U2840 ( .S0(n173), .S1(n172), .A0(guid3[62]), .A1(guid2[62]), .A2(guid1[62]), .A3(guid0[62]), .Z(n747));
Q_MX02 U2841 ( .S(n172), .A0(stitcher_out[6]), .A1(buffer[6]), .Z(n748));
Q_MX03 U2842 ( .S0(n566), .S1(n557), .A0(n754), .A1(n753), .A2(n749), .Z(fifo_in[61]));
Q_MX03 U2843 ( .S0(n172), .S1(n171), .A0(n750), .A1(n751), .A2(n752), .Z(n749));
Q_AN02 U2844 ( .A0(n173), .A1(debug_cmd[29]), .Z(n750));
Q_MX02 U2845 ( .S(n173), .A0(kme_internal_word0[61]), .A1(n1666), .Z(n751));
Q_MX04 U2846 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[61]), .A1(kme_internal_dek_kim_word[61]), .A2(iv1[61]), .A3(iv0[61]), .Z(n752));
Q_MX04 U2847 ( .S0(n173), .S1(n172), .A0(guid3[61]), .A1(guid2[61]), .A2(guid1[61]), .A3(guid0[61]), .Z(n753));
Q_MX02 U2848 ( .S(n172), .A0(stitcher_out[5]), .A1(buffer[5]), .Z(n754));
Q_MX03 U2849 ( .S0(n566), .S1(n557), .A0(n760), .A1(n759), .A2(n755), .Z(fifo_in[60]));
Q_MX03 U2850 ( .S0(n172), .S1(n171), .A0(n756), .A1(n757), .A2(n758), .Z(n755));
Q_AN02 U2851 ( .A0(n173), .A1(debug_cmd[28]), .Z(n756));
Q_MX02 U2852 ( .S(n173), .A0(kme_internal_word0[60]), .A1(n1667), .Z(n757));
Q_MX04 U2853 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[60]), .A1(kme_internal_dek_kim_word[60]), .A2(iv1[60]), .A3(iv0[60]), .Z(n758));
Q_MX04 U2854 ( .S0(n173), .S1(n172), .A0(guid3[60]), .A1(guid2[60]), .A2(guid1[60]), .A3(guid0[60]), .Z(n759));
Q_MX02 U2855 ( .S(n172), .A0(stitcher_out[4]), .A1(buffer[4]), .Z(n760));
Q_MX03 U2856 ( .S0(n566), .S1(n557), .A0(n766), .A1(n765), .A2(n761), .Z(fifo_in[59]));
Q_MX03 U2857 ( .S0(n172), .S1(n171), .A0(n762), .A1(n763), .A2(n764), .Z(n761));
Q_AN02 U2858 ( .A0(n173), .A1(debug_cmd[27]), .Z(n762));
Q_MX02 U2859 ( .S(n173), .A0(kme_internal_word0[59]), .A1(n1668), .Z(n763));
Q_MX04 U2860 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[59]), .A1(kme_internal_dek_kim_word[59]), .A2(iv1[59]), .A3(iv0[59]), .Z(n764));
Q_MX04 U2861 ( .S0(n173), .S1(n172), .A0(guid3[59]), .A1(guid2[59]), .A2(guid1[59]), .A3(guid0[59]), .Z(n765));
Q_MX02 U2862 ( .S(n172), .A0(stitcher_out[3]), .A1(buffer[3]), .Z(n766));
Q_MX03 U2863 ( .S0(n566), .S1(n557), .A0(n772), .A1(n771), .A2(n767), .Z(fifo_in[58]));
Q_MX03 U2864 ( .S0(n172), .S1(n171), .A0(n768), .A1(n769), .A2(n770), .Z(n767));
Q_AN02 U2865 ( .A0(n173), .A1(debug_cmd[26]), .Z(n768));
Q_MX02 U2866 ( .S(n173), .A0(kme_internal_word0[58]), .A1(n1669), .Z(n769));
Q_MX04 U2867 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[58]), .A1(kme_internal_dek_kim_word[58]), .A2(iv1[58]), .A3(iv0[58]), .Z(n770));
Q_MX04 U2868 ( .S0(n173), .S1(n172), .A0(guid3[58]), .A1(guid2[58]), .A2(guid1[58]), .A3(guid0[58]), .Z(n771));
Q_MX02 U2869 ( .S(n172), .A0(stitcher_out[2]), .A1(buffer[2]), .Z(n772));
Q_MX03 U2870 ( .S0(n566), .S1(n557), .A0(n778), .A1(n777), .A2(n773), .Z(fifo_in[57]));
Q_MX03 U2871 ( .S0(n172), .S1(n171), .A0(n774), .A1(n775), .A2(n776), .Z(n773));
Q_AN02 U2872 ( .A0(n173), .A1(debug_cmd[25]), .Z(n774));
Q_MX02 U2873 ( .S(n173), .A0(kme_internal_word0[57]), .A1(n1670), .Z(n775));
Q_MX04 U2874 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[57]), .A1(kme_internal_dek_kim_word[57]), .A2(iv1[57]), .A3(iv0[57]), .Z(n776));
Q_MX04 U2875 ( .S0(n173), .S1(n172), .A0(guid3[57]), .A1(guid2[57]), .A2(guid1[57]), .A3(guid0[57]), .Z(n777));
Q_MX02 U2876 ( .S(n172), .A0(stitcher_out[1]), .A1(buffer[1]), .Z(n778));
Q_MX03 U2877 ( .S0(n566), .S1(n557), .A0(n784), .A1(n783), .A2(n779), .Z(fifo_in[56]));
Q_MX03 U2878 ( .S0(n172), .S1(n171), .A0(n780), .A1(n781), .A2(n782), .Z(n779));
Q_AN02 U2879 ( .A0(n173), .A1(debug_cmd[24]), .Z(n780));
Q_MX02 U2880 ( .S(n173), .A0(kme_internal_word0[56]), .A1(n1671), .Z(n781));
Q_MX04 U2881 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[56]), .A1(kme_internal_dek_kim_word[56]), .A2(iv1[56]), .A3(iv0[56]), .Z(n782));
Q_MX04 U2882 ( .S0(n173), .S1(n172), .A0(guid3[56]), .A1(guid2[56]), .A2(guid1[56]), .A3(guid0[56]), .Z(n783));
Q_MX02 U2883 ( .S(n172), .A0(stitcher_out[0]), .A1(buffer[0]), .Z(n784));
Q_MX03 U2884 ( .S0(n566), .S1(n557), .A0(n790), .A1(n789), .A2(n785), .Z(fifo_in[55]));
Q_MX03 U2885 ( .S0(n172), .S1(n171), .A0(n786), .A1(n787), .A2(n788), .Z(n785));
Q_AN02 U2886 ( .A0(n173), .A1(debug_cmd[23]), .Z(n786));
Q_MX02 U2887 ( .S(n173), .A0(kme_internal_word0[55]), .A1(n1672), .Z(n787));
Q_MX04 U2888 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[55]), .A1(kme_internal_dek_kim_word[55]), .A2(iv1[55]), .A3(iv0[55]), .Z(n788));
Q_MX04 U2889 ( .S0(n173), .S1(n172), .A0(guid3[55]), .A1(guid2[55]), .A2(guid1[55]), .A3(guid0[55]), .Z(n789));
Q_MX02 U2890 ( .S(n172), .A0(stitcher_out[15]), .A1(buffer[15]), .Z(n790));
Q_MX03 U2891 ( .S0(n566), .S1(n557), .A0(n796), .A1(n795), .A2(n791), .Z(fifo_in[54]));
Q_MX03 U2892 ( .S0(n172), .S1(n171), .A0(n792), .A1(n793), .A2(n794), .Z(n791));
Q_AN02 U2893 ( .A0(n173), .A1(debug_cmd[22]), .Z(n792));
Q_MX02 U2894 ( .S(n173), .A0(kme_internal_word0[54]), .A1(n1673), .Z(n793));
Q_MX04 U2895 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[54]), .A1(kme_internal_dek_kim_word[54]), .A2(iv1[54]), .A3(iv0[54]), .Z(n794));
Q_MX04 U2896 ( .S0(n173), .S1(n172), .A0(guid3[54]), .A1(guid2[54]), .A2(guid1[54]), .A3(guid0[54]), .Z(n795));
Q_MX02 U2897 ( .S(n172), .A0(stitcher_out[14]), .A1(buffer[14]), .Z(n796));
Q_MX03 U2898 ( .S0(n566), .S1(n557), .A0(n802), .A1(n801), .A2(n797), .Z(fifo_in[53]));
Q_MX03 U2899 ( .S0(n172), .S1(n171), .A0(n798), .A1(n799), .A2(n800), .Z(n797));
Q_AN02 U2900 ( .A0(n173), .A1(debug_cmd[21]), .Z(n798));
Q_MX02 U2901 ( .S(n173), .A0(kme_internal_word0[53]), .A1(n1674), .Z(n799));
Q_MX04 U2902 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[53]), .A1(kme_internal_dek_kim_word[53]), .A2(iv1[53]), .A3(iv0[53]), .Z(n800));
Q_MX04 U2903 ( .S0(n173), .S1(n172), .A0(guid3[53]), .A1(guid2[53]), .A2(guid1[53]), .A3(guid0[53]), .Z(n801));
Q_MX02 U2904 ( .S(n172), .A0(stitcher_out[13]), .A1(buffer[13]), .Z(n802));
Q_MX03 U2905 ( .S0(n566), .S1(n557), .A0(n808), .A1(n807), .A2(n803), .Z(fifo_in[52]));
Q_MX03 U2906 ( .S0(n172), .S1(n171), .A0(n804), .A1(n805), .A2(n806), .Z(n803));
Q_AN02 U2907 ( .A0(n173), .A1(debug_cmd[20]), .Z(n804));
Q_MX02 U2908 ( .S(n173), .A0(kme_internal_word0[52]), .A1(n1675), .Z(n805));
Q_MX04 U2909 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[52]), .A1(kme_internal_dek_kim_word[52]), .A2(iv1[52]), .A3(iv0[52]), .Z(n806));
Q_MX04 U2910 ( .S0(n173), .S1(n172), .A0(guid3[52]), .A1(guid2[52]), .A2(guid1[52]), .A3(guid0[52]), .Z(n807));
Q_MX02 U2911 ( .S(n172), .A0(stitcher_out[12]), .A1(buffer[12]), .Z(n808));
Q_MX03 U2912 ( .S0(n566), .S1(n557), .A0(n814), .A1(n813), .A2(n809), .Z(fifo_in[51]));
Q_MX03 U2913 ( .S0(n172), .S1(n171), .A0(n810), .A1(n811), .A2(n812), .Z(n809));
Q_AN02 U2914 ( .A0(n173), .A1(debug_cmd[19]), .Z(n810));
Q_MX02 U2915 ( .S(n173), .A0(kme_internal_word0[51]), .A1(n1676), .Z(n811));
Q_MX04 U2916 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[51]), .A1(kme_internal_dek_kim_word[51]), .A2(iv1[51]), .A3(iv0[51]), .Z(n812));
Q_MX04 U2917 ( .S0(n173), .S1(n172), .A0(guid3[51]), .A1(guid2[51]), .A2(guid1[51]), .A3(guid0[51]), .Z(n813));
Q_MX02 U2918 ( .S(n172), .A0(stitcher_out[11]), .A1(buffer[11]), .Z(n814));
Q_MX03 U2919 ( .S0(n566), .S1(n557), .A0(n820), .A1(n819), .A2(n815), .Z(fifo_in[50]));
Q_MX03 U2920 ( .S0(n172), .S1(n171), .A0(n816), .A1(n817), .A2(n818), .Z(n815));
Q_AN02 U2921 ( .A0(n173), .A1(debug_cmd[18]), .Z(n816));
Q_MX02 U2922 ( .S(n173), .A0(kme_internal_word0[50]), .A1(n1677), .Z(n817));
Q_MX04 U2923 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[50]), .A1(kme_internal_dek_kim_word[50]), .A2(iv1[50]), .A3(iv0[50]), .Z(n818));
Q_MX04 U2924 ( .S0(n173), .S1(n172), .A0(guid3[50]), .A1(guid2[50]), .A2(guid1[50]), .A3(guid0[50]), .Z(n819));
Q_MX02 U2925 ( .S(n172), .A0(stitcher_out[10]), .A1(buffer[10]), .Z(n820));
Q_MX03 U2926 ( .S0(n566), .S1(n557), .A0(n826), .A1(n825), .A2(n821), .Z(fifo_in[49]));
Q_MX03 U2927 ( .S0(n172), .S1(n171), .A0(n822), .A1(n823), .A2(n824), .Z(n821));
Q_AN02 U2928 ( .A0(n173), .A1(debug_cmd[17]), .Z(n822));
Q_MX02 U2929 ( .S(n173), .A0(kme_internal_word0[49]), .A1(n1678), .Z(n823));
Q_MX04 U2930 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[49]), .A1(kme_internal_dek_kim_word[49]), .A2(iv1[49]), .A3(iv0[49]), .Z(n824));
Q_MX04 U2931 ( .S0(n173), .S1(n172), .A0(guid3[49]), .A1(guid2[49]), .A2(guid1[49]), .A3(guid0[49]), .Z(n825));
Q_MX02 U2932 ( .S(n172), .A0(stitcher_out[9]), .A1(buffer[9]), .Z(n826));
Q_MX03 U2933 ( .S0(n566), .S1(n557), .A0(n832), .A1(n831), .A2(n827), .Z(fifo_in[48]));
Q_MX03 U2934 ( .S0(n172), .S1(n171), .A0(n828), .A1(n829), .A2(n830), .Z(n827));
Q_AN02 U2935 ( .A0(n173), .A1(debug_cmd[16]), .Z(n828));
Q_MX02 U2936 ( .S(n173), .A0(n1707), .A1(n1679), .Z(n829));
Q_MX04 U2937 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[48]), .A1(kme_internal_dek_kim_word[48]), .A2(iv1[48]), .A3(iv0[48]), .Z(n830));
Q_MX04 U2938 ( .S0(n173), .S1(n172), .A0(guid3[48]), .A1(guid2[48]), .A2(guid1[48]), .A3(guid0[48]), .Z(n831));
Q_MX02 U2939 ( .S(n172), .A0(stitcher_out[8]), .A1(buffer[8]), .Z(n832));
Q_MX03 U2940 ( .S0(n566), .S1(n557), .A0(n838), .A1(n837), .A2(n833), .Z(fifo_in[47]));
Q_MX03 U2941 ( .S0(n172), .S1(n171), .A0(n834), .A1(n835), .A2(n836), .Z(n833));
Q_AN02 U2942 ( .A0(n173), .A1(debug_cmd[15]), .Z(n834));
Q_MX02 U2943 ( .S(n173), .A0(n1696), .A1(n1680), .Z(n835));
Q_MX04 U2944 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[47]), .A1(kme_internal_dek_kim_word[47]), .A2(iv1[47]), .A3(iv0[47]), .Z(n836));
Q_MX04 U2945 ( .S0(n173), .S1(n172), .A0(guid3[47]), .A1(guid2[47]), .A2(guid1[47]), .A3(guid0[47]), .Z(n837));
Q_MX02 U2946 ( .S(n172), .A0(stitcher_out[23]), .A1(buffer[23]), .Z(n838));
Q_MX03 U2947 ( .S0(n566), .S1(n557), .A0(n844), .A1(n843), .A2(n839), .Z(fifo_in[46]));
Q_MX03 U2948 ( .S0(n172), .S1(n171), .A0(n840), .A1(n841), .A2(n842), .Z(n839));
Q_AN02 U2949 ( .A0(n173), .A1(debug_cmd[14]), .Z(n840));
Q_MX02 U2950 ( .S(n173), .A0(n175), .A1(n1681), .Z(n841));
Q_MX04 U2951 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[46]), .A1(kme_internal_dek_kim_word[46]), .A2(iv1[46]), .A3(iv0[46]), .Z(n842));
Q_MX04 U2952 ( .S0(n173), .S1(n172), .A0(guid3[46]), .A1(guid2[46]), .A2(guid1[46]), .A3(guid0[46]), .Z(n843));
Q_MX02 U2953 ( .S(n172), .A0(stitcher_out[22]), .A1(buffer[22]), .Z(n844));
Q_MX03 U2954 ( .S0(n566), .S1(n557), .A0(n850), .A1(n849), .A2(n845), .Z(fifo_in[45]));
Q_MX03 U2955 ( .S0(n172), .S1(n171), .A0(n846), .A1(n847), .A2(n848), .Z(n845));
Q_AN02 U2956 ( .A0(n173), .A1(debug_cmd[13]), .Z(n846));
Q_MX02 U2957 ( .S(n173), .A0(n174), .A1(n1682), .Z(n847));
Q_MX04 U2958 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[45]), .A1(kme_internal_dek_kim_word[45]), .A2(iv1[45]), .A3(iv0[45]), .Z(n848));
Q_MX04 U2959 ( .S0(n173), .S1(n172), .A0(guid3[45]), .A1(guid2[45]), .A2(guid1[45]), .A3(guid0[45]), .Z(n849));
Q_MX02 U2960 ( .S(n172), .A0(stitcher_out[21]), .A1(buffer[21]), .Z(n850));
Q_MX03 U2961 ( .S0(n566), .S1(n557), .A0(n856), .A1(n855), .A2(n851), .Z(fifo_in[44]));
Q_MX03 U2962 ( .S0(n172), .S1(n171), .A0(n852), .A1(n853), .A2(n854), .Z(n851));
Q_AN02 U2963 ( .A0(n173), .A1(debug_cmd[12]), .Z(n852));
Q_MX02 U2964 ( .S(n173), .A0(stitcher_out[62]), .A1(n1683), .Z(n853));
Q_MX04 U2965 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[44]), .A1(kme_internal_dek_kim_word[44]), .A2(iv1[44]), .A3(iv0[44]), .Z(n854));
Q_MX04 U2966 ( .S0(n173), .S1(n172), .A0(guid3[44]), .A1(guid2[44]), .A2(guid1[44]), .A3(guid0[44]), .Z(n855));
Q_MX02 U2967 ( .S(n172), .A0(stitcher_out[20]), .A1(buffer[20]), .Z(n856));
Q_MX03 U2968 ( .S0(n566), .S1(n557), .A0(n862), .A1(n861), .A2(n857), .Z(fifo_in[43]));
Q_MX03 U2969 ( .S0(n172), .S1(n171), .A0(n858), .A1(n859), .A2(n860), .Z(n857));
Q_AN02 U2970 ( .A0(n173), .A1(debug_cmd[11]), .Z(n858));
Q_MX02 U2971 ( .S(n173), .A0(stitcher_out[61]), .A1(n1684), .Z(n859));
Q_MX04 U2972 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[43]), .A1(kme_internal_dek_kim_word[43]), .A2(iv1[43]), .A3(iv0[43]), .Z(n860));
Q_MX04 U2973 ( .S0(n173), .S1(n172), .A0(guid3[43]), .A1(guid2[43]), .A2(guid1[43]), .A3(guid0[43]), .Z(n861));
Q_MX02 U2974 ( .S(n172), .A0(stitcher_out[19]), .A1(buffer[19]), .Z(n862));
Q_MX03 U2975 ( .S0(n566), .S1(n557), .A0(n868), .A1(n867), .A2(n863), .Z(fifo_in[42]));
Q_MX03 U2976 ( .S0(n172), .S1(n171), .A0(n864), .A1(n865), .A2(n866), .Z(n863));
Q_AN02 U2977 ( .A0(n173), .A1(debug_cmd[10]), .Z(n864));
Q_MX02 U2978 ( .S(n173), .A0(stitcher_out[60]), .A1(n1685), .Z(n865));
Q_MX04 U2979 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[42]), .A1(kme_internal_dek_kim_word[42]), .A2(iv1[42]), .A3(iv0[42]), .Z(n866));
Q_MX04 U2980 ( .S0(n173), .S1(n172), .A0(guid3[42]), .A1(guid2[42]), .A2(guid1[42]), .A3(guid0[42]), .Z(n867));
Q_MX02 U2981 ( .S(n172), .A0(stitcher_out[18]), .A1(buffer[18]), .Z(n868));
Q_MX03 U2982 ( .S0(n566), .S1(n557), .A0(n874), .A1(n873), .A2(n869), .Z(fifo_in[41]));
Q_MX03 U2983 ( .S0(n172), .S1(n171), .A0(n870), .A1(n871), .A2(n872), .Z(n869));
Q_AN02 U2984 ( .A0(n173), .A1(debug_cmd[9]), .Z(n870));
Q_MX02 U2985 ( .S(n173), .A0(stitcher_out[59]), .A1(n1686), .Z(n871));
Q_MX04 U2986 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[41]), .A1(kme_internal_dek_kim_word[41]), .A2(iv1[41]), .A3(iv0[41]), .Z(n872));
Q_MX04 U2987 ( .S0(n173), .S1(n172), .A0(guid3[41]), .A1(guid2[41]), .A2(guid1[41]), .A3(guid0[41]), .Z(n873));
Q_MX02 U2988 ( .S(n172), .A0(stitcher_out[17]), .A1(buffer[17]), .Z(n874));
Q_MX03 U2989 ( .S0(n566), .S1(n557), .A0(n880), .A1(n879), .A2(n875), .Z(fifo_in[40]));
Q_MX03 U2990 ( .S0(n172), .S1(n171), .A0(n876), .A1(n877), .A2(n878), .Z(n875));
Q_AN02 U2991 ( .A0(n173), .A1(debug_cmd[8]), .Z(n876));
Q_MX02 U2992 ( .S(n173), .A0(stitcher_out[58]), .A1(n1687), .Z(n877));
Q_MX04 U2993 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[40]), .A1(kme_internal_dek_kim_word[40]), .A2(iv1[40]), .A3(iv0[40]), .Z(n878));
Q_MX04 U2994 ( .S0(n173), .S1(n172), .A0(guid3[40]), .A1(guid2[40]), .A2(guid1[40]), .A3(guid0[40]), .Z(n879));
Q_MX02 U2995 ( .S(n172), .A0(stitcher_out[16]), .A1(buffer[16]), .Z(n880));
Q_MX03 U2996 ( .S0(n566), .S1(n557), .A0(n886), .A1(n885), .A2(n881), .Z(fifo_in[39]));
Q_MX03 U2997 ( .S0(n172), .S1(n171), .A0(n882), .A1(n883), .A2(n884), .Z(n881));
Q_AN02 U2998 ( .A0(n173), .A1(debug_cmd[7]), .Z(n882));
Q_MX02 U2999 ( .S(n173), .A0(stitcher_out[57]), .A1(n1688), .Z(n883));
Q_MX04 U3000 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[39]), .A1(kme_internal_dek_kim_word[39]), .A2(iv1[39]), .A3(iv0[39]), .Z(n884));
Q_MX04 U3001 ( .S0(n173), .S1(n172), .A0(guid3[39]), .A1(guid2[39]), .A2(guid1[39]), .A3(guid0[39]), .Z(n885));
Q_MX02 U3002 ( .S(n172), .A0(stitcher_out[31]), .A1(buffer[31]), .Z(n886));
Q_MX03 U3003 ( .S0(n566), .S1(n557), .A0(n892), .A1(n891), .A2(n887), .Z(fifo_in[38]));
Q_MX03 U3004 ( .S0(n172), .S1(n171), .A0(n888), .A1(n889), .A2(n890), .Z(n887));
Q_AN02 U3005 ( .A0(n173), .A1(debug_cmd[6]), .Z(n888));
Q_MX02 U3006 ( .S(n173), .A0(kme_internal_word0[38]), .A1(n1689), .Z(n889));
Q_MX04 U3007 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[38]), .A1(kme_internal_dek_kim_word[38]), .A2(iv1[38]), .A3(iv0[38]), .Z(n890));
Q_MX04 U3008 ( .S0(n173), .S1(n172), .A0(guid3[38]), .A1(guid2[38]), .A2(guid1[38]), .A3(guid0[38]), .Z(n891));
Q_MX02 U3009 ( .S(n172), .A0(stitcher_out[30]), .A1(buffer[30]), .Z(n892));
Q_MX03 U3010 ( .S0(n566), .S1(n557), .A0(n898), .A1(n897), .A2(n893), .Z(fifo_in[37]));
Q_MX03 U3011 ( .S0(n172), .S1(n171), .A0(n894), .A1(n895), .A2(n896), .Z(n893));
Q_AN02 U3012 ( .A0(n173), .A1(debug_cmd[5]), .Z(n894));
Q_MX02 U3013 ( .S(n173), .A0(kme_internal_word0[37]), .A1(n1690), .Z(n895));
Q_MX04 U3014 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[37]), .A1(kme_internal_dek_kim_word[37]), .A2(iv1[37]), .A3(iv0[37]), .Z(n896));
Q_MX04 U3015 ( .S0(n173), .S1(n172), .A0(guid3[37]), .A1(guid2[37]), .A2(guid1[37]), .A3(guid0[37]), .Z(n897));
Q_MX02 U3016 ( .S(n172), .A0(stitcher_out[29]), .A1(buffer[29]), .Z(n898));
Q_MX03 U3017 ( .S0(n566), .S1(n557), .A0(n904), .A1(n903), .A2(n899), .Z(fifo_in[36]));
Q_MX03 U3018 ( .S0(n172), .S1(n171), .A0(n900), .A1(n901), .A2(n902), .Z(n899));
Q_AN02 U3019 ( .A0(n173), .A1(debug_cmd[4]), .Z(n900));
Q_MX02 U3020 ( .S(n173), .A0(kme_internal_word0[36]), .A1(n1691), .Z(n901));
Q_MX04 U3021 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[36]), .A1(kme_internal_dek_kim_word[36]), .A2(iv1[36]), .A3(iv0[36]), .Z(n902));
Q_MX04 U3022 ( .S0(n173), .S1(n172), .A0(guid3[36]), .A1(guid2[36]), .A2(guid1[36]), .A3(guid0[36]), .Z(n903));
Q_MX02 U3023 ( .S(n172), .A0(stitcher_out[28]), .A1(buffer[28]), .Z(n904));
Q_MX03 U3024 ( .S0(n566), .S1(n557), .A0(n910), .A1(n909), .A2(n905), .Z(fifo_in[35]));
Q_MX03 U3025 ( .S0(n172), .S1(n171), .A0(n906), .A1(n907), .A2(n908), .Z(n905));
Q_AN02 U3026 ( .A0(n173), .A1(debug_cmd[3]), .Z(n906));
Q_MX02 U3027 ( .S(n173), .A0(kme_internal_word0[35]), .A1(n1692), .Z(n907));
Q_MX04 U3028 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[35]), .A1(kme_internal_dek_kim_word[35]), .A2(iv1[35]), .A3(iv0[35]), .Z(n908));
Q_MX04 U3029 ( .S0(n173), .S1(n172), .A0(guid3[35]), .A1(guid2[35]), .A2(guid1[35]), .A3(guid0[35]), .Z(n909));
Q_MX02 U3030 ( .S(n172), .A0(stitcher_out[27]), .A1(buffer[27]), .Z(n910));
Q_MX03 U3031 ( .S0(n566), .S1(n557), .A0(n916), .A1(n915), .A2(n911), .Z(fifo_in[34]));
Q_MX03 U3032 ( .S0(n172), .S1(n171), .A0(n912), .A1(n913), .A2(n914), .Z(n911));
Q_AN02 U3033 ( .A0(n173), .A1(debug_cmd[2]), .Z(n912));
Q_MX02 U3034 ( .S(n173), .A0(kme_internal_word0[34]), .A1(n1693), .Z(n913));
Q_MX04 U3035 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[34]), .A1(kme_internal_dek_kim_word[34]), .A2(iv1[34]), .A3(iv0[34]), .Z(n914));
Q_MX04 U3036 ( .S0(n173), .S1(n172), .A0(guid3[34]), .A1(guid2[34]), .A2(guid1[34]), .A3(guid0[34]), .Z(n915));
Q_MX02 U3037 ( .S(n172), .A0(stitcher_out[26]), .A1(buffer[26]), .Z(n916));
Q_MX03 U3038 ( .S0(n566), .S1(n557), .A0(n922), .A1(n921), .A2(n917), .Z(fifo_in[33]));
Q_MX03 U3039 ( .S0(n172), .S1(n171), .A0(n918), .A1(n919), .A2(n920), .Z(n917));
Q_AN02 U3040 ( .A0(n173), .A1(debug_cmd[1]), .Z(n918));
Q_MX02 U3041 ( .S(n173), .A0(kme_internal_word0[33]), .A1(n1694), .Z(n919));
Q_MX04 U3042 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[33]), .A1(kme_internal_dek_kim_word[33]), .A2(iv1[33]), .A3(iv0[33]), .Z(n920));
Q_MX04 U3043 ( .S0(n173), .S1(n172), .A0(guid3[33]), .A1(guid2[33]), .A2(guid1[33]), .A3(guid0[33]), .Z(n921));
Q_MX02 U3044 ( .S(n172), .A0(stitcher_out[25]), .A1(buffer[25]), .Z(n922));
Q_MX03 U3045 ( .S0(n566), .S1(n557), .A0(n928), .A1(n927), .A2(n923), .Z(fifo_in[32]));
Q_MX03 U3046 ( .S0(n172), .S1(n171), .A0(n924), .A1(n925), .A2(n926), .Z(n923));
Q_AN02 U3047 ( .A0(n173), .A1(debug_cmd[0]), .Z(n924));
Q_MX02 U3048 ( .S(n173), .A0(kme_internal_word0[32]), .A1(n1695), .Z(n925));
Q_MX04 U3049 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[32]), .A1(kme_internal_dek_kim_word[32]), .A2(iv1[32]), .A3(iv0[32]), .Z(n926));
Q_MX04 U3050 ( .S0(n173), .S1(n172), .A0(guid3[32]), .A1(guid2[32]), .A2(guid1[32]), .A3(guid0[32]), .Z(n927));
Q_MX02 U3051 ( .S(n172), .A0(stitcher_out[24]), .A1(buffer[24]), .Z(n928));
Q_MX03 U3052 ( .S0(n566), .S1(n557), .A0(n934), .A1(n933), .A2(n929), .Z(fifo_in[31]));
Q_MX03 U3053 ( .S0(n172), .S1(n171), .A0(n930), .A1(n931), .A2(n932), .Z(n929));
Q_AN02 U3054 ( .A0(n173), .A1(stitcher_out[31]), .Z(n930));
Q_AN02 U3055 ( .A0(n1153), .A1(kme_internal_word0[31]), .Z(n931));
Q_MX04 U3056 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[31]), .A1(kme_internal_dek_kim_word[31]), .A2(iv1[31]), .A3(iv0[31]), .Z(n932));
Q_MX04 U3057 ( .S0(n173), .S1(n172), .A0(guid3[31]), .A1(guid2[31]), .A2(guid1[31]), .A3(guid0[31]), .Z(n933));
Q_MX02 U3058 ( .S(n172), .A0(n935), .A1(stitcher_out[7]), .Z(n934));
Q_AN02 U3059 ( .A0(n1153), .A1(stitcher_out[39]), .Z(n935));
Q_MX03 U3060 ( .S0(n566), .S1(n557), .A0(n941), .A1(n940), .A2(n936), .Z(fifo_in[30]));
Q_MX03 U3061 ( .S0(n172), .S1(n171), .A0(n937), .A1(n938), .A2(n939), .Z(n936));
Q_AN02 U3062 ( .A0(n173), .A1(stitcher_out[30]), .Z(n937));
Q_AN02 U3063 ( .A0(n1153), .A1(kme_internal_word0[30]), .Z(n938));
Q_MX04 U3064 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[30]), .A1(kme_internal_dek_kim_word[30]), .A2(iv1[30]), .A3(iv0[30]), .Z(n939));
Q_MX04 U3065 ( .S0(n173), .S1(n172), .A0(guid3[30]), .A1(guid2[30]), .A2(guid1[30]), .A3(guid0[30]), .Z(n940));
Q_MX02 U3066 ( .S(n172), .A0(n942), .A1(stitcher_out[6]), .Z(n941));
Q_AN02 U3067 ( .A0(n1153), .A1(stitcher_out[38]), .Z(n942));
Q_MX03 U3068 ( .S0(n566), .S1(n557), .A0(n948), .A1(n947), .A2(n943), .Z(fifo_in[29]));
Q_MX03 U3069 ( .S0(n172), .S1(n171), .A0(n944), .A1(n945), .A2(n946), .Z(n943));
Q_AN02 U3070 ( .A0(n173), .A1(stitcher_out[29]), .Z(n944));
Q_AN02 U3071 ( .A0(n1153), .A1(kme_internal_word0[29]), .Z(n945));
Q_MX04 U3072 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[29]), .A1(kme_internal_dek_kim_word[29]), .A2(iv1[29]), .A3(iv0[29]), .Z(n946));
Q_MX04 U3073 ( .S0(n173), .S1(n172), .A0(guid3[29]), .A1(guid2[29]), .A2(guid1[29]), .A3(guid0[29]), .Z(n947));
Q_MX02 U3074 ( .S(n172), .A0(n949), .A1(stitcher_out[5]), .Z(n948));
Q_AN02 U3075 ( .A0(n1153), .A1(stitcher_out[37]), .Z(n949));
Q_MX03 U3076 ( .S0(n566), .S1(n557), .A0(n955), .A1(n954), .A2(n950), .Z(fifo_in[28]));
Q_MX03 U3077 ( .S0(n172), .S1(n171), .A0(n951), .A1(n952), .A2(n953), .Z(n950));
Q_AN02 U3078 ( .A0(n173), .A1(stitcher_out[28]), .Z(n951));
Q_AN02 U3079 ( .A0(n1153), .A1(kme_internal_word0[28]), .Z(n952));
Q_MX04 U3080 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[28]), .A1(kme_internal_dek_kim_word[28]), .A2(iv1[28]), .A3(iv0[28]), .Z(n953));
Q_MX04 U3081 ( .S0(n173), .S1(n172), .A0(guid3[28]), .A1(guid2[28]), .A2(guid1[28]), .A3(guid0[28]), .Z(n954));
Q_MX02 U3082 ( .S(n172), .A0(n956), .A1(stitcher_out[4]), .Z(n955));
Q_AN02 U3083 ( .A0(n1153), .A1(stitcher_out[36]), .Z(n956));
Q_MX03 U3084 ( .S0(n566), .S1(n557), .A0(n962), .A1(n961), .A2(n957), .Z(fifo_in[27]));
Q_MX03 U3085 ( .S0(n172), .S1(n171), .A0(n958), .A1(n959), .A2(n960), .Z(n957));
Q_AN02 U3086 ( .A0(n173), .A1(stitcher_out[27]), .Z(n958));
Q_AN02 U3087 ( .A0(n1153), .A1(kme_internal_word0[27]), .Z(n959));
Q_MX04 U3088 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[27]), .A1(kme_internal_dek_kim_word[27]), .A2(iv1[27]), .A3(iv0[27]), .Z(n960));
Q_MX04 U3089 ( .S0(n173), .S1(n172), .A0(guid3[27]), .A1(guid2[27]), .A2(guid1[27]), .A3(guid0[27]), .Z(n961));
Q_MX02 U3090 ( .S(n172), .A0(n963), .A1(stitcher_out[3]), .Z(n962));
Q_AN02 U3091 ( .A0(n1153), .A1(stitcher_out[35]), .Z(n963));
Q_MX03 U3092 ( .S0(n566), .S1(n557), .A0(n969), .A1(n968), .A2(n964), .Z(fifo_in[26]));
Q_MX03 U3093 ( .S0(n172), .S1(n171), .A0(n965), .A1(n966), .A2(n967), .Z(n964));
Q_AN02 U3094 ( .A0(n173), .A1(stitcher_out[26]), .Z(n965));
Q_AN02 U3095 ( .A0(n1153), .A1(kme_internal_word0[26]), .Z(n966));
Q_MX04 U3096 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[26]), .A1(kme_internal_dek_kim_word[26]), .A2(iv1[26]), .A3(iv0[26]), .Z(n967));
Q_MX04 U3097 ( .S0(n173), .S1(n172), .A0(guid3[26]), .A1(guid2[26]), .A2(guid1[26]), .A3(guid0[26]), .Z(n968));
Q_MX02 U3098 ( .S(n172), .A0(n970), .A1(stitcher_out[2]), .Z(n969));
Q_AN02 U3099 ( .A0(n1153), .A1(stitcher_out[34]), .Z(n970));
Q_MX03 U3100 ( .S0(n566), .S1(n557), .A0(n976), .A1(n975), .A2(n971), .Z(fifo_in[25]));
Q_MX03 U3101 ( .S0(n172), .S1(n171), .A0(n972), .A1(n973), .A2(n974), .Z(n971));
Q_AN02 U3102 ( .A0(n173), .A1(stitcher_out[25]), .Z(n972));
Q_AN02 U3103 ( .A0(n1153), .A1(kme_internal_word0[25]), .Z(n973));
Q_MX04 U3104 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[25]), .A1(kme_internal_dek_kim_word[25]), .A2(iv1[25]), .A3(iv0[25]), .Z(n974));
Q_MX04 U3105 ( .S0(n173), .S1(n172), .A0(guid3[25]), .A1(guid2[25]), .A2(guid1[25]), .A3(guid0[25]), .Z(n975));
Q_MX02 U3106 ( .S(n172), .A0(n977), .A1(stitcher_out[1]), .Z(n976));
Q_AN02 U3107 ( .A0(n1153), .A1(stitcher_out[33]), .Z(n977));
Q_MX03 U3108 ( .S0(n566), .S1(n557), .A0(n983), .A1(n982), .A2(n978), .Z(fifo_in[24]));
Q_MX03 U3109 ( .S0(n172), .S1(n171), .A0(n979), .A1(n980), .A2(n981), .Z(n978));
Q_AN02 U3110 ( .A0(n173), .A1(stitcher_out[24]), .Z(n979));
Q_AN02 U3111 ( .A0(n1153), .A1(kme_internal_word0[24]), .Z(n980));
Q_MX04 U3112 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[24]), .A1(kme_internal_dek_kim_word[24]), .A2(iv1[24]), .A3(iv0[24]), .Z(n981));
Q_MX04 U3113 ( .S0(n173), .S1(n172), .A0(guid3[24]), .A1(guid2[24]), .A2(guid1[24]), .A3(guid0[24]), .Z(n982));
Q_MX02 U3114 ( .S(n172), .A0(n984), .A1(stitcher_out[0]), .Z(n983));
Q_AN02 U3115 ( .A0(n1153), .A1(stitcher_out[32]), .Z(n984));
Q_MX03 U3116 ( .S0(n566), .S1(n557), .A0(n990), .A1(n989), .A2(n985), .Z(fifo_in[23]));
Q_MX03 U3117 ( .S0(n172), .S1(n171), .A0(n986), .A1(n987), .A2(n988), .Z(n985));
Q_AN02 U3118 ( .A0(n173), .A1(stitcher_out[23]), .Z(n986));
Q_AN02 U3119 ( .A0(n1153), .A1(kme_internal_word0[23]), .Z(n987));
Q_MX04 U3120 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[23]), .A1(kme_internal_dek_kim_word[23]), .A2(iv1[23]), .A3(iv0[23]), .Z(n988));
Q_MX04 U3121 ( .S0(n173), .S1(n172), .A0(guid3[23]), .A1(guid2[23]), .A2(guid1[23]), .A3(guid0[23]), .Z(n989));
Q_MX02 U3122 ( .S(n172), .A0(n991), .A1(stitcher_out[15]), .Z(n990));
Q_AN02 U3123 ( .A0(n1153), .A1(stitcher_out[47]), .Z(n991));
Q_MX03 U3124 ( .S0(n566), .S1(n557), .A0(n997), .A1(n996), .A2(n992), .Z(fifo_in[22]));
Q_MX03 U3125 ( .S0(n172), .S1(n171), .A0(n993), .A1(n994), .A2(n995), .Z(n992));
Q_AN02 U3126 ( .A0(n173), .A1(stitcher_out[22]), .Z(n993));
Q_AN02 U3127 ( .A0(n1153), .A1(kme_internal_word0[22]), .Z(n994));
Q_MX04 U3128 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[22]), .A1(kme_internal_dek_kim_word[22]), .A2(iv1[22]), .A3(iv0[22]), .Z(n995));
Q_MX04 U3129 ( .S0(n173), .S1(n172), .A0(guid3[22]), .A1(guid2[22]), .A2(guid1[22]), .A3(guid0[22]), .Z(n996));
Q_MX02 U3130 ( .S(n172), .A0(n998), .A1(stitcher_out[14]), .Z(n997));
Q_AN02 U3131 ( .A0(n1153), .A1(stitcher_out[46]), .Z(n998));
Q_MX03 U3132 ( .S0(n566), .S1(n557), .A0(n1004), .A1(n1003), .A2(n999), .Z(fifo_in[21]));
Q_MX03 U3133 ( .S0(n172), .S1(n171), .A0(n1000), .A1(n1001), .A2(n1002), .Z(n999));
Q_AN02 U3134 ( .A0(n173), .A1(stitcher_out[21]), .Z(n1000));
Q_AN02 U3135 ( .A0(n1153), .A1(kme_internal_word0[21]), .Z(n1001));
Q_MX04 U3136 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[21]), .A1(kme_internal_dek_kim_word[21]), .A2(iv1[21]), .A3(iv0[21]), .Z(n1002));
Q_MX04 U3137 ( .S0(n173), .S1(n172), .A0(guid3[21]), .A1(guid2[21]), .A2(guid1[21]), .A3(guid0[21]), .Z(n1003));
Q_MX02 U3138 ( .S(n172), .A0(n1005), .A1(stitcher_out[13]), .Z(n1004));
Q_AN02 U3139 ( .A0(n1153), .A1(stitcher_out[45]), .Z(n1005));
Q_MX03 U3140 ( .S0(n566), .S1(n557), .A0(n1011), .A1(n1010), .A2(n1006), .Z(fifo_in[20]));
Q_MX03 U3141 ( .S0(n172), .S1(n171), .A0(n1007), .A1(n1008), .A2(n1009), .Z(n1006));
Q_AN02 U3142 ( .A0(n173), .A1(stitcher_out[20]), .Z(n1007));
Q_AN02 U3143 ( .A0(n1153), .A1(kme_internal_word0[20]), .Z(n1008));
Q_MX04 U3144 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[20]), .A1(kme_internal_dek_kim_word[20]), .A2(iv1[20]), .A3(iv0[20]), .Z(n1009));
Q_MX04 U3145 ( .S0(n173), .S1(n172), .A0(guid3[20]), .A1(guid2[20]), .A2(guid1[20]), .A3(guid0[20]), .Z(n1010));
Q_MX02 U3146 ( .S(n172), .A0(n1012), .A1(stitcher_out[12]), .Z(n1011));
Q_AN02 U3147 ( .A0(n1153), .A1(stitcher_out[44]), .Z(n1012));
Q_MX03 U3148 ( .S0(n566), .S1(n557), .A0(n1018), .A1(n1017), .A2(n1013), .Z(fifo_in[19]));
Q_MX03 U3149 ( .S0(n172), .S1(n171), .A0(n1014), .A1(n1015), .A2(n1016), .Z(n1013));
Q_AN02 U3150 ( .A0(n173), .A1(stitcher_out[19]), .Z(n1014));
Q_AN02 U3151 ( .A0(n1153), .A1(kme_internal_word0[19]), .Z(n1015));
Q_MX04 U3152 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[19]), .A1(kme_internal_dek_kim_word[19]), .A2(iv1[19]), .A3(iv0[19]), .Z(n1016));
Q_MX04 U3153 ( .S0(n173), .S1(n172), .A0(guid3[19]), .A1(guid2[19]), .A2(guid1[19]), .A3(guid0[19]), .Z(n1017));
Q_MX02 U3154 ( .S(n172), .A0(n1019), .A1(stitcher_out[11]), .Z(n1018));
Q_AN02 U3155 ( .A0(n1153), .A1(stitcher_out[43]), .Z(n1019));
Q_MX03 U3156 ( .S0(n566), .S1(n557), .A0(n1025), .A1(n1024), .A2(n1020), .Z(fifo_in[18]));
Q_MX03 U3157 ( .S0(n172), .S1(n171), .A0(n1021), .A1(n1022), .A2(n1023), .Z(n1020));
Q_AN02 U3158 ( .A0(n173), .A1(stitcher_out[18]), .Z(n1021));
Q_AN02 U3159 ( .A0(n1153), .A1(kme_internal_word0[18]), .Z(n1022));
Q_MX04 U3160 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[18]), .A1(kme_internal_dek_kim_word[18]), .A2(iv1[18]), .A3(iv0[18]), .Z(n1023));
Q_MX04 U3161 ( .S0(n173), .S1(n172), .A0(guid3[18]), .A1(guid2[18]), .A2(guid1[18]), .A3(guid0[18]), .Z(n1024));
Q_MX02 U3162 ( .S(n172), .A0(n1026), .A1(stitcher_out[10]), .Z(n1025));
Q_AN02 U3163 ( .A0(n1153), .A1(stitcher_out[42]), .Z(n1026));
Q_MX03 U3164 ( .S0(n566), .S1(n557), .A0(n1032), .A1(n1031), .A2(n1027), .Z(fifo_in[17]));
Q_MX03 U3165 ( .S0(n172), .S1(n171), .A0(n1028), .A1(n1029), .A2(n1030), .Z(n1027));
Q_AN02 U3166 ( .A0(n173), .A1(stitcher_out[17]), .Z(n1028));
Q_AN02 U3167 ( .A0(n1153), .A1(kme_internal_word0[17]), .Z(n1029));
Q_MX04 U3168 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[17]), .A1(kme_internal_dek_kim_word[17]), .A2(iv1[17]), .A3(iv0[17]), .Z(n1030));
Q_MX04 U3169 ( .S0(n173), .S1(n172), .A0(guid3[17]), .A1(guid2[17]), .A2(guid1[17]), .A3(guid0[17]), .Z(n1031));
Q_MX02 U3170 ( .S(n172), .A0(n1033), .A1(stitcher_out[9]), .Z(n1032));
Q_AN02 U3171 ( .A0(n1153), .A1(stitcher_out[41]), .Z(n1033));
Q_MX03 U3172 ( .S0(n566), .S1(n557), .A0(n1039), .A1(n1038), .A2(n1034), .Z(fifo_in[16]));
Q_MX03 U3173 ( .S0(n172), .S1(n171), .A0(n1035), .A1(n1036), .A2(n1037), .Z(n1034));
Q_AN02 U3174 ( .A0(n173), .A1(stitcher_out[16]), .Z(n1035));
Q_AN02 U3175 ( .A0(n1153), .A1(kme_internal_word0[16]), .Z(n1036));
Q_MX04 U3176 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[16]), .A1(kme_internal_dek_kim_word[16]), .A2(iv1[16]), .A3(iv0[16]), .Z(n1037));
Q_MX04 U3177 ( .S0(n173), .S1(n172), .A0(guid3[16]), .A1(guid2[16]), .A2(guid1[16]), .A3(guid0[16]), .Z(n1038));
Q_MX02 U3178 ( .S(n172), .A0(n1040), .A1(stitcher_out[8]), .Z(n1039));
Q_AN02 U3179 ( .A0(n1153), .A1(stitcher_out[40]), .Z(n1040));
Q_MX03 U3180 ( .S0(n566), .S1(n557), .A0(n1046), .A1(n1045), .A2(n1041), .Z(fifo_in[15]));
Q_MX03 U3181 ( .S0(n172), .S1(n171), .A0(n1042), .A1(n1043), .A2(n1044), .Z(n1041));
Q_AN02 U3182 ( .A0(n173), .A1(stitcher_out[15]), .Z(n1042));
Q_AN02 U3183 ( .A0(n1153), .A1(kme_internal_word0[15]), .Z(n1043));
Q_MX04 U3184 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[15]), .A1(kme_internal_dek_kim_word[15]), .A2(iv1[15]), .A3(iv0[15]), .Z(n1044));
Q_MX04 U3185 ( .S0(n173), .S1(n172), .A0(guid3[15]), .A1(guid2[15]), .A2(guid1[15]), .A3(guid0[15]), .Z(n1045));
Q_MX02 U3186 ( .S(n172), .A0(n1047), .A1(stitcher_out[23]), .Z(n1046));
Q_AN02 U3187 ( .A0(n1153), .A1(stitcher_out[55]), .Z(n1047));
Q_MX03 U3188 ( .S0(n566), .S1(n557), .A0(n1053), .A1(n1052), .A2(n1048), .Z(fifo_in[14]));
Q_MX03 U3189 ( .S0(n172), .S1(n171), .A0(n1049), .A1(n1050), .A2(n1051), .Z(n1048));
Q_AN02 U3190 ( .A0(n173), .A1(stitcher_out[14]), .Z(n1049));
Q_AN02 U3191 ( .A0(n1153), .A1(kme_internal_word0[14]), .Z(n1050));
Q_MX04 U3192 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[14]), .A1(kme_internal_dek_kim_word[14]), .A2(iv1[14]), .A3(iv0[14]), .Z(n1051));
Q_MX04 U3193 ( .S0(n173), .S1(n172), .A0(guid3[14]), .A1(guid2[14]), .A2(guid1[14]), .A3(guid0[14]), .Z(n1052));
Q_MX02 U3194 ( .S(n172), .A0(n1054), .A1(stitcher_out[22]), .Z(n1053));
Q_AN02 U3195 ( .A0(n1153), .A1(stitcher_out[54]), .Z(n1054));
Q_MX03 U3196 ( .S0(n566), .S1(n557), .A0(n1060), .A1(n1059), .A2(n1055), .Z(fifo_in[13]));
Q_MX03 U3197 ( .S0(n172), .S1(n171), .A0(n1056), .A1(n1057), .A2(n1058), .Z(n1055));
Q_AN02 U3198 ( .A0(n173), .A1(stitcher_out[13]), .Z(n1056));
Q_AN02 U3199 ( .A0(n1153), .A1(kme_internal_word0[13]), .Z(n1057));
Q_MX04 U3200 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[13]), .A1(kme_internal_dek_kim_word[13]), .A2(iv1[13]), .A3(iv0[13]), .Z(n1058));
Q_MX04 U3201 ( .S0(n173), .S1(n172), .A0(guid3[13]), .A1(guid2[13]), .A2(guid1[13]), .A3(guid0[13]), .Z(n1059));
Q_MX02 U3202 ( .S(n172), .A0(n1061), .A1(stitcher_out[21]), .Z(n1060));
Q_AN02 U3203 ( .A0(n1153), .A1(stitcher_out[53]), .Z(n1061));
Q_MX03 U3204 ( .S0(n566), .S1(n557), .A0(n1067), .A1(n1066), .A2(n1062), .Z(fifo_in[12]));
Q_MX03 U3205 ( .S0(n172), .S1(n171), .A0(n1063), .A1(n1064), .A2(n1065), .Z(n1062));
Q_AN02 U3206 ( .A0(n173), .A1(stitcher_out[12]), .Z(n1063));
Q_AN02 U3207 ( .A0(n1153), .A1(kme_internal_word0[12]), .Z(n1064));
Q_MX04 U3208 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[12]), .A1(kme_internal_dek_kim_word[12]), .A2(iv1[12]), .A3(iv0[12]), .Z(n1065));
Q_MX04 U3209 ( .S0(n173), .S1(n172), .A0(guid3[12]), .A1(guid2[12]), .A2(guid1[12]), .A3(guid0[12]), .Z(n1066));
Q_MX02 U3210 ( .S(n172), .A0(n1068), .A1(stitcher_out[20]), .Z(n1067));
Q_AN02 U3211 ( .A0(n1153), .A1(stitcher_out[52]), .Z(n1068));
Q_MX03 U3212 ( .S0(n566), .S1(n557), .A0(n1074), .A1(n1073), .A2(n1069), .Z(fifo_in[11]));
Q_MX03 U3213 ( .S0(n172), .S1(n171), .A0(n1070), .A1(n1071), .A2(n1072), .Z(n1069));
Q_AN02 U3214 ( .A0(n173), .A1(stitcher_out[11]), .Z(n1070));
Q_AN02 U3215 ( .A0(n1153), .A1(kme_internal_word0[11]), .Z(n1071));
Q_MX04 U3216 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[11]), .A1(kme_internal_dek_kim_word[11]), .A2(iv1[11]), .A3(iv0[11]), .Z(n1072));
Q_MX04 U3217 ( .S0(n173), .S1(n172), .A0(guid3[11]), .A1(guid2[11]), .A2(guid1[11]), .A3(guid0[11]), .Z(n1073));
Q_MX02 U3218 ( .S(n172), .A0(n1075), .A1(stitcher_out[19]), .Z(n1074));
Q_AN02 U3219 ( .A0(n1153), .A1(stitcher_out[51]), .Z(n1075));
Q_MX03 U3220 ( .S0(n566), .S1(n557), .A0(n1081), .A1(n1080), .A2(n1076), .Z(fifo_in[10]));
Q_MX03 U3221 ( .S0(n172), .S1(n171), .A0(n1077), .A1(n1078), .A2(n1079), .Z(n1076));
Q_AN02 U3222 ( .A0(n173), .A1(stitcher_out[10]), .Z(n1077));
Q_AN02 U3223 ( .A0(n1153), .A1(kme_internal_word0[10]), .Z(n1078));
Q_MX04 U3224 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[10]), .A1(kme_internal_dek_kim_word[10]), .A2(iv1[10]), .A3(iv0[10]), .Z(n1079));
Q_MX04 U3225 ( .S0(n173), .S1(n172), .A0(guid3[10]), .A1(guid2[10]), .A2(guid1[10]), .A3(guid0[10]), .Z(n1080));
Q_MX02 U3226 ( .S(n172), .A0(n1082), .A1(stitcher_out[18]), .Z(n1081));
Q_AN02 U3227 ( .A0(n1153), .A1(stitcher_out[50]), .Z(n1082));
Q_MX03 U3228 ( .S0(n566), .S1(n557), .A0(n1088), .A1(n1087), .A2(n1083), .Z(fifo_in[9]));
Q_MX03 U3229 ( .S0(n172), .S1(n171), .A0(n1084), .A1(n1085), .A2(n1086), .Z(n1083));
Q_AN02 U3230 ( .A0(n173), .A1(stitcher_out[9]), .Z(n1084));
Q_AN02 U3231 ( .A0(n1153), .A1(kme_internal_word0[9]), .Z(n1085));
Q_MX04 U3232 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[9]), .A1(kme_internal_dek_kim_word[9]), .A2(iv1[9]), .A3(iv0[9]), .Z(n1086));
Q_MX04 U3233 ( .S0(n173), .S1(n172), .A0(guid3[9]), .A1(guid2[9]), .A2(guid1[9]), .A3(guid0[9]), .Z(n1087));
Q_MX02 U3234 ( .S(n172), .A0(n1089), .A1(stitcher_out[17]), .Z(n1088));
Q_AN02 U3235 ( .A0(n1153), .A1(stitcher_out[49]), .Z(n1089));
Q_MX03 U3236 ( .S0(n566), .S1(n557), .A0(n1095), .A1(n1094), .A2(n1090), .Z(fifo_in[8]));
Q_MX03 U3237 ( .S0(n172), .S1(n171), .A0(n1091), .A1(n1092), .A2(n1093), .Z(n1090));
Q_AN02 U3238 ( .A0(n173), .A1(stitcher_out[8]), .Z(n1091));
Q_AN02 U3239 ( .A0(n1153), .A1(kme_internal_word0[8]), .Z(n1092));
Q_MX04 U3240 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[8]), .A1(kme_internal_dek_kim_word[8]), .A2(iv1[8]), .A3(iv0[8]), .Z(n1093));
Q_MX04 U3241 ( .S0(n173), .S1(n172), .A0(guid3[8]), .A1(guid2[8]), .A2(guid1[8]), .A3(guid0[8]), .Z(n1094));
Q_MX02 U3242 ( .S(n172), .A0(n1096), .A1(stitcher_out[16]), .Z(n1095));
Q_AN02 U3243 ( .A0(n1153), .A1(stitcher_out[48]), .Z(n1096));
Q_MX03 U3244 ( .S0(n566), .S1(n557), .A0(n1102), .A1(n1101), .A2(n1097), .Z(fifo_in[7]));
Q_MX03 U3245 ( .S0(n172), .S1(n171), .A0(n1098), .A1(n1099), .A2(n1100), .Z(n1097));
Q_AN02 U3246 ( .A0(n173), .A1(stitcher_out[7]), .Z(n1098));
Q_AN02 U3247 ( .A0(n1153), .A1(kme_internal_word0[7]), .Z(n1099));
Q_MX04 U3248 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[7]), .A1(kme_internal_dek_kim_word[7]), .A2(iv1[7]), .A3(iv0[7]), .Z(n1100));
Q_MX04 U3249 ( .S0(n173), .S1(n172), .A0(guid3[7]), .A1(guid2[7]), .A2(guid1[7]), .A3(guid0[7]), .Z(n1101));
Q_MX02 U3250 ( .S(n172), .A0(n1103), .A1(stitcher_out[31]), .Z(n1102));
Q_AN02 U3251 ( .A0(n1153), .A1(stitcher_out[63]), .Z(n1103));
Q_MX03 U3252 ( .S0(n566), .S1(n557), .A0(n1109), .A1(n1108), .A2(n1104), .Z(fifo_in[6]));
Q_MX03 U3253 ( .S0(n172), .S1(n171), .A0(n1105), .A1(n1106), .A2(n1107), .Z(n1104));
Q_AN02 U3254 ( .A0(n173), .A1(stitcher_out[6]), .Z(n1105));
Q_AN02 U3255 ( .A0(n1153), .A1(kme_internal_word0[6]), .Z(n1106));
Q_MX04 U3256 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[6]), .A1(kme_internal_dek_kim_word[6]), .A2(iv1[6]), .A3(iv0[6]), .Z(n1107));
Q_MX04 U3257 ( .S0(n173), .S1(n172), .A0(guid3[6]), .A1(guid2[6]), .A2(guid1[6]), .A3(guid0[6]), .Z(n1108));
Q_MX02 U3258 ( .S(n172), .A0(n1110), .A1(stitcher_out[30]), .Z(n1109));
Q_AN02 U3259 ( .A0(n1153), .A1(stitcher_out[62]), .Z(n1110));
Q_MX03 U3260 ( .S0(n566), .S1(n557), .A0(n1116), .A1(n1115), .A2(n1111), .Z(fifo_in[5]));
Q_MX03 U3261 ( .S0(n172), .S1(n171), .A0(n1112), .A1(n1113), .A2(n1114), .Z(n1111));
Q_AN02 U3262 ( .A0(n173), .A1(stitcher_out[5]), .Z(n1112));
Q_AN02 U3263 ( .A0(n1153), .A1(kme_internal_word0[5]), .Z(n1113));
Q_MX04 U3264 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[5]), .A1(kme_internal_dek_kim_word[5]), .A2(iv1[5]), .A3(iv0[5]), .Z(n1114));
Q_MX04 U3265 ( .S0(n173), .S1(n172), .A0(guid3[5]), .A1(guid2[5]), .A2(guid1[5]), .A3(guid0[5]), .Z(n1115));
Q_MX02 U3266 ( .S(n172), .A0(n1117), .A1(stitcher_out[29]), .Z(n1116));
Q_AN02 U3267 ( .A0(n1153), .A1(stitcher_out[61]), .Z(n1117));
Q_MX03 U3268 ( .S0(n566), .S1(n557), .A0(n1123), .A1(n1122), .A2(n1118), .Z(fifo_in[4]));
Q_MX03 U3269 ( .S0(n172), .S1(n171), .A0(n1119), .A1(n1120), .A2(n1121), .Z(n1118));
Q_AN02 U3270 ( .A0(n173), .A1(stitcher_out[4]), .Z(n1119));
Q_AN02 U3271 ( .A0(n1153), .A1(kme_internal_word0[4]), .Z(n1120));
Q_MX04 U3272 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[4]), .A1(kme_internal_dek_kim_word[4]), .A2(iv1[4]), .A3(iv0[4]), .Z(n1121));
Q_MX04 U3273 ( .S0(n173), .S1(n172), .A0(guid3[4]), .A1(guid2[4]), .A2(guid1[4]), .A3(guid0[4]), .Z(n1122));
Q_MX02 U3274 ( .S(n172), .A0(n1124), .A1(stitcher_out[28]), .Z(n1123));
Q_AN02 U3275 ( .A0(n1153), .A1(stitcher_out[60]), .Z(n1124));
Q_MX03 U3276 ( .S0(n566), .S1(n557), .A0(n1130), .A1(n1129), .A2(n1125), .Z(fifo_in[3]));
Q_MX03 U3277 ( .S0(n172), .S1(n171), .A0(n1126), .A1(n1127), .A2(n1128), .Z(n1125));
Q_AN02 U3278 ( .A0(n173), .A1(stitcher_out[3]), .Z(n1126));
Q_AN02 U3279 ( .A0(n1153), .A1(kme_internal_word0[3]), .Z(n1127));
Q_MX04 U3280 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[3]), .A1(kme_internal_dek_kim_word[3]), .A2(iv1[3]), .A3(iv0[3]), .Z(n1128));
Q_MX04 U3281 ( .S0(n173), .S1(n172), .A0(guid3[3]), .A1(guid2[3]), .A2(guid1[3]), .A3(guid0[3]), .Z(n1129));
Q_MX02 U3282 ( .S(n172), .A0(n1131), .A1(stitcher_out[27]), .Z(n1130));
Q_AN02 U3283 ( .A0(n1153), .A1(stitcher_out[59]), .Z(n1131));
Q_MX03 U3284 ( .S0(n566), .S1(n557), .A0(n1137), .A1(n1136), .A2(n1132), .Z(fifo_in[2]));
Q_MX03 U3285 ( .S0(n172), .S1(n171), .A0(n1133), .A1(n1134), .A2(n1135), .Z(n1132));
Q_AN02 U3286 ( .A0(n173), .A1(stitcher_out[2]), .Z(n1133));
Q_AN02 U3287 ( .A0(n1153), .A1(kme_internal_word0[2]), .Z(n1134));
Q_MX04 U3288 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[2]), .A1(kme_internal_dek_kim_word[2]), .A2(iv1[2]), .A3(iv0[2]), .Z(n1135));
Q_MX04 U3289 ( .S0(n173), .S1(n172), .A0(guid3[2]), .A1(guid2[2]), .A2(guid1[2]), .A3(guid0[2]), .Z(n1136));
Q_MX02 U3290 ( .S(n172), .A0(n1138), .A1(stitcher_out[26]), .Z(n1137));
Q_AN02 U3291 ( .A0(n1153), .A1(stitcher_out[58]), .Z(n1138));
Q_MX03 U3292 ( .S0(n566), .S1(n557), .A0(n1144), .A1(n1143), .A2(n1139), .Z(fifo_in[1]));
Q_MX03 U3293 ( .S0(n172), .S1(n171), .A0(n1140), .A1(n1141), .A2(n1142), .Z(n1139));
Q_AN02 U3294 ( .A0(n173), .A1(stitcher_out[1]), .Z(n1140));
Q_AN02 U3295 ( .A0(n1153), .A1(kme_internal_word0[1]), .Z(n1141));
Q_MX04 U3296 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[1]), .A1(kme_internal_dek_kim_word[1]), .A2(iv1[1]), .A3(iv0[1]), .Z(n1142));
Q_MX04 U3297 ( .S0(n173), .S1(n172), .A0(guid3[1]), .A1(guid2[1]), .A2(guid1[1]), .A3(guid0[1]), .Z(n1143));
Q_MX02 U3298 ( .S(n172), .A0(n1145), .A1(stitcher_out[25]), .Z(n1144));
Q_AN02 U3299 ( .A0(n1153), .A1(stitcher_out[57]), .Z(n1145));
Q_MX03 U3300 ( .S0(n566), .S1(n557), .A0(n1151), .A1(n1150), .A2(n1146), .Z(fifo_in[0]));
Q_MX03 U3301 ( .S0(n172), .S1(n171), .A0(n1147), .A1(n1148), .A2(n1149), .Z(n1146));
Q_AN02 U3302 ( .A0(n173), .A1(stitcher_out[0]), .Z(n1147));
Q_AN02 U3303 ( .A0(n1153), .A1(kme_internal_word0[0]), .Z(n1148));
Q_MX04 U3304 ( .S0(n173), .S1(n172), .A0(kme_internal_dak_kim_word[0]), .A1(kme_internal_dek_kim_word[0]), .A2(iv1[0]), .A3(iv0[0]), .Z(n1149));
Q_MX04 U3305 ( .S0(n173), .S1(n172), .A0(guid3[0]), .A1(guid2[0]), .A2(guid1[0]), .A3(guid0[0]), .Z(n1150));
Q_MX02 U3306 ( .S(n172), .A0(n1152), .A1(stitcher_out[24]), .Z(n1151));
Q_AN02 U3307 ( .A0(n1153), .A1(stitcher_out[56]), .Z(n1152));
Q_INV U3308 ( .A(n173), .Z(n1153));
Q_AN02 U3309 ( .A0(n146), .A1(kme_internal_dek_kim_word[63]), .Z(nxt_kme_internal_dek_kim_word[63]));
Q_AN02 U3310 ( .A0(n146), .A1(kme_internal_dek_kim_word[62]), .Z(nxt_kme_internal_dek_kim_word[62]));
Q_AN02 U3311 ( .A0(n146), .A1(kme_internal_dek_kim_word[61]), .Z(nxt_kme_internal_dek_kim_word[61]));
Q_AN02 U3312 ( .A0(n146), .A1(kme_internal_dek_kim_word[60]), .Z(nxt_kme_internal_dek_kim_word[60]));
Q_AN02 U3313 ( .A0(n146), .A1(kme_internal_dek_kim_word[59]), .Z(nxt_kme_internal_dek_kim_word[59]));
Q_AN02 U3314 ( .A0(n146), .A1(kme_internal_dek_kim_word[58]), .Z(nxt_kme_internal_dek_kim_word[58]));
Q_AN02 U3315 ( .A0(n146), .A1(kme_internal_dek_kim_word[57]), .Z(nxt_kme_internal_dek_kim_word[57]));
Q_AN02 U3316 ( .A0(n146), .A1(kme_internal_dek_kim_word[56]), .Z(nxt_kme_internal_dek_kim_word[56]));
Q_AN02 U3317 ( .A0(n146), .A1(kme_internal_dek_kim_word[55]), .Z(nxt_kme_internal_dek_kim_word[55]));
Q_AN02 U3318 ( .A0(n146), .A1(kme_internal_dek_kim_word[54]), .Z(nxt_kme_internal_dek_kim_word[54]));
Q_AN02 U3319 ( .A0(n146), .A1(kme_internal_dek_kim_word[53]), .Z(nxt_kme_internal_dek_kim_word[53]));
Q_AN02 U3320 ( .A0(n146), .A1(kme_internal_dek_kim_word[52]), .Z(nxt_kme_internal_dek_kim_word[52]));
Q_AN02 U3321 ( .A0(n146), .A1(kme_internal_dek_kim_word[51]), .Z(nxt_kme_internal_dek_kim_word[51]));
Q_AN02 U3322 ( .A0(n146), .A1(kme_internal_dek_kim_word[50]), .Z(nxt_kme_internal_dek_kim_word[50]));
Q_AN02 U3323 ( .A0(n146), .A1(kme_internal_dek_kim_word[49]), .Z(nxt_kme_internal_dek_kim_word[49]));
Q_AN02 U3324 ( .A0(n146), .A1(kme_internal_dek_kim_word[48]), .Z(nxt_kme_internal_dek_kim_word[48]));
Q_AN02 U3325 ( .A0(n146), .A1(kme_internal_dek_kim_word[47]), .Z(nxt_kme_internal_dek_kim_word[47]));
Q_AN02 U3326 ( .A0(n146), .A1(kme_internal_dek_kim_word[46]), .Z(nxt_kme_internal_dek_kim_word[46]));
Q_AN02 U3327 ( .A0(n146), .A1(kme_internal_dek_kim_word[45]), .Z(nxt_kme_internal_dek_kim_word[45]));
Q_AN02 U3328 ( .A0(n146), .A1(kme_internal_dek_kim_word[44]), .Z(nxt_kme_internal_dek_kim_word[44]));
Q_AN02 U3329 ( .A0(n146), .A1(kme_internal_dek_kim_word[43]), .Z(nxt_kme_internal_dek_kim_word[43]));
Q_AN02 U3330 ( .A0(n146), .A1(kme_internal_dek_kim_word[42]), .Z(nxt_kme_internal_dek_kim_word[42]));
Q_AN02 U3331 ( .A0(n146), .A1(kme_internal_dek_kim_word[41]), .Z(nxt_kme_internal_dek_kim_word[41]));
Q_AN02 U3332 ( .A0(n146), .A1(kme_internal_dek_kim_word[40]), .Z(nxt_kme_internal_dek_kim_word[40]));
Q_AN02 U3333 ( .A0(n146), .A1(kme_internal_dek_kim_word[39]), .Z(nxt_kme_internal_dek_kim_word[39]));
Q_AN02 U3334 ( .A0(n146), .A1(kme_internal_dek_kim_word[38]), .Z(nxt_kme_internal_dek_kim_word[38]));
Q_AN02 U3335 ( .A0(n146), .A1(kme_internal_dek_kim_word[37]), .Z(nxt_kme_internal_dek_kim_word[37]));
Q_AN02 U3336 ( .A0(n146), .A1(kme_internal_dek_kim_word[36]), .Z(nxt_kme_internal_dek_kim_word[36]));
Q_AN02 U3337 ( .A0(n146), .A1(kme_internal_dek_kim_word[35]), .Z(nxt_kme_internal_dek_kim_word[35]));
Q_AN02 U3338 ( .A0(n146), .A1(kme_internal_dek_kim_word[34]), .Z(nxt_kme_internal_dek_kim_word[34]));
Q_AN02 U3339 ( .A0(n146), .A1(kme_internal_dek_kim_word[33]), .Z(nxt_kme_internal_dek_kim_word[33]));
Q_AN02 U3340 ( .A0(n146), .A1(kme_internal_dek_kim_word[32]), .Z(nxt_kme_internal_dek_kim_word[32]));
Q_AN02 U3341 ( .A0(n146), .A1(kme_internal_dek_kim_word[31]), .Z(nxt_kme_internal_dek_kim_word[31]));
Q_AN02 U3342 ( .A0(n146), .A1(kme_internal_dek_kim_word[30]), .Z(nxt_kme_internal_dek_kim_word[30]));
Q_AN02 U3343 ( .A0(n146), .A1(kme_internal_dek_kim_word[29]), .Z(nxt_kme_internal_dek_kim_word[29]));
Q_AN02 U3344 ( .A0(n146), .A1(kme_internal_dek_kim_word[28]), .Z(nxt_kme_internal_dek_kim_word[28]));
Q_AN02 U3345 ( .A0(n146), .A1(kme_internal_dek_kim_word[27]), .Z(nxt_kme_internal_dek_kim_word[27]));
Q_AN02 U3346 ( .A0(n146), .A1(kme_internal_dek_kim_word[26]), .Z(nxt_kme_internal_dek_kim_word[26]));
Q_AN02 U3347 ( .A0(n146), .A1(kme_internal_dek_kim_word[25]), .Z(nxt_kme_internal_dek_kim_word[25]));
Q_AN02 U3348 ( .A0(n146), .A1(kme_internal_dek_kim_word[24]), .Z(nxt_kme_internal_dek_kim_word[24]));
Q_AN02 U3349 ( .A0(n146), .A1(kme_internal_dek_kim_word[23]), .Z(nxt_kme_internal_dek_kim_word[23]));
Q_AN02 U3350 ( .A0(n146), .A1(kme_internal_dek_kim_word[22]), .Z(nxt_kme_internal_dek_kim_word[22]));
Q_AN02 U3351 ( .A0(n146), .A1(kme_internal_dek_kim_word[21]), .Z(nxt_kme_internal_dek_kim_word[21]));
Q_AN02 U3352 ( .A0(n146), .A1(kme_internal_dek_kim_word[20]), .Z(nxt_kme_internal_dek_kim_word[20]));
Q_MX02 U3353 ( .S(n192), .A0(n1154), .A1(n1710), .Z(nxt_kme_internal_dek_kim_word[19]));
Q_AN02 U3354 ( .A0(n147), .A1(kme_internal_dek_kim_word[19]), .Z(n1154));
Q_MX02 U3355 ( .S(n192), .A0(n1155), .A1(n1712), .Z(nxt_kme_internal_dek_kim_word[18]));
Q_AN02 U3356 ( .A0(n147), .A1(kme_internal_dek_kim_word[18]), .Z(n1155));
Q_MX02 U3357 ( .S(n146), .A0(stitcher_out[55]), .A1(kme_internal_dek_kim_word[16]), .Z(nxt_kme_internal_dek_kim_word[16]));
Q_MX02 U3358 ( .S(n149), .A0(n1156), .A1(kme_internal_dek_kim_word[15]), .Z(nxt_kme_internal_dek_kim_word[15]));
Q_MX02 U3359 ( .S(n149), .A0(n1157), .A1(kme_internal_dek_kim_word[14]), .Z(nxt_kme_internal_dek_kim_word[14]));
Q_MX02 U3360 ( .S(n149), .A0(n1158), .A1(kme_internal_dek_kim_word[13]), .Z(nxt_kme_internal_dek_kim_word[13]));
Q_MX02 U3361 ( .S(n149), .A0(n1159), .A1(kme_internal_dek_kim_word[12]), .Z(nxt_kme_internal_dek_kim_word[12]));
Q_MX02 U3362 ( .S(n149), .A0(n1160), .A1(kme_internal_dek_kim_word[11]), .Z(nxt_kme_internal_dek_kim_word[11]));
Q_MX02 U3363 ( .S(n149), .A0(n1161), .A1(kme_internal_dek_kim_word[10]), .Z(nxt_kme_internal_dek_kim_word[10]));
Q_MX02 U3364 ( .S(n149), .A0(n1162), .A1(kme_internal_dek_kim_word[9]), .Z(nxt_kme_internal_dek_kim_word[9]));
Q_MX02 U3365 ( .S(n149), .A0(n1163), .A1(kme_internal_dek_kim_word[8]), .Z(nxt_kme_internal_dek_kim_word[8]));
Q_MX02 U3366 ( .S(n149), .A0(n1164), .A1(kme_internal_dek_kim_word[7]), .Z(nxt_kme_internal_dek_kim_word[7]));
Q_MX02 U3367 ( .S(n149), .A0(n1165), .A1(kme_internal_dek_kim_word[6]), .Z(nxt_kme_internal_dek_kim_word[6]));
Q_MX02 U3368 ( .S(n149), .A0(n1166), .A1(kme_internal_dek_kim_word[5]), .Z(nxt_kme_internal_dek_kim_word[5]));
Q_MX02 U3369 ( .S(n149), .A0(n1167), .A1(kme_internal_dek_kim_word[4]), .Z(nxt_kme_internal_dek_kim_word[4]));
Q_MX02 U3370 ( .S(n149), .A0(n1168), .A1(kme_internal_dek_kim_word[3]), .Z(nxt_kme_internal_dek_kim_word[3]));
Q_MX02 U3371 ( .S(n149), .A0(n1169), .A1(kme_internal_dek_kim_word[2]), .Z(nxt_kme_internal_dek_kim_word[2]));
Q_MX02 U3372 ( .S(n149), .A0(n1170), .A1(kme_internal_dek_kim_word[1]), .Z(nxt_kme_internal_dek_kim_word[1]));
Q_MX02 U3373 ( .S(n149), .A0(n1171), .A1(kme_internal_dek_kim_word[0]), .Z(nxt_kme_internal_dek_kim_word[0]));
Q_AN02 U3374 ( .A0(n146), .A1(kme_internal_dak_kim_word[63]), .Z(nxt_kme_internal_dak_kim_word[63]));
Q_AN02 U3375 ( .A0(n146), .A1(kme_internal_dak_kim_word[62]), .Z(nxt_kme_internal_dak_kim_word[62]));
Q_AN02 U3376 ( .A0(n146), .A1(kme_internal_dak_kim_word[61]), .Z(nxt_kme_internal_dak_kim_word[61]));
Q_AN02 U3377 ( .A0(n146), .A1(kme_internal_dak_kim_word[60]), .Z(nxt_kme_internal_dak_kim_word[60]));
Q_AN02 U3378 ( .A0(n146), .A1(kme_internal_dak_kim_word[59]), .Z(nxt_kme_internal_dak_kim_word[59]));
Q_AN02 U3379 ( .A0(n146), .A1(kme_internal_dak_kim_word[58]), .Z(nxt_kme_internal_dak_kim_word[58]));
Q_AN02 U3380 ( .A0(n146), .A1(kme_internal_dak_kim_word[57]), .Z(nxt_kme_internal_dak_kim_word[57]));
Q_AN02 U3381 ( .A0(n146), .A1(kme_internal_dak_kim_word[56]), .Z(nxt_kme_internal_dak_kim_word[56]));
Q_AN02 U3382 ( .A0(n146), .A1(kme_internal_dak_kim_word[55]), .Z(nxt_kme_internal_dak_kim_word[55]));
Q_AN02 U3383 ( .A0(n146), .A1(kme_internal_dak_kim_word[54]), .Z(nxt_kme_internal_dak_kim_word[54]));
Q_AN02 U3384 ( .A0(n146), .A1(kme_internal_dak_kim_word[53]), .Z(nxt_kme_internal_dak_kim_word[53]));
Q_AN02 U3385 ( .A0(n146), .A1(kme_internal_dak_kim_word[52]), .Z(nxt_kme_internal_dak_kim_word[52]));
Q_AN02 U3386 ( .A0(n146), .A1(kme_internal_dak_kim_word[51]), .Z(nxt_kme_internal_dak_kim_word[51]));
Q_AN02 U3387 ( .A0(n146), .A1(kme_internal_dak_kim_word[50]), .Z(nxt_kme_internal_dak_kim_word[50]));
Q_AN02 U3388 ( .A0(n146), .A1(kme_internal_dak_kim_word[49]), .Z(nxt_kme_internal_dak_kim_word[49]));
Q_AN02 U3389 ( .A0(n146), .A1(kme_internal_dak_kim_word[48]), .Z(nxt_kme_internal_dak_kim_word[48]));
Q_AN02 U3390 ( .A0(n146), .A1(kme_internal_dak_kim_word[47]), .Z(nxt_kme_internal_dak_kim_word[47]));
Q_AN02 U3391 ( .A0(n146), .A1(kme_internal_dak_kim_word[46]), .Z(nxt_kme_internal_dak_kim_word[46]));
Q_AN02 U3392 ( .A0(n146), .A1(kme_internal_dak_kim_word[45]), .Z(nxt_kme_internal_dak_kim_word[45]));
Q_AN02 U3393 ( .A0(n146), .A1(kme_internal_dak_kim_word[44]), .Z(nxt_kme_internal_dak_kim_word[44]));
Q_AN02 U3394 ( .A0(n146), .A1(kme_internal_dak_kim_word[43]), .Z(nxt_kme_internal_dak_kim_word[43]));
Q_AN02 U3395 ( .A0(n146), .A1(kme_internal_dak_kim_word[42]), .Z(nxt_kme_internal_dak_kim_word[42]));
Q_AN02 U3396 ( .A0(n146), .A1(kme_internal_dak_kim_word[41]), .Z(nxt_kme_internal_dak_kim_word[41]));
Q_AN02 U3397 ( .A0(n146), .A1(kme_internal_dak_kim_word[40]), .Z(nxt_kme_internal_dak_kim_word[40]));
Q_AN02 U3398 ( .A0(n146), .A1(kme_internal_dak_kim_word[39]), .Z(nxt_kme_internal_dak_kim_word[39]));
Q_AN02 U3399 ( .A0(n146), .A1(kme_internal_dak_kim_word[38]), .Z(nxt_kme_internal_dak_kim_word[38]));
Q_AN02 U3400 ( .A0(n146), .A1(kme_internal_dak_kim_word[37]), .Z(nxt_kme_internal_dak_kim_word[37]));
Q_AN02 U3401 ( .A0(n146), .A1(kme_internal_dak_kim_word[36]), .Z(nxt_kme_internal_dak_kim_word[36]));
Q_AN02 U3402 ( .A0(n146), .A1(kme_internal_dak_kim_word[35]), .Z(nxt_kme_internal_dak_kim_word[35]));
Q_AN02 U3403 ( .A0(n146), .A1(kme_internal_dak_kim_word[34]), .Z(nxt_kme_internal_dak_kim_word[34]));
Q_AN02 U3404 ( .A0(n146), .A1(kme_internal_dak_kim_word[33]), .Z(nxt_kme_internal_dak_kim_word[33]));
Q_AN02 U3405 ( .A0(n146), .A1(kme_internal_dak_kim_word[32]), .Z(nxt_kme_internal_dak_kim_word[32]));
Q_AN02 U3406 ( .A0(n146), .A1(kme_internal_dak_kim_word[31]), .Z(nxt_kme_internal_dak_kim_word[31]));
Q_AN02 U3407 ( .A0(n146), .A1(kme_internal_dak_kim_word[30]), .Z(nxt_kme_internal_dak_kim_word[30]));
Q_AN02 U3408 ( .A0(n146), .A1(kme_internal_dak_kim_word[29]), .Z(nxt_kme_internal_dak_kim_word[29]));
Q_AN02 U3409 ( .A0(n146), .A1(kme_internal_dak_kim_word[28]), .Z(nxt_kme_internal_dak_kim_word[28]));
Q_AN02 U3410 ( .A0(n146), .A1(kme_internal_dak_kim_word[27]), .Z(nxt_kme_internal_dak_kim_word[27]));
Q_AN02 U3411 ( .A0(n146), .A1(kme_internal_dak_kim_word[26]), .Z(nxt_kme_internal_dak_kim_word[26]));
Q_AN02 U3412 ( .A0(n146), .A1(kme_internal_dak_kim_word[25]), .Z(nxt_kme_internal_dak_kim_word[25]));
Q_AN02 U3413 ( .A0(n146), .A1(kme_internal_dak_kim_word[24]), .Z(nxt_kme_internal_dak_kim_word[24]));
Q_AN02 U3414 ( .A0(n146), .A1(kme_internal_dak_kim_word[23]), .Z(nxt_kme_internal_dak_kim_word[23]));
Q_AN02 U3415 ( .A0(n146), .A1(kme_internal_dak_kim_word[22]), .Z(nxt_kme_internal_dak_kim_word[22]));
Q_AN02 U3416 ( .A0(n146), .A1(kme_internal_dak_kim_word[21]), .Z(nxt_kme_internal_dak_kim_word[21]));
Q_AN02 U3417 ( .A0(n146), .A1(kme_internal_dak_kim_word[20]), .Z(nxt_kme_internal_dak_kim_word[20]));
Q_AN02 U3418 ( .A0(n146), .A1(kme_internal_dak_kim_word[19]), .Z(nxt_kme_internal_dak_kim_word[19]));
Q_AN02 U3419 ( .A0(n146), .A1(kme_internal_dak_kim_word[18]), .Z(nxt_kme_internal_dak_kim_word[18]));
Q_MX02 U3420 ( .S(n146), .A0(stitcher_out[55]), .A1(kme_internal_dak_kim_word[16]), .Z(nxt_kme_internal_dak_kim_word[16]));
Q_MX02 U3421 ( .S(n149), .A0(n1156), .A1(kme_internal_dak_kim_word[15]), .Z(nxt_kme_internal_dak_kim_word[15]));
Q_AN02 U3422 ( .A0(n198), .A1(stitcher_out[63]), .Z(n1156));
Q_MX02 U3423 ( .S(n149), .A0(n1157), .A1(kme_internal_dak_kim_word[14]), .Z(nxt_kme_internal_dak_kim_word[14]));
Q_AN02 U3424 ( .A0(n198), .A1(stitcher_out[62]), .Z(n1157));
Q_MX02 U3425 ( .S(n149), .A0(n1158), .A1(kme_internal_dak_kim_word[13]), .Z(nxt_kme_internal_dak_kim_word[13]));
Q_AN02 U3426 ( .A0(n198), .A1(stitcher_out[61]), .Z(n1158));
Q_MX02 U3427 ( .S(n149), .A0(n1159), .A1(kme_internal_dak_kim_word[12]), .Z(nxt_kme_internal_dak_kim_word[12]));
Q_AN02 U3428 ( .A0(n198), .A1(stitcher_out[60]), .Z(n1159));
Q_MX02 U3429 ( .S(n149), .A0(n1160), .A1(kme_internal_dak_kim_word[11]), .Z(nxt_kme_internal_dak_kim_word[11]));
Q_AN02 U3430 ( .A0(n198), .A1(stitcher_out[59]), .Z(n1160));
Q_MX02 U3431 ( .S(n149), .A0(n1161), .A1(kme_internal_dak_kim_word[10]), .Z(nxt_kme_internal_dak_kim_word[10]));
Q_AN02 U3432 ( .A0(n198), .A1(stitcher_out[58]), .Z(n1161));
Q_MX02 U3433 ( .S(n149), .A0(n1162), .A1(kme_internal_dak_kim_word[9]), .Z(nxt_kme_internal_dak_kim_word[9]));
Q_AN02 U3434 ( .A0(n198), .A1(stitcher_out[57]), .Z(n1162));
Q_MX02 U3435 ( .S(n149), .A0(n1163), .A1(kme_internal_dak_kim_word[8]), .Z(nxt_kme_internal_dak_kim_word[8]));
Q_AN02 U3436 ( .A0(n198), .A1(stitcher_out[56]), .Z(n1163));
Q_MX02 U3437 ( .S(n149), .A0(n1164), .A1(kme_internal_dak_kim_word[7]), .Z(nxt_kme_internal_dak_kim_word[7]));
Q_AN02 U3438 ( .A0(n198), .A1(stitcher_out[55]), .Z(n1164));
Q_MX02 U3439 ( .S(n149), .A0(n1165), .A1(kme_internal_dak_kim_word[6]), .Z(nxt_kme_internal_dak_kim_word[6]));
Q_AN02 U3440 ( .A0(n198), .A1(stitcher_out[54]), .Z(n1165));
Q_MX02 U3441 ( .S(n149), .A0(n1166), .A1(kme_internal_dak_kim_word[5]), .Z(nxt_kme_internal_dak_kim_word[5]));
Q_AN02 U3442 ( .A0(n198), .A1(stitcher_out[53]), .Z(n1166));
Q_MX02 U3443 ( .S(n149), .A0(n1167), .A1(kme_internal_dak_kim_word[4]), .Z(nxt_kme_internal_dak_kim_word[4]));
Q_AN02 U3444 ( .A0(n198), .A1(stitcher_out[52]), .Z(n1167));
Q_MX02 U3445 ( .S(n149), .A0(n1168), .A1(kme_internal_dak_kim_word[3]), .Z(nxt_kme_internal_dak_kim_word[3]));
Q_AN02 U3446 ( .A0(n198), .A1(stitcher_out[51]), .Z(n1168));
Q_MX02 U3447 ( .S(n149), .A0(n1169), .A1(kme_internal_dak_kim_word[2]), .Z(nxt_kme_internal_dak_kim_word[2]));
Q_AN02 U3448 ( .A0(n198), .A1(stitcher_out[50]), .Z(n1169));
Q_MX02 U3449 ( .S(n149), .A0(n1170), .A1(kme_internal_dak_kim_word[1]), .Z(nxt_kme_internal_dak_kim_word[1]));
Q_AN02 U3450 ( .A0(n198), .A1(stitcher_out[49]), .Z(n1170));
Q_MX02 U3451 ( .S(n149), .A0(n1171), .A1(kme_internal_dak_kim_word[0]), .Z(nxt_kme_internal_dak_kim_word[0]));
Q_AN02 U3452 ( .A0(n198), .A1(stitcher_out[48]), .Z(n1171));
Q_AN02 U3453 ( .A0(n150), .A1(n1172), .Z(nxt_tlv_type[7]));
Q_MX02 U3454 ( .S(n205), .A0(stitcher_out[7]), .A1(tlv_type[7]), .Z(n1172));
Q_AN02 U3455 ( .A0(n150), .A1(n1173), .Z(nxt_tlv_type[6]));
Q_MX02 U3456 ( .S(n205), .A0(stitcher_out[6]), .A1(tlv_type[6]), .Z(n1173));
Q_AN02 U3457 ( .A0(n150), .A1(n1174), .Z(nxt_tlv_type[5]));
Q_MX02 U3458 ( .S(n205), .A0(stitcher_out[5]), .A1(tlv_type[5]), .Z(n1174));
Q_OR02 U3459 ( .A0(n1176), .A1(n1175), .Z(nxt_tlv_type[4]));
Q_MX02 U3460 ( .S(n205), .A0(stitcher_out[4]), .A1(tlv_type[4]), .Z(n1175));
Q_OR02 U3461 ( .A0(n1176), .A1(n1177), .Z(nxt_tlv_type[3]));
Q_INV U3462 ( .A(n150), .Z(n1176));
Q_MX02 U3463 ( .S(n205), .A0(stitcher_out[3]), .A1(tlv_type[3]), .Z(n1177));
Q_AN02 U3464 ( .A0(n150), .A1(n1178), .Z(nxt_tlv_type[2]));
Q_MX02 U3465 ( .S(n205), .A0(stitcher_out[2]), .A1(tlv_type[2]), .Z(n1178));
Q_AN02 U3466 ( .A0(n150), .A1(n1179), .Z(nxt_tlv_type[1]));
Q_MX02 U3467 ( .S(n205), .A0(stitcher_out[1]), .A1(tlv_type[1]), .Z(n1179));
Q_MX02 U3468 ( .S(n150), .A0(n205), .A1(n1180), .Z(nxt_tlv_type[0]));
Q_MX02 U3469 ( .S(n205), .A0(stitcher_out[0]), .A1(tlv_type[0]), .Z(n1180));
Q_MX02 U3470 ( .S(n631), .A0(stitcher_out[62]), .A1(n1181), .Z(nxt_aux_key_type[5]));
Q_AN02 U3471 ( .A0(n169), .A1(aux_key_type[5]), .Z(n1181));
Q_MX02 U3472 ( .S(n631), .A0(stitcher_out[61]), .A1(n1182), .Z(nxt_aux_key_type[4]));
Q_AN02 U3473 ( .A0(n169), .A1(aux_key_type[4]), .Z(n1182));
Q_MX02 U3474 ( .S(n631), .A0(stitcher_out[60]), .A1(n1183), .Z(nxt_aux_key_type[3]));
Q_AN02 U3475 ( .A0(n169), .A1(aux_key_type[3]), .Z(n1183));
Q_MX02 U3476 ( .S(n631), .A0(stitcher_out[59]), .A1(n1184), .Z(nxt_aux_key_type[2]));
Q_AN02 U3477 ( .A0(n169), .A1(aux_key_type[2]), .Z(n1184));
Q_MX02 U3478 ( .S(n631), .A0(stitcher_out[58]), .A1(n1185), .Z(nxt_aux_key_type[1]));
Q_AN02 U3479 ( .A0(n169), .A1(aux_key_type[1]), .Z(n1185));
Q_MX02 U3480 ( .S(n631), .A0(stitcher_out[57]), .A1(n1186), .Z(nxt_aux_key_type[0]));
Q_AN02 U3481 ( .A0(n169), .A1(aux_key_type[0]), .Z(n1186));
Q_MX02 U3482 ( .S(n631), .A0(stitcher_out[53]), .A1(n1187), .Z(nxt_aux_iv_op[1]));
Q_AN02 U3483 ( .A0(n169), .A1(aux_iv_op[1]), .Z(n1187));
Q_MX02 U3484 ( .S(n631), .A0(stitcher_out[52]), .A1(n1188), .Z(nxt_aux_iv_op[0]));
Q_AN02 U3485 ( .A0(n169), .A1(aux_iv_op[0]), .Z(n1188));
Q_MX02 U3486 ( .S(n631), .A0(stitcher_out[43]), .A1(n1189), .Z(nxt_aux_cipher_op[3]));
Q_AN02 U3487 ( .A0(n169), .A1(aux_cipher_op[3]), .Z(n1189));
Q_MX02 U3488 ( .S(n631), .A0(stitcher_out[42]), .A1(n1190), .Z(nxt_aux_cipher_op[2]));
Q_AN02 U3489 ( .A0(n169), .A1(aux_cipher_op[2]), .Z(n1190));
Q_MX02 U3490 ( .S(n631), .A0(stitcher_out[41]), .A1(n1191), .Z(nxt_aux_cipher_op[1]));
Q_AN02 U3491 ( .A0(n169), .A1(aux_cipher_op[1]), .Z(n1191));
Q_MX02 U3492 ( .S(n631), .A0(stitcher_out[40]), .A1(n1192), .Z(nxt_aux_cipher_op[0]));
Q_AN02 U3493 ( .A0(n169), .A1(aux_cipher_op[0]), .Z(n1192));
Q_MX02 U3494 ( .S(n631), .A0(stitcher_out[39]), .A1(n1193), .Z(nxt_aux_auth_op[3]));
Q_AN02 U3495 ( .A0(n169), .A1(aux_auth_op[3]), .Z(n1193));
Q_MX02 U3496 ( .S(n631), .A0(stitcher_out[38]), .A1(n1194), .Z(nxt_aux_auth_op[2]));
Q_AN02 U3497 ( .A0(n169), .A1(aux_auth_op[2]), .Z(n1194));
Q_MX02 U3498 ( .S(n631), .A0(stitcher_out[37]), .A1(n1195), .Z(nxt_aux_auth_op[1]));
Q_AN02 U3499 ( .A0(n169), .A1(aux_auth_op[1]), .Z(n1195));
Q_MX02 U3500 ( .S(n631), .A0(stitcher_out[36]), .A1(n1196), .Z(nxt_aux_auth_op[0]));
Q_AN02 U3501 ( .A0(n169), .A1(aux_auth_op[0]), .Z(n1196));
Q_MX02 U3502 ( .S(n631), .A0(stitcher_out[35]), .A1(n1197), .Z(nxt_aux_raw_auth_op[3]));
Q_AN02 U3503 ( .A0(n169), .A1(aux_raw_auth_op[3]), .Z(n1197));
Q_MX02 U3504 ( .S(n631), .A0(stitcher_out[34]), .A1(n1198), .Z(nxt_aux_raw_auth_op[2]));
Q_AN02 U3505 ( .A0(n169), .A1(aux_raw_auth_op[2]), .Z(n1198));
Q_MX02 U3506 ( .S(n631), .A0(stitcher_out[33]), .A1(n1199), .Z(nxt_aux_raw_auth_op[1]));
Q_AN02 U3507 ( .A0(n169), .A1(aux_raw_auth_op[1]), .Z(n1199));
Q_MX02 U3508 ( .S(n631), .A0(stitcher_out[32]), .A1(n1200), .Z(nxt_aux_raw_auth_op[0]));
Q_AN02 U3509 ( .A0(n169), .A1(aux_raw_auth_op[0]), .Z(n1200));
Q_MX02 U3510 ( .S(n207), .A0(n1201), .A1(stitcher_out[63]), .Z(nxt_debug_cmd[31]));
Q_AN02 U3511 ( .A0(n151), .A1(debug_cmd[31]), .Z(n1201));
Q_MX02 U3512 ( .S(n207), .A0(n1202), .A1(stitcher_out[62]), .Z(nxt_debug_cmd[30]));
Q_AN02 U3513 ( .A0(n151), .A1(debug_cmd[30]), .Z(n1202));
Q_MX02 U3514 ( .S(n207), .A0(n1203), .A1(stitcher_out[61]), .Z(nxt_debug_cmd[29]));
Q_AN02 U3515 ( .A0(n151), .A1(debug_cmd[29]), .Z(n1203));
Q_MX02 U3516 ( .S(n207), .A0(n1204), .A1(stitcher_out[60]), .Z(nxt_debug_cmd[28]));
Q_AN02 U3517 ( .A0(n151), .A1(debug_cmd[28]), .Z(n1204));
Q_MX02 U3518 ( .S(n207), .A0(n1205), .A1(stitcher_out[59]), .Z(nxt_debug_cmd[27]));
Q_AN02 U3519 ( .A0(n151), .A1(debug_cmd[27]), .Z(n1205));
Q_MX02 U3520 ( .S(n207), .A0(n1206), .A1(stitcher_out[58]), .Z(nxt_debug_cmd[26]));
Q_AN02 U3521 ( .A0(n151), .A1(debug_cmd[26]), .Z(n1206));
Q_MX02 U3522 ( .S(n207), .A0(n1207), .A1(stitcher_out[57]), .Z(nxt_debug_cmd[25]));
Q_AN02 U3523 ( .A0(n151), .A1(debug_cmd[25]), .Z(n1207));
Q_MX02 U3524 ( .S(n207), .A0(n1208), .A1(stitcher_out[56]), .Z(nxt_debug_cmd[24]));
Q_AN02 U3525 ( .A0(n151), .A1(debug_cmd[24]), .Z(n1208));
Q_MX02 U3526 ( .S(n207), .A0(n1209), .A1(stitcher_out[55]), .Z(nxt_debug_cmd[23]));
Q_AN02 U3527 ( .A0(n151), .A1(debug_cmd[23]), .Z(n1209));
Q_MX02 U3528 ( .S(n207), .A0(n1210), .A1(stitcher_out[54]), .Z(nxt_debug_cmd[22]));
Q_AN02 U3529 ( .A0(n151), .A1(debug_cmd[22]), .Z(n1210));
Q_MX02 U3530 ( .S(n207), .A0(n1211), .A1(stitcher_out[53]), .Z(nxt_debug_cmd[21]));
Q_AN02 U3531 ( .A0(n151), .A1(debug_cmd[21]), .Z(n1211));
Q_MX02 U3532 ( .S(n207), .A0(n1212), .A1(stitcher_out[52]), .Z(nxt_debug_cmd[20]));
Q_AN02 U3533 ( .A0(n151), .A1(debug_cmd[20]), .Z(n1212));
Q_MX02 U3534 ( .S(n207), .A0(n1213), .A1(stitcher_out[51]), .Z(nxt_debug_cmd[19]));
Q_AN02 U3535 ( .A0(n151), .A1(debug_cmd[19]), .Z(n1213));
Q_MX02 U3536 ( .S(n207), .A0(n1214), .A1(stitcher_out[50]), .Z(nxt_debug_cmd[18]));
Q_AN02 U3537 ( .A0(n151), .A1(debug_cmd[18]), .Z(n1214));
Q_MX02 U3538 ( .S(n207), .A0(n1215), .A1(stitcher_out[49]), .Z(nxt_debug_cmd[17]));
Q_AN02 U3539 ( .A0(n151), .A1(debug_cmd[17]), .Z(n1215));
Q_MX02 U3540 ( .S(n207), .A0(n1216), .A1(stitcher_out[48]), .Z(nxt_debug_cmd[16]));
Q_AN02 U3541 ( .A0(n151), .A1(debug_cmd[16]), .Z(n1216));
Q_MX02 U3542 ( .S(n207), .A0(n1217), .A1(stitcher_out[47]), .Z(nxt_debug_cmd[15]));
Q_AN02 U3543 ( .A0(n151), .A1(debug_cmd[15]), .Z(n1217));
Q_MX02 U3544 ( .S(n207), .A0(n1218), .A1(stitcher_out[46]), .Z(nxt_debug_cmd[14]));
Q_AN02 U3545 ( .A0(n151), .A1(debug_cmd[14]), .Z(n1218));
Q_MX02 U3546 ( .S(n207), .A0(n1219), .A1(stitcher_out[45]), .Z(nxt_debug_cmd[13]));
Q_AN02 U3547 ( .A0(n151), .A1(debug_cmd[13]), .Z(n1219));
Q_MX02 U3548 ( .S(n207), .A0(n1220), .A1(stitcher_out[44]), .Z(nxt_debug_cmd[12]));
Q_AN02 U3549 ( .A0(n151), .A1(debug_cmd[12]), .Z(n1220));
Q_MX02 U3550 ( .S(n207), .A0(n1221), .A1(stitcher_out[43]), .Z(nxt_debug_cmd[11]));
Q_AN02 U3551 ( .A0(n151), .A1(debug_cmd[11]), .Z(n1221));
Q_MX02 U3552 ( .S(n207), .A0(n1222), .A1(stitcher_out[42]), .Z(nxt_debug_cmd[10]));
Q_AN02 U3553 ( .A0(n151), .A1(debug_cmd[10]), .Z(n1222));
Q_MX02 U3554 ( .S(n207), .A0(n1223), .A1(stitcher_out[41]), .Z(nxt_debug_cmd[9]));
Q_AN02 U3555 ( .A0(n151), .A1(debug_cmd[9]), .Z(n1223));
Q_MX02 U3556 ( .S(n207), .A0(n1224), .A1(stitcher_out[40]), .Z(nxt_debug_cmd[8]));
Q_AN02 U3557 ( .A0(n151), .A1(debug_cmd[8]), .Z(n1224));
Q_MX02 U3558 ( .S(n207), .A0(n1225), .A1(stitcher_out[39]), .Z(nxt_debug_cmd[7]));
Q_AN02 U3559 ( .A0(n151), .A1(debug_cmd[7]), .Z(n1225));
Q_MX02 U3560 ( .S(n207), .A0(n1226), .A1(stitcher_out[38]), .Z(nxt_debug_cmd[6]));
Q_AN02 U3561 ( .A0(n151), .A1(debug_cmd[6]), .Z(n1226));
Q_MX02 U3562 ( .S(n207), .A0(n1227), .A1(stitcher_out[37]), .Z(nxt_debug_cmd[5]));
Q_AN02 U3563 ( .A0(n151), .A1(debug_cmd[5]), .Z(n1227));
Q_MX02 U3564 ( .S(n207), .A0(n1228), .A1(stitcher_out[36]), .Z(nxt_debug_cmd[4]));
Q_AN02 U3565 ( .A0(n151), .A1(debug_cmd[4]), .Z(n1228));
Q_MX02 U3566 ( .S(n207), .A0(n1229), .A1(stitcher_out[35]), .Z(nxt_debug_cmd[3]));
Q_AN02 U3567 ( .A0(n151), .A1(debug_cmd[3]), .Z(n1229));
Q_MX02 U3568 ( .S(n207), .A0(n1230), .A1(stitcher_out[34]), .Z(nxt_debug_cmd[2]));
Q_AN02 U3569 ( .A0(n151), .A1(debug_cmd[2]), .Z(n1230));
Q_MX02 U3570 ( .S(n207), .A0(n1231), .A1(stitcher_out[33]), .Z(nxt_debug_cmd[1]));
Q_AN02 U3571 ( .A0(n151), .A1(debug_cmd[1]), .Z(n1231));
Q_MX02 U3572 ( .S(n207), .A0(n1232), .A1(stitcher_out[32]), .Z(nxt_debug_cmd[0]));
Q_AN02 U3573 ( .A0(n151), .A1(debug_cmd[0]), .Z(n1232));
Q_MX02 U3574 ( .S(n268), .A0(skip[6]), .A1(n152), .Z(nxt_skip[6]));
Q_MX02 U3575 ( .S(n299), .A0(skip[5]), .A1(n153), .Z(nxt_skip[5]));
Q_MX02 U3576 ( .S(n308), .A0(skip[4]), .A1(n154), .Z(nxt_skip[4]));
Q_AO21 U3577 ( .A0(n1234), .A1(skip[0]), .B0(n1239), .Z(nxt_skip[0]));
Q_AN02 U3578 ( .A0(n1234), .A1(skip[1]), .Z(n1233));
Q_AO21 U3579 ( .A0(n1234), .A1(skip[2]), .B0(n1237), .Z(nxt_skip[2]));
Q_AO21 U3580 ( .A0(n1234), .A1(skip[3]), .B0(n1235), .Z(nxt_skip[3]));
Q_AN02 U3581 ( .A0(n156), .A1(n155), .Z(n1234));
Q_MX02 U3582 ( .S(n387), .A0(n155), .A1(n1234), .Z(n1236));
Q_INV U3583 ( .A(n1236), .Z(n1235));
Q_NR02 U3584 ( .A0(n157), .A1(n156), .Z(n1237));
Q_AO21 U3585 ( .A0(n157), .A1(n156), .B0(n1233), .Z(nxt_skip[1]));
Q_XNR2 U3586 ( .A0(n156), .A1(n155), .Z(n1238));
Q_NR02 U3587 ( .A0(n157), .A1(n1238), .Z(n1239));
Q_MX02 U3588 ( .S(n388), .A0(n1240), .A1(stitcher_out[7]), .Z(nxt_guid0[63]));
Q_AN02 U3589 ( .A0(n158), .A1(guid0[63]), .Z(n1240));
Q_MX02 U3590 ( .S(n388), .A0(n1241), .A1(stitcher_out[6]), .Z(nxt_guid0[62]));
Q_AN02 U3591 ( .A0(n158), .A1(guid0[62]), .Z(n1241));
Q_MX02 U3592 ( .S(n388), .A0(n1242), .A1(stitcher_out[5]), .Z(nxt_guid0[61]));
Q_AN02 U3593 ( .A0(n158), .A1(guid0[61]), .Z(n1242));
Q_MX02 U3594 ( .S(n388), .A0(n1243), .A1(stitcher_out[4]), .Z(nxt_guid0[60]));
Q_AN02 U3595 ( .A0(n158), .A1(guid0[60]), .Z(n1243));
Q_MX02 U3596 ( .S(n388), .A0(n1244), .A1(stitcher_out[3]), .Z(nxt_guid0[59]));
Q_AN02 U3597 ( .A0(n158), .A1(guid0[59]), .Z(n1244));
Q_MX02 U3598 ( .S(n388), .A0(n1245), .A1(stitcher_out[2]), .Z(nxt_guid0[58]));
Q_AN02 U3599 ( .A0(n158), .A1(guid0[58]), .Z(n1245));
Q_MX02 U3600 ( .S(n388), .A0(n1246), .A1(stitcher_out[1]), .Z(nxt_guid0[57]));
Q_AN02 U3601 ( .A0(n158), .A1(guid0[57]), .Z(n1246));
Q_MX02 U3602 ( .S(n388), .A0(n1247), .A1(stitcher_out[0]), .Z(nxt_guid0[56]));
Q_AN02 U3603 ( .A0(n158), .A1(guid0[56]), .Z(n1247));
Q_MX02 U3604 ( .S(n388), .A0(n1248), .A1(stitcher_out[15]), .Z(nxt_guid0[55]));
Q_AN02 U3605 ( .A0(n158), .A1(guid0[55]), .Z(n1248));
Q_MX02 U3606 ( .S(n388), .A0(n1249), .A1(stitcher_out[14]), .Z(nxt_guid0[54]));
Q_AN02 U3607 ( .A0(n158), .A1(guid0[54]), .Z(n1249));
Q_MX02 U3608 ( .S(n388), .A0(n1250), .A1(stitcher_out[13]), .Z(nxt_guid0[53]));
Q_AN02 U3609 ( .A0(n158), .A1(guid0[53]), .Z(n1250));
Q_MX02 U3610 ( .S(n388), .A0(n1251), .A1(stitcher_out[12]), .Z(nxt_guid0[52]));
Q_AN02 U3611 ( .A0(n158), .A1(guid0[52]), .Z(n1251));
Q_MX02 U3612 ( .S(n388), .A0(n1252), .A1(stitcher_out[11]), .Z(nxt_guid0[51]));
Q_AN02 U3613 ( .A0(n158), .A1(guid0[51]), .Z(n1252));
Q_MX02 U3614 ( .S(n388), .A0(n1253), .A1(stitcher_out[10]), .Z(nxt_guid0[50]));
Q_AN02 U3615 ( .A0(n158), .A1(guid0[50]), .Z(n1253));
Q_MX02 U3616 ( .S(n388), .A0(n1254), .A1(stitcher_out[9]), .Z(nxt_guid0[49]));
Q_AN02 U3617 ( .A0(n158), .A1(guid0[49]), .Z(n1254));
Q_MX02 U3618 ( .S(n388), .A0(n1255), .A1(stitcher_out[8]), .Z(nxt_guid0[48]));
Q_AN02 U3619 ( .A0(n158), .A1(guid0[48]), .Z(n1255));
Q_MX02 U3620 ( .S(n388), .A0(n1256), .A1(stitcher_out[23]), .Z(nxt_guid0[47]));
Q_AN02 U3621 ( .A0(n158), .A1(guid0[47]), .Z(n1256));
Q_MX02 U3622 ( .S(n388), .A0(n1257), .A1(stitcher_out[22]), .Z(nxt_guid0[46]));
Q_AN02 U3623 ( .A0(n158), .A1(guid0[46]), .Z(n1257));
Q_MX02 U3624 ( .S(n388), .A0(n1258), .A1(stitcher_out[21]), .Z(nxt_guid0[45]));
Q_AN02 U3625 ( .A0(n158), .A1(guid0[45]), .Z(n1258));
Q_MX02 U3626 ( .S(n388), .A0(n1259), .A1(stitcher_out[20]), .Z(nxt_guid0[44]));
Q_AN02 U3627 ( .A0(n158), .A1(guid0[44]), .Z(n1259));
Q_MX02 U3628 ( .S(n388), .A0(n1260), .A1(stitcher_out[19]), .Z(nxt_guid0[43]));
Q_AN02 U3629 ( .A0(n158), .A1(guid0[43]), .Z(n1260));
Q_MX02 U3630 ( .S(n388), .A0(n1261), .A1(stitcher_out[18]), .Z(nxt_guid0[42]));
Q_AN02 U3631 ( .A0(n158), .A1(guid0[42]), .Z(n1261));
Q_MX02 U3632 ( .S(n388), .A0(n1262), .A1(stitcher_out[17]), .Z(nxt_guid0[41]));
Q_AN02 U3633 ( .A0(n158), .A1(guid0[41]), .Z(n1262));
Q_MX02 U3634 ( .S(n388), .A0(n1263), .A1(stitcher_out[16]), .Z(nxt_guid0[40]));
Q_AN02 U3635 ( .A0(n158), .A1(guid0[40]), .Z(n1263));
Q_MX02 U3636 ( .S(n388), .A0(n1264), .A1(stitcher_out[31]), .Z(nxt_guid0[39]));
Q_AN02 U3637 ( .A0(n158), .A1(guid0[39]), .Z(n1264));
Q_MX02 U3638 ( .S(n388), .A0(n1265), .A1(stitcher_out[30]), .Z(nxt_guid0[38]));
Q_AN02 U3639 ( .A0(n158), .A1(guid0[38]), .Z(n1265));
Q_MX02 U3640 ( .S(n388), .A0(n1266), .A1(stitcher_out[29]), .Z(nxt_guid0[37]));
Q_AN02 U3641 ( .A0(n158), .A1(guid0[37]), .Z(n1266));
Q_MX02 U3642 ( .S(n388), .A0(n1267), .A1(stitcher_out[28]), .Z(nxt_guid0[36]));
Q_AN02 U3643 ( .A0(n158), .A1(guid0[36]), .Z(n1267));
Q_MX02 U3644 ( .S(n388), .A0(n1268), .A1(stitcher_out[27]), .Z(nxt_guid0[35]));
Q_AN02 U3645 ( .A0(n158), .A1(guid0[35]), .Z(n1268));
Q_MX02 U3646 ( .S(n388), .A0(n1269), .A1(stitcher_out[26]), .Z(nxt_guid0[34]));
Q_AN02 U3647 ( .A0(n158), .A1(guid0[34]), .Z(n1269));
Q_MX02 U3648 ( .S(n388), .A0(n1270), .A1(stitcher_out[25]), .Z(nxt_guid0[33]));
Q_AN02 U3649 ( .A0(n158), .A1(guid0[33]), .Z(n1270));
Q_MX02 U3650 ( .S(n388), .A0(n1271), .A1(stitcher_out[24]), .Z(nxt_guid0[32]));
Q_AN02 U3651 ( .A0(n158), .A1(guid0[32]), .Z(n1271));
Q_MX02 U3652 ( .S(n388), .A0(n1272), .A1(stitcher_out[39]), .Z(nxt_guid0[31]));
Q_AN02 U3653 ( .A0(n158), .A1(guid0[31]), .Z(n1272));
Q_MX02 U3654 ( .S(n388), .A0(n1273), .A1(stitcher_out[38]), .Z(nxt_guid0[30]));
Q_AN02 U3655 ( .A0(n158), .A1(guid0[30]), .Z(n1273));
Q_MX02 U3656 ( .S(n388), .A0(n1274), .A1(stitcher_out[37]), .Z(nxt_guid0[29]));
Q_AN02 U3657 ( .A0(n158), .A1(guid0[29]), .Z(n1274));
Q_MX02 U3658 ( .S(n388), .A0(n1275), .A1(stitcher_out[36]), .Z(nxt_guid0[28]));
Q_AN02 U3659 ( .A0(n158), .A1(guid0[28]), .Z(n1275));
Q_MX02 U3660 ( .S(n388), .A0(n1276), .A1(stitcher_out[35]), .Z(nxt_guid0[27]));
Q_AN02 U3661 ( .A0(n158), .A1(guid0[27]), .Z(n1276));
Q_MX02 U3662 ( .S(n388), .A0(n1277), .A1(stitcher_out[34]), .Z(nxt_guid0[26]));
Q_AN02 U3663 ( .A0(n158), .A1(guid0[26]), .Z(n1277));
Q_MX02 U3664 ( .S(n388), .A0(n1278), .A1(stitcher_out[33]), .Z(nxt_guid0[25]));
Q_AN02 U3665 ( .A0(n158), .A1(guid0[25]), .Z(n1278));
Q_MX02 U3666 ( .S(n388), .A0(n1279), .A1(stitcher_out[32]), .Z(nxt_guid0[24]));
Q_AN02 U3667 ( .A0(n158), .A1(guid0[24]), .Z(n1279));
Q_MX02 U3668 ( .S(n388), .A0(n1280), .A1(stitcher_out[47]), .Z(nxt_guid0[23]));
Q_AN02 U3669 ( .A0(n158), .A1(guid0[23]), .Z(n1280));
Q_MX02 U3670 ( .S(n388), .A0(n1281), .A1(stitcher_out[46]), .Z(nxt_guid0[22]));
Q_AN02 U3671 ( .A0(n158), .A1(guid0[22]), .Z(n1281));
Q_MX02 U3672 ( .S(n388), .A0(n1282), .A1(stitcher_out[45]), .Z(nxt_guid0[21]));
Q_AN02 U3673 ( .A0(n158), .A1(guid0[21]), .Z(n1282));
Q_MX02 U3674 ( .S(n388), .A0(n1283), .A1(stitcher_out[44]), .Z(nxt_guid0[20]));
Q_AN02 U3675 ( .A0(n158), .A1(guid0[20]), .Z(n1283));
Q_MX02 U3676 ( .S(n388), .A0(n1284), .A1(stitcher_out[43]), .Z(nxt_guid0[19]));
Q_AN02 U3677 ( .A0(n158), .A1(guid0[19]), .Z(n1284));
Q_MX02 U3678 ( .S(n388), .A0(n1285), .A1(stitcher_out[42]), .Z(nxt_guid0[18]));
Q_AN02 U3679 ( .A0(n158), .A1(guid0[18]), .Z(n1285));
Q_MX02 U3680 ( .S(n388), .A0(n1286), .A1(stitcher_out[41]), .Z(nxt_guid0[17]));
Q_AN02 U3681 ( .A0(n158), .A1(guid0[17]), .Z(n1286));
Q_MX02 U3682 ( .S(n388), .A0(n1287), .A1(stitcher_out[40]), .Z(nxt_guid0[16]));
Q_AN02 U3683 ( .A0(n158), .A1(guid0[16]), .Z(n1287));
Q_MX02 U3684 ( .S(n388), .A0(n1288), .A1(stitcher_out[55]), .Z(nxt_guid0[15]));
Q_AN02 U3685 ( .A0(n158), .A1(guid0[15]), .Z(n1288));
Q_MX02 U3686 ( .S(n388), .A0(n1289), .A1(stitcher_out[54]), .Z(nxt_guid0[14]));
Q_AN02 U3687 ( .A0(n158), .A1(guid0[14]), .Z(n1289));
Q_MX02 U3688 ( .S(n388), .A0(n1290), .A1(stitcher_out[53]), .Z(nxt_guid0[13]));
Q_AN02 U3689 ( .A0(n158), .A1(guid0[13]), .Z(n1290));
Q_MX02 U3690 ( .S(n388), .A0(n1291), .A1(stitcher_out[52]), .Z(nxt_guid0[12]));
Q_AN02 U3691 ( .A0(n158), .A1(guid0[12]), .Z(n1291));
Q_MX02 U3692 ( .S(n388), .A0(n1292), .A1(stitcher_out[51]), .Z(nxt_guid0[11]));
Q_AN02 U3693 ( .A0(n158), .A1(guid0[11]), .Z(n1292));
Q_MX02 U3694 ( .S(n388), .A0(n1293), .A1(stitcher_out[50]), .Z(nxt_guid0[10]));
Q_AN02 U3695 ( .A0(n158), .A1(guid0[10]), .Z(n1293));
Q_MX02 U3696 ( .S(n388), .A0(n1294), .A1(stitcher_out[49]), .Z(nxt_guid0[9]));
Q_AN02 U3697 ( .A0(n158), .A1(guid0[9]), .Z(n1294));
Q_MX02 U3698 ( .S(n388), .A0(n1295), .A1(stitcher_out[48]), .Z(nxt_guid0[8]));
Q_AN02 U3699 ( .A0(n158), .A1(guid0[8]), .Z(n1295));
Q_MX02 U3700 ( .S(n388), .A0(n1296), .A1(stitcher_out[63]), .Z(nxt_guid0[7]));
Q_AN02 U3701 ( .A0(n158), .A1(guid0[7]), .Z(n1296));
Q_MX02 U3702 ( .S(n388), .A0(n1297), .A1(stitcher_out[62]), .Z(nxt_guid0[6]));
Q_AN02 U3703 ( .A0(n158), .A1(guid0[6]), .Z(n1297));
Q_MX02 U3704 ( .S(n388), .A0(n1298), .A1(stitcher_out[61]), .Z(nxt_guid0[5]));
Q_AN02 U3705 ( .A0(n158), .A1(guid0[5]), .Z(n1298));
Q_MX02 U3706 ( .S(n388), .A0(n1299), .A1(stitcher_out[60]), .Z(nxt_guid0[4]));
Q_AN02 U3707 ( .A0(n158), .A1(guid0[4]), .Z(n1299));
Q_MX02 U3708 ( .S(n388), .A0(n1300), .A1(stitcher_out[59]), .Z(nxt_guid0[3]));
Q_AN02 U3709 ( .A0(n158), .A1(guid0[3]), .Z(n1300));
Q_MX02 U3710 ( .S(n388), .A0(n1301), .A1(stitcher_out[58]), .Z(nxt_guid0[2]));
Q_AN02 U3711 ( .A0(n158), .A1(guid0[2]), .Z(n1301));
Q_MX02 U3712 ( .S(n388), .A0(n1302), .A1(stitcher_out[57]), .Z(nxt_guid0[1]));
Q_AN02 U3713 ( .A0(n158), .A1(guid0[1]), .Z(n1302));
Q_MX02 U3714 ( .S(n388), .A0(n1303), .A1(stitcher_out[56]), .Z(nxt_guid0[0]));
Q_AN02 U3715 ( .A0(n158), .A1(guid0[0]), .Z(n1303));
Q_MX02 U3716 ( .S(n391), .A0(n1304), .A1(stitcher_out[7]), .Z(nxt_guid1[63]));
Q_AN02 U3717 ( .A0(n159), .A1(guid1[63]), .Z(n1304));
Q_MX02 U3718 ( .S(n391), .A0(n1305), .A1(stitcher_out[6]), .Z(nxt_guid1[62]));
Q_AN02 U3719 ( .A0(n159), .A1(guid1[62]), .Z(n1305));
Q_MX02 U3720 ( .S(n391), .A0(n1306), .A1(stitcher_out[5]), .Z(nxt_guid1[61]));
Q_AN02 U3721 ( .A0(n159), .A1(guid1[61]), .Z(n1306));
Q_MX02 U3722 ( .S(n391), .A0(n1307), .A1(stitcher_out[4]), .Z(nxt_guid1[60]));
Q_AN02 U3723 ( .A0(n159), .A1(guid1[60]), .Z(n1307));
Q_MX02 U3724 ( .S(n391), .A0(n1308), .A1(stitcher_out[3]), .Z(nxt_guid1[59]));
Q_AN02 U3725 ( .A0(n159), .A1(guid1[59]), .Z(n1308));
Q_MX02 U3726 ( .S(n391), .A0(n1309), .A1(stitcher_out[2]), .Z(nxt_guid1[58]));
Q_AN02 U3727 ( .A0(n159), .A1(guid1[58]), .Z(n1309));
Q_MX02 U3728 ( .S(n391), .A0(n1310), .A1(stitcher_out[1]), .Z(nxt_guid1[57]));
Q_AN02 U3729 ( .A0(n159), .A1(guid1[57]), .Z(n1310));
Q_MX02 U3730 ( .S(n391), .A0(n1311), .A1(stitcher_out[0]), .Z(nxt_guid1[56]));
Q_AN02 U3731 ( .A0(n159), .A1(guid1[56]), .Z(n1311));
Q_MX02 U3732 ( .S(n391), .A0(n1312), .A1(stitcher_out[15]), .Z(nxt_guid1[55]));
Q_AN02 U3733 ( .A0(n159), .A1(guid1[55]), .Z(n1312));
Q_MX02 U3734 ( .S(n391), .A0(n1313), .A1(stitcher_out[14]), .Z(nxt_guid1[54]));
Q_AN02 U3735 ( .A0(n159), .A1(guid1[54]), .Z(n1313));
Q_MX02 U3736 ( .S(n391), .A0(n1314), .A1(stitcher_out[13]), .Z(nxt_guid1[53]));
Q_AN02 U3737 ( .A0(n159), .A1(guid1[53]), .Z(n1314));
Q_MX02 U3738 ( .S(n391), .A0(n1315), .A1(stitcher_out[12]), .Z(nxt_guid1[52]));
Q_AN02 U3739 ( .A0(n159), .A1(guid1[52]), .Z(n1315));
Q_MX02 U3740 ( .S(n391), .A0(n1316), .A1(stitcher_out[11]), .Z(nxt_guid1[51]));
Q_AN02 U3741 ( .A0(n159), .A1(guid1[51]), .Z(n1316));
Q_MX02 U3742 ( .S(n391), .A0(n1317), .A1(stitcher_out[10]), .Z(nxt_guid1[50]));
Q_AN02 U3743 ( .A0(n159), .A1(guid1[50]), .Z(n1317));
Q_MX02 U3744 ( .S(n391), .A0(n1318), .A1(stitcher_out[9]), .Z(nxt_guid1[49]));
Q_AN02 U3745 ( .A0(n159), .A1(guid1[49]), .Z(n1318));
Q_MX02 U3746 ( .S(n391), .A0(n1319), .A1(stitcher_out[8]), .Z(nxt_guid1[48]));
Q_AN02 U3747 ( .A0(n159), .A1(guid1[48]), .Z(n1319));
Q_MX02 U3748 ( .S(n391), .A0(n1320), .A1(stitcher_out[23]), .Z(nxt_guid1[47]));
Q_AN02 U3749 ( .A0(n159), .A1(guid1[47]), .Z(n1320));
Q_MX02 U3750 ( .S(n391), .A0(n1321), .A1(stitcher_out[22]), .Z(nxt_guid1[46]));
Q_AN02 U3751 ( .A0(n159), .A1(guid1[46]), .Z(n1321));
Q_MX02 U3752 ( .S(n391), .A0(n1322), .A1(stitcher_out[21]), .Z(nxt_guid1[45]));
Q_AN02 U3753 ( .A0(n159), .A1(guid1[45]), .Z(n1322));
Q_MX02 U3754 ( .S(n391), .A0(n1323), .A1(stitcher_out[20]), .Z(nxt_guid1[44]));
Q_AN02 U3755 ( .A0(n159), .A1(guid1[44]), .Z(n1323));
Q_MX02 U3756 ( .S(n391), .A0(n1324), .A1(stitcher_out[19]), .Z(nxt_guid1[43]));
Q_AN02 U3757 ( .A0(n159), .A1(guid1[43]), .Z(n1324));
Q_MX02 U3758 ( .S(n391), .A0(n1325), .A1(stitcher_out[18]), .Z(nxt_guid1[42]));
Q_AN02 U3759 ( .A0(n159), .A1(guid1[42]), .Z(n1325));
Q_MX02 U3760 ( .S(n391), .A0(n1326), .A1(stitcher_out[17]), .Z(nxt_guid1[41]));
Q_AN02 U3761 ( .A0(n159), .A1(guid1[41]), .Z(n1326));
Q_MX02 U3762 ( .S(n391), .A0(n1327), .A1(stitcher_out[16]), .Z(nxt_guid1[40]));
Q_AN02 U3763 ( .A0(n159), .A1(guid1[40]), .Z(n1327));
Q_MX02 U3764 ( .S(n391), .A0(n1328), .A1(stitcher_out[31]), .Z(nxt_guid1[39]));
Q_AN02 U3765 ( .A0(n159), .A1(guid1[39]), .Z(n1328));
Q_MX02 U3766 ( .S(n391), .A0(n1329), .A1(stitcher_out[30]), .Z(nxt_guid1[38]));
Q_AN02 U3767 ( .A0(n159), .A1(guid1[38]), .Z(n1329));
Q_MX02 U3768 ( .S(n391), .A0(n1330), .A1(stitcher_out[29]), .Z(nxt_guid1[37]));
Q_AN02 U3769 ( .A0(n159), .A1(guid1[37]), .Z(n1330));
Q_MX02 U3770 ( .S(n391), .A0(n1331), .A1(stitcher_out[28]), .Z(nxt_guid1[36]));
Q_AN02 U3771 ( .A0(n159), .A1(guid1[36]), .Z(n1331));
Q_MX02 U3772 ( .S(n391), .A0(n1332), .A1(stitcher_out[27]), .Z(nxt_guid1[35]));
Q_AN02 U3773 ( .A0(n159), .A1(guid1[35]), .Z(n1332));
Q_MX02 U3774 ( .S(n391), .A0(n1333), .A1(stitcher_out[26]), .Z(nxt_guid1[34]));
Q_AN02 U3775 ( .A0(n159), .A1(guid1[34]), .Z(n1333));
Q_MX02 U3776 ( .S(n391), .A0(n1334), .A1(stitcher_out[25]), .Z(nxt_guid1[33]));
Q_AN02 U3777 ( .A0(n159), .A1(guid1[33]), .Z(n1334));
Q_MX02 U3778 ( .S(n391), .A0(n1335), .A1(stitcher_out[24]), .Z(nxt_guid1[32]));
Q_AN02 U3779 ( .A0(n159), .A1(guid1[32]), .Z(n1335));
Q_MX02 U3780 ( .S(n391), .A0(n1336), .A1(stitcher_out[39]), .Z(nxt_guid1[31]));
Q_AN02 U3781 ( .A0(n159), .A1(guid1[31]), .Z(n1336));
Q_MX02 U3782 ( .S(n391), .A0(n1337), .A1(stitcher_out[38]), .Z(nxt_guid1[30]));
Q_AN02 U3783 ( .A0(n159), .A1(guid1[30]), .Z(n1337));
Q_MX02 U3784 ( .S(n391), .A0(n1338), .A1(stitcher_out[37]), .Z(nxt_guid1[29]));
Q_AN02 U3785 ( .A0(n159), .A1(guid1[29]), .Z(n1338));
Q_MX02 U3786 ( .S(n391), .A0(n1339), .A1(stitcher_out[36]), .Z(nxt_guid1[28]));
Q_AN02 U3787 ( .A0(n159), .A1(guid1[28]), .Z(n1339));
Q_MX02 U3788 ( .S(n391), .A0(n1340), .A1(stitcher_out[35]), .Z(nxt_guid1[27]));
Q_AN02 U3789 ( .A0(n159), .A1(guid1[27]), .Z(n1340));
Q_MX02 U3790 ( .S(n391), .A0(n1341), .A1(stitcher_out[34]), .Z(nxt_guid1[26]));
Q_AN02 U3791 ( .A0(n159), .A1(guid1[26]), .Z(n1341));
Q_MX02 U3792 ( .S(n391), .A0(n1342), .A1(stitcher_out[33]), .Z(nxt_guid1[25]));
Q_AN02 U3793 ( .A0(n159), .A1(guid1[25]), .Z(n1342));
Q_MX02 U3794 ( .S(n391), .A0(n1343), .A1(stitcher_out[32]), .Z(nxt_guid1[24]));
Q_AN02 U3795 ( .A0(n159), .A1(guid1[24]), .Z(n1343));
Q_MX02 U3796 ( .S(n391), .A0(n1344), .A1(stitcher_out[47]), .Z(nxt_guid1[23]));
Q_AN02 U3797 ( .A0(n159), .A1(guid1[23]), .Z(n1344));
Q_MX02 U3798 ( .S(n391), .A0(n1345), .A1(stitcher_out[46]), .Z(nxt_guid1[22]));
Q_AN02 U3799 ( .A0(n159), .A1(guid1[22]), .Z(n1345));
Q_MX02 U3800 ( .S(n391), .A0(n1346), .A1(stitcher_out[45]), .Z(nxt_guid1[21]));
Q_AN02 U3801 ( .A0(n159), .A1(guid1[21]), .Z(n1346));
Q_MX02 U3802 ( .S(n391), .A0(n1347), .A1(stitcher_out[44]), .Z(nxt_guid1[20]));
Q_AN02 U3803 ( .A0(n159), .A1(guid1[20]), .Z(n1347));
Q_MX02 U3804 ( .S(n391), .A0(n1348), .A1(stitcher_out[43]), .Z(nxt_guid1[19]));
Q_AN02 U3805 ( .A0(n159), .A1(guid1[19]), .Z(n1348));
Q_MX02 U3806 ( .S(n391), .A0(n1349), .A1(stitcher_out[42]), .Z(nxt_guid1[18]));
Q_AN02 U3807 ( .A0(n159), .A1(guid1[18]), .Z(n1349));
Q_MX02 U3808 ( .S(n391), .A0(n1350), .A1(stitcher_out[41]), .Z(nxt_guid1[17]));
Q_AN02 U3809 ( .A0(n159), .A1(guid1[17]), .Z(n1350));
Q_MX02 U3810 ( .S(n391), .A0(n1351), .A1(stitcher_out[40]), .Z(nxt_guid1[16]));
Q_AN02 U3811 ( .A0(n159), .A1(guid1[16]), .Z(n1351));
Q_MX02 U3812 ( .S(n391), .A0(n1352), .A1(stitcher_out[55]), .Z(nxt_guid1[15]));
Q_AN02 U3813 ( .A0(n159), .A1(guid1[15]), .Z(n1352));
Q_MX02 U3814 ( .S(n391), .A0(n1353), .A1(stitcher_out[54]), .Z(nxt_guid1[14]));
Q_AN02 U3815 ( .A0(n159), .A1(guid1[14]), .Z(n1353));
Q_MX02 U3816 ( .S(n391), .A0(n1354), .A1(stitcher_out[53]), .Z(nxt_guid1[13]));
Q_AN02 U3817 ( .A0(n159), .A1(guid1[13]), .Z(n1354));
Q_MX02 U3818 ( .S(n391), .A0(n1355), .A1(stitcher_out[52]), .Z(nxt_guid1[12]));
Q_AN02 U3819 ( .A0(n159), .A1(guid1[12]), .Z(n1355));
Q_MX02 U3820 ( .S(n391), .A0(n1356), .A1(stitcher_out[51]), .Z(nxt_guid1[11]));
Q_AN02 U3821 ( .A0(n159), .A1(guid1[11]), .Z(n1356));
Q_MX02 U3822 ( .S(n391), .A0(n1357), .A1(stitcher_out[50]), .Z(nxt_guid1[10]));
Q_AN02 U3823 ( .A0(n159), .A1(guid1[10]), .Z(n1357));
Q_MX02 U3824 ( .S(n391), .A0(n1358), .A1(stitcher_out[49]), .Z(nxt_guid1[9]));
Q_AN02 U3825 ( .A0(n159), .A1(guid1[9]), .Z(n1358));
Q_MX02 U3826 ( .S(n391), .A0(n1359), .A1(stitcher_out[48]), .Z(nxt_guid1[8]));
Q_AN02 U3827 ( .A0(n159), .A1(guid1[8]), .Z(n1359));
Q_MX02 U3828 ( .S(n391), .A0(n1360), .A1(stitcher_out[63]), .Z(nxt_guid1[7]));
Q_AN02 U3829 ( .A0(n159), .A1(guid1[7]), .Z(n1360));
Q_MX02 U3830 ( .S(n391), .A0(n1361), .A1(stitcher_out[62]), .Z(nxt_guid1[6]));
Q_AN02 U3831 ( .A0(n159), .A1(guid1[6]), .Z(n1361));
Q_MX02 U3832 ( .S(n391), .A0(n1362), .A1(stitcher_out[61]), .Z(nxt_guid1[5]));
Q_AN02 U3833 ( .A0(n159), .A1(guid1[5]), .Z(n1362));
Q_MX02 U3834 ( .S(n391), .A0(n1363), .A1(stitcher_out[60]), .Z(nxt_guid1[4]));
Q_AN02 U3835 ( .A0(n159), .A1(guid1[4]), .Z(n1363));
Q_MX02 U3836 ( .S(n391), .A0(n1364), .A1(stitcher_out[59]), .Z(nxt_guid1[3]));
Q_AN02 U3837 ( .A0(n159), .A1(guid1[3]), .Z(n1364));
Q_MX02 U3838 ( .S(n391), .A0(n1365), .A1(stitcher_out[58]), .Z(nxt_guid1[2]));
Q_AN02 U3839 ( .A0(n159), .A1(guid1[2]), .Z(n1365));
Q_MX02 U3840 ( .S(n391), .A0(n1366), .A1(stitcher_out[57]), .Z(nxt_guid1[1]));
Q_AN02 U3841 ( .A0(n159), .A1(guid1[1]), .Z(n1366));
Q_MX02 U3842 ( .S(n391), .A0(n1367), .A1(stitcher_out[56]), .Z(nxt_guid1[0]));
Q_AN02 U3843 ( .A0(n159), .A1(guid1[0]), .Z(n1367));
Q_MX02 U3844 ( .S(n396), .A0(n1368), .A1(stitcher_out[7]), .Z(nxt_guid2[63]));
Q_AN02 U3845 ( .A0(n160), .A1(guid2[63]), .Z(n1368));
Q_MX02 U3846 ( .S(n396), .A0(n1369), .A1(stitcher_out[6]), .Z(nxt_guid2[62]));
Q_AN02 U3847 ( .A0(n160), .A1(guid2[62]), .Z(n1369));
Q_MX02 U3848 ( .S(n396), .A0(n1370), .A1(stitcher_out[5]), .Z(nxt_guid2[61]));
Q_AN02 U3849 ( .A0(n160), .A1(guid2[61]), .Z(n1370));
Q_MX02 U3850 ( .S(n396), .A0(n1371), .A1(stitcher_out[4]), .Z(nxt_guid2[60]));
Q_AN02 U3851 ( .A0(n160), .A1(guid2[60]), .Z(n1371));
Q_MX02 U3852 ( .S(n396), .A0(n1372), .A1(stitcher_out[3]), .Z(nxt_guid2[59]));
Q_AN02 U3853 ( .A0(n160), .A1(guid2[59]), .Z(n1372));
Q_MX02 U3854 ( .S(n396), .A0(n1373), .A1(stitcher_out[2]), .Z(nxt_guid2[58]));
Q_AN02 U3855 ( .A0(n160), .A1(guid2[58]), .Z(n1373));
Q_MX02 U3856 ( .S(n396), .A0(n1374), .A1(stitcher_out[1]), .Z(nxt_guid2[57]));
Q_AN02 U3857 ( .A0(n160), .A1(guid2[57]), .Z(n1374));
Q_MX02 U3858 ( .S(n396), .A0(n1375), .A1(stitcher_out[0]), .Z(nxt_guid2[56]));
Q_AN02 U3859 ( .A0(n160), .A1(guid2[56]), .Z(n1375));
Q_MX02 U3860 ( .S(n396), .A0(n1376), .A1(stitcher_out[15]), .Z(nxt_guid2[55]));
Q_AN02 U3861 ( .A0(n160), .A1(guid2[55]), .Z(n1376));
Q_MX02 U3862 ( .S(n396), .A0(n1377), .A1(stitcher_out[14]), .Z(nxt_guid2[54]));
Q_AN02 U3863 ( .A0(n160), .A1(guid2[54]), .Z(n1377));
Q_MX02 U3864 ( .S(n396), .A0(n1378), .A1(stitcher_out[13]), .Z(nxt_guid2[53]));
Q_AN02 U3865 ( .A0(n160), .A1(guid2[53]), .Z(n1378));
Q_MX02 U3866 ( .S(n396), .A0(n1379), .A1(stitcher_out[12]), .Z(nxt_guid2[52]));
Q_AN02 U3867 ( .A0(n160), .A1(guid2[52]), .Z(n1379));
Q_MX02 U3868 ( .S(n396), .A0(n1380), .A1(stitcher_out[11]), .Z(nxt_guid2[51]));
Q_AN02 U3869 ( .A0(n160), .A1(guid2[51]), .Z(n1380));
Q_MX02 U3870 ( .S(n396), .A0(n1381), .A1(stitcher_out[10]), .Z(nxt_guid2[50]));
Q_AN02 U3871 ( .A0(n160), .A1(guid2[50]), .Z(n1381));
Q_MX02 U3872 ( .S(n396), .A0(n1382), .A1(stitcher_out[9]), .Z(nxt_guid2[49]));
Q_AN02 U3873 ( .A0(n160), .A1(guid2[49]), .Z(n1382));
Q_MX02 U3874 ( .S(n396), .A0(n1383), .A1(stitcher_out[8]), .Z(nxt_guid2[48]));
Q_AN02 U3875 ( .A0(n160), .A1(guid2[48]), .Z(n1383));
Q_MX02 U3876 ( .S(n396), .A0(n1384), .A1(stitcher_out[23]), .Z(nxt_guid2[47]));
Q_AN02 U3877 ( .A0(n160), .A1(guid2[47]), .Z(n1384));
Q_MX02 U3878 ( .S(n396), .A0(n1385), .A1(stitcher_out[22]), .Z(nxt_guid2[46]));
Q_AN02 U3879 ( .A0(n160), .A1(guid2[46]), .Z(n1385));
Q_MX02 U3880 ( .S(n396), .A0(n1386), .A1(stitcher_out[21]), .Z(nxt_guid2[45]));
Q_AN02 U3881 ( .A0(n160), .A1(guid2[45]), .Z(n1386));
Q_MX02 U3882 ( .S(n396), .A0(n1387), .A1(stitcher_out[20]), .Z(nxt_guid2[44]));
Q_AN02 U3883 ( .A0(n160), .A1(guid2[44]), .Z(n1387));
Q_MX02 U3884 ( .S(n396), .A0(n1388), .A1(stitcher_out[19]), .Z(nxt_guid2[43]));
Q_AN02 U3885 ( .A0(n160), .A1(guid2[43]), .Z(n1388));
Q_MX02 U3886 ( .S(n396), .A0(n1389), .A1(stitcher_out[18]), .Z(nxt_guid2[42]));
Q_AN02 U3887 ( .A0(n160), .A1(guid2[42]), .Z(n1389));
Q_MX02 U3888 ( .S(n396), .A0(n1390), .A1(stitcher_out[17]), .Z(nxt_guid2[41]));
Q_AN02 U3889 ( .A0(n160), .A1(guid2[41]), .Z(n1390));
Q_MX02 U3890 ( .S(n396), .A0(n1391), .A1(stitcher_out[16]), .Z(nxt_guid2[40]));
Q_AN02 U3891 ( .A0(n160), .A1(guid2[40]), .Z(n1391));
Q_MX02 U3892 ( .S(n396), .A0(n1392), .A1(stitcher_out[31]), .Z(nxt_guid2[39]));
Q_AN02 U3893 ( .A0(n160), .A1(guid2[39]), .Z(n1392));
Q_MX02 U3894 ( .S(n396), .A0(n1393), .A1(stitcher_out[30]), .Z(nxt_guid2[38]));
Q_AN02 U3895 ( .A0(n160), .A1(guid2[38]), .Z(n1393));
Q_MX02 U3896 ( .S(n396), .A0(n1394), .A1(stitcher_out[29]), .Z(nxt_guid2[37]));
Q_AN02 U3897 ( .A0(n160), .A1(guid2[37]), .Z(n1394));
Q_MX02 U3898 ( .S(n396), .A0(n1395), .A1(stitcher_out[28]), .Z(nxt_guid2[36]));
Q_AN02 U3899 ( .A0(n160), .A1(guid2[36]), .Z(n1395));
Q_MX02 U3900 ( .S(n396), .A0(n1396), .A1(stitcher_out[27]), .Z(nxt_guid2[35]));
Q_AN02 U3901 ( .A0(n160), .A1(guid2[35]), .Z(n1396));
Q_MX02 U3902 ( .S(n396), .A0(n1397), .A1(stitcher_out[26]), .Z(nxt_guid2[34]));
Q_AN02 U3903 ( .A0(n160), .A1(guid2[34]), .Z(n1397));
Q_MX02 U3904 ( .S(n396), .A0(n1398), .A1(stitcher_out[25]), .Z(nxt_guid2[33]));
Q_AN02 U3905 ( .A0(n160), .A1(guid2[33]), .Z(n1398));
Q_MX02 U3906 ( .S(n396), .A0(n1399), .A1(stitcher_out[24]), .Z(nxt_guid2[32]));
Q_AN02 U3907 ( .A0(n160), .A1(guid2[32]), .Z(n1399));
Q_MX02 U3908 ( .S(n396), .A0(n1400), .A1(stitcher_out[39]), .Z(nxt_guid2[31]));
Q_AN02 U3909 ( .A0(n160), .A1(guid2[31]), .Z(n1400));
Q_MX02 U3910 ( .S(n396), .A0(n1401), .A1(stitcher_out[38]), .Z(nxt_guid2[30]));
Q_AN02 U3911 ( .A0(n160), .A1(guid2[30]), .Z(n1401));
Q_MX02 U3912 ( .S(n396), .A0(n1402), .A1(stitcher_out[37]), .Z(nxt_guid2[29]));
Q_AN02 U3913 ( .A0(n160), .A1(guid2[29]), .Z(n1402));
Q_MX02 U3914 ( .S(n396), .A0(n1403), .A1(stitcher_out[36]), .Z(nxt_guid2[28]));
Q_AN02 U3915 ( .A0(n160), .A1(guid2[28]), .Z(n1403));
Q_MX02 U3916 ( .S(n396), .A0(n1404), .A1(stitcher_out[35]), .Z(nxt_guid2[27]));
Q_AN02 U3917 ( .A0(n160), .A1(guid2[27]), .Z(n1404));
Q_MX02 U3918 ( .S(n396), .A0(n1405), .A1(stitcher_out[34]), .Z(nxt_guid2[26]));
Q_AN02 U3919 ( .A0(n160), .A1(guid2[26]), .Z(n1405));
Q_MX02 U3920 ( .S(n396), .A0(n1406), .A1(stitcher_out[33]), .Z(nxt_guid2[25]));
Q_AN02 U3921 ( .A0(n160), .A1(guid2[25]), .Z(n1406));
Q_MX02 U3922 ( .S(n396), .A0(n1407), .A1(stitcher_out[32]), .Z(nxt_guid2[24]));
Q_AN02 U3923 ( .A0(n160), .A1(guid2[24]), .Z(n1407));
Q_MX02 U3924 ( .S(n396), .A0(n1408), .A1(stitcher_out[47]), .Z(nxt_guid2[23]));
Q_AN02 U3925 ( .A0(n160), .A1(guid2[23]), .Z(n1408));
Q_MX02 U3926 ( .S(n396), .A0(n1409), .A1(stitcher_out[46]), .Z(nxt_guid2[22]));
Q_AN02 U3927 ( .A0(n160), .A1(guid2[22]), .Z(n1409));
Q_MX02 U3928 ( .S(n396), .A0(n1410), .A1(stitcher_out[45]), .Z(nxt_guid2[21]));
Q_AN02 U3929 ( .A0(n160), .A1(guid2[21]), .Z(n1410));
Q_MX02 U3930 ( .S(n396), .A0(n1411), .A1(stitcher_out[44]), .Z(nxt_guid2[20]));
Q_AN02 U3931 ( .A0(n160), .A1(guid2[20]), .Z(n1411));
Q_MX02 U3932 ( .S(n396), .A0(n1412), .A1(stitcher_out[43]), .Z(nxt_guid2[19]));
Q_AN02 U3933 ( .A0(n160), .A1(guid2[19]), .Z(n1412));
Q_MX02 U3934 ( .S(n396), .A0(n1413), .A1(stitcher_out[42]), .Z(nxt_guid2[18]));
Q_AN02 U3935 ( .A0(n160), .A1(guid2[18]), .Z(n1413));
Q_MX02 U3936 ( .S(n396), .A0(n1414), .A1(stitcher_out[41]), .Z(nxt_guid2[17]));
Q_AN02 U3937 ( .A0(n160), .A1(guid2[17]), .Z(n1414));
Q_MX02 U3938 ( .S(n396), .A0(n1415), .A1(stitcher_out[40]), .Z(nxt_guid2[16]));
Q_AN02 U3939 ( .A0(n160), .A1(guid2[16]), .Z(n1415));
Q_MX02 U3940 ( .S(n396), .A0(n1416), .A1(stitcher_out[55]), .Z(nxt_guid2[15]));
Q_AN02 U3941 ( .A0(n160), .A1(guid2[15]), .Z(n1416));
Q_MX02 U3942 ( .S(n396), .A0(n1417), .A1(stitcher_out[54]), .Z(nxt_guid2[14]));
Q_AN02 U3943 ( .A0(n160), .A1(guid2[14]), .Z(n1417));
Q_MX02 U3944 ( .S(n396), .A0(n1418), .A1(stitcher_out[53]), .Z(nxt_guid2[13]));
Q_AN02 U3945 ( .A0(n160), .A1(guid2[13]), .Z(n1418));
Q_MX02 U3946 ( .S(n396), .A0(n1419), .A1(stitcher_out[52]), .Z(nxt_guid2[12]));
Q_AN02 U3947 ( .A0(n160), .A1(guid2[12]), .Z(n1419));
Q_MX02 U3948 ( .S(n396), .A0(n1420), .A1(stitcher_out[51]), .Z(nxt_guid2[11]));
Q_AN02 U3949 ( .A0(n160), .A1(guid2[11]), .Z(n1420));
Q_MX02 U3950 ( .S(n396), .A0(n1421), .A1(stitcher_out[50]), .Z(nxt_guid2[10]));
Q_AN02 U3951 ( .A0(n160), .A1(guid2[10]), .Z(n1421));
Q_MX02 U3952 ( .S(n396), .A0(n1422), .A1(stitcher_out[49]), .Z(nxt_guid2[9]));
Q_AN02 U3953 ( .A0(n160), .A1(guid2[9]), .Z(n1422));
Q_MX02 U3954 ( .S(n396), .A0(n1423), .A1(stitcher_out[48]), .Z(nxt_guid2[8]));
Q_AN02 U3955 ( .A0(n160), .A1(guid2[8]), .Z(n1423));
Q_MX02 U3956 ( .S(n396), .A0(n1424), .A1(stitcher_out[63]), .Z(nxt_guid2[7]));
Q_AN02 U3957 ( .A0(n160), .A1(guid2[7]), .Z(n1424));
Q_MX02 U3958 ( .S(n396), .A0(n1425), .A1(stitcher_out[62]), .Z(nxt_guid2[6]));
Q_AN02 U3959 ( .A0(n160), .A1(guid2[6]), .Z(n1425));
Q_MX02 U3960 ( .S(n396), .A0(n1426), .A1(stitcher_out[61]), .Z(nxt_guid2[5]));
Q_AN02 U3961 ( .A0(n160), .A1(guid2[5]), .Z(n1426));
Q_MX02 U3962 ( .S(n396), .A0(n1427), .A1(stitcher_out[60]), .Z(nxt_guid2[4]));
Q_AN02 U3963 ( .A0(n160), .A1(guid2[4]), .Z(n1427));
Q_MX02 U3964 ( .S(n396), .A0(n1428), .A1(stitcher_out[59]), .Z(nxt_guid2[3]));
Q_AN02 U3965 ( .A0(n160), .A1(guid2[3]), .Z(n1428));
Q_MX02 U3966 ( .S(n396), .A0(n1429), .A1(stitcher_out[58]), .Z(nxt_guid2[2]));
Q_AN02 U3967 ( .A0(n160), .A1(guid2[2]), .Z(n1429));
Q_MX02 U3968 ( .S(n396), .A0(n1430), .A1(stitcher_out[57]), .Z(nxt_guid2[1]));
Q_AN02 U3969 ( .A0(n160), .A1(guid2[1]), .Z(n1430));
Q_MX02 U3970 ( .S(n396), .A0(n1431), .A1(stitcher_out[56]), .Z(nxt_guid2[0]));
Q_AN02 U3971 ( .A0(n160), .A1(guid2[0]), .Z(n1431));
Q_MX02 U3972 ( .S(n401), .A0(n1432), .A1(stitcher_out[7]), .Z(nxt_guid3[63]));
Q_AN02 U3973 ( .A0(n161), .A1(guid3[63]), .Z(n1432));
Q_MX02 U3974 ( .S(n401), .A0(n1433), .A1(stitcher_out[6]), .Z(nxt_guid3[62]));
Q_AN02 U3975 ( .A0(n161), .A1(guid3[62]), .Z(n1433));
Q_MX02 U3976 ( .S(n401), .A0(n1434), .A1(stitcher_out[5]), .Z(nxt_guid3[61]));
Q_AN02 U3977 ( .A0(n161), .A1(guid3[61]), .Z(n1434));
Q_MX02 U3978 ( .S(n401), .A0(n1435), .A1(stitcher_out[4]), .Z(nxt_guid3[60]));
Q_AN02 U3979 ( .A0(n161), .A1(guid3[60]), .Z(n1435));
Q_MX02 U3980 ( .S(n401), .A0(n1436), .A1(stitcher_out[3]), .Z(nxt_guid3[59]));
Q_AN02 U3981 ( .A0(n161), .A1(guid3[59]), .Z(n1436));
Q_MX02 U3982 ( .S(n401), .A0(n1437), .A1(stitcher_out[2]), .Z(nxt_guid3[58]));
Q_AN02 U3983 ( .A0(n161), .A1(guid3[58]), .Z(n1437));
Q_MX02 U3984 ( .S(n401), .A0(n1438), .A1(stitcher_out[1]), .Z(nxt_guid3[57]));
Q_AN02 U3985 ( .A0(n161), .A1(guid3[57]), .Z(n1438));
Q_MX02 U3986 ( .S(n401), .A0(n1439), .A1(stitcher_out[0]), .Z(nxt_guid3[56]));
Q_AN02 U3987 ( .A0(n161), .A1(guid3[56]), .Z(n1439));
Q_MX02 U3988 ( .S(n401), .A0(n1440), .A1(stitcher_out[15]), .Z(nxt_guid3[55]));
Q_AN02 U3989 ( .A0(n161), .A1(guid3[55]), .Z(n1440));
Q_MX02 U3990 ( .S(n401), .A0(n1441), .A1(stitcher_out[14]), .Z(nxt_guid3[54]));
Q_AN02 U3991 ( .A0(n161), .A1(guid3[54]), .Z(n1441));
Q_MX02 U3992 ( .S(n401), .A0(n1442), .A1(stitcher_out[13]), .Z(nxt_guid3[53]));
Q_AN02 U3993 ( .A0(n161), .A1(guid3[53]), .Z(n1442));
Q_MX02 U3994 ( .S(n401), .A0(n1443), .A1(stitcher_out[12]), .Z(nxt_guid3[52]));
Q_AN02 U3995 ( .A0(n161), .A1(guid3[52]), .Z(n1443));
Q_MX02 U3996 ( .S(n401), .A0(n1444), .A1(stitcher_out[11]), .Z(nxt_guid3[51]));
Q_AN02 U3997 ( .A0(n161), .A1(guid3[51]), .Z(n1444));
Q_MX02 U3998 ( .S(n401), .A0(n1445), .A1(stitcher_out[10]), .Z(nxt_guid3[50]));
Q_AN02 U3999 ( .A0(n161), .A1(guid3[50]), .Z(n1445));
Q_MX02 U4000 ( .S(n401), .A0(n1446), .A1(stitcher_out[9]), .Z(nxt_guid3[49]));
Q_AN02 U4001 ( .A0(n161), .A1(guid3[49]), .Z(n1446));
Q_MX02 U4002 ( .S(n401), .A0(n1447), .A1(stitcher_out[8]), .Z(nxt_guid3[48]));
Q_AN02 U4003 ( .A0(n161), .A1(guid3[48]), .Z(n1447));
Q_MX02 U4004 ( .S(n401), .A0(n1448), .A1(stitcher_out[23]), .Z(nxt_guid3[47]));
Q_AN02 U4005 ( .A0(n161), .A1(guid3[47]), .Z(n1448));
Q_MX02 U4006 ( .S(n401), .A0(n1449), .A1(stitcher_out[22]), .Z(nxt_guid3[46]));
Q_AN02 U4007 ( .A0(n161), .A1(guid3[46]), .Z(n1449));
Q_MX02 U4008 ( .S(n401), .A0(n1450), .A1(stitcher_out[21]), .Z(nxt_guid3[45]));
Q_AN02 U4009 ( .A0(n161), .A1(guid3[45]), .Z(n1450));
Q_MX02 U4010 ( .S(n401), .A0(n1451), .A1(stitcher_out[20]), .Z(nxt_guid3[44]));
Q_AN02 U4011 ( .A0(n161), .A1(guid3[44]), .Z(n1451));
Q_MX02 U4012 ( .S(n401), .A0(n1452), .A1(stitcher_out[19]), .Z(nxt_guid3[43]));
Q_AN02 U4013 ( .A0(n161), .A1(guid3[43]), .Z(n1452));
Q_MX02 U4014 ( .S(n401), .A0(n1453), .A1(stitcher_out[18]), .Z(nxt_guid3[42]));
Q_AN02 U4015 ( .A0(n161), .A1(guid3[42]), .Z(n1453));
Q_MX02 U4016 ( .S(n401), .A0(n1454), .A1(stitcher_out[17]), .Z(nxt_guid3[41]));
Q_AN02 U4017 ( .A0(n161), .A1(guid3[41]), .Z(n1454));
Q_MX02 U4018 ( .S(n401), .A0(n1455), .A1(stitcher_out[16]), .Z(nxt_guid3[40]));
Q_AN02 U4019 ( .A0(n161), .A1(guid3[40]), .Z(n1455));
Q_MX02 U4020 ( .S(n401), .A0(n1456), .A1(stitcher_out[31]), .Z(nxt_guid3[39]));
Q_AN02 U4021 ( .A0(n161), .A1(guid3[39]), .Z(n1456));
Q_MX02 U4022 ( .S(n401), .A0(n1457), .A1(stitcher_out[30]), .Z(nxt_guid3[38]));
Q_AN02 U4023 ( .A0(n161), .A1(guid3[38]), .Z(n1457));
Q_MX02 U4024 ( .S(n401), .A0(n1458), .A1(stitcher_out[29]), .Z(nxt_guid3[37]));
Q_AN02 U4025 ( .A0(n161), .A1(guid3[37]), .Z(n1458));
Q_MX02 U4026 ( .S(n401), .A0(n1459), .A1(stitcher_out[28]), .Z(nxt_guid3[36]));
Q_AN02 U4027 ( .A0(n161), .A1(guid3[36]), .Z(n1459));
Q_MX02 U4028 ( .S(n401), .A0(n1460), .A1(stitcher_out[27]), .Z(nxt_guid3[35]));
Q_AN02 U4029 ( .A0(n161), .A1(guid3[35]), .Z(n1460));
Q_MX02 U4030 ( .S(n401), .A0(n1461), .A1(stitcher_out[26]), .Z(nxt_guid3[34]));
Q_AN02 U4031 ( .A0(n161), .A1(guid3[34]), .Z(n1461));
Q_MX02 U4032 ( .S(n401), .A0(n1462), .A1(stitcher_out[25]), .Z(nxt_guid3[33]));
Q_AN02 U4033 ( .A0(n161), .A1(guid3[33]), .Z(n1462));
Q_MX02 U4034 ( .S(n401), .A0(n1463), .A1(stitcher_out[24]), .Z(nxt_guid3[32]));
Q_AN02 U4035 ( .A0(n161), .A1(guid3[32]), .Z(n1463));
Q_MX02 U4036 ( .S(n401), .A0(n1464), .A1(stitcher_out[39]), .Z(nxt_guid3[31]));
Q_AN02 U4037 ( .A0(n161), .A1(guid3[31]), .Z(n1464));
Q_MX02 U4038 ( .S(n401), .A0(n1465), .A1(stitcher_out[38]), .Z(nxt_guid3[30]));
Q_AN02 U4039 ( .A0(n161), .A1(guid3[30]), .Z(n1465));
Q_MX02 U4040 ( .S(n401), .A0(n1466), .A1(stitcher_out[37]), .Z(nxt_guid3[29]));
Q_AN02 U4041 ( .A0(n161), .A1(guid3[29]), .Z(n1466));
Q_MX02 U4042 ( .S(n401), .A0(n1467), .A1(stitcher_out[36]), .Z(nxt_guid3[28]));
Q_AN02 U4043 ( .A0(n161), .A1(guid3[28]), .Z(n1467));
Q_MX02 U4044 ( .S(n401), .A0(n1468), .A1(stitcher_out[35]), .Z(nxt_guid3[27]));
Q_AN02 U4045 ( .A0(n161), .A1(guid3[27]), .Z(n1468));
Q_MX02 U4046 ( .S(n401), .A0(n1469), .A1(stitcher_out[34]), .Z(nxt_guid3[26]));
Q_AN02 U4047 ( .A0(n161), .A1(guid3[26]), .Z(n1469));
Q_MX02 U4048 ( .S(n401), .A0(n1470), .A1(stitcher_out[33]), .Z(nxt_guid3[25]));
Q_AN02 U4049 ( .A0(n161), .A1(guid3[25]), .Z(n1470));
Q_MX02 U4050 ( .S(n401), .A0(n1471), .A1(stitcher_out[32]), .Z(nxt_guid3[24]));
Q_AN02 U4051 ( .A0(n161), .A1(guid3[24]), .Z(n1471));
Q_MX02 U4052 ( .S(n401), .A0(n1472), .A1(stitcher_out[47]), .Z(nxt_guid3[23]));
Q_AN02 U4053 ( .A0(n161), .A1(guid3[23]), .Z(n1472));
Q_MX02 U4054 ( .S(n401), .A0(n1473), .A1(stitcher_out[46]), .Z(nxt_guid3[22]));
Q_AN02 U4055 ( .A0(n161), .A1(guid3[22]), .Z(n1473));
Q_MX02 U4056 ( .S(n401), .A0(n1474), .A1(stitcher_out[45]), .Z(nxt_guid3[21]));
Q_AN02 U4057 ( .A0(n161), .A1(guid3[21]), .Z(n1474));
Q_MX02 U4058 ( .S(n401), .A0(n1475), .A1(stitcher_out[44]), .Z(nxt_guid3[20]));
Q_AN02 U4059 ( .A0(n161), .A1(guid3[20]), .Z(n1475));
Q_MX02 U4060 ( .S(n401), .A0(n1476), .A1(stitcher_out[43]), .Z(nxt_guid3[19]));
Q_AN02 U4061 ( .A0(n161), .A1(guid3[19]), .Z(n1476));
Q_MX02 U4062 ( .S(n401), .A0(n1477), .A1(stitcher_out[42]), .Z(nxt_guid3[18]));
Q_AN02 U4063 ( .A0(n161), .A1(guid3[18]), .Z(n1477));
Q_MX02 U4064 ( .S(n401), .A0(n1478), .A1(stitcher_out[41]), .Z(nxt_guid3[17]));
Q_AN02 U4065 ( .A0(n161), .A1(guid3[17]), .Z(n1478));
Q_MX02 U4066 ( .S(n401), .A0(n1479), .A1(stitcher_out[40]), .Z(nxt_guid3[16]));
Q_AN02 U4067 ( .A0(n161), .A1(guid3[16]), .Z(n1479));
Q_MX02 U4068 ( .S(n401), .A0(n1480), .A1(stitcher_out[55]), .Z(nxt_guid3[15]));
Q_AN02 U4069 ( .A0(n161), .A1(guid3[15]), .Z(n1480));
Q_MX02 U4070 ( .S(n401), .A0(n1481), .A1(stitcher_out[54]), .Z(nxt_guid3[14]));
Q_AN02 U4071 ( .A0(n161), .A1(guid3[14]), .Z(n1481));
Q_MX02 U4072 ( .S(n401), .A0(n1482), .A1(stitcher_out[53]), .Z(nxt_guid3[13]));
Q_AN02 U4073 ( .A0(n161), .A1(guid3[13]), .Z(n1482));
Q_MX02 U4074 ( .S(n401), .A0(n1483), .A1(stitcher_out[52]), .Z(nxt_guid3[12]));
Q_AN02 U4075 ( .A0(n161), .A1(guid3[12]), .Z(n1483));
Q_MX02 U4076 ( .S(n401), .A0(n1484), .A1(stitcher_out[51]), .Z(nxt_guid3[11]));
Q_AN02 U4077 ( .A0(n161), .A1(guid3[11]), .Z(n1484));
Q_MX02 U4078 ( .S(n401), .A0(n1485), .A1(stitcher_out[50]), .Z(nxt_guid3[10]));
Q_AN02 U4079 ( .A0(n161), .A1(guid3[10]), .Z(n1485));
Q_MX02 U4080 ( .S(n401), .A0(n1486), .A1(stitcher_out[49]), .Z(nxt_guid3[9]));
Q_AN02 U4081 ( .A0(n161), .A1(guid3[9]), .Z(n1486));
Q_MX02 U4082 ( .S(n401), .A0(n1487), .A1(stitcher_out[48]), .Z(nxt_guid3[8]));
Q_AN02 U4083 ( .A0(n161), .A1(guid3[8]), .Z(n1487));
Q_MX02 U4084 ( .S(n401), .A0(n1488), .A1(stitcher_out[63]), .Z(nxt_guid3[7]));
Q_AN02 U4085 ( .A0(n161), .A1(guid3[7]), .Z(n1488));
Q_MX02 U4086 ( .S(n401), .A0(n1489), .A1(stitcher_out[62]), .Z(nxt_guid3[6]));
Q_AN02 U4087 ( .A0(n161), .A1(guid3[6]), .Z(n1489));
Q_MX02 U4088 ( .S(n401), .A0(n1490), .A1(stitcher_out[61]), .Z(nxt_guid3[5]));
Q_AN02 U4089 ( .A0(n161), .A1(guid3[5]), .Z(n1490));
Q_MX02 U4090 ( .S(n401), .A0(n1491), .A1(stitcher_out[60]), .Z(nxt_guid3[4]));
Q_AN02 U4091 ( .A0(n161), .A1(guid3[4]), .Z(n1491));
Q_MX02 U4092 ( .S(n401), .A0(n1492), .A1(stitcher_out[59]), .Z(nxt_guid3[3]));
Q_AN02 U4093 ( .A0(n161), .A1(guid3[3]), .Z(n1492));
Q_MX02 U4094 ( .S(n401), .A0(n1493), .A1(stitcher_out[58]), .Z(nxt_guid3[2]));
Q_AN02 U4095 ( .A0(n161), .A1(guid3[2]), .Z(n1493));
Q_MX02 U4096 ( .S(n401), .A0(n1494), .A1(stitcher_out[57]), .Z(nxt_guid3[1]));
Q_AN02 U4097 ( .A0(n161), .A1(guid3[1]), .Z(n1494));
Q_MX02 U4098 ( .S(n401), .A0(n1495), .A1(stitcher_out[56]), .Z(nxt_guid3[0]));
Q_AN02 U4099 ( .A0(n161), .A1(guid3[0]), .Z(n1495));
Q_MX02 U4100 ( .S(n413), .A0(n1496), .A1(stitcher_out[63]), .Z(nxt_iv0[63]));
Q_AN02 U4101 ( .A0(n162), .A1(iv0[63]), .Z(n1496));
Q_MX02 U4102 ( .S(n413), .A0(n1497), .A1(stitcher_out[62]), .Z(nxt_iv0[62]));
Q_AN02 U4103 ( .A0(n162), .A1(iv0[62]), .Z(n1497));
Q_MX02 U4104 ( .S(n413), .A0(n1498), .A1(stitcher_out[61]), .Z(nxt_iv0[61]));
Q_AN02 U4105 ( .A0(n162), .A1(iv0[61]), .Z(n1498));
Q_MX02 U4106 ( .S(n413), .A0(n1499), .A1(stitcher_out[60]), .Z(nxt_iv0[60]));
Q_AN02 U4107 ( .A0(n162), .A1(iv0[60]), .Z(n1499));
Q_MX02 U4108 ( .S(n413), .A0(n1500), .A1(stitcher_out[59]), .Z(nxt_iv0[59]));
Q_AN02 U4109 ( .A0(n162), .A1(iv0[59]), .Z(n1500));
Q_MX02 U4110 ( .S(n413), .A0(n1501), .A1(stitcher_out[58]), .Z(nxt_iv0[58]));
Q_AN02 U4111 ( .A0(n162), .A1(iv0[58]), .Z(n1501));
Q_MX02 U4112 ( .S(n413), .A0(n1502), .A1(stitcher_out[57]), .Z(nxt_iv0[57]));
Q_AN02 U4113 ( .A0(n162), .A1(iv0[57]), .Z(n1502));
Q_MX02 U4114 ( .S(n413), .A0(n1503), .A1(stitcher_out[56]), .Z(nxt_iv0[56]));
Q_AN02 U4115 ( .A0(n162), .A1(iv0[56]), .Z(n1503));
Q_MX02 U4116 ( .S(n413), .A0(n1504), .A1(stitcher_out[55]), .Z(nxt_iv0[55]));
Q_AN02 U4117 ( .A0(n162), .A1(iv0[55]), .Z(n1504));
Q_MX02 U4118 ( .S(n413), .A0(n1505), .A1(stitcher_out[54]), .Z(nxt_iv0[54]));
Q_AN02 U4119 ( .A0(n162), .A1(iv0[54]), .Z(n1505));
Q_MX02 U4120 ( .S(n413), .A0(n1506), .A1(stitcher_out[53]), .Z(nxt_iv0[53]));
Q_AN02 U4121 ( .A0(n162), .A1(iv0[53]), .Z(n1506));
Q_MX02 U4122 ( .S(n413), .A0(n1507), .A1(stitcher_out[52]), .Z(nxt_iv0[52]));
Q_AN02 U4123 ( .A0(n162), .A1(iv0[52]), .Z(n1507));
Q_MX02 U4124 ( .S(n413), .A0(n1508), .A1(stitcher_out[51]), .Z(nxt_iv0[51]));
Q_AN02 U4125 ( .A0(n162), .A1(iv0[51]), .Z(n1508));
Q_MX02 U4126 ( .S(n413), .A0(n1509), .A1(stitcher_out[50]), .Z(nxt_iv0[50]));
Q_AN02 U4127 ( .A0(n162), .A1(iv0[50]), .Z(n1509));
Q_MX02 U4128 ( .S(n413), .A0(n1510), .A1(stitcher_out[49]), .Z(nxt_iv0[49]));
Q_AN02 U4129 ( .A0(n162), .A1(iv0[49]), .Z(n1510));
Q_MX02 U4130 ( .S(n413), .A0(n1511), .A1(stitcher_out[48]), .Z(nxt_iv0[48]));
Q_AN02 U4131 ( .A0(n162), .A1(iv0[48]), .Z(n1511));
Q_MX02 U4132 ( .S(n413), .A0(n1512), .A1(stitcher_out[47]), .Z(nxt_iv0[47]));
Q_AN02 U4133 ( .A0(n162), .A1(iv0[47]), .Z(n1512));
Q_MX02 U4134 ( .S(n413), .A0(n1513), .A1(stitcher_out[46]), .Z(nxt_iv0[46]));
Q_AN02 U4135 ( .A0(n162), .A1(iv0[46]), .Z(n1513));
Q_MX02 U4136 ( .S(n413), .A0(n1514), .A1(stitcher_out[45]), .Z(nxt_iv0[45]));
Q_AN02 U4137 ( .A0(n162), .A1(iv0[45]), .Z(n1514));
Q_MX02 U4138 ( .S(n413), .A0(n1515), .A1(stitcher_out[44]), .Z(nxt_iv0[44]));
Q_AN02 U4139 ( .A0(n162), .A1(iv0[44]), .Z(n1515));
Q_MX02 U4140 ( .S(n413), .A0(n1516), .A1(stitcher_out[43]), .Z(nxt_iv0[43]));
Q_AN02 U4141 ( .A0(n162), .A1(iv0[43]), .Z(n1516));
Q_MX02 U4142 ( .S(n413), .A0(n1517), .A1(stitcher_out[42]), .Z(nxt_iv0[42]));
Q_AN02 U4143 ( .A0(n162), .A1(iv0[42]), .Z(n1517));
Q_MX02 U4144 ( .S(n413), .A0(n1518), .A1(stitcher_out[41]), .Z(nxt_iv0[41]));
Q_AN02 U4145 ( .A0(n162), .A1(iv0[41]), .Z(n1518));
Q_MX02 U4146 ( .S(n413), .A0(n1519), .A1(stitcher_out[40]), .Z(nxt_iv0[40]));
Q_AN02 U4147 ( .A0(n162), .A1(iv0[40]), .Z(n1519));
Q_MX02 U4148 ( .S(n413), .A0(n1520), .A1(stitcher_out[39]), .Z(nxt_iv0[39]));
Q_AN02 U4149 ( .A0(n162), .A1(iv0[39]), .Z(n1520));
Q_MX02 U4150 ( .S(n413), .A0(n1521), .A1(stitcher_out[38]), .Z(nxt_iv0[38]));
Q_AN02 U4151 ( .A0(n162), .A1(iv0[38]), .Z(n1521));
Q_MX02 U4152 ( .S(n413), .A0(n1522), .A1(stitcher_out[37]), .Z(nxt_iv0[37]));
Q_AN02 U4153 ( .A0(n162), .A1(iv0[37]), .Z(n1522));
Q_MX02 U4154 ( .S(n413), .A0(n1523), .A1(stitcher_out[36]), .Z(nxt_iv0[36]));
Q_AN02 U4155 ( .A0(n162), .A1(iv0[36]), .Z(n1523));
Q_MX02 U4156 ( .S(n413), .A0(n1524), .A1(stitcher_out[35]), .Z(nxt_iv0[35]));
Q_AN02 U4157 ( .A0(n162), .A1(iv0[35]), .Z(n1524));
Q_MX02 U4158 ( .S(n413), .A0(n1525), .A1(stitcher_out[34]), .Z(nxt_iv0[34]));
Q_AN02 U4159 ( .A0(n162), .A1(iv0[34]), .Z(n1525));
Q_MX02 U4160 ( .S(n413), .A0(n1526), .A1(stitcher_out[33]), .Z(nxt_iv0[33]));
Q_AN02 U4161 ( .A0(n162), .A1(iv0[33]), .Z(n1526));
Q_MX02 U4162 ( .S(n413), .A0(n1527), .A1(stitcher_out[32]), .Z(nxt_iv0[32]));
Q_AN02 U4163 ( .A0(n162), .A1(iv0[32]), .Z(n1527));
Q_MX02 U4164 ( .S(n413), .A0(n1528), .A1(stitcher_out[31]), .Z(nxt_iv0[31]));
Q_AN02 U4165 ( .A0(n162), .A1(iv0[31]), .Z(n1528));
Q_MX02 U4166 ( .S(n413), .A0(n1529), .A1(stitcher_out[30]), .Z(nxt_iv0[30]));
Q_AN02 U4167 ( .A0(n162), .A1(iv0[30]), .Z(n1529));
Q_MX02 U4168 ( .S(n413), .A0(n1530), .A1(stitcher_out[29]), .Z(nxt_iv0[29]));
Q_AN02 U4169 ( .A0(n162), .A1(iv0[29]), .Z(n1530));
Q_MX02 U4170 ( .S(n413), .A0(n1531), .A1(stitcher_out[28]), .Z(nxt_iv0[28]));
Q_AN02 U4171 ( .A0(n162), .A1(iv0[28]), .Z(n1531));
Q_MX02 U4172 ( .S(n413), .A0(n1532), .A1(stitcher_out[27]), .Z(nxt_iv0[27]));
Q_AN02 U4173 ( .A0(n162), .A1(iv0[27]), .Z(n1532));
Q_MX02 U4174 ( .S(n413), .A0(n1533), .A1(stitcher_out[26]), .Z(nxt_iv0[26]));
Q_AN02 U4175 ( .A0(n162), .A1(iv0[26]), .Z(n1533));
Q_MX02 U4176 ( .S(n413), .A0(n1534), .A1(stitcher_out[25]), .Z(nxt_iv0[25]));
Q_AN02 U4177 ( .A0(n162), .A1(iv0[25]), .Z(n1534));
Q_MX02 U4178 ( .S(n413), .A0(n1535), .A1(stitcher_out[24]), .Z(nxt_iv0[24]));
Q_AN02 U4179 ( .A0(n162), .A1(iv0[24]), .Z(n1535));
Q_MX02 U4180 ( .S(n413), .A0(n1536), .A1(stitcher_out[23]), .Z(nxt_iv0[23]));
Q_AN02 U4181 ( .A0(n162), .A1(iv0[23]), .Z(n1536));
Q_MX02 U4182 ( .S(n413), .A0(n1537), .A1(stitcher_out[22]), .Z(nxt_iv0[22]));
Q_AN02 U4183 ( .A0(n162), .A1(iv0[22]), .Z(n1537));
Q_MX02 U4184 ( .S(n413), .A0(n1538), .A1(stitcher_out[21]), .Z(nxt_iv0[21]));
Q_AN02 U4185 ( .A0(n162), .A1(iv0[21]), .Z(n1538));
Q_MX02 U4186 ( .S(n413), .A0(n1539), .A1(stitcher_out[20]), .Z(nxt_iv0[20]));
Q_AN02 U4187 ( .A0(n162), .A1(iv0[20]), .Z(n1539));
Q_MX02 U4188 ( .S(n413), .A0(n1540), .A1(stitcher_out[19]), .Z(nxt_iv0[19]));
Q_AN02 U4189 ( .A0(n162), .A1(iv0[19]), .Z(n1540));
Q_MX02 U4190 ( .S(n413), .A0(n1541), .A1(stitcher_out[18]), .Z(nxt_iv0[18]));
Q_AN02 U4191 ( .A0(n162), .A1(iv0[18]), .Z(n1541));
Q_MX02 U4192 ( .S(n413), .A0(n1542), .A1(stitcher_out[17]), .Z(nxt_iv0[17]));
Q_AN02 U4193 ( .A0(n162), .A1(iv0[17]), .Z(n1542));
Q_MX02 U4194 ( .S(n413), .A0(n1543), .A1(stitcher_out[16]), .Z(nxt_iv0[16]));
Q_AN02 U4195 ( .A0(n162), .A1(iv0[16]), .Z(n1543));
Q_MX02 U4196 ( .S(n413), .A0(n1544), .A1(stitcher_out[15]), .Z(nxt_iv0[15]));
Q_AN02 U4197 ( .A0(n162), .A1(iv0[15]), .Z(n1544));
Q_MX02 U4198 ( .S(n413), .A0(n1545), .A1(stitcher_out[14]), .Z(nxt_iv0[14]));
Q_AN02 U4199 ( .A0(n162), .A1(iv0[14]), .Z(n1545));
Q_MX02 U4200 ( .S(n413), .A0(n1546), .A1(stitcher_out[13]), .Z(nxt_iv0[13]));
Q_AN02 U4201 ( .A0(n162), .A1(iv0[13]), .Z(n1546));
Q_MX02 U4202 ( .S(n413), .A0(n1547), .A1(stitcher_out[12]), .Z(nxt_iv0[12]));
Q_AN02 U4203 ( .A0(n162), .A1(iv0[12]), .Z(n1547));
Q_MX02 U4204 ( .S(n413), .A0(n1548), .A1(stitcher_out[11]), .Z(nxt_iv0[11]));
Q_AN02 U4205 ( .A0(n162), .A1(iv0[11]), .Z(n1548));
Q_MX02 U4206 ( .S(n413), .A0(n1549), .A1(stitcher_out[10]), .Z(nxt_iv0[10]));
Q_AN02 U4207 ( .A0(n162), .A1(iv0[10]), .Z(n1549));
Q_MX02 U4208 ( .S(n413), .A0(n1550), .A1(stitcher_out[9]), .Z(nxt_iv0[9]));
Q_AN02 U4209 ( .A0(n162), .A1(iv0[9]), .Z(n1550));
Q_MX02 U4210 ( .S(n413), .A0(n1551), .A1(stitcher_out[8]), .Z(nxt_iv0[8]));
Q_AN02 U4211 ( .A0(n162), .A1(iv0[8]), .Z(n1551));
Q_MX02 U4212 ( .S(n413), .A0(n1552), .A1(stitcher_out[7]), .Z(nxt_iv0[7]));
Q_AN02 U4213 ( .A0(n162), .A1(iv0[7]), .Z(n1552));
Q_MX02 U4214 ( .S(n413), .A0(n1553), .A1(stitcher_out[6]), .Z(nxt_iv0[6]));
Q_AN02 U4215 ( .A0(n162), .A1(iv0[6]), .Z(n1553));
Q_MX02 U4216 ( .S(n413), .A0(n1554), .A1(stitcher_out[5]), .Z(nxt_iv0[5]));
Q_AN02 U4217 ( .A0(n162), .A1(iv0[5]), .Z(n1554));
Q_MX02 U4218 ( .S(n413), .A0(n1555), .A1(stitcher_out[4]), .Z(nxt_iv0[4]));
Q_AN02 U4219 ( .A0(n162), .A1(iv0[4]), .Z(n1555));
Q_MX02 U4220 ( .S(n413), .A0(n1556), .A1(stitcher_out[3]), .Z(nxt_iv0[3]));
Q_AN02 U4221 ( .A0(n162), .A1(iv0[3]), .Z(n1556));
Q_MX02 U4222 ( .S(n413), .A0(n1557), .A1(stitcher_out[2]), .Z(nxt_iv0[2]));
Q_AN02 U4223 ( .A0(n162), .A1(iv0[2]), .Z(n1557));
Q_MX02 U4224 ( .S(n413), .A0(n1558), .A1(stitcher_out[1]), .Z(nxt_iv0[1]));
Q_AN02 U4225 ( .A0(n162), .A1(iv0[1]), .Z(n1558));
Q_MX02 U4226 ( .S(n413), .A0(n1559), .A1(stitcher_out[0]), .Z(nxt_iv0[0]));
Q_AN02 U4227 ( .A0(n162), .A1(iv0[0]), .Z(n1559));
Q_MX02 U4228 ( .S(n421), .A0(n1560), .A1(stitcher_out[63]), .Z(nxt_iv1[63]));
Q_AN02 U4229 ( .A0(n163), .A1(iv1[63]), .Z(n1560));
Q_MX02 U4230 ( .S(n421), .A0(n1561), .A1(stitcher_out[62]), .Z(nxt_iv1[62]));
Q_AN02 U4231 ( .A0(n163), .A1(iv1[62]), .Z(n1561));
Q_MX02 U4232 ( .S(n421), .A0(n1562), .A1(stitcher_out[61]), .Z(nxt_iv1[61]));
Q_AN02 U4233 ( .A0(n163), .A1(iv1[61]), .Z(n1562));
Q_MX02 U4234 ( .S(n421), .A0(n1563), .A1(stitcher_out[60]), .Z(nxt_iv1[60]));
Q_AN02 U4235 ( .A0(n163), .A1(iv1[60]), .Z(n1563));
Q_MX02 U4236 ( .S(n421), .A0(n1564), .A1(stitcher_out[59]), .Z(nxt_iv1[59]));
Q_AN02 U4237 ( .A0(n163), .A1(iv1[59]), .Z(n1564));
Q_MX02 U4238 ( .S(n421), .A0(n1565), .A1(stitcher_out[58]), .Z(nxt_iv1[58]));
Q_AN02 U4239 ( .A0(n163), .A1(iv1[58]), .Z(n1565));
Q_MX02 U4240 ( .S(n421), .A0(n1566), .A1(stitcher_out[57]), .Z(nxt_iv1[57]));
Q_AN02 U4241 ( .A0(n163), .A1(iv1[57]), .Z(n1566));
Q_MX02 U4242 ( .S(n421), .A0(n1567), .A1(stitcher_out[56]), .Z(nxt_iv1[56]));
Q_AN02 U4243 ( .A0(n163), .A1(iv1[56]), .Z(n1567));
Q_MX02 U4244 ( .S(n421), .A0(n1568), .A1(stitcher_out[55]), .Z(nxt_iv1[55]));
Q_AN02 U4245 ( .A0(n163), .A1(iv1[55]), .Z(n1568));
Q_MX02 U4246 ( .S(n421), .A0(n1569), .A1(stitcher_out[54]), .Z(nxt_iv1[54]));
Q_AN02 U4247 ( .A0(n163), .A1(iv1[54]), .Z(n1569));
Q_MX02 U4248 ( .S(n421), .A0(n1570), .A1(stitcher_out[53]), .Z(nxt_iv1[53]));
Q_AN02 U4249 ( .A0(n163), .A1(iv1[53]), .Z(n1570));
Q_MX02 U4250 ( .S(n421), .A0(n1571), .A1(stitcher_out[52]), .Z(nxt_iv1[52]));
Q_AN02 U4251 ( .A0(n163), .A1(iv1[52]), .Z(n1571));
Q_MX02 U4252 ( .S(n421), .A0(n1572), .A1(stitcher_out[51]), .Z(nxt_iv1[51]));
Q_AN02 U4253 ( .A0(n163), .A1(iv1[51]), .Z(n1572));
Q_MX02 U4254 ( .S(n421), .A0(n1573), .A1(stitcher_out[50]), .Z(nxt_iv1[50]));
Q_AN02 U4255 ( .A0(n163), .A1(iv1[50]), .Z(n1573));
Q_MX02 U4256 ( .S(n421), .A0(n1574), .A1(stitcher_out[49]), .Z(nxt_iv1[49]));
Q_AN02 U4257 ( .A0(n163), .A1(iv1[49]), .Z(n1574));
Q_MX02 U4258 ( .S(n421), .A0(n1575), .A1(stitcher_out[48]), .Z(nxt_iv1[48]));
Q_AN02 U4259 ( .A0(n163), .A1(iv1[48]), .Z(n1575));
Q_MX02 U4260 ( .S(n421), .A0(n1576), .A1(stitcher_out[47]), .Z(nxt_iv1[47]));
Q_AN02 U4261 ( .A0(n163), .A1(iv1[47]), .Z(n1576));
Q_MX02 U4262 ( .S(n421), .A0(n1577), .A1(stitcher_out[46]), .Z(nxt_iv1[46]));
Q_AN02 U4263 ( .A0(n163), .A1(iv1[46]), .Z(n1577));
Q_MX02 U4264 ( .S(n421), .A0(n1578), .A1(stitcher_out[45]), .Z(nxt_iv1[45]));
Q_AN02 U4265 ( .A0(n163), .A1(iv1[45]), .Z(n1578));
Q_MX02 U4266 ( .S(n421), .A0(n1579), .A1(stitcher_out[44]), .Z(nxt_iv1[44]));
Q_AN02 U4267 ( .A0(n163), .A1(iv1[44]), .Z(n1579));
Q_MX02 U4268 ( .S(n421), .A0(n1580), .A1(stitcher_out[43]), .Z(nxt_iv1[43]));
Q_AN02 U4269 ( .A0(n163), .A1(iv1[43]), .Z(n1580));
Q_MX02 U4270 ( .S(n421), .A0(n1581), .A1(stitcher_out[42]), .Z(nxt_iv1[42]));
Q_AN02 U4271 ( .A0(n163), .A1(iv1[42]), .Z(n1581));
Q_MX02 U4272 ( .S(n421), .A0(n1582), .A1(stitcher_out[41]), .Z(nxt_iv1[41]));
Q_AN02 U4273 ( .A0(n163), .A1(iv1[41]), .Z(n1582));
Q_MX02 U4274 ( .S(n421), .A0(n1583), .A1(stitcher_out[40]), .Z(nxt_iv1[40]));
Q_AN02 U4275 ( .A0(n163), .A1(iv1[40]), .Z(n1583));
Q_MX02 U4276 ( .S(n421), .A0(n1584), .A1(stitcher_out[39]), .Z(nxt_iv1[39]));
Q_AN02 U4277 ( .A0(n163), .A1(iv1[39]), .Z(n1584));
Q_MX02 U4278 ( .S(n421), .A0(n1585), .A1(stitcher_out[38]), .Z(nxt_iv1[38]));
Q_AN02 U4279 ( .A0(n163), .A1(iv1[38]), .Z(n1585));
Q_MX02 U4280 ( .S(n421), .A0(n1586), .A1(stitcher_out[37]), .Z(nxt_iv1[37]));
Q_AN02 U4281 ( .A0(n163), .A1(iv1[37]), .Z(n1586));
Q_MX02 U4282 ( .S(n421), .A0(n1587), .A1(stitcher_out[36]), .Z(nxt_iv1[36]));
Q_AN02 U4283 ( .A0(n163), .A1(iv1[36]), .Z(n1587));
Q_MX02 U4284 ( .S(n421), .A0(n1588), .A1(stitcher_out[35]), .Z(nxt_iv1[35]));
Q_AN02 U4285 ( .A0(n163), .A1(iv1[35]), .Z(n1588));
Q_MX02 U4286 ( .S(n421), .A0(n1589), .A1(stitcher_out[34]), .Z(nxt_iv1[34]));
Q_AN02 U4287 ( .A0(n163), .A1(iv1[34]), .Z(n1589));
Q_MX02 U4288 ( .S(n421), .A0(n1590), .A1(stitcher_out[33]), .Z(nxt_iv1[33]));
Q_AN02 U4289 ( .A0(n163), .A1(iv1[33]), .Z(n1590));
Q_MX02 U4290 ( .S(n421), .A0(n1591), .A1(stitcher_out[32]), .Z(nxt_iv1[32]));
Q_AN02 U4291 ( .A0(n163), .A1(iv1[32]), .Z(n1591));
Q_MX02 U4292 ( .S(n421), .A0(n1592), .A1(stitcher_out[31]), .Z(nxt_iv1[31]));
Q_AN02 U4293 ( .A0(n163), .A1(iv1[31]), .Z(n1592));
Q_MX02 U4294 ( .S(n421), .A0(n1593), .A1(stitcher_out[30]), .Z(nxt_iv1[30]));
Q_AN02 U4295 ( .A0(n163), .A1(iv1[30]), .Z(n1593));
Q_MX02 U4296 ( .S(n421), .A0(n1594), .A1(stitcher_out[29]), .Z(nxt_iv1[29]));
Q_AN02 U4297 ( .A0(n163), .A1(iv1[29]), .Z(n1594));
Q_MX02 U4298 ( .S(n421), .A0(n1595), .A1(stitcher_out[28]), .Z(nxt_iv1[28]));
Q_AN02 U4299 ( .A0(n163), .A1(iv1[28]), .Z(n1595));
Q_MX02 U4300 ( .S(n421), .A0(n1596), .A1(stitcher_out[27]), .Z(nxt_iv1[27]));
Q_AN02 U4301 ( .A0(n163), .A1(iv1[27]), .Z(n1596));
Q_MX02 U4302 ( .S(n421), .A0(n1597), .A1(stitcher_out[26]), .Z(nxt_iv1[26]));
Q_AN02 U4303 ( .A0(n163), .A1(iv1[26]), .Z(n1597));
Q_MX02 U4304 ( .S(n421), .A0(n1598), .A1(stitcher_out[25]), .Z(nxt_iv1[25]));
Q_AN02 U4305 ( .A0(n163), .A1(iv1[25]), .Z(n1598));
Q_MX02 U4306 ( .S(n421), .A0(n1599), .A1(stitcher_out[24]), .Z(nxt_iv1[24]));
Q_AN02 U4307 ( .A0(n163), .A1(iv1[24]), .Z(n1599));
Q_MX02 U4308 ( .S(n421), .A0(n1600), .A1(stitcher_out[23]), .Z(nxt_iv1[23]));
Q_AN02 U4309 ( .A0(n163), .A1(iv1[23]), .Z(n1600));
Q_MX02 U4310 ( .S(n421), .A0(n1601), .A1(stitcher_out[22]), .Z(nxt_iv1[22]));
Q_AN02 U4311 ( .A0(n163), .A1(iv1[22]), .Z(n1601));
Q_MX02 U4312 ( .S(n421), .A0(n1602), .A1(stitcher_out[21]), .Z(nxt_iv1[21]));
Q_AN02 U4313 ( .A0(n163), .A1(iv1[21]), .Z(n1602));
Q_MX02 U4314 ( .S(n421), .A0(n1603), .A1(stitcher_out[20]), .Z(nxt_iv1[20]));
Q_AN02 U4315 ( .A0(n163), .A1(iv1[20]), .Z(n1603));
Q_MX02 U4316 ( .S(n421), .A0(n1604), .A1(stitcher_out[19]), .Z(nxt_iv1[19]));
Q_AN02 U4317 ( .A0(n163), .A1(iv1[19]), .Z(n1604));
Q_MX02 U4318 ( .S(n421), .A0(n1605), .A1(stitcher_out[18]), .Z(nxt_iv1[18]));
Q_AN02 U4319 ( .A0(n163), .A1(iv1[18]), .Z(n1605));
Q_MX02 U4320 ( .S(n421), .A0(n1606), .A1(stitcher_out[17]), .Z(nxt_iv1[17]));
Q_AN02 U4321 ( .A0(n163), .A1(iv1[17]), .Z(n1606));
Q_MX02 U4322 ( .S(n421), .A0(n1607), .A1(stitcher_out[16]), .Z(nxt_iv1[16]));
Q_AN02 U4323 ( .A0(n163), .A1(iv1[16]), .Z(n1607));
Q_MX02 U4324 ( .S(n421), .A0(n1608), .A1(stitcher_out[15]), .Z(nxt_iv1[15]));
Q_AN02 U4325 ( .A0(n163), .A1(iv1[15]), .Z(n1608));
Q_MX02 U4326 ( .S(n421), .A0(n1609), .A1(stitcher_out[14]), .Z(nxt_iv1[14]));
Q_AN02 U4327 ( .A0(n163), .A1(iv1[14]), .Z(n1609));
Q_MX02 U4328 ( .S(n421), .A0(n1610), .A1(stitcher_out[13]), .Z(nxt_iv1[13]));
Q_AN02 U4329 ( .A0(n163), .A1(iv1[13]), .Z(n1610));
Q_MX02 U4330 ( .S(n421), .A0(n1611), .A1(stitcher_out[12]), .Z(nxt_iv1[12]));
Q_AN02 U4331 ( .A0(n163), .A1(iv1[12]), .Z(n1611));
Q_MX02 U4332 ( .S(n421), .A0(n1612), .A1(stitcher_out[11]), .Z(nxt_iv1[11]));
Q_AN02 U4333 ( .A0(n163), .A1(iv1[11]), .Z(n1612));
Q_MX02 U4334 ( .S(n421), .A0(n1613), .A1(stitcher_out[10]), .Z(nxt_iv1[10]));
Q_AN02 U4335 ( .A0(n163), .A1(iv1[10]), .Z(n1613));
Q_MX02 U4336 ( .S(n421), .A0(n1614), .A1(stitcher_out[9]), .Z(nxt_iv1[9]));
Q_AN02 U4337 ( .A0(n163), .A1(iv1[9]), .Z(n1614));
Q_MX02 U4338 ( .S(n421), .A0(n1615), .A1(stitcher_out[8]), .Z(nxt_iv1[8]));
Q_AN02 U4339 ( .A0(n163), .A1(iv1[8]), .Z(n1615));
Q_MX02 U4340 ( .S(n421), .A0(n1616), .A1(stitcher_out[7]), .Z(nxt_iv1[7]));
Q_AN02 U4341 ( .A0(n163), .A1(iv1[7]), .Z(n1616));
Q_MX02 U4342 ( .S(n421), .A0(n1617), .A1(stitcher_out[6]), .Z(nxt_iv1[6]));
Q_AN02 U4343 ( .A0(n163), .A1(iv1[6]), .Z(n1617));
Q_MX02 U4344 ( .S(n421), .A0(n1618), .A1(stitcher_out[5]), .Z(nxt_iv1[5]));
Q_AN02 U4345 ( .A0(n163), .A1(iv1[5]), .Z(n1618));
Q_MX02 U4346 ( .S(n421), .A0(n1619), .A1(stitcher_out[4]), .Z(nxt_iv1[4]));
Q_AN02 U4347 ( .A0(n163), .A1(iv1[4]), .Z(n1619));
Q_MX02 U4348 ( .S(n421), .A0(n1620), .A1(stitcher_out[3]), .Z(nxt_iv1[3]));
Q_AN02 U4349 ( .A0(n163), .A1(iv1[3]), .Z(n1620));
Q_MX02 U4350 ( .S(n421), .A0(n1621), .A1(stitcher_out[2]), .Z(nxt_iv1[2]));
Q_AN02 U4351 ( .A0(n163), .A1(iv1[2]), .Z(n1621));
Q_MX02 U4352 ( .S(n421), .A0(n1622), .A1(stitcher_out[1]), .Z(nxt_iv1[1]));
Q_AN02 U4353 ( .A0(n163), .A1(iv1[1]), .Z(n1622));
Q_MX02 U4354 ( .S(n421), .A0(n1623), .A1(stitcher_out[0]), .Z(nxt_iv1[0]));
Q_AN02 U4355 ( .A0(n163), .A1(iv1[0]), .Z(n1623));
Q_MX03 U4356 ( .S0(n164), .S1(n435), .A0(debug_cmd[31]), .A1(buffer[31]), .A2(stitcher_out[63]), .Z(nxt_buffer[31]));
Q_MX03 U4357 ( .S0(n164), .S1(n435), .A0(debug_cmd[30]), .A1(buffer[30]), .A2(stitcher_out[62]), .Z(nxt_buffer[30]));
Q_MX03 U4358 ( .S0(n164), .S1(n435), .A0(debug_cmd[29]), .A1(buffer[29]), .A2(stitcher_out[61]), .Z(nxt_buffer[29]));
Q_MX03 U4359 ( .S0(n164), .S1(n435), .A0(debug_cmd[28]), .A1(buffer[28]), .A2(stitcher_out[60]), .Z(nxt_buffer[28]));
Q_MX03 U4360 ( .S0(n164), .S1(n435), .A0(debug_cmd[27]), .A1(buffer[27]), .A2(stitcher_out[59]), .Z(nxt_buffer[27]));
Q_MX03 U4361 ( .S0(n164), .S1(n435), .A0(debug_cmd[26]), .A1(buffer[26]), .A2(stitcher_out[58]), .Z(nxt_buffer[26]));
Q_MX03 U4362 ( .S0(n164), .S1(n435), .A0(debug_cmd[25]), .A1(buffer[25]), .A2(stitcher_out[57]), .Z(nxt_buffer[25]));
Q_MX03 U4363 ( .S0(n164), .S1(n435), .A0(debug_cmd[24]), .A1(buffer[24]), .A2(stitcher_out[56]), .Z(nxt_buffer[24]));
Q_MX03 U4364 ( .S0(n164), .S1(n435), .A0(debug_cmd[23]), .A1(buffer[23]), .A2(stitcher_out[55]), .Z(nxt_buffer[23]));
Q_MX03 U4365 ( .S0(n164), .S1(n435), .A0(debug_cmd[22]), .A1(buffer[22]), .A2(stitcher_out[54]), .Z(nxt_buffer[22]));
Q_MX03 U4366 ( .S0(n164), .S1(n435), .A0(debug_cmd[21]), .A1(buffer[21]), .A2(stitcher_out[53]), .Z(nxt_buffer[21]));
Q_MX03 U4367 ( .S0(n164), .S1(n435), .A0(debug_cmd[20]), .A1(buffer[20]), .A2(stitcher_out[52]), .Z(nxt_buffer[20]));
Q_MX03 U4368 ( .S0(n164), .S1(n435), .A0(debug_cmd[19]), .A1(buffer[19]), .A2(stitcher_out[51]), .Z(nxt_buffer[19]));
Q_MX03 U4369 ( .S0(n164), .S1(n435), .A0(debug_cmd[18]), .A1(buffer[18]), .A2(stitcher_out[50]), .Z(nxt_buffer[18]));
Q_MX03 U4370 ( .S0(n164), .S1(n435), .A0(debug_cmd[17]), .A1(buffer[17]), .A2(stitcher_out[49]), .Z(nxt_buffer[17]));
Q_MX03 U4371 ( .S0(n164), .S1(n435), .A0(debug_cmd[16]), .A1(buffer[16]), .A2(stitcher_out[48]), .Z(nxt_buffer[16]));
Q_MX03 U4372 ( .S0(n164), .S1(n435), .A0(debug_cmd[15]), .A1(buffer[15]), .A2(stitcher_out[47]), .Z(nxt_buffer[15]));
Q_MX03 U4373 ( .S0(n164), .S1(n435), .A0(debug_cmd[14]), .A1(buffer[14]), .A2(stitcher_out[46]), .Z(nxt_buffer[14]));
Q_MX03 U4374 ( .S0(n164), .S1(n435), .A0(debug_cmd[13]), .A1(buffer[13]), .A2(stitcher_out[45]), .Z(nxt_buffer[13]));
Q_MX03 U4375 ( .S0(n164), .S1(n435), .A0(debug_cmd[12]), .A1(buffer[12]), .A2(stitcher_out[44]), .Z(nxt_buffer[12]));
Q_MX03 U4376 ( .S0(n164), .S1(n435), .A0(debug_cmd[11]), .A1(buffer[11]), .A2(stitcher_out[43]), .Z(nxt_buffer[11]));
Q_MX03 U4377 ( .S0(n164), .S1(n435), .A0(debug_cmd[10]), .A1(buffer[10]), .A2(stitcher_out[42]), .Z(nxt_buffer[10]));
Q_MX03 U4378 ( .S0(n164), .S1(n435), .A0(debug_cmd[9]), .A1(buffer[9]), .A2(stitcher_out[41]), .Z(nxt_buffer[9]));
Q_MX03 U4379 ( .S0(n164), .S1(n435), .A0(debug_cmd[8]), .A1(buffer[8]), .A2(stitcher_out[40]), .Z(nxt_buffer[8]));
Q_MX03 U4380 ( .S0(n164), .S1(n435), .A0(debug_cmd[7]), .A1(buffer[7]), .A2(stitcher_out[39]), .Z(nxt_buffer[7]));
Q_MX03 U4381 ( .S0(n164), .S1(n435), .A0(debug_cmd[6]), .A1(buffer[6]), .A2(stitcher_out[38]), .Z(nxt_buffer[6]));
Q_MX03 U4382 ( .S0(n164), .S1(n435), .A0(debug_cmd[5]), .A1(buffer[5]), .A2(stitcher_out[37]), .Z(nxt_buffer[5]));
Q_MX03 U4383 ( .S0(n164), .S1(n435), .A0(debug_cmd[4]), .A1(buffer[4]), .A2(stitcher_out[36]), .Z(nxt_buffer[4]));
Q_MX03 U4384 ( .S0(n164), .S1(n435), .A0(debug_cmd[3]), .A1(buffer[3]), .A2(stitcher_out[35]), .Z(nxt_buffer[3]));
Q_MX03 U4385 ( .S0(n164), .S1(n435), .A0(debug_cmd[2]), .A1(buffer[2]), .A2(stitcher_out[34]), .Z(nxt_buffer[2]));
Q_MX03 U4386 ( .S0(n164), .S1(n435), .A0(debug_cmd[1]), .A1(buffer[1]), .A2(stitcher_out[33]), .Z(nxt_buffer[1]));
Q_MX03 U4387 ( .S0(n164), .S1(n435), .A0(debug_cmd[0]), .A1(buffer[0]), .A2(stitcher_out[32]), .Z(nxt_buffer[0]));
Q_MX02 U4388 ( .S(n591), .A0(stitcher_out[31]), .A1(n1624), .Z(nxt_aux_key_header[31]));
Q_AN02 U4389 ( .A0(n167), .A1(aux_key_header[31]), .Z(n1624));
Q_MX02 U4390 ( .S(n591), .A0(stitcher_out[30]), .A1(n1625), .Z(nxt_aux_key_header[30]));
Q_AN02 U4391 ( .A0(n167), .A1(aux_key_header[30]), .Z(n1625));
Q_MX02 U4392 ( .S(n591), .A0(stitcher_out[29]), .A1(n1626), .Z(nxt_aux_key_header[29]));
Q_AN02 U4393 ( .A0(n167), .A1(aux_key_header[29]), .Z(n1626));
Q_MX02 U4394 ( .S(n591), .A0(stitcher_out[28]), .A1(n1627), .Z(nxt_aux_key_header[28]));
Q_AN02 U4395 ( .A0(n167), .A1(aux_key_header[28]), .Z(n1627));
Q_MX02 U4396 ( .S(n591), .A0(stitcher_out[27]), .A1(n1628), .Z(nxt_aux_key_header[27]));
Q_AN02 U4397 ( .A0(n167), .A1(aux_key_header[27]), .Z(n1628));
Q_MX02 U4398 ( .S(n591), .A0(stitcher_out[26]), .A1(n1629), .Z(nxt_aux_key_header[26]));
Q_AN02 U4399 ( .A0(n167), .A1(aux_key_header[26]), .Z(n1629));
Q_MX02 U4400 ( .S(n591), .A0(stitcher_out[25]), .A1(n1630), .Z(nxt_aux_key_header[25]));
Q_AN02 U4401 ( .A0(n167), .A1(aux_key_header[25]), .Z(n1630));
Q_MX02 U4402 ( .S(n591), .A0(stitcher_out[24]), .A1(n1631), .Z(nxt_aux_key_header[24]));
Q_AN02 U4403 ( .A0(n167), .A1(aux_key_header[24]), .Z(n1631));
Q_MX02 U4404 ( .S(n591), .A0(stitcher_out[23]), .A1(n1632), .Z(nxt_aux_key_header[23]));
Q_AN02 U4405 ( .A0(n167), .A1(aux_key_header[23]), .Z(n1632));
Q_MX02 U4406 ( .S(n591), .A0(stitcher_out[22]), .A1(n1633), .Z(nxt_aux_key_header[22]));
Q_AN02 U4407 ( .A0(n167), .A1(aux_key_header[22]), .Z(n1633));
Q_MX02 U4408 ( .S(n591), .A0(stitcher_out[21]), .A1(n1634), .Z(nxt_aux_key_header[21]));
Q_AN02 U4409 ( .A0(n167), .A1(aux_key_header[21]), .Z(n1634));
Q_MX02 U4410 ( .S(n591), .A0(stitcher_out[20]), .A1(n1635), .Z(nxt_aux_key_header[20]));
Q_AN02 U4411 ( .A0(n167), .A1(aux_key_header[20]), .Z(n1635));
Q_MX02 U4412 ( .S(n591), .A0(stitcher_out[19]), .A1(n1636), .Z(nxt_aux_key_header[19]));
Q_AN02 U4413 ( .A0(n167), .A1(aux_key_header[19]), .Z(n1636));
Q_MX02 U4414 ( .S(n591), .A0(stitcher_out[18]), .A1(n1637), .Z(nxt_aux_key_header[18]));
Q_AN02 U4415 ( .A0(n167), .A1(aux_key_header[18]), .Z(n1637));
Q_MX02 U4416 ( .S(n591), .A0(stitcher_out[17]), .A1(n1638), .Z(nxt_aux_key_header[17]));
Q_AN02 U4417 ( .A0(n167), .A1(aux_key_header[17]), .Z(n1638));
Q_MX02 U4418 ( .S(n591), .A0(stitcher_out[16]), .A1(n1639), .Z(nxt_aux_key_header[16]));
Q_AN02 U4419 ( .A0(n167), .A1(aux_key_header[16]), .Z(n1639));
Q_MX02 U4420 ( .S(n591), .A0(stitcher_out[15]), .A1(n1640), .Z(nxt_aux_key_header[15]));
Q_AN02 U4421 ( .A0(n167), .A1(aux_key_header[15]), .Z(n1640));
Q_MX02 U4422 ( .S(n591), .A0(stitcher_out[14]), .A1(n1641), .Z(nxt_aux_key_header[14]));
Q_AN02 U4423 ( .A0(n167), .A1(aux_key_header[14]), .Z(n1641));
Q_MX02 U4424 ( .S(n591), .A0(stitcher_out[13]), .A1(n1642), .Z(nxt_aux_key_header[13]));
Q_AN02 U4425 ( .A0(n167), .A1(aux_key_header[13]), .Z(n1642));
Q_MX02 U4426 ( .S(n591), .A0(stitcher_out[12]), .A1(n1643), .Z(nxt_aux_key_header[12]));
Q_AN02 U4427 ( .A0(n167), .A1(aux_key_header[12]), .Z(n1643));
Q_MX02 U4428 ( .S(n591), .A0(stitcher_out[11]), .A1(n1644), .Z(nxt_aux_key_header[11]));
Q_AN02 U4429 ( .A0(n167), .A1(aux_key_header[11]), .Z(n1644));
Q_MX02 U4430 ( .S(n591), .A0(stitcher_out[10]), .A1(n1645), .Z(nxt_aux_key_header[10]));
Q_AN02 U4431 ( .A0(n167), .A1(aux_key_header[10]), .Z(n1645));
Q_MX02 U4432 ( .S(n591), .A0(stitcher_out[9]), .A1(n1646), .Z(nxt_aux_key_header[9]));
Q_AN02 U4433 ( .A0(n167), .A1(aux_key_header[9]), .Z(n1646));
Q_MX02 U4434 ( .S(n591), .A0(stitcher_out[8]), .A1(n1647), .Z(nxt_aux_key_header[8]));
Q_AN02 U4435 ( .A0(n167), .A1(aux_key_header[8]), .Z(n1647));
Q_MX02 U4436 ( .S(n591), .A0(stitcher_out[7]), .A1(n1648), .Z(nxt_aux_key_header[7]));
Q_AN02 U4437 ( .A0(n167), .A1(aux_key_header[7]), .Z(n1648));
Q_MX02 U4438 ( .S(n591), .A0(stitcher_out[6]), .A1(n1649), .Z(nxt_aux_key_header[6]));
Q_AN02 U4439 ( .A0(n167), .A1(aux_key_header[6]), .Z(n1649));
Q_MX02 U4440 ( .S(n591), .A0(stitcher_out[5]), .A1(n1650), .Z(nxt_aux_key_header[5]));
Q_AN02 U4441 ( .A0(n167), .A1(aux_key_header[5]), .Z(n1650));
Q_MX02 U4442 ( .S(n591), .A0(stitcher_out[4]), .A1(n1651), .Z(nxt_aux_key_header[4]));
Q_AN02 U4443 ( .A0(n167), .A1(aux_key_header[4]), .Z(n1651));
Q_MX02 U4444 ( .S(n591), .A0(stitcher_out[3]), .A1(n1652), .Z(nxt_aux_key_header[3]));
Q_AN02 U4445 ( .A0(n167), .A1(aux_key_header[3]), .Z(n1652));
Q_MX02 U4446 ( .S(n591), .A0(stitcher_out[2]), .A1(n1653), .Z(nxt_aux_key_header[2]));
Q_AN02 U4447 ( .A0(n167), .A1(aux_key_header[2]), .Z(n1653));
Q_MX02 U4448 ( .S(n591), .A0(stitcher_out[1]), .A1(n1654), .Z(nxt_aux_key_header[1]));
Q_AN02 U4449 ( .A0(n167), .A1(aux_key_header[1]), .Z(n1654));
Q_MX02 U4450 ( .S(n591), .A0(stitcher_out[0]), .A1(n1655), .Z(nxt_aux_key_header[0]));
Q_AN02 U4451 ( .A0(n167), .A1(aux_key_header[0]), .Z(n1655));
Q_MX02 U4452 ( .S(n170), .A0(stitcher_out[7]), .A1(kme_internal_word0[7]), .Z(nxt_kme_internal_word0[7]));
Q_MX02 U4453 ( .S(n170), .A0(stitcher_out[6]), .A1(kme_internal_word0[6]), .Z(nxt_kme_internal_word0[6]));
Q_MX02 U4454 ( .S(n170), .A0(stitcher_out[5]), .A1(kme_internal_word0[5]), .Z(nxt_kme_internal_word0[5]));
Q_MX02 U4455 ( .S(n170), .A0(stitcher_out[4]), .A1(kme_internal_word0[4]), .Z(nxt_kme_internal_word0[4]));
Q_MX02 U4456 ( .S(n170), .A0(stitcher_out[3]), .A1(kme_internal_word0[3]), .Z(nxt_kme_internal_word0[3]));
Q_MX02 U4457 ( .S(n170), .A0(stitcher_out[2]), .A1(kme_internal_word0[2]), .Z(nxt_kme_internal_word0[2]));
Q_MX02 U4458 ( .S(n170), .A0(stitcher_out[1]), .A1(kme_internal_word0[1]), .Z(nxt_kme_internal_word0[1]));
Q_MX02 U4459 ( .S(n170), .A0(stitcher_out[0]), .A1(kme_internal_word0[0]), .Z(nxt_kme_internal_word0[0]));
Q_AN02 U4460 ( .A0(n170), .A1(kme_internal_word0[15]), .Z(nxt_kme_internal_word0[15]));
Q_AN02 U4461 ( .A0(n170), .A1(kme_internal_word0[14]), .Z(nxt_kme_internal_word0[14]));
Q_AN02 U4462 ( .A0(n170), .A1(kme_internal_word0[13]), .Z(nxt_kme_internal_word0[13]));
Q_AN02 U4463 ( .A0(n170), .A1(kme_internal_word0[12]), .Z(nxt_kme_internal_word0[12]));
Q_AN02 U4464 ( .A0(n170), .A1(kme_internal_word0[11]), .Z(nxt_kme_internal_word0[11]));
Q_AN02 U4465 ( .A0(n170), .A1(kme_internal_word0[10]), .Z(nxt_kme_internal_word0[10]));
Q_AN02 U4466 ( .A0(n170), .A1(kme_internal_word0[9]), .Z(nxt_kme_internal_word0[9]));
Q_AN02 U4467 ( .A0(n170), .A1(kme_internal_word0[8]), .Z(nxt_kme_internal_word0[8]));
Q_MX02 U4468 ( .S(n170), .A0(stitcher_out[23]), .A1(kme_internal_word0[23]), .Z(nxt_kme_internal_word0[23]));
Q_MX02 U4469 ( .S(n170), .A0(stitcher_out[22]), .A1(kme_internal_word0[22]), .Z(nxt_kme_internal_word0[22]));
Q_MX02 U4470 ( .S(n170), .A0(stitcher_out[21]), .A1(kme_internal_word0[21]), .Z(nxt_kme_internal_word0[21]));
Q_MX02 U4471 ( .S(n170), .A0(stitcher_out[20]), .A1(kme_internal_word0[20]), .Z(nxt_kme_internal_word0[20]));
Q_MX02 U4472 ( .S(n170), .A0(stitcher_out[19]), .A1(kme_internal_word0[19]), .Z(nxt_kme_internal_word0[19]));
Q_MX02 U4473 ( .S(n170), .A0(stitcher_out[18]), .A1(kme_internal_word0[18]), .Z(nxt_kme_internal_word0[18]));
Q_MX02 U4474 ( .S(n170), .A0(stitcher_out[17]), .A1(kme_internal_word0[17]), .Z(nxt_kme_internal_word0[17]));
Q_MX02 U4475 ( .S(n170), .A0(stitcher_out[16]), .A1(kme_internal_word0[16]), .Z(nxt_kme_internal_word0[16]));
Q_MX02 U4476 ( .S(n170), .A0(stitcher_out[27]), .A1(kme_internal_word0[27]), .Z(nxt_kme_internal_word0[27]));
Q_MX02 U4477 ( .S(n170), .A0(stitcher_out[26]), .A1(kme_internal_word0[26]), .Z(nxt_kme_internal_word0[26]));
Q_MX02 U4478 ( .S(n170), .A0(stitcher_out[25]), .A1(kme_internal_word0[25]), .Z(nxt_kme_internal_word0[25]));
Q_MX02 U4479 ( .S(n170), .A0(stitcher_out[24]), .A1(kme_internal_word0[24]), .Z(nxt_kme_internal_word0[24]));
Q_MX02 U4480 ( .S(n170), .A0(stitcher_out[42]), .A1(kme_internal_word0[38]), .Z(nxt_kme_internal_word0[38]));
Q_MX02 U4481 ( .S(n170), .A0(stitcher_out[41]), .A1(kme_internal_word0[37]), .Z(nxt_kme_internal_word0[37]));
Q_MX02 U4482 ( .S(n170), .A0(stitcher_out[40]), .A1(kme_internal_word0[36]), .Z(nxt_kme_internal_word0[36]));
Q_MX02 U4483 ( .S(n170), .A0(stitcher_out[39]), .A1(kme_internal_word0[35]), .Z(nxt_kme_internal_word0[35]));
Q_MX02 U4484 ( .S(n170), .A0(stitcher_out[38]), .A1(kme_internal_word0[34]), .Z(nxt_kme_internal_word0[34]));
Q_MX02 U4485 ( .S(n170), .A0(stitcher_out[37]), .A1(kme_internal_word0[33]), .Z(nxt_kme_internal_word0[33]));
Q_MX02 U4486 ( .S(n170), .A0(stitcher_out[36]), .A1(kme_internal_word0[32]), .Z(nxt_kme_internal_word0[32]));
Q_MX02 U4487 ( .S(n170), .A0(stitcher_out[35]), .A1(kme_internal_word0[31]), .Z(nxt_kme_internal_word0[31]));
Q_MX02 U4488 ( .S(n170), .A0(stitcher_out[34]), .A1(kme_internal_word0[30]), .Z(nxt_kme_internal_word0[30]));
Q_MX02 U4489 ( .S(n170), .A0(stitcher_out[33]), .A1(kme_internal_word0[29]), .Z(nxt_kme_internal_word0[29]));
Q_MX02 U4490 ( .S(n170), .A0(stitcher_out[32]), .A1(kme_internal_word0[28]), .Z(nxt_kme_internal_word0[28]));
Q_MX02 U4491 ( .S(n631), .A0(stitcher_out[62]), .A1(n1656), .Z(nxt_kme_internal_word0[44]));
Q_AN02 U4492 ( .A0(n169), .A1(kme_internal_word0[44]), .Z(n1656));
Q_MX02 U4493 ( .S(n631), .A0(stitcher_out[61]), .A1(n1657), .Z(nxt_kme_internal_word0[43]));
Q_AN02 U4494 ( .A0(n169), .A1(kme_internal_word0[43]), .Z(n1657));
Q_MX02 U4495 ( .S(n631), .A0(stitcher_out[60]), .A1(n1658), .Z(nxt_kme_internal_word0[42]));
Q_AN02 U4496 ( .A0(n169), .A1(kme_internal_word0[42]), .Z(n1658));
Q_MX02 U4497 ( .S(n631), .A0(stitcher_out[59]), .A1(n1659), .Z(nxt_kme_internal_word0[41]));
Q_AN02 U4498 ( .A0(n169), .A1(kme_internal_word0[41]), .Z(n1659));
Q_MX02 U4499 ( .S(n631), .A0(stitcher_out[58]), .A1(n1660), .Z(nxt_kme_internal_word0[40]));
Q_AN02 U4500 ( .A0(n169), .A1(kme_internal_word0[40]), .Z(n1660));
Q_MX02 U4501 ( .S(n631), .A0(stitcher_out[57]), .A1(n1661), .Z(nxt_kme_internal_word0[39]));
Q_AN02 U4502 ( .A0(n169), .A1(kme_internal_word0[39]), .Z(n1661));
Q_MX02 U4503 ( .S(n631), .A0(n1696), .A1(n1662), .Z(nxt_kme_internal_word0[47]));
Q_AN02 U4504 ( .A0(n169), .A1(kme_internal_word0[47]), .Z(n1662));
Q_MX02 U4505 ( .S(n631), .A0(n1707), .A1(n1663), .Z(nxt_kme_internal_word0[48]));
Q_AN02 U4506 ( .A0(n169), .A1(kme_internal_word0[48]), .Z(n1663));
Q_AN02 U4507 ( .A0(n170), .A1(kme_internal_word0[63]), .Z(nxt_kme_internal_word0[63]));
Q_AN02 U4508 ( .A0(n170), .A1(kme_internal_word0[62]), .Z(nxt_kme_internal_word0[62]));
Q_AN02 U4509 ( .A0(n170), .A1(kme_internal_word0[61]), .Z(nxt_kme_internal_word0[61]));
Q_AN02 U4510 ( .A0(n170), .A1(kme_internal_word0[60]), .Z(nxt_kme_internal_word0[60]));
Q_AN02 U4511 ( .A0(n170), .A1(kme_internal_word0[59]), .Z(nxt_kme_internal_word0[59]));
Q_AN02 U4512 ( .A0(n170), .A1(kme_internal_word0[58]), .Z(nxt_kme_internal_word0[58]));
Q_AN02 U4513 ( .A0(n170), .A1(kme_internal_word0[57]), .Z(nxt_kme_internal_word0[57]));
Q_AN02 U4514 ( .A0(n170), .A1(kme_internal_word0[56]), .Z(nxt_kme_internal_word0[56]));
Q_AN02 U4515 ( .A0(n170), .A1(kme_internal_word0[55]), .Z(nxt_kme_internal_word0[55]));
Q_AN02 U4516 ( .A0(n170), .A1(kme_internal_word0[54]), .Z(nxt_kme_internal_word0[54]));
Q_AN02 U4517 ( .A0(n170), .A1(kme_internal_word0[53]), .Z(nxt_kme_internal_word0[53]));
Q_AN02 U4518 ( .A0(n170), .A1(kme_internal_word0[52]), .Z(nxt_kme_internal_word0[52]));
Q_AN02 U4519 ( .A0(n170), .A1(kme_internal_word0[51]), .Z(nxt_kme_internal_word0[51]));
Q_AN02 U4520 ( .A0(n170), .A1(kme_internal_word0[50]), .Z(nxt_kme_internal_word0[50]));
Q_AN02 U4521 ( .A0(n170), .A1(kme_internal_word0[49]), .Z(nxt_kme_internal_word0[49]));
Q_MX02 U4522 ( .S(skip[4]), .A0(buffer[31]), .A1(buffer[7]), .Z(n1664));
Q_MX02 U4523 ( .S(skip[4]), .A0(buffer[30]), .A1(buffer[6]), .Z(n1665));
Q_MX02 U4524 ( .S(skip[4]), .A0(buffer[29]), .A1(buffer[5]), .Z(n1666));
Q_MX02 U4525 ( .S(skip[4]), .A0(buffer[28]), .A1(buffer[4]), .Z(n1667));
Q_MX02 U4526 ( .S(skip[4]), .A0(buffer[27]), .A1(buffer[3]), .Z(n1668));
Q_MX02 U4527 ( .S(skip[4]), .A0(buffer[26]), .A1(buffer[2]), .Z(n1669));
Q_MX02 U4528 ( .S(skip[4]), .A0(buffer[25]), .A1(buffer[1]), .Z(n1670));
Q_MX02 U4529 ( .S(skip[4]), .A0(buffer[24]), .A1(buffer[0]), .Z(n1671));
Q_MX02 U4530 ( .S(skip[4]), .A0(buffer[23]), .A1(buffer[15]), .Z(n1672));
Q_MX02 U4531 ( .S(skip[4]), .A0(buffer[22]), .A1(buffer[14]), .Z(n1673));
Q_MX02 U4532 ( .S(skip[4]), .A0(buffer[21]), .A1(buffer[13]), .Z(n1674));
Q_MX02 U4533 ( .S(skip[4]), .A0(buffer[20]), .A1(buffer[12]), .Z(n1675));
Q_MX02 U4534 ( .S(skip[4]), .A0(buffer[19]), .A1(buffer[11]), .Z(n1676));
Q_MX02 U4535 ( .S(skip[4]), .A0(buffer[18]), .A1(buffer[10]), .Z(n1677));
Q_MX02 U4536 ( .S(skip[4]), .A0(buffer[17]), .A1(buffer[9]), .Z(n1678));
Q_MX02 U4537 ( .S(skip[4]), .A0(buffer[16]), .A1(buffer[8]), .Z(n1679));
Q_MX02 U4538 ( .S(skip[4]), .A0(buffer[15]), .A1(buffer[23]), .Z(n1680));
Q_MX02 U4539 ( .S(skip[4]), .A0(buffer[14]), .A1(buffer[22]), .Z(n1681));
Q_MX02 U4540 ( .S(skip[4]), .A0(buffer[13]), .A1(buffer[21]), .Z(n1682));
Q_MX02 U4541 ( .S(skip[4]), .A0(buffer[12]), .A1(buffer[20]), .Z(n1683));
Q_MX02 U4542 ( .S(skip[4]), .A0(buffer[11]), .A1(buffer[19]), .Z(n1684));
Q_MX02 U4543 ( .S(skip[4]), .A0(buffer[10]), .A1(buffer[18]), .Z(n1685));
Q_MX02 U4544 ( .S(skip[4]), .A0(buffer[9]), .A1(buffer[17]), .Z(n1686));
Q_MX02 U4545 ( .S(skip[4]), .A0(buffer[8]), .A1(buffer[16]), .Z(n1687));
Q_MX02 U4546 ( .S(skip[4]), .A0(buffer[7]), .A1(buffer[31]), .Z(n1688));
Q_MX02 U4547 ( .S(skip[4]), .A0(buffer[6]), .A1(buffer[30]), .Z(n1689));
Q_MX02 U4548 ( .S(skip[4]), .A0(buffer[5]), .A1(buffer[29]), .Z(n1690));
Q_MX02 U4549 ( .S(skip[4]), .A0(buffer[4]), .A1(buffer[28]), .Z(n1691));
Q_MX02 U4550 ( .S(skip[4]), .A0(buffer[3]), .A1(buffer[27]), .Z(n1692));
Q_MX02 U4551 ( .S(skip[4]), .A0(buffer[2]), .A1(buffer[26]), .Z(n1693));
Q_MX02 U4552 ( .S(skip[4]), .A0(buffer[1]), .A1(buffer[25]), .Z(n1694));
Q_MX02 U4553 ( .S(skip[4]), .A0(buffer[0]), .A1(buffer[24]), .Z(n1695));
Q_LDN0 _zyL492_tfiRv78_REG  ( .G(n631), .D(n1707), .Q(_zyL492_tfiRv78), .QN( ));
Q_AN02 U4555 ( .A0(n145), .A1(n140), .Z(n1696));
Q_OR02 U4556 ( .A0(stitcher_out[32]), .A1(n1698), .Z(n1697));
Q_OR03 U4557 ( .A0(stitcher_out[35]), .A1(stitcher_out[34]), .A2(n1699), .Z(n1698));
Q_INV U4558 ( .A(stitcher_out[33]), .Z(n1699));
Q_OA21 U4559 ( .A0(stitcher_out[36]), .A1(n1700), .B0(n1697), .Z(n140));
Q_OR03 U4560 ( .A0(stitcher_out[39]), .A1(stitcher_out[38]), .A2(n1701), .Z(n1700));
Q_INV U4561 ( .A(stitcher_out[37]), .Z(n1701));
Q_INV U4562 ( .A(n1702), .Z(n145));
Q_OR03 U4563 ( .A0(n1704), .A1(n1707), .A2(n1703), .Z(n1702));
Q_AN02 U4564 ( .A0(stitcher_out[40]), .A1(n32), .Z(n1703));
Q_NR02 U4565 ( .A0(n1706), .A1(n1705), .Z(n1704));
Q_OR03 U4566 ( .A0(stitcher_out[43]), .A1(stitcher_out[42]), .A2(stitcher_out[41]), .Z(n1705));
Q_INV U4567 ( .A(stitcher_out[40]), .Z(n1706));
Q_NR02 U4568 ( .A0(stitcher_out[40]), .A1(n1708), .Z(n1707));
Q_OR03 U4569 ( .A0(stitcher_out[43]), .A1(stitcher_out[42]), .A2(n1709), .Z(n1708));
Q_INV U4570 ( .A(stitcher_out[41]), .Z(n1709));
Q_AN03 U4571 ( .A0(n1711), .A1(n2040), .A2(n1717), .Z(n1710));
Q_ND02 U4572 ( .A0(n2053), .A1(n2035), .Z(n1711));
Q_AN03 U4573 ( .A0(n1715), .A1(n1714), .A2(n1713), .Z(n1712));
Q_OR02 U4574 ( .A0(n2051), .A1(n2093), .Z(n1713));
Q_OR02 U4575 ( .A0(aux_key_header[14]), .A1(aux_key_header[31]), .Z(n1714));
Q_OR02 U4576 ( .A0(n2052), .A1(n2042), .Z(n1715));
Q_OA21 U4577 ( .A0(n2051), .A1(n1994), .B0(n1716), .Z(n142));
Q_INV U4578 ( .A(n1717), .Z(n1716));
Q_OR03 U4579 ( .A0(n2106), .A1(n2110), .A2(n1718), .Z(n1717));
Q_AN02 U4580 ( .A0(aux_cipher_op[0]), .A1(n33), .Z(n1718));
Q_INV U4581 ( .A(n1719), .Z(n135));
Q_OR03 U4582 ( .A0(tlv_type[1]), .A1(n2056), .A2(n2037), .Z(n1719));
Q_OR02 U4583 ( .A0(n2057), .A1(n2056), .Z(n1720));
Q_OR03 U4584 ( .A0(stitcher_out[61]), .A1(stitcher_out[62]), .A2(always_validate_kim_ref), .Z(n141));
Q_INV U4585 ( .A(n1721), .Z(n136));
Q_OR02 U4586 ( .A0(n2056), .A1(n2055), .Z(n1721));
Q_INV U4587 ( .A(n1722), .Z(n137));
Q_OR02 U4588 ( .A0(n1723), .A1(n2036), .Z(n1722));
Q_OR03 U4589 ( .A0(tlv_type[4]), .A1(tlv_type[3]), .A2(tlv_type[2]), .Z(n1723));
Q_OR02 U4590 ( .A0(n1726), .A1(n1725), .Z(n1724));
Q_OR03 U4591 ( .A0(stitcher_out[1]), .A1(stitcher_out[0]), .A2(n1727), .Z(n1725));
Q_OR03 U4592 ( .A0(stitcher_out[4]), .A1(stitcher_out[3]), .A2(stitcher_out[2]), .Z(n1726));
Q_OR03 U4593 ( .A0(stitcher_out[7]), .A1(stitcher_out[6]), .A2(stitcher_out[5]), .Z(n1727));
Q_OR02 U4594 ( .A0(always_validate_kim_ref), .A1(n1728), .Z(n143));
Q_INV U4595 ( .A(n1728), .Z(n138));
Q_OR02 U4596 ( .A0(aux_key_type[4]), .A1(aux_key_type[5]), .Z(n1728));
Q_AN02 U4597 ( .A0(n1733), .A1(n1729), .Z(n139));
Q_AN03 U4598 ( .A0(n1730), .A1(n1731), .A2(n1732), .Z(n1729));
Q_XNR2 U4599 ( .A0(fifo_in[67]), .A1(skip[3]), .Z(n1730));
Q_XNR2 U4600 ( .A0(fifo_in[66]), .A1(skip[2]), .Z(n1731));
Q_XNR2 U4601 ( .A0(fifo_in[65]), .A1(skip[1]), .Z(n1732));
Q_XNR2 U4602 ( .A0(fifo_in[64]), .A1(skip[0]), .Z(n1733));
Q_AN02 U4603 ( .A0(n1734), .A1(skip[6]), .Z(n144));
Q_NR03 U4604 ( .A0(stitcher_empty), .A1(fifo_in_stall), .A2(skip[6]), .Z(stitcher_rd));
Q_INV U4605 ( .A(fifo_in_stall), .Z(n1734));
Q_FDP1 \tlv_type_REG[7] ( .CK(clk), .R(rst_n), .D(nxt_tlv_type[7]), .Q(tlv_type[7]), .QN( ));
Q_FDP1 \tlv_type_REG[6] ( .CK(clk), .R(rst_n), .D(nxt_tlv_type[6]), .Q(tlv_type[6]), .QN( ));
Q_FDP1 \tlv_type_REG[5] ( .CK(clk), .R(rst_n), .D(nxt_tlv_type[5]), .Q(tlv_type[5]), .QN( ));
Q_FDP1 \tlv_type_REG[4] ( .CK(clk), .R(rst_n), .D(nxt_tlv_type[4]), .Q(tlv_type[4]), .QN(n2057));
Q_FDP1 \tlv_type_REG[3] ( .CK(clk), .R(rst_n), .D(nxt_tlv_type[3]), .Q(tlv_type[3]), .QN(n2044));
Q_FDP1 \tlv_type_REG[2] ( .CK(clk), .R(rst_n), .D(nxt_tlv_type[2]), .Q(tlv_type[2]), .QN(n2058));
Q_FDP1 \tlv_type_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_tlv_type[1]), .Q(tlv_type[1]), .QN(n409));
Q_FDP1 \tlv_type_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_tlv_type[0]), .Q(tlv_type[0]), .QN(n2059));
Q_FDP1 \aux_key_type_REG[5] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_type[5]), .Q(aux_key_type[5]), .QN( ));
Q_FDP1 \aux_key_type_REG[4] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_type[4]), .Q(aux_key_type[4]), .QN( ));
Q_FDP1 \aux_key_type_REG[3] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_type[3]), .Q(aux_key_type[3]), .QN(n2071));
Q_FDP1 \aux_key_type_REG[2] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_type[2]), .Q(aux_key_type[2]), .QN(n1960));
Q_FDP1 \aux_key_type_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_type[1]), .Q(aux_key_type[1]), .QN(n1972));
Q_FDP1 \aux_key_type_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_type[0]), .Q(aux_key_type[0]), .QN(n2098));
Q_FDP1 \aux_iv_op_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_aux_iv_op[1]), .Q(aux_iv_op[1]), .QN( ));
Q_FDP1 \aux_iv_op_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_aux_iv_op[0]), .Q(aux_iv_op[0]), .QN(n2041));
Q_FDP1 \aux_cipher_op_REG[3] ( .CK(clk), .R(rst_n), .D(nxt_aux_cipher_op[3]), .Q(aux_cipher_op[3]), .QN( ));
Q_FDP1 \aux_cipher_op_REG[2] ( .CK(clk), .R(rst_n), .D(nxt_aux_cipher_op[2]), .Q(aux_cipher_op[2]), .QN( ));
Q_FDP1 \aux_cipher_op_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_aux_cipher_op[1]), .Q(aux_cipher_op[1]), .QN(n2113));
Q_FDP1 \aux_cipher_op_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_aux_cipher_op[0]), .Q(aux_cipher_op[0]), .QN(n2108));
Q_FDP1 \aux_auth_op_REG[3] ( .CK(clk), .R(rst_n), .D(nxt_aux_auth_op[3]), .Q(aux_auth_op[3]), .QN( ));
Q_FDP1 \aux_auth_op_REG[2] ( .CK(clk), .R(rst_n), .D(nxt_aux_auth_op[2]), .Q(aux_auth_op[2]), .QN( ));
Q_FDP1 \aux_auth_op_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_aux_auth_op[1]), .Q(aux_auth_op[1]), .QN(n2130));
Q_FDP1 \aux_auth_op_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_aux_auth_op[0]), .Q(aux_auth_op[0]), .QN(n2089));
Q_FDP1 \aux_raw_auth_op_REG[3] ( .CK(clk), .R(rst_n), .D(nxt_aux_raw_auth_op[3]), .Q(aux_raw_auth_op[3]), .QN( ));
Q_FDP1 \aux_raw_auth_op_REG[2] ( .CK(clk), .R(rst_n), .D(nxt_aux_raw_auth_op[2]), .Q(aux_raw_auth_op[2]), .QN( ));
Q_FDP1 \aux_raw_auth_op_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_aux_raw_auth_op[1]), .Q(aux_raw_auth_op[1]), .QN(n2126));
Q_FDP1 \aux_raw_auth_op_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_aux_raw_auth_op[0]), .Q(aux_raw_auth_op[0]), .QN(n2086));
Q_FDP1 \kme_internal_word0_REG[63] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[63]), .Q(kme_internal_word0[63]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[62] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[62]), .Q(kme_internal_word0[62]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[61] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[61]), .Q(kme_internal_word0[61]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[60] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[60]), .Q(kme_internal_word0[60]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[59] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[59]), .Q(kme_internal_word0[59]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[58] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[58]), .Q(kme_internal_word0[58]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[57] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[57]), .Q(kme_internal_word0[57]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[56] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[56]), .Q(kme_internal_word0[56]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[55] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[55]), .Q(kme_internal_word0[55]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[54] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[54]), .Q(kme_internal_word0[54]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[53] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[53]), .Q(kme_internal_word0[53]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[52] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[52]), .Q(kme_internal_word0[52]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[51] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[51]), .Q(kme_internal_word0[51]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[50] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[50]), .Q(kme_internal_word0[50]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[49] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[49]), .Q(kme_internal_word0[49]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[48] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[48]), .Q(kme_internal_word0[48]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[47] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[47]), .Q(kme_internal_word0[47]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[46] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[46]), .Q(kme_internal_word0[46]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[45] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[45]), .Q(kme_internal_word0[45]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[44] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[44]), .Q(kme_internal_word0[44]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[43] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[43]), .Q(kme_internal_word0[43]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[42] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[42]), .Q(kme_internal_word0[42]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[41] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[41]), .Q(kme_internal_word0[41]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[40] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[40]), .Q(kme_internal_word0[40]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[39] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[39]), .Q(kme_internal_word0[39]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[38] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[38]), .Q(kme_internal_word0[38]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[37] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[37]), .Q(kme_internal_word0[37]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[36] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[36]), .Q(kme_internal_word0[36]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[35] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[35]), .Q(kme_internal_word0[35]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[34] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[34]), .Q(kme_internal_word0[34]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[33] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[33]), .Q(kme_internal_word0[33]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[32] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[32]), .Q(kme_internal_word0[32]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[31] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[31]), .Q(kme_internal_word0[31]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[30] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[30]), .Q(kme_internal_word0[30]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[29] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[29]), .Q(kme_internal_word0[29]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[28] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[28]), .Q(kme_internal_word0[28]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[27] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[27]), .Q(kme_internal_word0[27]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[26] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[26]), .Q(kme_internal_word0[26]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[25] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[25]), .Q(kme_internal_word0[25]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[24] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[24]), .Q(kme_internal_word0[24]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[23] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[23]), .Q(kme_internal_word0[23]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[22] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[22]), .Q(kme_internal_word0[22]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[21] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[21]), .Q(kme_internal_word0[21]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[20] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[20]), .Q(kme_internal_word0[20]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[19] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[19]), .Q(kme_internal_word0[19]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[18] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[18]), .Q(kme_internal_word0[18]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[17] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[17]), .Q(kme_internal_word0[17]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[16] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[16]), .Q(kme_internal_word0[16]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[15] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[15]), .Q(kme_internal_word0[15]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[14] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[14]), .Q(kme_internal_word0[14]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[13] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[13]), .Q(kme_internal_word0[13]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[12] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[12]), .Q(kme_internal_word0[12]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[11] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[11]), .Q(kme_internal_word0[11]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[10] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[10]), .Q(kme_internal_word0[10]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[9] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[9]), .Q(kme_internal_word0[9]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[8] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[8]), .Q(kme_internal_word0[8]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[7] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[7]), .Q(kme_internal_word0[7]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[6] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[6]), .Q(kme_internal_word0[6]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[5] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[5]), .Q(kme_internal_word0[5]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[4] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[4]), .Q(kme_internal_word0[4]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[3] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[3]), .Q(kme_internal_word0[3]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[2] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[2]), .Q(kme_internal_word0[2]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[1]), .Q(kme_internal_word0[1]), .QN( ));
Q_FDP1 \kme_internal_word0_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_word0[0]), .Q(kme_internal_word0[0]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[63] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[63]), .Q(kme_internal_dek_kim_word[63]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[62] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[62]), .Q(kme_internal_dek_kim_word[62]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[61] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[61]), .Q(kme_internal_dek_kim_word[61]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[60] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[60]), .Q(kme_internal_dek_kim_word[60]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[59] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[59]), .Q(kme_internal_dek_kim_word[59]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[58] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[58]), .Q(kme_internal_dek_kim_word[58]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[57] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[57]), .Q(kme_internal_dek_kim_word[57]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[56] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[56]), .Q(kme_internal_dek_kim_word[56]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[55] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[55]), .Q(kme_internal_dek_kim_word[55]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[54] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[54]), .Q(kme_internal_dek_kim_word[54]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[53] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[53]), .Q(kme_internal_dek_kim_word[53]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[52] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[52]), .Q(kme_internal_dek_kim_word[52]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[51] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[51]), .Q(kme_internal_dek_kim_word[51]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[50] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[50]), .Q(kme_internal_dek_kim_word[50]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[49] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[49]), .Q(kme_internal_dek_kim_word[49]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[48] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[48]), .Q(kme_internal_dek_kim_word[48]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[47] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[47]), .Q(kme_internal_dek_kim_word[47]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[46] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[46]), .Q(kme_internal_dek_kim_word[46]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[45] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[45]), .Q(kme_internal_dek_kim_word[45]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[44] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[44]), .Q(kme_internal_dek_kim_word[44]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[43] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[43]), .Q(kme_internal_dek_kim_word[43]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[42] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[42]), .Q(kme_internal_dek_kim_word[42]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[41] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[41]), .Q(kme_internal_dek_kim_word[41]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[40] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[40]), .Q(kme_internal_dek_kim_word[40]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[39] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[39]), .Q(kme_internal_dek_kim_word[39]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[38] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[38]), .Q(kme_internal_dek_kim_word[38]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[37] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[37]), .Q(kme_internal_dek_kim_word[37]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[36] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[36]), .Q(kme_internal_dek_kim_word[36]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[35] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[35]), .Q(kme_internal_dek_kim_word[35]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[34] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[34]), .Q(kme_internal_dek_kim_word[34]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[33] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[33]), .Q(kme_internal_dek_kim_word[33]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[32] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[32]), .Q(kme_internal_dek_kim_word[32]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[31] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[31]), .Q(kme_internal_dek_kim_word[31]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[30] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[30]), .Q(kme_internal_dek_kim_word[30]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[29] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[29]), .Q(kme_internal_dek_kim_word[29]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[28] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[28]), .Q(kme_internal_dek_kim_word[28]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[27] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[27]), .Q(kme_internal_dek_kim_word[27]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[26] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[26]), .Q(kme_internal_dek_kim_word[26]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[25] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[25]), .Q(kme_internal_dek_kim_word[25]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[24] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[24]), .Q(kme_internal_dek_kim_word[24]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[23] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[23]), .Q(kme_internal_dek_kim_word[23]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[22] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[22]), .Q(kme_internal_dek_kim_word[22]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[21] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[21]), .Q(kme_internal_dek_kim_word[21]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[20] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[20]), .Q(kme_internal_dek_kim_word[20]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[19] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[19]), .Q(kme_internal_dek_kim_word[19]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[18] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[18]), .Q(kme_internal_dek_kim_word[18]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[17] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[17]), .Q(kme_internal_dek_kim_word[17]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[16] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[16]), .Q(kme_internal_dek_kim_word[16]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[15] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[15]), .Q(kme_internal_dek_kim_word[15]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[14] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[14]), .Q(kme_internal_dek_kim_word[14]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[13] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[13]), .Q(kme_internal_dek_kim_word[13]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[12] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[12]), .Q(kme_internal_dek_kim_word[12]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[11] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[11]), .Q(kme_internal_dek_kim_word[11]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[10] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[10]), .Q(kme_internal_dek_kim_word[10]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[9] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[9]), .Q(kme_internal_dek_kim_word[9]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[8] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[8]), .Q(kme_internal_dek_kim_word[8]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[7] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[7]), .Q(kme_internal_dek_kim_word[7]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[6] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[6]), .Q(kme_internal_dek_kim_word[6]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[5] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[5]), .Q(kme_internal_dek_kim_word[5]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[4] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[4]), .Q(kme_internal_dek_kim_word[4]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[3] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[3]), .Q(kme_internal_dek_kim_word[3]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[2] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[2]), .Q(kme_internal_dek_kim_word[2]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[1]), .Q(kme_internal_dek_kim_word[1]), .QN( ));
Q_FDP1 \kme_internal_dek_kim_word_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dek_kim_word[0]), .Q(kme_internal_dek_kim_word[0]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[63] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[63]), .Q(kme_internal_dak_kim_word[63]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[62] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[62]), .Q(kme_internal_dak_kim_word[62]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[61] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[61]), .Q(kme_internal_dak_kim_word[61]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[60] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[60]), .Q(kme_internal_dak_kim_word[60]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[59] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[59]), .Q(kme_internal_dak_kim_word[59]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[58] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[58]), .Q(kme_internal_dak_kim_word[58]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[57] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[57]), .Q(kme_internal_dak_kim_word[57]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[56] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[56]), .Q(kme_internal_dak_kim_word[56]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[55] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[55]), .Q(kme_internal_dak_kim_word[55]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[54] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[54]), .Q(kme_internal_dak_kim_word[54]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[53] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[53]), .Q(kme_internal_dak_kim_word[53]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[52] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[52]), .Q(kme_internal_dak_kim_word[52]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[51] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[51]), .Q(kme_internal_dak_kim_word[51]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[50] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[50]), .Q(kme_internal_dak_kim_word[50]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[49] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[49]), .Q(kme_internal_dak_kim_word[49]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[48] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[48]), .Q(kme_internal_dak_kim_word[48]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[47] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[47]), .Q(kme_internal_dak_kim_word[47]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[46] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[46]), .Q(kme_internal_dak_kim_word[46]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[45] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[45]), .Q(kme_internal_dak_kim_word[45]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[44] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[44]), .Q(kme_internal_dak_kim_word[44]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[43] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[43]), .Q(kme_internal_dak_kim_word[43]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[42] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[42]), .Q(kme_internal_dak_kim_word[42]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[41] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[41]), .Q(kme_internal_dak_kim_word[41]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[40] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[40]), .Q(kme_internal_dak_kim_word[40]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[39] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[39]), .Q(kme_internal_dak_kim_word[39]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[38] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[38]), .Q(kme_internal_dak_kim_word[38]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[37] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[37]), .Q(kme_internal_dak_kim_word[37]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[36] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[36]), .Q(kme_internal_dak_kim_word[36]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[35] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[35]), .Q(kme_internal_dak_kim_word[35]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[34] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[34]), .Q(kme_internal_dak_kim_word[34]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[33] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[33]), .Q(kme_internal_dak_kim_word[33]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[32] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[32]), .Q(kme_internal_dak_kim_word[32]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[31] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[31]), .Q(kme_internal_dak_kim_word[31]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[30] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[30]), .Q(kme_internal_dak_kim_word[30]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[29] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[29]), .Q(kme_internal_dak_kim_word[29]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[28] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[28]), .Q(kme_internal_dak_kim_word[28]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[27] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[27]), .Q(kme_internal_dak_kim_word[27]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[26] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[26]), .Q(kme_internal_dak_kim_word[26]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[25] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[25]), .Q(kme_internal_dak_kim_word[25]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[24] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[24]), .Q(kme_internal_dak_kim_word[24]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[23] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[23]), .Q(kme_internal_dak_kim_word[23]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[22] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[22]), .Q(kme_internal_dak_kim_word[22]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[21] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[21]), .Q(kme_internal_dak_kim_word[21]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[20] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[20]), .Q(kme_internal_dak_kim_word[20]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[19] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[19]), .Q(kme_internal_dak_kim_word[19]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[18] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[18]), .Q(kme_internal_dak_kim_word[18]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[17] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[17]), .Q(kme_internal_dak_kim_word[17]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[16] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[16]), .Q(kme_internal_dak_kim_word[16]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[15] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[15]), .Q(kme_internal_dak_kim_word[15]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[14] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[14]), .Q(kme_internal_dak_kim_word[14]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[13] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[13]), .Q(kme_internal_dak_kim_word[13]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[12] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[12]), .Q(kme_internal_dak_kim_word[12]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[11] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[11]), .Q(kme_internal_dak_kim_word[11]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[10] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[10]), .Q(kme_internal_dak_kim_word[10]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[9] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[9]), .Q(kme_internal_dak_kim_word[9]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[8] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[8]), .Q(kme_internal_dak_kim_word[8]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[7] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[7]), .Q(kme_internal_dak_kim_word[7]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[6] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[6]), .Q(kme_internal_dak_kim_word[6]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[5] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[5]), .Q(kme_internal_dak_kim_word[5]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[4] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[4]), .Q(kme_internal_dak_kim_word[4]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[3] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[3]), .Q(kme_internal_dak_kim_word[3]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[2] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[2]), .Q(kme_internal_dak_kim_word[2]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[1]), .Q(kme_internal_dak_kim_word[1]), .QN( ));
Q_FDP1 \kme_internal_dak_kim_word_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_kme_internal_dak_kim_word[0]), .Q(kme_internal_dak_kim_word[0]), .QN( ));
Q_FDP1 \debug_cmd_REG[31] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[31]), .Q(debug_cmd[31]), .QN( ));
Q_FDP1 \debug_cmd_REG[30] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[30]), .Q(debug_cmd[30]), .QN( ));
Q_FDP1 \debug_cmd_REG[29] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[29]), .Q(debug_cmd[29]), .QN( ));
Q_FDP1 \debug_cmd_REG[28] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[28]), .Q(debug_cmd[28]), .QN( ));
Q_FDP1 \debug_cmd_REG[27] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[27]), .Q(debug_cmd[27]), .QN( ));
Q_FDP1 \debug_cmd_REG[26] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[26]), .Q(debug_cmd[26]), .QN( ));
Q_FDP1 \debug_cmd_REG[25] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[25]), .Q(debug_cmd[25]), .QN( ));
Q_FDP1 \debug_cmd_REG[24] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[24]), .Q(debug_cmd[24]), .QN( ));
Q_FDP1 \debug_cmd_REG[23] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[23]), .Q(debug_cmd[23]), .QN( ));
Q_FDP1 \debug_cmd_REG[22] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[22]), .Q(debug_cmd[22]), .QN( ));
Q_FDP1 \debug_cmd_REG[21] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[21]), .Q(debug_cmd[21]), .QN( ));
Q_FDP1 \debug_cmd_REG[20] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[20]), .Q(debug_cmd[20]), .QN( ));
Q_FDP1 \debug_cmd_REG[19] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[19]), .Q(debug_cmd[19]), .QN( ));
Q_FDP1 \debug_cmd_REG[18] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[18]), .Q(debug_cmd[18]), .QN( ));
Q_FDP1 \debug_cmd_REG[17] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[17]), .Q(debug_cmd[17]), .QN( ));
Q_FDP1 \debug_cmd_REG[16] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[16]), .Q(debug_cmd[16]), .QN( ));
Q_FDP1 \debug_cmd_REG[15] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[15]), .Q(debug_cmd[15]), .QN( ));
Q_FDP1 \debug_cmd_REG[14] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[14]), .Q(debug_cmd[14]), .QN( ));
Q_FDP1 \debug_cmd_REG[13] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[13]), .Q(debug_cmd[13]), .QN( ));
Q_FDP1 \debug_cmd_REG[12] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[12]), .Q(debug_cmd[12]), .QN( ));
Q_FDP1 \debug_cmd_REG[11] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[11]), .Q(debug_cmd[11]), .QN( ));
Q_FDP1 \debug_cmd_REG[10] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[10]), .Q(debug_cmd[10]), .QN( ));
Q_FDP1 \debug_cmd_REG[9] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[9]), .Q(debug_cmd[9]), .QN( ));
Q_FDP1 \debug_cmd_REG[8] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[8]), .Q(debug_cmd[8]), .QN( ));
Q_FDP1 \debug_cmd_REG[7] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[7]), .Q(debug_cmd[7]), .QN( ));
Q_FDP1 \debug_cmd_REG[6] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[6]), .Q(debug_cmd[6]), .QN( ));
Q_FDP1 \debug_cmd_REG[5] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[5]), .Q(debug_cmd[5]), .QN( ));
Q_FDP1 \debug_cmd_REG[4] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[4]), .Q(debug_cmd[4]), .QN( ));
Q_FDP1 \debug_cmd_REG[3] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[3]), .Q(debug_cmd[3]), .QN( ));
Q_FDP1 \debug_cmd_REG[2] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[2]), .Q(debug_cmd[2]), .QN( ));
Q_FDP1 \debug_cmd_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[1]), .Q(debug_cmd[1]), .QN( ));
Q_FDP1 \debug_cmd_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_debug_cmd[0]), .Q(debug_cmd[0]), .QN( ));
Q_FDP1 \aux_key_header_REG[31] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[31]), .Q(aux_key_header[31]), .QN(n2050));
Q_FDP1 \aux_key_header_REG[30] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[30]), .Q(aux_key_header[30]), .QN( ));
Q_FDP1 \aux_key_header_REG[29] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[29]), .Q(aux_key_header[29]), .QN( ));
Q_FDP1 \aux_key_header_REG[28] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[28]), .Q(aux_key_header[28]), .QN( ));
Q_FDP1 \aux_key_header_REG[27] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[27]), .Q(aux_key_header[27]), .QN( ));
Q_FDP1 \aux_key_header_REG[26] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[26]), .Q(aux_key_header[26]), .QN( ));
Q_FDP1 \aux_key_header_REG[25] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[25]), .Q(aux_key_header[25]), .QN( ));
Q_FDP1 \aux_key_header_REG[24] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[24]), .Q(aux_key_header[24]), .QN( ));
Q_FDP1 \aux_key_header_REG[23] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[23]), .Q(aux_key_header[23]), .QN( ));
Q_FDP1 \aux_key_header_REG[22] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[22]), .Q(aux_key_header[22]), .QN( ));
Q_FDP1 \aux_key_header_REG[21] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[21]), .Q(aux_key_header[21]), .QN( ));
Q_FDP1 \aux_key_header_REG[20] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[20]), .Q(aux_key_header[20]), .QN( ));
Q_FDP1 \aux_key_header_REG[19] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[19]), .Q(aux_key_header[19]), .QN( ));
Q_FDP1 \aux_key_header_REG[18] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[18]), .Q(aux_key_header[18]), .QN( ));
Q_FDP1 \aux_key_header_REG[17] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[17]), .Q(aux_key_header[17]), .QN( ));
Q_FDP1 \aux_key_header_REG[16] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[16]), .Q(aux_key_header[16]), .QN(n1995));
Q_FDP1 \aux_key_header_REG[15] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[15]), .Q(aux_key_header[15]), .QN(n2094));
Q_FDP1 \aux_key_header_REG[14] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[14]), .Q(aux_key_header[14]), .QN(n2048));
Q_FDP1 \aux_key_header_REG[13] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[13]), .Q(aux_key_header[13]), .QN( ));
Q_FDP1 \aux_key_header_REG[12] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[12]), .Q(aux_key_header[12]), .QN( ));
Q_FDP1 \aux_key_header_REG[11] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[11]), .Q(aux_key_header[11]), .QN( ));
Q_FDP1 \aux_key_header_REG[10] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[10]), .Q(aux_key_header[10]), .QN( ));
Q_FDP1 \aux_key_header_REG[9] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[9]), .Q(aux_key_header[9]), .QN( ));
Q_FDP1 \aux_key_header_REG[8] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[8]), .Q(aux_key_header[8]), .QN( ));
Q_FDP1 \aux_key_header_REG[7] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[7]), .Q(aux_key_header[7]), .QN( ));
Q_FDP1 \aux_key_header_REG[6] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[6]), .Q(aux_key_header[6]), .QN( ));
Q_FDP1 \aux_key_header_REG[5] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[5]), .Q(aux_key_header[5]), .QN( ));
Q_FDP1 \aux_key_header_REG[4] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[4]), .Q(aux_key_header[4]), .QN( ));
Q_FDP1 \aux_key_header_REG[3] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[3]), .Q(aux_key_header[3]), .QN( ));
Q_FDP1 \aux_key_header_REG[2] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[2]), .Q(aux_key_header[2]), .QN( ));
Q_FDP1 \aux_key_header_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[1]), .Q(aux_key_header[1]), .QN( ));
Q_FDP1 \aux_key_header_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_aux_key_header[0]), .Q(aux_key_header[0]), .QN( ));
Q_FDP1 \skip_REG[6] ( .CK(clk), .R(rst_n), .D(nxt_skip[6]), .Q(skip[6]), .QN( ));
Q_FDP1 \skip_REG[5] ( .CK(clk), .R(rst_n), .D(nxt_skip[5]), .Q(skip[5]), .QN( ));
Q_FDP1 \skip_REG[4] ( .CK(clk), .R(rst_n), .D(nxt_skip[4]), .Q(skip[4]), .QN( ));
Q_FDP1 \skip_REG[3] ( .CK(clk), .R(rst_n), .D(nxt_skip[3]), .Q(skip[3]), .QN( ));
Q_FDP1 \skip_REG[2] ( .CK(clk), .R(rst_n), .D(nxt_skip[2]), .Q(skip[2]), .QN( ));
Q_FDP1 \skip_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_skip[1]), .Q(skip[1]), .QN( ));
Q_FDP1 \skip_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_skip[0]), .Q(skip[0]), .QN( ));
Q_FDP1 \guid0_REG[63] ( .CK(clk), .R(rst_n), .D(nxt_guid0[63]), .Q(guid0[63]), .QN( ));
Q_FDP1 \guid0_REG[62] ( .CK(clk), .R(rst_n), .D(nxt_guid0[62]), .Q(guid0[62]), .QN( ));
Q_FDP1 \guid0_REG[61] ( .CK(clk), .R(rst_n), .D(nxt_guid0[61]), .Q(guid0[61]), .QN( ));
Q_FDP1 \guid0_REG[60] ( .CK(clk), .R(rst_n), .D(nxt_guid0[60]), .Q(guid0[60]), .QN( ));
Q_FDP1 \guid0_REG[59] ( .CK(clk), .R(rst_n), .D(nxt_guid0[59]), .Q(guid0[59]), .QN( ));
Q_FDP1 \guid0_REG[58] ( .CK(clk), .R(rst_n), .D(nxt_guid0[58]), .Q(guid0[58]), .QN( ));
Q_FDP1 \guid0_REG[57] ( .CK(clk), .R(rst_n), .D(nxt_guid0[57]), .Q(guid0[57]), .QN( ));
Q_FDP1 \guid0_REG[56] ( .CK(clk), .R(rst_n), .D(nxt_guid0[56]), .Q(guid0[56]), .QN( ));
Q_FDP1 \guid0_REG[55] ( .CK(clk), .R(rst_n), .D(nxt_guid0[55]), .Q(guid0[55]), .QN( ));
Q_FDP1 \guid0_REG[54] ( .CK(clk), .R(rst_n), .D(nxt_guid0[54]), .Q(guid0[54]), .QN( ));
Q_FDP1 \guid0_REG[53] ( .CK(clk), .R(rst_n), .D(nxt_guid0[53]), .Q(guid0[53]), .QN( ));
Q_FDP1 \guid0_REG[52] ( .CK(clk), .R(rst_n), .D(nxt_guid0[52]), .Q(guid0[52]), .QN( ));
Q_FDP1 \guid0_REG[51] ( .CK(clk), .R(rst_n), .D(nxt_guid0[51]), .Q(guid0[51]), .QN( ));
Q_FDP1 \guid0_REG[50] ( .CK(clk), .R(rst_n), .D(nxt_guid0[50]), .Q(guid0[50]), .QN( ));
Q_FDP1 \guid0_REG[49] ( .CK(clk), .R(rst_n), .D(nxt_guid0[49]), .Q(guid0[49]), .QN( ));
Q_FDP1 \guid0_REG[48] ( .CK(clk), .R(rst_n), .D(nxt_guid0[48]), .Q(guid0[48]), .QN( ));
Q_FDP1 \guid0_REG[47] ( .CK(clk), .R(rst_n), .D(nxt_guid0[47]), .Q(guid0[47]), .QN( ));
Q_FDP1 \guid0_REG[46] ( .CK(clk), .R(rst_n), .D(nxt_guid0[46]), .Q(guid0[46]), .QN( ));
Q_FDP1 \guid0_REG[45] ( .CK(clk), .R(rst_n), .D(nxt_guid0[45]), .Q(guid0[45]), .QN( ));
Q_FDP1 \guid0_REG[44] ( .CK(clk), .R(rst_n), .D(nxt_guid0[44]), .Q(guid0[44]), .QN( ));
Q_FDP1 \guid0_REG[43] ( .CK(clk), .R(rst_n), .D(nxt_guid0[43]), .Q(guid0[43]), .QN( ));
Q_FDP1 \guid0_REG[42] ( .CK(clk), .R(rst_n), .D(nxt_guid0[42]), .Q(guid0[42]), .QN( ));
Q_FDP1 \guid0_REG[41] ( .CK(clk), .R(rst_n), .D(nxt_guid0[41]), .Q(guid0[41]), .QN( ));
Q_FDP1 \guid0_REG[40] ( .CK(clk), .R(rst_n), .D(nxt_guid0[40]), .Q(guid0[40]), .QN( ));
Q_FDP1 \guid0_REG[39] ( .CK(clk), .R(rst_n), .D(nxt_guid0[39]), .Q(guid0[39]), .QN( ));
Q_FDP1 \guid0_REG[38] ( .CK(clk), .R(rst_n), .D(nxt_guid0[38]), .Q(guid0[38]), .QN( ));
Q_FDP1 \guid0_REG[37] ( .CK(clk), .R(rst_n), .D(nxt_guid0[37]), .Q(guid0[37]), .QN( ));
Q_FDP1 \guid0_REG[36] ( .CK(clk), .R(rst_n), .D(nxt_guid0[36]), .Q(guid0[36]), .QN( ));
Q_FDP1 \guid0_REG[35] ( .CK(clk), .R(rst_n), .D(nxt_guid0[35]), .Q(guid0[35]), .QN( ));
Q_FDP1 \guid0_REG[34] ( .CK(clk), .R(rst_n), .D(nxt_guid0[34]), .Q(guid0[34]), .QN( ));
Q_FDP1 \guid0_REG[33] ( .CK(clk), .R(rst_n), .D(nxt_guid0[33]), .Q(guid0[33]), .QN( ));
Q_FDP1 \guid0_REG[32] ( .CK(clk), .R(rst_n), .D(nxt_guid0[32]), .Q(guid0[32]), .QN( ));
Q_FDP1 \guid0_REG[31] ( .CK(clk), .R(rst_n), .D(nxt_guid0[31]), .Q(guid0[31]), .QN( ));
Q_FDP1 \guid0_REG[30] ( .CK(clk), .R(rst_n), .D(nxt_guid0[30]), .Q(guid0[30]), .QN( ));
Q_FDP1 \guid0_REG[29] ( .CK(clk), .R(rst_n), .D(nxt_guid0[29]), .Q(guid0[29]), .QN( ));
Q_FDP1 \guid0_REG[28] ( .CK(clk), .R(rst_n), .D(nxt_guid0[28]), .Q(guid0[28]), .QN( ));
Q_FDP1 \guid0_REG[27] ( .CK(clk), .R(rst_n), .D(nxt_guid0[27]), .Q(guid0[27]), .QN( ));
Q_FDP1 \guid0_REG[26] ( .CK(clk), .R(rst_n), .D(nxt_guid0[26]), .Q(guid0[26]), .QN( ));
Q_FDP1 \guid0_REG[25] ( .CK(clk), .R(rst_n), .D(nxt_guid0[25]), .Q(guid0[25]), .QN( ));
Q_FDP1 \guid0_REG[24] ( .CK(clk), .R(rst_n), .D(nxt_guid0[24]), .Q(guid0[24]), .QN( ));
Q_FDP1 \guid0_REG[23] ( .CK(clk), .R(rst_n), .D(nxt_guid0[23]), .Q(guid0[23]), .QN( ));
Q_FDP1 \guid0_REG[22] ( .CK(clk), .R(rst_n), .D(nxt_guid0[22]), .Q(guid0[22]), .QN( ));
Q_FDP1 \guid0_REG[21] ( .CK(clk), .R(rst_n), .D(nxt_guid0[21]), .Q(guid0[21]), .QN( ));
Q_FDP1 \guid0_REG[20] ( .CK(clk), .R(rst_n), .D(nxt_guid0[20]), .Q(guid0[20]), .QN( ));
Q_FDP1 \guid0_REG[19] ( .CK(clk), .R(rst_n), .D(nxt_guid0[19]), .Q(guid0[19]), .QN( ));
Q_FDP1 \guid0_REG[18] ( .CK(clk), .R(rst_n), .D(nxt_guid0[18]), .Q(guid0[18]), .QN( ));
Q_FDP1 \guid0_REG[17] ( .CK(clk), .R(rst_n), .D(nxt_guid0[17]), .Q(guid0[17]), .QN( ));
Q_FDP1 \guid0_REG[16] ( .CK(clk), .R(rst_n), .D(nxt_guid0[16]), .Q(guid0[16]), .QN( ));
Q_FDP1 \guid0_REG[15] ( .CK(clk), .R(rst_n), .D(nxt_guid0[15]), .Q(guid0[15]), .QN( ));
Q_FDP1 \guid0_REG[14] ( .CK(clk), .R(rst_n), .D(nxt_guid0[14]), .Q(guid0[14]), .QN( ));
Q_FDP1 \guid0_REG[13] ( .CK(clk), .R(rst_n), .D(nxt_guid0[13]), .Q(guid0[13]), .QN( ));
Q_FDP1 \guid0_REG[12] ( .CK(clk), .R(rst_n), .D(nxt_guid0[12]), .Q(guid0[12]), .QN( ));
Q_FDP1 \guid0_REG[11] ( .CK(clk), .R(rst_n), .D(nxt_guid0[11]), .Q(guid0[11]), .QN( ));
Q_FDP1 \guid0_REG[10] ( .CK(clk), .R(rst_n), .D(nxt_guid0[10]), .Q(guid0[10]), .QN( ));
Q_FDP1 \guid0_REG[9] ( .CK(clk), .R(rst_n), .D(nxt_guid0[9]), .Q(guid0[9]), .QN( ));
Q_FDP1 \guid0_REG[8] ( .CK(clk), .R(rst_n), .D(nxt_guid0[8]), .Q(guid0[8]), .QN( ));
Q_FDP1 \guid0_REG[7] ( .CK(clk), .R(rst_n), .D(nxt_guid0[7]), .Q(guid0[7]), .QN( ));
Q_FDP1 \guid0_REG[6] ( .CK(clk), .R(rst_n), .D(nxt_guid0[6]), .Q(guid0[6]), .QN( ));
Q_FDP1 \guid0_REG[5] ( .CK(clk), .R(rst_n), .D(nxt_guid0[5]), .Q(guid0[5]), .QN( ));
Q_FDP1 \guid0_REG[4] ( .CK(clk), .R(rst_n), .D(nxt_guid0[4]), .Q(guid0[4]), .QN( ));
Q_FDP1 \guid0_REG[3] ( .CK(clk), .R(rst_n), .D(nxt_guid0[3]), .Q(guid0[3]), .QN( ));
Q_FDP1 \guid0_REG[2] ( .CK(clk), .R(rst_n), .D(nxt_guid0[2]), .Q(guid0[2]), .QN( ));
Q_FDP1 \guid0_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_guid0[1]), .Q(guid0[1]), .QN( ));
Q_FDP1 \guid0_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_guid0[0]), .Q(guid0[0]), .QN( ));
Q_FDP1 \guid1_REG[63] ( .CK(clk), .R(rst_n), .D(nxt_guid1[63]), .Q(guid1[63]), .QN( ));
Q_FDP1 \guid1_REG[62] ( .CK(clk), .R(rst_n), .D(nxt_guid1[62]), .Q(guid1[62]), .QN( ));
Q_FDP1 \guid1_REG[61] ( .CK(clk), .R(rst_n), .D(nxt_guid1[61]), .Q(guid1[61]), .QN( ));
Q_FDP1 \guid1_REG[60] ( .CK(clk), .R(rst_n), .D(nxt_guid1[60]), .Q(guid1[60]), .QN( ));
Q_FDP1 \guid1_REG[59] ( .CK(clk), .R(rst_n), .D(nxt_guid1[59]), .Q(guid1[59]), .QN( ));
Q_FDP1 \guid1_REG[58] ( .CK(clk), .R(rst_n), .D(nxt_guid1[58]), .Q(guid1[58]), .QN( ));
Q_FDP1 \guid1_REG[57] ( .CK(clk), .R(rst_n), .D(nxt_guid1[57]), .Q(guid1[57]), .QN( ));
Q_FDP1 \guid1_REG[56] ( .CK(clk), .R(rst_n), .D(nxt_guid1[56]), .Q(guid1[56]), .QN( ));
Q_FDP1 \guid1_REG[55] ( .CK(clk), .R(rst_n), .D(nxt_guid1[55]), .Q(guid1[55]), .QN( ));
Q_FDP1 \guid1_REG[54] ( .CK(clk), .R(rst_n), .D(nxt_guid1[54]), .Q(guid1[54]), .QN( ));
Q_FDP1 \guid1_REG[53] ( .CK(clk), .R(rst_n), .D(nxt_guid1[53]), .Q(guid1[53]), .QN( ));
Q_FDP1 \guid1_REG[52] ( .CK(clk), .R(rst_n), .D(nxt_guid1[52]), .Q(guid1[52]), .QN( ));
Q_FDP1 \guid1_REG[51] ( .CK(clk), .R(rst_n), .D(nxt_guid1[51]), .Q(guid1[51]), .QN( ));
Q_FDP1 \guid1_REG[50] ( .CK(clk), .R(rst_n), .D(nxt_guid1[50]), .Q(guid1[50]), .QN( ));
Q_FDP1 \guid1_REG[49] ( .CK(clk), .R(rst_n), .D(nxt_guid1[49]), .Q(guid1[49]), .QN( ));
Q_FDP1 \guid1_REG[48] ( .CK(clk), .R(rst_n), .D(nxt_guid1[48]), .Q(guid1[48]), .QN( ));
Q_FDP1 \guid1_REG[47] ( .CK(clk), .R(rst_n), .D(nxt_guid1[47]), .Q(guid1[47]), .QN( ));
Q_FDP1 \guid1_REG[46] ( .CK(clk), .R(rst_n), .D(nxt_guid1[46]), .Q(guid1[46]), .QN( ));
Q_FDP1 \guid1_REG[45] ( .CK(clk), .R(rst_n), .D(nxt_guid1[45]), .Q(guid1[45]), .QN( ));
Q_FDP1 \guid1_REG[44] ( .CK(clk), .R(rst_n), .D(nxt_guid1[44]), .Q(guid1[44]), .QN( ));
Q_FDP1 \guid1_REG[43] ( .CK(clk), .R(rst_n), .D(nxt_guid1[43]), .Q(guid1[43]), .QN( ));
Q_FDP1 \guid1_REG[42] ( .CK(clk), .R(rst_n), .D(nxt_guid1[42]), .Q(guid1[42]), .QN( ));
Q_FDP1 \guid1_REG[41] ( .CK(clk), .R(rst_n), .D(nxt_guid1[41]), .Q(guid1[41]), .QN( ));
Q_FDP1 \guid1_REG[40] ( .CK(clk), .R(rst_n), .D(nxt_guid1[40]), .Q(guid1[40]), .QN( ));
Q_FDP1 \guid1_REG[39] ( .CK(clk), .R(rst_n), .D(nxt_guid1[39]), .Q(guid1[39]), .QN( ));
Q_FDP1 \guid1_REG[38] ( .CK(clk), .R(rst_n), .D(nxt_guid1[38]), .Q(guid1[38]), .QN( ));
Q_FDP1 \guid1_REG[37] ( .CK(clk), .R(rst_n), .D(nxt_guid1[37]), .Q(guid1[37]), .QN( ));
Q_FDP1 \guid1_REG[36] ( .CK(clk), .R(rst_n), .D(nxt_guid1[36]), .Q(guid1[36]), .QN( ));
Q_FDP1 \guid1_REG[35] ( .CK(clk), .R(rst_n), .D(nxt_guid1[35]), .Q(guid1[35]), .QN( ));
Q_FDP1 \guid1_REG[34] ( .CK(clk), .R(rst_n), .D(nxt_guid1[34]), .Q(guid1[34]), .QN( ));
Q_FDP1 \guid1_REG[33] ( .CK(clk), .R(rst_n), .D(nxt_guid1[33]), .Q(guid1[33]), .QN( ));
Q_FDP1 \guid1_REG[32] ( .CK(clk), .R(rst_n), .D(nxt_guid1[32]), .Q(guid1[32]), .QN( ));
Q_FDP1 \guid1_REG[31] ( .CK(clk), .R(rst_n), .D(nxt_guid1[31]), .Q(guid1[31]), .QN( ));
Q_FDP1 \guid1_REG[30] ( .CK(clk), .R(rst_n), .D(nxt_guid1[30]), .Q(guid1[30]), .QN( ));
Q_FDP1 \guid1_REG[29] ( .CK(clk), .R(rst_n), .D(nxt_guid1[29]), .Q(guid1[29]), .QN( ));
Q_FDP1 \guid1_REG[28] ( .CK(clk), .R(rst_n), .D(nxt_guid1[28]), .Q(guid1[28]), .QN( ));
Q_FDP1 \guid1_REG[27] ( .CK(clk), .R(rst_n), .D(nxt_guid1[27]), .Q(guid1[27]), .QN( ));
Q_FDP1 \guid1_REG[26] ( .CK(clk), .R(rst_n), .D(nxt_guid1[26]), .Q(guid1[26]), .QN( ));
Q_FDP1 \guid1_REG[25] ( .CK(clk), .R(rst_n), .D(nxt_guid1[25]), .Q(guid1[25]), .QN( ));
Q_FDP1 \guid1_REG[24] ( .CK(clk), .R(rst_n), .D(nxt_guid1[24]), .Q(guid1[24]), .QN( ));
Q_FDP1 \guid1_REG[23] ( .CK(clk), .R(rst_n), .D(nxt_guid1[23]), .Q(guid1[23]), .QN( ));
Q_FDP1 \guid1_REG[22] ( .CK(clk), .R(rst_n), .D(nxt_guid1[22]), .Q(guid1[22]), .QN( ));
Q_FDP1 \guid1_REG[21] ( .CK(clk), .R(rst_n), .D(nxt_guid1[21]), .Q(guid1[21]), .QN( ));
Q_FDP1 \guid1_REG[20] ( .CK(clk), .R(rst_n), .D(nxt_guid1[20]), .Q(guid1[20]), .QN( ));
Q_FDP1 \guid1_REG[19] ( .CK(clk), .R(rst_n), .D(nxt_guid1[19]), .Q(guid1[19]), .QN( ));
Q_FDP1 \guid1_REG[18] ( .CK(clk), .R(rst_n), .D(nxt_guid1[18]), .Q(guid1[18]), .QN( ));
Q_FDP1 \guid1_REG[17] ( .CK(clk), .R(rst_n), .D(nxt_guid1[17]), .Q(guid1[17]), .QN( ));
Q_FDP1 \guid1_REG[16] ( .CK(clk), .R(rst_n), .D(nxt_guid1[16]), .Q(guid1[16]), .QN( ));
Q_FDP1 \guid1_REG[15] ( .CK(clk), .R(rst_n), .D(nxt_guid1[15]), .Q(guid1[15]), .QN( ));
Q_FDP1 \guid1_REG[14] ( .CK(clk), .R(rst_n), .D(nxt_guid1[14]), .Q(guid1[14]), .QN( ));
Q_FDP1 \guid1_REG[13] ( .CK(clk), .R(rst_n), .D(nxt_guid1[13]), .Q(guid1[13]), .QN( ));
Q_FDP1 \guid1_REG[12] ( .CK(clk), .R(rst_n), .D(nxt_guid1[12]), .Q(guid1[12]), .QN( ));
Q_FDP1 \guid1_REG[11] ( .CK(clk), .R(rst_n), .D(nxt_guid1[11]), .Q(guid1[11]), .QN( ));
Q_FDP1 \guid1_REG[10] ( .CK(clk), .R(rst_n), .D(nxt_guid1[10]), .Q(guid1[10]), .QN( ));
Q_FDP1 \guid1_REG[9] ( .CK(clk), .R(rst_n), .D(nxt_guid1[9]), .Q(guid1[9]), .QN( ));
Q_FDP1 \guid1_REG[8] ( .CK(clk), .R(rst_n), .D(nxt_guid1[8]), .Q(guid1[8]), .QN( ));
Q_FDP1 \guid1_REG[7] ( .CK(clk), .R(rst_n), .D(nxt_guid1[7]), .Q(guid1[7]), .QN( ));
Q_FDP1 \guid1_REG[6] ( .CK(clk), .R(rst_n), .D(nxt_guid1[6]), .Q(guid1[6]), .QN( ));
Q_FDP1 \guid1_REG[5] ( .CK(clk), .R(rst_n), .D(nxt_guid1[5]), .Q(guid1[5]), .QN( ));
Q_FDP1 \guid1_REG[4] ( .CK(clk), .R(rst_n), .D(nxt_guid1[4]), .Q(guid1[4]), .QN( ));
Q_FDP1 \guid1_REG[3] ( .CK(clk), .R(rst_n), .D(nxt_guid1[3]), .Q(guid1[3]), .QN( ));
Q_FDP1 \guid1_REG[2] ( .CK(clk), .R(rst_n), .D(nxt_guid1[2]), .Q(guid1[2]), .QN( ));
Q_FDP1 \guid1_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_guid1[1]), .Q(guid1[1]), .QN( ));
Q_FDP1 \guid1_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_guid1[0]), .Q(guid1[0]), .QN( ));
Q_FDP1 \guid2_REG[63] ( .CK(clk), .R(rst_n), .D(nxt_guid2[63]), .Q(guid2[63]), .QN( ));
Q_FDP1 \guid2_REG[62] ( .CK(clk), .R(rst_n), .D(nxt_guid2[62]), .Q(guid2[62]), .QN( ));
Q_FDP1 \guid2_REG[61] ( .CK(clk), .R(rst_n), .D(nxt_guid2[61]), .Q(guid2[61]), .QN( ));
Q_FDP1 \guid2_REG[60] ( .CK(clk), .R(rst_n), .D(nxt_guid2[60]), .Q(guid2[60]), .QN( ));
Q_FDP1 \guid2_REG[59] ( .CK(clk), .R(rst_n), .D(nxt_guid2[59]), .Q(guid2[59]), .QN( ));
Q_FDP1 \guid2_REG[58] ( .CK(clk), .R(rst_n), .D(nxt_guid2[58]), .Q(guid2[58]), .QN( ));
Q_FDP1 \guid2_REG[57] ( .CK(clk), .R(rst_n), .D(nxt_guid2[57]), .Q(guid2[57]), .QN( ));
Q_FDP1 \guid2_REG[56] ( .CK(clk), .R(rst_n), .D(nxt_guid2[56]), .Q(guid2[56]), .QN( ));
Q_FDP1 \guid2_REG[55] ( .CK(clk), .R(rst_n), .D(nxt_guid2[55]), .Q(guid2[55]), .QN( ));
Q_FDP1 \guid2_REG[54] ( .CK(clk), .R(rst_n), .D(nxt_guid2[54]), .Q(guid2[54]), .QN( ));
Q_FDP1 \guid2_REG[53] ( .CK(clk), .R(rst_n), .D(nxt_guid2[53]), .Q(guid2[53]), .QN( ));
Q_FDP1 \guid2_REG[52] ( .CK(clk), .R(rst_n), .D(nxt_guid2[52]), .Q(guid2[52]), .QN( ));
Q_FDP1 \guid2_REG[51] ( .CK(clk), .R(rst_n), .D(nxt_guid2[51]), .Q(guid2[51]), .QN( ));
Q_FDP1 \guid2_REG[50] ( .CK(clk), .R(rst_n), .D(nxt_guid2[50]), .Q(guid2[50]), .QN( ));
Q_FDP1 \guid2_REG[49] ( .CK(clk), .R(rst_n), .D(nxt_guid2[49]), .Q(guid2[49]), .QN( ));
Q_FDP1 \guid2_REG[48] ( .CK(clk), .R(rst_n), .D(nxt_guid2[48]), .Q(guid2[48]), .QN( ));
Q_FDP1 \guid2_REG[47] ( .CK(clk), .R(rst_n), .D(nxt_guid2[47]), .Q(guid2[47]), .QN( ));
Q_FDP1 \guid2_REG[46] ( .CK(clk), .R(rst_n), .D(nxt_guid2[46]), .Q(guid2[46]), .QN( ));
Q_FDP1 \guid2_REG[45] ( .CK(clk), .R(rst_n), .D(nxt_guid2[45]), .Q(guid2[45]), .QN( ));
Q_FDP1 \guid2_REG[44] ( .CK(clk), .R(rst_n), .D(nxt_guid2[44]), .Q(guid2[44]), .QN( ));
Q_FDP1 \guid2_REG[43] ( .CK(clk), .R(rst_n), .D(nxt_guid2[43]), .Q(guid2[43]), .QN( ));
Q_FDP1 \guid2_REG[42] ( .CK(clk), .R(rst_n), .D(nxt_guid2[42]), .Q(guid2[42]), .QN( ));
Q_FDP1 \guid2_REG[41] ( .CK(clk), .R(rst_n), .D(nxt_guid2[41]), .Q(guid2[41]), .QN( ));
Q_FDP1 \guid2_REG[40] ( .CK(clk), .R(rst_n), .D(nxt_guid2[40]), .Q(guid2[40]), .QN( ));
Q_FDP1 \guid2_REG[39] ( .CK(clk), .R(rst_n), .D(nxt_guid2[39]), .Q(guid2[39]), .QN( ));
Q_FDP1 \guid2_REG[38] ( .CK(clk), .R(rst_n), .D(nxt_guid2[38]), .Q(guid2[38]), .QN( ));
Q_FDP1 \guid2_REG[37] ( .CK(clk), .R(rst_n), .D(nxt_guid2[37]), .Q(guid2[37]), .QN( ));
Q_FDP1 \guid2_REG[36] ( .CK(clk), .R(rst_n), .D(nxt_guid2[36]), .Q(guid2[36]), .QN( ));
Q_FDP1 \guid2_REG[35] ( .CK(clk), .R(rst_n), .D(nxt_guid2[35]), .Q(guid2[35]), .QN( ));
Q_FDP1 \guid2_REG[34] ( .CK(clk), .R(rst_n), .D(nxt_guid2[34]), .Q(guid2[34]), .QN( ));
Q_FDP1 \guid2_REG[33] ( .CK(clk), .R(rst_n), .D(nxt_guid2[33]), .Q(guid2[33]), .QN( ));
Q_FDP1 \guid2_REG[32] ( .CK(clk), .R(rst_n), .D(nxt_guid2[32]), .Q(guid2[32]), .QN( ));
Q_FDP1 \guid2_REG[31] ( .CK(clk), .R(rst_n), .D(nxt_guid2[31]), .Q(guid2[31]), .QN( ));
Q_FDP1 \guid2_REG[30] ( .CK(clk), .R(rst_n), .D(nxt_guid2[30]), .Q(guid2[30]), .QN( ));
Q_FDP1 \guid2_REG[29] ( .CK(clk), .R(rst_n), .D(nxt_guid2[29]), .Q(guid2[29]), .QN( ));
Q_FDP1 \guid2_REG[28] ( .CK(clk), .R(rst_n), .D(nxt_guid2[28]), .Q(guid2[28]), .QN( ));
Q_FDP1 \guid2_REG[27] ( .CK(clk), .R(rst_n), .D(nxt_guid2[27]), .Q(guid2[27]), .QN( ));
Q_FDP1 \guid2_REG[26] ( .CK(clk), .R(rst_n), .D(nxt_guid2[26]), .Q(guid2[26]), .QN( ));
Q_FDP1 \guid2_REG[25] ( .CK(clk), .R(rst_n), .D(nxt_guid2[25]), .Q(guid2[25]), .QN( ));
Q_FDP1 \guid2_REG[24] ( .CK(clk), .R(rst_n), .D(nxt_guid2[24]), .Q(guid2[24]), .QN( ));
Q_FDP1 \guid2_REG[23] ( .CK(clk), .R(rst_n), .D(nxt_guid2[23]), .Q(guid2[23]), .QN( ));
Q_FDP1 \guid2_REG[22] ( .CK(clk), .R(rst_n), .D(nxt_guid2[22]), .Q(guid2[22]), .QN( ));
Q_FDP1 \guid2_REG[21] ( .CK(clk), .R(rst_n), .D(nxt_guid2[21]), .Q(guid2[21]), .QN( ));
Q_FDP1 \guid2_REG[20] ( .CK(clk), .R(rst_n), .D(nxt_guid2[20]), .Q(guid2[20]), .QN( ));
Q_FDP1 \guid2_REG[19] ( .CK(clk), .R(rst_n), .D(nxt_guid2[19]), .Q(guid2[19]), .QN( ));
Q_FDP1 \guid2_REG[18] ( .CK(clk), .R(rst_n), .D(nxt_guid2[18]), .Q(guid2[18]), .QN( ));
Q_FDP1 \guid2_REG[17] ( .CK(clk), .R(rst_n), .D(nxt_guid2[17]), .Q(guid2[17]), .QN( ));
Q_FDP1 \guid2_REG[16] ( .CK(clk), .R(rst_n), .D(nxt_guid2[16]), .Q(guid2[16]), .QN( ));
Q_FDP1 \guid2_REG[15] ( .CK(clk), .R(rst_n), .D(nxt_guid2[15]), .Q(guid2[15]), .QN( ));
Q_FDP1 \guid2_REG[14] ( .CK(clk), .R(rst_n), .D(nxt_guid2[14]), .Q(guid2[14]), .QN( ));
Q_FDP1 \guid2_REG[13] ( .CK(clk), .R(rst_n), .D(nxt_guid2[13]), .Q(guid2[13]), .QN( ));
Q_FDP1 \guid2_REG[12] ( .CK(clk), .R(rst_n), .D(nxt_guid2[12]), .Q(guid2[12]), .QN( ));
Q_FDP1 \guid2_REG[11] ( .CK(clk), .R(rst_n), .D(nxt_guid2[11]), .Q(guid2[11]), .QN( ));
Q_FDP1 \guid2_REG[10] ( .CK(clk), .R(rst_n), .D(nxt_guid2[10]), .Q(guid2[10]), .QN( ));
Q_FDP1 \guid2_REG[9] ( .CK(clk), .R(rst_n), .D(nxt_guid2[9]), .Q(guid2[9]), .QN( ));
Q_FDP1 \guid2_REG[8] ( .CK(clk), .R(rst_n), .D(nxt_guid2[8]), .Q(guid2[8]), .QN( ));
Q_FDP1 \guid2_REG[7] ( .CK(clk), .R(rst_n), .D(nxt_guid2[7]), .Q(guid2[7]), .QN( ));
Q_FDP1 \guid2_REG[6] ( .CK(clk), .R(rst_n), .D(nxt_guid2[6]), .Q(guid2[6]), .QN( ));
Q_FDP1 \guid2_REG[5] ( .CK(clk), .R(rst_n), .D(nxt_guid2[5]), .Q(guid2[5]), .QN( ));
Q_FDP1 \guid2_REG[4] ( .CK(clk), .R(rst_n), .D(nxt_guid2[4]), .Q(guid2[4]), .QN( ));
Q_FDP1 \guid2_REG[3] ( .CK(clk), .R(rst_n), .D(nxt_guid2[3]), .Q(guid2[3]), .QN( ));
Q_FDP1 \guid2_REG[2] ( .CK(clk), .R(rst_n), .D(nxt_guid2[2]), .Q(guid2[2]), .QN( ));
Q_FDP1 \guid2_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_guid2[1]), .Q(guid2[1]), .QN( ));
Q_FDP1 \guid2_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_guid2[0]), .Q(guid2[0]), .QN( ));
Q_FDP1 \guid3_REG[63] ( .CK(clk), .R(rst_n), .D(nxt_guid3[63]), .Q(guid3[63]), .QN( ));
Q_FDP1 \guid3_REG[62] ( .CK(clk), .R(rst_n), .D(nxt_guid3[62]), .Q(guid3[62]), .QN( ));
Q_FDP1 \guid3_REG[61] ( .CK(clk), .R(rst_n), .D(nxt_guid3[61]), .Q(guid3[61]), .QN( ));
Q_FDP1 \guid3_REG[60] ( .CK(clk), .R(rst_n), .D(nxt_guid3[60]), .Q(guid3[60]), .QN( ));
Q_FDP1 \guid3_REG[59] ( .CK(clk), .R(rst_n), .D(nxt_guid3[59]), .Q(guid3[59]), .QN( ));
Q_FDP1 \guid3_REG[58] ( .CK(clk), .R(rst_n), .D(nxt_guid3[58]), .Q(guid3[58]), .QN( ));
Q_FDP1 \guid3_REG[57] ( .CK(clk), .R(rst_n), .D(nxt_guid3[57]), .Q(guid3[57]), .QN( ));
Q_FDP1 \guid3_REG[56] ( .CK(clk), .R(rst_n), .D(nxt_guid3[56]), .Q(guid3[56]), .QN( ));
Q_FDP1 \guid3_REG[55] ( .CK(clk), .R(rst_n), .D(nxt_guid3[55]), .Q(guid3[55]), .QN( ));
Q_FDP1 \guid3_REG[54] ( .CK(clk), .R(rst_n), .D(nxt_guid3[54]), .Q(guid3[54]), .QN( ));
Q_FDP1 \guid3_REG[53] ( .CK(clk), .R(rst_n), .D(nxt_guid3[53]), .Q(guid3[53]), .QN( ));
Q_FDP1 \guid3_REG[52] ( .CK(clk), .R(rst_n), .D(nxt_guid3[52]), .Q(guid3[52]), .QN( ));
Q_FDP1 \guid3_REG[51] ( .CK(clk), .R(rst_n), .D(nxt_guid3[51]), .Q(guid3[51]), .QN( ));
Q_FDP1 \guid3_REG[50] ( .CK(clk), .R(rst_n), .D(nxt_guid3[50]), .Q(guid3[50]), .QN( ));
Q_FDP1 \guid3_REG[49] ( .CK(clk), .R(rst_n), .D(nxt_guid3[49]), .Q(guid3[49]), .QN( ));
Q_FDP1 \guid3_REG[48] ( .CK(clk), .R(rst_n), .D(nxt_guid3[48]), .Q(guid3[48]), .QN( ));
Q_FDP1 \guid3_REG[47] ( .CK(clk), .R(rst_n), .D(nxt_guid3[47]), .Q(guid3[47]), .QN( ));
Q_FDP1 \guid3_REG[46] ( .CK(clk), .R(rst_n), .D(nxt_guid3[46]), .Q(guid3[46]), .QN( ));
Q_FDP1 \guid3_REG[45] ( .CK(clk), .R(rst_n), .D(nxt_guid3[45]), .Q(guid3[45]), .QN( ));
Q_FDP1 \guid3_REG[44] ( .CK(clk), .R(rst_n), .D(nxt_guid3[44]), .Q(guid3[44]), .QN( ));
Q_FDP1 \guid3_REG[43] ( .CK(clk), .R(rst_n), .D(nxt_guid3[43]), .Q(guid3[43]), .QN( ));
Q_FDP1 \guid3_REG[42] ( .CK(clk), .R(rst_n), .D(nxt_guid3[42]), .Q(guid3[42]), .QN( ));
Q_FDP1 \guid3_REG[41] ( .CK(clk), .R(rst_n), .D(nxt_guid3[41]), .Q(guid3[41]), .QN( ));
Q_FDP1 \guid3_REG[40] ( .CK(clk), .R(rst_n), .D(nxt_guid3[40]), .Q(guid3[40]), .QN( ));
Q_FDP1 \guid3_REG[39] ( .CK(clk), .R(rst_n), .D(nxt_guid3[39]), .Q(guid3[39]), .QN( ));
Q_FDP1 \guid3_REG[38] ( .CK(clk), .R(rst_n), .D(nxt_guid3[38]), .Q(guid3[38]), .QN( ));
Q_FDP1 \guid3_REG[37] ( .CK(clk), .R(rst_n), .D(nxt_guid3[37]), .Q(guid3[37]), .QN( ));
Q_FDP1 \guid3_REG[36] ( .CK(clk), .R(rst_n), .D(nxt_guid3[36]), .Q(guid3[36]), .QN( ));
Q_FDP1 \guid3_REG[35] ( .CK(clk), .R(rst_n), .D(nxt_guid3[35]), .Q(guid3[35]), .QN( ));
Q_FDP1 \guid3_REG[34] ( .CK(clk), .R(rst_n), .D(nxt_guid3[34]), .Q(guid3[34]), .QN( ));
Q_FDP1 \guid3_REG[33] ( .CK(clk), .R(rst_n), .D(nxt_guid3[33]), .Q(guid3[33]), .QN( ));
Q_FDP1 \guid3_REG[32] ( .CK(clk), .R(rst_n), .D(nxt_guid3[32]), .Q(guid3[32]), .QN( ));
Q_FDP1 \guid3_REG[31] ( .CK(clk), .R(rst_n), .D(nxt_guid3[31]), .Q(guid3[31]), .QN( ));
Q_FDP1 \guid3_REG[30] ( .CK(clk), .R(rst_n), .D(nxt_guid3[30]), .Q(guid3[30]), .QN( ));
Q_FDP1 \guid3_REG[29] ( .CK(clk), .R(rst_n), .D(nxt_guid3[29]), .Q(guid3[29]), .QN( ));
Q_FDP1 \guid3_REG[28] ( .CK(clk), .R(rst_n), .D(nxt_guid3[28]), .Q(guid3[28]), .QN( ));
Q_FDP1 \guid3_REG[27] ( .CK(clk), .R(rst_n), .D(nxt_guid3[27]), .Q(guid3[27]), .QN( ));
Q_FDP1 \guid3_REG[26] ( .CK(clk), .R(rst_n), .D(nxt_guid3[26]), .Q(guid3[26]), .QN( ));
Q_FDP1 \guid3_REG[25] ( .CK(clk), .R(rst_n), .D(nxt_guid3[25]), .Q(guid3[25]), .QN( ));
Q_FDP1 \guid3_REG[24] ( .CK(clk), .R(rst_n), .D(nxt_guid3[24]), .Q(guid3[24]), .QN( ));
Q_FDP1 \guid3_REG[23] ( .CK(clk), .R(rst_n), .D(nxt_guid3[23]), .Q(guid3[23]), .QN( ));
Q_FDP1 \guid3_REG[22] ( .CK(clk), .R(rst_n), .D(nxt_guid3[22]), .Q(guid3[22]), .QN( ));
Q_FDP1 \guid3_REG[21] ( .CK(clk), .R(rst_n), .D(nxt_guid3[21]), .Q(guid3[21]), .QN( ));
Q_FDP1 \guid3_REG[20] ( .CK(clk), .R(rst_n), .D(nxt_guid3[20]), .Q(guid3[20]), .QN( ));
Q_FDP1 \guid3_REG[19] ( .CK(clk), .R(rst_n), .D(nxt_guid3[19]), .Q(guid3[19]), .QN( ));
Q_FDP1 \guid3_REG[18] ( .CK(clk), .R(rst_n), .D(nxt_guid3[18]), .Q(guid3[18]), .QN( ));
Q_FDP1 \guid3_REG[17] ( .CK(clk), .R(rst_n), .D(nxt_guid3[17]), .Q(guid3[17]), .QN( ));
Q_FDP1 \guid3_REG[16] ( .CK(clk), .R(rst_n), .D(nxt_guid3[16]), .Q(guid3[16]), .QN( ));
Q_FDP1 \guid3_REG[15] ( .CK(clk), .R(rst_n), .D(nxt_guid3[15]), .Q(guid3[15]), .QN( ));
Q_FDP1 \guid3_REG[14] ( .CK(clk), .R(rst_n), .D(nxt_guid3[14]), .Q(guid3[14]), .QN( ));
Q_FDP1 \guid3_REG[13] ( .CK(clk), .R(rst_n), .D(nxt_guid3[13]), .Q(guid3[13]), .QN( ));
Q_FDP1 \guid3_REG[12] ( .CK(clk), .R(rst_n), .D(nxt_guid3[12]), .Q(guid3[12]), .QN( ));
Q_FDP1 \guid3_REG[11] ( .CK(clk), .R(rst_n), .D(nxt_guid3[11]), .Q(guid3[11]), .QN( ));
Q_FDP1 \guid3_REG[10] ( .CK(clk), .R(rst_n), .D(nxt_guid3[10]), .Q(guid3[10]), .QN( ));
Q_FDP1 \guid3_REG[9] ( .CK(clk), .R(rst_n), .D(nxt_guid3[9]), .Q(guid3[9]), .QN( ));
Q_FDP1 \guid3_REG[8] ( .CK(clk), .R(rst_n), .D(nxt_guid3[8]), .Q(guid3[8]), .QN( ));
Q_FDP1 \guid3_REG[7] ( .CK(clk), .R(rst_n), .D(nxt_guid3[7]), .Q(guid3[7]), .QN( ));
Q_FDP1 \guid3_REG[6] ( .CK(clk), .R(rst_n), .D(nxt_guid3[6]), .Q(guid3[6]), .QN( ));
Q_FDP1 \guid3_REG[5] ( .CK(clk), .R(rst_n), .D(nxt_guid3[5]), .Q(guid3[5]), .QN( ));
Q_FDP1 \guid3_REG[4] ( .CK(clk), .R(rst_n), .D(nxt_guid3[4]), .Q(guid3[4]), .QN( ));
Q_FDP1 \guid3_REG[3] ( .CK(clk), .R(rst_n), .D(nxt_guid3[3]), .Q(guid3[3]), .QN( ));
Q_FDP1 \guid3_REG[2] ( .CK(clk), .R(rst_n), .D(nxt_guid3[2]), .Q(guid3[2]), .QN( ));
Q_FDP1 \guid3_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_guid3[1]), .Q(guid3[1]), .QN( ));
Q_FDP1 \guid3_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_guid3[0]), .Q(guid3[0]), .QN( ));
Q_FDP1 \iv0_REG[63] ( .CK(clk), .R(rst_n), .D(nxt_iv0[63]), .Q(iv0[63]), .QN( ));
Q_FDP1 \iv0_REG[62] ( .CK(clk), .R(rst_n), .D(nxt_iv0[62]), .Q(iv0[62]), .QN( ));
Q_FDP1 \iv0_REG[61] ( .CK(clk), .R(rst_n), .D(nxt_iv0[61]), .Q(iv0[61]), .QN( ));
Q_FDP1 \iv0_REG[60] ( .CK(clk), .R(rst_n), .D(nxt_iv0[60]), .Q(iv0[60]), .QN( ));
Q_FDP1 \iv0_REG[59] ( .CK(clk), .R(rst_n), .D(nxt_iv0[59]), .Q(iv0[59]), .QN( ));
Q_FDP1 \iv0_REG[58] ( .CK(clk), .R(rst_n), .D(nxt_iv0[58]), .Q(iv0[58]), .QN( ));
Q_FDP1 \iv0_REG[57] ( .CK(clk), .R(rst_n), .D(nxt_iv0[57]), .Q(iv0[57]), .QN( ));
Q_FDP1 \iv0_REG[56] ( .CK(clk), .R(rst_n), .D(nxt_iv0[56]), .Q(iv0[56]), .QN( ));
Q_FDP1 \iv0_REG[55] ( .CK(clk), .R(rst_n), .D(nxt_iv0[55]), .Q(iv0[55]), .QN( ));
Q_FDP1 \iv0_REG[54] ( .CK(clk), .R(rst_n), .D(nxt_iv0[54]), .Q(iv0[54]), .QN( ));
Q_FDP1 \iv0_REG[53] ( .CK(clk), .R(rst_n), .D(nxt_iv0[53]), .Q(iv0[53]), .QN( ));
Q_FDP1 \iv0_REG[52] ( .CK(clk), .R(rst_n), .D(nxt_iv0[52]), .Q(iv0[52]), .QN( ));
Q_FDP1 \iv0_REG[51] ( .CK(clk), .R(rst_n), .D(nxt_iv0[51]), .Q(iv0[51]), .QN( ));
Q_FDP1 \iv0_REG[50] ( .CK(clk), .R(rst_n), .D(nxt_iv0[50]), .Q(iv0[50]), .QN( ));
Q_FDP1 \iv0_REG[49] ( .CK(clk), .R(rst_n), .D(nxt_iv0[49]), .Q(iv0[49]), .QN( ));
Q_FDP1 \iv0_REG[48] ( .CK(clk), .R(rst_n), .D(nxt_iv0[48]), .Q(iv0[48]), .QN( ));
Q_FDP1 \iv0_REG[47] ( .CK(clk), .R(rst_n), .D(nxt_iv0[47]), .Q(iv0[47]), .QN( ));
Q_FDP1 \iv0_REG[46] ( .CK(clk), .R(rst_n), .D(nxt_iv0[46]), .Q(iv0[46]), .QN( ));
Q_FDP1 \iv0_REG[45] ( .CK(clk), .R(rst_n), .D(nxt_iv0[45]), .Q(iv0[45]), .QN( ));
Q_FDP1 \iv0_REG[44] ( .CK(clk), .R(rst_n), .D(nxt_iv0[44]), .Q(iv0[44]), .QN( ));
Q_FDP1 \iv0_REG[43] ( .CK(clk), .R(rst_n), .D(nxt_iv0[43]), .Q(iv0[43]), .QN( ));
Q_FDP1 \iv0_REG[42] ( .CK(clk), .R(rst_n), .D(nxt_iv0[42]), .Q(iv0[42]), .QN( ));
Q_FDP1 \iv0_REG[41] ( .CK(clk), .R(rst_n), .D(nxt_iv0[41]), .Q(iv0[41]), .QN( ));
Q_FDP1 \iv0_REG[40] ( .CK(clk), .R(rst_n), .D(nxt_iv0[40]), .Q(iv0[40]), .QN( ));
Q_FDP1 \iv0_REG[39] ( .CK(clk), .R(rst_n), .D(nxt_iv0[39]), .Q(iv0[39]), .QN( ));
Q_FDP1 \iv0_REG[38] ( .CK(clk), .R(rst_n), .D(nxt_iv0[38]), .Q(iv0[38]), .QN( ));
Q_FDP1 \iv0_REG[37] ( .CK(clk), .R(rst_n), .D(nxt_iv0[37]), .Q(iv0[37]), .QN( ));
Q_FDP1 \iv0_REG[36] ( .CK(clk), .R(rst_n), .D(nxt_iv0[36]), .Q(iv0[36]), .QN( ));
Q_FDP1 \iv0_REG[35] ( .CK(clk), .R(rst_n), .D(nxt_iv0[35]), .Q(iv0[35]), .QN( ));
Q_FDP1 \iv0_REG[34] ( .CK(clk), .R(rst_n), .D(nxt_iv0[34]), .Q(iv0[34]), .QN( ));
Q_FDP1 \iv0_REG[33] ( .CK(clk), .R(rst_n), .D(nxt_iv0[33]), .Q(iv0[33]), .QN( ));
Q_FDP1 \iv0_REG[32] ( .CK(clk), .R(rst_n), .D(nxt_iv0[32]), .Q(iv0[32]), .QN( ));
Q_FDP1 \iv0_REG[31] ( .CK(clk), .R(rst_n), .D(nxt_iv0[31]), .Q(iv0[31]), .QN( ));
Q_FDP1 \iv0_REG[30] ( .CK(clk), .R(rst_n), .D(nxt_iv0[30]), .Q(iv0[30]), .QN( ));
Q_FDP1 \iv0_REG[29] ( .CK(clk), .R(rst_n), .D(nxt_iv0[29]), .Q(iv0[29]), .QN( ));
Q_FDP1 \iv0_REG[28] ( .CK(clk), .R(rst_n), .D(nxt_iv0[28]), .Q(iv0[28]), .QN( ));
Q_FDP1 \iv0_REG[27] ( .CK(clk), .R(rst_n), .D(nxt_iv0[27]), .Q(iv0[27]), .QN( ));
Q_FDP1 \iv0_REG[26] ( .CK(clk), .R(rst_n), .D(nxt_iv0[26]), .Q(iv0[26]), .QN( ));
Q_FDP1 \iv0_REG[25] ( .CK(clk), .R(rst_n), .D(nxt_iv0[25]), .Q(iv0[25]), .QN( ));
Q_FDP1 \iv0_REG[24] ( .CK(clk), .R(rst_n), .D(nxt_iv0[24]), .Q(iv0[24]), .QN( ));
Q_FDP1 \iv0_REG[23] ( .CK(clk), .R(rst_n), .D(nxt_iv0[23]), .Q(iv0[23]), .QN( ));
Q_FDP1 \iv0_REG[22] ( .CK(clk), .R(rst_n), .D(nxt_iv0[22]), .Q(iv0[22]), .QN( ));
Q_FDP1 \iv0_REG[21] ( .CK(clk), .R(rst_n), .D(nxt_iv0[21]), .Q(iv0[21]), .QN( ));
Q_FDP1 \iv0_REG[20] ( .CK(clk), .R(rst_n), .D(nxt_iv0[20]), .Q(iv0[20]), .QN( ));
Q_FDP1 \iv0_REG[19] ( .CK(clk), .R(rst_n), .D(nxt_iv0[19]), .Q(iv0[19]), .QN( ));
Q_FDP1 \iv0_REG[18] ( .CK(clk), .R(rst_n), .D(nxt_iv0[18]), .Q(iv0[18]), .QN( ));
Q_FDP1 \iv0_REG[17] ( .CK(clk), .R(rst_n), .D(nxt_iv0[17]), .Q(iv0[17]), .QN( ));
Q_FDP1 \iv0_REG[16] ( .CK(clk), .R(rst_n), .D(nxt_iv0[16]), .Q(iv0[16]), .QN( ));
Q_FDP1 \iv0_REG[15] ( .CK(clk), .R(rst_n), .D(nxt_iv0[15]), .Q(iv0[15]), .QN( ));
Q_FDP1 \iv0_REG[14] ( .CK(clk), .R(rst_n), .D(nxt_iv0[14]), .Q(iv0[14]), .QN( ));
Q_FDP1 \iv0_REG[13] ( .CK(clk), .R(rst_n), .D(nxt_iv0[13]), .Q(iv0[13]), .QN( ));
Q_FDP1 \iv0_REG[12] ( .CK(clk), .R(rst_n), .D(nxt_iv0[12]), .Q(iv0[12]), .QN( ));
Q_FDP1 \iv0_REG[11] ( .CK(clk), .R(rst_n), .D(nxt_iv0[11]), .Q(iv0[11]), .QN( ));
Q_FDP1 \iv0_REG[10] ( .CK(clk), .R(rst_n), .D(nxt_iv0[10]), .Q(iv0[10]), .QN( ));
Q_FDP1 \iv0_REG[9] ( .CK(clk), .R(rst_n), .D(nxt_iv0[9]), .Q(iv0[9]), .QN( ));
Q_FDP1 \iv0_REG[8] ( .CK(clk), .R(rst_n), .D(nxt_iv0[8]), .Q(iv0[8]), .QN( ));
Q_FDP1 \iv0_REG[7] ( .CK(clk), .R(rst_n), .D(nxt_iv0[7]), .Q(iv0[7]), .QN( ));
Q_FDP1 \iv0_REG[6] ( .CK(clk), .R(rst_n), .D(nxt_iv0[6]), .Q(iv0[6]), .QN( ));
Q_FDP1 \iv0_REG[5] ( .CK(clk), .R(rst_n), .D(nxt_iv0[5]), .Q(iv0[5]), .QN( ));
Q_FDP1 \iv0_REG[4] ( .CK(clk), .R(rst_n), .D(nxt_iv0[4]), .Q(iv0[4]), .QN( ));
Q_FDP1 \iv0_REG[3] ( .CK(clk), .R(rst_n), .D(nxt_iv0[3]), .Q(iv0[3]), .QN( ));
Q_FDP1 \iv0_REG[2] ( .CK(clk), .R(rst_n), .D(nxt_iv0[2]), .Q(iv0[2]), .QN( ));
Q_FDP1 \iv0_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_iv0[1]), .Q(iv0[1]), .QN( ));
Q_FDP1 \iv0_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_iv0[0]), .Q(iv0[0]), .QN( ));
Q_FDP1 \iv1_REG[63] ( .CK(clk), .R(rst_n), .D(nxt_iv1[63]), .Q(iv1[63]), .QN( ));
Q_FDP1 \iv1_REG[62] ( .CK(clk), .R(rst_n), .D(nxt_iv1[62]), .Q(iv1[62]), .QN( ));
Q_FDP1 \iv1_REG[61] ( .CK(clk), .R(rst_n), .D(nxt_iv1[61]), .Q(iv1[61]), .QN( ));
Q_FDP1 \iv1_REG[60] ( .CK(clk), .R(rst_n), .D(nxt_iv1[60]), .Q(iv1[60]), .QN( ));
Q_FDP1 \iv1_REG[59] ( .CK(clk), .R(rst_n), .D(nxt_iv1[59]), .Q(iv1[59]), .QN( ));
Q_FDP1 \iv1_REG[58] ( .CK(clk), .R(rst_n), .D(nxt_iv1[58]), .Q(iv1[58]), .QN( ));
Q_FDP1 \iv1_REG[57] ( .CK(clk), .R(rst_n), .D(nxt_iv1[57]), .Q(iv1[57]), .QN( ));
Q_FDP1 \iv1_REG[56] ( .CK(clk), .R(rst_n), .D(nxt_iv1[56]), .Q(iv1[56]), .QN( ));
Q_FDP1 \iv1_REG[55] ( .CK(clk), .R(rst_n), .D(nxt_iv1[55]), .Q(iv1[55]), .QN( ));
Q_FDP1 \iv1_REG[54] ( .CK(clk), .R(rst_n), .D(nxt_iv1[54]), .Q(iv1[54]), .QN( ));
Q_FDP1 \iv1_REG[53] ( .CK(clk), .R(rst_n), .D(nxt_iv1[53]), .Q(iv1[53]), .QN( ));
Q_FDP1 \iv1_REG[52] ( .CK(clk), .R(rst_n), .D(nxt_iv1[52]), .Q(iv1[52]), .QN( ));
Q_FDP1 \iv1_REG[51] ( .CK(clk), .R(rst_n), .D(nxt_iv1[51]), .Q(iv1[51]), .QN( ));
Q_FDP1 \iv1_REG[50] ( .CK(clk), .R(rst_n), .D(nxt_iv1[50]), .Q(iv1[50]), .QN( ));
Q_FDP1 \iv1_REG[49] ( .CK(clk), .R(rst_n), .D(nxt_iv1[49]), .Q(iv1[49]), .QN( ));
Q_FDP1 \iv1_REG[48] ( .CK(clk), .R(rst_n), .D(nxt_iv1[48]), .Q(iv1[48]), .QN( ));
Q_FDP1 \iv1_REG[47] ( .CK(clk), .R(rst_n), .D(nxt_iv1[47]), .Q(iv1[47]), .QN( ));
Q_FDP1 \iv1_REG[46] ( .CK(clk), .R(rst_n), .D(nxt_iv1[46]), .Q(iv1[46]), .QN( ));
Q_FDP1 \iv1_REG[45] ( .CK(clk), .R(rst_n), .D(nxt_iv1[45]), .Q(iv1[45]), .QN( ));
Q_FDP1 \iv1_REG[44] ( .CK(clk), .R(rst_n), .D(nxt_iv1[44]), .Q(iv1[44]), .QN( ));
Q_FDP1 \iv1_REG[43] ( .CK(clk), .R(rst_n), .D(nxt_iv1[43]), .Q(iv1[43]), .QN( ));
Q_FDP1 \iv1_REG[42] ( .CK(clk), .R(rst_n), .D(nxt_iv1[42]), .Q(iv1[42]), .QN( ));
Q_FDP1 \iv1_REG[41] ( .CK(clk), .R(rst_n), .D(nxt_iv1[41]), .Q(iv1[41]), .QN( ));
Q_FDP1 \iv1_REG[40] ( .CK(clk), .R(rst_n), .D(nxt_iv1[40]), .Q(iv1[40]), .QN( ));
Q_FDP1 \iv1_REG[39] ( .CK(clk), .R(rst_n), .D(nxt_iv1[39]), .Q(iv1[39]), .QN( ));
Q_FDP1 \iv1_REG[38] ( .CK(clk), .R(rst_n), .D(nxt_iv1[38]), .Q(iv1[38]), .QN( ));
Q_FDP1 \iv1_REG[37] ( .CK(clk), .R(rst_n), .D(nxt_iv1[37]), .Q(iv1[37]), .QN( ));
Q_FDP1 \iv1_REG[36] ( .CK(clk), .R(rst_n), .D(nxt_iv1[36]), .Q(iv1[36]), .QN( ));
Q_FDP1 \iv1_REG[35] ( .CK(clk), .R(rst_n), .D(nxt_iv1[35]), .Q(iv1[35]), .QN( ));
Q_FDP1 \iv1_REG[34] ( .CK(clk), .R(rst_n), .D(nxt_iv1[34]), .Q(iv1[34]), .QN( ));
Q_FDP1 \iv1_REG[33] ( .CK(clk), .R(rst_n), .D(nxt_iv1[33]), .Q(iv1[33]), .QN( ));
Q_FDP1 \iv1_REG[32] ( .CK(clk), .R(rst_n), .D(nxt_iv1[32]), .Q(iv1[32]), .QN( ));
Q_FDP1 \iv1_REG[31] ( .CK(clk), .R(rst_n), .D(nxt_iv1[31]), .Q(iv1[31]), .QN( ));
Q_FDP1 \iv1_REG[30] ( .CK(clk), .R(rst_n), .D(nxt_iv1[30]), .Q(iv1[30]), .QN( ));
Q_FDP1 \iv1_REG[29] ( .CK(clk), .R(rst_n), .D(nxt_iv1[29]), .Q(iv1[29]), .QN( ));
Q_FDP1 \iv1_REG[28] ( .CK(clk), .R(rst_n), .D(nxt_iv1[28]), .Q(iv1[28]), .QN( ));
Q_FDP1 \iv1_REG[27] ( .CK(clk), .R(rst_n), .D(nxt_iv1[27]), .Q(iv1[27]), .QN( ));
Q_FDP1 \iv1_REG[26] ( .CK(clk), .R(rst_n), .D(nxt_iv1[26]), .Q(iv1[26]), .QN( ));
Q_FDP1 \iv1_REG[25] ( .CK(clk), .R(rst_n), .D(nxt_iv1[25]), .Q(iv1[25]), .QN( ));
Q_FDP1 \iv1_REG[24] ( .CK(clk), .R(rst_n), .D(nxt_iv1[24]), .Q(iv1[24]), .QN( ));
Q_FDP1 \iv1_REG[23] ( .CK(clk), .R(rst_n), .D(nxt_iv1[23]), .Q(iv1[23]), .QN( ));
Q_FDP1 \iv1_REG[22] ( .CK(clk), .R(rst_n), .D(nxt_iv1[22]), .Q(iv1[22]), .QN( ));
Q_FDP1 \iv1_REG[21] ( .CK(clk), .R(rst_n), .D(nxt_iv1[21]), .Q(iv1[21]), .QN( ));
Q_FDP1 \iv1_REG[20] ( .CK(clk), .R(rst_n), .D(nxt_iv1[20]), .Q(iv1[20]), .QN( ));
Q_FDP1 \iv1_REG[19] ( .CK(clk), .R(rst_n), .D(nxt_iv1[19]), .Q(iv1[19]), .QN( ));
Q_FDP1 \iv1_REG[18] ( .CK(clk), .R(rst_n), .D(nxt_iv1[18]), .Q(iv1[18]), .QN( ));
Q_FDP1 \iv1_REG[17] ( .CK(clk), .R(rst_n), .D(nxt_iv1[17]), .Q(iv1[17]), .QN( ));
Q_FDP1 \iv1_REG[16] ( .CK(clk), .R(rst_n), .D(nxt_iv1[16]), .Q(iv1[16]), .QN( ));
Q_FDP1 \iv1_REG[15] ( .CK(clk), .R(rst_n), .D(nxt_iv1[15]), .Q(iv1[15]), .QN( ));
Q_FDP1 \iv1_REG[14] ( .CK(clk), .R(rst_n), .D(nxt_iv1[14]), .Q(iv1[14]), .QN( ));
Q_FDP1 \iv1_REG[13] ( .CK(clk), .R(rst_n), .D(nxt_iv1[13]), .Q(iv1[13]), .QN( ));
Q_FDP1 \iv1_REG[12] ( .CK(clk), .R(rst_n), .D(nxt_iv1[12]), .Q(iv1[12]), .QN( ));
Q_FDP1 \iv1_REG[11] ( .CK(clk), .R(rst_n), .D(nxt_iv1[11]), .Q(iv1[11]), .QN( ));
Q_FDP1 \iv1_REG[10] ( .CK(clk), .R(rst_n), .D(nxt_iv1[10]), .Q(iv1[10]), .QN( ));
Q_FDP1 \iv1_REG[9] ( .CK(clk), .R(rst_n), .D(nxt_iv1[9]), .Q(iv1[9]), .QN( ));
Q_FDP1 \iv1_REG[8] ( .CK(clk), .R(rst_n), .D(nxt_iv1[8]), .Q(iv1[8]), .QN( ));
Q_FDP1 \iv1_REG[7] ( .CK(clk), .R(rst_n), .D(nxt_iv1[7]), .Q(iv1[7]), .QN( ));
Q_FDP1 \iv1_REG[6] ( .CK(clk), .R(rst_n), .D(nxt_iv1[6]), .Q(iv1[6]), .QN( ));
Q_FDP1 \iv1_REG[5] ( .CK(clk), .R(rst_n), .D(nxt_iv1[5]), .Q(iv1[5]), .QN( ));
Q_FDP1 \iv1_REG[4] ( .CK(clk), .R(rst_n), .D(nxt_iv1[4]), .Q(iv1[4]), .QN( ));
Q_FDP1 \iv1_REG[3] ( .CK(clk), .R(rst_n), .D(nxt_iv1[3]), .Q(iv1[3]), .QN( ));
Q_FDP1 \iv1_REG[2] ( .CK(clk), .R(rst_n), .D(nxt_iv1[2]), .Q(iv1[2]), .QN( ));
Q_FDP1 \iv1_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_iv1[1]), .Q(iv1[1]), .QN( ));
Q_FDP1 \iv1_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_iv1[0]), .Q(iv1[0]), .QN( ));
Q_FDP1 \buffer_REG[31] ( .CK(clk), .R(rst_n), .D(nxt_buffer[31]), .Q(buffer[31]), .QN( ));
Q_FDP1 \buffer_REG[30] ( .CK(clk), .R(rst_n), .D(nxt_buffer[30]), .Q(buffer[30]), .QN( ));
Q_FDP1 \buffer_REG[29] ( .CK(clk), .R(rst_n), .D(nxt_buffer[29]), .Q(buffer[29]), .QN( ));
Q_FDP1 \buffer_REG[28] ( .CK(clk), .R(rst_n), .D(nxt_buffer[28]), .Q(buffer[28]), .QN( ));
Q_FDP1 \buffer_REG[27] ( .CK(clk), .R(rst_n), .D(nxt_buffer[27]), .Q(buffer[27]), .QN( ));
Q_FDP1 \buffer_REG[26] ( .CK(clk), .R(rst_n), .D(nxt_buffer[26]), .Q(buffer[26]), .QN( ));
Q_FDP1 \buffer_REG[25] ( .CK(clk), .R(rst_n), .D(nxt_buffer[25]), .Q(buffer[25]), .QN( ));
Q_FDP1 \buffer_REG[24] ( .CK(clk), .R(rst_n), .D(nxt_buffer[24]), .Q(buffer[24]), .QN( ));
Q_FDP1 \buffer_REG[23] ( .CK(clk), .R(rst_n), .D(nxt_buffer[23]), .Q(buffer[23]), .QN( ));
Q_FDP1 \buffer_REG[22] ( .CK(clk), .R(rst_n), .D(nxt_buffer[22]), .Q(buffer[22]), .QN( ));
Q_FDP1 \buffer_REG[21] ( .CK(clk), .R(rst_n), .D(nxt_buffer[21]), .Q(buffer[21]), .QN( ));
Q_FDP1 \buffer_REG[20] ( .CK(clk), .R(rst_n), .D(nxt_buffer[20]), .Q(buffer[20]), .QN( ));
Q_FDP1 \buffer_REG[19] ( .CK(clk), .R(rst_n), .D(nxt_buffer[19]), .Q(buffer[19]), .QN( ));
Q_FDP1 \buffer_REG[18] ( .CK(clk), .R(rst_n), .D(nxt_buffer[18]), .Q(buffer[18]), .QN( ));
Q_FDP1 \buffer_REG[17] ( .CK(clk), .R(rst_n), .D(nxt_buffer[17]), .Q(buffer[17]), .QN( ));
Q_FDP1 \buffer_REG[16] ( .CK(clk), .R(rst_n), .D(nxt_buffer[16]), .Q(buffer[16]), .QN( ));
Q_FDP1 \buffer_REG[15] ( .CK(clk), .R(rst_n), .D(nxt_buffer[15]), .Q(buffer[15]), .QN( ));
Q_FDP1 \buffer_REG[14] ( .CK(clk), .R(rst_n), .D(nxt_buffer[14]), .Q(buffer[14]), .QN( ));
Q_FDP1 \buffer_REG[13] ( .CK(clk), .R(rst_n), .D(nxt_buffer[13]), .Q(buffer[13]), .QN( ));
Q_FDP1 \buffer_REG[12] ( .CK(clk), .R(rst_n), .D(nxt_buffer[12]), .Q(buffer[12]), .QN( ));
Q_FDP1 \buffer_REG[11] ( .CK(clk), .R(rst_n), .D(nxt_buffer[11]), .Q(buffer[11]), .QN( ));
Q_FDP1 \buffer_REG[10] ( .CK(clk), .R(rst_n), .D(nxt_buffer[10]), .Q(buffer[10]), .QN( ));
Q_FDP1 \buffer_REG[9] ( .CK(clk), .R(rst_n), .D(nxt_buffer[9]), .Q(buffer[9]), .QN( ));
Q_FDP1 \buffer_REG[8] ( .CK(clk), .R(rst_n), .D(nxt_buffer[8]), .Q(buffer[8]), .QN( ));
Q_FDP1 \buffer_REG[7] ( .CK(clk), .R(rst_n), .D(nxt_buffer[7]), .Q(buffer[7]), .QN( ));
Q_FDP1 \buffer_REG[6] ( .CK(clk), .R(rst_n), .D(nxt_buffer[6]), .Q(buffer[6]), .QN( ));
Q_FDP1 \buffer_REG[5] ( .CK(clk), .R(rst_n), .D(nxt_buffer[5]), .Q(buffer[5]), .QN( ));
Q_FDP1 \buffer_REG[4] ( .CK(clk), .R(rst_n), .D(nxt_buffer[4]), .Q(buffer[4]), .QN( ));
Q_FDP1 \buffer_REG[3] ( .CK(clk), .R(rst_n), .D(nxt_buffer[3]), .Q(buffer[3]), .QN( ));
Q_FDP1 \buffer_REG[2] ( .CK(clk), .R(rst_n), .D(nxt_buffer[2]), .Q(buffer[2]), .QN( ));
Q_FDP1 \buffer_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_buffer[1]), .Q(buffer[1]), .QN( ));
Q_FDP1 \buffer_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_buffer[0]), .Q(buffer[0]), .QN( ));
Q_FDP1 \fifo_in_REG[67] ( .CK(clk), .R(rst_n), .D(nxt_fifo_in_id[3]), .Q(fifo_in[67]), .QN( ));
Q_FDP1 \fifo_in_REG[66] ( .CK(clk), .R(rst_n), .D(nxt_fifo_in_id[2]), .Q(fifo_in[66]), .QN( ));
Q_FDP1 \fifo_in_REG[65] ( .CK(clk), .R(rst_n), .D(nxt_fifo_in_id[1]), .Q(fifo_in[65]), .QN( ));
Q_FDP1 \fifo_in_REG[64] ( .CK(clk), .R(rst_n), .D(nxt_fifo_in_id[0]), .Q(fifo_in[64]), .QN( ));
Q_AN02 U5317 ( .A0(n2139), .A1(n1741), .Z(n1736));
Q_AN02 U5318 ( .A0(n2139), .A1(n1743), .Z(n1737));
Q_AN02 U5319 ( .A0(n2139), .A1(n1745), .Z(n1738));
Q_AN02 U5320 ( .A0(n2139), .A1(n1747), .Z(n1739));
Q_AN02 U5321 ( .A0(n2139), .A1(n1748), .Z(n1740));
Q_XOR2 U5322 ( .A0(tlv_counter[4]), .A1(n1742), .Z(n1741));
Q_AD01HF U5323 ( .A0(tlv_counter[3]), .B0(n1744), .S(n1743), .CO(n1742));
Q_AD01HF U5324 ( .A0(tlv_counter[2]), .B0(n1746), .S(n1745), .CO(n1744));
Q_AD01HF U5325 ( .A0(tlv_counter[1]), .B0(tlv_counter[0]), .S(n1747), .CO(n1746));
Q_AN02 U5326 ( .A0(rst_n), .A1(_zy_sva_b177), .Z(n1749));
Q_AN02 U5327 ( .A0(rst_n), .A1(_zy_sva_b176), .Z(n1750));
Q_AN02 U5328 ( .A0(rst_n), .A1(_zy_sva_b175), .Z(n1751));
Q_AN02 U5329 ( .A0(rst_n), .A1(_zy_sva_b174), .Z(n1752));
Q_AN02 U5330 ( .A0(rst_n), .A1(_zy_sva_b173), .Z(n1753));
Q_AN02 U5331 ( .A0(rst_n), .A1(_zy_sva_b172), .Z(n1754));
Q_AN02 U5332 ( .A0(rst_n), .A1(_zy_sva_b171), .Z(n1755));
Q_AN02 U5333 ( .A0(rst_n), .A1(_zy_sva_b170), .Z(n1756));
Q_AN02 U5334 ( .A0(rst_n), .A1(_zy_sva_b169), .Z(n1757));
Q_AN02 U5335 ( .A0(rst_n), .A1(_zy_sva_b168), .Z(n1758));
Q_AN02 U5336 ( .A0(rst_n), .A1(_zy_sva_b167), .Z(n1759));
Q_AN02 U5337 ( .A0(rst_n), .A1(_zy_sva_b166), .Z(n1760));
Q_AN02 U5338 ( .A0(rst_n), .A1(_zy_sva_b165), .Z(n1761));
Q_AN02 U5339 ( .A0(rst_n), .A1(_zy_sva_b164), .Z(n1762));
Q_AN02 U5340 ( .A0(rst_n), .A1(_zy_sva_b163), .Z(n1763));
Q_AN02 U5341 ( .A0(rst_n), .A1(_zy_sva_b162), .Z(n1764));
Q_AN02 U5342 ( .A0(rst_n), .A1(_zy_sva_b161), .Z(n1765));
Q_AN02 U5343 ( .A0(rst_n), .A1(_zy_sva_b160), .Z(n1766));
Q_AN02 U5344 ( .A0(rst_n), .A1(_zy_sva_b159), .Z(n1767));
Q_AN02 U5345 ( .A0(rst_n), .A1(_zy_sva_b158), .Z(n1768));
Q_AN02 U5346 ( .A0(rst_n), .A1(_zy_sva_b157), .Z(n1769));
Q_AN02 U5347 ( .A0(rst_n), .A1(_zy_sva_b156), .Z(n1770));
Q_AN02 U5348 ( .A0(rst_n), .A1(_zy_sva_b155), .Z(n1771));
Q_AN02 U5349 ( .A0(rst_n), .A1(_zy_sva_b154), .Z(n1772));
Q_AN02 U5350 ( .A0(rst_n), .A1(_zy_sva_b153), .Z(n1773));
Q_AN02 U5351 ( .A0(rst_n), .A1(_zy_sva_b152), .Z(n1774));
Q_AN02 U5352 ( .A0(rst_n), .A1(_zy_sva_b151), .Z(n1775));
Q_AN02 U5353 ( .A0(rst_n), .A1(_zy_sva_b150), .Z(n1776));
Q_AN02 U5354 ( .A0(rst_n), .A1(_zy_sva_b149), .Z(n1777));
Q_AN02 U5355 ( .A0(rst_n), .A1(_zy_sva_b148), .Z(n1778));
Q_AN02 U5356 ( .A0(rst_n), .A1(_zy_sva_b147), .Z(n1779));
Q_AN02 U5357 ( .A0(rst_n), .A1(_zy_sva_b146), .Z(n1780));
Q_AN02 U5358 ( .A0(rst_n), .A1(_zy_sva_b145), .Z(n1781));
Q_AN02 U5359 ( .A0(rst_n), .A1(_zy_sva_b144), .Z(n1782));
Q_AN02 U5360 ( .A0(rst_n), .A1(_zy_sva_b143), .Z(n1783));
Q_AN02 U5361 ( .A0(rst_n), .A1(_zy_sva_b142), .Z(n1784));
Q_AN02 U5362 ( .A0(rst_n), .A1(_zy_sva_b141), .Z(n1785));
Q_AN02 U5363 ( .A0(rst_n), .A1(_zy_sva_b140), .Z(n1786));
Q_AN02 U5364 ( .A0(rst_n), .A1(_zy_sva_b139), .Z(n1787));
Q_AN02 U5365 ( .A0(rst_n), .A1(_zy_sva_b138), .Z(n1788));
Q_AN02 U5366 ( .A0(rst_n), .A1(_zy_sva_b137), .Z(n1789));
Q_AN02 U5367 ( .A0(rst_n), .A1(_zy_sva_b136), .Z(n1790));
Q_AN02 U5368 ( .A0(rst_n), .A1(_zy_sva_b135), .Z(n1791));
Q_AN02 U5369 ( .A0(rst_n), .A1(_zy_sva_b134), .Z(n1792));
Q_AN02 U5370 ( .A0(rst_n), .A1(_zy_sva_b133), .Z(n1793));
Q_AN02 U5371 ( .A0(rst_n), .A1(_zy_sva_b132), .Z(n1794));
Q_AN02 U5372 ( .A0(rst_n), .A1(_zy_sva_b131), .Z(n1795));
Q_AN02 U5373 ( .A0(rst_n), .A1(_zy_sva_b130), .Z(n1796));
Q_AN02 U5374 ( .A0(rst_n), .A1(_zy_sva_b129), .Z(n1797));
Q_AN02 U5375 ( .A0(rst_n), .A1(_zy_sva_b128), .Z(n1798));
Q_AN02 U5376 ( .A0(rst_n), .A1(_zy_sva_b127), .Z(n1799));
Q_AN02 U5377 ( .A0(rst_n), .A1(_zy_sva_b126), .Z(n1800));
Q_AN02 U5378 ( .A0(rst_n), .A1(_zy_sva_b125), .Z(n1801));
Q_AN02 U5379 ( .A0(rst_n), .A1(_zy_sva_b124), .Z(n1802));
Q_AN02 U5380 ( .A0(rst_n), .A1(_zy_sva_b123), .Z(n1803));
Q_AN02 U5381 ( .A0(rst_n), .A1(_zy_sva_b122), .Z(n1804));
Q_AN02 U5382 ( .A0(rst_n), .A1(_zy_sva_b121), .Z(n1805));
Q_AN02 U5383 ( .A0(rst_n), .A1(_zy_sva_b120), .Z(n1806));
Q_AN02 U5384 ( .A0(rst_n), .A1(_zy_sva_b119), .Z(n1807));
Q_AN02 U5385 ( .A0(rst_n), .A1(_zy_sva_b118), .Z(n1808));
Q_AN02 U5386 ( .A0(rst_n), .A1(_zy_sva_b117), .Z(n1809));
Q_AN02 U5387 ( .A0(rst_n), .A1(_zy_sva_b116), .Z(n1810));
Q_AN02 U5388 ( .A0(rst_n), .A1(_zy_sva_b115), .Z(n1811));
Q_AN02 U5389 ( .A0(rst_n), .A1(_zy_sva_b114), .Z(n1812));
Q_AN02 U5390 ( .A0(rst_n), .A1(_zy_sva_b113), .Z(n1813));
Q_AN02 U5391 ( .A0(rst_n), .A1(_zy_sva_b112), .Z(n1814));
Q_AN02 U5392 ( .A0(rst_n), .A1(_zy_sva_b111), .Z(n1815));
Q_AN02 U5393 ( .A0(rst_n), .A1(_zy_sva_b110), .Z(n1816));
Q_AN02 U5394 ( .A0(rst_n), .A1(_zy_sva_b109), .Z(n1817));
Q_AN02 U5395 ( .A0(rst_n), .A1(_zy_sva_b108), .Z(n1818));
Q_AN02 U5396 ( .A0(rst_n), .A1(_zy_sva_b107), .Z(n1819));
Q_AN02 U5397 ( .A0(rst_n), .A1(_zy_sva_b106), .Z(n1820));
Q_AN02 U5398 ( .A0(rst_n), .A1(_zy_sva_b105), .Z(n1821));
Q_AN02 U5399 ( .A0(rst_n), .A1(_zy_sva_b104), .Z(n1822));
Q_AN02 U5400 ( .A0(rst_n), .A1(_zy_sva_b103), .Z(n1823));
Q_AN02 U5401 ( .A0(rst_n), .A1(_zy_sva_b102), .Z(n1824));
Q_AN02 U5402 ( .A0(rst_n), .A1(_zy_sva_b101), .Z(n1825));
Q_AN02 U5403 ( .A0(rst_n), .A1(_zy_sva_b100), .Z(n1826));
Q_AN02 U5404 ( .A0(rst_n), .A1(_zy_sva_b99), .Z(n1827));
Q_AN02 U5405 ( .A0(rst_n), .A1(_zy_sva_b98), .Z(n1828));
Q_AN02 U5406 ( .A0(rst_n), .A1(_zy_sva_b97), .Z(n1829));
Q_AN02 U5407 ( .A0(rst_n), .A1(_zy_sva_b96), .Z(n1830));
Q_AN02 U5408 ( .A0(rst_n), .A1(_zy_sva_b95), .Z(n1831));
Q_AN02 U5409 ( .A0(rst_n), .A1(_zy_sva_b94), .Z(n1832));
Q_AN02 U5410 ( .A0(rst_n), .A1(_zy_sva_b93), .Z(n1833));
Q_AN02 U5411 ( .A0(rst_n), .A1(_zy_sva_b92), .Z(n1834));
Q_AN02 U5412 ( .A0(rst_n), .A1(_zy_sva_b91), .Z(n1835));
Q_AN02 U5413 ( .A0(rst_n), .A1(_zy_sva_b90), .Z(n1836));
Q_AN02 U5414 ( .A0(rst_n), .A1(_zy_sva_b89), .Z(n1837));
Q_AN02 U5415 ( .A0(rst_n), .A1(_zy_sva_b88), .Z(n1838));
Q_AN02 U5416 ( .A0(rst_n), .A1(_zy_sva_b87), .Z(n1839));
Q_AN02 U5417 ( .A0(rst_n), .A1(_zy_sva_b86), .Z(n1840));
Q_AN02 U5418 ( .A0(rst_n), .A1(_zy_sva_b85), .Z(n1841));
Q_AN02 U5419 ( .A0(rst_n), .A1(_zy_sva_b84), .Z(n1842));
Q_AN02 U5420 ( .A0(rst_n), .A1(_zy_sva_b83), .Z(n1843));
Q_AN02 U5421 ( .A0(rst_n), .A1(_zy_sva_b82), .Z(n1844));
Q_AN02 U5422 ( .A0(rst_n), .A1(_zy_sva_b81), .Z(n1845));
Q_AN02 U5423 ( .A0(rst_n), .A1(_zy_sva_b80), .Z(n1846));
Q_AN02 U5424 ( .A0(rst_n), .A1(_zy_sva_b79), .Z(n1847));
Q_AN02 U5425 ( .A0(rst_n), .A1(_zy_sva_b78), .Z(n1848));
Q_AN02 U5426 ( .A0(rst_n), .A1(_zy_sva_b77), .Z(n1849));
Q_AN02 U5427 ( .A0(rst_n), .A1(_zy_sva_b76), .Z(n1850));
Q_AN02 U5428 ( .A0(rst_n), .A1(_zy_sva_b75), .Z(n1851));
Q_AN02 U5429 ( .A0(rst_n), .A1(_zy_sva_b74), .Z(n1852));
Q_AN02 U5430 ( .A0(rst_n), .A1(_zy_sva_b73), .Z(n1853));
Q_AN02 U5431 ( .A0(rst_n), .A1(_zy_sva_b72), .Z(n1854));
Q_AN02 U5432 ( .A0(rst_n), .A1(_zy_sva_b71), .Z(n1855));
Q_AN02 U5433 ( .A0(rst_n), .A1(_zy_sva_b70), .Z(n1856));
Q_AN02 U5434 ( .A0(rst_n), .A1(_zy_sva_b69), .Z(n1857));
Q_AN02 U5435 ( .A0(rst_n), .A1(_zy_sva_b68), .Z(n1858));
Q_AN02 U5436 ( .A0(rst_n), .A1(_zy_sva_b67), .Z(n1859));
Q_AN02 U5437 ( .A0(rst_n), .A1(_zy_sva_b66), .Z(n1860));
Q_AN02 U5438 ( .A0(rst_n), .A1(_zy_sva_b65), .Z(n1861));
Q_AN02 U5439 ( .A0(rst_n), .A1(_zy_sva_b64), .Z(n1862));
Q_AN02 U5440 ( .A0(rst_n), .A1(_zy_sva_b63), .Z(n1863));
Q_AN02 U5441 ( .A0(rst_n), .A1(_zy_sva_b62), .Z(n1864));
Q_AN02 U5442 ( .A0(rst_n), .A1(_zy_sva_b61), .Z(n1865));
Q_AN02 U5443 ( .A0(rst_n), .A1(_zy_sva_b60), .Z(n1866));
Q_AN02 U5444 ( .A0(rst_n), .A1(_zy_sva_b59), .Z(n1867));
Q_AN02 U5445 ( .A0(rst_n), .A1(_zy_sva_b58), .Z(n1868));
Q_AN02 U5446 ( .A0(rst_n), .A1(_zy_sva_b57), .Z(n1869));
Q_AN02 U5447 ( .A0(rst_n), .A1(_zy_sva_b56), .Z(n1870));
Q_AN02 U5448 ( .A0(rst_n), .A1(_zy_sva_b55), .Z(n1871));
Q_AN02 U5449 ( .A0(rst_n), .A1(_zy_sva_b54), .Z(n1872));
Q_AN02 U5450 ( .A0(rst_n), .A1(_zy_sva_b53), .Z(n1873));
Q_AN02 U5451 ( .A0(rst_n), .A1(_zy_sva_b52), .Z(n1874));
Q_AN02 U5452 ( .A0(rst_n), .A1(_zy_sva_b51), .Z(n1875));
Q_AN02 U5453 ( .A0(rst_n), .A1(_zy_sva_b50), .Z(n1876));
Q_AN02 U5454 ( .A0(rst_n), .A1(_zy_sva_b49), .Z(n1877));
Q_AN02 U5455 ( .A0(rst_n), .A1(_zy_sva_b48), .Z(n1878));
Q_AN02 U5456 ( .A0(rst_n), .A1(_zy_sva_b47), .Z(n1879));
Q_AN02 U5457 ( .A0(rst_n), .A1(_zy_sva_b46), .Z(n1880));
Q_AN02 U5458 ( .A0(rst_n), .A1(_zy_sva_b45), .Z(n1881));
Q_AN02 U5459 ( .A0(rst_n), .A1(_zy_sva_b44), .Z(n1882));
Q_AN02 U5460 ( .A0(rst_n), .A1(_zy_sva_b43), .Z(n1883));
Q_AN02 U5461 ( .A0(rst_n), .A1(_zy_sva_b42), .Z(n1884));
Q_AN02 U5462 ( .A0(rst_n), .A1(_zy_sva_b41), .Z(n1885));
Q_AN02 U5463 ( .A0(rst_n), .A1(_zy_sva_b40), .Z(n1886));
Q_AN02 U5464 ( .A0(rst_n), .A1(_zy_sva_b39), .Z(n1887));
Q_AN02 U5465 ( .A0(rst_n), .A1(_zy_sva_b38), .Z(n1888));
Q_AN02 U5466 ( .A0(rst_n), .A1(_zy_sva_b37), .Z(n1889));
Q_AN02 U5467 ( .A0(rst_n), .A1(_zy_sva_b36), .Z(n1890));
Q_AN02 U5468 ( .A0(rst_n), .A1(_zy_sva_b35), .Z(n1891));
Q_AN02 U5469 ( .A0(rst_n), .A1(_zy_sva_b34), .Z(n1892));
Q_AN02 U5470 ( .A0(rst_n), .A1(_zy_sva_b33), .Z(n1893));
Q_AN02 U5471 ( .A0(rst_n), .A1(_zy_sva_b32), .Z(n1894));
Q_AN02 U5472 ( .A0(rst_n), .A1(_zy_sva_b31), .Z(n1895));
Q_AN02 U5473 ( .A0(rst_n), .A1(_zy_sva_b30), .Z(n1896));
Q_AN02 U5474 ( .A0(rst_n), .A1(_zy_sva_b29), .Z(n1897));
Q_AN02 U5475 ( .A0(rst_n), .A1(_zy_sva_b28), .Z(n1898));
Q_AN02 U5476 ( .A0(rst_n), .A1(_zy_sva_b27), .Z(n1899));
Q_AN02 U5477 ( .A0(rst_n), .A1(_zy_sva_b26), .Z(n1900));
Q_AN02 U5478 ( .A0(rst_n), .A1(_zy_sva_b25), .Z(n1901));
Q_AN02 U5479 ( .A0(rst_n), .A1(_zy_sva_b24), .Z(n1902));
Q_AN02 U5480 ( .A0(rst_n), .A1(_zy_sva_b23), .Z(n1903));
Q_AN02 U5481 ( .A0(rst_n), .A1(_zy_sva_b22), .Z(n1904));
Q_AN02 U5482 ( .A0(rst_n), .A1(_zy_sva_b21), .Z(n1905));
Q_AN02 U5483 ( .A0(rst_n), .A1(_zy_sva_b20), .Z(n1906));
Q_AN02 U5484 ( .A0(rst_n), .A1(_zy_sva_b19), .Z(n1907));
Q_AN02 U5485 ( .A0(rst_n), .A1(_zy_sva_b18), .Z(n1908));
Q_AN02 U5486 ( .A0(rst_n), .A1(_zy_sva_b17), .Z(n1909));
Q_AN02 U5487 ( .A0(rst_n), .A1(_zy_sva_b16), .Z(n1910));
Q_AN02 U5488 ( .A0(rst_n), .A1(_zy_sva_b15), .Z(n1911));
Q_AN02 U5489 ( .A0(rst_n), .A1(_zy_sva_b14), .Z(n1912));
Q_AN02 U5490 ( .A0(rst_n), .A1(_zy_sva_b13), .Z(n1913));
Q_AN02 U5491 ( .A0(rst_n), .A1(_zy_sva_b12), .Z(n1914));
Q_AN02 U5492 ( .A0(rst_n), .A1(_zy_sva_b11), .Z(n1915));
Q_AN02 U5493 ( .A0(rst_n), .A1(_zy_sva_b10), .Z(n1916));
Q_AN02 U5494 ( .A0(rst_n), .A1(_zy_sva_b9), .Z(n1917));
Q_AN02 U5495 ( .A0(rst_n), .A1(_zy_sva_b8), .Z(n1918));
Q_AN02 U5496 ( .A0(rst_n), .A1(_zy_sva_b7), .Z(n1919));
Q_AN02 U5497 ( .A0(rst_n), .A1(_zy_sva_b6), .Z(n1920));
Q_AN02 U5498 ( .A0(rst_n), .A1(_zy_sva_b5), .Z(n1921));
Q_AN02 U5499 ( .A0(rst_n), .A1(_zy_sva_b4), .Z(n1922));
Q_AN02 U5500 ( .A0(rst_n), .A1(_zy_sva_b3), .Z(n1923));
Q_AN02 U5501 ( .A0(rst_n), .A1(_zy_sva_b2), .Z(n1924));
Q_AN02 U5502 ( .A0(rst_n), .A1(_zy_sva_b1), .Z(n1925));
Q_AN02 U5503 ( .A0(rst_n), .A1(_zy_sva_b0), .Z(n1926));
Q_INV U5504 ( .A(stitcher_out[64]), .Z(n2145));
Q_OR03 U5505 ( .A0(stitcher_out[71]), .A1(stitcher_out[70]), .A2(stitcher_out[69]), .Z(n2144));
Q_OR03 U5506 ( .A0(stitcher_out[68]), .A1(stitcher_out[67]), .A2(stitcher_out[66]), .Z(n2143));
Q_OR03 U5507 ( .A0(stitcher_out[65]), .A1(n2145), .A2(n2144), .Z(n2142));
Q_NR02 U5508 ( .A0(n2143), .A1(n2142), .Z(stitcher_sot));
Q_INV U5509 ( .A(stitcher_out[65]), .Z(n2141));
Q_OR03 U5510 ( .A0(n2141), .A1(stitcher_out[64]), .A2(n2144), .Z(n2140));
Q_OR02 U5511 ( .A0(n2143), .A1(n2140), .Z(n2139));
Q_INV U5512 ( .A(n2139), .Z(stitcher_eot));
Q_OR03 U5513 ( .A0(tlv_counter[4]), .A1(tlv_counter[3]), .A2(tlv_counter[2]), .Z(n2138));
Q_NR03 U5514 ( .A0(tlv_counter[1]), .A1(tlv_counter[0]), .A2(n2138), .Z(n2137));
Q_AN02 U5515 ( .A0(stitcher_empty), .A1(n2137), .Z(tlv_parser_idle));
Q_AN02 U5516 ( .A0(fifo_in_valid), .A1(fifo_in[70]), .Z(tlv_parser_int_tlv_start_pulse));
ixc_assign _zz_strnp_0 ( _zy_simnet_stitcher_rd_0_w$, stitcher_rd);
ixc_assign_71 _zz_strnp_1 ( _zy_simnet_parser_kimreader_data_1_w$[0:70], 
	parser_kimreader_data[70:0]);
ixc_assign_71 _zz_strnp_2 ( parser_kimreader_data[70:0], 
	_zy_simnet_parser_kimreader_data_2_w$[0:70]);
ixc_assign_71 _zz_strnp_3 ( _zy_simnet_fifo_in_5_w$[0:70], fifo_in[70:0]);
ixc_assign _zz_strnp_4 ( _zy_simnet_fifo_in_valid_6_w$, fifo_in_valid);
Q_INV U5522 ( .A(rst_n), .Z(_zy_sva_key_type0_line4_1_reset_or));
Q_OR03 U5523 ( .A0(int_tlv_counter[5]), .A1(int_tlv_counter[4]), .A2(int_tlv_counter[3]), .Z(n2134));
Q_OR03 U5524 ( .A0(n2135), .A1(n2136), .A2(int_tlv_counter[0]), .Z(n2133));
Q_OR02 U5525 ( .A0(n2134), .A1(n2133), .Z(n2132));
Q_INV U5526 ( .A(n2132), .Z(n2131));
Q_OR03 U5527 ( .A0(aux_auth_op[3]), .A1(aux_auth_op[2]), .A2(n2130), .Z(n2129));
Q_OR02 U5528 ( .A0(aux_auth_op[0]), .A1(n2129), .Z(n2128));
Q_INV U5529 ( .A(n2128), .Z(n2127));
Q_OR03 U5530 ( .A0(aux_raw_auth_op[3]), .A1(aux_raw_auth_op[2]), .A2(n2126), .Z(n2125));
Q_OR02 U5531 ( .A0(aux_raw_auth_op[0]), .A1(n2125), .Z(n2124));
Q_INV U5532 ( .A(n2124), .Z(n2123));
Q_ND02 U5533 ( .A0(n2128), .A1(n2124), .Z(n2122));
Q_OR03 U5534 ( .A0(aux_cipher_op[3]), .A1(aux_cipher_op[2]), .A2(aux_cipher_op[1]), .Z(n2121));
Q_OR02 U5535 ( .A0(aux_cipher_op[0]), .A1(n2121), .Z(n2120));
Q_INV U5536 ( .A(n2120), .Z(n2119));
Q_OR03 U5537 ( .A0(aux_key_type[5]), .A1(aux_key_type[4]), .A2(aux_key_type[3]), .Z(n2118));
Q_OR03 U5538 ( .A0(aux_key_type[2]), .A1(aux_key_type[1]), .A2(aux_key_type[0]), .Z(n2117));
Q_OR02 U5539 ( .A0(n2118), .A1(n2117), .Z(n2116));
Q_INV U5540 ( .A(n2116), .Z(n2115));
Q_NR03 U5541 ( .A0(n2116), .A1(n2120), .A2(n2132), .Z(n2114));
Q_AN02 U5542 ( .A0(n2122), .A1(n2114), .Z(_zy_sva_b0_t));
Q_OR03 U5543 ( .A0(aux_cipher_op[3]), .A1(aux_cipher_op[2]), .A2(n2113), .Z(n2112));
Q_OR02 U5544 ( .A0(aux_cipher_op[0]), .A1(n2112), .Z(n2111));
Q_INV U5545 ( .A(n2111), .Z(n2110));
Q_AN03 U5546 ( .A0(n2115), .A1(n2110), .A2(n2124), .Z(n2109));
Q_AN03 U5547 ( .A0(n2128), .A1(n2131), .A2(n2109), .Z(_zy_sva_b1_t));
Q_OR02 U5548 ( .A0(n2108), .A1(n2121), .Z(n2107));
Q_INV U5549 ( .A(n2107), .Z(n2106));
Q_AN03 U5550 ( .A0(n2115), .A1(n2106), .A2(n2124), .Z(n2105));
Q_AN03 U5551 ( .A0(n2128), .A1(n2131), .A2(n2105), .Z(_zy_sva_b2_t));
Q_OR03 U5552 ( .A0(aux_auth_op[3]), .A1(aux_auth_op[2]), .A2(aux_auth_op[1]), .Z(n2104));
Q_OR02 U5553 ( .A0(aux_auth_op[0]), .A1(n2104), .Z(n2103));
Q_INV U5554 ( .A(n2103), .Z(n2102));
Q_OR03 U5555 ( .A0(aux_raw_auth_op[3]), .A1(aux_raw_auth_op[2]), .A2(aux_raw_auth_op[1]), .Z(n2101));
Q_OR02 U5556 ( .A0(aux_raw_auth_op[0]), .A1(n2101), .Z(n2100));
Q_INV U5557 ( .A(n2100), .Z(n2099));
Q_OR03 U5558 ( .A0(aux_key_type[2]), .A1(aux_key_type[1]), .A2(n2098), .Z(n2097));
Q_OR02 U5559 ( .A0(n2118), .A1(n2097), .Z(n2096));
Q_INV U5560 ( .A(n2096), .Z(n2095));
Q_AN02 U5561 ( .A0(n2094), .A1(aux_key_header[16]), .Z(n2093));
Q_AN02 U5562 ( .A0(aux_key_header[15]), .A1(aux_key_header[16]), .Z(n2092));
Q_NR03 U5563 ( .A0(n2092), .A1(n2093), .A2(n2096), .Z(n2091));
Q_NR03 U5564 ( .A0(n2120), .A1(n2100), .A2(n2103), .Z(n2090));
Q_AN03 U5565 ( .A0(n2131), .A1(n2091), .A2(n2090), .Z(_zy_sva_b3_t));
Q_OR02 U5566 ( .A0(n2089), .A1(n2104), .Z(n2088));
Q_INV U5567 ( .A(n2088), .Z(n2087));
Q_OR02 U5568 ( .A0(n2086), .A1(n2101), .Z(n2085));
Q_INV U5569 ( .A(n2085), .Z(n2084));
Q_NR03 U5570 ( .A0(n2120), .A1(n2085), .A2(n2088), .Z(n2083));
Q_AN03 U5571 ( .A0(n2131), .A1(n2091), .A2(n2083), .Z(_zy_sva_b4_t));
Q_AN03 U5572 ( .A0(aux_key_header[16]), .A1(n2095), .A2(n2119), .Z(n2082));
Q_NR03 U5573 ( .A0(n2100), .A1(n2103), .A2(n2132), .Z(n2081));
Q_AN02 U5574 ( .A0(n2082), .A1(n2081), .Z(_zy_sva_b5_t));
Q_NR03 U5575 ( .A0(n2085), .A1(n2088), .A2(n2132), .Z(n2080));
Q_AN02 U5576 ( .A0(n2082), .A1(n2080), .Z(_zy_sva_b6_t));
Q_NR03 U5577 ( .A0(n2120), .A1(n2124), .A2(n2128), .Z(n2079));
Q_AN03 U5578 ( .A0(n2131), .A1(n2091), .A2(n2079), .Z(_zy_sva_b7_t));
Q_NR03 U5579 ( .A0(n2124), .A1(n2128), .A2(n2132), .Z(n2078));
Q_AN02 U5580 ( .A0(n2082), .A1(n2078), .Z(_zy_sva_b8_t));
Q_NR03 U5581 ( .A0(n2096), .A1(n2107), .A2(n2100), .Z(n2077));
Q_AN03 U5582 ( .A0(n2102), .A1(n2131), .A2(n2077), .Z(_zy_sva_b9_t));
Q_NR03 U5583 ( .A0(n2096), .A1(n2111), .A2(n2100), .Z(n2076));
Q_AN03 U5584 ( .A0(n2102), .A1(n2131), .A2(n2076), .Z(_zy_sva_b10_t));
Q_NR03 U5585 ( .A0(n2096), .A1(n2107), .A2(n2085), .Z(n2075));
Q_AN03 U5586 ( .A0(n2087), .A1(n2131), .A2(n2075), .Z(_zy_sva_b11_t));
Q_NR03 U5587 ( .A0(n2096), .A1(n2111), .A2(n2085), .Z(n2074));
Q_AN03 U5588 ( .A0(n2087), .A1(n2131), .A2(n2074), .Z(_zy_sva_b12_t));
Q_NR03 U5589 ( .A0(n2096), .A1(n2107), .A2(n2124), .Z(n2073));
Q_AN03 U5590 ( .A0(n2127), .A1(n2131), .A2(n2073), .Z(_zy_sva_b13_t));
Q_NR03 U5591 ( .A0(n2096), .A1(n2111), .A2(n2124), .Z(n2072));
Q_AN03 U5592 ( .A0(n2127), .A1(n2131), .A2(n2072), .Z(_zy_sva_b14_t));
Q_OR03 U5593 ( .A0(aux_key_type[5]), .A1(aux_key_type[4]), .A2(n2071), .Z(n2070));
Q_OR02 U5594 ( .A0(n2070), .A1(n2097), .Z(n2069));
Q_INV U5595 ( .A(n2069), .Z(n2068));
Q_NR03 U5596 ( .A0(n2092), .A1(n2093), .A2(n2069), .Z(n2067));
Q_AN03 U5597 ( .A0(n2131), .A1(n2067), .A2(n2079), .Z(_zy_sva_b15_t));
Q_AN03 U5598 ( .A0(aux_key_header[16]), .A1(n2068), .A2(n2119), .Z(n2066));
Q_AN02 U5599 ( .A0(n2066), .A1(n2078), .Z(_zy_sva_b16_t));
Q_NR03 U5600 ( .A0(n2069), .A1(n2107), .A2(n2124), .Z(n2065));
Q_AN03 U5601 ( .A0(n2127), .A1(n2131), .A2(n2065), .Z(_zy_sva_b17_t));
Q_NR03 U5602 ( .A0(n2069), .A1(n2111), .A2(n2124), .Z(n2064));
Q_AN03 U5603 ( .A0(n2127), .A1(n2131), .A2(n2064), .Z(_zy_sva_b18_t));
Q_AN03 U5604 ( .A0(n2131), .A1(n2067), .A2(n2090), .Z(_zy_sva_b19_t));
Q_AN03 U5605 ( .A0(n2131), .A1(n2067), .A2(n2083), .Z(_zy_sva_b20_t));
Q_AN02 U5606 ( .A0(n2066), .A1(n2081), .Z(_zy_sva_b21_t));
Q_AN02 U5607 ( .A0(n2066), .A1(n2080), .Z(_zy_sva_b22_t));
Q_NR03 U5608 ( .A0(n2069), .A1(n2107), .A2(n2100), .Z(n2063));
Q_AN03 U5609 ( .A0(n2102), .A1(n2131), .A2(n2063), .Z(_zy_sva_b23_t));
Q_NR03 U5610 ( .A0(n2069), .A1(n2107), .A2(n2085), .Z(n2062));
Q_AN03 U5611 ( .A0(n2087), .A1(n2131), .A2(n2062), .Z(_zy_sva_b24_t));
Q_NR03 U5612 ( .A0(n2069), .A1(n2111), .A2(n2100), .Z(n2061));
Q_AN03 U5613 ( .A0(n2102), .A1(n2131), .A2(n2061), .Z(_zy_sva_b25_t));
Q_NR03 U5614 ( .A0(n2069), .A1(n2111), .A2(n2085), .Z(n2060));
Q_AN03 U5615 ( .A0(n2087), .A1(n2131), .A2(n2060), .Z(_zy_sva_b26_t));
Q_OR03 U5616 ( .A0(tlv_type[7]), .A1(tlv_type[6]), .A2(tlv_type[5]), .Z(n2056));
Q_OR03 U5617 ( .A0(n2057), .A1(tlv_type[3]), .A2(n2058), .Z(n2055));
Q_OR03 U5618 ( .A0(tlv_type[1]), .A1(n2059), .A2(n2056), .Z(n2054));
Q_OR02 U5619 ( .A0(n2055), .A1(n2054), .Z(n2053));
Q_INV U5620 ( .A(n2053), .Z(n2052));
Q_NR02 U5621 ( .A0(aux_key_header[15]), .A1(aux_key_header[16]), .Z(n2051));
Q_AN03 U5622 ( .A0(n2050), .A1(aux_key_header[14]), .A2(n2051), .Z(n2049));
Q_AN03 U5623 ( .A0(n2131), .A1(n2049), .A2(n2052), .Z(_zy_sva_b27_t));
Q_AN03 U5624 ( .A0(aux_key_header[31]), .A1(n2048), .A2(n2051), .Z(n2047));
Q_AN03 U5625 ( .A0(n2131), .A1(n2047), .A2(n2052), .Z(_zy_sva_b28_t));
Q_AN03 U5626 ( .A0(n2050), .A1(aux_key_header[14]), .A2(n2093), .Z(n2046));
Q_AN03 U5627 ( .A0(n2131), .A1(n2046), .A2(n2052), .Z(_zy_sva_b29_t));
Q_AN03 U5628 ( .A0(aux_key_header[31]), .A1(n2048), .A2(n2093), .Z(n2045));
Q_AN03 U5629 ( .A0(n2131), .A1(n2045), .A2(n2052), .Z(_zy_sva_b30_t));
Q_AN03 U5630 ( .A0(tlv_type[1]), .A1(tlv_type[0]), .A2(n41), .Z(n2043));
Q_AN02 U5631 ( .A0(n40), .A1(n2043), .Z(n2042));
Q_AN03 U5632 ( .A0(n2131), .A1(n2049), .A2(n2042), .Z(_zy_sva_b31_t));
Q_AN03 U5633 ( .A0(n2131), .A1(n2047), .A2(n2042), .Z(_zy_sva_b32_t));
Q_AN03 U5634 ( .A0(n2131), .A1(n2046), .A2(n2042), .Z(_zy_sva_b33_t));
Q_AN03 U5635 ( .A0(n2131), .A1(n2045), .A2(n2042), .Z(_zy_sva_b34_t));
Q_AN02 U5636 ( .A0(n2041), .A1(aux_iv_op[1]), .Z(n2040));
Q_AN03 U5637 ( .A0(n2040), .A1(n2106), .A2(n2131), .Z(n2039));
Q_AN02 U5638 ( .A0(n2052), .A1(n2039), .Z(_zy_sva_b35_t));
Q_AN03 U5639 ( .A0(n2040), .A1(n2110), .A2(n2131), .Z(n2038));
Q_AN02 U5640 ( .A0(n2052), .A1(n2038), .Z(_zy_sva_b36_t));
Q_OR03 U5641 ( .A0(n2057), .A1(n2044), .A2(tlv_type[2]), .Z(n2037));
Q_OR03 U5642 ( .A0(tlv_type[1]), .A1(tlv_type[0]), .A2(n2056), .Z(n2036));
Q_OR02 U5643 ( .A0(n2037), .A1(n2036), .Z(n2035));
Q_INV U5644 ( .A(n2035), .Z(n2034));
Q_AN02 U5645 ( .A0(n2034), .A1(n2038), .Z(_zy_sva_b37_t));
Q_OR03 U5646 ( .A0(fifo_in[67]), .A1(fifo_in[66]), .A2(fifo_in[65]), .Z(n2033));
Q_OR02 U5647 ( .A0(fifo_in[64]), .A1(n2033), .Z(n2032));
Q_INV U5648 ( .A(n2032), .Z(n2031));
Q_OR03 U5649 ( .A0(stitcher_out[62]), .A1(stitcher_out[61]), .A2(stitcher_out[60]), .Z(n2030));
Q_OR03 U5650 ( .A0(stitcher_out[59]), .A1(stitcher_out[58]), .A2(stitcher_out[57]), .Z(n2029));
Q_OR02 U5651 ( .A0(n2030), .A1(n2029), .Z(n2028));
Q_NR03 U5652 ( .A0(n190), .A1(n2028), .A2(n2032), .Z(_zy_sva_b42_t));
Q_AN02 U5653 ( .A0(n2052), .A1(_zy_sva_b42_t), .Z(_zy_sva_b38_t));
Q_AN02 U5654 ( .A0(n2042), .A1(_zy_sva_b42_t), .Z(_zy_sva_b39_t));
Q_AN02 U5655 ( .A0(n2034), .A1(_zy_sva_b42_t), .Z(_zy_sva_b40_t));
Q_NR02 U5656 ( .A0(n2037), .A1(n2054), .Z(n2027));
Q_AN02 U5657 ( .A0(n2027), .A1(_zy_sva_b42_t), .Z(_zy_sva_b41_t));
Q_INV U5658 ( .A(stitcher_out[57]), .Z(n2026));
Q_OR03 U5659 ( .A0(stitcher_out[59]), .A1(stitcher_out[58]), .A2(n2026), .Z(n2025));
Q_OR02 U5660 ( .A0(n2030), .A1(n2025), .Z(n2024));
Q_NR03 U5661 ( .A0(n190), .A1(n2024), .A2(n2032), .Z(_zy_sva_b47_t));
Q_AN02 U5662 ( .A0(n2052), .A1(_zy_sva_b47_t), .Z(_zy_sva_b43_t));
Q_AN02 U5663 ( .A0(n2042), .A1(_zy_sva_b47_t), .Z(_zy_sva_b44_t));
Q_AN02 U5664 ( .A0(n2034), .A1(_zy_sva_b47_t), .Z(_zy_sva_b45_t));
Q_AN02 U5665 ( .A0(n2027), .A1(_zy_sva_b47_t), .Z(_zy_sva_b46_t));
Q_INV U5666 ( .A(stitcher_out[58]), .Z(n2023));
Q_OR03 U5667 ( .A0(stitcher_out[59]), .A1(n2023), .A2(stitcher_out[57]), .Z(n2022));
Q_OR02 U5668 ( .A0(n2030), .A1(n2022), .Z(n2021));
Q_NR03 U5669 ( .A0(n190), .A1(n2021), .A2(n2032), .Z(_zy_sva_b52_t));
Q_AN02 U5670 ( .A0(n2052), .A1(_zy_sva_b52_t), .Z(_zy_sva_b48_t));
Q_AN02 U5671 ( .A0(n2042), .A1(_zy_sva_b52_t), .Z(_zy_sva_b49_t));
Q_AN02 U5672 ( .A0(n2034), .A1(_zy_sva_b52_t), .Z(_zy_sva_b50_t));
Q_AN02 U5673 ( .A0(n2027), .A1(_zy_sva_b52_t), .Z(_zy_sva_b51_t));
Q_OR03 U5674 ( .A0(stitcher_out[59]), .A1(n2023), .A2(n2026), .Z(n2020));
Q_OR02 U5675 ( .A0(n2030), .A1(n2020), .Z(n2019));
Q_NR03 U5676 ( .A0(n190), .A1(n2019), .A2(n2032), .Z(_zy_sva_b57_t));
Q_AN02 U5677 ( .A0(n2052), .A1(_zy_sva_b57_t), .Z(_zy_sva_b53_t));
Q_AN02 U5678 ( .A0(n2042), .A1(_zy_sva_b57_t), .Z(_zy_sva_b54_t));
Q_AN02 U5679 ( .A0(n2034), .A1(_zy_sva_b57_t), .Z(_zy_sva_b55_t));
Q_AN02 U5680 ( .A0(n2027), .A1(_zy_sva_b57_t), .Z(_zy_sva_b56_t));
Q_INV U5681 ( .A(stitcher_out[59]), .Z(n2018));
Q_OR03 U5682 ( .A0(n2018), .A1(stitcher_out[58]), .A2(stitcher_out[57]), .Z(n2017));
Q_OR02 U5683 ( .A0(n2030), .A1(n2017), .Z(n2016));
Q_NR03 U5684 ( .A0(n190), .A1(n2016), .A2(n2032), .Z(_zy_sva_b62_t));
Q_AN02 U5685 ( .A0(n2052), .A1(_zy_sva_b62_t), .Z(_zy_sva_b58_t));
Q_AN02 U5686 ( .A0(n2042), .A1(_zy_sva_b62_t), .Z(_zy_sva_b59_t));
Q_AN02 U5687 ( .A0(n2034), .A1(_zy_sva_b62_t), .Z(_zy_sva_b60_t));
Q_AN02 U5688 ( .A0(n2027), .A1(_zy_sva_b62_t), .Z(_zy_sva_b61_t));
Q_OR03 U5689 ( .A0(n2018), .A1(stitcher_out[58]), .A2(n2026), .Z(n2015));
Q_OR02 U5690 ( .A0(n2030), .A1(n2015), .Z(n2014));
Q_NR03 U5691 ( .A0(n190), .A1(n2014), .A2(n2032), .Z(_zy_sva_b67_t));
Q_AN02 U5692 ( .A0(n2052), .A1(_zy_sva_b67_t), .Z(_zy_sva_b63_t));
Q_AN02 U5693 ( .A0(n2042), .A1(_zy_sva_b67_t), .Z(_zy_sva_b64_t));
Q_AN02 U5694 ( .A0(n2034), .A1(_zy_sva_b67_t), .Z(_zy_sva_b65_t));
Q_AN02 U5695 ( .A0(n2027), .A1(_zy_sva_b67_t), .Z(_zy_sva_b66_t));
Q_OR03 U5696 ( .A0(n2018), .A1(n2023), .A2(stitcher_out[57]), .Z(n2013));
Q_OR02 U5697 ( .A0(n2030), .A1(n2013), .Z(n2012));
Q_NR03 U5698 ( .A0(n190), .A1(n2012), .A2(n2032), .Z(_zy_sva_b72_t));
Q_AN02 U5699 ( .A0(n2052), .A1(_zy_sva_b72_t), .Z(_zy_sva_b68_t));
Q_AN02 U5700 ( .A0(n2042), .A1(_zy_sva_b72_t), .Z(_zy_sva_b69_t));
Q_AN02 U5701 ( .A0(n2034), .A1(_zy_sva_b72_t), .Z(_zy_sva_b70_t));
Q_AN02 U5702 ( .A0(n2027), .A1(_zy_sva_b72_t), .Z(_zy_sva_b71_t));
Q_INV U5703 ( .A(stitcher_out[60]), .Z(n2011));
Q_AN03 U5704 ( .A0(stitcher_out[59]), .A1(stitcher_out[58]), .A2(stitcher_out[57]), .Z(n2010));
Q_AN02 U5705 ( .A0(n37), .A1(n2010), .Z(n2009));
Q_AN03 U5706 ( .A0(fifo_in_valid), .A1(n2009), .A2(n2031), .Z(_zy_sva_b77_t));
Q_AN02 U5707 ( .A0(n2052), .A1(_zy_sva_b77_t), .Z(_zy_sva_b73_t));
Q_AN02 U5708 ( .A0(n2042), .A1(_zy_sva_b77_t), .Z(_zy_sva_b74_t));
Q_AN02 U5709 ( .A0(n2034), .A1(_zy_sva_b77_t), .Z(_zy_sva_b75_t));
Q_AN02 U5710 ( .A0(n2027), .A1(_zy_sva_b77_t), .Z(_zy_sva_b76_t));
Q_OR03 U5711 ( .A0(stitcher_out[62]), .A1(stitcher_out[61]), .A2(n2011), .Z(n2008));
Q_OR02 U5712 ( .A0(n2008), .A1(n2029), .Z(n2007));
Q_NR03 U5713 ( .A0(n190), .A1(n2007), .A2(n2032), .Z(_zy_sva_b82_t));
Q_AN02 U5714 ( .A0(n2052), .A1(_zy_sva_b82_t), .Z(_zy_sva_b78_t));
Q_AN02 U5715 ( .A0(n2042), .A1(_zy_sva_b82_t), .Z(_zy_sva_b79_t));
Q_AN02 U5716 ( .A0(n2034), .A1(_zy_sva_b82_t), .Z(_zy_sva_b80_t));
Q_AN02 U5717 ( .A0(n2027), .A1(_zy_sva_b82_t), .Z(_zy_sva_b81_t));
Q_OR02 U5718 ( .A0(n2008), .A1(n2025), .Z(n2006));
Q_NR03 U5719 ( .A0(n190), .A1(n2006), .A2(n2032), .Z(_zy_sva_b87_t));
Q_AN02 U5720 ( .A0(n2052), .A1(_zy_sva_b87_t), .Z(_zy_sva_b83_t));
Q_AN02 U5721 ( .A0(n2042), .A1(_zy_sva_b87_t), .Z(_zy_sva_b84_t));
Q_AN02 U5722 ( .A0(n2034), .A1(_zy_sva_b87_t), .Z(_zy_sva_b85_t));
Q_AN02 U5723 ( .A0(n2027), .A1(_zy_sva_b87_t), .Z(_zy_sva_b86_t));
Q_OR02 U5724 ( .A0(n2008), .A1(n2022), .Z(n2005));
Q_NR03 U5725 ( .A0(n190), .A1(n2005), .A2(n2032), .Z(_zy_sva_b92_t));
Q_AN02 U5726 ( .A0(n2052), .A1(_zy_sva_b92_t), .Z(_zy_sva_b88_t));
Q_AN02 U5727 ( .A0(n2042), .A1(_zy_sva_b92_t), .Z(_zy_sva_b89_t));
Q_AN02 U5728 ( .A0(n2034), .A1(_zy_sva_b92_t), .Z(_zy_sva_b90_t));
Q_AN02 U5729 ( .A0(n2027), .A1(_zy_sva_b92_t), .Z(_zy_sva_b91_t));
Q_NR02 U5730 ( .A0(n2008), .A1(n2020), .Z(n2004));
Q_AN03 U5731 ( .A0(fifo_in_valid), .A1(n2004), .A2(n2031), .Z(_zy_sva_b97_t));
Q_AN02 U5732 ( .A0(n2052), .A1(_zy_sva_b97_t), .Z(_zy_sva_b93_t));
Q_AN02 U5733 ( .A0(n2042), .A1(_zy_sva_b97_t), .Z(_zy_sva_b94_t));
Q_AN02 U5734 ( .A0(n2034), .A1(_zy_sva_b97_t), .Z(_zy_sva_b95_t));
Q_AN02 U5735 ( .A0(n2027), .A1(_zy_sva_b97_t), .Z(_zy_sva_b96_t));
Q_OR02 U5736 ( .A0(n2008), .A1(n2017), .Z(n2003));
Q_NR03 U5737 ( .A0(n190), .A1(n2003), .A2(n2032), .Z(_zy_sva_b102_t));
Q_AN02 U5738 ( .A0(n2052), .A1(_zy_sva_b102_t), .Z(_zy_sva_b98_t));
Q_AN02 U5739 ( .A0(n2042), .A1(_zy_sva_b102_t), .Z(_zy_sva_b99_t));
Q_AN02 U5740 ( .A0(n2034), .A1(_zy_sva_b102_t), .Z(_zy_sva_b100_t));
Q_AN02 U5741 ( .A0(n2027), .A1(_zy_sva_b102_t), .Z(_zy_sva_b101_t));
Q_NR02 U5742 ( .A0(n2008), .A1(n2015), .Z(n2002));
Q_AN03 U5743 ( .A0(fifo_in_valid), .A1(n2002), .A2(n2031), .Z(_zy_sva_b107_t));
Q_AN02 U5744 ( .A0(n2052), .A1(_zy_sva_b107_t), .Z(_zy_sva_b103_t));
Q_AN02 U5745 ( .A0(n2042), .A1(_zy_sva_b107_t), .Z(_zy_sva_b104_t));
Q_AN02 U5746 ( .A0(n2034), .A1(_zy_sva_b107_t), .Z(_zy_sva_b105_t));
Q_AN02 U5747 ( .A0(n2027), .A1(_zy_sva_b107_t), .Z(_zy_sva_b106_t));
Q_AN03 U5748 ( .A0(fifo_in[67]), .A1(fifo_in[66]), .A2(fifo_in[65]), .Z(n2001));
Q_AN02 U5749 ( .A0(fifo_in[64]), .A1(n2001), .Z(n2000));
Q_NR03 U5750 ( .A0(aux_key_header[31]), .A1(aux_key_header[14]), .A2(n190), .Z(n1999));
Q_AN03 U5751 ( .A0(n2051), .A1(n1999), .A2(n2000), .Z(_zy_sva_b108_t));
Q_AN03 U5752 ( .A0(aux_key_header[31]), .A1(n2048), .A2(fifo_in_valid), .Z(n1998));
Q_AN03 U5753 ( .A0(n2051), .A1(n1998), .A2(n2000), .Z(_zy_sva_b109_t));
Q_AN03 U5754 ( .A0(n2050), .A1(aux_key_header[14]), .A2(fifo_in_valid), .Z(n1997));
Q_AN03 U5755 ( .A0(n2051), .A1(n1997), .A2(n2000), .Z(_zy_sva_b110_t));
Q_AN03 U5756 ( .A0(aux_key_header[31]), .A1(aux_key_header[14]), .A2(fifo_in_valid), .Z(n1996));
Q_AN03 U5757 ( .A0(n2051), .A1(n1996), .A2(n2000), .Z(_zy_sva_b111_t));
Q_AN02 U5758 ( .A0(aux_key_header[15]), .A1(n1995), .Z(n1994));
Q_AN03 U5759 ( .A0(n1994), .A1(n1999), .A2(n2000), .Z(_zy_sva_b112_t));
Q_AN03 U5760 ( .A0(n1994), .A1(n1998), .A2(n2000), .Z(_zy_sva_b113_t));
Q_AN03 U5761 ( .A0(n1994), .A1(n1997), .A2(n2000), .Z(_zy_sva_b114_t));
Q_AN03 U5762 ( .A0(n1994), .A1(n1996), .A2(n2000), .Z(_zy_sva_b115_t));
Q_AN03 U5763 ( .A0(n2093), .A1(n1999), .A2(n2000), .Z(_zy_sva_b116_t));
Q_AN03 U5764 ( .A0(n2093), .A1(n1998), .A2(n2000), .Z(_zy_sva_b117_t));
Q_AN03 U5765 ( .A0(n2093), .A1(n1997), .A2(n2000), .Z(_zy_sva_b118_t));
Q_AN03 U5766 ( .A0(n2093), .A1(n1996), .A2(n2000), .Z(_zy_sva_b119_t));
Q_AN03 U5767 ( .A0(n2092), .A1(n1999), .A2(n2000), .Z(_zy_sva_b120_t));
Q_AN03 U5768 ( .A0(n2092), .A1(n1998), .A2(n2000), .Z(_zy_sva_b121_t));
Q_AN03 U5769 ( .A0(n2092), .A1(n1997), .A2(n2000), .Z(_zy_sva_b122_t));
Q_AN03 U5770 ( .A0(n2092), .A1(n1996), .A2(n2000), .Z(_zy_sva_b123_t));
Q_AN03 U5771 ( .A0(aux_key_type[2]), .A1(aux_key_type[1]), .A2(aux_key_type[0]), .Z(n1993));
Q_AN02 U5772 ( .A0(n38), .A1(n1993), .Z(n1992));
Q_AN03 U5773 ( .A0(n1992), .A1(n2106), .A2(n2099), .Z(n1991));
Q_AN03 U5774 ( .A0(n2102), .A1(n2131), .A2(n1991), .Z(_zy_sva_b124_t));
Q_AN03 U5775 ( .A0(n1992), .A1(n2106), .A2(n2084), .Z(n1990));
Q_AN03 U5776 ( .A0(n2087), .A1(n2131), .A2(n1990), .Z(_zy_sva_b125_t));
Q_AN03 U5777 ( .A0(n1992), .A1(n2110), .A2(n2099), .Z(n1989));
Q_AN03 U5778 ( .A0(n2102), .A1(n2131), .A2(n1989), .Z(_zy_sva_b126_t));
Q_AN03 U5779 ( .A0(n1992), .A1(n2110), .A2(n2084), .Z(n1988));
Q_AN03 U5780 ( .A0(n2087), .A1(n2131), .A2(n1988), .Z(_zy_sva_b127_t));
Q_AN03 U5781 ( .A0(n1992), .A1(n2119), .A2(n2099), .Z(n1987));
Q_AN03 U5782 ( .A0(n2102), .A1(n2131), .A2(n1987), .Z(_zy_sva_b128_t));
Q_AN03 U5783 ( .A0(n1992), .A1(n2119), .A2(n2084), .Z(n1986));
Q_AN03 U5784 ( .A0(n2087), .A1(n2131), .A2(n1986), .Z(_zy_sva_b129_t));
Q_AN03 U5785 ( .A0(n1992), .A1(n2106), .A2(n2123), .Z(n1985));
Q_AN03 U5786 ( .A0(n2127), .A1(n2131), .A2(n1985), .Z(_zy_sva_b130_t));
Q_AN03 U5787 ( .A0(n1992), .A1(n2110), .A2(n2123), .Z(n1984));
Q_AN03 U5788 ( .A0(n2127), .A1(n2131), .A2(n1984), .Z(_zy_sva_b131_t));
Q_AN03 U5789 ( .A0(n1992), .A1(n2119), .A2(n2123), .Z(n1983));
Q_AN03 U5790 ( .A0(n2127), .A1(n2131), .A2(n1983), .Z(_zy_sva_b132_t));
Q_OR02 U5791 ( .A0(n2070), .A1(n2117), .Z(n1982));
Q_NR03 U5792 ( .A0(n1982), .A1(n2107), .A2(n2100), .Z(n1981));
Q_AN03 U5793 ( .A0(n2102), .A1(n2131), .A2(n1981), .Z(_zy_sva_b133_t));
Q_NR03 U5794 ( .A0(n1982), .A1(n2107), .A2(n2085), .Z(n1980));
Q_AN03 U5795 ( .A0(n2087), .A1(n2131), .A2(n1980), .Z(_zy_sva_b134_t));
Q_NR03 U5796 ( .A0(n1982), .A1(n2111), .A2(n2100), .Z(n1979));
Q_AN03 U5797 ( .A0(n2102), .A1(n2131), .A2(n1979), .Z(_zy_sva_b135_t));
Q_NR03 U5798 ( .A0(n1982), .A1(n2111), .A2(n2085), .Z(n1978));
Q_AN03 U5799 ( .A0(n2087), .A1(n2131), .A2(n1978), .Z(_zy_sva_b136_t));
Q_NR03 U5800 ( .A0(n1982), .A1(n2120), .A2(n2100), .Z(n1977));
Q_AN03 U5801 ( .A0(n2102), .A1(n2131), .A2(n1977), .Z(_zy_sva_b137_t));
Q_NR03 U5802 ( .A0(n1982), .A1(n2120), .A2(n2085), .Z(n1976));
Q_AN03 U5803 ( .A0(n2087), .A1(n2131), .A2(n1976), .Z(_zy_sva_b138_t));
Q_NR03 U5804 ( .A0(n1982), .A1(n2107), .A2(n2124), .Z(n1975));
Q_AN03 U5805 ( .A0(n2127), .A1(n2131), .A2(n1975), .Z(_zy_sva_b139_t));
Q_NR03 U5806 ( .A0(n1982), .A1(n2111), .A2(n2124), .Z(n1974));
Q_AN03 U5807 ( .A0(n2127), .A1(n2131), .A2(n1974), .Z(_zy_sva_b140_t));
Q_NR03 U5808 ( .A0(n1982), .A1(n2120), .A2(n2124), .Z(n1973));
Q_AN03 U5809 ( .A0(n2127), .A1(n2131), .A2(n1973), .Z(_zy_sva_b141_t));
Q_OR03 U5810 ( .A0(aux_key_type[2]), .A1(n1972), .A2(aux_key_type[0]), .Z(n1971));
Q_OR02 U5811 ( .A0(n2070), .A1(n1971), .Z(n1970));
Q_NR03 U5812 ( .A0(n1970), .A1(n2107), .A2(n2100), .Z(n1969));
Q_AN03 U5813 ( .A0(n2102), .A1(n2131), .A2(n1969), .Z(_zy_sva_b142_t));
Q_NR03 U5814 ( .A0(n1970), .A1(n2107), .A2(n2085), .Z(n1968));
Q_AN03 U5815 ( .A0(n2087), .A1(n2131), .A2(n1968), .Z(_zy_sva_b143_t));
Q_NR03 U5816 ( .A0(n1970), .A1(n2111), .A2(n2100), .Z(n1967));
Q_AN03 U5817 ( .A0(n2102), .A1(n2131), .A2(n1967), .Z(_zy_sva_b144_t));
Q_NR03 U5818 ( .A0(n1970), .A1(n2111), .A2(n2085), .Z(n1966));
Q_AN03 U5819 ( .A0(n2087), .A1(n2131), .A2(n1966), .Z(_zy_sva_b145_t));
Q_NR03 U5820 ( .A0(n1970), .A1(n2120), .A2(n2100), .Z(n1965));
Q_AN03 U5821 ( .A0(n2102), .A1(n2131), .A2(n1965), .Z(_zy_sva_b146_t));
Q_NR03 U5822 ( .A0(n1970), .A1(n2120), .A2(n2085), .Z(n1964));
Q_AN03 U5823 ( .A0(n2087), .A1(n2131), .A2(n1964), .Z(_zy_sva_b147_t));
Q_NR03 U5824 ( .A0(n1970), .A1(n2107), .A2(n2124), .Z(n1963));
Q_AN03 U5825 ( .A0(n2127), .A1(n2131), .A2(n1963), .Z(_zy_sva_b148_t));
Q_NR03 U5826 ( .A0(n1970), .A1(n2111), .A2(n2124), .Z(n1962));
Q_AN03 U5827 ( .A0(n2127), .A1(n2131), .A2(n1962), .Z(_zy_sva_b149_t));
Q_NR03 U5828 ( .A0(n1970), .A1(n2120), .A2(n2124), .Z(n1961));
Q_AN03 U5829 ( .A0(n2127), .A1(n2131), .A2(n1961), .Z(_zy_sva_b150_t));
Q_AN03 U5830 ( .A0(n1960), .A1(aux_key_type[1]), .A2(aux_key_type[0]), .Z(n1959));
Q_AN02 U5831 ( .A0(n39), .A1(n1959), .Z(n1958));
Q_AN03 U5832 ( .A0(n1958), .A1(n2106), .A2(n2099), .Z(n1957));
Q_AN03 U5833 ( .A0(n2102), .A1(n2131), .A2(n1957), .Z(_zy_sva_b151_t));
Q_AN03 U5834 ( .A0(n1958), .A1(n2106), .A2(n2084), .Z(n1956));
Q_AN03 U5835 ( .A0(n2087), .A1(n2131), .A2(n1956), .Z(_zy_sva_b152_t));
Q_AN03 U5836 ( .A0(n1958), .A1(n2110), .A2(n2099), .Z(n1955));
Q_AN03 U5837 ( .A0(n2102), .A1(n2131), .A2(n1955), .Z(_zy_sva_b153_t));
Q_AN03 U5838 ( .A0(n1958), .A1(n2110), .A2(n2084), .Z(n1954));
Q_AN03 U5839 ( .A0(n2087), .A1(n2131), .A2(n1954), .Z(_zy_sva_b154_t));
Q_AN03 U5840 ( .A0(n1958), .A1(n2119), .A2(n2099), .Z(n1953));
Q_AN03 U5841 ( .A0(n2102), .A1(n2131), .A2(n1953), .Z(_zy_sva_b155_t));
Q_AN03 U5842 ( .A0(n1958), .A1(n2119), .A2(n2084), .Z(n1952));
Q_AN03 U5843 ( .A0(n2087), .A1(n2131), .A2(n1952), .Z(_zy_sva_b156_t));
Q_AN03 U5844 ( .A0(n1958), .A1(n2106), .A2(n2123), .Z(n1951));
Q_AN03 U5845 ( .A0(n2127), .A1(n2131), .A2(n1951), .Z(_zy_sva_b157_t));
Q_AN03 U5846 ( .A0(n1958), .A1(n2110), .A2(n2123), .Z(n1950));
Q_AN03 U5847 ( .A0(n2127), .A1(n2131), .A2(n1950), .Z(_zy_sva_b158_t));
Q_AN03 U5848 ( .A0(n1958), .A1(n2119), .A2(n2123), .Z(n1949));
Q_AN03 U5849 ( .A0(n2127), .A1(n2131), .A2(n1949), .Z(_zy_sva_b159_t));
Q_OR03 U5850 ( .A0(n1960), .A1(aux_key_type[1]), .A2(aux_key_type[0]), .Z(n1948));
Q_OR02 U5851 ( .A0(n2070), .A1(n1948), .Z(n1947));
Q_NR03 U5852 ( .A0(n1947), .A1(n2107), .A2(n2100), .Z(n1946));
Q_AN03 U5853 ( .A0(n2102), .A1(n2131), .A2(n1946), .Z(_zy_sva_b160_t));
Q_NR03 U5854 ( .A0(n1947), .A1(n2107), .A2(n2085), .Z(n1945));
Q_AN03 U5855 ( .A0(n2087), .A1(n2131), .A2(n1945), .Z(_zy_sva_b161_t));
Q_NR03 U5856 ( .A0(n1947), .A1(n2111), .A2(n2100), .Z(n1944));
Q_AN03 U5857 ( .A0(n2102), .A1(n2131), .A2(n1944), .Z(_zy_sva_b162_t));
Q_NR03 U5858 ( .A0(n1947), .A1(n2111), .A2(n2085), .Z(n1943));
Q_AN03 U5859 ( .A0(n2087), .A1(n2131), .A2(n1943), .Z(_zy_sva_b163_t));
Q_NR03 U5860 ( .A0(n1947), .A1(n2120), .A2(n2100), .Z(n1942));
Q_AN03 U5861 ( .A0(n2102), .A1(n2131), .A2(n1942), .Z(_zy_sva_b164_t));
Q_NR03 U5862 ( .A0(n1947), .A1(n2120), .A2(n2085), .Z(n1941));
Q_AN03 U5863 ( .A0(n2087), .A1(n2131), .A2(n1941), .Z(_zy_sva_b165_t));
Q_NR03 U5864 ( .A0(n1947), .A1(n2107), .A2(n2124), .Z(n1940));
Q_AN03 U5865 ( .A0(n2127), .A1(n2131), .A2(n1940), .Z(_zy_sva_b166_t));
Q_NR03 U5866 ( .A0(n1947), .A1(n2111), .A2(n2124), .Z(n1939));
Q_AN03 U5867 ( .A0(n2127), .A1(n2131), .A2(n1939), .Z(_zy_sva_b167_t));
Q_NR03 U5868 ( .A0(n1947), .A1(n2120), .A2(n2124), .Z(n1938));
Q_AN03 U5869 ( .A0(n2127), .A1(n2131), .A2(n1938), .Z(_zy_sva_b168_t));
Q_AN03 U5870 ( .A0(aux_key_type[2]), .A1(n1972), .A2(aux_key_type[0]), .Z(n1937));
Q_AN02 U5871 ( .A0(n39), .A1(n1937), .Z(n1936));
Q_AN03 U5872 ( .A0(n1936), .A1(n2106), .A2(n2099), .Z(n1935));
Q_AN03 U5873 ( .A0(n2102), .A1(n2131), .A2(n1935), .Z(_zy_sva_b169_t));
Q_AN03 U5874 ( .A0(n1936), .A1(n2106), .A2(n2084), .Z(n1934));
Q_AN03 U5875 ( .A0(n2087), .A1(n2131), .A2(n1934), .Z(_zy_sva_b170_t));
Q_AN03 U5876 ( .A0(n1936), .A1(n2110), .A2(n2099), .Z(n1933));
Q_AN03 U5877 ( .A0(n2102), .A1(n2131), .A2(n1933), .Z(_zy_sva_b171_t));
Q_AN03 U5878 ( .A0(n1936), .A1(n2110), .A2(n2084), .Z(n1932));
Q_AN03 U5879 ( .A0(n2087), .A1(n2131), .A2(n1932), .Z(_zy_sva_b172_t));
Q_AN03 U5880 ( .A0(n1936), .A1(n2119), .A2(n2099), .Z(n1931));
Q_AN03 U5881 ( .A0(n2102), .A1(n2131), .A2(n1931), .Z(_zy_sva_b173_t));
Q_AN03 U5882 ( .A0(n1936), .A1(n2119), .A2(n2084), .Z(n1930));
Q_AN03 U5883 ( .A0(n2087), .A1(n2131), .A2(n1930), .Z(_zy_sva_b174_t));
Q_AN03 U5884 ( .A0(n1936), .A1(n2106), .A2(n2123), .Z(n1929));
Q_AN03 U5885 ( .A0(n2127), .A1(n2131), .A2(n1929), .Z(_zy_sva_b175_t));
Q_AN03 U5886 ( .A0(n1936), .A1(n2110), .A2(n2123), .Z(n1928));
Q_AN03 U5887 ( .A0(n2127), .A1(n2131), .A2(n1928), .Z(_zy_sva_b176_t));
Q_AN03 U5888 ( .A0(n1936), .A1(n2119), .A2(n2123), .Z(n1927));
Q_AN03 U5889 ( .A0(n2127), .A1(n2131), .A2(n1927), .Z(_zy_sva_b177_t));
ixc_sample_logic_1_3 _zz_zy_sva_b0 ( _zy_sva_b0, _zy_sva_b0_t);
ixc_sample_logic_1_3 _zz_zy_sva_b1 ( _zy_sva_b1, _zy_sva_b1_t);
ixc_sample_logic_1_3 _zz_zy_sva_b2 ( _zy_sva_b2, _zy_sva_b2_t);
ixc_sample_logic_1_3 _zz_zy_sva_b3 ( _zy_sva_b3, _zy_sva_b3_t);
ixc_sample_logic_1_3 _zz_zy_sva_b4 ( _zy_sva_b4, _zy_sva_b4_t);
ixc_sample_logic_1_3 _zz_zy_sva_b5 ( _zy_sva_b5, _zy_sva_b5_t);
ixc_sample_logic_1_3 _zz_zy_sva_b6 ( _zy_sva_b6, _zy_sva_b6_t);
ixc_sample_logic_1_3 _zz_zy_sva_b7 ( _zy_sva_b7, _zy_sva_b7_t);
ixc_sample_logic_1_3 _zz_zy_sva_b8 ( _zy_sva_b8, _zy_sva_b8_t);
ixc_sample_logic_1_3 _zz_zy_sva_b9 ( _zy_sva_b9, _zy_sva_b9_t);
ixc_sample_logic_1_3 _zz_zy_sva_b10 ( _zy_sva_b10, _zy_sva_b10_t);
ixc_sample_logic_1_3 _zz_zy_sva_b11 ( _zy_sva_b11, _zy_sva_b11_t);
ixc_sample_logic_1_3 _zz_zy_sva_b12 ( _zy_sva_b12, _zy_sva_b12_t);
ixc_sample_logic_1_3 _zz_zy_sva_b13 ( _zy_sva_b13, _zy_sva_b13_t);
ixc_sample_logic_1_3 _zz_zy_sva_b14 ( _zy_sva_b14, _zy_sva_b14_t);
ixc_sample_logic_1_3 _zz_zy_sva_b15 ( _zy_sva_b15, _zy_sva_b15_t);
ixc_sample_logic_1_3 _zz_zy_sva_b16 ( _zy_sva_b16, _zy_sva_b16_t);
ixc_sample_logic_1_3 _zz_zy_sva_b17 ( _zy_sva_b17, _zy_sva_b17_t);
ixc_sample_logic_1_3 _zz_zy_sva_b18 ( _zy_sva_b18, _zy_sva_b18_t);
ixc_sample_logic_1_3 _zz_zy_sva_b19 ( _zy_sva_b19, _zy_sva_b19_t);
ixc_sample_logic_1_3 _zz_zy_sva_b20 ( _zy_sva_b20, _zy_sva_b20_t);
ixc_sample_logic_1_3 _zz_zy_sva_b21 ( _zy_sva_b21, _zy_sva_b21_t);
ixc_sample_logic_1_3 _zz_zy_sva_b22 ( _zy_sva_b22, _zy_sva_b22_t);
ixc_sample_logic_1_3 _zz_zy_sva_b23 ( _zy_sva_b23, _zy_sva_b23_t);
ixc_sample_logic_1_3 _zz_zy_sva_b24 ( _zy_sva_b24, _zy_sva_b24_t);
ixc_sample_logic_1_3 _zz_zy_sva_b25 ( _zy_sva_b25, _zy_sva_b25_t);
ixc_sample_logic_1_3 _zz_zy_sva_b26 ( _zy_sva_b26, _zy_sva_b26_t);
ixc_sample_logic_1_3 _zz_zy_sva_b27 ( _zy_sva_b27, _zy_sva_b27_t);
ixc_sample_logic_1_3 _zz_zy_sva_b28 ( _zy_sva_b28, _zy_sva_b28_t);
ixc_sample_logic_1_3 _zz_zy_sva_b29 ( _zy_sva_b29, _zy_sva_b29_t);
ixc_sample_logic_1_3 _zz_zy_sva_b30 ( _zy_sva_b30, _zy_sva_b30_t);
ixc_sample_logic_1_3 _zz_zy_sva_b31 ( _zy_sva_b31, _zy_sva_b31_t);
ixc_sample_logic_1_3 _zz_zy_sva_b32 ( _zy_sva_b32, _zy_sva_b32_t);
ixc_sample_logic_1_3 _zz_zy_sva_b33 ( _zy_sva_b33, _zy_sva_b33_t);
ixc_sample_logic_1_3 _zz_zy_sva_b34 ( _zy_sva_b34, _zy_sva_b34_t);
ixc_sample_logic_1_3 _zz_zy_sva_b35 ( _zy_sva_b35, _zy_sva_b35_t);
ixc_sample_logic_1_3 _zz_zy_sva_b36 ( _zy_sva_b36, _zy_sva_b36_t);
ixc_sample_logic_1_3 _zz_zy_sva_b37 ( _zy_sva_b37, _zy_sva_b37_t);
ixc_sample_logic_1_3 _zz_zy_sva_b38 ( _zy_sva_b38, _zy_sva_b38_t);
ixc_sample_logic_1_3 _zz_zy_sva_b39 ( _zy_sva_b39, _zy_sva_b39_t);
ixc_sample_logic_1_3 _zz_zy_sva_b40 ( _zy_sva_b40, _zy_sva_b40_t);
ixc_sample_logic_1_3 _zz_zy_sva_b41 ( _zy_sva_b41, _zy_sva_b41_t);
ixc_sample_logic_1_3 _zz_zy_sva_b42 ( _zy_sva_b42, _zy_sva_b42_t);
ixc_sample_logic_1_3 _zz_zy_sva_b43 ( _zy_sva_b43, _zy_sva_b43_t);
ixc_sample_logic_1_3 _zz_zy_sva_b44 ( _zy_sva_b44, _zy_sva_b44_t);
ixc_sample_logic_1_3 _zz_zy_sva_b45 ( _zy_sva_b45, _zy_sva_b45_t);
ixc_sample_logic_1_3 _zz_zy_sva_b46 ( _zy_sva_b46, _zy_sva_b46_t);
ixc_sample_logic_1_3 _zz_zy_sva_b47 ( _zy_sva_b47, _zy_sva_b47_t);
ixc_sample_logic_1_3 _zz_zy_sva_b48 ( _zy_sva_b48, _zy_sva_b48_t);
ixc_sample_logic_1_3 _zz_zy_sva_b49 ( _zy_sva_b49, _zy_sva_b49_t);
ixc_sample_logic_1_3 _zz_zy_sva_b50 ( _zy_sva_b50, _zy_sva_b50_t);
ixc_sample_logic_1_3 _zz_zy_sva_b51 ( _zy_sva_b51, _zy_sva_b51_t);
ixc_sample_logic_1_3 _zz_zy_sva_b52 ( _zy_sva_b52, _zy_sva_b52_t);
ixc_sample_logic_1_3 _zz_zy_sva_b53 ( _zy_sva_b53, _zy_sva_b53_t);
ixc_sample_logic_1_3 _zz_zy_sva_b54 ( _zy_sva_b54, _zy_sva_b54_t);
ixc_sample_logic_1_3 _zz_zy_sva_b55 ( _zy_sva_b55, _zy_sva_b55_t);
ixc_sample_logic_1_3 _zz_zy_sva_b56 ( _zy_sva_b56, _zy_sva_b56_t);
ixc_sample_logic_1_3 _zz_zy_sva_b57 ( _zy_sva_b57, _zy_sva_b57_t);
ixc_sample_logic_1_3 _zz_zy_sva_b58 ( _zy_sva_b58, _zy_sva_b58_t);
ixc_sample_logic_1_3 _zz_zy_sva_b59 ( _zy_sva_b59, _zy_sva_b59_t);
ixc_sample_logic_1_3 _zz_zy_sva_b60 ( _zy_sva_b60, _zy_sva_b60_t);
ixc_sample_logic_1_3 _zz_zy_sva_b61 ( _zy_sva_b61, _zy_sva_b61_t);
ixc_sample_logic_1_3 _zz_zy_sva_b62 ( _zy_sva_b62, _zy_sva_b62_t);
ixc_sample_logic_1_3 _zz_zy_sva_b63 ( _zy_sva_b63, _zy_sva_b63_t);
ixc_sample_logic_1_3 _zz_zy_sva_b64 ( _zy_sva_b64, _zy_sva_b64_t);
ixc_sample_logic_1_3 _zz_zy_sva_b65 ( _zy_sva_b65, _zy_sva_b65_t);
ixc_sample_logic_1_3 _zz_zy_sva_b66 ( _zy_sva_b66, _zy_sva_b66_t);
ixc_sample_logic_1_3 _zz_zy_sva_b67 ( _zy_sva_b67, _zy_sva_b67_t);
ixc_sample_logic_1_3 _zz_zy_sva_b68 ( _zy_sva_b68, _zy_sva_b68_t);
ixc_sample_logic_1_3 _zz_zy_sva_b69 ( _zy_sva_b69, _zy_sva_b69_t);
ixc_sample_logic_1_3 _zz_zy_sva_b70 ( _zy_sva_b70, _zy_sva_b70_t);
ixc_sample_logic_1_3 _zz_zy_sva_b71 ( _zy_sva_b71, _zy_sva_b71_t);
ixc_sample_logic_1_3 _zz_zy_sva_b72 ( _zy_sva_b72, _zy_sva_b72_t);
ixc_sample_logic_1_3 _zz_zy_sva_b73 ( _zy_sva_b73, _zy_sva_b73_t);
ixc_sample_logic_1_3 _zz_zy_sva_b74 ( _zy_sva_b74, _zy_sva_b74_t);
ixc_sample_logic_1_3 _zz_zy_sva_b75 ( _zy_sva_b75, _zy_sva_b75_t);
ixc_sample_logic_1_3 _zz_zy_sva_b76 ( _zy_sva_b76, _zy_sva_b76_t);
ixc_sample_logic_1_3 _zz_zy_sva_b77 ( _zy_sva_b77, _zy_sva_b77_t);
ixc_sample_logic_1_3 _zz_zy_sva_b78 ( _zy_sva_b78, _zy_sva_b78_t);
ixc_sample_logic_1_3 _zz_zy_sva_b79 ( _zy_sva_b79, _zy_sva_b79_t);
ixc_sample_logic_1_3 _zz_zy_sva_b80 ( _zy_sva_b80, _zy_sva_b80_t);
ixc_sample_logic_1_3 _zz_zy_sva_b81 ( _zy_sva_b81, _zy_sva_b81_t);
ixc_sample_logic_1_3 _zz_zy_sva_b82 ( _zy_sva_b82, _zy_sva_b82_t);
ixc_sample_logic_1_3 _zz_zy_sva_b83 ( _zy_sva_b83, _zy_sva_b83_t);
ixc_sample_logic_1_3 _zz_zy_sva_b84 ( _zy_sva_b84, _zy_sva_b84_t);
ixc_sample_logic_1_3 _zz_zy_sva_b85 ( _zy_sva_b85, _zy_sva_b85_t);
ixc_sample_logic_1_3 _zz_zy_sva_b86 ( _zy_sva_b86, _zy_sva_b86_t);
ixc_sample_logic_1_3 _zz_zy_sva_b87 ( _zy_sva_b87, _zy_sva_b87_t);
ixc_sample_logic_1_3 _zz_zy_sva_b88 ( _zy_sva_b88, _zy_sva_b88_t);
ixc_sample_logic_1_3 _zz_zy_sva_b89 ( _zy_sva_b89, _zy_sva_b89_t);
ixc_sample_logic_1_3 _zz_zy_sva_b90 ( _zy_sva_b90, _zy_sva_b90_t);
ixc_sample_logic_1_3 _zz_zy_sva_b91 ( _zy_sva_b91, _zy_sva_b91_t);
ixc_sample_logic_1_3 _zz_zy_sva_b92 ( _zy_sva_b92, _zy_sva_b92_t);
ixc_sample_logic_1_3 _zz_zy_sva_b93 ( _zy_sva_b93, _zy_sva_b93_t);
ixc_sample_logic_1_3 _zz_zy_sva_b94 ( _zy_sva_b94, _zy_sva_b94_t);
ixc_sample_logic_1_3 _zz_zy_sva_b95 ( _zy_sva_b95, _zy_sva_b95_t);
ixc_sample_logic_1_3 _zz_zy_sva_b96 ( _zy_sva_b96, _zy_sva_b96_t);
ixc_sample_logic_1_3 _zz_zy_sva_b97 ( _zy_sva_b97, _zy_sva_b97_t);
ixc_sample_logic_1_3 _zz_zy_sva_b98 ( _zy_sva_b98, _zy_sva_b98_t);
ixc_sample_logic_1_3 _zz_zy_sva_b99 ( _zy_sva_b99, _zy_sva_b99_t);
ixc_sample_logic_1_3 _zz_zy_sva_b100 ( _zy_sva_b100, _zy_sva_b100_t);
ixc_sample_logic_1_3 _zz_zy_sva_b101 ( _zy_sva_b101, _zy_sva_b101_t);
ixc_sample_logic_1_3 _zz_zy_sva_b102 ( _zy_sva_b102, _zy_sva_b102_t);
ixc_sample_logic_1_3 _zz_zy_sva_b103 ( _zy_sva_b103, _zy_sva_b103_t);
ixc_sample_logic_1_3 _zz_zy_sva_b104 ( _zy_sva_b104, _zy_sva_b104_t);
ixc_sample_logic_1_3 _zz_zy_sva_b105 ( _zy_sva_b105, _zy_sva_b105_t);
ixc_sample_logic_1_3 _zz_zy_sva_b106 ( _zy_sva_b106, _zy_sva_b106_t);
ixc_sample_logic_1_3 _zz_zy_sva_b107 ( _zy_sva_b107, _zy_sva_b107_t);
ixc_sample_logic_1_3 _zz_zy_sva_b108 ( _zy_sva_b108, _zy_sva_b108_t);
ixc_sample_logic_1_3 _zz_zy_sva_b109 ( _zy_sva_b109, _zy_sva_b109_t);
ixc_sample_logic_1_3 _zz_zy_sva_b110 ( _zy_sva_b110, _zy_sva_b110_t);
ixc_sample_logic_1_3 _zz_zy_sva_b111 ( _zy_sva_b111, _zy_sva_b111_t);
ixc_sample_logic_1_3 _zz_zy_sva_b112 ( _zy_sva_b112, _zy_sva_b112_t);
ixc_sample_logic_1_3 _zz_zy_sva_b113 ( _zy_sva_b113, _zy_sva_b113_t);
ixc_sample_logic_1_3 _zz_zy_sva_b114 ( _zy_sva_b114, _zy_sva_b114_t);
ixc_sample_logic_1_3 _zz_zy_sva_b115 ( _zy_sva_b115, _zy_sva_b115_t);
ixc_sample_logic_1_3 _zz_zy_sva_b116 ( _zy_sva_b116, _zy_sva_b116_t);
ixc_sample_logic_1_3 _zz_zy_sva_b117 ( _zy_sva_b117, _zy_sva_b117_t);
ixc_sample_logic_1_3 _zz_zy_sva_b118 ( _zy_sva_b118, _zy_sva_b118_t);
ixc_sample_logic_1_3 _zz_zy_sva_b119 ( _zy_sva_b119, _zy_sva_b119_t);
ixc_sample_logic_1_3 _zz_zy_sva_b120 ( _zy_sva_b120, _zy_sva_b120_t);
ixc_sample_logic_1_3 _zz_zy_sva_b121 ( _zy_sva_b121, _zy_sva_b121_t);
ixc_sample_logic_1_3 _zz_zy_sva_b122 ( _zy_sva_b122, _zy_sva_b122_t);
ixc_sample_logic_1_3 _zz_zy_sva_b123 ( _zy_sva_b123, _zy_sva_b123_t);
ixc_sample_logic_1_3 _zz_zy_sva_b124 ( _zy_sva_b124, _zy_sva_b124_t);
ixc_sample_logic_1_3 _zz_zy_sva_b125 ( _zy_sva_b125, _zy_sva_b125_t);
ixc_sample_logic_1_3 _zz_zy_sva_b126 ( _zy_sva_b126, _zy_sva_b126_t);
ixc_sample_logic_1_3 _zz_zy_sva_b127 ( _zy_sva_b127, _zy_sva_b127_t);
ixc_sample_logic_1_3 _zz_zy_sva_b128 ( _zy_sva_b128, _zy_sva_b128_t);
ixc_sample_logic_1_3 _zz_zy_sva_b129 ( _zy_sva_b129, _zy_sva_b129_t);
ixc_sample_logic_1_3 _zz_zy_sva_b130 ( _zy_sva_b130, _zy_sva_b130_t);
ixc_sample_logic_1_3 _zz_zy_sva_b131 ( _zy_sva_b131, _zy_sva_b131_t);
ixc_sample_logic_1_3 _zz_zy_sva_b132 ( _zy_sva_b132, _zy_sva_b132_t);
ixc_sample_logic_1_3 _zz_zy_sva_b133 ( _zy_sva_b133, _zy_sva_b133_t);
ixc_sample_logic_1_3 _zz_zy_sva_b134 ( _zy_sva_b134, _zy_sva_b134_t);
ixc_sample_logic_1_3 _zz_zy_sva_b135 ( _zy_sva_b135, _zy_sva_b135_t);
ixc_sample_logic_1_3 _zz_zy_sva_b136 ( _zy_sva_b136, _zy_sva_b136_t);
ixc_sample_logic_1_3 _zz_zy_sva_b137 ( _zy_sva_b137, _zy_sva_b137_t);
ixc_sample_logic_1_3 _zz_zy_sva_b138 ( _zy_sva_b138, _zy_sva_b138_t);
ixc_sample_logic_1_3 _zz_zy_sva_b139 ( _zy_sva_b139, _zy_sva_b139_t);
ixc_sample_logic_1_3 _zz_zy_sva_b140 ( _zy_sva_b140, _zy_sva_b140_t);
ixc_sample_logic_1_3 _zz_zy_sva_b141 ( _zy_sva_b141, _zy_sva_b141_t);
ixc_sample_logic_1_3 _zz_zy_sva_b142 ( _zy_sva_b142, _zy_sva_b142_t);
ixc_sample_logic_1_3 _zz_zy_sva_b143 ( _zy_sva_b143, _zy_sva_b143_t);
ixc_sample_logic_1_3 _zz_zy_sva_b144 ( _zy_sva_b144, _zy_sva_b144_t);
ixc_sample_logic_1_3 _zz_zy_sva_b145 ( _zy_sva_b145, _zy_sva_b145_t);
ixc_sample_logic_1_3 _zz_zy_sva_b146 ( _zy_sva_b146, _zy_sva_b146_t);
ixc_sample_logic_1_3 _zz_zy_sva_b147 ( _zy_sva_b147, _zy_sva_b147_t);
ixc_sample_logic_1_3 _zz_zy_sva_b148 ( _zy_sva_b148, _zy_sva_b148_t);
ixc_sample_logic_1_3 _zz_zy_sva_b149 ( _zy_sva_b149, _zy_sva_b149_t);
ixc_sample_logic_1_3 _zz_zy_sva_b150 ( _zy_sva_b150, _zy_sva_b150_t);
ixc_sample_logic_1_3 _zz_zy_sva_b151 ( _zy_sva_b151, _zy_sva_b151_t);
ixc_sample_logic_1_3 _zz_zy_sva_b152 ( _zy_sva_b152, _zy_sva_b152_t);
ixc_sample_logic_1_3 _zz_zy_sva_b153 ( _zy_sva_b153, _zy_sva_b153_t);
ixc_sample_logic_1_3 _zz_zy_sva_b154 ( _zy_sva_b154, _zy_sva_b154_t);
ixc_sample_logic_1_3 _zz_zy_sva_b155 ( _zy_sva_b155, _zy_sva_b155_t);
ixc_sample_logic_1_3 _zz_zy_sva_b156 ( _zy_sva_b156, _zy_sva_b156_t);
ixc_sample_logic_1_3 _zz_zy_sva_b157 ( _zy_sva_b157, _zy_sva_b157_t);
ixc_sample_logic_1_3 _zz_zy_sva_b158 ( _zy_sva_b158, _zy_sva_b158_t);
ixc_sample_logic_1_3 _zz_zy_sva_b159 ( _zy_sva_b159, _zy_sva_b159_t);
ixc_sample_logic_1_3 _zz_zy_sva_b160 ( _zy_sva_b160, _zy_sva_b160_t);
ixc_sample_logic_1_3 _zz_zy_sva_b161 ( _zy_sva_b161, _zy_sva_b161_t);
ixc_sample_logic_1_3 _zz_zy_sva_b162 ( _zy_sva_b162, _zy_sva_b162_t);
ixc_sample_logic_1_3 _zz_zy_sva_b163 ( _zy_sva_b163, _zy_sva_b163_t);
ixc_sample_logic_1_3 _zz_zy_sva_b164 ( _zy_sva_b164, _zy_sva_b164_t);
ixc_sample_logic_1_3 _zz_zy_sva_b165 ( _zy_sva_b165, _zy_sva_b165_t);
ixc_sample_logic_1_3 _zz_zy_sva_b166 ( _zy_sva_b166, _zy_sva_b166_t);
ixc_sample_logic_1_3 _zz_zy_sva_b167 ( _zy_sva_b167, _zy_sva_b167_t);
ixc_sample_logic_1_3 _zz_zy_sva_b168 ( _zy_sva_b168, _zy_sva_b168_t);
ixc_sample_logic_1_3 _zz_zy_sva_b169 ( _zy_sva_b169, _zy_sva_b169_t);
ixc_sample_logic_1_3 _zz_zy_sva_b170 ( _zy_sva_b170, _zy_sva_b170_t);
ixc_sample_logic_1_3 _zz_zy_sva_b171 ( _zy_sva_b171, _zy_sva_b171_t);
ixc_sample_logic_1_3 _zz_zy_sva_b172 ( _zy_sva_b172, _zy_sva_b172_t);
ixc_sample_logic_1_3 _zz_zy_sva_b173 ( _zy_sva_b173, _zy_sva_b173_t);
ixc_sample_logic_1_3 _zz_zy_sva_b174 ( _zy_sva_b174, _zy_sva_b174_t);
ixc_sample_logic_1_3 _zz_zy_sva_b175 ( _zy_sva_b175, _zy_sva_b175_t);
ixc_sample_logic_1_3 _zz_zy_sva_b176 ( _zy_sva_b176, _zy_sva_b176_t);
ixc_sample_logic_1_3 _zz_zy_sva_b177 ( _zy_sva_b177, _zy_sva_b177_t);
cr_kme_fifo_xcm57 parser_fifo ( .fifo_in_stall( fifo_in_stall), .fifo_out( 
	_zy_simnet_parser_kimreader_data_2_w$[0:70]), .fifo_out_valid( 
	parser_kimreader_valid), .fifo_overflow( _zy_simnet_dio_3), 
	.fifo_underflow( _zy_simnet_dio_4), .clk( clk), .rst_n( rst_n), 
	.fifo_in( _zy_simnet_fifo_in_5_w$[0:70]), .fifo_in_valid( 
	_zy_simnet_fifo_in_valid_6_w$), .fifo_out_ack( kimreader_parser_ack), 
	.fifo_in_stall_override( _zy_simnet_cio_7));
wire [2:0] n2147 = 3'b000;
Q_ASSERT \key_type_0_.brcm_aux_cmd  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_39_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_39_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2147[0]));
// pragma CVASTRPROP INSTANCE "\key_type_0_.brcm_aux_cmd " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_0_.brcm_aux_cmd " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_0_.brcm_aux_cmd " ASSERT_LINE 889
wire [2:0] n2148 = 3'b000;
Q_ASSERT \key_type_0_.brcm_aux_cmd_iv  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_iv_40_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_iv_40_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2148[0]));
// pragma CVASTRPROP INSTANCE "\key_type_0_.brcm_aux_cmd_iv " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_0_.brcm_aux_cmd_iv " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_0_.brcm_aux_cmd_iv " ASSERT_LINE 890
wire [2:0] n2149 = 3'b000;
Q_ASSERT \key_type_0_.brcm_aux_cmd_guid  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_guid_41_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_guid_41_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2149[0]));
// pragma CVASTRPROP INSTANCE "\key_type_0_.brcm_aux_cmd_guid " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_0_.brcm_aux_cmd_guid " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_0_.brcm_aux_cmd_guid " ASSERT_LINE 891
wire [2:0] n2150 = 3'b000;
Q_ASSERT \key_type_0_.brcm_aux_cmd_guid_iv  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_guid_iv_42_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_guid_iv_42_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2150[0]));
// pragma CVASTRPROP INSTANCE "\key_type_0_.brcm_aux_cmd_guid_iv " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_0_.brcm_aux_cmd_guid_iv " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_0_.brcm_aux_cmd_guid_iv " ASSERT_LINE 892
wire [2:0] n2151 = 3'b000;
Q_ASSERT \key_type_0_.brcm_key_type  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_key_type_43_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_key_type_43_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2151[0]));
// pragma CVASTRPROP INSTANCE "\key_type_0_.brcm_key_type " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_0_.brcm_key_type " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_0_.brcm_key_type " ASSERT_LINE 893
wire [2:0] n2152 = 3'b000;
Q_ASSERT \key_type_1_.brcm_aux_cmd  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_44_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_44_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2152[0]));
// pragma CVASTRPROP INSTANCE "\key_type_1_.brcm_aux_cmd " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_1_.brcm_aux_cmd " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_1_.brcm_aux_cmd " ASSERT_LINE 889
wire [2:0] n2153 = 3'b000;
Q_ASSERT \key_type_1_.brcm_aux_cmd_iv  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_iv_45_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_iv_45_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2153[0]));
// pragma CVASTRPROP INSTANCE "\key_type_1_.brcm_aux_cmd_iv " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_1_.brcm_aux_cmd_iv " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_1_.brcm_aux_cmd_iv " ASSERT_LINE 890
wire [2:0] n2154 = 3'b000;
Q_ASSERT \key_type_1_.brcm_aux_cmd_guid  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_guid_46_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_guid_46_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2154[0]));
// pragma CVASTRPROP INSTANCE "\key_type_1_.brcm_aux_cmd_guid " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_1_.brcm_aux_cmd_guid " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_1_.brcm_aux_cmd_guid " ASSERT_LINE 891
wire [2:0] n2155 = 3'b000;
Q_ASSERT \key_type_1_.brcm_aux_cmd_guid_iv  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_guid_iv_47_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_guid_iv_47_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2155[0]));
// pragma CVASTRPROP INSTANCE "\key_type_1_.brcm_aux_cmd_guid_iv " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_1_.brcm_aux_cmd_guid_iv " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_1_.brcm_aux_cmd_guid_iv " ASSERT_LINE 892
wire [2:0] n2156 = 3'b000;
Q_ASSERT \key_type_1_.brcm_key_type  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_key_type_48_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_key_type_48_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2156[0]));
// pragma CVASTRPROP INSTANCE "\key_type_1_.brcm_key_type " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_1_.brcm_key_type " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_1_.brcm_key_type " ASSERT_LINE 893
wire [2:0] n2157 = 3'b000;
Q_ASSERT \key_type_2_.brcm_aux_cmd  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_49_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_49_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2157[0]));
// pragma CVASTRPROP INSTANCE "\key_type_2_.brcm_aux_cmd " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_2_.brcm_aux_cmd " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_2_.brcm_aux_cmd " ASSERT_LINE 889
wire [2:0] n2158 = 3'b000;
Q_ASSERT \key_type_2_.brcm_aux_cmd_iv  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_iv_50_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_iv_50_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2158[0]));
// pragma CVASTRPROP INSTANCE "\key_type_2_.brcm_aux_cmd_iv " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_2_.brcm_aux_cmd_iv " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_2_.brcm_aux_cmd_iv " ASSERT_LINE 890
wire [2:0] n2159 = 3'b000;
Q_ASSERT \key_type_2_.brcm_aux_cmd_guid  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_guid_51_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_guid_51_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2159[0]));
// pragma CVASTRPROP INSTANCE "\key_type_2_.brcm_aux_cmd_guid " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_2_.brcm_aux_cmd_guid " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_2_.brcm_aux_cmd_guid " ASSERT_LINE 891
wire [2:0] n2160 = 3'b000;
Q_ASSERT \key_type_2_.brcm_aux_cmd_guid_iv  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_guid_iv_52_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_guid_iv_52_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2160[0]));
// pragma CVASTRPROP INSTANCE "\key_type_2_.brcm_aux_cmd_guid_iv " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_2_.brcm_aux_cmd_guid_iv " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_2_.brcm_aux_cmd_guid_iv " ASSERT_LINE 892
wire [2:0] n2161 = 3'b000;
Q_ASSERT \key_type_2_.brcm_key_type  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_key_type_53_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_key_type_53_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2161[0]));
// pragma CVASTRPROP INSTANCE "\key_type_2_.brcm_key_type " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_2_.brcm_key_type " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_2_.brcm_key_type " ASSERT_LINE 893
wire [2:0] n2162 = 3'b000;
Q_ASSERT \key_type_3_.brcm_aux_cmd  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_54_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_54_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2162[0]));
// pragma CVASTRPROP INSTANCE "\key_type_3_.brcm_aux_cmd " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_3_.brcm_aux_cmd " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_3_.brcm_aux_cmd " ASSERT_LINE 889
wire [2:0] n2163 = 3'b000;
Q_ASSERT \key_type_3_.brcm_aux_cmd_iv  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_iv_55_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_iv_55_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2163[0]));
// pragma CVASTRPROP INSTANCE "\key_type_3_.brcm_aux_cmd_iv " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_3_.brcm_aux_cmd_iv " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_3_.brcm_aux_cmd_iv " ASSERT_LINE 890
wire [2:0] n2164 = 3'b000;
Q_ASSERT \key_type_3_.brcm_aux_cmd_guid  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_guid_56_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_guid_56_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2164[0]));
// pragma CVASTRPROP INSTANCE "\key_type_3_.brcm_aux_cmd_guid " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_3_.brcm_aux_cmd_guid " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_3_.brcm_aux_cmd_guid " ASSERT_LINE 891
wire [2:0] n2165 = 3'b000;
Q_ASSERT \key_type_3_.brcm_aux_cmd_guid_iv  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_guid_iv_57_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_guid_iv_57_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2165[0]));
// pragma CVASTRPROP INSTANCE "\key_type_3_.brcm_aux_cmd_guid_iv " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_3_.brcm_aux_cmd_guid_iv " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_3_.brcm_aux_cmd_guid_iv " ASSERT_LINE 892
wire [2:0] n2166 = 3'b000;
Q_ASSERT \key_type_3_.brcm_key_type  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_key_type_58_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_key_type_58_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2166[0]));
// pragma CVASTRPROP INSTANCE "\key_type_3_.brcm_key_type " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_3_.brcm_key_type " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_3_.brcm_key_type " ASSERT_LINE 893
wire [2:0] n2167 = 3'b000;
Q_ASSERT \key_type_4_.brcm_aux_cmd  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_59_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_59_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2167[0]));
// pragma CVASTRPROP INSTANCE "\key_type_4_.brcm_aux_cmd " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_4_.brcm_aux_cmd " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_4_.brcm_aux_cmd " ASSERT_LINE 889
wire [2:0] n2168 = 3'b000;
Q_ASSERT \key_type_4_.brcm_aux_cmd_iv  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_iv_60_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_iv_60_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2168[0]));
// pragma CVASTRPROP INSTANCE "\key_type_4_.brcm_aux_cmd_iv " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_4_.brcm_aux_cmd_iv " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_4_.brcm_aux_cmd_iv " ASSERT_LINE 890
wire [2:0] n2169 = 3'b000;
Q_ASSERT \key_type_4_.brcm_aux_cmd_guid  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_guid_61_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_guid_61_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2169[0]));
// pragma CVASTRPROP INSTANCE "\key_type_4_.brcm_aux_cmd_guid " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_4_.brcm_aux_cmd_guid " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_4_.brcm_aux_cmd_guid " ASSERT_LINE 891
wire [2:0] n2170 = 3'b000;
Q_ASSERT \key_type_4_.brcm_aux_cmd_guid_iv  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_guid_iv_62_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_guid_iv_62_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2170[0]));
// pragma CVASTRPROP INSTANCE "\key_type_4_.brcm_aux_cmd_guid_iv " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_4_.brcm_aux_cmd_guid_iv " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_4_.brcm_aux_cmd_guid_iv " ASSERT_LINE 892
wire [2:0] n2171 = 3'b000;
Q_ASSERT \key_type_4_.brcm_key_type  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_key_type_63_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_key_type_63_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2171[0]));
// pragma CVASTRPROP INSTANCE "\key_type_4_.brcm_key_type " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_4_.brcm_key_type " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_4_.brcm_key_type " ASSERT_LINE 893
wire [2:0] n2172 = 3'b000;
Q_ASSERT \key_type_5_.brcm_aux_cmd  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_64_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_64_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2172[0]));
// pragma CVASTRPROP INSTANCE "\key_type_5_.brcm_aux_cmd " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_5_.brcm_aux_cmd " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_5_.brcm_aux_cmd " ASSERT_LINE 889
wire [2:0] n2173 = 3'b000;
Q_ASSERT \key_type_5_.brcm_aux_cmd_iv  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_iv_65_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_iv_65_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2173[0]));
// pragma CVASTRPROP INSTANCE "\key_type_5_.brcm_aux_cmd_iv " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_5_.brcm_aux_cmd_iv " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_5_.brcm_aux_cmd_iv " ASSERT_LINE 890
wire [2:0] n2174 = 3'b000;
Q_ASSERT \key_type_5_.brcm_aux_cmd_guid  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_guid_66_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_guid_66_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2174[0]));
// pragma CVASTRPROP INSTANCE "\key_type_5_.brcm_aux_cmd_guid " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_5_.brcm_aux_cmd_guid " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_5_.brcm_aux_cmd_guid " ASSERT_LINE 891
wire [2:0] n2175 = 3'b000;
Q_ASSERT \key_type_5_.brcm_aux_cmd_guid_iv  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_guid_iv_67_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_guid_iv_67_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2175[0]));
// pragma CVASTRPROP INSTANCE "\key_type_5_.brcm_aux_cmd_guid_iv " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_5_.brcm_aux_cmd_guid_iv " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_5_.brcm_aux_cmd_guid_iv " ASSERT_LINE 892
wire [2:0] n2176 = 3'b000;
Q_ASSERT \key_type_5_.brcm_key_type  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_key_type_68_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_key_type_68_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2176[0]));
// pragma CVASTRPROP INSTANCE "\key_type_5_.brcm_key_type " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_5_.brcm_key_type " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_5_.brcm_key_type " ASSERT_LINE 893
wire [2:0] n2177 = 3'b000;
Q_ASSERT \key_type_6_.brcm_aux_cmd  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_69_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_69_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2177[0]));
// pragma CVASTRPROP INSTANCE "\key_type_6_.brcm_aux_cmd " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_6_.brcm_aux_cmd " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_6_.brcm_aux_cmd " ASSERT_LINE 889
wire [2:0] n2178 = 3'b000;
Q_ASSERT \key_type_6_.brcm_aux_cmd_iv  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_iv_70_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_iv_70_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2178[0]));
// pragma CVASTRPROP INSTANCE "\key_type_6_.brcm_aux_cmd_iv " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_6_.brcm_aux_cmd_iv " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_6_.brcm_aux_cmd_iv " ASSERT_LINE 890
wire [2:0] n2179 = 3'b000;
Q_ASSERT \key_type_6_.brcm_aux_cmd_guid  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_guid_71_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_guid_71_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2179[0]));
// pragma CVASTRPROP INSTANCE "\key_type_6_.brcm_aux_cmd_guid " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_6_.brcm_aux_cmd_guid " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_6_.brcm_aux_cmd_guid " ASSERT_LINE 891
wire [2:0] n2180 = 3'b000;
Q_ASSERT \key_type_6_.brcm_aux_cmd_guid_iv  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_guid_iv_72_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_guid_iv_72_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2180[0]));
// pragma CVASTRPROP INSTANCE "\key_type_6_.brcm_aux_cmd_guid_iv " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_6_.brcm_aux_cmd_guid_iv " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_6_.brcm_aux_cmd_guid_iv " ASSERT_LINE 892
wire [2:0] n2181 = 3'b000;
Q_ASSERT \key_type_6_.brcm_key_type  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_key_type_73_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_key_type_73_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2181[0]));
// pragma CVASTRPROP INSTANCE "\key_type_6_.brcm_key_type " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_6_.brcm_key_type " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_6_.brcm_key_type " ASSERT_LINE 893
wire [2:0] n2182 = 3'b000;
Q_ASSERT \key_type_7_.brcm_aux_cmd  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_74_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_74_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2182[0]));
// pragma CVASTRPROP INSTANCE "\key_type_7_.brcm_aux_cmd " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_7_.brcm_aux_cmd " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_7_.brcm_aux_cmd " ASSERT_LINE 889
wire [2:0] n2183 = 3'b000;
Q_ASSERT \key_type_7_.brcm_aux_cmd_iv  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_iv_75_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_iv_75_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2183[0]));
// pragma CVASTRPROP INSTANCE "\key_type_7_.brcm_aux_cmd_iv " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_7_.brcm_aux_cmd_iv " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_7_.brcm_aux_cmd_iv " ASSERT_LINE 890
wire [2:0] n2184 = 3'b000;
Q_ASSERT \key_type_7_.brcm_aux_cmd_guid  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_guid_76_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_guid_76_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2184[0]));
// pragma CVASTRPROP INSTANCE "\key_type_7_.brcm_aux_cmd_guid " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_7_.brcm_aux_cmd_guid " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_7_.brcm_aux_cmd_guid " ASSERT_LINE 891
wire [2:0] n2185 = 3'b000;
Q_ASSERT \key_type_7_.brcm_aux_cmd_guid_iv  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_guid_iv_77_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_guid_iv_77_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2185[0]));
// pragma CVASTRPROP INSTANCE "\key_type_7_.brcm_aux_cmd_guid_iv " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_7_.brcm_aux_cmd_guid_iv " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_7_.brcm_aux_cmd_guid_iv " ASSERT_LINE 892
wire [2:0] n2186 = 3'b000;
Q_ASSERT \key_type_7_.brcm_key_type  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_key_type_78_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_key_type_78_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2186[0]));
// pragma CVASTRPROP INSTANCE "\key_type_7_.brcm_key_type " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_7_.brcm_key_type " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_7_.brcm_key_type " ASSERT_LINE 893
wire [2:0] n2187 = 3'b000;
Q_ASSERT \key_type_8_.brcm_aux_cmd  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_79_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_79_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2187[0]));
// pragma CVASTRPROP INSTANCE "\key_type_8_.brcm_aux_cmd " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_8_.brcm_aux_cmd " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_8_.brcm_aux_cmd " ASSERT_LINE 889
wire [2:0] n2188 = 3'b000;
Q_ASSERT \key_type_8_.brcm_aux_cmd_iv  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_iv_80_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_iv_80_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2188[0]));
// pragma CVASTRPROP INSTANCE "\key_type_8_.brcm_aux_cmd_iv " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_8_.brcm_aux_cmd_iv " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_8_.brcm_aux_cmd_iv " ASSERT_LINE 890
wire [2:0] n2189 = 3'b000;
Q_ASSERT \key_type_8_.brcm_aux_cmd_guid  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_guid_81_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_guid_81_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2189[0]));
// pragma CVASTRPROP INSTANCE "\key_type_8_.brcm_aux_cmd_guid " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_8_.brcm_aux_cmd_guid " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_8_.brcm_aux_cmd_guid " ASSERT_LINE 891
wire [2:0] n2190 = 3'b000;
Q_ASSERT \key_type_8_.brcm_aux_cmd_guid_iv  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_guid_iv_82_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_guid_iv_82_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2190[0]));
// pragma CVASTRPROP INSTANCE "\key_type_8_.brcm_aux_cmd_guid_iv " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_8_.brcm_aux_cmd_guid_iv " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_8_.brcm_aux_cmd_guid_iv " ASSERT_LINE 892
wire [2:0] n2191 = 3'b000;
Q_ASSERT \key_type_8_.brcm_key_type  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_key_type_83_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_key_type_83_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2191[0]));
// pragma CVASTRPROP INSTANCE "\key_type_8_.brcm_key_type " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_8_.brcm_key_type " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_8_.brcm_key_type " ASSERT_LINE 893
wire [2:0] n2192 = 3'b000;
Q_ASSERT \key_type_9_.brcm_aux_cmd  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_84_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_84_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2192[0]));
// pragma CVASTRPROP INSTANCE "\key_type_9_.brcm_aux_cmd " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_9_.brcm_aux_cmd " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_9_.brcm_aux_cmd " ASSERT_LINE 889
wire [2:0] n2193 = 3'b000;
Q_ASSERT \key_type_9_.brcm_aux_cmd_iv  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_iv_85_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_iv_85_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2193[0]));
// pragma CVASTRPROP INSTANCE "\key_type_9_.brcm_aux_cmd_iv " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_9_.brcm_aux_cmd_iv " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_9_.brcm_aux_cmd_iv " ASSERT_LINE 890
wire [2:0] n2194 = 3'b000;
Q_ASSERT \key_type_9_.brcm_aux_cmd_guid  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_guid_86_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_guid_86_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2194[0]));
// pragma CVASTRPROP INSTANCE "\key_type_9_.brcm_aux_cmd_guid " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_9_.brcm_aux_cmd_guid " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_9_.brcm_aux_cmd_guid " ASSERT_LINE 891
wire [2:0] n2195 = 3'b000;
Q_ASSERT \key_type_9_.brcm_aux_cmd_guid_iv  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_guid_iv_87_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_guid_iv_87_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2195[0]));
// pragma CVASTRPROP INSTANCE "\key_type_9_.brcm_aux_cmd_guid_iv " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_9_.brcm_aux_cmd_guid_iv " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_9_.brcm_aux_cmd_guid_iv " ASSERT_LINE 892
wire [2:0] n2196 = 3'b000;
Q_ASSERT \key_type_9_.brcm_key_type  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_key_type_88_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_key_type_88_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2196[0]));
// pragma CVASTRPROP INSTANCE "\key_type_9_.brcm_key_type " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_9_.brcm_key_type " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_9_.brcm_key_type " ASSERT_LINE 893
wire [2:0] n2197 = 3'b000;
Q_ASSERT \key_type_10_.brcm_aux_cmd  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_89_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_89_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2197[0]));
// pragma CVASTRPROP INSTANCE "\key_type_10_.brcm_aux_cmd " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_10_.brcm_aux_cmd " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_10_.brcm_aux_cmd " ASSERT_LINE 889
wire [2:0] n2198 = 3'b000;
Q_ASSERT \key_type_10_.brcm_aux_cmd_iv  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_iv_90_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_iv_90_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2198[0]));
// pragma CVASTRPROP INSTANCE "\key_type_10_.brcm_aux_cmd_iv " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_10_.brcm_aux_cmd_iv " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_10_.brcm_aux_cmd_iv " ASSERT_LINE 890
wire [2:0] n2199 = 3'b000;
Q_ASSERT \key_type_10_.brcm_aux_cmd_guid  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_guid_91_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_guid_91_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2199[0]));
// pragma CVASTRPROP INSTANCE "\key_type_10_.brcm_aux_cmd_guid " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_10_.brcm_aux_cmd_guid " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_10_.brcm_aux_cmd_guid " ASSERT_LINE 891
wire [2:0] n2200 = 3'b000;
Q_ASSERT \key_type_10_.brcm_aux_cmd_guid_iv  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_guid_iv_92_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_guid_iv_92_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2200[0]));
// pragma CVASTRPROP INSTANCE "\key_type_10_.brcm_aux_cmd_guid_iv " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_10_.brcm_aux_cmd_guid_iv " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_10_.brcm_aux_cmd_guid_iv " ASSERT_LINE 892
wire [2:0] n2201 = 3'b000;
Q_ASSERT \key_type_10_.brcm_key_type  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_key_type_93_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_key_type_93_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2201[0]));
// pragma CVASTRPROP INSTANCE "\key_type_10_.brcm_key_type " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_10_.brcm_key_type " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_10_.brcm_key_type " ASSERT_LINE 893
wire [2:0] n2202 = 3'b000;
Q_ASSERT \key_type_11_.brcm_aux_cmd  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_94_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_94_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2202[0]));
// pragma CVASTRPROP INSTANCE "\key_type_11_.brcm_aux_cmd " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_11_.brcm_aux_cmd " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_11_.brcm_aux_cmd " ASSERT_LINE 889
wire [2:0] n2203 = 3'b000;
Q_ASSERT \key_type_11_.brcm_aux_cmd_iv  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_iv_95_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_iv_95_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2203[0]));
// pragma CVASTRPROP INSTANCE "\key_type_11_.brcm_aux_cmd_iv " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_11_.brcm_aux_cmd_iv " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_11_.brcm_aux_cmd_iv " ASSERT_LINE 890
wire [2:0] n2204 = 3'b000;
Q_ASSERT \key_type_11_.brcm_aux_cmd_guid  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_guid_96_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_guid_96_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2204[0]));
// pragma CVASTRPROP INSTANCE "\key_type_11_.brcm_aux_cmd_guid " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_11_.brcm_aux_cmd_guid " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_11_.brcm_aux_cmd_guid " ASSERT_LINE 891
wire [2:0] n2205 = 3'b000;
Q_ASSERT \key_type_11_.brcm_aux_cmd_guid_iv  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_guid_iv_97_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_guid_iv_97_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2205[0]));
// pragma CVASTRPROP INSTANCE "\key_type_11_.brcm_aux_cmd_guid_iv " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_11_.brcm_aux_cmd_guid_iv " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_11_.brcm_aux_cmd_guid_iv " ASSERT_LINE 892
wire [2:0] n2206 = 3'b000;
Q_ASSERT \key_type_11_.brcm_key_type  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_key_type_98_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_key_type_98_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2206[0]));
// pragma CVASTRPROP INSTANCE "\key_type_11_.brcm_key_type " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_11_.brcm_key_type " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_11_.brcm_key_type " ASSERT_LINE 893
wire [2:0] n2207 = 3'b000;
Q_ASSERT \key_type_12_.brcm_aux_cmd  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_99_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_99_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2207[0]));
// pragma CVASTRPROP INSTANCE "\key_type_12_.brcm_aux_cmd " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_12_.brcm_aux_cmd " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_12_.brcm_aux_cmd " ASSERT_LINE 889
wire [2:0] n2208 = 3'b000;
Q_ASSERT \key_type_12_.brcm_aux_cmd_iv  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_iv_100_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_iv_100_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2208[0]));
// pragma CVASTRPROP INSTANCE "\key_type_12_.brcm_aux_cmd_iv " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_12_.brcm_aux_cmd_iv " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_12_.brcm_aux_cmd_iv " ASSERT_LINE 890
wire [2:0] n2209 = 3'b000;
Q_ASSERT \key_type_12_.brcm_aux_cmd_guid  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_guid_101_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_guid_101_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2209[0]));
// pragma CVASTRPROP INSTANCE "\key_type_12_.brcm_aux_cmd_guid " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_12_.brcm_aux_cmd_guid " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_12_.brcm_aux_cmd_guid " ASSERT_LINE 891
wire [2:0] n2210 = 3'b000;
Q_ASSERT \key_type_12_.brcm_aux_cmd_guid_iv  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_guid_iv_102_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_guid_iv_102_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2210[0]));
// pragma CVASTRPROP INSTANCE "\key_type_12_.brcm_aux_cmd_guid_iv " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_12_.brcm_aux_cmd_guid_iv " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_12_.brcm_aux_cmd_guid_iv " ASSERT_LINE 892
wire [2:0] n2211 = 3'b000;
Q_ASSERT \key_type_12_.brcm_key_type  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_key_type_103_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_key_type_103_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2211[0]));
// pragma CVASTRPROP INSTANCE "\key_type_12_.brcm_key_type " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_12_.brcm_key_type " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_12_.brcm_key_type " ASSERT_LINE 893
wire [2:0] n2212 = 3'b000;
Q_ASSERT \key_type_13_.brcm_aux_cmd  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_104_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_104_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2212[0]));
// pragma CVASTRPROP INSTANCE "\key_type_13_.brcm_aux_cmd " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_13_.brcm_aux_cmd " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_13_.brcm_aux_cmd " ASSERT_LINE 889
wire [2:0] n2213 = 3'b000;
Q_ASSERT \key_type_13_.brcm_aux_cmd_iv  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_iv_105_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_iv_105_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2213[0]));
// pragma CVASTRPROP INSTANCE "\key_type_13_.brcm_aux_cmd_iv " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_13_.brcm_aux_cmd_iv " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_13_.brcm_aux_cmd_iv " ASSERT_LINE 890
wire [2:0] n2214 = 3'b000;
Q_ASSERT \key_type_13_.brcm_aux_cmd_guid  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_guid_106_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_guid_106_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2214[0]));
// pragma CVASTRPROP INSTANCE "\key_type_13_.brcm_aux_cmd_guid " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_13_.brcm_aux_cmd_guid " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_13_.brcm_aux_cmd_guid " ASSERT_LINE 891
wire [2:0] n2215 = 3'b000;
Q_ASSERT \key_type_13_.brcm_aux_cmd_guid_iv  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_aux_cmd_guid_iv_107_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_aux_cmd_guid_iv_107_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2215[0]));
// pragma CVASTRPROP INSTANCE "\key_type_13_.brcm_aux_cmd_guid_iv " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_13_.brcm_aux_cmd_guid_iv " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_13_.brcm_aux_cmd_guid_iv " ASSERT_LINE 892
wire [2:0] n2216 = 3'b000;
Q_ASSERT \key_type_13_.brcm_key_type  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_key_type_108_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_key_type_108_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2216[0]));
// pragma CVASTRPROP INSTANCE "\key_type_13_.brcm_key_type " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_13_.brcm_key_type " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_13_.brcm_key_type " ASSERT_LINE 893
wire [2:0] n2217 = 3'b000;
Q_ASSERT \kdf_mode_0_.dek_op_0_.dak_op_0_.brcm_kdf_ops  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_ops_109_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_ops_109_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2217[0]));
// pragma CVASTRPROP INSTANCE "\kdf_mode_0_.dek_op_0_.dak_op_0_.brcm_kdf_ops " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\kdf_mode_0_.dek_op_0_.dak_op_0_.brcm_kdf_ops " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\kdf_mode_0_.dek_op_0_.dak_op_0_.brcm_kdf_ops " ASSERT_LINE 902
wire [2:0] n2218 = 3'b000;
Q_ASSERT \kdf_mode_0_.dek_op_0_.dak_op_1_.brcm_kdf_ops  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_ops_110_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_ops_110_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2218[0]));
// pragma CVASTRPROP INSTANCE "\kdf_mode_0_.dek_op_0_.dak_op_1_.brcm_kdf_ops " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\kdf_mode_0_.dek_op_0_.dak_op_1_.brcm_kdf_ops " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\kdf_mode_0_.dek_op_0_.dak_op_1_.brcm_kdf_ops " ASSERT_LINE 902
wire [2:0] n2219 = 3'b000;
Q_ASSERT \kdf_mode_0_.dek_op_1_.dak_op_0_.brcm_kdf_ops  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_ops_111_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_ops_111_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2219[0]));
// pragma CVASTRPROP INSTANCE "\kdf_mode_0_.dek_op_1_.dak_op_0_.brcm_kdf_ops " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\kdf_mode_0_.dek_op_1_.dak_op_0_.brcm_kdf_ops " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\kdf_mode_0_.dek_op_1_.dak_op_0_.brcm_kdf_ops " ASSERT_LINE 902
wire [2:0] n2220 = 3'b000;
Q_ASSERT \kdf_mode_0_.dek_op_1_.dak_op_1_.brcm_kdf_ops  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_ops_112_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_ops_112_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2220[0]));
// pragma CVASTRPROP INSTANCE "\kdf_mode_0_.dek_op_1_.dak_op_1_.brcm_kdf_ops " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\kdf_mode_0_.dek_op_1_.dak_op_1_.brcm_kdf_ops " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\kdf_mode_0_.dek_op_1_.dak_op_1_.brcm_kdf_ops " ASSERT_LINE 902
wire [2:0] n2221 = 3'b000;
Q_ASSERT \kdf_mode_1_.dek_op_0_.dak_op_0_.brcm_kdf_ops  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_ops_113_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_ops_113_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2221[0]));
// pragma CVASTRPROP INSTANCE "\kdf_mode_1_.dek_op_0_.dak_op_0_.brcm_kdf_ops " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\kdf_mode_1_.dek_op_0_.dak_op_0_.brcm_kdf_ops " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\kdf_mode_1_.dek_op_0_.dak_op_0_.brcm_kdf_ops " ASSERT_LINE 902
wire [2:0] n2222 = 3'b000;
Q_ASSERT \kdf_mode_1_.dek_op_0_.dak_op_1_.brcm_kdf_ops  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_ops_114_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_ops_114_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2222[0]));
// pragma CVASTRPROP INSTANCE "\kdf_mode_1_.dek_op_0_.dak_op_1_.brcm_kdf_ops " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\kdf_mode_1_.dek_op_0_.dak_op_1_.brcm_kdf_ops " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\kdf_mode_1_.dek_op_0_.dak_op_1_.brcm_kdf_ops " ASSERT_LINE 902
wire [2:0] n2223 = 3'b000;
Q_ASSERT \kdf_mode_1_.dek_op_1_.dak_op_0_.brcm_kdf_ops  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_ops_115_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_ops_115_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2223[0]));
// pragma CVASTRPROP INSTANCE "\kdf_mode_1_.dek_op_1_.dak_op_0_.brcm_kdf_ops " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\kdf_mode_1_.dek_op_1_.dak_op_0_.brcm_kdf_ops " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\kdf_mode_1_.dek_op_1_.dak_op_0_.brcm_kdf_ops " ASSERT_LINE 902
wire [2:0] n2224 = 3'b000;
Q_ASSERT \kdf_mode_1_.dek_op_1_.dak_op_1_.brcm_kdf_ops  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_ops_116_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_ops_116_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2224[0]));
// pragma CVASTRPROP INSTANCE "\kdf_mode_1_.dek_op_1_.dak_op_1_.brcm_kdf_ops " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\kdf_mode_1_.dek_op_1_.dak_op_1_.brcm_kdf_ops " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\kdf_mode_1_.dek_op_1_.dak_op_1_.brcm_kdf_ops " ASSERT_LINE 902
wire [2:0] n2225 = 3'b000;
Q_ASSERT \kdf_mode_2_.dek_op_0_.dak_op_0_.brcm_kdf_ops  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_ops_117_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_ops_117_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2225[0]));
// pragma CVASTRPROP INSTANCE "\kdf_mode_2_.dek_op_0_.dak_op_0_.brcm_kdf_ops " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\kdf_mode_2_.dek_op_0_.dak_op_0_.brcm_kdf_ops " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\kdf_mode_2_.dek_op_0_.dak_op_0_.brcm_kdf_ops " ASSERT_LINE 902
wire [2:0] n2226 = 3'b000;
Q_ASSERT \kdf_mode_2_.dek_op_0_.dak_op_1_.brcm_kdf_ops  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_ops_118_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_ops_118_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2226[0]));
// pragma CVASTRPROP INSTANCE "\kdf_mode_2_.dek_op_0_.dak_op_1_.brcm_kdf_ops " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\kdf_mode_2_.dek_op_0_.dak_op_1_.brcm_kdf_ops " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\kdf_mode_2_.dek_op_0_.dak_op_1_.brcm_kdf_ops " ASSERT_LINE 902
wire [2:0] n2227 = 3'b000;
Q_ASSERT \kdf_mode_2_.dek_op_1_.dak_op_0_.brcm_kdf_ops  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_ops_119_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_ops_119_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2227[0]));
// pragma CVASTRPROP INSTANCE "\kdf_mode_2_.dek_op_1_.dak_op_0_.brcm_kdf_ops " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\kdf_mode_2_.dek_op_1_.dak_op_0_.brcm_kdf_ops " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\kdf_mode_2_.dek_op_1_.dak_op_0_.brcm_kdf_ops " ASSERT_LINE 902
wire [2:0] n2228 = 3'b000;
Q_ASSERT \kdf_mode_2_.dek_op_1_.dak_op_1_.brcm_kdf_ops  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_ops_120_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_ops_120_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2228[0]));
// pragma CVASTRPROP INSTANCE "\kdf_mode_2_.dek_op_1_.dak_op_1_.brcm_kdf_ops " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\kdf_mode_2_.dek_op_1_.dak_op_1_.brcm_kdf_ops " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\kdf_mode_2_.dek_op_1_.dak_op_1_.brcm_kdf_ops " ASSERT_LINE 902
wire [2:0] n2229 = 3'b000;
Q_ASSERT \kdf_mode_3_.dek_op_0_.dak_op_0_.brcm_kdf_ops  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_ops_121_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_ops_121_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2229[0]));
// pragma CVASTRPROP INSTANCE "\kdf_mode_3_.dek_op_0_.dak_op_0_.brcm_kdf_ops " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\kdf_mode_3_.dek_op_0_.dak_op_0_.brcm_kdf_ops " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\kdf_mode_3_.dek_op_0_.dak_op_0_.brcm_kdf_ops " ASSERT_LINE 902
wire [2:0] n2230 = 3'b000;
Q_ASSERT \kdf_mode_3_.dek_op_0_.dak_op_1_.brcm_kdf_ops  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_ops_122_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_ops_122_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2230[0]));
// pragma CVASTRPROP INSTANCE "\kdf_mode_3_.dek_op_0_.dak_op_1_.brcm_kdf_ops " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\kdf_mode_3_.dek_op_0_.dak_op_1_.brcm_kdf_ops " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\kdf_mode_3_.dek_op_0_.dak_op_1_.brcm_kdf_ops " ASSERT_LINE 902
wire [2:0] n2231 = 3'b000;
Q_ASSERT \kdf_mode_3_.dek_op_1_.dak_op_0_.brcm_kdf_ops  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_ops_123_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_ops_123_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2231[0]));
// pragma CVASTRPROP INSTANCE "\kdf_mode_3_.dek_op_1_.dak_op_0_.brcm_kdf_ops " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\kdf_mode_3_.dek_op_1_.dak_op_0_.brcm_kdf_ops " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\kdf_mode_3_.dek_op_1_.dak_op_0_.brcm_kdf_ops " ASSERT_LINE 902
wire [2:0] n2232 = 3'b000;
Q_ASSERT \kdf_mode_3_.dek_op_1_.dak_op_1_.brcm_kdf_ops  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_ops_124_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_ops_124_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2232[0]));
// pragma CVASTRPROP INSTANCE "\kdf_mode_3_.dek_op_1_.dak_op_1_.brcm_kdf_ops " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\kdf_mode_3_.dek_op_1_.dak_op_1_.brcm_kdf_ops " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\kdf_mode_3_.dek_op_1_.dak_op_1_.brcm_kdf_ops " ASSERT_LINE 902
wire [2:0] n2233 = 3'b000;
Q_ASSERT \key_type_enc_dek_7_.null_gcm  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_null_gcm_125_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_null_gcm_125_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2233[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_7_.null_gcm " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_7_.null_gcm " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_7_.null_gcm " ASSERT_LINE 1114
wire [2:0] n2234 = 3'b000;
Q_ASSERT \key_type_enc_dek_7_.sha_gcm  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_sha_gcm_126_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_sha_gcm_126_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2234[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_7_.sha_gcm " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_7_.sha_gcm " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_7_.sha_gcm " ASSERT_LINE 1121
wire [2:0] n2235 = 3'b000;
Q_ASSERT \key_type_enc_dek_7_.null_xts  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_null_xts_127_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_null_xts_127_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2235[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_7_.null_xts " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_7_.null_xts " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_7_.null_xts " ASSERT_LINE 1127
wire [2:0] n2236 = 3'b000;
Q_ASSERT \key_type_enc_dek_7_.sha_xts  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_sha_xts_128_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_sha_xts_128_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2236[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_7_.sha_xts " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_7_.sha_xts " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_7_.sha_xts " ASSERT_LINE 1133
wire [2:0] n2237 = 3'b000;
Q_ASSERT \key_type_enc_dek_7_.null_null  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_null_null_129_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_null_null_129_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2237[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_7_.null_null " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_7_.null_null " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_7_.null_null " ASSERT_LINE 1139
wire [2:0] n2238 = 3'b000;
Q_ASSERT \key_type_enc_dek_7_.sha_null  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_sha_null_130_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_sha_null_130_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2238[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_7_.sha_null " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_7_.sha_null " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_7_.sha_null " ASSERT_LINE 1145
wire [2:0] n2239 = 3'b000;
Q_ASSERT \key_type_enc_dek_7_.hmac_gcm  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_hmac_gcm_131_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_hmac_gcm_131_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2239[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_7_.hmac_gcm " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_7_.hmac_gcm " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_7_.hmac_gcm " ASSERT_LINE 1152
wire [2:0] n2240 = 3'b000;
Q_ASSERT \key_type_enc_dek_7_.hmac_xts  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_hmac_xts_132_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_hmac_xts_132_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2240[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_7_.hmac_xts " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_7_.hmac_xts " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_7_.hmac_xts " ASSERT_LINE 1158
wire [2:0] n2241 = 3'b000;
Q_ASSERT \key_type_enc_dek_7_.hmac_null  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_hmac_null_133_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_hmac_null_133_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2241[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_7_.hmac_null " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_7_.hmac_null " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_7_.hmac_null " ASSERT_LINE 1164
wire [2:0] n2242 = 3'b000;
Q_ASSERT \key_type_enc_dek_8_.null_gcm  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_null_gcm_134_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_null_gcm_134_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2242[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_8_.null_gcm " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_8_.null_gcm " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_8_.null_gcm " ASSERT_LINE 1114
wire [2:0] n2243 = 3'b000;
Q_ASSERT \key_type_enc_dek_8_.sha_gcm  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_sha_gcm_135_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_sha_gcm_135_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2243[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_8_.sha_gcm " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_8_.sha_gcm " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_8_.sha_gcm " ASSERT_LINE 1121
wire [2:0] n2244 = 3'b000;
Q_ASSERT \key_type_enc_dek_8_.null_xts  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_null_xts_136_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_null_xts_136_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2244[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_8_.null_xts " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_8_.null_xts " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_8_.null_xts " ASSERT_LINE 1127
wire [2:0] n2245 = 3'b000;
Q_ASSERT \key_type_enc_dek_8_.sha_xts  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_sha_xts_137_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_sha_xts_137_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2245[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_8_.sha_xts " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_8_.sha_xts " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_8_.sha_xts " ASSERT_LINE 1133
wire [2:0] n2246 = 3'b000;
Q_ASSERT \key_type_enc_dek_8_.null_null  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_null_null_138_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_null_null_138_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2246[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_8_.null_null " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_8_.null_null " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_8_.null_null " ASSERT_LINE 1139
wire [2:0] n2247 = 3'b000;
Q_ASSERT \key_type_enc_dek_8_.sha_null  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_sha_null_139_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_sha_null_139_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2247[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_8_.sha_null " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_8_.sha_null " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_8_.sha_null " ASSERT_LINE 1145
wire [2:0] n2248 = 3'b000;
Q_ASSERT \key_type_enc_dek_8_.hmac_gcm  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_hmac_gcm_140_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_hmac_gcm_140_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2248[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_8_.hmac_gcm " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_8_.hmac_gcm " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_8_.hmac_gcm " ASSERT_LINE 1152
wire [2:0] n2249 = 3'b000;
Q_ASSERT \key_type_enc_dek_8_.hmac_xts  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_hmac_xts_141_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_hmac_xts_141_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2249[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_8_.hmac_xts " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_8_.hmac_xts " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_8_.hmac_xts " ASSERT_LINE 1158
wire [2:0] n2250 = 3'b000;
Q_ASSERT \key_type_enc_dek_8_.hmac_null  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_hmac_null_142_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_hmac_null_142_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2250[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_8_.hmac_null " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_8_.hmac_null " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_8_.hmac_null " ASSERT_LINE 1164
wire [2:0] n2251 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_10_.null_gcm  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_null_gcm_143_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_null_gcm_143_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2251[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_10_.null_gcm " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_10_.null_gcm " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_10_.null_gcm " ASSERT_LINE 1175
wire [2:0] n2252 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_10_.sha_gcm  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_sha_gcm_144_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_sha_gcm_144_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2252[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_10_.sha_gcm " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_10_.sha_gcm " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_10_.sha_gcm " ASSERT_LINE 1182
wire [2:0] n2253 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_10_.null_xts  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_null_xts_145_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_null_xts_145_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2253[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_10_.null_xts " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_10_.null_xts " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_10_.null_xts " ASSERT_LINE 1188
wire [2:0] n2254 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_10_.sha_xts  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_sha_xts_146_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_sha_xts_146_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2254[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_10_.sha_xts " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_10_.sha_xts " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_10_.sha_xts " ASSERT_LINE 1194
wire [2:0] n2255 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_10_.null_null  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_null_null_147_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_null_null_147_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2255[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_10_.null_null " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_10_.null_null " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_10_.null_null " ASSERT_LINE 1200
wire [2:0] n2256 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_10_.sha_null  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_sha_null_148_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_sha_null_148_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2256[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_10_.sha_null " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_10_.sha_null " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_10_.sha_null " ASSERT_LINE 1206
wire [2:0] n2257 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_10_.hmac_gcm  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_hmac_gcm_149_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_hmac_gcm_149_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2257[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_10_.hmac_gcm " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_10_.hmac_gcm " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_10_.hmac_gcm " ASSERT_LINE 1213
wire [2:0] n2258 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_10_.hmac_xts  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_hmac_xts_150_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_hmac_xts_150_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2258[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_10_.hmac_xts " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_10_.hmac_xts " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_10_.hmac_xts " ASSERT_LINE 1219
wire [2:0] n2259 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_10_.hmac_null  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_hmac_null_151_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_hmac_null_151_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2259[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_10_.hmac_null " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_10_.hmac_null " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_10_.hmac_null " ASSERT_LINE 1225
wire [2:0] n2260 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_11_.null_gcm  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_null_gcm_152_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_null_gcm_152_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2260[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_11_.null_gcm " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_11_.null_gcm " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_11_.null_gcm " ASSERT_LINE 1175
wire [2:0] n2261 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_11_.sha_gcm  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_sha_gcm_153_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_sha_gcm_153_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2261[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_11_.sha_gcm " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_11_.sha_gcm " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_11_.sha_gcm " ASSERT_LINE 1182
wire [2:0] n2262 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_11_.null_xts  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_null_xts_154_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_null_xts_154_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2262[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_11_.null_xts " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_11_.null_xts " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_11_.null_xts " ASSERT_LINE 1188
wire [2:0] n2263 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_11_.sha_xts  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_sha_xts_155_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_sha_xts_155_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2263[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_11_.sha_xts " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_11_.sha_xts " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_11_.sha_xts " ASSERT_LINE 1194
wire [2:0] n2264 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_11_.null_null  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_null_null_156_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_null_null_156_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2264[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_11_.null_null " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_11_.null_null " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_11_.null_null " ASSERT_LINE 1200
wire [2:0] n2265 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_11_.sha_null  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_sha_null_157_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_sha_null_157_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2265[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_11_.sha_null " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_11_.sha_null " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_11_.sha_null " ASSERT_LINE 1206
wire [2:0] n2266 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_11_.hmac_gcm  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_hmac_gcm_158_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_hmac_gcm_158_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2266[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_11_.hmac_gcm " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_11_.hmac_gcm " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_11_.hmac_gcm " ASSERT_LINE 1213
wire [2:0] n2267 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_11_.hmac_xts  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_hmac_xts_159_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_hmac_xts_159_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2267[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_11_.hmac_xts " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_11_.hmac_xts " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_11_.hmac_xts " ASSERT_LINE 1219
wire [2:0] n2268 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_11_.hmac_null  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_hmac_null_160_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_hmac_null_160_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2268[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_11_.hmac_null " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_11_.hmac_null " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_11_.hmac_null " ASSERT_LINE 1225
wire [2:0] n2269 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_12_.null_gcm  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_null_gcm_161_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_null_gcm_161_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2269[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_12_.null_gcm " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_12_.null_gcm " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_12_.null_gcm " ASSERT_LINE 1175
wire [2:0] n2270 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_12_.sha_gcm  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_sha_gcm_162_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_sha_gcm_162_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2270[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_12_.sha_gcm " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_12_.sha_gcm " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_12_.sha_gcm " ASSERT_LINE 1182
wire [2:0] n2271 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_12_.null_xts  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_null_xts_163_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_null_xts_163_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2271[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_12_.null_xts " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_12_.null_xts " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_12_.null_xts " ASSERT_LINE 1188
wire [2:0] n2272 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_12_.sha_xts  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_sha_xts_164_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_sha_xts_164_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2272[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_12_.sha_xts " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_12_.sha_xts " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_12_.sha_xts " ASSERT_LINE 1194
wire [2:0] n2273 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_12_.null_null  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_null_null_165_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_null_null_165_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2273[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_12_.null_null " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_12_.null_null " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_12_.null_null " ASSERT_LINE 1200
wire [2:0] n2274 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_12_.sha_null  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_sha_null_166_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_sha_null_166_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2274[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_12_.sha_null " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_12_.sha_null " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_12_.sha_null " ASSERT_LINE 1206
wire [2:0] n2275 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_12_.hmac_gcm  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_hmac_gcm_167_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_hmac_gcm_167_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2275[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_12_.hmac_gcm " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_12_.hmac_gcm " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_12_.hmac_gcm " ASSERT_LINE 1213
wire [2:0] n2276 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_12_.hmac_xts  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_hmac_xts_168_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_hmac_xts_168_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2276[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_12_.hmac_xts " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_12_.hmac_xts " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_12_.hmac_xts " ASSERT_LINE 1219
wire [2:0] n2277 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_12_.hmac_null  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_hmac_null_169_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_hmac_null_169_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2277[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_12_.hmac_null " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_12_.hmac_null " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_12_.hmac_null " ASSERT_LINE 1225
wire [2:0] n2278 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_13_.null_gcm  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_null_gcm_170_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_null_gcm_170_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2278[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_13_.null_gcm " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_13_.null_gcm " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_13_.null_gcm " ASSERT_LINE 1175
wire [2:0] n2279 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_13_.sha_gcm  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_sha_gcm_171_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_sha_gcm_171_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2279[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_13_.sha_gcm " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_13_.sha_gcm " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_13_.sha_gcm " ASSERT_LINE 1182
wire [2:0] n2280 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_13_.null_xts  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_null_xts_172_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_null_xts_172_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2280[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_13_.null_xts " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_13_.null_xts " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_13_.null_xts " ASSERT_LINE 1188
wire [2:0] n2281 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_13_.sha_xts  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_sha_xts_173_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_sha_xts_173_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2281[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_13_.sha_xts " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_13_.sha_xts " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_13_.sha_xts " ASSERT_LINE 1194
wire [2:0] n2282 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_13_.null_null  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_null_null_174_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_null_null_174_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2282[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_13_.null_null " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_13_.null_null " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_13_.null_null " ASSERT_LINE 1200
wire [2:0] n2283 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_13_.sha_null  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_sha_null_175_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_sha_null_175_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2283[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_13_.sha_null " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_13_.sha_null " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_13_.sha_null " ASSERT_LINE 1206
wire [2:0] n2284 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_13_.hmac_gcm  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_hmac_gcm_176_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_hmac_gcm_176_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2284[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_13_.hmac_gcm " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_13_.hmac_gcm " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_13_.hmac_gcm " ASSERT_LINE 1213
wire [2:0] n2285 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_13_.hmac_xts  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_hmac_xts_177_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_hmac_xts_177_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2285[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_13_.hmac_xts " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_13_.hmac_xts " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_13_.hmac_xts " ASSERT_LINE 1219
wire [2:0] n2286 = 3'b000;
Q_ASSERT \key_type_enc_dek_dak_13_.hmac_null  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_hmac_null_178_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_hmac_null_178_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2286[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_13_.hmac_null " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_dak_13_.hmac_null " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_dak_13_.hmac_null " ASSERT_LINE 1225
wire [2:0] n2287 = 3'b000;
Q_ASSERT key_type0_line4 ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_key_type0_line4_1_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_key_type0_line4_1_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2287[0]));
// pragma CVASTRPROP INSTANCE "key_type0_line4" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "key_type0_line4" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "key_type0_line4" ASSERT_LINE 914
wire [2:0] n2288 = 3'b000;
Q_ASSERT key_type0_line5a ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_key_type0_line5a_2_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_key_type0_line5a_2_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2288[0]));
// pragma CVASTRPROP INSTANCE "key_type0_line5a" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "key_type0_line5a" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "key_type0_line5a" ASSERT_LINE 920
wire [2:0] n2289 = 3'b000;
Q_ASSERT key_type0_line5b ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_key_type0_line5b_3_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_key_type0_line5b_3_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2289[0]));
// pragma CVASTRPROP INSTANCE "key_type0_line5b" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "key_type0_line5b" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "key_type0_line5b" ASSERT_LINE 926
wire [2:0] n2290 = 3'b000;
Q_ASSERT key_type1_line7a ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_key_type1_line7a_4_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_key_type1_line7a_4_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2290[0]));
// pragma CVASTRPROP INSTANCE "key_type1_line7a" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "key_type1_line7a" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "key_type1_line7a" ASSERT_LINE 936
wire [2:0] n2291 = 3'b000;
Q_ASSERT key_type1_line7b ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_key_type1_line7b_5_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_key_type1_line7b_5_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2291[0]));
// pragma CVASTRPROP INSTANCE "key_type1_line7b" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "key_type1_line7b" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "key_type1_line7b" ASSERT_LINE 944
wire [2:0] n2292 = 3'b000;
Q_ASSERT key_type1_line8a ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_key_type1_line8a_6_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_key_type1_line8a_6_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2292[0]));
// pragma CVASTRPROP INSTANCE "key_type1_line8a" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "key_type1_line8a" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "key_type1_line8a" ASSERT_LINE 952
wire [2:0] n2293 = 3'b000;
Q_ASSERT key_type1_line8b ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_key_type1_line8b_7_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_key_type1_line8b_7_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2293[0]));
// pragma CVASTRPROP INSTANCE "key_type1_line8b" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "key_type1_line8b" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "key_type1_line8b" ASSERT_LINE 960
wire [2:0] n2294 = 3'b000;
Q_ASSERT key_type1_line9 ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_key_type1_line9_8_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_key_type1_line9_8_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2294[0]));
// pragma CVASTRPROP INSTANCE "key_type1_line9" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "key_type1_line9" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "key_type1_line9" ASSERT_LINE 969
wire [2:0] n2295 = 3'b000;
Q_ASSERT key_type1_line10 ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_key_type1_line10_9_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_key_type1_line10_9_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2295[0]));
// pragma CVASTRPROP INSTANCE "key_type1_line10" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "key_type1_line10" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "key_type1_line10" ASSERT_LINE 977
wire [2:0] n2296 = 3'b000;
Q_ASSERT key_type1_line11a ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_key_type1_line11a_10_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_key_type1_line11a_10_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2296[0]));
// pragma CVASTRPROP INSTANCE "key_type1_line11a" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "key_type1_line11a" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "key_type1_line11a" ASSERT_LINE 983
wire [2:0] n2297 = 3'b000;
Q_ASSERT key_type1_line11b ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_key_type1_line11b_11_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_key_type1_line11b_11_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2297[0]));
// pragma CVASTRPROP INSTANCE "key_type1_line11b" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "key_type1_line11b" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "key_type1_line11b" ASSERT_LINE 989
wire [2:0] n2298 = 3'b000;
Q_ASSERT key_type1_line11c ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_key_type1_line11c_12_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_key_type1_line11c_12_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2298[0]));
// pragma CVASTRPROP INSTANCE "key_type1_line11c" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "key_type1_line11c" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "key_type1_line11c" ASSERT_LINE 995
wire [2:0] n2299 = 3'b000;
Q_ASSERT key_type1_line11d ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_key_type1_line11d_13_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_key_type1_line11d_13_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2299[0]));
// pragma CVASTRPROP INSTANCE "key_type1_line11d" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "key_type1_line11d" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "key_type1_line11d" ASSERT_LINE 1001
wire [2:0] n2300 = 3'b000;
Q_ASSERT key_type1_line12a ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_key_type1_line12a_14_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_key_type1_line12a_14_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2300[0]));
// pragma CVASTRPROP INSTANCE "key_type1_line12a" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "key_type1_line12a" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "key_type1_line12a" ASSERT_LINE 1007
wire [2:0] n2301 = 3'b000;
Q_ASSERT key_type1_line12b ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_key_type1_line12b_15_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_key_type1_line12b_15_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2301[0]));
// pragma CVASTRPROP INSTANCE "key_type1_line12b" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "key_type1_line12b" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "key_type1_line12b" ASSERT_LINE 1014
wire [2:0] n2302 = 3'b000;
Q_ASSERT key_type9_line14 ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_key_type9_line14_16_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_key_type9_line14_16_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2302[0]));
// pragma CVASTRPROP INSTANCE "key_type9_line14" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "key_type9_line14" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "key_type9_line14" ASSERT_LINE 1023
wire [2:0] n2303 = 3'b000;
Q_ASSERT key_type9_line15 ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_key_type9_line15_17_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_key_type9_line15_17_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2303[0]));
// pragma CVASTRPROP INSTANCE "key_type9_line15" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "key_type9_line15" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "key_type9_line15" ASSERT_LINE 1030
wire [2:0] n2304 = 3'b000;
Q_ASSERT key_type9_line16a ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_key_type9_line16a_18_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_key_type9_line16a_18_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2304[0]));
// pragma CVASTRPROP INSTANCE "key_type9_line16a" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "key_type9_line16a" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "key_type9_line16a" ASSERT_LINE 1036
wire [2:0] n2305 = 3'b000;
Q_ASSERT key_type9_line16b ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_key_type9_line16b_19_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_key_type9_line16b_19_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2305[0]));
// pragma CVASTRPROP INSTANCE "key_type9_line16b" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "key_type9_line16b" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "key_type9_line16b" ASSERT_LINE 1042
wire [2:0] n2306 = 3'b000;
Q_ASSERT key_type9_line17a ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_key_type9_line17a_20_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_key_type9_line17a_20_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2306[0]));
// pragma CVASTRPROP INSTANCE "key_type9_line17a" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "key_type9_line17a" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "key_type9_line17a" ASSERT_LINE 1050
wire [2:0] n2307 = 3'b000;
Q_ASSERT key_type9_line17b ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_key_type9_line17b_21_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_key_type9_line17b_21_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2307[0]));
// pragma CVASTRPROP INSTANCE "key_type9_line17b" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "key_type9_line17b" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "key_type9_line17b" ASSERT_LINE 1059
wire [2:0] n2308 = 3'b000;
Q_ASSERT key_type9_line18a ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_key_type9_line18a_22_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_key_type9_line18a_22_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2308[0]));
// pragma CVASTRPROP INSTANCE "key_type9_line18a" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "key_type9_line18a" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "key_type9_line18a" ASSERT_LINE 1066
wire [2:0] n2309 = 3'b000;
Q_ASSERT key_type9_line18b ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_key_type9_line18b_23_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_key_type9_line18b_23_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2309[0]));
// pragma CVASTRPROP INSTANCE "key_type9_line18b" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "key_type9_line18b" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "key_type9_line18b" ASSERT_LINE 1074
wire [2:0] n2310 = 3'b000;
Q_ASSERT key_type9_line19a ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_key_type9_line19a_24_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_key_type9_line19a_24_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2310[0]));
// pragma CVASTRPROP INSTANCE "key_type9_line19a" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "key_type9_line19a" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "key_type9_line19a" ASSERT_LINE 1081
wire [2:0] n2311 = 3'b000;
Q_ASSERT key_type9_line19b ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_key_type9_line19b_25_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_key_type9_line19b_25_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2311[0]));
// pragma CVASTRPROP INSTANCE "key_type9_line19b" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "key_type9_line19b" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "key_type9_line19b" ASSERT_LINE 1088
wire [2:0] n2312 = 3'b000;
Q_ASSERT key_type9_line19c ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_key_type9_line19c_26_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_key_type9_line19c_26_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2312[0]));
// pragma CVASTRPROP INSTANCE "key_type9_line19c" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "key_type9_line19c" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "key_type9_line19c" ASSERT_LINE 1094
wire [2:0] n2313 = 3'b000;
Q_ASSERT key_type9_line19d ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_key_type9_line19d_27_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_key_type9_line19d_27_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2313[0]));
// pragma CVASTRPROP INSTANCE "key_type9_line19d" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "key_type9_line19d" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "key_type9_line19d" ASSERT_LINE 1101
wire [2:0] n2314 = 3'b000;
Q_ASSERT guid_miss_aux_cmd_0 ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_guid_miss_aux_cmd_0_28_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_guid_miss_aux_cmd_0_28_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2314[0]));
// pragma CVASTRPROP INSTANCE "guid_miss_aux_cmd_0" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "guid_miss_aux_cmd_0" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "guid_miss_aux_cmd_0" ASSERT_LINE 1234
wire [2:0] n2315 = 3'b000;
Q_ASSERT guid_miss_aux_cmd_1 ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_guid_miss_aux_cmd_1_29_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_guid_miss_aux_cmd_1_29_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2315[0]));
// pragma CVASTRPROP INSTANCE "guid_miss_aux_cmd_1" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "guid_miss_aux_cmd_1" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "guid_miss_aux_cmd_1" ASSERT_LINE 1240
wire [2:0] n2316 = 3'b000;
Q_ASSERT guid_miss_aux_cmd_2 ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_guid_miss_aux_cmd_2_30_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_guid_miss_aux_cmd_2_30_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2316[0]));
// pragma CVASTRPROP INSTANCE "guid_miss_aux_cmd_2" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "guid_miss_aux_cmd_2" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "guid_miss_aux_cmd_2" ASSERT_LINE 1246
wire [2:0] n2317 = 3'b000;
Q_ASSERT guid_miss_aux_cmd_3 ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_guid_miss_aux_cmd_3_31_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_guid_miss_aux_cmd_3_31_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2317[0]));
// pragma CVASTRPROP INSTANCE "guid_miss_aux_cmd_3" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "guid_miss_aux_cmd_3" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "guid_miss_aux_cmd_3" ASSERT_LINE 1252
wire [2:0] n2318 = 3'b000;
Q_ASSERT guid_miss_aux_cmd_iv_0 ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_guid_miss_aux_cmd_iv_0_32_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_guid_miss_aux_cmd_iv_0_32_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2318[0]));
// pragma CVASTRPROP INSTANCE "guid_miss_aux_cmd_iv_0" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "guid_miss_aux_cmd_iv_0" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "guid_miss_aux_cmd_iv_0" ASSERT_LINE 1258
wire [2:0] n2319 = 3'b000;
Q_ASSERT guid_miss_aux_cmd_iv_1 ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_guid_miss_aux_cmd_iv_1_33_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_guid_miss_aux_cmd_iv_1_33_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2319[0]));
// pragma CVASTRPROP INSTANCE "guid_miss_aux_cmd_iv_1" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "guid_miss_aux_cmd_iv_1" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "guid_miss_aux_cmd_iv_1" ASSERT_LINE 1264
wire [2:0] n2320 = 3'b000;
Q_ASSERT guid_miss_aux_cmd_iv_2 ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_guid_miss_aux_cmd_iv_2_34_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_guid_miss_aux_cmd_iv_2_34_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2320[0]));
// pragma CVASTRPROP INSTANCE "guid_miss_aux_cmd_iv_2" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "guid_miss_aux_cmd_iv_2" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "guid_miss_aux_cmd_iv_2" ASSERT_LINE 1270
wire [2:0] n2321 = 3'b000;
Q_ASSERT guid_miss_aux_cmd_iv_3 ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_guid_miss_aux_cmd_iv_3_35_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_guid_miss_aux_cmd_iv_3_35_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2321[0]));
// pragma CVASTRPROP INSTANCE "guid_miss_aux_cmd_iv_3" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "guid_miss_aux_cmd_iv_3" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "guid_miss_aux_cmd_iv_3" ASSERT_LINE 1276
wire [2:0] n2322 = 3'b000;
Q_ASSERT iv_miss_aux_cmd_0 ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_iv_miss_aux_cmd_0_36_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_iv_miss_aux_cmd_0_36_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2322[0]));
// pragma CVASTRPROP INSTANCE "iv_miss_aux_cmd_0" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "iv_miss_aux_cmd_0" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "iv_miss_aux_cmd_0" ASSERT_LINE 1282
wire [2:0] n2323 = 3'b000;
Q_ASSERT iv_miss_aux_cmd_1 ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_iv_miss_aux_cmd_1_37_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_iv_miss_aux_cmd_1_37_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2323[0]));
// pragma CVASTRPROP INSTANCE "iv_miss_aux_cmd_1" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "iv_miss_aux_cmd_1" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "iv_miss_aux_cmd_1" ASSERT_LINE 1287
wire [2:0] n2324 = 3'b000;
Q_ASSERT iv_miss_aux_cmd_guid ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_iv_miss_aux_cmd_guid_38_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_iv_miss_aux_cmd_guid_38_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2324[0]));
// pragma CVASTRPROP INSTANCE "iv_miss_aux_cmd_guid" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "iv_miss_aux_cmd_guid" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v"
//pragma CVAINTPROP INSTANCE "iv_miss_aux_cmd_guid" ASSERT_LINE 1292
Q_XOR2 U6247 ( .A0(int_tlv_counter[1]), .A1(int_tlv_counter[0]), .Z(n134));
Q_FDP4EP \_zy_sva_key_type0_line4_1_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_key_type0_line4_1_ccheck[0]));
Q_FDP4EP \_zy_sva_key_type0_line4_1_cpass_REG[0] ( .CK(clk), .CE(n1926), .R(n1735), .D(n47), .Q(_zy_sva_key_type0_line4_1_cpass[0]));
Q_FDP4EP \_zy_sva_key_type0_line5a_2_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_key_type0_line5a_2_ccheck[0]));
Q_FDP4EP \_zy_sva_key_type0_line5a_2_cpass_REG[0] ( .CK(clk), .CE(n1925), .R(n1735), .D(n47), .Q(_zy_sva_key_type0_line5a_2_cpass[0]));
Q_FDP4EP \_zy_sva_key_type0_line5b_3_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_key_type0_line5b_3_ccheck[0]));
Q_FDP4EP \_zy_sva_key_type0_line5b_3_cpass_REG[0] ( .CK(clk), .CE(n1924), .R(n1735), .D(n47), .Q(_zy_sva_key_type0_line5b_3_cpass[0]));
Q_FDP4EP \_zy_sva_key_type1_line7a_4_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_key_type1_line7a_4_ccheck[0]));
Q_FDP4EP \_zy_sva_key_type1_line7a_4_cpass_REG[0] ( .CK(clk), .CE(n1923), .R(n1735), .D(n47), .Q(_zy_sva_key_type1_line7a_4_cpass[0]));
Q_FDP4EP \_zy_sva_key_type1_line7b_5_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_key_type1_line7b_5_ccheck[0]));
Q_FDP4EP \_zy_sva_key_type1_line7b_5_cpass_REG[0] ( .CK(clk), .CE(n1922), .R(n1735), .D(n47), .Q(_zy_sva_key_type1_line7b_5_cpass[0]));
Q_FDP4EP \_zy_sva_key_type1_line8a_6_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_key_type1_line8a_6_ccheck[0]));
Q_FDP4EP \_zy_sva_key_type1_line8a_6_cpass_REG[0] ( .CK(clk), .CE(n1921), .R(n1735), .D(n47), .Q(_zy_sva_key_type1_line8a_6_cpass[0]));
Q_FDP4EP \_zy_sva_key_type1_line8b_7_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_key_type1_line8b_7_ccheck[0]));
Q_FDP4EP \_zy_sva_key_type1_line8b_7_cpass_REG[0] ( .CK(clk), .CE(n1920), .R(n1735), .D(n47), .Q(_zy_sva_key_type1_line8b_7_cpass[0]));
Q_FDP4EP \_zy_sva_key_type1_line9_8_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_key_type1_line9_8_ccheck[0]));
Q_FDP4EP \_zy_sva_key_type1_line9_8_cpass_REG[0] ( .CK(clk), .CE(n1919), .R(n1735), .D(n47), .Q(_zy_sva_key_type1_line9_8_cpass[0]));
Q_FDP4EP \_zy_sva_key_type1_line10_9_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_key_type1_line10_9_ccheck[0]));
Q_FDP4EP \_zy_sva_key_type1_line10_9_cpass_REG[0] ( .CK(clk), .CE(n1918), .R(n1735), .D(n47), .Q(_zy_sva_key_type1_line10_9_cpass[0]));
Q_FDP4EP \_zy_sva_key_type1_line11a_10_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_key_type1_line11a_10_ccheck[0]));
Q_FDP4EP \_zy_sva_key_type1_line11a_10_cpass_REG[0] ( .CK(clk), .CE(n1917), .R(n1735), .D(n47), .Q(_zy_sva_key_type1_line11a_10_cpass[0]));
Q_FDP4EP \_zy_sva_key_type1_line11b_11_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_key_type1_line11b_11_ccheck[0]));
Q_FDP4EP \_zy_sva_key_type1_line11b_11_cpass_REG[0] ( .CK(clk), .CE(n1916), .R(n1735), .D(n47), .Q(_zy_sva_key_type1_line11b_11_cpass[0]));
Q_FDP4EP \_zy_sva_key_type1_line11c_12_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_key_type1_line11c_12_ccheck[0]));
Q_FDP4EP \_zy_sva_key_type1_line11c_12_cpass_REG[0] ( .CK(clk), .CE(n1915), .R(n1735), .D(n47), .Q(_zy_sva_key_type1_line11c_12_cpass[0]));
Q_FDP4EP \_zy_sva_key_type1_line11d_13_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_key_type1_line11d_13_ccheck[0]));
Q_FDP4EP \_zy_sva_key_type1_line11d_13_cpass_REG[0] ( .CK(clk), .CE(n1914), .R(n1735), .D(n47), .Q(_zy_sva_key_type1_line11d_13_cpass[0]));
Q_FDP4EP \_zy_sva_key_type1_line12a_14_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_key_type1_line12a_14_ccheck[0]));
Q_FDP4EP \_zy_sva_key_type1_line12a_14_cpass_REG[0] ( .CK(clk), .CE(n1913), .R(n1735), .D(n47), .Q(_zy_sva_key_type1_line12a_14_cpass[0]));
Q_FDP4EP \_zy_sva_key_type1_line12b_15_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_key_type1_line12b_15_ccheck[0]));
Q_FDP4EP \_zy_sva_key_type1_line12b_15_cpass_REG[0] ( .CK(clk), .CE(n1912), .R(n1735), .D(n47), .Q(_zy_sva_key_type1_line12b_15_cpass[0]));
Q_FDP4EP \_zy_sva_key_type9_line14_16_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_key_type9_line14_16_ccheck[0]));
Q_FDP4EP \_zy_sva_key_type9_line14_16_cpass_REG[0] ( .CK(clk), .CE(n1911), .R(n1735), .D(n47), .Q(_zy_sva_key_type9_line14_16_cpass[0]));
Q_FDP4EP \_zy_sva_key_type9_line15_17_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_key_type9_line15_17_ccheck[0]));
Q_FDP4EP \_zy_sva_key_type9_line15_17_cpass_REG[0] ( .CK(clk), .CE(n1910), .R(n1735), .D(n47), .Q(_zy_sva_key_type9_line15_17_cpass[0]));
Q_FDP4EP \_zy_sva_key_type9_line16a_18_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_key_type9_line16a_18_ccheck[0]));
Q_FDP4EP \_zy_sva_key_type9_line16a_18_cpass_REG[0] ( .CK(clk), .CE(n1909), .R(n1735), .D(n47), .Q(_zy_sva_key_type9_line16a_18_cpass[0]));
Q_FDP4EP \_zy_sva_key_type9_line16b_19_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_key_type9_line16b_19_ccheck[0]));
Q_FDP4EP \_zy_sva_key_type9_line16b_19_cpass_REG[0] ( .CK(clk), .CE(n1908), .R(n1735), .D(n47), .Q(_zy_sva_key_type9_line16b_19_cpass[0]));
Q_FDP4EP \_zy_sva_key_type9_line17a_20_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_key_type9_line17a_20_ccheck[0]));
Q_FDP4EP \_zy_sva_key_type9_line17a_20_cpass_REG[0] ( .CK(clk), .CE(n1907), .R(n1735), .D(n47), .Q(_zy_sva_key_type9_line17a_20_cpass[0]));
Q_FDP4EP \_zy_sva_key_type9_line17b_21_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_key_type9_line17b_21_ccheck[0]));
Q_FDP4EP \_zy_sva_key_type9_line17b_21_cpass_REG[0] ( .CK(clk), .CE(n1906), .R(n1735), .D(n47), .Q(_zy_sva_key_type9_line17b_21_cpass[0]));
Q_FDP4EP \_zy_sva_key_type9_line18a_22_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_key_type9_line18a_22_ccheck[0]));
Q_FDP4EP \_zy_sva_key_type9_line18a_22_cpass_REG[0] ( .CK(clk), .CE(n1905), .R(n1735), .D(n47), .Q(_zy_sva_key_type9_line18a_22_cpass[0]));
Q_FDP4EP \_zy_sva_key_type9_line18b_23_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_key_type9_line18b_23_ccheck[0]));
Q_FDP4EP \_zy_sva_key_type9_line18b_23_cpass_REG[0] ( .CK(clk), .CE(n1904), .R(n1735), .D(n47), .Q(_zy_sva_key_type9_line18b_23_cpass[0]));
Q_FDP4EP \_zy_sva_key_type9_line19a_24_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_key_type9_line19a_24_ccheck[0]));
Q_FDP4EP \_zy_sva_key_type9_line19a_24_cpass_REG[0] ( .CK(clk), .CE(n1903), .R(n1735), .D(n47), .Q(_zy_sva_key_type9_line19a_24_cpass[0]));
Q_FDP4EP \_zy_sva_key_type9_line19b_25_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_key_type9_line19b_25_ccheck[0]));
Q_FDP4EP \_zy_sva_key_type9_line19b_25_cpass_REG[0] ( .CK(clk), .CE(n1902), .R(n1735), .D(n47), .Q(_zy_sva_key_type9_line19b_25_cpass[0]));
Q_FDP4EP \_zy_sva_key_type9_line19c_26_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_key_type9_line19c_26_ccheck[0]));
Q_FDP4EP \_zy_sva_key_type9_line19c_26_cpass_REG[0] ( .CK(clk), .CE(n1901), .R(n1735), .D(n47), .Q(_zy_sva_key_type9_line19c_26_cpass[0]));
Q_FDP4EP \_zy_sva_key_type9_line19d_27_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_key_type9_line19d_27_ccheck[0]));
Q_FDP4EP \_zy_sva_key_type9_line19d_27_cpass_REG[0] ( .CK(clk), .CE(n1900), .R(n1735), .D(n47), .Q(_zy_sva_key_type9_line19d_27_cpass[0]));
Q_FDP4EP \_zy_sva_guid_miss_aux_cmd_0_28_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_guid_miss_aux_cmd_0_28_ccheck[0]));
Q_FDP4EP \_zy_sva_guid_miss_aux_cmd_0_28_cpass_REG[0] ( .CK(clk), .CE(n1899), .R(n1735), .D(n47), .Q(_zy_sva_guid_miss_aux_cmd_0_28_cpass[0]));
Q_FDP4EP \_zy_sva_guid_miss_aux_cmd_1_29_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_guid_miss_aux_cmd_1_29_ccheck[0]));
Q_FDP4EP \_zy_sva_guid_miss_aux_cmd_1_29_cpass_REG[0] ( .CK(clk), .CE(n1898), .R(n1735), .D(n47), .Q(_zy_sva_guid_miss_aux_cmd_1_29_cpass[0]));
Q_FDP4EP \_zy_sva_guid_miss_aux_cmd_2_30_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_guid_miss_aux_cmd_2_30_ccheck[0]));
Q_FDP4EP \_zy_sva_guid_miss_aux_cmd_2_30_cpass_REG[0] ( .CK(clk), .CE(n1897), .R(n1735), .D(n47), .Q(_zy_sva_guid_miss_aux_cmd_2_30_cpass[0]));
Q_FDP4EP \_zy_sva_guid_miss_aux_cmd_3_31_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_guid_miss_aux_cmd_3_31_ccheck[0]));
Q_FDP4EP \_zy_sva_guid_miss_aux_cmd_3_31_cpass_REG[0] ( .CK(clk), .CE(n1896), .R(n1735), .D(n47), .Q(_zy_sva_guid_miss_aux_cmd_3_31_cpass[0]));
Q_FDP4EP \_zy_sva_guid_miss_aux_cmd_iv_0_32_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_guid_miss_aux_cmd_iv_0_32_ccheck[0]));
Q_FDP4EP \_zy_sva_guid_miss_aux_cmd_iv_0_32_cpass_REG[0] ( .CK(clk), .CE(n1895), .R(n1735), .D(n47), .Q(_zy_sva_guid_miss_aux_cmd_iv_0_32_cpass[0]));
Q_FDP4EP \_zy_sva_guid_miss_aux_cmd_iv_1_33_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_guid_miss_aux_cmd_iv_1_33_ccheck[0]));
Q_FDP4EP \_zy_sva_guid_miss_aux_cmd_iv_1_33_cpass_REG[0] ( .CK(clk), .CE(n1894), .R(n1735), .D(n47), .Q(_zy_sva_guid_miss_aux_cmd_iv_1_33_cpass[0]));
Q_FDP4EP \_zy_sva_guid_miss_aux_cmd_iv_2_34_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_guid_miss_aux_cmd_iv_2_34_ccheck[0]));
Q_FDP4EP \_zy_sva_guid_miss_aux_cmd_iv_2_34_cpass_REG[0] ( .CK(clk), .CE(n1893), .R(n1735), .D(n47), .Q(_zy_sva_guid_miss_aux_cmd_iv_2_34_cpass[0]));
Q_FDP4EP \_zy_sva_guid_miss_aux_cmd_iv_3_35_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_guid_miss_aux_cmd_iv_3_35_ccheck[0]));
Q_FDP4EP \_zy_sva_guid_miss_aux_cmd_iv_3_35_cpass_REG[0] ( .CK(clk), .CE(n1892), .R(n1735), .D(n47), .Q(_zy_sva_guid_miss_aux_cmd_iv_3_35_cpass[0]));
Q_FDP4EP \_zy_sva_iv_miss_aux_cmd_0_36_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_iv_miss_aux_cmd_0_36_ccheck[0]));
Q_FDP4EP \_zy_sva_iv_miss_aux_cmd_0_36_cpass_REG[0] ( .CK(clk), .CE(n1891), .R(n1735), .D(n47), .Q(_zy_sva_iv_miss_aux_cmd_0_36_cpass[0]));
Q_FDP4EP \_zy_sva_iv_miss_aux_cmd_1_37_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_iv_miss_aux_cmd_1_37_ccheck[0]));
Q_FDP4EP \_zy_sva_iv_miss_aux_cmd_1_37_cpass_REG[0] ( .CK(clk), .CE(n1890), .R(n1735), .D(n47), .Q(_zy_sva_iv_miss_aux_cmd_1_37_cpass[0]));
Q_FDP4EP \_zy_sva_iv_miss_aux_cmd_guid_38_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_iv_miss_aux_cmd_guid_38_ccheck[0]));
Q_FDP4EP \_zy_sva_iv_miss_aux_cmd_guid_38_cpass_REG[0] ( .CK(clk), .CE(n1889), .R(n1735), .D(n47), .Q(_zy_sva_iv_miss_aux_cmd_guid_38_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_39_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_39_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_39_cpass_REG[0] ( .CK(clk), .CE(n1888), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_39_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_iv_40_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_iv_40_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_iv_40_cpass_REG[0] ( .CK(clk), .CE(n1887), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_iv_40_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_41_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_41_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_41_cpass_REG[0] ( .CK(clk), .CE(n1886), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_41_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_iv_42_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_iv_42_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_iv_42_cpass_REG[0] ( .CK(clk), .CE(n1885), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_iv_42_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_key_type_43_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_key_type_43_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_key_type_43_cpass_REG[0] ( .CK(clk), .CE(n1884), .R(n1735), .D(n47), .Q(_zy_sva_brcm_key_type_43_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_44_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_44_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_44_cpass_REG[0] ( .CK(clk), .CE(n1883), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_44_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_iv_45_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_iv_45_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_iv_45_cpass_REG[0] ( .CK(clk), .CE(n1882), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_iv_45_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_46_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_46_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_46_cpass_REG[0] ( .CK(clk), .CE(n1881), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_46_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_iv_47_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_iv_47_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_iv_47_cpass_REG[0] ( .CK(clk), .CE(n1880), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_iv_47_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_key_type_48_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_key_type_48_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_key_type_48_cpass_REG[0] ( .CK(clk), .CE(n1879), .R(n1735), .D(n47), .Q(_zy_sva_brcm_key_type_48_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_49_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_49_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_49_cpass_REG[0] ( .CK(clk), .CE(n1878), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_49_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_iv_50_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_iv_50_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_iv_50_cpass_REG[0] ( .CK(clk), .CE(n1877), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_iv_50_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_51_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_51_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_51_cpass_REG[0] ( .CK(clk), .CE(n1876), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_51_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_iv_52_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_iv_52_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_iv_52_cpass_REG[0] ( .CK(clk), .CE(n1875), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_iv_52_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_key_type_53_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_key_type_53_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_key_type_53_cpass_REG[0] ( .CK(clk), .CE(n1874), .R(n1735), .D(n47), .Q(_zy_sva_brcm_key_type_53_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_54_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_54_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_54_cpass_REG[0] ( .CK(clk), .CE(n1873), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_54_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_iv_55_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_iv_55_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_iv_55_cpass_REG[0] ( .CK(clk), .CE(n1872), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_iv_55_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_56_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_56_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_56_cpass_REG[0] ( .CK(clk), .CE(n1871), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_56_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_iv_57_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_iv_57_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_iv_57_cpass_REG[0] ( .CK(clk), .CE(n1870), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_iv_57_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_key_type_58_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_key_type_58_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_key_type_58_cpass_REG[0] ( .CK(clk), .CE(n1869), .R(n1735), .D(n47), .Q(_zy_sva_brcm_key_type_58_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_59_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_59_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_59_cpass_REG[0] ( .CK(clk), .CE(n1868), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_59_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_iv_60_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_iv_60_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_iv_60_cpass_REG[0] ( .CK(clk), .CE(n1867), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_iv_60_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_61_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_61_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_61_cpass_REG[0] ( .CK(clk), .CE(n1866), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_61_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_iv_62_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_iv_62_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_iv_62_cpass_REG[0] ( .CK(clk), .CE(n1865), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_iv_62_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_key_type_63_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_key_type_63_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_key_type_63_cpass_REG[0] ( .CK(clk), .CE(n1864), .R(n1735), .D(n47), .Q(_zy_sva_brcm_key_type_63_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_64_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_64_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_64_cpass_REG[0] ( .CK(clk), .CE(n1863), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_64_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_iv_65_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_iv_65_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_iv_65_cpass_REG[0] ( .CK(clk), .CE(n1862), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_iv_65_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_66_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_66_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_66_cpass_REG[0] ( .CK(clk), .CE(n1861), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_66_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_iv_67_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_iv_67_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_iv_67_cpass_REG[0] ( .CK(clk), .CE(n1860), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_iv_67_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_key_type_68_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_key_type_68_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_key_type_68_cpass_REG[0] ( .CK(clk), .CE(n1859), .R(n1735), .D(n47), .Q(_zy_sva_brcm_key_type_68_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_69_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_69_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_69_cpass_REG[0] ( .CK(clk), .CE(n1858), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_69_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_iv_70_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_iv_70_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_iv_70_cpass_REG[0] ( .CK(clk), .CE(n1857), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_iv_70_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_71_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_71_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_71_cpass_REG[0] ( .CK(clk), .CE(n1856), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_71_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_iv_72_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_iv_72_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_iv_72_cpass_REG[0] ( .CK(clk), .CE(n1855), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_iv_72_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_key_type_73_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_key_type_73_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_key_type_73_cpass_REG[0] ( .CK(clk), .CE(n1854), .R(n1735), .D(n47), .Q(_zy_sva_brcm_key_type_73_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_74_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_74_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_74_cpass_REG[0] ( .CK(clk), .CE(n1853), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_74_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_iv_75_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_iv_75_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_iv_75_cpass_REG[0] ( .CK(clk), .CE(n1852), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_iv_75_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_76_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_76_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_76_cpass_REG[0] ( .CK(clk), .CE(n1851), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_76_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_iv_77_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_iv_77_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_iv_77_cpass_REG[0] ( .CK(clk), .CE(n1850), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_iv_77_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_key_type_78_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_key_type_78_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_key_type_78_cpass_REG[0] ( .CK(clk), .CE(n1849), .R(n1735), .D(n47), .Q(_zy_sva_brcm_key_type_78_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_79_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_79_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_79_cpass_REG[0] ( .CK(clk), .CE(n1848), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_79_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_iv_80_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_iv_80_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_iv_80_cpass_REG[0] ( .CK(clk), .CE(n1847), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_iv_80_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_81_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_81_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_81_cpass_REG[0] ( .CK(clk), .CE(n1846), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_81_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_iv_82_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_iv_82_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_iv_82_cpass_REG[0] ( .CK(clk), .CE(n1845), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_iv_82_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_key_type_83_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_key_type_83_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_key_type_83_cpass_REG[0] ( .CK(clk), .CE(n1844), .R(n1735), .D(n47), .Q(_zy_sva_brcm_key_type_83_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_84_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_84_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_84_cpass_REG[0] ( .CK(clk), .CE(n1843), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_84_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_iv_85_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_iv_85_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_iv_85_cpass_REG[0] ( .CK(clk), .CE(n1842), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_iv_85_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_86_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_86_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_86_cpass_REG[0] ( .CK(clk), .CE(n1841), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_86_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_iv_87_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_iv_87_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_iv_87_cpass_REG[0] ( .CK(clk), .CE(n1840), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_iv_87_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_key_type_88_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_key_type_88_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_key_type_88_cpass_REG[0] ( .CK(clk), .CE(n1839), .R(n1735), .D(n47), .Q(_zy_sva_brcm_key_type_88_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_89_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_89_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_89_cpass_REG[0] ( .CK(clk), .CE(n1838), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_89_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_iv_90_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_iv_90_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_iv_90_cpass_REG[0] ( .CK(clk), .CE(n1837), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_iv_90_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_91_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_91_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_91_cpass_REG[0] ( .CK(clk), .CE(n1836), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_91_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_iv_92_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_iv_92_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_iv_92_cpass_REG[0] ( .CK(clk), .CE(n1835), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_iv_92_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_key_type_93_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_key_type_93_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_key_type_93_cpass_REG[0] ( .CK(clk), .CE(n1834), .R(n1735), .D(n47), .Q(_zy_sva_brcm_key_type_93_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_94_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_94_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_94_cpass_REG[0] ( .CK(clk), .CE(n1833), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_94_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_iv_95_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_iv_95_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_iv_95_cpass_REG[0] ( .CK(clk), .CE(n1832), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_iv_95_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_96_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_96_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_96_cpass_REG[0] ( .CK(clk), .CE(n1831), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_96_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_iv_97_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_iv_97_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_iv_97_cpass_REG[0] ( .CK(clk), .CE(n1830), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_iv_97_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_key_type_98_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_key_type_98_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_key_type_98_cpass_REG[0] ( .CK(clk), .CE(n1829), .R(n1735), .D(n47), .Q(_zy_sva_brcm_key_type_98_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_99_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_99_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_99_cpass_REG[0] ( .CK(clk), .CE(n1828), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_99_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_iv_100_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_iv_100_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_iv_100_cpass_REG[0] ( .CK(clk), .CE(n1827), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_iv_100_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_101_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_101_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_101_cpass_REG[0] ( .CK(clk), .CE(n1826), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_101_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_iv_102_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_iv_102_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_iv_102_cpass_REG[0] ( .CK(clk), .CE(n1825), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_iv_102_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_key_type_103_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_key_type_103_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_key_type_103_cpass_REG[0] ( .CK(clk), .CE(n1824), .R(n1735), .D(n47), .Q(_zy_sva_brcm_key_type_103_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_104_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_104_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_104_cpass_REG[0] ( .CK(clk), .CE(n1823), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_104_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_iv_105_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_iv_105_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_iv_105_cpass_REG[0] ( .CK(clk), .CE(n1822), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_iv_105_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_106_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_106_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_106_cpass_REG[0] ( .CK(clk), .CE(n1821), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_106_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_iv_107_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_iv_107_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_aux_cmd_guid_iv_107_cpass_REG[0] ( .CK(clk), .CE(n1820), .R(n1735), .D(n47), .Q(_zy_sva_brcm_aux_cmd_guid_iv_107_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_key_type_108_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_key_type_108_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_key_type_108_cpass_REG[0] ( .CK(clk), .CE(n1819), .R(n1735), .D(n47), .Q(_zy_sva_brcm_key_type_108_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_109_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_109_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_109_cpass_REG[0] ( .CK(clk), .CE(n1818), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_109_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_110_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_110_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_110_cpass_REG[0] ( .CK(clk), .CE(n1817), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_110_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_111_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_111_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_111_cpass_REG[0] ( .CK(clk), .CE(n1816), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_111_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_112_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_112_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_112_cpass_REG[0] ( .CK(clk), .CE(n1815), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_112_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_113_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_113_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_113_cpass_REG[0] ( .CK(clk), .CE(n1814), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_113_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_114_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_114_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_114_cpass_REG[0] ( .CK(clk), .CE(n1813), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_114_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_115_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_115_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_115_cpass_REG[0] ( .CK(clk), .CE(n1812), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_115_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_116_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_116_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_116_cpass_REG[0] ( .CK(clk), .CE(n1811), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_116_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_117_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_117_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_117_cpass_REG[0] ( .CK(clk), .CE(n1810), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_117_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_118_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_118_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_118_cpass_REG[0] ( .CK(clk), .CE(n1809), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_118_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_119_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_119_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_119_cpass_REG[0] ( .CK(clk), .CE(n1808), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_119_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_120_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_120_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_120_cpass_REG[0] ( .CK(clk), .CE(n1807), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_120_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_121_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_121_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_121_cpass_REG[0] ( .CK(clk), .CE(n1806), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_121_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_122_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_122_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_122_cpass_REG[0] ( .CK(clk), .CE(n1805), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_122_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_123_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_123_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_123_cpass_REG[0] ( .CK(clk), .CE(n1804), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_123_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_124_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_124_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_ops_124_cpass_REG[0] ( .CK(clk), .CE(n1803), .R(n1735), .D(n47), .Q(_zy_sva_brcm_kdf_ops_124_cpass[0]));
Q_FDP4EP \_zy_sva_null_gcm_125_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_null_gcm_125_ccheck[0]));
Q_FDP4EP \_zy_sva_null_gcm_125_cpass_REG[0] ( .CK(clk), .CE(n1802), .R(n1735), .D(n47), .Q(_zy_sva_null_gcm_125_cpass[0]));
Q_FDP4EP \_zy_sva_sha_gcm_126_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_sha_gcm_126_ccheck[0]));
Q_FDP4EP \_zy_sva_sha_gcm_126_cpass_REG[0] ( .CK(clk), .CE(n1801), .R(n1735), .D(n47), .Q(_zy_sva_sha_gcm_126_cpass[0]));
Q_FDP4EP \_zy_sva_null_xts_127_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_null_xts_127_ccheck[0]));
Q_FDP4EP \_zy_sva_null_xts_127_cpass_REG[0] ( .CK(clk), .CE(n1800), .R(n1735), .D(n47), .Q(_zy_sva_null_xts_127_cpass[0]));
Q_FDP4EP \_zy_sva_sha_xts_128_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_sha_xts_128_ccheck[0]));
Q_FDP4EP \_zy_sva_sha_xts_128_cpass_REG[0] ( .CK(clk), .CE(n1799), .R(n1735), .D(n47), .Q(_zy_sva_sha_xts_128_cpass[0]));
Q_FDP4EP \_zy_sva_null_null_129_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_null_null_129_ccheck[0]));
Q_FDP4EP \_zy_sva_null_null_129_cpass_REG[0] ( .CK(clk), .CE(n1798), .R(n1735), .D(n47), .Q(_zy_sva_null_null_129_cpass[0]));
Q_FDP4EP \_zy_sva_sha_null_130_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_sha_null_130_ccheck[0]));
Q_FDP4EP \_zy_sva_sha_null_130_cpass_REG[0] ( .CK(clk), .CE(n1797), .R(n1735), .D(n47), .Q(_zy_sva_sha_null_130_cpass[0]));
Q_FDP4EP \_zy_sva_hmac_gcm_131_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_hmac_gcm_131_ccheck[0]));
Q_FDP4EP \_zy_sva_hmac_gcm_131_cpass_REG[0] ( .CK(clk), .CE(n1796), .R(n1735), .D(n47), .Q(_zy_sva_hmac_gcm_131_cpass[0]));
Q_FDP4EP \_zy_sva_hmac_xts_132_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_hmac_xts_132_ccheck[0]));
Q_FDP4EP \_zy_sva_hmac_xts_132_cpass_REG[0] ( .CK(clk), .CE(n1795), .R(n1735), .D(n47), .Q(_zy_sva_hmac_xts_132_cpass[0]));
Q_FDP4EP \_zy_sva_hmac_null_133_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_hmac_null_133_ccheck[0]));
Q_FDP4EP \_zy_sva_hmac_null_133_cpass_REG[0] ( .CK(clk), .CE(n1794), .R(n1735), .D(n47), .Q(_zy_sva_hmac_null_133_cpass[0]));
Q_FDP4EP \_zy_sva_null_gcm_134_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_null_gcm_134_ccheck[0]));
Q_FDP4EP \_zy_sva_null_gcm_134_cpass_REG[0] ( .CK(clk), .CE(n1793), .R(n1735), .D(n47), .Q(_zy_sva_null_gcm_134_cpass[0]));
Q_FDP4EP \_zy_sva_sha_gcm_135_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_sha_gcm_135_ccheck[0]));
Q_FDP4EP \_zy_sva_sha_gcm_135_cpass_REG[0] ( .CK(clk), .CE(n1792), .R(n1735), .D(n47), .Q(_zy_sva_sha_gcm_135_cpass[0]));
Q_FDP4EP \_zy_sva_null_xts_136_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_null_xts_136_ccheck[0]));
Q_FDP4EP \_zy_sva_null_xts_136_cpass_REG[0] ( .CK(clk), .CE(n1791), .R(n1735), .D(n47), .Q(_zy_sva_null_xts_136_cpass[0]));
Q_FDP4EP \_zy_sva_sha_xts_137_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_sha_xts_137_ccheck[0]));
Q_FDP4EP \_zy_sva_sha_xts_137_cpass_REG[0] ( .CK(clk), .CE(n1790), .R(n1735), .D(n47), .Q(_zy_sva_sha_xts_137_cpass[0]));
Q_FDP4EP \_zy_sva_null_null_138_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_null_null_138_ccheck[0]));
Q_FDP4EP \_zy_sva_null_null_138_cpass_REG[0] ( .CK(clk), .CE(n1789), .R(n1735), .D(n47), .Q(_zy_sva_null_null_138_cpass[0]));
Q_FDP4EP \_zy_sva_sha_null_139_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_sha_null_139_ccheck[0]));
Q_FDP4EP \_zy_sva_sha_null_139_cpass_REG[0] ( .CK(clk), .CE(n1788), .R(n1735), .D(n47), .Q(_zy_sva_sha_null_139_cpass[0]));
Q_FDP4EP \_zy_sva_hmac_gcm_140_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_hmac_gcm_140_ccheck[0]));
Q_FDP4EP \_zy_sva_hmac_gcm_140_cpass_REG[0] ( .CK(clk), .CE(n1787), .R(n1735), .D(n47), .Q(_zy_sva_hmac_gcm_140_cpass[0]));
Q_FDP4EP \_zy_sva_hmac_xts_141_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_hmac_xts_141_ccheck[0]));
Q_FDP4EP \_zy_sva_hmac_xts_141_cpass_REG[0] ( .CK(clk), .CE(n1786), .R(n1735), .D(n47), .Q(_zy_sva_hmac_xts_141_cpass[0]));
Q_FDP4EP \_zy_sva_hmac_null_142_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_hmac_null_142_ccheck[0]));
Q_FDP4EP \_zy_sva_hmac_null_142_cpass_REG[0] ( .CK(clk), .CE(n1785), .R(n1735), .D(n47), .Q(_zy_sva_hmac_null_142_cpass[0]));
Q_FDP4EP \_zy_sva_null_gcm_143_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_null_gcm_143_ccheck[0]));
Q_FDP4EP \_zy_sva_null_gcm_143_cpass_REG[0] ( .CK(clk), .CE(n1784), .R(n1735), .D(n47), .Q(_zy_sva_null_gcm_143_cpass[0]));
Q_FDP4EP \_zy_sva_sha_gcm_144_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_sha_gcm_144_ccheck[0]));
Q_FDP4EP \_zy_sva_sha_gcm_144_cpass_REG[0] ( .CK(clk), .CE(n1783), .R(n1735), .D(n47), .Q(_zy_sva_sha_gcm_144_cpass[0]));
Q_FDP4EP \_zy_sva_null_xts_145_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_null_xts_145_ccheck[0]));
Q_FDP4EP \_zy_sva_null_xts_145_cpass_REG[0] ( .CK(clk), .CE(n1782), .R(n1735), .D(n47), .Q(_zy_sva_null_xts_145_cpass[0]));
Q_FDP4EP \_zy_sva_sha_xts_146_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_sha_xts_146_ccheck[0]));
Q_FDP4EP \_zy_sva_sha_xts_146_cpass_REG[0] ( .CK(clk), .CE(n1781), .R(n1735), .D(n47), .Q(_zy_sva_sha_xts_146_cpass[0]));
Q_FDP4EP \_zy_sva_null_null_147_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_null_null_147_ccheck[0]));
Q_FDP4EP \_zy_sva_null_null_147_cpass_REG[0] ( .CK(clk), .CE(n1780), .R(n1735), .D(n47), .Q(_zy_sva_null_null_147_cpass[0]));
Q_FDP4EP \_zy_sva_sha_null_148_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_sha_null_148_ccheck[0]));
Q_FDP4EP \_zy_sva_sha_null_148_cpass_REG[0] ( .CK(clk), .CE(n1779), .R(n1735), .D(n47), .Q(_zy_sva_sha_null_148_cpass[0]));
Q_FDP4EP \_zy_sva_hmac_gcm_149_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_hmac_gcm_149_ccheck[0]));
Q_FDP4EP \_zy_sva_hmac_gcm_149_cpass_REG[0] ( .CK(clk), .CE(n1778), .R(n1735), .D(n47), .Q(_zy_sva_hmac_gcm_149_cpass[0]));
Q_FDP4EP \_zy_sva_hmac_xts_150_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_hmac_xts_150_ccheck[0]));
Q_FDP4EP \_zy_sva_hmac_xts_150_cpass_REG[0] ( .CK(clk), .CE(n1777), .R(n1735), .D(n47), .Q(_zy_sva_hmac_xts_150_cpass[0]));
Q_FDP4EP \_zy_sva_hmac_null_151_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_hmac_null_151_ccheck[0]));
Q_FDP4EP \_zy_sva_hmac_null_151_cpass_REG[0] ( .CK(clk), .CE(n1776), .R(n1735), .D(n47), .Q(_zy_sva_hmac_null_151_cpass[0]));
Q_FDP4EP \_zy_sva_null_gcm_152_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_null_gcm_152_ccheck[0]));
Q_FDP4EP \_zy_sva_null_gcm_152_cpass_REG[0] ( .CK(clk), .CE(n1775), .R(n1735), .D(n47), .Q(_zy_sva_null_gcm_152_cpass[0]));
Q_FDP4EP \_zy_sva_sha_gcm_153_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_sha_gcm_153_ccheck[0]));
Q_FDP4EP \_zy_sva_sha_gcm_153_cpass_REG[0] ( .CK(clk), .CE(n1774), .R(n1735), .D(n47), .Q(_zy_sva_sha_gcm_153_cpass[0]));
Q_FDP4EP \_zy_sva_null_xts_154_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_null_xts_154_ccheck[0]));
Q_FDP4EP \_zy_sva_null_xts_154_cpass_REG[0] ( .CK(clk), .CE(n1773), .R(n1735), .D(n47), .Q(_zy_sva_null_xts_154_cpass[0]));
Q_FDP4EP \_zy_sva_sha_xts_155_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_sha_xts_155_ccheck[0]));
Q_FDP4EP \_zy_sva_sha_xts_155_cpass_REG[0] ( .CK(clk), .CE(n1772), .R(n1735), .D(n47), .Q(_zy_sva_sha_xts_155_cpass[0]));
Q_FDP4EP \_zy_sva_null_null_156_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_null_null_156_ccheck[0]));
Q_FDP4EP \_zy_sva_null_null_156_cpass_REG[0] ( .CK(clk), .CE(n1771), .R(n1735), .D(n47), .Q(_zy_sva_null_null_156_cpass[0]));
Q_FDP4EP \_zy_sva_sha_null_157_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_sha_null_157_ccheck[0]));
Q_FDP4EP \_zy_sva_sha_null_157_cpass_REG[0] ( .CK(clk), .CE(n1770), .R(n1735), .D(n47), .Q(_zy_sva_sha_null_157_cpass[0]));
Q_FDP4EP \_zy_sva_hmac_gcm_158_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_hmac_gcm_158_ccheck[0]));
Q_FDP4EP \_zy_sva_hmac_gcm_158_cpass_REG[0] ( .CK(clk), .CE(n1769), .R(n1735), .D(n47), .Q(_zy_sva_hmac_gcm_158_cpass[0]));
Q_FDP4EP \_zy_sva_hmac_xts_159_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_hmac_xts_159_ccheck[0]));
Q_FDP4EP \_zy_sva_hmac_xts_159_cpass_REG[0] ( .CK(clk), .CE(n1768), .R(n1735), .D(n47), .Q(_zy_sva_hmac_xts_159_cpass[0]));
Q_FDP4EP \_zy_sva_hmac_null_160_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_hmac_null_160_ccheck[0]));
Q_FDP4EP \_zy_sva_hmac_null_160_cpass_REG[0] ( .CK(clk), .CE(n1767), .R(n1735), .D(n47), .Q(_zy_sva_hmac_null_160_cpass[0]));
Q_FDP4EP \_zy_sva_null_gcm_161_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_null_gcm_161_ccheck[0]));
Q_FDP4EP \_zy_sva_null_gcm_161_cpass_REG[0] ( .CK(clk), .CE(n1766), .R(n1735), .D(n47), .Q(_zy_sva_null_gcm_161_cpass[0]));
Q_FDP4EP \_zy_sva_sha_gcm_162_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_sha_gcm_162_ccheck[0]));
Q_FDP4EP \_zy_sva_sha_gcm_162_cpass_REG[0] ( .CK(clk), .CE(n1765), .R(n1735), .D(n47), .Q(_zy_sva_sha_gcm_162_cpass[0]));
Q_FDP4EP \_zy_sva_null_xts_163_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_null_xts_163_ccheck[0]));
Q_FDP4EP \_zy_sva_null_xts_163_cpass_REG[0] ( .CK(clk), .CE(n1764), .R(n1735), .D(n47), .Q(_zy_sva_null_xts_163_cpass[0]));
Q_FDP4EP \_zy_sva_sha_xts_164_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_sha_xts_164_ccheck[0]));
Q_FDP4EP \_zy_sva_sha_xts_164_cpass_REG[0] ( .CK(clk), .CE(n1763), .R(n1735), .D(n47), .Q(_zy_sva_sha_xts_164_cpass[0]));
Q_FDP4EP \_zy_sva_null_null_165_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_null_null_165_ccheck[0]));
Q_FDP4EP \_zy_sva_null_null_165_cpass_REG[0] ( .CK(clk), .CE(n1762), .R(n1735), .D(n47), .Q(_zy_sva_null_null_165_cpass[0]));
Q_FDP4EP \_zy_sva_sha_null_166_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_sha_null_166_ccheck[0]));
Q_FDP4EP \_zy_sva_sha_null_166_cpass_REG[0] ( .CK(clk), .CE(n1761), .R(n1735), .D(n47), .Q(_zy_sva_sha_null_166_cpass[0]));
Q_FDP4EP \_zy_sva_hmac_gcm_167_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_hmac_gcm_167_ccheck[0]));
Q_FDP4EP \_zy_sva_hmac_gcm_167_cpass_REG[0] ( .CK(clk), .CE(n1760), .R(n1735), .D(n47), .Q(_zy_sva_hmac_gcm_167_cpass[0]));
Q_FDP4EP \_zy_sva_hmac_xts_168_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_hmac_xts_168_ccheck[0]));
Q_FDP4EP \_zy_sva_hmac_xts_168_cpass_REG[0] ( .CK(clk), .CE(n1759), .R(n1735), .D(n47), .Q(_zy_sva_hmac_xts_168_cpass[0]));
Q_FDP4EP \_zy_sva_hmac_null_169_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_hmac_null_169_ccheck[0]));
Q_FDP4EP \_zy_sva_hmac_null_169_cpass_REG[0] ( .CK(clk), .CE(n1758), .R(n1735), .D(n47), .Q(_zy_sva_hmac_null_169_cpass[0]));
Q_FDP4EP \_zy_sva_null_gcm_170_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_null_gcm_170_ccheck[0]));
Q_FDP4EP \_zy_sva_null_gcm_170_cpass_REG[0] ( .CK(clk), .CE(n1757), .R(n1735), .D(n47), .Q(_zy_sva_null_gcm_170_cpass[0]));
Q_FDP4EP \_zy_sva_sha_gcm_171_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_sha_gcm_171_ccheck[0]));
Q_FDP4EP \_zy_sva_sha_gcm_171_cpass_REG[0] ( .CK(clk), .CE(n1756), .R(n1735), .D(n47), .Q(_zy_sva_sha_gcm_171_cpass[0]));
Q_FDP4EP \_zy_sva_null_xts_172_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_null_xts_172_ccheck[0]));
Q_FDP4EP \_zy_sva_null_xts_172_cpass_REG[0] ( .CK(clk), .CE(n1755), .R(n1735), .D(n47), .Q(_zy_sva_null_xts_172_cpass[0]));
Q_FDP4EP \_zy_sva_sha_xts_173_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_sha_xts_173_ccheck[0]));
Q_FDP4EP \_zy_sva_sha_xts_173_cpass_REG[0] ( .CK(clk), .CE(n1754), .R(n1735), .D(n47), .Q(_zy_sva_sha_xts_173_cpass[0]));
Q_FDP4EP \_zy_sva_null_null_174_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_null_null_174_ccheck[0]));
Q_FDP4EP \_zy_sva_null_null_174_cpass_REG[0] ( .CK(clk), .CE(n1753), .R(n1735), .D(n47), .Q(_zy_sva_null_null_174_cpass[0]));
Q_FDP4EP \_zy_sva_sha_null_175_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_sha_null_175_ccheck[0]));
Q_FDP4EP \_zy_sva_sha_null_175_cpass_REG[0] ( .CK(clk), .CE(n1752), .R(n1735), .D(n47), .Q(_zy_sva_sha_null_175_cpass[0]));
Q_FDP4EP \_zy_sva_hmac_gcm_176_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_hmac_gcm_176_ccheck[0]));
Q_FDP4EP \_zy_sva_hmac_gcm_176_cpass_REG[0] ( .CK(clk), .CE(n1751), .R(n1735), .D(n47), .Q(_zy_sva_hmac_gcm_176_cpass[0]));
Q_FDP4EP \_zy_sva_hmac_xts_177_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_hmac_xts_177_ccheck[0]));
Q_FDP4EP \_zy_sva_hmac_xts_177_cpass_REG[0] ( .CK(clk), .CE(n1750), .R(n1735), .D(n47), .Q(_zy_sva_hmac_xts_177_cpass[0]));
Q_FDP4EP \_zy_sva_hmac_null_178_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n1735), .D(n47), .Q(_zy_sva_hmac_null_178_ccheck[0]));
Q_FDP4EP \_zy_sva_hmac_null_178_cpass_REG[0] ( .CK(clk), .CE(n1749), .R(n1735), .D(n47), .Q(_zy_sva_hmac_null_178_cpass[0]));
Q_FDP4EP \tlv_counter_REG[4] ( .CK(clk), .CE(stitcher_rd), .R(n2146), .D(n1736), .Q(tlv_counter[4]));
Q_INV U6605 ( .A(rst_n), .Z(n2146));
Q_FDP4EP \tlv_counter_REG[3] ( .CK(clk), .CE(stitcher_rd), .R(n2146), .D(n1737), .Q(tlv_counter[3]));
Q_INV U6607 ( .A(tlv_counter[3]), .Z(n538));
Q_FDP4EP \tlv_counter_REG[2] ( .CK(clk), .CE(stitcher_rd), .R(n2146), .D(n1738), .Q(tlv_counter[2]));
Q_INV U6609 ( .A(tlv_counter[2]), .Z(n444));
Q_FDP4EP \tlv_counter_REG[1] ( .CK(clk), .CE(stitcher_rd), .R(n2146), .D(n1739), .Q(tlv_counter[1]));
Q_INV U6611 ( .A(tlv_counter[1]), .Z(n534));
Q_FDP4EP \tlv_counter_REG[0] ( .CK(clk), .CE(stitcher_rd), .R(n2146), .D(n1740), .Q(tlv_counter[0]));
Q_INV U6613 ( .A(tlv_counter[0]), .Z(n1748));
Q_FDP4EP \int_tlv_counter_REG[5] ( .CK(clk), .CE(fifo_in_valid), .R(n2146), .D(n121), .Q(int_tlv_counter[5]));
Q_INV U6615 ( .A(int_tlv_counter[5]), .Z(n706));
Q_FDP4EP \int_tlv_counter_REG[4] ( .CK(clk), .CE(fifo_in_valid), .R(n2146), .D(n122), .Q(int_tlv_counter[4]));
Q_INV U6617 ( .A(int_tlv_counter[4]), .Z(n688));
Q_FDP4EP \int_tlv_counter_REG[3] ( .CK(clk), .CE(fifo_in_valid), .R(n2146), .D(n123), .Q(int_tlv_counter[3]));
Q_INV U6619 ( .A(int_tlv_counter[3]), .Z(n697));
Q_FDP4EP \int_tlv_counter_REG[2] ( .CK(clk), .CE(fifo_in_valid), .R(n2146), .D(n124), .Q(int_tlv_counter[2]));
Q_INV U6621 ( .A(int_tlv_counter[2]), .Z(n2135));
Q_FDP4EP \int_tlv_counter_REG[1] ( .CK(clk), .CE(fifo_in_valid), .R(n2146), .D(n125), .Q(int_tlv_counter[1]));
Q_INV U6623 ( .A(int_tlv_counter[1]), .Z(n2136));
Q_FDP4EP \int_tlv_counter_REG[0] ( .CK(clk), .CE(fifo_in_valid), .R(n2146), .D(n126), .Q(int_tlv_counter[0]));
Q_INV U6625 ( .A(int_tlv_counter[0]), .Z(n682));
Q_FDP4EP \fifo_in_REG[68] ( .CK(clk), .CE(n110), .R(n2146), .D(n45), .Q(fifo_in[68]));
Q_FDP4EP key_blob_region_REG  ( .CK(clk), .CE(n109), .R(n2146), .D(n111), .Q(key_blob_region));
Q_INV U6628 ( .A(key_blob_region), .Z(n617));
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "\parser_kimreader_data.sot  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m2 "\parser_kimreader_data.eoi  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m3 "\parser_kimreader_data.eot  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m4 "\parser_kimreader_data.id  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m5 "\parser_kimreader_data.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m6 "\stitcher_out.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m7 "\stitcher_out.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m8 "\stitcher_out.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m9 "\stitcher_out.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m10 "\fifo_in.sot  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m11 "\fifo_in.eoi  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m12 "\fifo_in.eot  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m13 "\fifo_in.id  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m14 "\fifo_in.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m15 "\tlv_word0.tlv_bip2  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m16 "\tlv_word0.frame_size  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m17 "\tlv_word0.trace  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m18 "\tlv_word0.unused  (1,0) 1 10 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m19 "\tlv_word0.tlv_frame_num  (1,0) 1 10 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m20 "\tlv_word0.resv0  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m21 "\tlv_word0.tlv_eng_id  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m22 "\tlv_word0.tlv_seq_num  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m23 "\tlv_word0.tlv_len  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m24 "\tlv_word0.tlv_type  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m25 "\tlv_word1.pf_number  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m26 "\tlv_word1.vf_number  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m27 "\tlv_word1.scheduler_handle  (1,0) 1 15 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m28 "\tlv_word1.src_data_len  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m29 "\tlv_word2.key_type  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m30 "\tlv_word2.rsvd1  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m31 "\tlv_word2.cipher_pad  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m32 "\tlv_word2.iv_op  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m33 "\tlv_word2.aad_len  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m34 "\tlv_word2.cipher_op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m35 "\tlv_word2.auth_op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m36 "\tlv_word2.raw_auth_op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m37 "\tlv_word2.rsvd0  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m38 "\tlv_word2.chu_comp_thrsh  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m39 "\tlv_word2.xp10_crc_mode  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m40 "\tlv_word2.xp10_user_prefix_size  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m41 "\tlv_word2.xp10_prefix_mode  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m42 "\tlv_word2.lz77_max_symb_len  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m43 "\tlv_word2.lz77_min_match_len  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m44 "\tlv_word2.lz77_dly_match_win  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m45 "\tlv_word2.lz77_win_size  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m46 "\tlv_word2.comp_mode  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m47 "\frame_word.debug.tlvp_corrupt  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m48 "\frame_word.debug.cmd_mode  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m49 "\frame_word.debug.module_id  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m50 "\frame_word.debug.cmd_type  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m51 "\frame_word.debug.tlv_num  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m52 "\frame_word.debug.byte_num  (1,0) 1 9 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m53 "\frame_word.debug.byte_msk  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m54 "\frame_word.frmd_out_type  (1,0) 1 6 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m55 "\frame_word.md_op  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m56 "\frame_word.md_type  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m57 "\frame_word.frmd_in_type  (1,0) 1 6 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m58 "\frame_word.frmd_in_aux  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m59 "\frame_word.frmd_crc_in  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m60 "\frame_word.src_guid_present  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m61 "\frame_word.compound_cmd_frm_size  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m62 "\kme_internal_word0.tlv_bip2  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m63 "\kme_internal_word0.resv0  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m64 "\kme_internal_word0.kdf_dek_iter  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m65 "\kme_internal_word0.keyless_algos  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m66 "\kme_internal_word0.needs_dek  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m67 "\kme_internal_word0.needs_dak  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m68 "\kme_internal_word0.key_type  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m69 "\kme_internal_word0.tlv_frame_num  (1,0) 1 10 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m70 "\kme_internal_word0.tlv_eng_id  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m71 "\kme_internal_word0.tlv_seq_num  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m72 "\kme_internal_word0.tlv_len  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m73 "\kme_internal_word0.tlv_type  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m74 "\nxt_kme_internal_word0.tlv_bip2  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m75 "\nxt_kme_internal_word0.resv0  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m76 "\nxt_kme_internal_word0.kdf_dek_iter  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m77 "\nxt_kme_internal_word0.keyless_algos  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m78 "\nxt_kme_internal_word0.needs_dek  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m79 "\nxt_kme_internal_word0.needs_dak  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m80 "\nxt_kme_internal_word0.key_type  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m81 "\nxt_kme_internal_word0.tlv_frame_num  (1,0) 1 10 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m82 "\nxt_kme_internal_word0.tlv_eng_id  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m83 "\nxt_kme_internal_word0.tlv_seq_num  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m84 "\nxt_kme_internal_word0.tlv_len  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m85 "\nxt_kme_internal_word0.tlv_type  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m86 "\kme_internal_dek_kim_word.dek_kim_entry.valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m87 "\kme_internal_dek_kim_word.dek_kim_entry.label_index  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m88 "\kme_internal_dek_kim_word.dek_kim_entry.ckv_length  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m89 "\kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer  (1,0) 1 14 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m90 "\kme_internal_dek_kim_word.dek_kim_entry.pf_num  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m91 "\kme_internal_dek_kim_word.dek_kim_entry.vf_num  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m92 "\kme_internal_dek_kim_word.dek_kim_entry.vf_valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m93 "\kme_internal_dek_kim_word.unused  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m94 "\kme_internal_dek_kim_word.missing_iv  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m95 "\kme_internal_dek_kim_word.missing_guid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m96 "\kme_internal_dek_kim_word.validate_dek  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m97 "\kme_internal_dek_kim_word.vf_valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m98 "\kme_internal_dek_kim_word.pf_num  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m99 "\kme_internal_dek_kim_word.vf_num  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m100 "\nxt_kme_internal_dek_kim_word.dek_kim_entry.valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m101 "\nxt_kme_internal_dek_kim_word.dek_kim_entry.label_index  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m102 "\nxt_kme_internal_dek_kim_word.dek_kim_entry.ckv_length  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m103 "\nxt_kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer  (1,0) 1 14 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m104 "\nxt_kme_internal_dek_kim_word.dek_kim_entry.pf_num  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m105 "\nxt_kme_internal_dek_kim_word.dek_kim_entry.vf_num  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m106 "\nxt_kme_internal_dek_kim_word.dek_kim_entry.vf_valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m107 "\nxt_kme_internal_dek_kim_word.unused  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m108 "\nxt_kme_internal_dek_kim_word.missing_iv  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m109 "\nxt_kme_internal_dek_kim_word.missing_guid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m110 "\nxt_kme_internal_dek_kim_word.validate_dek  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m111 "\nxt_kme_internal_dek_kim_word.vf_valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m112 "\nxt_kme_internal_dek_kim_word.pf_num  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m113 "\nxt_kme_internal_dek_kim_word.vf_num  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m114 "\kme_internal_dak_kim_word.dak_kim_entry.valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m115 "\kme_internal_dak_kim_word.dak_kim_entry.label_index  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m116 "\kme_internal_dak_kim_word.dak_kim_entry.ckv_length  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m117 "\kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer  (1,0) 1 14 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m118 "\kme_internal_dak_kim_word.dak_kim_entry.pf_num  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m119 "\kme_internal_dak_kim_word.dak_kim_entry.vf_num  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m120 "\kme_internal_dak_kim_word.dak_kim_entry.vf_valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m121 "\kme_internal_dak_kim_word.unused  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m122 "\kme_internal_dak_kim_word.validate_dak  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m123 "\kme_internal_dak_kim_word.vf_valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m124 "\kme_internal_dak_kim_word.pf_num  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m125 "\kme_internal_dak_kim_word.vf_num  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m126 "\nxt_kme_internal_dak_kim_word.dak_kim_entry.valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m127 "\nxt_kme_internal_dak_kim_word.dak_kim_entry.label_index  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m128 "\nxt_kme_internal_dak_kim_word.dak_kim_entry.ckv_length  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m129 "\nxt_kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer  (1,0) 1 14 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m130 "\nxt_kme_internal_dak_kim_word.dak_kim_entry.pf_num  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m131 "\nxt_kme_internal_dak_kim_word.dak_kim_entry.vf_num  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m132 "\nxt_kme_internal_dak_kim_word.dak_kim_entry.vf_valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m133 "\nxt_kme_internal_dak_kim_word.unused  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m134 "\nxt_kme_internal_dak_kim_word.validate_dak  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m135 "\nxt_kme_internal_dak_kim_word.vf_valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m136 "\nxt_kme_internal_dak_kim_word.pf_num  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m137 "\nxt_kme_internal_dak_kim_word.vf_num  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m138 "\debug_cmd.tlvp_corrupt  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m139 "\debug_cmd.cmd_mode  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m140 "\debug_cmd.module_id  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m141 "\debug_cmd.cmd_type  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m142 "\debug_cmd.tlv_num  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m143 "\debug_cmd.byte_num  (1,0) 1 9 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m144 "\debug_cmd.byte_msk  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m145 "\nxt_debug_cmd.tlvp_corrupt  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m146 "\nxt_debug_cmd.cmd_mode  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m147 "\nxt_debug_cmd.module_id  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m148 "\nxt_debug_cmd.cmd_type  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m149 "\nxt_debug_cmd.tlv_num  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m150 "\nxt_debug_cmd.byte_num  (1,0) 1 9 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m151 "\nxt_debug_cmd.byte_msk  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m152 "\aux_key_header.dak_key_op  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m153 "\aux_key_header.dak_key_ref  (1,0) 1 13 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m154 "\aux_key_header.kdf_mode  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m155 "\aux_key_header.dek_key_op  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m156 "\aux_key_header.dek_key_ref  (1,0) 1 13 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m157 "\nxt_aux_key_header.dak_key_op  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m158 "\nxt_aux_key_header.dak_key_ref  (1,0) 1 13 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m159 "\nxt_aux_key_header.kdf_mode  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m160 "\nxt_aux_key_header.dek_key_op  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m161 "\nxt_aux_key_header.dek_key_ref  (1,0) 1 13 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m162 "\skip.start  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m163 "\skip.partial  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m164 "\skip.endian_swap  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m165 "\skip.till  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m166 "\nxt_skip.start  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m167 "\nxt_skip.partial  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m168 "\nxt_skip.endian_swap  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m169 "\nxt_skip.till  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "169"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r1 "parser_kimreader_data 5 \parser_kimreader_data.sot  \parser_kimreader_data.eoi  \parser_kimreader_data.eot  \parser_kimreader_data.id  \parser_kimreader_data.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r2 "stitcher_out 6 \stitcher_out.tvalid  \stitcher_out.tlast  \stitcher_out.tid  \stitcher_out.tstrb  \stitcher_out.tuser  \stitcher_out.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r3 "fifo_in 5 \fifo_in.sot  \fifo_in.eoi  \fifo_in.eot  \fifo_in.id  \fifo_in.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r4 "tlv_word0 13 \tlv_word0.tlv_bip2  \tlv_word0.no_data  \tlv_word0.aux_frmd_crc  \tlv_word0.frame_size  \tlv_word0.vf_valid  \tlv_word0.trace  \tlv_word0.unused  \tlv_word0.tlv_frame_num  \tlv_word0.resv0  \tlv_word0.tlv_eng_id  \tlv_word0.tlv_seq_num  \tlv_word0.tlv_len  \tlv_word0.tlv_type "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r5 "tlv_word1 4 \tlv_word1.pf_number  \tlv_word1.vf_number  \tlv_word1.scheduler_handle  \tlv_word1.src_data_len "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r6 "tlv_word2 19 \tlv_word2.rsvd2  \tlv_word2.key_type  \tlv_word2.rsvd1  \tlv_word2.cipher_pad  \tlv_word2.iv_op  \tlv_word2.aad_len  \tlv_word2.cipher_op  \tlv_word2.auth_op  \tlv_word2.raw_auth_op  \tlv_word2.rsvd0  \tlv_word2.chu_comp_thrsh  \tlv_word2.xp10_crc_mode  \tlv_word2.xp10_user_prefix_size  \tlv_word2.xp10_prefix_mode  \tlv_word2.lz77_max_symb_len  \tlv_word2.lz77_min_match_len  \tlv_word2.lz77_dly_match_win  \tlv_word2.lz77_win_size  \tlv_word2.comp_mode "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r7 "frame_word 11 \frame_word.debug  { \frame_word.debug.tlvp_corrupt  \frame_word.debug.cmd_mode  \frame_word.debug.module_id  \frame_word.debug.cmd_type  \frame_word.debug.tlv_num  \frame_word.debug.byte_num  \frame_word.debug.byte_msk  } \frame_word.trace  \frame_word.dst_guid_present  \frame_word.frmd_out_type  \frame_word.md_op  \frame_word.md_type  \frame_word.frmd_in_type  \frame_word.frmd_in_aux  \frame_word.frmd_crc_in  \frame_word.src_guid_present  \frame_word.compound_cmd_frm_size "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r8 "kme_internal_word0 12 \kme_internal_word0.tlv_bip2  \kme_internal_word0.resv0  \kme_internal_word0.kdf_dek_iter  \kme_internal_word0.keyless_algos  \kme_internal_word0.needs_dek  \kme_internal_word0.needs_dak  \kme_internal_word0.key_type  \kme_internal_word0.tlv_frame_num  \kme_internal_word0.tlv_eng_id  \kme_internal_word0.tlv_seq_num  \kme_internal_word0.tlv_len  \kme_internal_word0.tlv_type "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r9 "nxt_kme_internal_word0 12 \nxt_kme_internal_word0.tlv_bip2  \nxt_kme_internal_word0.resv0  \nxt_kme_internal_word0.kdf_dek_iter  \nxt_kme_internal_word0.keyless_algos  \nxt_kme_internal_word0.needs_dek  \nxt_kme_internal_word0.needs_dak  \nxt_kme_internal_word0.key_type  \nxt_kme_internal_word0.tlv_frame_num  \nxt_kme_internal_word0.tlv_eng_id  \nxt_kme_internal_word0.tlv_seq_num  \nxt_kme_internal_word0.tlv_len  \nxt_kme_internal_word0.tlv_type "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r10 "kme_internal_dek_kim_word 8 \kme_internal_dek_kim_word.dek_kim_entry  { \kme_internal_dek_kim_word.dek_kim_entry.valid  \kme_internal_dek_kim_word.dek_kim_entry.label_index  \kme_internal_dek_kim_word.dek_kim_entry.ckv_length  \kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer  \kme_internal_dek_kim_word.dek_kim_entry.pf_num  \kme_internal_dek_kim_word.dek_kim_entry.vf_num  \kme_internal_dek_kim_word.dek_kim_entry.vf_valid  } \kme_internal_dek_kim_word.unused  \kme_internal_dek_kim_word.missing_iv  \kme_internal_dek_kim_word.missing_guid  \kme_internal_dek_kim_word.validate_dek  \kme_internal_dek_kim_word.vf_valid  \kme_internal_dek_kim_word.pf_num  \kme_internal_dek_kim_word.vf_num "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r11 "nxt_kme_internal_dek_kim_word 8 \nxt_kme_internal_dek_kim_word.dek_kim_entry  { \nxt_kme_internal_dek_kim_word.dek_kim_entry.valid  \nxt_kme_internal_dek_kim_word.dek_kim_entry.label_index  \nxt_kme_internal_dek_kim_word.dek_kim_entry.ckv_length  \nxt_kme_internal_dek_kim_word.dek_kim_entry.ckv_pointer  \nxt_kme_internal_dek_kim_word.dek_kim_entry.pf_num  \nxt_kme_internal_dek_kim_word.dek_kim_entry.vf_num  \nxt_kme_internal_dek_kim_word.dek_kim_entry.vf_valid  } \nxt_kme_internal_dek_kim_word.unused  \nxt_kme_internal_dek_kim_word.missing_iv  \nxt_kme_internal_dek_kim_word.missing_guid  \nxt_kme_internal_dek_kim_word.validate_dek  \nxt_kme_internal_dek_kim_word.vf_valid  \nxt_kme_internal_dek_kim_word.pf_num  \nxt_kme_internal_dek_kim_word.vf_num "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r12 "kme_internal_dak_kim_word 6 \kme_internal_dak_kim_word.dak_kim_entry  { \kme_internal_dak_kim_word.dak_kim_entry.valid  \kme_internal_dak_kim_word.dak_kim_entry.label_index  \kme_internal_dak_kim_word.dak_kim_entry.ckv_length  \kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer  \kme_internal_dak_kim_word.dak_kim_entry.pf_num  \kme_internal_dak_kim_word.dak_kim_entry.vf_num  \kme_internal_dak_kim_word.dak_kim_entry.vf_valid  } \kme_internal_dak_kim_word.unused  \kme_internal_dak_kim_word.validate_dak  \kme_internal_dak_kim_word.vf_valid  \kme_internal_dak_kim_word.pf_num  \kme_internal_dak_kim_word.vf_num "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r13 "nxt_kme_internal_dak_kim_word 6 \nxt_kme_internal_dak_kim_word.dak_kim_entry  { \nxt_kme_internal_dak_kim_word.dak_kim_entry.valid  \nxt_kme_internal_dak_kim_word.dak_kim_entry.label_index  \nxt_kme_internal_dak_kim_word.dak_kim_entry.ckv_length  \nxt_kme_internal_dak_kim_word.dak_kim_entry.ckv_pointer  \nxt_kme_internal_dak_kim_word.dak_kim_entry.pf_num  \nxt_kme_internal_dak_kim_word.dak_kim_entry.vf_num  \nxt_kme_internal_dak_kim_word.dak_kim_entry.vf_valid  } \nxt_kme_internal_dak_kim_word.unused  \nxt_kme_internal_dak_kim_word.validate_dak  \nxt_kme_internal_dak_kim_word.vf_valid  \nxt_kme_internal_dak_kim_word.pf_num  \nxt_kme_internal_dak_kim_word.vf_num "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r14 "debug_cmd 7 \debug_cmd.tlvp_corrupt  \debug_cmd.cmd_mode  \debug_cmd.module_id  \debug_cmd.cmd_type  \debug_cmd.tlv_num  \debug_cmd.byte_num  \debug_cmd.byte_msk "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r15 "nxt_debug_cmd 7 \nxt_debug_cmd.tlvp_corrupt  \nxt_debug_cmd.cmd_mode  \nxt_debug_cmd.module_id  \nxt_debug_cmd.cmd_type  \nxt_debug_cmd.tlv_num  \nxt_debug_cmd.byte_num  \nxt_debug_cmd.byte_msk "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r16 "aux_key_header 5 \aux_key_header.dak_key_op  \aux_key_header.dak_key_ref  \aux_key_header.kdf_mode  \aux_key_header.dek_key_op  \aux_key_header.dek_key_ref "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r17 "nxt_aux_key_header 5 \nxt_aux_key_header.dak_key_op  \nxt_aux_key_header.dak_key_ref  \nxt_aux_key_header.kdf_mode  \nxt_aux_key_header.dek_key_op  \nxt_aux_key_header.dek_key_ref "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r18 "skip 4 \skip.start  \skip.partial  \skip.endian_swap  \skip.till "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r19 "nxt_skip 4 \nxt_skip.start  \nxt_skip.partial  \nxt_skip.endian_swap  \nxt_skip.till "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_NUM "19"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_5 "-1 key_type_enc_dek_dak 10 13 "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_4 "-1 key_type_enc_dek 7 8 "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_3 "2 dak_op 0 1 "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_2 "1 dek_op 0 1 "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_1 "-1 kdf_mode 0 3 "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_0 "-1 key_type 0 13 "
// pragma CVASTRPROP MODULE HDLICE PROP_RANOFF TRUE
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type_enc_dek_dak[13]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type_enc_dek_dak[12]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type_enc_dek_dak[11]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type_enc_dek_dak[10]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type_enc_dek[8]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type_enc_dek[7]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[3].dek_op[1].dak_op[1]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[3].dek_op[1].dak_op[0]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[3].dek_op[1]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[3].dek_op[0].dak_op[1]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[3].dek_op[0].dak_op[0]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[3].dek_op[0]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[3]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[2].dek_op[1].dak_op[1]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[2].dek_op[1].dak_op[0]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[2].dek_op[1]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[2].dek_op[0].dak_op[1]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[2].dek_op[0].dak_op[0]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[2].dek_op[0]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[2]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[1].dek_op[1].dak_op[1]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[1].dek_op[1].dak_op[0]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[1].dek_op[1]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[1].dek_op[0].dak_op[1]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[1].dek_op[0].dak_op[0]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[1].dek_op[0]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[1]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[0].dek_op[1].dak_op[1]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[0].dek_op[1].dak_op[0]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[0].dek_op[1]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[0].dek_op[0].dak_op[1]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[0].dek_op[0].dak_op[0]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[0].dek_op[0]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[0]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type[13]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type[12]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type[11]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type[10]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type[9]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type[8]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type[7]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type[6]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type[5]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type[4]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type[3]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type[2]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type[1]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type[0]"
endmodule
