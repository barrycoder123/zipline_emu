
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
(* celldefine = 1 *) 
module nx_indirect_access_cntrl_xcm112 ( clk, rst_n, wr_stb, reg_addr, cmnd_op, 
	cmnd_addr, cmnd_table_id, stat_code, stat_datawords, stat_addr, 
	stat_table_id, capability_lst, capability_type, enable, .addr_limit( {
	\addr_limit[0][4] , \addr_limit[0][3] , \addr_limit[0][2] , 
	\addr_limit[0][1] , \addr_limit[0][0] } ), wr_dat, rd_dat, sw_cs, 
	sw_ce, sw_we, sw_add, sw_wdat, sw_rdat, sw_match, sw_aindex, grant, 
	yield, reset);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
input clk;
input rst_n;
input wr_stb;
input [10:0] reg_addr;
input [3:0] cmnd_op;
input [4:0] cmnd_addr;
input [0:0] cmnd_table_id;
output [2:0] stat_code;
output [4:0] stat_datawords;
output [4:0] stat_addr;
output [0:0] stat_table_id;
output [15:0] capability_lst;
output [3:0] capability_type;
output enable;
input \addr_limit[0][4] ;
input \addr_limit[0][3] ;
input \addr_limit[0][2] ;
input \addr_limit[0][1] ;
input \addr_limit[0][0] ;
input [63:0] wr_dat;
output [63:0] rd_dat;
output sw_cs;
output sw_ce;
output sw_we;
output [4:0] sw_add;
output [63:0] sw_wdat;
input [63:0] sw_rdat;
input sw_match;
input [3:0] sw_aindex;
input grant;
output yield;
output reset;
wire [0:2] _zy_simnet_stat_code_0_w$;
wire [0:4] _zy_simnet_stat_datawords_1_w$;
wire [0:4] _zy_simnet_stat_addr_2_w$;
wire _zy_simnet_stat_table_id_3_w$;
wire [0:15] _zy_simnet_capability_lst_4_w$;
wire [0:3] _zy_simnet_capability_type_5_w$;
wire _zy_simnet_enable_6_w$;
wire [0:63] _zy_simnet_rd_dat_7_w$;
wire _zy_simnet_sw_cs_8_w$;
wire _zy_simnet_sw_ce_9_w$;
wire _zy_simnet_sw_we_10_w$;
wire [0:4] _zy_simnet_sw_add_11_w$;
wire [0:63] _zy_simnet_sw_wdat_12_w$;
wire _zy_simnet_yield_13_w$;
wire _zy_simnet_reset_14_w$;
wire [3:0] cmnd;
wire init_r;
wire [0:0] inc_r;
wire init_inc_r;
wire sw_cs_r;
wire sw_ce_r;
wire rst_r;
wire rst_or_ini_r;
wire [4:0] rst_addr_r;
wire sw_we_r;
wire cmnd_rd_stb;
wire cmnd_wr_stb;
wire cmnd_ena_stb;
wire cmnd_dis_stb;
wire cmnd_rst_stb;
wire cmnd_ini_stb;
wire cmnd_inc_stb;
wire cmnd_sis_stb;
wire cmnd_tmo_stb;
wire cmnd_cmp_stb;
wire cmnd_issued;
wire ack_error;
wire unsupported_op;
wire [3:0] state_r;
wire [0:0] timer_r;
wire timeout;
wire sim_tmo_r;
wire [4:0] maxaddr;
wire badaddr;
wire igrant;
wire [2:0] stat;
supply0 n1;
supply1 n2;
Q_BUF U0 ( .A(timer_r[0]), .Z(timeout));
Q_BUF U1 ( .A(n2), .Z(stat_datawords[0]));
Q_BUF U2 ( .A(n1), .Z(stat_datawords[1]));
Q_BUF U3 ( .A(n1), .Z(stat_datawords[2]));
Q_BUF U4 ( .A(n1), .Z(stat_datawords[3]));
Q_BUF U5 ( .A(n1), .Z(stat_datawords[4]));
Q_BUF U6 ( .A(n1), .Z(capability_type[0]));
Q_BUF U7 ( .A(n2), .Z(capability_type[1]));
Q_BUF U8 ( .A(n1), .Z(capability_type[2]));
Q_BUF U9 ( .A(n1), .Z(capability_type[3]));
Q_BUF U10 ( .A(n2), .Z(capability_lst[0]));
Q_BUF U11 ( .A(n2), .Z(capability_lst[1]));
Q_BUF U12 ( .A(n1), .Z(capability_lst[2]));
Q_BUF U13 ( .A(n1), .Z(capability_lst[3]));
Q_BUF U14 ( .A(n1), .Z(capability_lst[4]));
Q_BUF U15 ( .A(n2), .Z(capability_lst[5]));
Q_BUF U16 ( .A(n1), .Z(capability_lst[6]));
Q_BUF U17 ( .A(n1), .Z(capability_lst[7]));
Q_BUF U18 ( .A(n1), .Z(capability_lst[8]));
Q_BUF U19 ( .A(n1), .Z(capability_lst[9]));
Q_BUF U20 ( .A(n1), .Z(capability_lst[10]));
Q_BUF U21 ( .A(n1), .Z(capability_lst[11]));
Q_BUF U22 ( .A(n1), .Z(capability_lst[12]));
Q_BUF U23 ( .A(n1), .Z(capability_lst[13]));
Q_BUF U24 ( .A(n1), .Z(capability_lst[14]));
Q_BUF U25 ( .A(n2), .Z(capability_lst[15]));
Q_BUF U26 ( .A(n1), .Z(stat_table_id[0]));
ixc_assign_3 _zz_strnp_7 ( stat[2:0], stat_code[2:0]);
ixc_assign_4 _zz_strnp_1 ( cmnd[3:0], cmnd_op[3:0]);
ixc_assign \genblk1._zz_strnp_0 ( reset, rst_r);
ixc_context_read_6 _zzixc_ctxrd_0 ( { stat_code[2], stat_code[1], 
	stat_code[0], stat[2], stat[1], stat[0]});
ixc_assign _zz_strnp_22 ( _zy_simnet_reset_14_w$, reset);
ixc_assign _zz_strnp_21 ( _zy_simnet_yield_13_w$, yield);
ixc_assign_64 _zz_strnp_20 ( _zy_simnet_sw_wdat_12_w$[0:63], sw_wdat[63:0]);
ixc_assign_5 _zz_strnp_19 ( _zy_simnet_sw_add_11_w$[0:4], sw_add[4:0]);
ixc_assign _zz_strnp_18 ( _zy_simnet_sw_we_10_w$, sw_we);
ixc_assign _zz_strnp_17 ( _zy_simnet_sw_ce_9_w$, sw_ce);
ixc_assign _zz_strnp_16 ( _zy_simnet_sw_cs_8_w$, sw_cs);
ixc_assign_64 _zz_strnp_15 ( _zy_simnet_rd_dat_7_w$[0:63], rd_dat[63:0]);
ixc_assign _zz_strnp_14 ( _zy_simnet_enable_6_w$, enable);
ixc_assign_4 _zz_strnp_13 ( _zy_simnet_capability_type_5_w$[0:3], { n1, n1, 
	n2, n1});
ixc_assign_16 _zz_strnp_12 ( _zy_simnet_capability_lst_4_w$[0:15], { n2, n1, 
	n1, n1, n1, n1, n1, n1, n1, n1, n2, n1, n1, n1, n2, n2});
ixc_assign _zz_strnp_11 ( _zy_simnet_stat_table_id_3_w$, n1);
ixc_assign_5 _zz_strnp_10 ( _zy_simnet_stat_addr_2_w$[0:4], stat_addr[4:0]);
ixc_assign_5 _zz_strnp_9 ( _zy_simnet_stat_datawords_1_w$[0:4], { n1, n1, n1, 
	n1, n2});
ixc_assign_3 _zz_strnp_8 ( _zy_simnet_stat_code_0_w$[0:2], stat_code[2:0]);
ixc_assign_5 _zz_strnp_6 ( stat_addr[4:0], maxaddr[4:0]);
Q_AN02 U47 ( .A0(n19), .A1(grant), .Z(igrant));
Q_AN02 U48 ( .A0(cmnd_issued), .A1(n18), .Z(badaddr));
Q_AO21 U49 ( .A0(n15), .A1(n17), .B0(n14), .Z(n18));
Q_AN02 U50 ( .A0(cmnd_addr[0]), .A1(n16), .Z(n17));
Q_INV U51 ( .A(maxaddr[0]), .Z(n16));
Q_OR03 U52 ( .A0(n11), .A1(n10), .A2(n13), .Z(n14));
Q_OA21 U53 ( .A0(cmnd_addr[1]), .A1(n7), .B0(n9), .Z(n15));
Q_AN03 U54 ( .A0(cmnd_addr[1]), .A1(n7), .A2(n9), .Z(n10));
Q_INV U55 ( .A(maxaddr[1]), .Z(n7));
Q_OA21 U56 ( .A0(cmnd_addr[2]), .A1(n6), .B0(n8), .Z(n9));
Q_AN03 U57 ( .A0(cmnd_addr[2]), .A1(n6), .A2(n8), .Z(n11));
Q_INV U58 ( .A(maxaddr[2]), .Z(n6));
Q_OA21 U59 ( .A0(cmnd_addr[3]), .A1(n5), .B0(n4), .Z(n8));
Q_AN03 U60 ( .A0(cmnd_addr[3]), .A1(n5), .A2(n4), .Z(n12));
Q_INV U61 ( .A(maxaddr[3]), .Z(n5));
Q_OR02 U62 ( .A0(cmnd_addr[4]), .A1(n3), .Z(n4));
Q_AO21 U63 ( .A0(cmnd_addr[4]), .A1(n3), .B0(n12), .Z(n13));
Q_INV U64 ( .A(maxaddr[4]), .Z(n3));
ixc_assign _zz_strnp_5 ( yield, timeout);
ixc_assign _zz_strnp_4 ( sw_we, sw_we_r);
ixc_assign _zz_strnp_3 ( sw_ce, sw_ce_r);
ixc_assign _zz_strnp_2 ( sw_cs, sw_cs_r);
Q_MX02 U69 ( .S(rst_or_ini_r), .A0(cmnd_addr[0]), .A1(rst_addr_r[0]), .Z(sw_add[0]));
Q_MX02 U70 ( .S(rst_or_ini_r), .A0(cmnd_addr[1]), .A1(rst_addr_r[1]), .Z(sw_add[1]));
Q_MX02 U71 ( .S(rst_or_ini_r), .A0(cmnd_addr[2]), .A1(rst_addr_r[2]), .Z(sw_add[2]));
Q_MX02 U72 ( .S(rst_or_ini_r), .A0(cmnd_addr[3]), .A1(rst_addr_r[3]), .Z(sw_add[3]));
Q_MX02 U73 ( .S(rst_or_ini_r), .A0(cmnd_addr[4]), .A1(rst_addr_r[4]), .Z(sw_add[4]));
Q_AN02 U74 ( .A0(enable), .A1(\addr_limit[0][0] ), .Z(maxaddr[0]));
Q_AN02 U75 ( .A0(enable), .A1(\addr_limit[0][1] ), .Z(maxaddr[1]));
Q_AN02 U76 ( .A0(enable), .A1(\addr_limit[0][2] ), .Z(maxaddr[2]));
Q_AN02 U77 ( .A0(enable), .A1(\addr_limit[0][3] ), .Z(maxaddr[3]));
Q_AN02 U78 ( .A0(enable), .A1(\addr_limit[0][4] ), .Z(maxaddr[4]));
Q_INV U79 ( .A(reg_addr[2]), .Z(n20));
Q_INV U80 ( .A(reg_addr[3]), .Z(n21));
Q_INV U81 ( .A(reg_addr[10]), .Z(n22));
Q_OR03 U82 ( .A0(n22), .A1(reg_addr[9]), .A2(reg_addr[8]), .Z(n23));
Q_OR03 U83 ( .A0(reg_addr[7]), .A1(reg_addr[6]), .A2(reg_addr[5]), .Z(n24));
Q_OR03 U84 ( .A0(reg_addr[4]), .A1(n21), .A2(n20), .Z(n25));
Q_OR03 U85 ( .A0(reg_addr[1]), .A1(reg_addr[0]), .A2(n23), .Z(n26));
Q_NR03 U86 ( .A0(n24), .A1(n25), .A2(n26), .Z(n27));
Q_AN02 U87 ( .A0(wr_stb), .A1(n27), .Z(n51));
Q_INV U88 ( .A(n46), .Z(cmnd_issued));
Q_INV U89 ( .A(unsupported_op), .Z(n45));
Q_OA21 U90 ( .A0(n29), .A1(n30), .B0(n28), .Z(unsupported_op));
Q_AN02 U91 ( .A0(n28), .A1(n31), .Z(ack_error));
Q_AO21 U92 ( .A0(n33), .A1(n34), .B0(n32), .Z(n46));
Q_INV U93 ( .A(n51), .Z(n32));
Q_MX02 U94 ( .S(cmnd[3]), .A0(n37), .A1(n35), .Z(n33));
Q_INV U95 ( .A(cmnd_cmp_stb), .Z(n47));
Q_AN02 U96 ( .A0(n28), .A1(n38), .Z(cmnd_cmp_stb));
Q_AN02 U97 ( .A0(n28), .A1(n39), .Z(cmnd_tmo_stb));
Q_AN03 U98 ( .A0(n28), .A1(n34), .A2(n37), .Z(cmnd_sis_stb));
Q_AN02 U99 ( .A0(n51), .A1(cmnd[3]), .Z(n28));
Q_AN02 U100 ( .A0(n40), .A1(n31), .Z(cmnd_inc_stb));
Q_AN02 U101 ( .A0(n35), .A1(cmnd[0]), .Z(n31));
Q_AN02 U102 ( .A0(n40), .A1(n39), .Z(cmnd_ini_stb));
Q_AN02 U103 ( .A0(n35), .A1(n34), .Z(n39));
Q_AN02 U104 ( .A0(cmnd[2]), .A1(cmnd[1]), .Z(n35));
Q_INV U105 ( .A(cmnd_rst_stb), .Z(n48));
Q_AN02 U106 ( .A0(n30), .A1(n41), .Z(cmnd_rst_stb));
Q_AN02 U107 ( .A0(n40), .A1(cmnd[0]), .Z(n41));
Q_AN02 U108 ( .A0(n30), .A1(n42), .Z(cmnd_dis_stb));
Q_AN02 U109 ( .A0(n40), .A1(n34), .Z(n42));
Q_AN02 U110 ( .A0(cmnd[2]), .A1(n43), .Z(n30));
Q_AN02 U111 ( .A0(n29), .A1(n41), .Z(cmnd_ena_stb));
Q_INV U112 ( .A(cmnd_wr_stb), .Z(n49));
Q_AN02 U113 ( .A0(n29), .A1(n42), .Z(cmnd_wr_stb));
Q_INV U114 ( .A(cmnd[0]), .Z(n34));
Q_AN02 U115 ( .A0(n44), .A1(cmnd[1]), .Z(n29));
Q_INV U116 ( .A(cmnd_rd_stb), .Z(n50));
Q_AN02 U117 ( .A0(n40), .A1(n38), .Z(cmnd_rd_stb));
Q_AN02 U118 ( .A0(n37), .A1(cmnd[0]), .Z(n38));
Q_NR02 U119 ( .A0(cmnd[2]), .A1(cmnd[1]), .Z(n37));
Q_INV U120 ( .A(cmnd[1]), .Z(n43));
Q_INV U121 ( .A(cmnd[2]), .Z(n44));
Q_AN02 U122 ( .A0(n51), .A1(n36), .Z(n40));
Q_INV U123 ( .A(cmnd[3]), .Z(n36));
Q_OR02 U124 ( .A0(cmnd_ini_stb), .A1(cmnd_inc_stb), .Z(n383));
Q_XNR2 U125 ( .A0(rst_addr_r[0]), .A1(cmnd_addr[0]), .Z(n53));
Q_XNR2 U126 ( .A0(rst_addr_r[1]), .A1(cmnd_addr[1]), .Z(n54));
Q_XNR2 U127 ( .A0(rst_addr_r[2]), .A1(cmnd_addr[2]), .Z(n55));
Q_XNR2 U128 ( .A0(rst_addr_r[3]), .A1(cmnd_addr[3]), .Z(n56));
Q_XNR2 U129 ( .A0(rst_addr_r[4]), .A1(cmnd_addr[4]), .Z(n57));
Q_AN03 U130 ( .A0(n57), .A1(n56), .A2(n55), .Z(n58));
Q_AN03 U131 ( .A0(n54), .A1(n53), .A2(n58), .Z(n384));
Q_AN02 U132 ( .A0(init_inc_r), .A1(igrant), .Z(n59));
Q_XOR2 U133 ( .A0(inc_r[0]), .A1(n59), .Z(n60));
Q_AD01HF U134 ( .A0(rst_addr_r[0]), .B0(igrant), .S(n61), .CO(n62));
Q_AD01HF U135 ( .A0(rst_addr_r[1]), .B0(n62), .S(n63), .CO(n64));
Q_AD01HF U136 ( .A0(rst_addr_r[2]), .B0(n64), .S(n65), .CO(n66));
Q_AD01HF U137 ( .A0(rst_addr_r[3]), .B0(n66), .S(n67), .CO(n68));
Q_XOR2 U138 ( .A0(rst_addr_r[4]), .A1(n68), .Z(n69));
Q_MX02 U139 ( .S(n302), .A0(n75), .A1(n71), .Z(n70));
Q_ND02 U140 ( .A0(n72), .A1(n73), .Z(n71));
Q_ND02 U141 ( .A0(n361), .A1(n267), .Z(n73));
Q_OR02 U142 ( .A0(n74), .A1(n267), .Z(n72));
Q_OR02 U143 ( .A0(n267), .A1(n363), .Z(n75));
Q_INV U144 ( .A(n76), .Z(n77));
Q_MX02 U145 ( .S(n302), .A0(n72), .A1(n78), .Z(n76));
Q_INV U146 ( .A(n79), .Z(n78));
Q_INV U147 ( .A(n80), .Z(n81));
Q_MX02 U148 ( .S(n302), .A0(n87), .A1(n82), .Z(n80));
Q_INV U149 ( .A(n83), .Z(n82));
Q_MX02 U150 ( .S(n267), .A0(n79), .A1(n84), .Z(n83));
Q_INV U151 ( .A(n85), .Z(n84));
Q_XOR2 U152 ( .A0(n361), .A1(n86), .Z(n79));
Q_OR02 U153 ( .A0(n362), .A1(n74), .Z(n87));
Q_OR02 U154 ( .A0(n361), .A1(n363), .Z(n74));
Q_NR02 U155 ( .A0(n364), .A1(n89), .Z(n88));
Q_MX02 U156 ( .S(n267), .A0(n85), .A1(n363), .Z(n89));
Q_OR02 U157 ( .A0(n361), .A1(n86), .Z(n85));
Q_INV U158 ( .A(n363), .Z(n86));
Q_AN03 U159 ( .A0(n362), .A1(n361), .A2(n364), .Z(n90));
Q_AO21 U160 ( .A0(n90), .A1(state_r[3]), .B0(n88), .Z(n388));
Q_AO21 U161 ( .A0(n90), .A1(state_r[2]), .B0(n81), .Z(n387));
Q_AO21 U162 ( .A0(n90), .A1(state_r[1]), .B0(n77), .Z(n386));
Q_AO21 U163 ( .A0(n90), .A1(state_r[0]), .B0(n70), .Z(n385));
Q_AN02 U164 ( .A0(n366), .A1(cmnd_addr[0]), .Z(n92));
Q_MX02 U165 ( .S(n367), .A0(n92), .A1(n61), .Z(n93));
Q_AN02 U166 ( .A0(n366), .A1(cmnd_addr[1]), .Z(n94));
Q_MX02 U167 ( .S(n367), .A0(n94), .A1(n63), .Z(n95));
Q_AN02 U168 ( .A0(n366), .A1(cmnd_addr[2]), .Z(n96));
Q_MX02 U169 ( .S(n367), .A0(n96), .A1(n65), .Z(n97));
Q_AN02 U170 ( .A0(n366), .A1(cmnd_addr[3]), .Z(n98));
Q_MX02 U171 ( .S(n367), .A0(n98), .A1(n67), .Z(n99));
Q_AN02 U172 ( .A0(n366), .A1(cmnd_addr[4]), .Z(n100));
Q_MX02 U173 ( .S(n367), .A0(n100), .A1(n69), .Z(n101));
Q_AN02 U174 ( .A0(n372), .A1(n60), .Z(n102));
Q_MX03 U175 ( .S0(n374), .S1(n375), .A0(sw_aindex[0]), .A1(wr_dat[0]), .A2(sw_rdat[0]), .Z(n103));
Q_MX03 U176 ( .S0(n374), .S1(n375), .A0(sw_aindex[1]), .A1(wr_dat[1]), .A2(sw_rdat[1]), .Z(n104));
Q_MX03 U177 ( .S0(n374), .S1(n375), .A0(sw_aindex[2]), .A1(wr_dat[2]), .A2(sw_rdat[2]), .Z(n105));
Q_MX03 U178 ( .S0(n374), .S1(n375), .A0(sw_aindex[3]), .A1(wr_dat[3]), .A2(sw_rdat[3]), .Z(n106));
Q_MX03 U179 ( .S0(n374), .S1(n375), .A0(sw_match), .A1(wr_dat[4]), .A2(sw_rdat[4]), .Z(n107));
Q_AN02 U180 ( .A0(n374), .A1(wr_dat[5]), .Z(n108));
Q_MX02 U181 ( .S(n375), .A0(n108), .A1(sw_rdat[5]), .Z(n109));
Q_AN02 U182 ( .A0(n374), .A1(wr_dat[6]), .Z(n110));
Q_MX02 U183 ( .S(n375), .A0(n110), .A1(sw_rdat[6]), .Z(n111));
Q_AN02 U184 ( .A0(n374), .A1(wr_dat[7]), .Z(n112));
Q_MX02 U185 ( .S(n375), .A0(n112), .A1(sw_rdat[7]), .Z(n113));
Q_AN02 U186 ( .A0(n374), .A1(wr_dat[8]), .Z(n114));
Q_MX02 U187 ( .S(n375), .A0(n114), .A1(sw_rdat[8]), .Z(n115));
Q_AN02 U188 ( .A0(n374), .A1(wr_dat[9]), .Z(n116));
Q_MX02 U189 ( .S(n375), .A0(n116), .A1(sw_rdat[9]), .Z(n117));
Q_AN02 U190 ( .A0(n374), .A1(wr_dat[10]), .Z(n118));
Q_MX02 U191 ( .S(n375), .A0(n118), .A1(sw_rdat[10]), .Z(n119));
Q_AN02 U192 ( .A0(n374), .A1(wr_dat[11]), .Z(n120));
Q_MX02 U193 ( .S(n375), .A0(n120), .A1(sw_rdat[11]), .Z(n121));
Q_AN02 U194 ( .A0(n374), .A1(wr_dat[12]), .Z(n122));
Q_MX02 U195 ( .S(n375), .A0(n122), .A1(sw_rdat[12]), .Z(n123));
Q_AN02 U196 ( .A0(n374), .A1(wr_dat[13]), .Z(n124));
Q_MX02 U197 ( .S(n375), .A0(n124), .A1(sw_rdat[13]), .Z(n125));
Q_AN02 U198 ( .A0(n374), .A1(wr_dat[14]), .Z(n126));
Q_MX02 U199 ( .S(n375), .A0(n126), .A1(sw_rdat[14]), .Z(n127));
Q_AN02 U200 ( .A0(n374), .A1(wr_dat[15]), .Z(n128));
Q_MX02 U201 ( .S(n375), .A0(n128), .A1(sw_rdat[15]), .Z(n129));
Q_AN02 U202 ( .A0(n374), .A1(wr_dat[16]), .Z(n130));
Q_MX02 U203 ( .S(n375), .A0(n130), .A1(sw_rdat[16]), .Z(n131));
Q_AN02 U204 ( .A0(n374), .A1(wr_dat[17]), .Z(n132));
Q_MX02 U205 ( .S(n375), .A0(n132), .A1(sw_rdat[17]), .Z(n133));
Q_AN02 U206 ( .A0(n374), .A1(wr_dat[18]), .Z(n134));
Q_MX02 U207 ( .S(n375), .A0(n134), .A1(sw_rdat[18]), .Z(n135));
Q_AN02 U208 ( .A0(n374), .A1(wr_dat[19]), .Z(n136));
Q_MX02 U209 ( .S(n375), .A0(n136), .A1(sw_rdat[19]), .Z(n137));
Q_AN02 U210 ( .A0(n374), .A1(wr_dat[20]), .Z(n138));
Q_MX02 U211 ( .S(n375), .A0(n138), .A1(sw_rdat[20]), .Z(n139));
Q_AN02 U212 ( .A0(n374), .A1(wr_dat[21]), .Z(n140));
Q_MX02 U213 ( .S(n375), .A0(n140), .A1(sw_rdat[21]), .Z(n141));
Q_AN02 U214 ( .A0(n374), .A1(wr_dat[22]), .Z(n142));
Q_MX02 U215 ( .S(n375), .A0(n142), .A1(sw_rdat[22]), .Z(n143));
Q_AN02 U216 ( .A0(n374), .A1(wr_dat[23]), .Z(n144));
Q_MX02 U217 ( .S(n375), .A0(n144), .A1(sw_rdat[23]), .Z(n145));
Q_AN02 U218 ( .A0(n374), .A1(wr_dat[24]), .Z(n146));
Q_MX02 U219 ( .S(n375), .A0(n146), .A1(sw_rdat[24]), .Z(n147));
Q_AN02 U220 ( .A0(n374), .A1(wr_dat[25]), .Z(n148));
Q_MX02 U221 ( .S(n375), .A0(n148), .A1(sw_rdat[25]), .Z(n149));
Q_AN02 U222 ( .A0(n374), .A1(wr_dat[26]), .Z(n150));
Q_MX02 U223 ( .S(n375), .A0(n150), .A1(sw_rdat[26]), .Z(n151));
Q_AN02 U224 ( .A0(n374), .A1(wr_dat[27]), .Z(n152));
Q_MX02 U225 ( .S(n375), .A0(n152), .A1(sw_rdat[27]), .Z(n153));
Q_AN02 U226 ( .A0(n374), .A1(wr_dat[28]), .Z(n154));
Q_MX02 U227 ( .S(n375), .A0(n154), .A1(sw_rdat[28]), .Z(n155));
Q_AN02 U228 ( .A0(n374), .A1(wr_dat[29]), .Z(n156));
Q_MX02 U229 ( .S(n375), .A0(n156), .A1(sw_rdat[29]), .Z(n157));
Q_AN02 U230 ( .A0(n374), .A1(wr_dat[30]), .Z(n158));
Q_MX02 U231 ( .S(n375), .A0(n158), .A1(sw_rdat[30]), .Z(n159));
Q_AN02 U232 ( .A0(n374), .A1(wr_dat[31]), .Z(n160));
Q_MX02 U233 ( .S(n375), .A0(n160), .A1(sw_rdat[31]), .Z(n161));
Q_AN02 U234 ( .A0(n374), .A1(wr_dat[32]), .Z(n162));
Q_MX02 U235 ( .S(n375), .A0(n162), .A1(sw_rdat[32]), .Z(n163));
Q_AN02 U236 ( .A0(n374), .A1(wr_dat[33]), .Z(n164));
Q_MX02 U237 ( .S(n375), .A0(n164), .A1(sw_rdat[33]), .Z(n165));
Q_AN02 U238 ( .A0(n374), .A1(wr_dat[34]), .Z(n166));
Q_MX02 U239 ( .S(n375), .A0(n166), .A1(sw_rdat[34]), .Z(n167));
Q_AN02 U240 ( .A0(n374), .A1(wr_dat[35]), .Z(n168));
Q_MX02 U241 ( .S(n375), .A0(n168), .A1(sw_rdat[35]), .Z(n169));
Q_AN02 U242 ( .A0(n374), .A1(wr_dat[36]), .Z(n170));
Q_MX02 U243 ( .S(n375), .A0(n170), .A1(sw_rdat[36]), .Z(n171));
Q_AN02 U244 ( .A0(n374), .A1(wr_dat[37]), .Z(n172));
Q_MX02 U245 ( .S(n375), .A0(n172), .A1(sw_rdat[37]), .Z(n173));
Q_AN02 U246 ( .A0(n374), .A1(wr_dat[38]), .Z(n174));
Q_MX02 U247 ( .S(n375), .A0(n174), .A1(sw_rdat[38]), .Z(n175));
Q_AN02 U248 ( .A0(n374), .A1(wr_dat[39]), .Z(n176));
Q_MX02 U249 ( .S(n375), .A0(n176), .A1(sw_rdat[39]), .Z(n177));
Q_AN02 U250 ( .A0(n374), .A1(wr_dat[40]), .Z(n178));
Q_MX02 U251 ( .S(n375), .A0(n178), .A1(sw_rdat[40]), .Z(n179));
Q_AN02 U252 ( .A0(n374), .A1(wr_dat[41]), .Z(n180));
Q_MX02 U253 ( .S(n375), .A0(n180), .A1(sw_rdat[41]), .Z(n181));
Q_AN02 U254 ( .A0(n374), .A1(wr_dat[42]), .Z(n182));
Q_MX02 U255 ( .S(n375), .A0(n182), .A1(sw_rdat[42]), .Z(n183));
Q_AN02 U256 ( .A0(n374), .A1(wr_dat[43]), .Z(n184));
Q_MX02 U257 ( .S(n375), .A0(n184), .A1(sw_rdat[43]), .Z(n185));
Q_AN02 U258 ( .A0(n374), .A1(wr_dat[44]), .Z(n186));
Q_MX02 U259 ( .S(n375), .A0(n186), .A1(sw_rdat[44]), .Z(n187));
Q_AN02 U260 ( .A0(n374), .A1(wr_dat[45]), .Z(n188));
Q_MX02 U261 ( .S(n375), .A0(n188), .A1(sw_rdat[45]), .Z(n189));
Q_AN02 U262 ( .A0(n374), .A1(wr_dat[46]), .Z(n190));
Q_MX02 U263 ( .S(n375), .A0(n190), .A1(sw_rdat[46]), .Z(n191));
Q_AN02 U264 ( .A0(n374), .A1(wr_dat[47]), .Z(n192));
Q_MX02 U265 ( .S(n375), .A0(n192), .A1(sw_rdat[47]), .Z(n193));
Q_AN02 U266 ( .A0(n374), .A1(wr_dat[48]), .Z(n194));
Q_MX02 U267 ( .S(n375), .A0(n194), .A1(sw_rdat[48]), .Z(n195));
Q_AN02 U268 ( .A0(n374), .A1(wr_dat[49]), .Z(n196));
Q_MX02 U269 ( .S(n375), .A0(n196), .A1(sw_rdat[49]), .Z(n197));
Q_AN02 U270 ( .A0(n374), .A1(wr_dat[50]), .Z(n198));
Q_MX02 U271 ( .S(n375), .A0(n198), .A1(sw_rdat[50]), .Z(n199));
Q_AN02 U272 ( .A0(n374), .A1(wr_dat[51]), .Z(n200));
Q_MX02 U273 ( .S(n375), .A0(n200), .A1(sw_rdat[51]), .Z(n201));
Q_AN02 U274 ( .A0(n374), .A1(wr_dat[52]), .Z(n202));
Q_MX02 U275 ( .S(n375), .A0(n202), .A1(sw_rdat[52]), .Z(n203));
Q_AN02 U276 ( .A0(n374), .A1(wr_dat[53]), .Z(n204));
Q_MX02 U277 ( .S(n375), .A0(n204), .A1(sw_rdat[53]), .Z(n205));
Q_AN02 U278 ( .A0(n374), .A1(wr_dat[54]), .Z(n206));
Q_MX02 U279 ( .S(n375), .A0(n206), .A1(sw_rdat[54]), .Z(n207));
Q_AN02 U280 ( .A0(n374), .A1(wr_dat[55]), .Z(n208));
Q_MX02 U281 ( .S(n375), .A0(n208), .A1(sw_rdat[55]), .Z(n209));
Q_AN02 U282 ( .A0(n374), .A1(wr_dat[56]), .Z(n210));
Q_MX02 U283 ( .S(n375), .A0(n210), .A1(sw_rdat[56]), .Z(n211));
Q_AN02 U284 ( .A0(n374), .A1(wr_dat[57]), .Z(n212));
Q_MX02 U285 ( .S(n375), .A0(n212), .A1(sw_rdat[57]), .Z(n213));
Q_AN02 U286 ( .A0(n374), .A1(wr_dat[58]), .Z(n214));
Q_MX02 U287 ( .S(n375), .A0(n214), .A1(sw_rdat[58]), .Z(n215));
Q_AN02 U288 ( .A0(n374), .A1(wr_dat[59]), .Z(n216));
Q_MX02 U289 ( .S(n375), .A0(n216), .A1(sw_rdat[59]), .Z(n217));
Q_AN02 U290 ( .A0(n374), .A1(wr_dat[60]), .Z(n218));
Q_MX02 U291 ( .S(n375), .A0(n218), .A1(sw_rdat[60]), .Z(n219));
Q_AN02 U292 ( .A0(n374), .A1(wr_dat[61]), .Z(n220));
Q_MX02 U293 ( .S(n375), .A0(n220), .A1(sw_rdat[61]), .Z(n221));
Q_AN02 U294 ( .A0(n374), .A1(wr_dat[62]), .Z(n222));
Q_MX02 U295 ( .S(n375), .A0(n222), .A1(sw_rdat[62]), .Z(n223));
Q_AN02 U296 ( .A0(n374), .A1(wr_dat[63]), .Z(n224));
Q_MX02 U297 ( .S(n375), .A0(n224), .A1(sw_rdat[63]), .Z(n225));
Q_FDP1 \state_r_REG[3] ( .CK(clk), .R(rst_n), .D(n388), .Q(state_r[3]), .QN(n242));
Q_FDP1 \state_r_REG[2] ( .CK(clk), .R(rst_n), .D(n387), .Q(state_r[2]), .QN(n350));
Q_FDP1 \state_r_REG[1] ( .CK(clk), .R(rst_n), .D(n386), .Q(state_r[1]), .QN(n258));
Q_FDP2 \state_r_REG[0] ( .CK(clk), .S(rst_n), .D(n385), .Q(state_r[0]), .QN(n247));
Q_FDP1 \timer_r_REG[0] ( .CK(clk), .R(rst_n), .D(n91), .Q(timer_r[0]), .QN(n52));
Q_ND02 U303 ( .A0(n227), .A1(n228), .Z(n226));
Q_ND02 U304 ( .A0(n229), .A1(n333), .Z(n228));
Q_OR02 U305 ( .A0(n230), .A1(n377), .Z(n229));
Q_INV U306 ( .A(n376), .Z(n230));
Q_ND02 U307 ( .A0(n227), .A1(n232), .Z(n231));
Q_ND02 U308 ( .A0(n376), .A1(n333), .Z(n232));
Q_OR03 U309 ( .A0(n376), .A1(n377), .A2(n333), .Z(n227));
Q_MX02 U310 ( .S(n333), .A0(n376), .A1(n377), .Z(n233));
Q_FDP1 sw_cs_r_REG  ( .CK(clk), .R(rst_n), .D(n371), .Q(sw_cs_r), .QN( ));
Q_FDP1 sw_ce_r_REG  ( .CK(clk), .R(rst_n), .D(n370), .Q(sw_ce_r), .QN( ));
Q_FDP1 rst_r_REG  ( .CK(clk), .R(rst_n), .D(n369), .Q(rst_r), .QN(n389));
Q_FDP1 rst_or_ini_r_REG  ( .CK(clk), .R(rst_n), .D(n368), .Q(rst_or_ini_r), .QN( ));
Q_FDP1 sw_we_r_REG  ( .CK(clk), .R(rst_n), .D(n365), .Q(sw_we_r), .QN( ));
Q_OA21 U316 ( .A0(n235), .A1(n236), .B0(n234), .Z(n361));
Q_OR03 U317 ( .A0(n238), .A1(n239), .A2(n237), .Z(n236));
Q_AN03 U318 ( .A0(n242), .A1(n243), .A2(n240), .Z(n241));
Q_AN02 U319 ( .A0(n49), .A1(cmnd_rd_stb), .Z(n243));
Q_AO21 U320 ( .A0(n242), .A1(n244), .B0(n241), .Z(n239));
Q_AN02 U321 ( .A0(n245), .A1(n246), .Z(n244));
Q_NR02 U322 ( .A0(state_r[0]), .A1(cmnd_ena_stb), .Z(n246));
Q_OA21 U323 ( .A0(n249), .A1(n250), .B0(n248), .Z(n238));
Q_AN03 U324 ( .A0(state_r[3]), .A1(n252), .A2(n251), .Z(n250));
Q_OA21 U325 ( .A0(n254), .A1(n255), .B0(n253), .Z(n249));
Q_NR02 U326 ( .A0(n259), .A1(igrant), .Z(n255));
Q_AN02 U327 ( .A0(n256), .A1(n257), .Z(n254));
Q_INV U328 ( .A(n384), .Z(n257));
Q_NR02 U329 ( .A0(state_r[1]), .A1(state_r[0]), .Z(n256));
Q_AN03 U330 ( .A0(n263), .A1(n47), .A2(n261), .Z(n262));
Q_AN02 U331 ( .A0(cmnd_rst_stb), .A1(n242), .Z(n263));
Q_OR03 U332 ( .A0(n264), .A1(n262), .A2(n260), .Z(n235));
Q_AN03 U333 ( .A0(n265), .A1(n266), .A2(n251), .Z(n264));
Q_INV U334 ( .A(n267), .Z(n362));
Q_OA21 U335 ( .A0(n268), .A1(n237), .B0(n234), .Z(n267));
Q_AO21 U336 ( .A0(n240), .A1(n270), .B0(n269), .Z(n268));
Q_AN02 U337 ( .A0(n242), .A1(cmnd_wr_stb), .Z(n270));
Q_AN02 U338 ( .A0(n272), .A1(n273), .Z(n274));
Q_NR02 U339 ( .A0(state_r[3]), .A1(n353), .Z(n273));
Q_MX02 U340 ( .S(state_r[1]), .A0(cmnd_ena_stb), .A1(n276), .Z(n272));
Q_OR03 U341 ( .A0(n277), .A1(n274), .A2(n271), .Z(n237));
Q_AN02 U342 ( .A0(n52), .A1(n46), .Z(n248));
Q_AN03 U343 ( .A0(n279), .A1(n280), .A2(n278), .Z(n277));
Q_NR02 U344 ( .A0(cmnd_dis_stb), .A1(unsupported_op), .Z(n280));
Q_OA21 U345 ( .A0(n281), .A1(n282), .B0(n248), .Z(n271));
Q_OA21 U346 ( .A0(n283), .A1(n284), .B0(state_r[3]), .Z(n282));
Q_AN02 U347 ( .A0(state_r[2]), .A1(n276), .Z(n284));
Q_AN02 U348 ( .A0(n253), .A1(igrant), .Z(n286));
Q_AN02 U349 ( .A0(n242), .A1(state_r[2]), .Z(n253));
Q_AO21 U350 ( .A0(n287), .A1(n259), .B0(n285), .Z(n281));
Q_OA21 U351 ( .A0(state_r[0]), .A1(n288), .B0(n286), .Z(n285));
Q_AN02 U352 ( .A0(n258), .A1(n384), .Z(n288));
Q_OR02 U353 ( .A0(n242), .A1(n276), .Z(n287));
Q_AN02 U354 ( .A0(ack_error), .A1(enable), .Z(n276));
Q_OA21 U355 ( .A0(n289), .A1(n290), .B0(n245), .Z(n269));
Q_AN02 U356 ( .A0(n292), .A1(n47), .Z(n291));
Q_AN03 U357 ( .A0(n293), .A1(n294), .A2(n291), .Z(n290));
Q_AN02 U358 ( .A0(n242), .A1(state_r[0]), .Z(n293));
Q_AN02 U359 ( .A0(n295), .A1(n296), .Z(n289));
Q_AN03 U360 ( .A0(n298), .A1(n299), .A2(n297), .Z(n363));
Q_AO21 U361 ( .A0(n292), .A1(n301), .B0(n300), .Z(n297));
Q_INV U362 ( .A(n300), .Z(n301));
Q_INV U363 ( .A(n302), .Z(n364));
Q_OA21 U364 ( .A0(n303), .A1(n260), .B0(n234), .Z(n302));
Q_AN03 U365 ( .A0(n300), .A1(n242), .A2(n299), .Z(n304));
Q_AN02 U366 ( .A0(n240), .A1(n49), .Z(n299));
Q_AO21 U367 ( .A0(n50), .A1(cmnd_cmp_stb), .B0(cmnd_rd_stb), .Z(n300));
Q_AN03 U368 ( .A0(n292), .A1(n306), .A2(n261), .Z(n305));
Q_NR02 U369 ( .A0(state_r[3]), .A1(cmnd_cmp_stb), .Z(n306));
Q_AO21 U370 ( .A0(n48), .A1(n383), .B0(cmnd_rst_stb), .Z(n292));
Q_AN02 U371 ( .A0(n295), .A1(n46), .Z(n308));
Q_AN03 U372 ( .A0(n265), .A1(n245), .A2(n308), .Z(n309));
Q_OR03 U373 ( .A0(n309), .A1(n307), .A2(n304), .Z(n303));
Q_AO21 U374 ( .A0(n310), .A1(n311), .B0(n305), .Z(n307));
Q_AN02 U375 ( .A0(igrant), .A1(n46), .Z(n266));
Q_AN02 U376 ( .A0(n312), .A1(n266), .Z(n310));
Q_AN02 U377 ( .A0(n313), .A1(n247), .Z(n311));
Q_NR02 U378 ( .A0(timeout), .A1(state_r[3]), .Z(n313));
Q_AN02 U379 ( .A0(ack_error), .A1(init_r), .Z(n315));
Q_AO21 U380 ( .A0(n278), .A1(n316), .B0(n314), .Z(n260));
Q_AN02 U381 ( .A0(n279), .A1(cmnd_dis_stb), .Z(n316));
Q_NR02 U382 ( .A0(cmnd_cmp_stb), .A1(n383), .Z(n279));
Q_AN02 U383 ( .A0(n317), .A1(n261), .Z(n278));
Q_AN02 U384 ( .A0(n240), .A1(n294), .Z(n261));
Q_NR02 U385 ( .A0(cmnd_wr_stb), .A1(cmnd_rd_stb), .Z(n294));
Q_NR02 U386 ( .A0(cmnd_rst_stb), .A1(state_r[3]), .Z(n317));
Q_OA21 U387 ( .A0(n318), .A1(n319), .B0(n315), .Z(n314));
Q_AN02 U388 ( .A0(n265), .A1(n46), .Z(n296));
Q_AN02 U389 ( .A0(n52), .A1(state_r[3]), .Z(n265));
Q_OA21 U390 ( .A0(state_r[2]), .A1(n259), .B0(n296), .Z(n318));
Q_AN02 U391 ( .A0(state_r[1]), .A1(state_r[0]), .Z(n259));
Q_AO21 U392 ( .A0(n247), .A1(igrant), .B0(state_r[0]), .Z(n295));
Q_AN03 U393 ( .A0(n252), .A1(n371), .A2(n52), .Z(n91));
Q_INV U394 ( .A(igrant), .Z(n252));
Q_OA21 U395 ( .A0(n321), .A1(n322), .B0(n320), .Z(n365));
Q_AN02 U396 ( .A0(cmnd_sis_stb), .A1(n323), .Z(n366));
Q_INV U397 ( .A(n367), .Z(n323));
Q_OA21 U398 ( .A0(n321), .A1(n324), .B0(n320), .Z(n368));
Q_AN02 U399 ( .A0(n322), .A1(n325), .Z(n324));
Q_AN02 U400 ( .A0(n387), .A1(n326), .Z(n322));
Q_AN02 U401 ( .A0(n320), .A1(n321), .Z(n369));
Q_AN02 U402 ( .A0(n327), .A1(n385), .Z(n321));
Q_OR03 U403 ( .A0(n369), .A1(n328), .A2(n370), .Z(n371));
Q_AN02 U404 ( .A0(n388), .A1(n329), .Z(n370));
Q_AN03 U405 ( .A0(n320), .A1(n387), .A2(n330), .Z(n328));
Q_INV U406 ( .A(n331), .Z(n330));
Q_INV U407 ( .A(n332), .Z(n372));
Q_AN02 U408 ( .A0(n312), .A1(n293), .Z(n375));
Q_AN02 U409 ( .A0(state_r[2]), .A1(state_r[1]), .Z(n312));
Q_AN02 U410 ( .A0(n335), .A1(n336), .Z(n337));
Q_INV U411 ( .A(n338), .Z(n335));
Q_OR03 U412 ( .A0(n339), .A1(n337), .A2(n334), .Z(n333));
Q_AN03 U413 ( .A0(n341), .A1(n45), .A2(n340), .Z(n334));
Q_OR02 U414 ( .A0(n331), .A1(n342), .Z(n339));
Q_AN02 U415 ( .A0(n386), .A1(n385), .Z(n331));
Q_INV U416 ( .A(n343), .Z(n342));
Q_AN02 U417 ( .A0(n320), .A1(n344), .Z(n336));
Q_NR02 U418 ( .A0(n387), .A1(n385), .Z(n344));
Q_OA21 U419 ( .A0(n346), .A1(n326), .B0(n336), .Z(n376));
Q_AN02 U420 ( .A0(n45), .A1(n386), .Z(n338));
Q_OA21 U421 ( .A0(n341), .A1(badaddr), .B0(n338), .Z(n346));
Q_AN02 U422 ( .A0(timeout), .A1(n234), .Z(n341));
Q_NR02 U423 ( .A0(n388), .A1(n387), .Z(n343));
Q_OA21 U424 ( .A0(n347), .A1(n326), .B0(n343), .Z(n377));
Q_AN03 U425 ( .A0(n386), .A1(n325), .A2(unsupported_op), .Z(n347));
Q_ND02 U426 ( .A0(n319), .A1(n340), .Z(n348));
Q_AN02 U427 ( .A0(n327), .A1(n349), .Z(n340));
Q_NR02 U428 ( .A0(n388), .A1(n385), .Z(n349));
Q_AN02 U429 ( .A0(n345), .A1(n386), .Z(n327));
Q_AN02 U430 ( .A0(n242), .A1(n283), .Z(n319));
Q_AN03 U431 ( .A0(n350), .A1(state_r[1]), .A2(n247), .Z(n283));
Q_OA21 U432 ( .A0(n374), .A1(n351), .B0(n234), .Z(n378));
Q_AN02 U433 ( .A0(n352), .A1(state_r[1]), .Z(n351));
Q_INV U434 ( .A(n373), .Z(n374));
Q_AN02 U435 ( .A0(n245), .A1(n247), .Z(n251));
Q_MX02 U436 ( .S(state_r[3]), .A0(n354), .A1(n275), .Z(n352));
Q_INV U437 ( .A(n353), .Z(n275));
Q_AN02 U438 ( .A0(state_r[2]), .A1(state_r[0]), .Z(n354));
Q_AN03 U439 ( .A0(n373), .A1(n320), .A2(n329), .Z(n355));
Q_AN02 U440 ( .A0(n356), .A1(n325), .Z(n329));
Q_INV U441 ( .A(n385), .Z(n325));
Q_NR02 U442 ( .A0(n387), .A1(n386), .Z(n356));
Q_INV U443 ( .A(n386), .Z(n326));
Q_INV U444 ( .A(n387), .Z(n345));
Q_INV U445 ( .A(n388), .Z(n320));
Q_AO21 U446 ( .A0(n298), .A1(n357), .B0(n355), .Z(n379));
Q_AN03 U447 ( .A0(n247), .A1(cmnd_ena_stb), .A2(n245), .Z(n357));
Q_OR03 U448 ( .A0(state_r[3]), .A1(state_r[1]), .A2(n353), .Z(n373));
Q_OR02 U449 ( .A0(state_r[2]), .A1(state_r[0]), .Z(n353));
Q_AN03 U450 ( .A0(n298), .A1(n258), .A2(n358), .Z(n380));
Q_AO21 U451 ( .A0(state_r[2]), .A1(n247), .B0(n332), .Z(n358));
Q_AN02 U452 ( .A0(n350), .A1(state_r[0]), .Z(n332));
Q_ND02 U453 ( .A0(n298), .A1(n240), .Z(n381));
Q_AN02 U454 ( .A0(n245), .A1(state_r[0]), .Z(n240));
Q_NR02 U455 ( .A0(state_r[2]), .A1(state_r[1]), .Z(n245));
Q_AN02 U456 ( .A0(n298), .A1(n247), .Z(n359));
Q_AN03 U457 ( .A0(state_r[2]), .A1(n258), .A2(n359), .Z(n367));
Q_NR02 U458 ( .A0(badaddr), .A1(state_r[3]), .Z(n298));
Q_INV U459 ( .A(badaddr), .Z(n234));
Q_OR03 U460 ( .A0(cmnd_rst_stb), .A1(cmnd_sis_stb), .A2(n367), .Z(n382));
Q_OR02 U461 ( .A0(cmnd_tmo_stb), .A1(timeout), .Z(n360));
Q_AN02 U462 ( .A0(n389), .A1(wr_dat[0]), .Z(sw_wdat[0]));
Q_AN02 U463 ( .A0(n389), .A1(wr_dat[1]), .Z(sw_wdat[1]));
Q_AN02 U464 ( .A0(n389), .A1(wr_dat[2]), .Z(sw_wdat[2]));
Q_AN02 U465 ( .A0(n389), .A1(wr_dat[3]), .Z(sw_wdat[3]));
Q_AN02 U466 ( .A0(n389), .A1(wr_dat[4]), .Z(sw_wdat[4]));
Q_AN02 U467 ( .A0(n389), .A1(wr_dat[5]), .Z(sw_wdat[5]));
Q_AN02 U468 ( .A0(n389), .A1(wr_dat[6]), .Z(sw_wdat[6]));
Q_AN02 U469 ( .A0(n389), .A1(wr_dat[7]), .Z(sw_wdat[7]));
Q_AN02 U470 ( .A0(n389), .A1(wr_dat[8]), .Z(sw_wdat[8]));
Q_AN02 U471 ( .A0(n389), .A1(wr_dat[9]), .Z(sw_wdat[9]));
Q_AN02 U472 ( .A0(n389), .A1(wr_dat[10]), .Z(sw_wdat[10]));
Q_AN02 U473 ( .A0(n389), .A1(wr_dat[11]), .Z(sw_wdat[11]));
Q_AN02 U474 ( .A0(n389), .A1(wr_dat[12]), .Z(sw_wdat[12]));
Q_AN02 U475 ( .A0(n389), .A1(wr_dat[13]), .Z(sw_wdat[13]));
Q_AN02 U476 ( .A0(n389), .A1(wr_dat[14]), .Z(sw_wdat[14]));
Q_AN02 U477 ( .A0(n389), .A1(wr_dat[15]), .Z(sw_wdat[15]));
Q_AN02 U478 ( .A0(n389), .A1(wr_dat[16]), .Z(sw_wdat[16]));
Q_AN02 U479 ( .A0(n389), .A1(wr_dat[17]), .Z(sw_wdat[17]));
Q_AN02 U480 ( .A0(n389), .A1(wr_dat[18]), .Z(sw_wdat[18]));
Q_AN02 U481 ( .A0(n389), .A1(wr_dat[19]), .Z(sw_wdat[19]));
Q_AN02 U482 ( .A0(n389), .A1(wr_dat[20]), .Z(sw_wdat[20]));
Q_AN02 U483 ( .A0(n389), .A1(wr_dat[21]), .Z(sw_wdat[21]));
Q_AN02 U484 ( .A0(n389), .A1(wr_dat[22]), .Z(sw_wdat[22]));
Q_AN02 U485 ( .A0(n389), .A1(wr_dat[23]), .Z(sw_wdat[23]));
Q_AN02 U486 ( .A0(n389), .A1(wr_dat[24]), .Z(sw_wdat[24]));
Q_AN02 U487 ( .A0(n389), .A1(wr_dat[25]), .Z(sw_wdat[25]));
Q_AN02 U488 ( .A0(n389), .A1(wr_dat[26]), .Z(sw_wdat[26]));
Q_AN02 U489 ( .A0(n389), .A1(wr_dat[27]), .Z(sw_wdat[27]));
Q_AN02 U490 ( .A0(n389), .A1(wr_dat[28]), .Z(sw_wdat[28]));
Q_AN02 U491 ( .A0(n389), .A1(wr_dat[29]), .Z(sw_wdat[29]));
Q_AN02 U492 ( .A0(n389), .A1(wr_dat[30]), .Z(sw_wdat[30]));
Q_AN02 U493 ( .A0(n389), .A1(wr_dat[31]), .Z(sw_wdat[31]));
Q_AN02 U494 ( .A0(n389), .A1(wr_dat[32]), .Z(sw_wdat[32]));
Q_AN02 U495 ( .A0(n389), .A1(wr_dat[33]), .Z(sw_wdat[33]));
Q_AN02 U496 ( .A0(n389), .A1(wr_dat[34]), .Z(sw_wdat[34]));
Q_AN02 U497 ( .A0(n389), .A1(wr_dat[35]), .Z(sw_wdat[35]));
Q_AN02 U498 ( .A0(n389), .A1(wr_dat[36]), .Z(sw_wdat[36]));
Q_AN02 U499 ( .A0(n389), .A1(wr_dat[37]), .Z(sw_wdat[37]));
Q_AN02 U500 ( .A0(n389), .A1(wr_dat[38]), .Z(sw_wdat[38]));
Q_AN02 U501 ( .A0(n389), .A1(wr_dat[39]), .Z(sw_wdat[39]));
Q_AN02 U502 ( .A0(n389), .A1(wr_dat[40]), .Z(sw_wdat[40]));
Q_AN02 U503 ( .A0(n389), .A1(wr_dat[41]), .Z(sw_wdat[41]));
Q_AN02 U504 ( .A0(n389), .A1(wr_dat[42]), .Z(sw_wdat[42]));
Q_AN02 U505 ( .A0(n389), .A1(wr_dat[43]), .Z(sw_wdat[43]));
Q_AN02 U506 ( .A0(n389), .A1(wr_dat[44]), .Z(sw_wdat[44]));
Q_AN02 U507 ( .A0(n389), .A1(wr_dat[45]), .Z(sw_wdat[45]));
Q_AN02 U508 ( .A0(n389), .A1(wr_dat[46]), .Z(sw_wdat[46]));
Q_AN02 U509 ( .A0(n389), .A1(wr_dat[47]), .Z(sw_wdat[47]));
Q_AN02 U510 ( .A0(n389), .A1(wr_dat[48]), .Z(sw_wdat[48]));
Q_AN02 U511 ( .A0(n389), .A1(wr_dat[49]), .Z(sw_wdat[49]));
Q_AN02 U512 ( .A0(n389), .A1(wr_dat[50]), .Z(sw_wdat[50]));
Q_AN02 U513 ( .A0(n389), .A1(wr_dat[51]), .Z(sw_wdat[51]));
Q_AN02 U514 ( .A0(n389), .A1(wr_dat[52]), .Z(sw_wdat[52]));
Q_AN02 U515 ( .A0(n389), .A1(wr_dat[53]), .Z(sw_wdat[53]));
Q_AN02 U516 ( .A0(n389), .A1(wr_dat[54]), .Z(sw_wdat[54]));
Q_AN02 U517 ( .A0(n389), .A1(wr_dat[55]), .Z(sw_wdat[55]));
Q_AN02 U518 ( .A0(n389), .A1(wr_dat[56]), .Z(sw_wdat[56]));
Q_AN02 U519 ( .A0(n389), .A1(wr_dat[57]), .Z(sw_wdat[57]));
Q_AN02 U520 ( .A0(n389), .A1(wr_dat[58]), .Z(sw_wdat[58]));
Q_AN02 U521 ( .A0(n389), .A1(wr_dat[59]), .Z(sw_wdat[59]));
Q_AN02 U522 ( .A0(n389), .A1(wr_dat[60]), .Z(sw_wdat[60]));
Q_AN02 U523 ( .A0(n389), .A1(wr_dat[61]), .Z(sw_wdat[61]));
Q_AN02 U524 ( .A0(n389), .A1(wr_dat[62]), .Z(sw_wdat[62]));
Q_AN02 U525 ( .A0(n389), .A1(wr_dat[63]), .Z(sw_wdat[63]));
Q_FDP4EP sim_tmo_r_REG  ( .CK(clk), .CE(n360), .R(n390), .D(cmnd_tmo_stb), .Q(sim_tmo_r));
Q_INV U527 ( .A(rst_n), .Z(n390));
Q_INV U528 ( .A(sim_tmo_r), .Z(n19));
Q_FDP4EP init_r_REG  ( .CK(clk), .CE(n379), .R(n390), .D(n373), .Q(init_r));
Q_INV U530 ( .A(init_r), .Z(enable));
Q_FDP4EP \stat_code_REG[0] ( .CK(clk), .CE(n348), .R(n390), .D(n226), .Q(stat_code[0]));
Q_FDP4EP \stat_code_REG[1] ( .CK(clk), .CE(n348), .R(n390), .D(n231), .Q(stat_code[1]));
Q_FDP4EP \stat_code_REG[2] ( .CK(clk), .CE(n348), .R(n390), .D(n233), .Q(stat_code[2]));
Q_FDP4EP \rst_addr_r_REG[0] ( .CK(clk), .CE(n382), .R(n390), .D(n93), .Q(rst_addr_r[0]));
Q_FDP4EP \rst_addr_r_REG[1] ( .CK(clk), .CE(n382), .R(n390), .D(n95), .Q(rst_addr_r[1]));
Q_FDP4EP \rst_addr_r_REG[2] ( .CK(clk), .CE(n382), .R(n390), .D(n97), .Q(rst_addr_r[2]));
Q_FDP4EP \rst_addr_r_REG[3] ( .CK(clk), .CE(n382), .R(n390), .D(n99), .Q(rst_addr_r[3]));
Q_FDP4EP \rst_addr_r_REG[4] ( .CK(clk), .CE(n382), .R(n390), .D(n101), .Q(rst_addr_r[4]));
Q_FDP4EP \inc_r_REG[0] ( .CK(clk), .CE(n380), .R(n390), .D(n102), .Q(inc_r[0]));
Q_FDP4EP \rd_dat_REG[0] ( .CK(clk), .CE(n378), .R(n390), .D(n103), .Q(rd_dat[0]));
Q_FDP4EP \rd_dat_REG[1] ( .CK(clk), .CE(n378), .R(n390), .D(n104), .Q(rd_dat[1]));
Q_FDP4EP \rd_dat_REG[2] ( .CK(clk), .CE(n378), .R(n390), .D(n105), .Q(rd_dat[2]));
Q_FDP4EP \rd_dat_REG[3] ( .CK(clk), .CE(n378), .R(n390), .D(n106), .Q(rd_dat[3]));
Q_FDP4EP \rd_dat_REG[4] ( .CK(clk), .CE(n378), .R(n390), .D(n107), .Q(rd_dat[4]));
Q_FDP4EP \rd_dat_REG[5] ( .CK(clk), .CE(n378), .R(n390), .D(n109), .Q(rd_dat[5]));
Q_FDP4EP \rd_dat_REG[6] ( .CK(clk), .CE(n378), .R(n390), .D(n111), .Q(rd_dat[6]));
Q_FDP4EP \rd_dat_REG[7] ( .CK(clk), .CE(n378), .R(n390), .D(n113), .Q(rd_dat[7]));
Q_FDP4EP \rd_dat_REG[8] ( .CK(clk), .CE(n378), .R(n390), .D(n115), .Q(rd_dat[8]));
Q_FDP4EP \rd_dat_REG[9] ( .CK(clk), .CE(n378), .R(n390), .D(n117), .Q(rd_dat[9]));
Q_FDP4EP \rd_dat_REG[10] ( .CK(clk), .CE(n378), .R(n390), .D(n119), .Q(rd_dat[10]));
Q_FDP4EP \rd_dat_REG[11] ( .CK(clk), .CE(n378), .R(n390), .D(n121), .Q(rd_dat[11]));
Q_FDP4EP \rd_dat_REG[12] ( .CK(clk), .CE(n378), .R(n390), .D(n123), .Q(rd_dat[12]));
Q_FDP4EP \rd_dat_REG[13] ( .CK(clk), .CE(n378), .R(n390), .D(n125), .Q(rd_dat[13]));
Q_FDP4EP \rd_dat_REG[14] ( .CK(clk), .CE(n378), .R(n390), .D(n127), .Q(rd_dat[14]));
Q_FDP4EP \rd_dat_REG[15] ( .CK(clk), .CE(n378), .R(n390), .D(n129), .Q(rd_dat[15]));
Q_FDP4EP \rd_dat_REG[16] ( .CK(clk), .CE(n378), .R(n390), .D(n131), .Q(rd_dat[16]));
Q_FDP4EP \rd_dat_REG[17] ( .CK(clk), .CE(n378), .R(n390), .D(n133), .Q(rd_dat[17]));
Q_FDP4EP \rd_dat_REG[18] ( .CK(clk), .CE(n378), .R(n390), .D(n135), .Q(rd_dat[18]));
Q_FDP4EP \rd_dat_REG[19] ( .CK(clk), .CE(n378), .R(n390), .D(n137), .Q(rd_dat[19]));
Q_FDP4EP \rd_dat_REG[20] ( .CK(clk), .CE(n378), .R(n390), .D(n139), .Q(rd_dat[20]));
Q_FDP4EP \rd_dat_REG[21] ( .CK(clk), .CE(n378), .R(n390), .D(n141), .Q(rd_dat[21]));
Q_FDP4EP \rd_dat_REG[22] ( .CK(clk), .CE(n378), .R(n390), .D(n143), .Q(rd_dat[22]));
Q_FDP4EP \rd_dat_REG[23] ( .CK(clk), .CE(n378), .R(n390), .D(n145), .Q(rd_dat[23]));
Q_FDP4EP \rd_dat_REG[24] ( .CK(clk), .CE(n378), .R(n390), .D(n147), .Q(rd_dat[24]));
Q_FDP4EP \rd_dat_REG[25] ( .CK(clk), .CE(n378), .R(n390), .D(n149), .Q(rd_dat[25]));
Q_FDP4EP \rd_dat_REG[26] ( .CK(clk), .CE(n378), .R(n390), .D(n151), .Q(rd_dat[26]));
Q_FDP4EP \rd_dat_REG[27] ( .CK(clk), .CE(n378), .R(n390), .D(n153), .Q(rd_dat[27]));
Q_FDP4EP \rd_dat_REG[28] ( .CK(clk), .CE(n378), .R(n390), .D(n155), .Q(rd_dat[28]));
Q_FDP4EP \rd_dat_REG[29] ( .CK(clk), .CE(n378), .R(n390), .D(n157), .Q(rd_dat[29]));
Q_FDP4EP \rd_dat_REG[30] ( .CK(clk), .CE(n378), .R(n390), .D(n159), .Q(rd_dat[30]));
Q_FDP4EP \rd_dat_REG[31] ( .CK(clk), .CE(n378), .R(n390), .D(n161), .Q(rd_dat[31]));
Q_FDP4EP \rd_dat_REG[32] ( .CK(clk), .CE(n378), .R(n390), .D(n163), .Q(rd_dat[32]));
Q_FDP4EP \rd_dat_REG[33] ( .CK(clk), .CE(n378), .R(n390), .D(n165), .Q(rd_dat[33]));
Q_FDP4EP \rd_dat_REG[34] ( .CK(clk), .CE(n378), .R(n390), .D(n167), .Q(rd_dat[34]));
Q_FDP4EP \rd_dat_REG[35] ( .CK(clk), .CE(n378), .R(n390), .D(n169), .Q(rd_dat[35]));
Q_FDP4EP \rd_dat_REG[36] ( .CK(clk), .CE(n378), .R(n390), .D(n171), .Q(rd_dat[36]));
Q_FDP4EP \rd_dat_REG[37] ( .CK(clk), .CE(n378), .R(n390), .D(n173), .Q(rd_dat[37]));
Q_FDP4EP \rd_dat_REG[38] ( .CK(clk), .CE(n378), .R(n390), .D(n175), .Q(rd_dat[38]));
Q_FDP4EP \rd_dat_REG[39] ( .CK(clk), .CE(n378), .R(n390), .D(n177), .Q(rd_dat[39]));
Q_FDP4EP \rd_dat_REG[40] ( .CK(clk), .CE(n378), .R(n390), .D(n179), .Q(rd_dat[40]));
Q_FDP4EP \rd_dat_REG[41] ( .CK(clk), .CE(n378), .R(n390), .D(n181), .Q(rd_dat[41]));
Q_FDP4EP \rd_dat_REG[42] ( .CK(clk), .CE(n378), .R(n390), .D(n183), .Q(rd_dat[42]));
Q_FDP4EP \rd_dat_REG[43] ( .CK(clk), .CE(n378), .R(n390), .D(n185), .Q(rd_dat[43]));
Q_FDP4EP \rd_dat_REG[44] ( .CK(clk), .CE(n378), .R(n390), .D(n187), .Q(rd_dat[44]));
Q_FDP4EP \rd_dat_REG[45] ( .CK(clk), .CE(n378), .R(n390), .D(n189), .Q(rd_dat[45]));
Q_FDP4EP \rd_dat_REG[46] ( .CK(clk), .CE(n378), .R(n390), .D(n191), .Q(rd_dat[46]));
Q_FDP4EP \rd_dat_REG[47] ( .CK(clk), .CE(n378), .R(n390), .D(n193), .Q(rd_dat[47]));
Q_FDP4EP \rd_dat_REG[48] ( .CK(clk), .CE(n378), .R(n390), .D(n195), .Q(rd_dat[48]));
Q_FDP4EP \rd_dat_REG[49] ( .CK(clk), .CE(n378), .R(n390), .D(n197), .Q(rd_dat[49]));
Q_FDP4EP \rd_dat_REG[50] ( .CK(clk), .CE(n378), .R(n390), .D(n199), .Q(rd_dat[50]));
Q_FDP4EP \rd_dat_REG[51] ( .CK(clk), .CE(n378), .R(n390), .D(n201), .Q(rd_dat[51]));
Q_FDP4EP \rd_dat_REG[52] ( .CK(clk), .CE(n378), .R(n390), .D(n203), .Q(rd_dat[52]));
Q_FDP4EP \rd_dat_REG[53] ( .CK(clk), .CE(n378), .R(n390), .D(n205), .Q(rd_dat[53]));
Q_FDP4EP \rd_dat_REG[54] ( .CK(clk), .CE(n378), .R(n390), .D(n207), .Q(rd_dat[54]));
Q_FDP4EP \rd_dat_REG[55] ( .CK(clk), .CE(n378), .R(n390), .D(n209), .Q(rd_dat[55]));
Q_FDP4EP \rd_dat_REG[56] ( .CK(clk), .CE(n378), .R(n390), .D(n211), .Q(rd_dat[56]));
Q_FDP4EP \rd_dat_REG[57] ( .CK(clk), .CE(n378), .R(n390), .D(n213), .Q(rd_dat[57]));
Q_FDP4EP \rd_dat_REG[58] ( .CK(clk), .CE(n378), .R(n390), .D(n215), .Q(rd_dat[58]));
Q_FDP4EP \rd_dat_REG[59] ( .CK(clk), .CE(n378), .R(n390), .D(n217), .Q(rd_dat[59]));
Q_FDP4EP \rd_dat_REG[60] ( .CK(clk), .CE(n378), .R(n390), .D(n219), .Q(rd_dat[60]));
Q_FDP4EP \rd_dat_REG[61] ( .CK(clk), .CE(n378), .R(n390), .D(n221), .Q(rd_dat[61]));
Q_FDP4EP \rd_dat_REG[62] ( .CK(clk), .CE(n378), .R(n390), .D(n223), .Q(rd_dat[62]));
Q_FDP4EP \rd_dat_REG[63] ( .CK(clk), .CE(n378), .R(n390), .D(n225), .Q(rd_dat[63]));
Q_INV U604 ( .A(n381), .Z(n391));
Q_FDP4EP init_inc_r_REG  ( .CK(clk), .CE(n391), .R(n390), .D(n1), .Q(init_inc_r));
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "addr_limit (2,0) 1 4 0 0 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "1"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_1 "-1 genblk2  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_0 "-1 genblk1  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "genblk2"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "genblk1"
endmodule
