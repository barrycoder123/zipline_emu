architecture module of ixc_dutexcl_s2h_port_sync is
  -- quickturn CVASTRPROP MODULE HDLICE PROP_IXCOM_MOD TRUE

begin
end module;
