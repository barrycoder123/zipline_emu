
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module cr_kme_regs_flops ( clk, i_reset_, i_sw_init, o_spare_config, 
	o_cceip0_out_ia_wdata_part0, o_cceip0_out_ia_wdata_part1, 
	o_cceip0_out_ia_wdata_part2, o_cceip0_out_ia_config, 
	o_cceip0_out_im_config, o_cceip0_out_im_read_done, 
	o_cceip1_out_ia_wdata_part0, o_cceip1_out_ia_wdata_part1, 
	o_cceip1_out_ia_wdata_part2, o_cceip1_out_ia_config, 
	o_cceip1_out_im_config, o_cceip1_out_im_read_done, 
	o_cceip2_out_ia_wdata_part0, o_cceip2_out_ia_wdata_part1, 
	o_cceip2_out_ia_wdata_part2, o_cceip2_out_ia_config, 
	o_cceip2_out_im_config, o_cceip2_out_im_read_done, 
	o_cceip3_out_ia_wdata_part0, o_cceip3_out_ia_wdata_part1, 
	o_cceip3_out_ia_wdata_part2, o_cceip3_out_ia_config, 
	o_cceip3_out_im_config, o_cceip3_out_im_read_done, 
	o_cddip0_out_ia_wdata_part0, o_cddip0_out_ia_wdata_part1, 
	o_cddip0_out_ia_wdata_part2, o_cddip0_out_ia_config, 
	o_cddip0_out_im_config, o_cddip0_out_im_read_done, 
	o_cddip1_out_ia_wdata_part0, o_cddip1_out_ia_wdata_part1, 
	o_cddip1_out_ia_wdata_part2, o_cddip1_out_ia_config, 
	o_cddip1_out_im_config, o_cddip1_out_im_read_done, 
	o_cddip2_out_ia_wdata_part0, o_cddip2_out_ia_wdata_part1, 
	o_cddip2_out_ia_wdata_part2, o_cddip2_out_ia_config, 
	o_cddip2_out_im_config, o_cddip2_out_im_read_done, 
	o_cddip3_out_ia_wdata_part0, o_cddip3_out_ia_wdata_part1, 
	o_cddip3_out_ia_wdata_part2, o_cddip3_out_ia_config, 
	o_cddip3_out_im_config, o_cddip3_out_im_read_done, 
	o_ckv_ia_wdata_part0, o_ckv_ia_wdata_part1, o_ckv_ia_config, 
	o_kim_ia_wdata_part0, o_kim_ia_wdata_part1, o_kim_ia_config, 
	o_label0_config, o_label0_data7, o_label0_data6, o_label0_data5, 
	o_label0_data4, o_label0_data3, o_label0_data2, o_label0_data1, 
	o_label0_data0, o_label1_config, o_label1_data7, o_label1_data6, 
	o_label1_data5, o_label1_data4, o_label1_data3, o_label1_data2, 
	o_label1_data1, o_label1_data0, o_label2_config, o_label2_data7, 
	o_label2_data6, o_label2_data5, o_label2_data4, o_label2_data3, 
	o_label2_data2, o_label2_data1, o_label2_data0, o_label3_config, 
	o_label3_data7, o_label3_data6, o_label3_data5, o_label3_data4, 
	o_label3_data3, o_label3_data2, o_label3_data1, o_label3_data0, 
	o_label4_config, o_label4_data7, o_label4_data6, o_label4_data5, 
	o_label4_data4, o_label4_data3, o_label4_data2, o_label4_data1, 
	o_label4_data0, o_label5_config, o_label5_data7, o_label5_data6, 
	o_label5_data5, o_label5_data4, o_label5_data3, o_label5_data2, 
	o_label5_data1, o_label5_data0, o_label6_config, o_label6_data7, 
	o_label6_data6, o_label6_data5, o_label6_data4, o_label6_data3, 
	o_label6_data2, o_label6_data1, o_label6_data0, o_label7_config, 
	o_label7_data7, o_label7_data6, o_label7_data5, o_label7_data4, 
	o_label7_data3, o_label7_data2, o_label7_data1, o_label7_data0, 
	o_kdf_drbg_ctrl, o_kdf_drbg_seed_0_state_key_31_0, 
	o_kdf_drbg_seed_0_state_key_63_32, o_kdf_drbg_seed_0_state_key_95_64, 
	o_kdf_drbg_seed_0_state_key_127_96, 
	o_kdf_drbg_seed_0_state_key_159_128, 
	o_kdf_drbg_seed_0_state_key_191_160, 
	o_kdf_drbg_seed_0_state_key_223_192, 
	o_kdf_drbg_seed_0_state_key_255_224, 
	o_kdf_drbg_seed_0_state_value_31_0, 
	o_kdf_drbg_seed_0_state_value_63_32, 
	o_kdf_drbg_seed_0_state_value_95_64, 
	o_kdf_drbg_seed_0_state_value_127_96, 
	o_kdf_drbg_seed_0_reseed_interval_0, 
	o_kdf_drbg_seed_0_reseed_interval_1, 
	o_kdf_drbg_seed_1_state_key_31_0, o_kdf_drbg_seed_1_state_key_63_32, 
	o_kdf_drbg_seed_1_state_key_95_64, 
	o_kdf_drbg_seed_1_state_key_127_96, 
	o_kdf_drbg_seed_1_state_key_159_128, 
	o_kdf_drbg_seed_1_state_key_191_160, 
	o_kdf_drbg_seed_1_state_key_223_192, 
	o_kdf_drbg_seed_1_state_key_255_224, 
	o_kdf_drbg_seed_1_state_value_31_0, 
	o_kdf_drbg_seed_1_state_value_63_32, 
	o_kdf_drbg_seed_1_state_value_95_64, 
	o_kdf_drbg_seed_1_state_value_127_96, 
	o_kdf_drbg_seed_1_reseed_interval_0, 
	o_kdf_drbg_seed_1_reseed_interval_1, o_interrupt_status, 
	o_interrupt_mask, o_engine_sticky_status, o_bimc_monitor_mask, 
	o_bimc_ecc_uncorrectable_error_cnt, o_bimc_ecc_correctable_error_cnt, 
	o_bimc_parity_error_cnt, o_bimc_global_config, o_bimc_eccpar_debug, 
	o_bimc_cmd2, o_bimc_cmd1, o_bimc_cmd0, o_bimc_rxcmd2, o_bimc_rxrsp2, 
	o_bimc_pollrsp2, o_bimc_dbgcmd2, o_im_consumed, o_tready_override, 
	o_regs_sa_ctrl, o_sa_snapshot_ia_wdata_part0, 
	o_sa_snapshot_ia_wdata_part1, o_sa_snapshot_ia_config, 
	o_sa_count_ia_wdata_part0, o_sa_count_ia_wdata_part1, 
	o_sa_count_ia_config, o_cceip_encrypt_kop_fifo_override, 
	o_cceip_validate_kop_fifo_override, 
	o_cddip_decrypt_kop_fifo_override, o_sa_global_ctrl, 
	o_sa_ctrl_ia_wdata_part0, o_sa_ctrl_ia_config, 
	o_kdf_test_key_size_config, w_load_spare_config, 
	w_load_cceip0_out_ia_wdata_part0, w_load_cceip0_out_ia_wdata_part1, 
	w_load_cceip0_out_ia_wdata_part2, w_load_cceip0_out_ia_config, 
	w_load_cceip0_out_im_config, w_load_cceip0_out_im_read_done, 
	w_load_cceip1_out_ia_wdata_part0, w_load_cceip1_out_ia_wdata_part1, 
	w_load_cceip1_out_ia_wdata_part2, w_load_cceip1_out_ia_config, 
	w_load_cceip1_out_im_config, w_load_cceip1_out_im_read_done, 
	w_load_cceip2_out_ia_wdata_part0, w_load_cceip2_out_ia_wdata_part1, 
	w_load_cceip2_out_ia_wdata_part2, w_load_cceip2_out_ia_config, 
	w_load_cceip2_out_im_config, w_load_cceip2_out_im_read_done, 
	w_load_cceip3_out_ia_wdata_part0, w_load_cceip3_out_ia_wdata_part1, 
	w_load_cceip3_out_ia_wdata_part2, w_load_cceip3_out_ia_config, 
	w_load_cceip3_out_im_config, w_load_cceip3_out_im_read_done, 
	w_load_cddip0_out_ia_wdata_part0, w_load_cddip0_out_ia_wdata_part1, 
	w_load_cddip0_out_ia_wdata_part2, w_load_cddip0_out_ia_config, 
	w_load_cddip0_out_im_config, w_load_cddip0_out_im_read_done, 
	w_load_cddip1_out_ia_wdata_part0, w_load_cddip1_out_ia_wdata_part1, 
	w_load_cddip1_out_ia_wdata_part2, w_load_cddip1_out_ia_config, 
	w_load_cddip1_out_im_config, w_load_cddip1_out_im_read_done, 
	w_load_cddip2_out_ia_wdata_part0, w_load_cddip2_out_ia_wdata_part1, 
	w_load_cddip2_out_ia_wdata_part2, w_load_cddip2_out_ia_config, 
	w_load_cddip2_out_im_config, w_load_cddip2_out_im_read_done, 
	w_load_cddip3_out_ia_wdata_part0, w_load_cddip3_out_ia_wdata_part1, 
	w_load_cddip3_out_ia_wdata_part2, w_load_cddip3_out_ia_config, 
	w_load_cddip3_out_im_config, w_load_cddip3_out_im_read_done, 
	w_load_ckv_ia_wdata_part0, w_load_ckv_ia_wdata_part1, 
	w_load_ckv_ia_config, w_load_kim_ia_wdata_part0, 
	w_load_kim_ia_wdata_part1, w_load_kim_ia_config, 
	w_load_label0_config, w_load_label0_data7, w_load_label0_data6, 
	w_load_label0_data5, w_load_label0_data4, w_load_label0_data3, 
	w_load_label0_data2, w_load_label0_data1, w_load_label0_data0, 
	w_load_label1_config, w_load_label1_data7, w_load_label1_data6, 
	w_load_label1_data5, w_load_label1_data4, w_load_label1_data3, 
	w_load_label1_data2, w_load_label1_data1, w_load_label1_data0, 
	w_load_label2_config, w_load_label2_data7, w_load_label2_data6, 
	w_load_label2_data5, w_load_label2_data4, w_load_label2_data3, 
	w_load_label2_data2, w_load_label2_data1, w_load_label2_data0, 
	w_load_label3_config, w_load_label3_data7, w_load_label3_data6, 
	w_load_label3_data5, w_load_label3_data4, w_load_label3_data3, 
	w_load_label3_data2, w_load_label3_data1, w_load_label3_data0, 
	w_load_label4_config, w_load_label4_data7, w_load_label4_data6, 
	w_load_label4_data5, w_load_label4_data4, w_load_label4_data3, 
	w_load_label4_data2, w_load_label4_data1, w_load_label4_data0, 
	w_load_label5_config, w_load_label5_data7, w_load_label5_data6, 
	w_load_label5_data5, w_load_label5_data4, w_load_label5_data3, 
	w_load_label5_data2, w_load_label5_data1, w_load_label5_data0, 
	w_load_label6_config, w_load_label6_data7, w_load_label6_data6, 
	w_load_label6_data5, w_load_label6_data4, w_load_label6_data3, 
	w_load_label6_data2, w_load_label6_data1, w_load_label6_data0, 
	w_load_label7_config, w_load_label7_data7, w_load_label7_data6, 
	w_load_label7_data5, w_load_label7_data4, w_load_label7_data3, 
	w_load_label7_data2, w_load_label7_data1, w_load_label7_data0, 
	w_load_kdf_drbg_ctrl, w_load_kdf_drbg_seed_0_state_key_31_0, 
	w_load_kdf_drbg_seed_0_state_key_63_32, 
	w_load_kdf_drbg_seed_0_state_key_95_64, 
	w_load_kdf_drbg_seed_0_state_key_127_96, 
	w_load_kdf_drbg_seed_0_state_key_159_128, 
	w_load_kdf_drbg_seed_0_state_key_191_160, 
	w_load_kdf_drbg_seed_0_state_key_223_192, 
	w_load_kdf_drbg_seed_0_state_key_255_224, 
	w_load_kdf_drbg_seed_0_state_value_31_0, 
	w_load_kdf_drbg_seed_0_state_value_63_32, 
	w_load_kdf_drbg_seed_0_state_value_95_64, 
	w_load_kdf_drbg_seed_0_state_value_127_96, 
	w_load_kdf_drbg_seed_0_reseed_interval_0, 
	w_load_kdf_drbg_seed_0_reseed_interval_1, 
	w_load_kdf_drbg_seed_1_state_key_31_0, 
	w_load_kdf_drbg_seed_1_state_key_63_32, 
	w_load_kdf_drbg_seed_1_state_key_95_64, 
	w_load_kdf_drbg_seed_1_state_key_127_96, 
	w_load_kdf_drbg_seed_1_state_key_159_128, 
	w_load_kdf_drbg_seed_1_state_key_191_160, 
	w_load_kdf_drbg_seed_1_state_key_223_192, 
	w_load_kdf_drbg_seed_1_state_key_255_224, 
	w_load_kdf_drbg_seed_1_state_value_31_0, 
	w_load_kdf_drbg_seed_1_state_value_63_32, 
	w_load_kdf_drbg_seed_1_state_value_95_64, 
	w_load_kdf_drbg_seed_1_state_value_127_96, 
	w_load_kdf_drbg_seed_1_reseed_interval_0, 
	w_load_kdf_drbg_seed_1_reseed_interval_1, w_load_interrupt_status, 
	w_load_interrupt_mask, w_load_engine_sticky_status, 
	w_load_bimc_monitor_mask, w_load_bimc_ecc_uncorrectable_error_cnt, 
	w_load_bimc_ecc_correctable_error_cnt, w_load_bimc_parity_error_cnt, 
	w_load_bimc_global_config, w_load_bimc_eccpar_debug, 
	w_load_bimc_cmd2, w_load_bimc_cmd1, w_load_bimc_cmd0, 
	w_load_bimc_rxcmd2, w_load_bimc_rxrsp2, w_load_bimc_pollrsp2, 
	w_load_bimc_dbgcmd2, w_load_im_consumed, w_load_tready_override, 
	w_load_regs_sa_ctrl, w_load_sa_snapshot_ia_wdata_part0, 
	w_load_sa_snapshot_ia_wdata_part1, w_load_sa_snapshot_ia_config, 
	w_load_sa_count_ia_wdata_part0, w_load_sa_count_ia_wdata_part1, 
	w_load_sa_count_ia_config, w_load_cceip_encrypt_kop_fifo_override, 
	w_load_cceip_validate_kop_fifo_override, 
	w_load_cddip_decrypt_kop_fifo_override, w_load_sa_global_ctrl, 
	w_load_sa_ctrl_ia_wdata_part0, w_load_sa_ctrl_ia_config, 
	w_load_kdf_test_key_size_config, f32_data);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
input clk;
input i_reset_;
input i_sw_init;
output [31:0] o_spare_config;
output [31:0] o_cceip0_out_ia_wdata_part0;
output [31:0] o_cceip0_out_ia_wdata_part1;
output [31:0] o_cceip0_out_ia_wdata_part2;
output [12:0] o_cceip0_out_ia_config;
output [11:0] o_cceip0_out_im_config;
output [1:0] o_cceip0_out_im_read_done;
output [31:0] o_cceip1_out_ia_wdata_part0;
output [31:0] o_cceip1_out_ia_wdata_part1;
output [31:0] o_cceip1_out_ia_wdata_part2;
output [12:0] o_cceip1_out_ia_config;
output [11:0] o_cceip1_out_im_config;
output [1:0] o_cceip1_out_im_read_done;
output [31:0] o_cceip2_out_ia_wdata_part0;
output [31:0] o_cceip2_out_ia_wdata_part1;
output [31:0] o_cceip2_out_ia_wdata_part2;
output [12:0] o_cceip2_out_ia_config;
output [11:0] o_cceip2_out_im_config;
output [1:0] o_cceip2_out_im_read_done;
output [31:0] o_cceip3_out_ia_wdata_part0;
output [31:0] o_cceip3_out_ia_wdata_part1;
output [31:0] o_cceip3_out_ia_wdata_part2;
output [12:0] o_cceip3_out_ia_config;
output [11:0] o_cceip3_out_im_config;
output [1:0] o_cceip3_out_im_read_done;
output [31:0] o_cddip0_out_ia_wdata_part0;
output [31:0] o_cddip0_out_ia_wdata_part1;
output [31:0] o_cddip0_out_ia_wdata_part2;
output [12:0] o_cddip0_out_ia_config;
output [11:0] o_cddip0_out_im_config;
output [1:0] o_cddip0_out_im_read_done;
output [31:0] o_cddip1_out_ia_wdata_part0;
output [31:0] o_cddip1_out_ia_wdata_part1;
output [31:0] o_cddip1_out_ia_wdata_part2;
output [12:0] o_cddip1_out_ia_config;
output [11:0] o_cddip1_out_im_config;
output [1:0] o_cddip1_out_im_read_done;
output [31:0] o_cddip2_out_ia_wdata_part0;
output [31:0] o_cddip2_out_ia_wdata_part1;
output [31:0] o_cddip2_out_ia_wdata_part2;
output [12:0] o_cddip2_out_ia_config;
output [11:0] o_cddip2_out_im_config;
output [1:0] o_cddip2_out_im_read_done;
output [31:0] o_cddip3_out_ia_wdata_part0;
output [31:0] o_cddip3_out_ia_wdata_part1;
output [31:0] o_cddip3_out_ia_wdata_part2;
output [12:0] o_cddip3_out_ia_config;
output [11:0] o_cddip3_out_im_config;
output [1:0] o_cddip3_out_im_read_done;
output [31:0] o_ckv_ia_wdata_part0;
output [31:0] o_ckv_ia_wdata_part1;
output [18:0] o_ckv_ia_config;
output [20:0] o_kim_ia_wdata_part0;
output [16:0] o_kim_ia_wdata_part1;
output [17:0] o_kim_ia_config;
output [15:0] o_label0_config;
output [31:0] o_label0_data7;
output [31:0] o_label0_data6;
output [31:0] o_label0_data5;
output [31:0] o_label0_data4;
output [31:0] o_label0_data3;
output [31:0] o_label0_data2;
output [31:0] o_label0_data1;
output [31:0] o_label0_data0;
output [15:0] o_label1_config;
output [31:0] o_label1_data7;
output [31:0] o_label1_data6;
output [31:0] o_label1_data5;
output [31:0] o_label1_data4;
output [31:0] o_label1_data3;
output [31:0] o_label1_data2;
output [31:0] o_label1_data1;
output [31:0] o_label1_data0;
output [15:0] o_label2_config;
output [31:0] o_label2_data7;
output [31:0] o_label2_data6;
output [31:0] o_label2_data5;
output [31:0] o_label2_data4;
output [31:0] o_label2_data3;
output [31:0] o_label2_data2;
output [31:0] o_label2_data1;
output [31:0] o_label2_data0;
output [15:0] o_label3_config;
output [31:0] o_label3_data7;
output [31:0] o_label3_data6;
output [31:0] o_label3_data5;
output [31:0] o_label3_data4;
output [31:0] o_label3_data3;
output [31:0] o_label3_data2;
output [31:0] o_label3_data1;
output [31:0] o_label3_data0;
output [15:0] o_label4_config;
output [31:0] o_label4_data7;
output [31:0] o_label4_data6;
output [31:0] o_label4_data5;
output [31:0] o_label4_data4;
output [31:0] o_label4_data3;
output [31:0] o_label4_data2;
output [31:0] o_label4_data1;
output [31:0] o_label4_data0;
output [15:0] o_label5_config;
output [31:0] o_label5_data7;
output [31:0] o_label5_data6;
output [31:0] o_label5_data5;
output [31:0] o_label5_data4;
output [31:0] o_label5_data3;
output [31:0] o_label5_data2;
output [31:0] o_label5_data1;
output [31:0] o_label5_data0;
output [15:0] o_label6_config;
output [31:0] o_label6_data7;
output [31:0] o_label6_data6;
output [31:0] o_label6_data5;
output [31:0] o_label6_data4;
output [31:0] o_label6_data3;
output [31:0] o_label6_data2;
output [31:0] o_label6_data1;
output [31:0] o_label6_data0;
output [15:0] o_label7_config;
output [31:0] o_label7_data7;
output [31:0] o_label7_data6;
output [31:0] o_label7_data5;
output [31:0] o_label7_data4;
output [31:0] o_label7_data3;
output [31:0] o_label7_data2;
output [31:0] o_label7_data1;
output [31:0] o_label7_data0;
output [1:0] o_kdf_drbg_ctrl;
output [31:0] o_kdf_drbg_seed_0_state_key_31_0;
output [31:0] o_kdf_drbg_seed_0_state_key_63_32;
output [31:0] o_kdf_drbg_seed_0_state_key_95_64;
output [31:0] o_kdf_drbg_seed_0_state_key_127_96;
output [31:0] o_kdf_drbg_seed_0_state_key_159_128;
output [31:0] o_kdf_drbg_seed_0_state_key_191_160;
output [31:0] o_kdf_drbg_seed_0_state_key_223_192;
output [31:0] o_kdf_drbg_seed_0_state_key_255_224;
output [31:0] o_kdf_drbg_seed_0_state_value_31_0;
output [31:0] o_kdf_drbg_seed_0_state_value_63_32;
output [31:0] o_kdf_drbg_seed_0_state_value_95_64;
output [31:0] o_kdf_drbg_seed_0_state_value_127_96;
output [31:0] o_kdf_drbg_seed_0_reseed_interval_0;
output [15:0] o_kdf_drbg_seed_0_reseed_interval_1;
output [31:0] o_kdf_drbg_seed_1_state_key_31_0;
output [31:0] o_kdf_drbg_seed_1_state_key_63_32;
output [31:0] o_kdf_drbg_seed_1_state_key_95_64;
output [31:0] o_kdf_drbg_seed_1_state_key_127_96;
output [31:0] o_kdf_drbg_seed_1_state_key_159_128;
output [31:0] o_kdf_drbg_seed_1_state_key_191_160;
output [31:0] o_kdf_drbg_seed_1_state_key_223_192;
output [31:0] o_kdf_drbg_seed_1_state_key_255_224;
output [31:0] o_kdf_drbg_seed_1_state_value_31_0;
output [31:0] o_kdf_drbg_seed_1_state_value_63_32;
output [31:0] o_kdf_drbg_seed_1_state_value_95_64;
output [31:0] o_kdf_drbg_seed_1_state_value_127_96;
output [31:0] o_kdf_drbg_seed_1_reseed_interval_0;
output [15:0] o_kdf_drbg_seed_1_reseed_interval_1;
output [4:0] o_interrupt_status;
output [4:0] o_interrupt_mask;
output [7:0] o_engine_sticky_status;
output [6:0] o_bimc_monitor_mask;
output [31:0] o_bimc_ecc_uncorrectable_error_cnt;
output [31:0] o_bimc_ecc_correctable_error_cnt;
output [31:0] o_bimc_parity_error_cnt;
output [31:0] o_bimc_global_config;
output [28:0] o_bimc_eccpar_debug;
output [10:0] o_bimc_cmd2;
output [31:0] o_bimc_cmd1;
output [31:0] o_bimc_cmd0;
output [9:0] o_bimc_rxcmd2;
output [9:0] o_bimc_rxrsp2;
output [9:0] o_bimc_pollrsp2;
output [9:0] o_bimc_dbgcmd2;
output [15:0] o_im_consumed;
output [8:0] o_tready_override;
output [31:0] o_regs_sa_ctrl;
output [31:0] o_sa_snapshot_ia_wdata_part0;
output [31:0] o_sa_snapshot_ia_wdata_part1;
output [8:0] o_sa_snapshot_ia_config;
output [31:0] o_sa_count_ia_wdata_part0;
output [31:0] o_sa_count_ia_wdata_part1;
output [8:0] o_sa_count_ia_config;
output [6:0] o_cceip_encrypt_kop_fifo_override;
output [6:0] o_cceip_validate_kop_fifo_override;
output [6:0] o_cddip_decrypt_kop_fifo_override;
output [31:0] o_sa_global_ctrl;
output [31:0] o_sa_ctrl_ia_wdata_part0;
output [8:0] o_sa_ctrl_ia_config;
output [31:0] o_kdf_test_key_size_config;
input w_load_spare_config;
input w_load_cceip0_out_ia_wdata_part0;
input w_load_cceip0_out_ia_wdata_part1;
input w_load_cceip0_out_ia_wdata_part2;
input w_load_cceip0_out_ia_config;
input w_load_cceip0_out_im_config;
input w_load_cceip0_out_im_read_done;
input w_load_cceip1_out_ia_wdata_part0;
input w_load_cceip1_out_ia_wdata_part1;
input w_load_cceip1_out_ia_wdata_part2;
input w_load_cceip1_out_ia_config;
input w_load_cceip1_out_im_config;
input w_load_cceip1_out_im_read_done;
input w_load_cceip2_out_ia_wdata_part0;
input w_load_cceip2_out_ia_wdata_part1;
input w_load_cceip2_out_ia_wdata_part2;
input w_load_cceip2_out_ia_config;
input w_load_cceip2_out_im_config;
input w_load_cceip2_out_im_read_done;
input w_load_cceip3_out_ia_wdata_part0;
input w_load_cceip3_out_ia_wdata_part1;
input w_load_cceip3_out_ia_wdata_part2;
input w_load_cceip3_out_ia_config;
input w_load_cceip3_out_im_config;
input w_load_cceip3_out_im_read_done;
input w_load_cddip0_out_ia_wdata_part0;
input w_load_cddip0_out_ia_wdata_part1;
input w_load_cddip0_out_ia_wdata_part2;
input w_load_cddip0_out_ia_config;
input w_load_cddip0_out_im_config;
input w_load_cddip0_out_im_read_done;
input w_load_cddip1_out_ia_wdata_part0;
input w_load_cddip1_out_ia_wdata_part1;
input w_load_cddip1_out_ia_wdata_part2;
input w_load_cddip1_out_ia_config;
input w_load_cddip1_out_im_config;
input w_load_cddip1_out_im_read_done;
input w_load_cddip2_out_ia_wdata_part0;
input w_load_cddip2_out_ia_wdata_part1;
input w_load_cddip2_out_ia_wdata_part2;
input w_load_cddip2_out_ia_config;
input w_load_cddip2_out_im_config;
input w_load_cddip2_out_im_read_done;
input w_load_cddip3_out_ia_wdata_part0;
input w_load_cddip3_out_ia_wdata_part1;
input w_load_cddip3_out_ia_wdata_part2;
input w_load_cddip3_out_ia_config;
input w_load_cddip3_out_im_config;
input w_load_cddip3_out_im_read_done;
input w_load_ckv_ia_wdata_part0;
input w_load_ckv_ia_wdata_part1;
input w_load_ckv_ia_config;
input w_load_kim_ia_wdata_part0;
input w_load_kim_ia_wdata_part1;
input w_load_kim_ia_config;
input w_load_label0_config;
input w_load_label0_data7;
input w_load_label0_data6;
input w_load_label0_data5;
input w_load_label0_data4;
input w_load_label0_data3;
input w_load_label0_data2;
input w_load_label0_data1;
input w_load_label0_data0;
input w_load_label1_config;
input w_load_label1_data7;
input w_load_label1_data6;
input w_load_label1_data5;
input w_load_label1_data4;
input w_load_label1_data3;
input w_load_label1_data2;
input w_load_label1_data1;
input w_load_label1_data0;
input w_load_label2_config;
input w_load_label2_data7;
input w_load_label2_data6;
input w_load_label2_data5;
input w_load_label2_data4;
input w_load_label2_data3;
input w_load_label2_data2;
input w_load_label2_data1;
input w_load_label2_data0;
input w_load_label3_config;
input w_load_label3_data7;
input w_load_label3_data6;
input w_load_label3_data5;
input w_load_label3_data4;
input w_load_label3_data3;
input w_load_label3_data2;
input w_load_label3_data1;
input w_load_label3_data0;
input w_load_label4_config;
input w_load_label4_data7;
input w_load_label4_data6;
input w_load_label4_data5;
input w_load_label4_data4;
input w_load_label4_data3;
input w_load_label4_data2;
input w_load_label4_data1;
input w_load_label4_data0;
input w_load_label5_config;
input w_load_label5_data7;
input w_load_label5_data6;
input w_load_label5_data5;
input w_load_label5_data4;
input w_load_label5_data3;
input w_load_label5_data2;
input w_load_label5_data1;
input w_load_label5_data0;
input w_load_label6_config;
input w_load_label6_data7;
input w_load_label6_data6;
input w_load_label6_data5;
input w_load_label6_data4;
input w_load_label6_data3;
input w_load_label6_data2;
input w_load_label6_data1;
input w_load_label6_data0;
input w_load_label7_config;
input w_load_label7_data7;
input w_load_label7_data6;
input w_load_label7_data5;
input w_load_label7_data4;
input w_load_label7_data3;
input w_load_label7_data2;
input w_load_label7_data1;
input w_load_label7_data0;
input w_load_kdf_drbg_ctrl;
input w_load_kdf_drbg_seed_0_state_key_31_0;
input w_load_kdf_drbg_seed_0_state_key_63_32;
input w_load_kdf_drbg_seed_0_state_key_95_64;
input w_load_kdf_drbg_seed_0_state_key_127_96;
input w_load_kdf_drbg_seed_0_state_key_159_128;
input w_load_kdf_drbg_seed_0_state_key_191_160;
input w_load_kdf_drbg_seed_0_state_key_223_192;
input w_load_kdf_drbg_seed_0_state_key_255_224;
input w_load_kdf_drbg_seed_0_state_value_31_0;
input w_load_kdf_drbg_seed_0_state_value_63_32;
input w_load_kdf_drbg_seed_0_state_value_95_64;
input w_load_kdf_drbg_seed_0_state_value_127_96;
input w_load_kdf_drbg_seed_0_reseed_interval_0;
input w_load_kdf_drbg_seed_0_reseed_interval_1;
input w_load_kdf_drbg_seed_1_state_key_31_0;
input w_load_kdf_drbg_seed_1_state_key_63_32;
input w_load_kdf_drbg_seed_1_state_key_95_64;
input w_load_kdf_drbg_seed_1_state_key_127_96;
input w_load_kdf_drbg_seed_1_state_key_159_128;
input w_load_kdf_drbg_seed_1_state_key_191_160;
input w_load_kdf_drbg_seed_1_state_key_223_192;
input w_load_kdf_drbg_seed_1_state_key_255_224;
input w_load_kdf_drbg_seed_1_state_value_31_0;
input w_load_kdf_drbg_seed_1_state_value_63_32;
input w_load_kdf_drbg_seed_1_state_value_95_64;
input w_load_kdf_drbg_seed_1_state_value_127_96;
input w_load_kdf_drbg_seed_1_reseed_interval_0;
input w_load_kdf_drbg_seed_1_reseed_interval_1;
input w_load_interrupt_status;
input w_load_interrupt_mask;
input w_load_engine_sticky_status;
input w_load_bimc_monitor_mask;
input w_load_bimc_ecc_uncorrectable_error_cnt;
input w_load_bimc_ecc_correctable_error_cnt;
input w_load_bimc_parity_error_cnt;
input w_load_bimc_global_config;
input w_load_bimc_eccpar_debug;
input w_load_bimc_cmd2;
input w_load_bimc_cmd1;
input w_load_bimc_cmd0;
input w_load_bimc_rxcmd2;
input w_load_bimc_rxrsp2;
input w_load_bimc_pollrsp2;
input w_load_bimc_dbgcmd2;
input w_load_im_consumed;
input w_load_tready_override;
input w_load_regs_sa_ctrl;
input w_load_sa_snapshot_ia_wdata_part0;
input w_load_sa_snapshot_ia_wdata_part1;
input w_load_sa_snapshot_ia_config;
input w_load_sa_count_ia_wdata_part0;
input w_load_sa_count_ia_wdata_part1;
input w_load_sa_count_ia_config;
input w_load_cceip_encrypt_kop_fifo_override;
input w_load_cceip_validate_kop_fifo_override;
input w_load_cddip_decrypt_kop_fifo_override;
input w_load_sa_global_ctrl;
input w_load_sa_ctrl_ia_wdata_part0;
input w_load_sa_ctrl_ia_config;
input w_load_kdf_test_key_size_config;
input [31:0] f32_data;
wire [0:31] _zy_simnet_o_spare_config_0_w$;
wire [0:31] _zy_simnet_o_cceip0_out_ia_wdata_part0_1_w$;
wire [0:31] _zy_simnet_o_cceip0_out_ia_wdata_part1_2_w$;
wire [0:31] _zy_simnet_o_cceip0_out_ia_wdata_part2_3_w$;
wire [0:12] _zy_simnet_o_cceip0_out_ia_config_4_w$;
wire [0:11] _zy_simnet_o_cceip0_out_im_config_5_w$;
wire [0:1] _zy_simnet_o_cceip0_out_im_read_done_6_w$;
wire [0:31] _zy_simnet_o_cceip1_out_ia_wdata_part0_7_w$;
wire [0:31] _zy_simnet_o_cceip1_out_ia_wdata_part1_8_w$;
wire [0:31] _zy_simnet_o_cceip1_out_ia_wdata_part2_9_w$;
wire [0:12] _zy_simnet_o_cceip1_out_ia_config_10_w$;
wire [0:11] _zy_simnet_o_cceip1_out_im_config_11_w$;
wire [0:1] _zy_simnet_o_cceip1_out_im_read_done_12_w$;
wire [0:31] _zy_simnet_o_cceip2_out_ia_wdata_part0_13_w$;
wire [0:31] _zy_simnet_o_cceip2_out_ia_wdata_part1_14_w$;
wire [0:31] _zy_simnet_o_cceip2_out_ia_wdata_part2_15_w$;
wire [0:12] _zy_simnet_o_cceip2_out_ia_config_16_w$;
wire [0:11] _zy_simnet_o_cceip2_out_im_config_17_w$;
wire [0:1] _zy_simnet_o_cceip2_out_im_read_done_18_w$;
wire [0:31] _zy_simnet_o_cceip3_out_ia_wdata_part0_19_w$;
wire [0:31] _zy_simnet_o_cceip3_out_ia_wdata_part1_20_w$;
wire [0:31] _zy_simnet_o_cceip3_out_ia_wdata_part2_21_w$;
wire [0:12] _zy_simnet_o_cceip3_out_ia_config_22_w$;
wire [0:11] _zy_simnet_o_cceip3_out_im_config_23_w$;
wire [0:1] _zy_simnet_o_cceip3_out_im_read_done_24_w$;
wire [0:31] _zy_simnet_o_cddip0_out_ia_wdata_part0_25_w$;
wire [0:31] _zy_simnet_o_cddip0_out_ia_wdata_part1_26_w$;
wire [0:31] _zy_simnet_o_cddip0_out_ia_wdata_part2_27_w$;
wire [0:12] _zy_simnet_o_cddip0_out_ia_config_28_w$;
wire [0:11] _zy_simnet_o_cddip0_out_im_config_29_w$;
wire [0:1] _zy_simnet_o_cddip0_out_im_read_done_30_w$;
wire [0:31] _zy_simnet_o_cddip1_out_ia_wdata_part0_31_w$;
wire [0:31] _zy_simnet_o_cddip1_out_ia_wdata_part1_32_w$;
wire [0:31] _zy_simnet_o_cddip1_out_ia_wdata_part2_33_w$;
wire [0:12] _zy_simnet_o_cddip1_out_ia_config_34_w$;
wire [0:11] _zy_simnet_o_cddip1_out_im_config_35_w$;
wire [0:1] _zy_simnet_o_cddip1_out_im_read_done_36_w$;
wire [0:31] _zy_simnet_o_cddip2_out_ia_wdata_part0_37_w$;
wire [0:31] _zy_simnet_o_cddip2_out_ia_wdata_part1_38_w$;
wire [0:31] _zy_simnet_o_cddip2_out_ia_wdata_part2_39_w$;
wire [0:12] _zy_simnet_o_cddip2_out_ia_config_40_w$;
wire [0:11] _zy_simnet_o_cddip2_out_im_config_41_w$;
wire [0:1] _zy_simnet_o_cddip2_out_im_read_done_42_w$;
wire [0:31] _zy_simnet_o_cddip3_out_ia_wdata_part0_43_w$;
wire [0:31] _zy_simnet_o_cddip3_out_ia_wdata_part1_44_w$;
wire [0:31] _zy_simnet_o_cddip3_out_ia_wdata_part2_45_w$;
wire [0:12] _zy_simnet_o_cddip3_out_ia_config_46_w$;
wire [0:11] _zy_simnet_o_cddip3_out_im_config_47_w$;
wire [0:1] _zy_simnet_o_cddip3_out_im_read_done_48_w$;
wire [0:31] _zy_simnet_o_ckv_ia_wdata_part0_49_w$;
wire [0:31] _zy_simnet_o_ckv_ia_wdata_part1_50_w$;
wire [0:18] _zy_simnet_o_ckv_ia_config_51_w$;
wire [0:20] _zy_simnet_o_kim_ia_wdata_part0_52_w$;
wire [0:16] _zy_simnet_o_kim_ia_wdata_part1_53_w$;
wire [0:17] _zy_simnet_o_kim_ia_config_54_w$;
wire [0:15] _zy_simnet_o_label0_config_55_w$;
wire [0:31] _zy_simnet_o_label0_data7_56_w$;
wire [0:31] _zy_simnet_o_label0_data6_57_w$;
wire [0:31] _zy_simnet_o_label0_data5_58_w$;
wire [0:31] _zy_simnet_o_label0_data4_59_w$;
wire [0:31] _zy_simnet_o_label0_data3_60_w$;
wire [0:31] _zy_simnet_o_label0_data2_61_w$;
wire [0:31] _zy_simnet_o_label0_data1_62_w$;
wire [0:31] _zy_simnet_o_label0_data0_63_w$;
wire [0:15] _zy_simnet_o_label1_config_64_w$;
wire [0:31] _zy_simnet_o_label1_data7_65_w$;
wire [0:31] _zy_simnet_o_label1_data6_66_w$;
wire [0:31] _zy_simnet_o_label1_data5_67_w$;
wire [0:31] _zy_simnet_o_label1_data4_68_w$;
wire [0:31] _zy_simnet_o_label1_data3_69_w$;
wire [0:31] _zy_simnet_o_label1_data2_70_w$;
wire [0:31] _zy_simnet_o_label1_data1_71_w$;
wire [0:31] _zy_simnet_o_label1_data0_72_w$;
wire [0:15] _zy_simnet_o_label2_config_73_w$;
wire [0:31] _zy_simnet_o_label2_data7_74_w$;
wire [0:31] _zy_simnet_o_label2_data6_75_w$;
wire [0:31] _zy_simnet_o_label2_data5_76_w$;
wire [0:31] _zy_simnet_o_label2_data4_77_w$;
wire [0:31] _zy_simnet_o_label2_data3_78_w$;
wire [0:31] _zy_simnet_o_label2_data2_79_w$;
wire [0:31] _zy_simnet_o_label2_data1_80_w$;
wire [0:31] _zy_simnet_o_label2_data0_81_w$;
wire [0:15] _zy_simnet_o_label3_config_82_w$;
wire [0:31] _zy_simnet_o_label3_data7_83_w$;
wire [0:31] _zy_simnet_o_label3_data6_84_w$;
wire [0:31] _zy_simnet_o_label3_data5_85_w$;
wire [0:31] _zy_simnet_o_label3_data4_86_w$;
wire [0:31] _zy_simnet_o_label3_data3_87_w$;
wire [0:31] _zy_simnet_o_label3_data2_88_w$;
wire [0:31] _zy_simnet_o_label3_data1_89_w$;
wire [0:31] _zy_simnet_o_label3_data0_90_w$;
wire [0:15] _zy_simnet_o_label4_config_91_w$;
wire [0:31] _zy_simnet_o_label4_data7_92_w$;
wire [0:31] _zy_simnet_o_label4_data6_93_w$;
wire [0:31] _zy_simnet_o_label4_data5_94_w$;
wire [0:31] _zy_simnet_o_label4_data4_95_w$;
wire [0:31] _zy_simnet_o_label4_data3_96_w$;
wire [0:31] _zy_simnet_o_label4_data2_97_w$;
wire [0:31] _zy_simnet_o_label4_data1_98_w$;
wire [0:31] _zy_simnet_o_label4_data0_99_w$;
wire [0:15] _zy_simnet_o_label5_config_100_w$;
wire [0:31] _zy_simnet_o_label5_data7_101_w$;
wire [0:31] _zy_simnet_o_label5_data6_102_w$;
wire [0:31] _zy_simnet_o_label5_data5_103_w$;
wire [0:31] _zy_simnet_o_label5_data4_104_w$;
wire [0:31] _zy_simnet_o_label5_data3_105_w$;
wire [0:31] _zy_simnet_o_label5_data2_106_w$;
wire [0:31] _zy_simnet_o_label5_data1_107_w$;
wire [0:31] _zy_simnet_o_label5_data0_108_w$;
wire [0:15] _zy_simnet_o_label6_config_109_w$;
wire [0:31] _zy_simnet_o_label6_data7_110_w$;
wire [0:31] _zy_simnet_o_label6_data6_111_w$;
wire [0:31] _zy_simnet_o_label6_data5_112_w$;
wire [0:31] _zy_simnet_o_label6_data4_113_w$;
wire [0:31] _zy_simnet_o_label6_data3_114_w$;
wire [0:31] _zy_simnet_o_label6_data2_115_w$;
wire [0:31] _zy_simnet_o_label6_data1_116_w$;
wire [0:31] _zy_simnet_o_label6_data0_117_w$;
wire [0:15] _zy_simnet_o_label7_config_118_w$;
wire [0:31] _zy_simnet_o_label7_data7_119_w$;
wire [0:31] _zy_simnet_o_label7_data6_120_w$;
wire [0:31] _zy_simnet_o_label7_data5_121_w$;
wire [0:31] _zy_simnet_o_label7_data4_122_w$;
wire [0:31] _zy_simnet_o_label7_data3_123_w$;
wire [0:31] _zy_simnet_o_label7_data2_124_w$;
wire [0:31] _zy_simnet_o_label7_data1_125_w$;
wire [0:31] _zy_simnet_o_label7_data0_126_w$;
wire [0:1] _zy_simnet_o_kdf_drbg_ctrl_127_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_key_31_0_128_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_key_63_32_129_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_key_95_64_130_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_key_127_96_131_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_key_159_128_132_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_key_191_160_133_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_key_223_192_134_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_key_255_224_135_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_value_31_0_136_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_value_63_32_137_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_value_95_64_138_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_value_127_96_139_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_reseed_interval_0_140_w$;
wire [0:15] _zy_simnet_o_kdf_drbg_seed_0_reseed_interval_1_141_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_key_31_0_142_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_key_63_32_143_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_key_95_64_144_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_key_127_96_145_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_key_159_128_146_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_key_191_160_147_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_key_223_192_148_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_key_255_224_149_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_value_31_0_150_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_value_63_32_151_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_value_95_64_152_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_value_127_96_153_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_reseed_interval_0_154_w$;
wire [0:15] _zy_simnet_o_kdf_drbg_seed_1_reseed_interval_1_155_w$;
wire [0:4] _zy_simnet_o_interrupt_status_156_w$;
wire [0:4] _zy_simnet_o_interrupt_mask_157_w$;
wire [0:7] _zy_simnet_o_engine_sticky_status_158_w$;
wire [0:6] _zy_simnet_o_bimc_monitor_mask_159_w$;
wire [0:31] _zy_simnet_o_bimc_ecc_uncorrectable_error_cnt_160_w$;
wire [0:31] _zy_simnet_o_bimc_ecc_correctable_error_cnt_161_w$;
wire [0:31] _zy_simnet_o_bimc_parity_error_cnt_162_w$;
wire [0:31] _zy_simnet_o_bimc_global_config_163_w$;
wire [0:28] _zy_simnet_o_bimc_eccpar_debug_164_w$;
wire [0:10] _zy_simnet_o_bimc_cmd2_165_w$;
wire [0:31] _zy_simnet_o_bimc_cmd1_166_w$;
wire [0:31] _zy_simnet_o_bimc_cmd0_167_w$;
wire [0:9] _zy_simnet_o_bimc_rxcmd2_168_w$;
wire [0:9] _zy_simnet_o_bimc_rxrsp2_169_w$;
wire [0:9] _zy_simnet_o_bimc_pollrsp2_170_w$;
wire [0:9] _zy_simnet_o_bimc_dbgcmd2_171_w$;
wire [0:15] _zy_simnet_o_im_consumed_172_w$;
wire [0:8] _zy_simnet_o_tready_override_173_w$;
wire [0:31] _zy_simnet_o_regs_sa_ctrl_174_w$;
wire [0:31] _zy_simnet_o_sa_snapshot_ia_wdata_part0_175_w$;
wire [0:31] _zy_simnet_o_sa_snapshot_ia_wdata_part1_176_w$;
wire [0:8] _zy_simnet_o_sa_snapshot_ia_config_177_w$;
wire [0:31] _zy_simnet_o_sa_count_ia_wdata_part0_178_w$;
wire [0:31] _zy_simnet_o_sa_count_ia_wdata_part1_179_w$;
wire [0:8] _zy_simnet_o_sa_count_ia_config_180_w$;
wire [0:6] _zy_simnet_o_cceip_encrypt_kop_fifo_override_181_w$;
wire [0:6] _zy_simnet_o_cceip_validate_kop_fifo_override_182_w$;
wire [0:6] _zy_simnet_o_cddip_decrypt_kop_fifo_override_183_w$;
wire [0:31] _zy_simnet_o_sa_global_ctrl_184_w$;
wire [0:31] _zy_simnet_o_sa_ctrl_ia_wdata_part0_185_w$;
wire [0:8] _zy_simnet_o_sa_ctrl_ia_config_186_w$;
wire [0:31] _zy_simnet_o_kdf_test_key_size_config_187_w$;
supply0 n260;
ixc_assign_32 _zz_strnp_187 ( 
	_zy_simnet_o_kdf_test_key_size_config_187_w$[0:31], 
	o_kdf_test_key_size_config[31:0]);
ixc_assign_9 _zz_strnp_186 ( _zy_simnet_o_sa_ctrl_ia_config_186_w$[0:8], 
	o_sa_ctrl_ia_config[8:0]);
ixc_assign_32 _zz_strnp_185 ( _zy_simnet_o_sa_ctrl_ia_wdata_part0_185_w$[0:31], 
	o_sa_ctrl_ia_wdata_part0[31:0]);
ixc_assign_32 _zz_strnp_184 ( _zy_simnet_o_sa_global_ctrl_184_w$[0:31], 
	o_sa_global_ctrl[31:0]);
ixc_assign_7 _zz_strnp_183 ( 
	_zy_simnet_o_cddip_decrypt_kop_fifo_override_183_w$[0:6], 
	o_cddip_decrypt_kop_fifo_override[6:0]);
ixc_assign_7 _zz_strnp_182 ( 
	_zy_simnet_o_cceip_validate_kop_fifo_override_182_w$[0:6], 
	o_cceip_validate_kop_fifo_override[6:0]);
ixc_assign_7 _zz_strnp_181 ( 
	_zy_simnet_o_cceip_encrypt_kop_fifo_override_181_w$[0:6], 
	o_cceip_encrypt_kop_fifo_override[6:0]);
ixc_assign_9 _zz_strnp_180 ( _zy_simnet_o_sa_count_ia_config_180_w$[0:8], 
	o_sa_count_ia_config[8:0]);
ixc_assign_32 _zz_strnp_179 ( 
	_zy_simnet_o_sa_count_ia_wdata_part1_179_w$[0:31], 
	o_sa_count_ia_wdata_part1[31:0]);
ixc_assign_32 _zz_strnp_178 ( 
	_zy_simnet_o_sa_count_ia_wdata_part0_178_w$[0:31], 
	o_sa_count_ia_wdata_part0[31:0]);
ixc_assign_9 _zz_strnp_177 ( _zy_simnet_o_sa_snapshot_ia_config_177_w$[0:8], 
	o_sa_snapshot_ia_config[8:0]);
ixc_assign_32 _zz_strnp_176 ( 
	_zy_simnet_o_sa_snapshot_ia_wdata_part1_176_w$[0:31], 
	o_sa_snapshot_ia_wdata_part1[31:0]);
ixc_assign_32 _zz_strnp_175 ( 
	_zy_simnet_o_sa_snapshot_ia_wdata_part0_175_w$[0:31], 
	o_sa_snapshot_ia_wdata_part0[31:0]);
ixc_assign_32 _zz_strnp_174 ( _zy_simnet_o_regs_sa_ctrl_174_w$[0:31], 
	o_regs_sa_ctrl[31:0]);
ixc_assign_9 _zz_strnp_173 ( _zy_simnet_o_tready_override_173_w$[0:8], 
	o_tready_override[8:0]);
ixc_assign_16 _zz_strnp_172 ( _zy_simnet_o_im_consumed_172_w$[0:15], 
	o_im_consumed[15:0]);
ixc_assign_10 _zz_strnp_171 ( _zy_simnet_o_bimc_dbgcmd2_171_w$[0:9], 
	o_bimc_dbgcmd2[9:0]);
ixc_assign_10 _zz_strnp_170 ( _zy_simnet_o_bimc_pollrsp2_170_w$[0:9], 
	o_bimc_pollrsp2[9:0]);
ixc_assign_10 _zz_strnp_169 ( _zy_simnet_o_bimc_rxrsp2_169_w$[0:9], 
	o_bimc_rxrsp2[9:0]);
ixc_assign_10 _zz_strnp_168 ( _zy_simnet_o_bimc_rxcmd2_168_w$[0:9], 
	o_bimc_rxcmd2[9:0]);
ixc_assign_32 _zz_strnp_167 ( _zy_simnet_o_bimc_cmd0_167_w$[0:31], 
	o_bimc_cmd0[31:0]);
ixc_assign_32 _zz_strnp_166 ( _zy_simnet_o_bimc_cmd1_166_w$[0:31], 
	o_bimc_cmd1[31:0]);
ixc_assign_11 _zz_strnp_165 ( _zy_simnet_o_bimc_cmd2_165_w$[0:10], 
	o_bimc_cmd2[10:0]);
ixc_assign_29 _zz_strnp_164 ( _zy_simnet_o_bimc_eccpar_debug_164_w$[0:28], 
	o_bimc_eccpar_debug[28:0]);
ixc_assign_32 _zz_strnp_163 ( _zy_simnet_o_bimc_global_config_163_w$[0:31], 
	o_bimc_global_config[31:0]);
ixc_assign_32 _zz_strnp_162 ( _zy_simnet_o_bimc_parity_error_cnt_162_w$[0:31], 
	o_bimc_parity_error_cnt[31:0]);
ixc_assign_32 _zz_strnp_161 ( 
	_zy_simnet_o_bimc_ecc_correctable_error_cnt_161_w$[0:31], 
	o_bimc_ecc_correctable_error_cnt[31:0]);
ixc_assign_32 _zz_strnp_160 ( 
	_zy_simnet_o_bimc_ecc_uncorrectable_error_cnt_160_w$[0:31], 
	o_bimc_ecc_uncorrectable_error_cnt[31:0]);
ixc_assign_7 _zz_strnp_159 ( _zy_simnet_o_bimc_monitor_mask_159_w$[0:6], 
	o_bimc_monitor_mask[6:0]);
ixc_assign_8 _zz_strnp_158 ( _zy_simnet_o_engine_sticky_status_158_w$[0:7], 
	o_engine_sticky_status[7:0]);
ixc_assign_5 _zz_strnp_157 ( _zy_simnet_o_interrupt_mask_157_w$[0:4], 
	o_interrupt_mask[4:0]);
ixc_assign_5 _zz_strnp_156 ( _zy_simnet_o_interrupt_status_156_w$[0:4], 
	o_interrupt_status[4:0]);
ixc_assign_16 _zz_strnp_155 ( 
	_zy_simnet_o_kdf_drbg_seed_1_reseed_interval_1_155_w$[0:15], 
	o_kdf_drbg_seed_1_reseed_interval_1[15:0]);
ixc_assign_32 _zz_strnp_154 ( 
	_zy_simnet_o_kdf_drbg_seed_1_reseed_interval_0_154_w$[0:31], 
	o_kdf_drbg_seed_1_reseed_interval_0[31:0]);
ixc_assign_32 _zz_strnp_153 ( 
	_zy_simnet_o_kdf_drbg_seed_1_state_value_127_96_153_w$[0:31], 
	o_kdf_drbg_seed_1_state_value_127_96[31:0]);
ixc_assign_32 _zz_strnp_152 ( 
	_zy_simnet_o_kdf_drbg_seed_1_state_value_95_64_152_w$[0:31], 
	o_kdf_drbg_seed_1_state_value_95_64[31:0]);
ixc_assign_32 _zz_strnp_151 ( 
	_zy_simnet_o_kdf_drbg_seed_1_state_value_63_32_151_w$[0:31], 
	o_kdf_drbg_seed_1_state_value_63_32[31:0]);
ixc_assign_32 _zz_strnp_150 ( 
	_zy_simnet_o_kdf_drbg_seed_1_state_value_31_0_150_w$[0:31], 
	o_kdf_drbg_seed_1_state_value_31_0[31:0]);
ixc_assign_32 _zz_strnp_149 ( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_255_224_149_w$[0:31], 
	o_kdf_drbg_seed_1_state_key_255_224[31:0]);
ixc_assign_32 _zz_strnp_148 ( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_223_192_148_w$[0:31], 
	o_kdf_drbg_seed_1_state_key_223_192[31:0]);
ixc_assign_32 _zz_strnp_147 ( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_191_160_147_w$[0:31], 
	o_kdf_drbg_seed_1_state_key_191_160[31:0]);
ixc_assign_32 _zz_strnp_146 ( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_159_128_146_w$[0:31], 
	o_kdf_drbg_seed_1_state_key_159_128[31:0]);
ixc_assign_32 _zz_strnp_145 ( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_127_96_145_w$[0:31], 
	o_kdf_drbg_seed_1_state_key_127_96[31:0]);
ixc_assign_32 _zz_strnp_144 ( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_95_64_144_w$[0:31], 
	o_kdf_drbg_seed_1_state_key_95_64[31:0]);
ixc_assign_32 _zz_strnp_143 ( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_63_32_143_w$[0:31], 
	o_kdf_drbg_seed_1_state_key_63_32[31:0]);
ixc_assign_32 _zz_strnp_142 ( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_31_0_142_w$[0:31], 
	o_kdf_drbg_seed_1_state_key_31_0[31:0]);
ixc_assign_16 _zz_strnp_141 ( 
	_zy_simnet_o_kdf_drbg_seed_0_reseed_interval_1_141_w$[0:15], 
	o_kdf_drbg_seed_0_reseed_interval_1[15:0]);
ixc_assign_32 _zz_strnp_140 ( 
	_zy_simnet_o_kdf_drbg_seed_0_reseed_interval_0_140_w$[0:31], 
	o_kdf_drbg_seed_0_reseed_interval_0[31:0]);
ixc_assign_32 _zz_strnp_139 ( 
	_zy_simnet_o_kdf_drbg_seed_0_state_value_127_96_139_w$[0:31], 
	o_kdf_drbg_seed_0_state_value_127_96[31:0]);
ixc_assign_32 _zz_strnp_138 ( 
	_zy_simnet_o_kdf_drbg_seed_0_state_value_95_64_138_w$[0:31], 
	o_kdf_drbg_seed_0_state_value_95_64[31:0]);
ixc_assign_32 _zz_strnp_137 ( 
	_zy_simnet_o_kdf_drbg_seed_0_state_value_63_32_137_w$[0:31], 
	o_kdf_drbg_seed_0_state_value_63_32[31:0]);
ixc_assign_32 _zz_strnp_136 ( 
	_zy_simnet_o_kdf_drbg_seed_0_state_value_31_0_136_w$[0:31], 
	o_kdf_drbg_seed_0_state_value_31_0[31:0]);
ixc_assign_32 _zz_strnp_135 ( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_255_224_135_w$[0:31], 
	o_kdf_drbg_seed_0_state_key_255_224[31:0]);
ixc_assign_32 _zz_strnp_134 ( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_223_192_134_w$[0:31], 
	o_kdf_drbg_seed_0_state_key_223_192[31:0]);
ixc_assign_32 _zz_strnp_133 ( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_191_160_133_w$[0:31], 
	o_kdf_drbg_seed_0_state_key_191_160[31:0]);
ixc_assign_32 _zz_strnp_132 ( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_159_128_132_w$[0:31], 
	o_kdf_drbg_seed_0_state_key_159_128[31:0]);
ixc_assign_32 _zz_strnp_131 ( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_127_96_131_w$[0:31], 
	o_kdf_drbg_seed_0_state_key_127_96[31:0]);
ixc_assign_32 _zz_strnp_130 ( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_95_64_130_w$[0:31], 
	o_kdf_drbg_seed_0_state_key_95_64[31:0]);
ixc_assign_32 _zz_strnp_129 ( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_63_32_129_w$[0:31], 
	o_kdf_drbg_seed_0_state_key_63_32[31:0]);
ixc_assign_32 _zz_strnp_128 ( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_31_0_128_w$[0:31], 
	o_kdf_drbg_seed_0_state_key_31_0[31:0]);
ixc_assign_2 _zz_strnp_127 ( _zy_simnet_o_kdf_drbg_ctrl_127_w$[0:1], 
	o_kdf_drbg_ctrl[1:0]);
ixc_assign_32 _zz_strnp_126 ( _zy_simnet_o_label7_data0_126_w$[0:31], 
	o_label7_data0[31:0]);
ixc_assign_32 _zz_strnp_125 ( _zy_simnet_o_label7_data1_125_w$[0:31], 
	o_label7_data1[31:0]);
ixc_assign_32 _zz_strnp_124 ( _zy_simnet_o_label7_data2_124_w$[0:31], 
	o_label7_data2[31:0]);
ixc_assign_32 _zz_strnp_123 ( _zy_simnet_o_label7_data3_123_w$[0:31], 
	o_label7_data3[31:0]);
ixc_assign_32 _zz_strnp_122 ( _zy_simnet_o_label7_data4_122_w$[0:31], 
	o_label7_data4[31:0]);
ixc_assign_32 _zz_strnp_121 ( _zy_simnet_o_label7_data5_121_w$[0:31], 
	o_label7_data5[31:0]);
ixc_assign_32 _zz_strnp_120 ( _zy_simnet_o_label7_data6_120_w$[0:31], 
	o_label7_data6[31:0]);
ixc_assign_32 _zz_strnp_119 ( _zy_simnet_o_label7_data7_119_w$[0:31], 
	o_label7_data7[31:0]);
ixc_assign_16 _zz_strnp_118 ( _zy_simnet_o_label7_config_118_w$[0:15], 
	o_label7_config[15:0]);
ixc_assign_32 _zz_strnp_117 ( _zy_simnet_o_label6_data0_117_w$[0:31], 
	o_label6_data0[31:0]);
ixc_assign_32 _zz_strnp_116 ( _zy_simnet_o_label6_data1_116_w$[0:31], 
	o_label6_data1[31:0]);
ixc_assign_32 _zz_strnp_115 ( _zy_simnet_o_label6_data2_115_w$[0:31], 
	o_label6_data2[31:0]);
ixc_assign_32 _zz_strnp_114 ( _zy_simnet_o_label6_data3_114_w$[0:31], 
	o_label6_data3[31:0]);
ixc_assign_32 _zz_strnp_113 ( _zy_simnet_o_label6_data4_113_w$[0:31], 
	o_label6_data4[31:0]);
ixc_assign_32 _zz_strnp_112 ( _zy_simnet_o_label6_data5_112_w$[0:31], 
	o_label6_data5[31:0]);
ixc_assign_32 _zz_strnp_111 ( _zy_simnet_o_label6_data6_111_w$[0:31], 
	o_label6_data6[31:0]);
ixc_assign_32 _zz_strnp_110 ( _zy_simnet_o_label6_data7_110_w$[0:31], 
	o_label6_data7[31:0]);
ixc_assign_16 _zz_strnp_109 ( _zy_simnet_o_label6_config_109_w$[0:15], 
	o_label6_config[15:0]);
ixc_assign_32 _zz_strnp_108 ( _zy_simnet_o_label5_data0_108_w$[0:31], 
	o_label5_data0[31:0]);
ixc_assign_32 _zz_strnp_107 ( _zy_simnet_o_label5_data1_107_w$[0:31], 
	o_label5_data1[31:0]);
ixc_assign_32 _zz_strnp_106 ( _zy_simnet_o_label5_data2_106_w$[0:31], 
	o_label5_data2[31:0]);
ixc_assign_32 _zz_strnp_105 ( _zy_simnet_o_label5_data3_105_w$[0:31], 
	o_label5_data3[31:0]);
ixc_assign_32 _zz_strnp_104 ( _zy_simnet_o_label5_data4_104_w$[0:31], 
	o_label5_data4[31:0]);
ixc_assign_32 _zz_strnp_103 ( _zy_simnet_o_label5_data5_103_w$[0:31], 
	o_label5_data5[31:0]);
ixc_assign_32 _zz_strnp_102 ( _zy_simnet_o_label5_data6_102_w$[0:31], 
	o_label5_data6[31:0]);
ixc_assign_32 _zz_strnp_101 ( _zy_simnet_o_label5_data7_101_w$[0:31], 
	o_label5_data7[31:0]);
ixc_assign_16 _zz_strnp_100 ( _zy_simnet_o_label5_config_100_w$[0:15], 
	o_label5_config[15:0]);
ixc_assign_32 _zz_strnp_99 ( _zy_simnet_o_label4_data0_99_w$[0:31], 
	o_label4_data0[31:0]);
ixc_assign_32 _zz_strnp_98 ( _zy_simnet_o_label4_data1_98_w$[0:31], 
	o_label4_data1[31:0]);
ixc_assign_32 _zz_strnp_97 ( _zy_simnet_o_label4_data2_97_w$[0:31], 
	o_label4_data2[31:0]);
ixc_assign_32 _zz_strnp_96 ( _zy_simnet_o_label4_data3_96_w$[0:31], 
	o_label4_data3[31:0]);
ixc_assign_32 _zz_strnp_95 ( _zy_simnet_o_label4_data4_95_w$[0:31], 
	o_label4_data4[31:0]);
ixc_assign_32 _zz_strnp_94 ( _zy_simnet_o_label4_data5_94_w$[0:31], 
	o_label4_data5[31:0]);
ixc_assign_32 _zz_strnp_93 ( _zy_simnet_o_label4_data6_93_w$[0:31], 
	o_label4_data6[31:0]);
ixc_assign_32 _zz_strnp_92 ( _zy_simnet_o_label4_data7_92_w$[0:31], 
	o_label4_data7[31:0]);
ixc_assign_16 _zz_strnp_91 ( _zy_simnet_o_label4_config_91_w$[0:15], 
	o_label4_config[15:0]);
ixc_assign_32 _zz_strnp_90 ( _zy_simnet_o_label3_data0_90_w$[0:31], 
	o_label3_data0[31:0]);
ixc_assign_32 _zz_strnp_89 ( _zy_simnet_o_label3_data1_89_w$[0:31], 
	o_label3_data1[31:0]);
ixc_assign_32 _zz_strnp_88 ( _zy_simnet_o_label3_data2_88_w$[0:31], 
	o_label3_data2[31:0]);
ixc_assign_32 _zz_strnp_87 ( _zy_simnet_o_label3_data3_87_w$[0:31], 
	o_label3_data3[31:0]);
ixc_assign_32 _zz_strnp_86 ( _zy_simnet_o_label3_data4_86_w$[0:31], 
	o_label3_data4[31:0]);
ixc_assign_32 _zz_strnp_85 ( _zy_simnet_o_label3_data5_85_w$[0:31], 
	o_label3_data5[31:0]);
ixc_assign_32 _zz_strnp_84 ( _zy_simnet_o_label3_data6_84_w$[0:31], 
	o_label3_data6[31:0]);
ixc_assign_32 _zz_strnp_83 ( _zy_simnet_o_label3_data7_83_w$[0:31], 
	o_label3_data7[31:0]);
ixc_assign_16 _zz_strnp_82 ( _zy_simnet_o_label3_config_82_w$[0:15], 
	o_label3_config[15:0]);
ixc_assign_32 _zz_strnp_81 ( _zy_simnet_o_label2_data0_81_w$[0:31], 
	o_label2_data0[31:0]);
ixc_assign_32 _zz_strnp_80 ( _zy_simnet_o_label2_data1_80_w$[0:31], 
	o_label2_data1[31:0]);
ixc_assign_32 _zz_strnp_79 ( _zy_simnet_o_label2_data2_79_w$[0:31], 
	o_label2_data2[31:0]);
ixc_assign_32 _zz_strnp_78 ( _zy_simnet_o_label2_data3_78_w$[0:31], 
	o_label2_data3[31:0]);
ixc_assign_32 _zz_strnp_77 ( _zy_simnet_o_label2_data4_77_w$[0:31], 
	o_label2_data4[31:0]);
ixc_assign_32 _zz_strnp_76 ( _zy_simnet_o_label2_data5_76_w$[0:31], 
	o_label2_data5[31:0]);
ixc_assign_32 _zz_strnp_75 ( _zy_simnet_o_label2_data6_75_w$[0:31], 
	o_label2_data6[31:0]);
ixc_assign_32 _zz_strnp_74 ( _zy_simnet_o_label2_data7_74_w$[0:31], 
	o_label2_data7[31:0]);
ixc_assign_16 _zz_strnp_73 ( _zy_simnet_o_label2_config_73_w$[0:15], 
	o_label2_config[15:0]);
ixc_assign_32 _zz_strnp_72 ( _zy_simnet_o_label1_data0_72_w$[0:31], 
	o_label1_data0[31:0]);
ixc_assign_32 _zz_strnp_71 ( _zy_simnet_o_label1_data1_71_w$[0:31], 
	o_label1_data1[31:0]);
ixc_assign_32 _zz_strnp_70 ( _zy_simnet_o_label1_data2_70_w$[0:31], 
	o_label1_data2[31:0]);
ixc_assign_32 _zz_strnp_69 ( _zy_simnet_o_label1_data3_69_w$[0:31], 
	o_label1_data3[31:0]);
ixc_assign_32 _zz_strnp_68 ( _zy_simnet_o_label1_data4_68_w$[0:31], 
	o_label1_data4[31:0]);
ixc_assign_32 _zz_strnp_67 ( _zy_simnet_o_label1_data5_67_w$[0:31], 
	o_label1_data5[31:0]);
ixc_assign_32 _zz_strnp_66 ( _zy_simnet_o_label1_data6_66_w$[0:31], 
	o_label1_data6[31:0]);
ixc_assign_32 _zz_strnp_65 ( _zy_simnet_o_label1_data7_65_w$[0:31], 
	o_label1_data7[31:0]);
ixc_assign_16 _zz_strnp_64 ( _zy_simnet_o_label1_config_64_w$[0:15], 
	o_label1_config[15:0]);
ixc_assign_32 _zz_strnp_63 ( _zy_simnet_o_label0_data0_63_w$[0:31], 
	o_label0_data0[31:0]);
ixc_assign_32 _zz_strnp_62 ( _zy_simnet_o_label0_data1_62_w$[0:31], 
	o_label0_data1[31:0]);
ixc_assign_32 _zz_strnp_61 ( _zy_simnet_o_label0_data2_61_w$[0:31], 
	o_label0_data2[31:0]);
ixc_assign_32 _zz_strnp_60 ( _zy_simnet_o_label0_data3_60_w$[0:31], 
	o_label0_data3[31:0]);
ixc_assign_32 _zz_strnp_59 ( _zy_simnet_o_label0_data4_59_w$[0:31], 
	o_label0_data4[31:0]);
ixc_assign_32 _zz_strnp_58 ( _zy_simnet_o_label0_data5_58_w$[0:31], 
	o_label0_data5[31:0]);
ixc_assign_32 _zz_strnp_57 ( _zy_simnet_o_label0_data6_57_w$[0:31], 
	o_label0_data6[31:0]);
ixc_assign_32 _zz_strnp_56 ( _zy_simnet_o_label0_data7_56_w$[0:31], 
	o_label0_data7[31:0]);
ixc_assign_16 _zz_strnp_55 ( _zy_simnet_o_label0_config_55_w$[0:15], 
	o_label0_config[15:0]);
ixc_assign_18 _zz_strnp_54 ( _zy_simnet_o_kim_ia_config_54_w$[0:17], 
	o_kim_ia_config[17:0]);
ixc_assign_17 _zz_strnp_53 ( _zy_simnet_o_kim_ia_wdata_part1_53_w$[0:16], 
	o_kim_ia_wdata_part1[16:0]);
ixc_assign_21 _zz_strnp_52 ( _zy_simnet_o_kim_ia_wdata_part0_52_w$[0:20], 
	o_kim_ia_wdata_part0[20:0]);
ixc_assign_19 _zz_strnp_51 ( _zy_simnet_o_ckv_ia_config_51_w$[0:18], 
	o_ckv_ia_config[18:0]);
ixc_assign_32 _zz_strnp_50 ( _zy_simnet_o_ckv_ia_wdata_part1_50_w$[0:31], 
	o_ckv_ia_wdata_part1[31:0]);
ixc_assign_32 _zz_strnp_49 ( _zy_simnet_o_ckv_ia_wdata_part0_49_w$[0:31], 
	o_ckv_ia_wdata_part0[31:0]);
ixc_assign_2 _zz_strnp_48 ( _zy_simnet_o_cddip3_out_im_read_done_48_w$[0:1], 
	o_cddip3_out_im_read_done[1:0]);
ixc_assign_12 _zz_strnp_47 ( _zy_simnet_o_cddip3_out_im_config_47_w$[0:11], 
	o_cddip3_out_im_config[11:0]);
ixc_assign_13 _zz_strnp_46 ( _zy_simnet_o_cddip3_out_ia_config_46_w$[0:12], 
	o_cddip3_out_ia_config[12:0]);
ixc_assign_32 _zz_strnp_45 ( 
	_zy_simnet_o_cddip3_out_ia_wdata_part2_45_w$[0:31], 
	o_cddip3_out_ia_wdata_part2[31:0]);
ixc_assign_32 _zz_strnp_44 ( 
	_zy_simnet_o_cddip3_out_ia_wdata_part1_44_w$[0:31], 
	o_cddip3_out_ia_wdata_part1[31:0]);
ixc_assign_32 _zz_strnp_43 ( 
	_zy_simnet_o_cddip3_out_ia_wdata_part0_43_w$[0:31], 
	o_cddip3_out_ia_wdata_part0[31:0]);
ixc_assign_2 _zz_strnp_42 ( _zy_simnet_o_cddip2_out_im_read_done_42_w$[0:1], 
	o_cddip2_out_im_read_done[1:0]);
ixc_assign_12 _zz_strnp_41 ( _zy_simnet_o_cddip2_out_im_config_41_w$[0:11], 
	o_cddip2_out_im_config[11:0]);
ixc_assign_13 _zz_strnp_40 ( _zy_simnet_o_cddip2_out_ia_config_40_w$[0:12], 
	o_cddip2_out_ia_config[12:0]);
ixc_assign_32 _zz_strnp_39 ( 
	_zy_simnet_o_cddip2_out_ia_wdata_part2_39_w$[0:31], 
	o_cddip2_out_ia_wdata_part2[31:0]);
ixc_assign_32 _zz_strnp_38 ( 
	_zy_simnet_o_cddip2_out_ia_wdata_part1_38_w$[0:31], 
	o_cddip2_out_ia_wdata_part1[31:0]);
ixc_assign_32 _zz_strnp_37 ( 
	_zy_simnet_o_cddip2_out_ia_wdata_part0_37_w$[0:31], 
	o_cddip2_out_ia_wdata_part0[31:0]);
ixc_assign_2 _zz_strnp_36 ( _zy_simnet_o_cddip1_out_im_read_done_36_w$[0:1], 
	o_cddip1_out_im_read_done[1:0]);
ixc_assign_12 _zz_strnp_35 ( _zy_simnet_o_cddip1_out_im_config_35_w$[0:11], 
	o_cddip1_out_im_config[11:0]);
ixc_assign_13 _zz_strnp_34 ( _zy_simnet_o_cddip1_out_ia_config_34_w$[0:12], 
	o_cddip1_out_ia_config[12:0]);
ixc_assign_32 _zz_strnp_33 ( 
	_zy_simnet_o_cddip1_out_ia_wdata_part2_33_w$[0:31], 
	o_cddip1_out_ia_wdata_part2[31:0]);
ixc_assign_32 _zz_strnp_32 ( 
	_zy_simnet_o_cddip1_out_ia_wdata_part1_32_w$[0:31], 
	o_cddip1_out_ia_wdata_part1[31:0]);
ixc_assign_32 _zz_strnp_31 ( 
	_zy_simnet_o_cddip1_out_ia_wdata_part0_31_w$[0:31], 
	o_cddip1_out_ia_wdata_part0[31:0]);
ixc_assign_2 _zz_strnp_30 ( _zy_simnet_o_cddip0_out_im_read_done_30_w$[0:1], 
	o_cddip0_out_im_read_done[1:0]);
ixc_assign_12 _zz_strnp_29 ( _zy_simnet_o_cddip0_out_im_config_29_w$[0:11], 
	o_cddip0_out_im_config[11:0]);
ixc_assign_13 _zz_strnp_28 ( _zy_simnet_o_cddip0_out_ia_config_28_w$[0:12], 
	o_cddip0_out_ia_config[12:0]);
ixc_assign_32 _zz_strnp_27 ( 
	_zy_simnet_o_cddip0_out_ia_wdata_part2_27_w$[0:31], 
	o_cddip0_out_ia_wdata_part2[31:0]);
ixc_assign_32 _zz_strnp_26 ( 
	_zy_simnet_o_cddip0_out_ia_wdata_part1_26_w$[0:31], 
	o_cddip0_out_ia_wdata_part1[31:0]);
ixc_assign_32 _zz_strnp_25 ( 
	_zy_simnet_o_cddip0_out_ia_wdata_part0_25_w$[0:31], 
	o_cddip0_out_ia_wdata_part0[31:0]);
ixc_assign_2 _zz_strnp_24 ( _zy_simnet_o_cceip3_out_im_read_done_24_w$[0:1], 
	o_cceip3_out_im_read_done[1:0]);
ixc_assign_12 _zz_strnp_23 ( _zy_simnet_o_cceip3_out_im_config_23_w$[0:11], 
	o_cceip3_out_im_config[11:0]);
ixc_assign_13 _zz_strnp_22 ( _zy_simnet_o_cceip3_out_ia_config_22_w$[0:12], 
	o_cceip3_out_ia_config[12:0]);
ixc_assign_32 _zz_strnp_21 ( 
	_zy_simnet_o_cceip3_out_ia_wdata_part2_21_w$[0:31], 
	o_cceip3_out_ia_wdata_part2[31:0]);
ixc_assign_32 _zz_strnp_20 ( 
	_zy_simnet_o_cceip3_out_ia_wdata_part1_20_w$[0:31], 
	o_cceip3_out_ia_wdata_part1[31:0]);
ixc_assign_32 _zz_strnp_19 ( 
	_zy_simnet_o_cceip3_out_ia_wdata_part0_19_w$[0:31], 
	o_cceip3_out_ia_wdata_part0[31:0]);
ixc_assign_2 _zz_strnp_18 ( _zy_simnet_o_cceip2_out_im_read_done_18_w$[0:1], 
	o_cceip2_out_im_read_done[1:0]);
ixc_assign_12 _zz_strnp_17 ( _zy_simnet_o_cceip2_out_im_config_17_w$[0:11], 
	o_cceip2_out_im_config[11:0]);
ixc_assign_13 _zz_strnp_16 ( _zy_simnet_o_cceip2_out_ia_config_16_w$[0:12], 
	o_cceip2_out_ia_config[12:0]);
ixc_assign_32 _zz_strnp_15 ( 
	_zy_simnet_o_cceip2_out_ia_wdata_part2_15_w$[0:31], 
	o_cceip2_out_ia_wdata_part2[31:0]);
ixc_assign_32 _zz_strnp_14 ( 
	_zy_simnet_o_cceip2_out_ia_wdata_part1_14_w$[0:31], 
	o_cceip2_out_ia_wdata_part1[31:0]);
ixc_assign_32 _zz_strnp_13 ( 
	_zy_simnet_o_cceip2_out_ia_wdata_part0_13_w$[0:31], 
	o_cceip2_out_ia_wdata_part0[31:0]);
ixc_assign_2 _zz_strnp_12 ( _zy_simnet_o_cceip1_out_im_read_done_12_w$[0:1], 
	o_cceip1_out_im_read_done[1:0]);
ixc_assign_12 _zz_strnp_11 ( _zy_simnet_o_cceip1_out_im_config_11_w$[0:11], 
	o_cceip1_out_im_config[11:0]);
ixc_assign_13 _zz_strnp_10 ( _zy_simnet_o_cceip1_out_ia_config_10_w$[0:12], 
	o_cceip1_out_ia_config[12:0]);
ixc_assign_32 _zz_strnp_9 ( _zy_simnet_o_cceip1_out_ia_wdata_part2_9_w$[0:31], 
	o_cceip1_out_ia_wdata_part2[31:0]);
ixc_assign_32 _zz_strnp_8 ( _zy_simnet_o_cceip1_out_ia_wdata_part1_8_w$[0:31], 
	o_cceip1_out_ia_wdata_part1[31:0]);
ixc_assign_32 _zz_strnp_7 ( _zy_simnet_o_cceip1_out_ia_wdata_part0_7_w$[0:31], 
	o_cceip1_out_ia_wdata_part0[31:0]);
ixc_assign_2 _zz_strnp_6 ( _zy_simnet_o_cceip0_out_im_read_done_6_w$[0:1], 
	o_cceip0_out_im_read_done[1:0]);
ixc_assign_12 _zz_strnp_5 ( _zy_simnet_o_cceip0_out_im_config_5_w$[0:11], 
	o_cceip0_out_im_config[11:0]);
ixc_assign_13 _zz_strnp_4 ( _zy_simnet_o_cceip0_out_ia_config_4_w$[0:12], 
	o_cceip0_out_ia_config[12:0]);
ixc_assign_32 _zz_strnp_3 ( _zy_simnet_o_cceip0_out_ia_wdata_part2_3_w$[0:31], 
	o_cceip0_out_ia_wdata_part2[31:0]);
ixc_assign_32 _zz_strnp_2 ( _zy_simnet_o_cceip0_out_ia_wdata_part1_2_w$[0:31], 
	o_cceip0_out_ia_wdata_part1[31:0]);
ixc_assign_32 _zz_strnp_1 ( _zy_simnet_o_cceip0_out_ia_wdata_part0_1_w$[0:31], 
	o_cceip0_out_ia_wdata_part0[31:0]);
ixc_assign_32 _zz_strnp_0 ( _zy_simnet_o_spare_config_0_w$[0:31], 
	o_spare_config[31:0]);
Q_OR02 U188 ( .A0(i_sw_init), .A1(f32_data[0]), .Z(n1));
Q_OR02 U189 ( .A0(i_sw_init), .A1(f32_data[8]), .Z(n2));
Q_OR02 U190 ( .A0(i_sw_init), .A1(f32_data[9]), .Z(n3));
Q_OR02 U191 ( .A0(i_sw_init), .A1(f32_data[30]), .Z(n4));
Q_OR02 U192 ( .A0(i_sw_init), .A1(f32_data[31]), .Z(n5));
Q_AN02 U193 ( .A0(n71), .A1(f32_data[0]), .Z(n6));
Q_AN02 U194 ( .A0(n71), .A1(f32_data[1]), .Z(n7));
Q_AN02 U195 ( .A0(n71), .A1(f32_data[2]), .Z(n8));
Q_AN02 U196 ( .A0(n71), .A1(f32_data[3]), .Z(n9));
Q_AN02 U197 ( .A0(n71), .A1(f32_data[4]), .Z(n10));
Q_AN02 U198 ( .A0(n71), .A1(f32_data[5]), .Z(n11));
Q_AN02 U199 ( .A0(n71), .A1(f32_data[6]), .Z(n12));
Q_AN02 U200 ( .A0(n71), .A1(f32_data[7]), .Z(n13));
Q_AN02 U201 ( .A0(n71), .A1(f32_data[8]), .Z(n14));
Q_AN02 U202 ( .A0(n71), .A1(f32_data[9]), .Z(n15));
Q_AN02 U203 ( .A0(n71), .A1(f32_data[10]), .Z(n16));
Q_AN02 U204 ( .A0(n71), .A1(f32_data[11]), .Z(n17));
Q_AN02 U205 ( .A0(n71), .A1(f32_data[12]), .Z(n18));
Q_AN02 U206 ( .A0(n71), .A1(f32_data[13]), .Z(n19));
Q_AN02 U207 ( .A0(n71), .A1(f32_data[14]), .Z(n20));
Q_AN02 U208 ( .A0(n71), .A1(f32_data[15]), .Z(n21));
Q_AN02 U209 ( .A0(n71), .A1(f32_data[16]), .Z(n22));
Q_AN02 U210 ( .A0(n71), .A1(f32_data[17]), .Z(n23));
Q_AN02 U211 ( .A0(n71), .A1(f32_data[18]), .Z(n24));
Q_AN02 U212 ( .A0(n71), .A1(f32_data[19]), .Z(n25));
Q_AN02 U213 ( .A0(n71), .A1(f32_data[20]), .Z(n26));
Q_AN02 U214 ( .A0(n71), .A1(f32_data[21]), .Z(n27));
Q_AN02 U215 ( .A0(n71), .A1(f32_data[22]), .Z(n28));
Q_AN02 U216 ( .A0(n71), .A1(f32_data[23]), .Z(n29));
Q_AN02 U217 ( .A0(n71), .A1(f32_data[24]), .Z(n30));
Q_AN02 U218 ( .A0(n71), .A1(f32_data[25]), .Z(n31));
Q_AN02 U219 ( .A0(n71), .A1(f32_data[26]), .Z(n32));
Q_AN02 U220 ( .A0(n71), .A1(f32_data[27]), .Z(n33));
Q_AN02 U221 ( .A0(n71), .A1(f32_data[28]), .Z(n34));
Q_AN02 U222 ( .A0(n71), .A1(f32_data[29]), .Z(n35));
Q_AN02 U223 ( .A0(n71), .A1(f32_data[30]), .Z(n36));
Q_AN02 U224 ( .A0(n71), .A1(f32_data[31]), .Z(n37));
Q_FDP2 \o_cceip0_out_im_config_REG[11] ( .CK(clk), .S(i_reset_), .D(n38), .Q(o_cceip0_out_im_config[11]), .QN( ));
Q_MX02 U226 ( .S(n77), .A0(o_cceip0_out_im_config[11]), .A1(n5), .Z(n38));
Q_FDP2 \o_cceip0_out_im_config_REG[10] ( .CK(clk), .S(i_reset_), .D(n39), .Q(o_cceip0_out_im_config[10]), .QN( ));
Q_MX02 U228 ( .S(n77), .A0(o_cceip0_out_im_config[10]), .A1(n4), .Z(n39));
Q_FDP2 \o_cceip0_out_im_config_REG[9] ( .CK(clk), .S(i_reset_), .D(n40), .Q(o_cceip0_out_im_config[9]), .QN( ));
Q_MX02 U230 ( .S(n77), .A0(o_cceip0_out_im_config[9]), .A1(n3), .Z(n40));
Q_FDP2 \o_cceip1_out_im_config_REG[11] ( .CK(clk), .S(i_reset_), .D(n41), .Q(o_cceip1_out_im_config[11]), .QN( ));
Q_MX02 U232 ( .S(n83), .A0(o_cceip1_out_im_config[11]), .A1(n5), .Z(n41));
Q_FDP2 \o_cceip1_out_im_config_REG[10] ( .CK(clk), .S(i_reset_), .D(n42), .Q(o_cceip1_out_im_config[10]), .QN( ));
Q_MX02 U234 ( .S(n83), .A0(o_cceip1_out_im_config[10]), .A1(n4), .Z(n42));
Q_FDP2 \o_cceip1_out_im_config_REG[9] ( .CK(clk), .S(i_reset_), .D(n43), .Q(o_cceip1_out_im_config[9]), .QN( ));
Q_MX02 U236 ( .S(n83), .A0(o_cceip1_out_im_config[9]), .A1(n3), .Z(n43));
Q_FDP2 \o_cceip2_out_im_config_REG[11] ( .CK(clk), .S(i_reset_), .D(n44), .Q(o_cceip2_out_im_config[11]), .QN( ));
Q_MX02 U238 ( .S(n89), .A0(o_cceip2_out_im_config[11]), .A1(n5), .Z(n44));
Q_FDP2 \o_cceip2_out_im_config_REG[10] ( .CK(clk), .S(i_reset_), .D(n45), .Q(o_cceip2_out_im_config[10]), .QN( ));
Q_MX02 U240 ( .S(n89), .A0(o_cceip2_out_im_config[10]), .A1(n4), .Z(n45));
Q_FDP2 \o_cceip2_out_im_config_REG[9] ( .CK(clk), .S(i_reset_), .D(n46), .Q(o_cceip2_out_im_config[9]), .QN( ));
Q_MX02 U242 ( .S(n89), .A0(o_cceip2_out_im_config[9]), .A1(n3), .Z(n46));
Q_FDP2 \o_cceip3_out_im_config_REG[11] ( .CK(clk), .S(i_reset_), .D(n47), .Q(o_cceip3_out_im_config[11]), .QN( ));
Q_MX02 U244 ( .S(n95), .A0(o_cceip3_out_im_config[11]), .A1(n5), .Z(n47));
Q_FDP2 \o_cceip3_out_im_config_REG[10] ( .CK(clk), .S(i_reset_), .D(n48), .Q(o_cceip3_out_im_config[10]), .QN( ));
Q_MX02 U246 ( .S(n95), .A0(o_cceip3_out_im_config[10]), .A1(n4), .Z(n48));
Q_FDP2 \o_cceip3_out_im_config_REG[9] ( .CK(clk), .S(i_reset_), .D(n49), .Q(o_cceip3_out_im_config[9]), .QN( ));
Q_MX02 U248 ( .S(n95), .A0(o_cceip3_out_im_config[9]), .A1(n3), .Z(n49));
Q_FDP2 \o_cddip0_out_im_config_REG[11] ( .CK(clk), .S(i_reset_), .D(n50), .Q(o_cddip0_out_im_config[11]), .QN( ));
Q_MX02 U250 ( .S(n101), .A0(o_cddip0_out_im_config[11]), .A1(n5), .Z(n50));
Q_FDP2 \o_cddip0_out_im_config_REG[10] ( .CK(clk), .S(i_reset_), .D(n51), .Q(o_cddip0_out_im_config[10]), .QN( ));
Q_MX02 U252 ( .S(n101), .A0(o_cddip0_out_im_config[10]), .A1(n4), .Z(n51));
Q_FDP2 \o_cddip0_out_im_config_REG[9] ( .CK(clk), .S(i_reset_), .D(n52), .Q(o_cddip0_out_im_config[9]), .QN( ));
Q_MX02 U254 ( .S(n101), .A0(o_cddip0_out_im_config[9]), .A1(n3), .Z(n52));
Q_FDP2 \o_cddip1_out_im_config_REG[11] ( .CK(clk), .S(i_reset_), .D(n53), .Q(o_cddip1_out_im_config[11]), .QN( ));
Q_MX02 U256 ( .S(n107), .A0(o_cddip1_out_im_config[11]), .A1(n5), .Z(n53));
Q_FDP2 \o_cddip1_out_im_config_REG[10] ( .CK(clk), .S(i_reset_), .D(n54), .Q(o_cddip1_out_im_config[10]), .QN( ));
Q_MX02 U258 ( .S(n107), .A0(o_cddip1_out_im_config[10]), .A1(n4), .Z(n54));
Q_FDP2 \o_cddip1_out_im_config_REG[9] ( .CK(clk), .S(i_reset_), .D(n55), .Q(o_cddip1_out_im_config[9]), .QN( ));
Q_MX02 U260 ( .S(n107), .A0(o_cddip1_out_im_config[9]), .A1(n3), .Z(n55));
Q_FDP2 \o_cddip2_out_im_config_REG[11] ( .CK(clk), .S(i_reset_), .D(n56), .Q(o_cddip2_out_im_config[11]), .QN( ));
Q_MX02 U262 ( .S(n113), .A0(o_cddip2_out_im_config[11]), .A1(n5), .Z(n56));
Q_FDP2 \o_cddip2_out_im_config_REG[10] ( .CK(clk), .S(i_reset_), .D(n57), .Q(o_cddip2_out_im_config[10]), .QN( ));
Q_MX02 U264 ( .S(n113), .A0(o_cddip2_out_im_config[10]), .A1(n4), .Z(n57));
Q_FDP2 \o_cddip2_out_im_config_REG[9] ( .CK(clk), .S(i_reset_), .D(n58), .Q(o_cddip2_out_im_config[9]), .QN( ));
Q_MX02 U266 ( .S(n113), .A0(o_cddip2_out_im_config[9]), .A1(n3), .Z(n58));
Q_FDP2 \o_cddip3_out_im_config_REG[11] ( .CK(clk), .S(i_reset_), .D(n59), .Q(o_cddip3_out_im_config[11]), .QN( ));
Q_MX02 U268 ( .S(n119), .A0(o_cddip3_out_im_config[11]), .A1(n5), .Z(n59));
Q_FDP2 \o_cddip3_out_im_config_REG[10] ( .CK(clk), .S(i_reset_), .D(n60), .Q(o_cddip3_out_im_config[10]), .QN( ));
Q_MX02 U270 ( .S(n119), .A0(o_cddip3_out_im_config[10]), .A1(n4), .Z(n60));
Q_FDP2 \o_cddip3_out_im_config_REG[9] ( .CK(clk), .S(i_reset_), .D(n61), .Q(o_cddip3_out_im_config[9]), .QN( ));
Q_MX02 U272 ( .S(n119), .A0(o_cddip3_out_im_config[9]), .A1(n3), .Z(n61));
Q_FDP2 \o_label0_config_REG[8] ( .CK(clk), .S(i_reset_), .D(n62), .Q(o_label0_config[8]), .QN( ));
Q_MX02 U274 ( .S(n127), .A0(o_label0_config[8]), .A1(n2), .Z(n62));
Q_FDP2 \o_label1_config_REG[8] ( .CK(clk), .S(i_reset_), .D(n63), .Q(o_label1_config[8]), .QN( ));
Q_MX02 U276 ( .S(n136), .A0(o_label1_config[8]), .A1(n2), .Z(n63));
Q_FDP2 \o_label2_config_REG[8] ( .CK(clk), .S(i_reset_), .D(n64), .Q(o_label2_config[8]), .QN( ));
Q_MX02 U278 ( .S(n145), .A0(o_label2_config[8]), .A1(n2), .Z(n64));
Q_FDP2 \o_label3_config_REG[8] ( .CK(clk), .S(i_reset_), .D(n65), .Q(o_label3_config[8]), .QN( ));
Q_MX02 U280 ( .S(n154), .A0(o_label3_config[8]), .A1(n2), .Z(n65));
Q_FDP2 \o_label4_config_REG[8] ( .CK(clk), .S(i_reset_), .D(n66), .Q(o_label4_config[8]), .QN( ));
Q_MX02 U282 ( .S(n163), .A0(o_label4_config[8]), .A1(n2), .Z(n66));
Q_FDP2 \o_label5_config_REG[8] ( .CK(clk), .S(i_reset_), .D(n67), .Q(o_label5_config[8]), .QN( ));
Q_MX02 U284 ( .S(n172), .A0(o_label5_config[8]), .A1(n2), .Z(n67));
Q_FDP2 \o_label6_config_REG[8] ( .CK(clk), .S(i_reset_), .D(n68), .Q(o_label6_config[8]), .QN( ));
Q_MX02 U286 ( .S(n181), .A0(o_label6_config[8]), .A1(n2), .Z(n68));
Q_FDP2 \o_label7_config_REG[8] ( .CK(clk), .S(i_reset_), .D(n69), .Q(o_label7_config[8]), .QN( ));
Q_MX02 U288 ( .S(n190), .A0(o_label7_config[8]), .A1(n2), .Z(n69));
Q_FDP2 \o_bimc_global_config_REG[0] ( .CK(clk), .S(i_reset_), .D(n70), .Q(o_bimc_global_config[0]), .QN( ));
Q_MX02 U290 ( .S(n235), .A0(o_bimc_global_config[0]), .A1(n1), .Z(n70));
Q_INV U291 ( .A(i_sw_init), .Z(n71));
Q_OR02 U292 ( .A0(i_sw_init), .A1(w_load_spare_config), .Z(n72));
Q_OR02 U293 ( .A0(i_sw_init), .A1(w_load_cceip0_out_ia_wdata_part0), .Z(n73));
Q_OR02 U294 ( .A0(i_sw_init), .A1(w_load_cceip0_out_ia_wdata_part1), .Z(n74));
Q_OR02 U295 ( .A0(i_sw_init), .A1(w_load_cceip0_out_ia_wdata_part2), .Z(n75));
Q_OR02 U296 ( .A0(i_sw_init), .A1(w_load_cceip0_out_ia_config), .Z(n76));
Q_OR02 U297 ( .A0(i_sw_init), .A1(w_load_cceip0_out_im_config), .Z(n77));
Q_OR02 U298 ( .A0(i_sw_init), .A1(w_load_cceip0_out_im_read_done), .Z(n78));
Q_OR02 U299 ( .A0(i_sw_init), .A1(w_load_cceip1_out_ia_wdata_part0), .Z(n79));
Q_OR02 U300 ( .A0(i_sw_init), .A1(w_load_cceip1_out_ia_wdata_part1), .Z(n80));
Q_OR02 U301 ( .A0(i_sw_init), .A1(w_load_cceip1_out_ia_wdata_part2), .Z(n81));
Q_OR02 U302 ( .A0(i_sw_init), .A1(w_load_cceip1_out_ia_config), .Z(n82));
Q_OR02 U303 ( .A0(i_sw_init), .A1(w_load_cceip1_out_im_config), .Z(n83));
Q_OR02 U304 ( .A0(i_sw_init), .A1(w_load_cceip1_out_im_read_done), .Z(n84));
Q_OR02 U305 ( .A0(i_sw_init), .A1(w_load_cceip2_out_ia_wdata_part0), .Z(n85));
Q_OR02 U306 ( .A0(i_sw_init), .A1(w_load_cceip2_out_ia_wdata_part1), .Z(n86));
Q_OR02 U307 ( .A0(i_sw_init), .A1(w_load_cceip2_out_ia_wdata_part2), .Z(n87));
Q_OR02 U308 ( .A0(i_sw_init), .A1(w_load_cceip2_out_ia_config), .Z(n88));
Q_OR02 U309 ( .A0(i_sw_init), .A1(w_load_cceip2_out_im_config), .Z(n89));
Q_OR02 U310 ( .A0(i_sw_init), .A1(w_load_cceip2_out_im_read_done), .Z(n90));
Q_OR02 U311 ( .A0(i_sw_init), .A1(w_load_cceip3_out_ia_wdata_part0), .Z(n91));
Q_OR02 U312 ( .A0(i_sw_init), .A1(w_load_cceip3_out_ia_wdata_part1), .Z(n92));
Q_OR02 U313 ( .A0(i_sw_init), .A1(w_load_cceip3_out_ia_wdata_part2), .Z(n93));
Q_OR02 U314 ( .A0(i_sw_init), .A1(w_load_cceip3_out_ia_config), .Z(n94));
Q_OR02 U315 ( .A0(i_sw_init), .A1(w_load_cceip3_out_im_config), .Z(n95));
Q_OR02 U316 ( .A0(i_sw_init), .A1(w_load_cceip3_out_im_read_done), .Z(n96));
Q_OR02 U317 ( .A0(i_sw_init), .A1(w_load_cddip0_out_ia_wdata_part0), .Z(n97));
Q_OR02 U318 ( .A0(i_sw_init), .A1(w_load_cddip0_out_ia_wdata_part1), .Z(n98));
Q_OR02 U319 ( .A0(i_sw_init), .A1(w_load_cddip0_out_ia_wdata_part2), .Z(n99));
Q_OR02 U320 ( .A0(i_sw_init), .A1(w_load_cddip0_out_ia_config), .Z(n100));
Q_OR02 U321 ( .A0(i_sw_init), .A1(w_load_cddip0_out_im_config), .Z(n101));
Q_OR02 U322 ( .A0(i_sw_init), .A1(w_load_cddip0_out_im_read_done), .Z(n102));
Q_OR02 U323 ( .A0(i_sw_init), .A1(w_load_cddip1_out_ia_wdata_part0), .Z(n103));
Q_OR02 U324 ( .A0(i_sw_init), .A1(w_load_cddip1_out_ia_wdata_part1), .Z(n104));
Q_OR02 U325 ( .A0(i_sw_init), .A1(w_load_cddip1_out_ia_wdata_part2), .Z(n105));
Q_OR02 U326 ( .A0(i_sw_init), .A1(w_load_cddip1_out_ia_config), .Z(n106));
Q_OR02 U327 ( .A0(i_sw_init), .A1(w_load_cddip1_out_im_config), .Z(n107));
Q_OR02 U328 ( .A0(i_sw_init), .A1(w_load_cddip1_out_im_read_done), .Z(n108));
Q_OR02 U329 ( .A0(i_sw_init), .A1(w_load_cddip2_out_ia_wdata_part0), .Z(n109));
Q_OR02 U330 ( .A0(i_sw_init), .A1(w_load_cddip2_out_ia_wdata_part1), .Z(n110));
Q_OR02 U331 ( .A0(i_sw_init), .A1(w_load_cddip2_out_ia_wdata_part2), .Z(n111));
Q_OR02 U332 ( .A0(i_sw_init), .A1(w_load_cddip2_out_ia_config), .Z(n112));
Q_OR02 U333 ( .A0(i_sw_init), .A1(w_load_cddip2_out_im_config), .Z(n113));
Q_OR02 U334 ( .A0(i_sw_init), .A1(w_load_cddip2_out_im_read_done), .Z(n114));
Q_OR02 U335 ( .A0(i_sw_init), .A1(w_load_cddip3_out_ia_wdata_part0), .Z(n115));
Q_OR02 U336 ( .A0(i_sw_init), .A1(w_load_cddip3_out_ia_wdata_part1), .Z(n116));
Q_OR02 U337 ( .A0(i_sw_init), .A1(w_load_cddip3_out_ia_wdata_part2), .Z(n117));
Q_OR02 U338 ( .A0(i_sw_init), .A1(w_load_cddip3_out_ia_config), .Z(n118));
Q_OR02 U339 ( .A0(i_sw_init), .A1(w_load_cddip3_out_im_config), .Z(n119));
Q_OR02 U340 ( .A0(i_sw_init), .A1(w_load_cddip3_out_im_read_done), .Z(n120));
Q_OR02 U341 ( .A0(i_sw_init), .A1(w_load_ckv_ia_wdata_part0), .Z(n121));
Q_OR02 U342 ( .A0(i_sw_init), .A1(w_load_ckv_ia_wdata_part1), .Z(n122));
Q_OR02 U343 ( .A0(i_sw_init), .A1(w_load_ckv_ia_config), .Z(n123));
Q_OR02 U344 ( .A0(i_sw_init), .A1(w_load_kim_ia_wdata_part0), .Z(n124));
Q_OR02 U345 ( .A0(i_sw_init), .A1(w_load_kim_ia_wdata_part1), .Z(n125));
Q_OR02 U346 ( .A0(i_sw_init), .A1(w_load_kim_ia_config), .Z(n126));
Q_OR02 U347 ( .A0(i_sw_init), .A1(w_load_label0_config), .Z(n127));
Q_OR02 U348 ( .A0(i_sw_init), .A1(w_load_label0_data7), .Z(n128));
Q_OR02 U349 ( .A0(i_sw_init), .A1(w_load_label0_data6), .Z(n129));
Q_OR02 U350 ( .A0(i_sw_init), .A1(w_load_label0_data5), .Z(n130));
Q_OR02 U351 ( .A0(i_sw_init), .A1(w_load_label0_data4), .Z(n131));
Q_OR02 U352 ( .A0(i_sw_init), .A1(w_load_label0_data3), .Z(n132));
Q_OR02 U353 ( .A0(i_sw_init), .A1(w_load_label0_data2), .Z(n133));
Q_OR02 U354 ( .A0(i_sw_init), .A1(w_load_label0_data1), .Z(n134));
Q_OR02 U355 ( .A0(i_sw_init), .A1(w_load_label0_data0), .Z(n135));
Q_OR02 U356 ( .A0(i_sw_init), .A1(w_load_label1_config), .Z(n136));
Q_OR02 U357 ( .A0(i_sw_init), .A1(w_load_label1_data7), .Z(n137));
Q_OR02 U358 ( .A0(i_sw_init), .A1(w_load_label1_data6), .Z(n138));
Q_OR02 U359 ( .A0(i_sw_init), .A1(w_load_label1_data5), .Z(n139));
Q_OR02 U360 ( .A0(i_sw_init), .A1(w_load_label1_data4), .Z(n140));
Q_OR02 U361 ( .A0(i_sw_init), .A1(w_load_label1_data3), .Z(n141));
Q_OR02 U362 ( .A0(i_sw_init), .A1(w_load_label1_data2), .Z(n142));
Q_OR02 U363 ( .A0(i_sw_init), .A1(w_load_label1_data1), .Z(n143));
Q_OR02 U364 ( .A0(i_sw_init), .A1(w_load_label1_data0), .Z(n144));
Q_OR02 U365 ( .A0(i_sw_init), .A1(w_load_label2_config), .Z(n145));
Q_OR02 U366 ( .A0(i_sw_init), .A1(w_load_label2_data7), .Z(n146));
Q_OR02 U367 ( .A0(i_sw_init), .A1(w_load_label2_data6), .Z(n147));
Q_OR02 U368 ( .A0(i_sw_init), .A1(w_load_label2_data5), .Z(n148));
Q_OR02 U369 ( .A0(i_sw_init), .A1(w_load_label2_data4), .Z(n149));
Q_OR02 U370 ( .A0(i_sw_init), .A1(w_load_label2_data3), .Z(n150));
Q_OR02 U371 ( .A0(i_sw_init), .A1(w_load_label2_data2), .Z(n151));
Q_OR02 U372 ( .A0(i_sw_init), .A1(w_load_label2_data1), .Z(n152));
Q_OR02 U373 ( .A0(i_sw_init), .A1(w_load_label2_data0), .Z(n153));
Q_OR02 U374 ( .A0(i_sw_init), .A1(w_load_label3_config), .Z(n154));
Q_OR02 U375 ( .A0(i_sw_init), .A1(w_load_label3_data7), .Z(n155));
Q_OR02 U376 ( .A0(i_sw_init), .A1(w_load_label3_data6), .Z(n156));
Q_OR02 U377 ( .A0(i_sw_init), .A1(w_load_label3_data5), .Z(n157));
Q_OR02 U378 ( .A0(i_sw_init), .A1(w_load_label3_data4), .Z(n158));
Q_OR02 U379 ( .A0(i_sw_init), .A1(w_load_label3_data3), .Z(n159));
Q_OR02 U380 ( .A0(i_sw_init), .A1(w_load_label3_data2), .Z(n160));
Q_OR02 U381 ( .A0(i_sw_init), .A1(w_load_label3_data1), .Z(n161));
Q_OR02 U382 ( .A0(i_sw_init), .A1(w_load_label3_data0), .Z(n162));
Q_OR02 U383 ( .A0(i_sw_init), .A1(w_load_label4_config), .Z(n163));
Q_OR02 U384 ( .A0(i_sw_init), .A1(w_load_label4_data7), .Z(n164));
Q_OR02 U385 ( .A0(i_sw_init), .A1(w_load_label4_data6), .Z(n165));
Q_OR02 U386 ( .A0(i_sw_init), .A1(w_load_label4_data5), .Z(n166));
Q_OR02 U387 ( .A0(i_sw_init), .A1(w_load_label4_data4), .Z(n167));
Q_OR02 U388 ( .A0(i_sw_init), .A1(w_load_label4_data3), .Z(n168));
Q_OR02 U389 ( .A0(i_sw_init), .A1(w_load_label4_data2), .Z(n169));
Q_OR02 U390 ( .A0(i_sw_init), .A1(w_load_label4_data1), .Z(n170));
Q_OR02 U391 ( .A0(i_sw_init), .A1(w_load_label4_data0), .Z(n171));
Q_OR02 U392 ( .A0(i_sw_init), .A1(w_load_label5_config), .Z(n172));
Q_OR02 U393 ( .A0(i_sw_init), .A1(w_load_label5_data7), .Z(n173));
Q_OR02 U394 ( .A0(i_sw_init), .A1(w_load_label5_data6), .Z(n174));
Q_OR02 U395 ( .A0(i_sw_init), .A1(w_load_label5_data5), .Z(n175));
Q_OR02 U396 ( .A0(i_sw_init), .A1(w_load_label5_data4), .Z(n176));
Q_OR02 U397 ( .A0(i_sw_init), .A1(w_load_label5_data3), .Z(n177));
Q_OR02 U398 ( .A0(i_sw_init), .A1(w_load_label5_data2), .Z(n178));
Q_OR02 U399 ( .A0(i_sw_init), .A1(w_load_label5_data1), .Z(n179));
Q_OR02 U400 ( .A0(i_sw_init), .A1(w_load_label5_data0), .Z(n180));
Q_OR02 U401 ( .A0(i_sw_init), .A1(w_load_label6_config), .Z(n181));
Q_OR02 U402 ( .A0(i_sw_init), .A1(w_load_label6_data7), .Z(n182));
Q_OR02 U403 ( .A0(i_sw_init), .A1(w_load_label6_data6), .Z(n183));
Q_OR02 U404 ( .A0(i_sw_init), .A1(w_load_label6_data5), .Z(n184));
Q_OR02 U405 ( .A0(i_sw_init), .A1(w_load_label6_data4), .Z(n185));
Q_OR02 U406 ( .A0(i_sw_init), .A1(w_load_label6_data3), .Z(n186));
Q_OR02 U407 ( .A0(i_sw_init), .A1(w_load_label6_data2), .Z(n187));
Q_OR02 U408 ( .A0(i_sw_init), .A1(w_load_label6_data1), .Z(n188));
Q_OR02 U409 ( .A0(i_sw_init), .A1(w_load_label6_data0), .Z(n189));
Q_OR02 U410 ( .A0(i_sw_init), .A1(w_load_label7_config), .Z(n190));
Q_OR02 U411 ( .A0(i_sw_init), .A1(w_load_label7_data7), .Z(n191));
Q_OR02 U412 ( .A0(i_sw_init), .A1(w_load_label7_data6), .Z(n192));
Q_OR02 U413 ( .A0(i_sw_init), .A1(w_load_label7_data5), .Z(n193));
Q_OR02 U414 ( .A0(i_sw_init), .A1(w_load_label7_data4), .Z(n194));
Q_OR02 U415 ( .A0(i_sw_init), .A1(w_load_label7_data3), .Z(n195));
Q_OR02 U416 ( .A0(i_sw_init), .A1(w_load_label7_data2), .Z(n196));
Q_OR02 U417 ( .A0(i_sw_init), .A1(w_load_label7_data1), .Z(n197));
Q_OR02 U418 ( .A0(i_sw_init), .A1(w_load_label7_data0), .Z(n198));
Q_OR02 U419 ( .A0(i_sw_init), .A1(w_load_kdf_drbg_ctrl), .Z(n199));
Q_OR02 U420 ( .A0(i_sw_init), .A1(w_load_kdf_drbg_seed_0_state_key_31_0), .Z(n200));
Q_OR02 U421 ( .A0(i_sw_init), .A1(w_load_kdf_drbg_seed_0_state_key_63_32), .Z(n201));
Q_OR02 U422 ( .A0(i_sw_init), .A1(w_load_kdf_drbg_seed_0_state_key_95_64), .Z(n202));
Q_OR02 U423 ( .A0(i_sw_init), .A1(w_load_kdf_drbg_seed_0_state_key_127_96), .Z(n203));
Q_OR02 U424 ( .A0(i_sw_init), .A1(w_load_kdf_drbg_seed_0_state_key_159_128), .Z(n204));
Q_OR02 U425 ( .A0(i_sw_init), .A1(w_load_kdf_drbg_seed_0_state_key_191_160), .Z(n205));
Q_OR02 U426 ( .A0(i_sw_init), .A1(w_load_kdf_drbg_seed_0_state_key_223_192), .Z(n206));
Q_OR02 U427 ( .A0(i_sw_init), .A1(w_load_kdf_drbg_seed_0_state_key_255_224), .Z(n207));
Q_OR02 U428 ( .A0(i_sw_init), .A1(w_load_kdf_drbg_seed_0_state_value_31_0), .Z(n208));
Q_OR02 U429 ( .A0(i_sw_init), .A1(w_load_kdf_drbg_seed_0_state_value_63_32), .Z(n209));
Q_OR02 U430 ( .A0(i_sw_init), .A1(w_load_kdf_drbg_seed_0_state_value_95_64), .Z(n210));
Q_OR02 U431 ( .A0(i_sw_init), .A1(w_load_kdf_drbg_seed_0_state_value_127_96), .Z(n211));
Q_OR02 U432 ( .A0(i_sw_init), .A1(w_load_kdf_drbg_seed_0_reseed_interval_0), .Z(n212));
Q_OR02 U433 ( .A0(i_sw_init), .A1(w_load_kdf_drbg_seed_0_reseed_interval_1), .Z(n213));
Q_OR02 U434 ( .A0(i_sw_init), .A1(w_load_kdf_drbg_seed_1_state_key_31_0), .Z(n214));
Q_OR02 U435 ( .A0(i_sw_init), .A1(w_load_kdf_drbg_seed_1_state_key_63_32), .Z(n215));
Q_OR02 U436 ( .A0(i_sw_init), .A1(w_load_kdf_drbg_seed_1_state_key_95_64), .Z(n216));
Q_OR02 U437 ( .A0(i_sw_init), .A1(w_load_kdf_drbg_seed_1_state_key_127_96), .Z(n217));
Q_OR02 U438 ( .A0(i_sw_init), .A1(w_load_kdf_drbg_seed_1_state_key_159_128), .Z(n218));
Q_OR02 U439 ( .A0(i_sw_init), .A1(w_load_kdf_drbg_seed_1_state_key_191_160), .Z(n219));
Q_OR02 U440 ( .A0(i_sw_init), .A1(w_load_kdf_drbg_seed_1_state_key_223_192), .Z(n220));
Q_OR02 U441 ( .A0(i_sw_init), .A1(w_load_kdf_drbg_seed_1_state_key_255_224), .Z(n221));
Q_OR02 U442 ( .A0(i_sw_init), .A1(w_load_kdf_drbg_seed_1_state_value_31_0), .Z(n222));
Q_OR02 U443 ( .A0(i_sw_init), .A1(w_load_kdf_drbg_seed_1_state_value_63_32), .Z(n223));
Q_OR02 U444 ( .A0(i_sw_init), .A1(w_load_kdf_drbg_seed_1_state_value_95_64), .Z(n224));
Q_OR02 U445 ( .A0(i_sw_init), .A1(w_load_kdf_drbg_seed_1_state_value_127_96), .Z(n225));
Q_OR02 U446 ( .A0(i_sw_init), .A1(w_load_kdf_drbg_seed_1_reseed_interval_0), .Z(n226));
Q_OR02 U447 ( .A0(i_sw_init), .A1(w_load_kdf_drbg_seed_1_reseed_interval_1), .Z(n227));
Q_OR02 U448 ( .A0(i_sw_init), .A1(w_load_interrupt_status), .Z(n228));
Q_OR02 U449 ( .A0(i_sw_init), .A1(w_load_interrupt_mask), .Z(n229));
Q_OR02 U450 ( .A0(i_sw_init), .A1(w_load_engine_sticky_status), .Z(n230));
Q_OR02 U451 ( .A0(i_sw_init), .A1(w_load_bimc_monitor_mask), .Z(n231));
Q_OR02 U452 ( .A0(i_sw_init), .A1(w_load_bimc_ecc_uncorrectable_error_cnt), .Z(n232));
Q_OR02 U453 ( .A0(i_sw_init), .A1(w_load_bimc_ecc_correctable_error_cnt), .Z(n233));
Q_OR02 U454 ( .A0(i_sw_init), .A1(w_load_bimc_parity_error_cnt), .Z(n234));
Q_OR02 U455 ( .A0(i_sw_init), .A1(w_load_bimc_global_config), .Z(n235));
Q_OR02 U456 ( .A0(i_sw_init), .A1(w_load_bimc_eccpar_debug), .Z(n236));
Q_OR02 U457 ( .A0(i_sw_init), .A1(w_load_bimc_cmd2), .Z(n237));
Q_OR02 U458 ( .A0(i_sw_init), .A1(w_load_bimc_cmd1), .Z(n238));
Q_OR02 U459 ( .A0(i_sw_init), .A1(w_load_bimc_cmd0), .Z(n239));
Q_OR02 U460 ( .A0(i_sw_init), .A1(w_load_bimc_rxcmd2), .Z(n240));
Q_OR02 U461 ( .A0(i_sw_init), .A1(w_load_bimc_rxrsp2), .Z(n241));
Q_OR02 U462 ( .A0(i_sw_init), .A1(w_load_bimc_pollrsp2), .Z(n242));
Q_OR02 U463 ( .A0(i_sw_init), .A1(w_load_bimc_dbgcmd2), .Z(n243));
Q_OR02 U464 ( .A0(i_sw_init), .A1(w_load_im_consumed), .Z(n244));
Q_OR02 U465 ( .A0(i_sw_init), .A1(w_load_tready_override), .Z(n245));
Q_OR02 U466 ( .A0(i_sw_init), .A1(w_load_regs_sa_ctrl), .Z(n246));
Q_OR02 U467 ( .A0(i_sw_init), .A1(w_load_sa_snapshot_ia_wdata_part0), .Z(n247));
Q_OR02 U468 ( .A0(i_sw_init), .A1(w_load_sa_snapshot_ia_wdata_part1), .Z(n248));
Q_OR02 U469 ( .A0(i_sw_init), .A1(w_load_sa_snapshot_ia_config), .Z(n249));
Q_OR02 U470 ( .A0(i_sw_init), .A1(w_load_sa_count_ia_wdata_part0), .Z(n250));
Q_OR02 U471 ( .A0(i_sw_init), .A1(w_load_sa_count_ia_wdata_part1), .Z(n251));
Q_OR02 U472 ( .A0(i_sw_init), .A1(w_load_sa_count_ia_config), .Z(n252));
Q_OR02 U473 ( .A0(i_sw_init), .A1(w_load_cceip_encrypt_kop_fifo_override), .Z(n253));
Q_OR02 U474 ( .A0(i_sw_init), .A1(w_load_cceip_validate_kop_fifo_override), .Z(n254));
Q_OR02 U475 ( .A0(i_sw_init), .A1(w_load_cddip_decrypt_kop_fifo_override), .Z(n255));
Q_OR02 U476 ( .A0(i_sw_init), .A1(w_load_sa_global_ctrl), .Z(n256));
Q_OR02 U477 ( .A0(i_sw_init), .A1(w_load_sa_ctrl_ia_wdata_part0), .Z(n257));
Q_OR02 U478 ( .A0(i_sw_init), .A1(w_load_sa_ctrl_ia_config), .Z(n258));
Q_OR02 U479 ( .A0(i_sw_init), .A1(w_load_kdf_test_key_size_config), .Z(n259));
Q_FDP4EP \o_bimc_dbgcmd2_REG[9] ( .CK(clk), .CE(w_load_bimc_dbgcmd2), .R(n260), .D(f32_data[9]), .Q(o_bimc_dbgcmd2[9]));
Q_FDP4EP \o_bimc_pollrsp2_REG[9] ( .CK(clk), .CE(w_load_bimc_pollrsp2), .R(n260), .D(f32_data[9]), .Q(o_bimc_pollrsp2[9]));
Q_FDP4EP \o_bimc_rxrsp2_REG[9] ( .CK(clk), .CE(w_load_bimc_rxrsp2), .R(n260), .D(f32_data[9]), .Q(o_bimc_rxrsp2[9]));
Q_FDP4EP \o_bimc_rxcmd2_REG[9] ( .CK(clk), .CE(w_load_bimc_rxcmd2), .R(n260), .D(f32_data[9]), .Q(o_bimc_rxcmd2[9]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[6] ( .CK(clk), .CE(w_load_cddip3_out_ia_wdata_part0), .R(n260), .D(f32_data[6]), .Q(o_cddip3_out_ia_wdata_part0[6]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[7] ( .CK(clk), .CE(w_load_cddip3_out_ia_wdata_part0), .R(n260), .D(f32_data[7]), .Q(o_cddip3_out_ia_wdata_part0[7]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[8] ( .CK(clk), .CE(w_load_cddip3_out_ia_wdata_part0), .R(n260), .D(f32_data[8]), .Q(o_cddip3_out_ia_wdata_part0[8]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[9] ( .CK(clk), .CE(w_load_cddip3_out_ia_wdata_part0), .R(n260), .D(f32_data[9]), .Q(o_cddip3_out_ia_wdata_part0[9]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[10] ( .CK(clk), .CE(w_load_cddip3_out_ia_wdata_part0), .R(n260), .D(f32_data[10]), .Q(o_cddip3_out_ia_wdata_part0[10]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[11] ( .CK(clk), .CE(w_load_cddip3_out_ia_wdata_part0), .R(n260), .D(f32_data[11]), .Q(o_cddip3_out_ia_wdata_part0[11]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[12] ( .CK(clk), .CE(w_load_cddip3_out_ia_wdata_part0), .R(n260), .D(f32_data[12]), .Q(o_cddip3_out_ia_wdata_part0[12]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[13] ( .CK(clk), .CE(w_load_cddip3_out_ia_wdata_part0), .R(n260), .D(f32_data[13]), .Q(o_cddip3_out_ia_wdata_part0[13]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[14] ( .CK(clk), .CE(w_load_cddip3_out_ia_wdata_part0), .R(n260), .D(f32_data[14]), .Q(o_cddip3_out_ia_wdata_part0[14]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[15] ( .CK(clk), .CE(w_load_cddip3_out_ia_wdata_part0), .R(n260), .D(f32_data[15]), .Q(o_cddip3_out_ia_wdata_part0[15]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[16] ( .CK(clk), .CE(w_load_cddip3_out_ia_wdata_part0), .R(n260), .D(f32_data[16]), .Q(o_cddip3_out_ia_wdata_part0[16]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[17] ( .CK(clk), .CE(w_load_cddip3_out_ia_wdata_part0), .R(n260), .D(f32_data[17]), .Q(o_cddip3_out_ia_wdata_part0[17]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[18] ( .CK(clk), .CE(w_load_cddip3_out_ia_wdata_part0), .R(n260), .D(f32_data[18]), .Q(o_cddip3_out_ia_wdata_part0[18]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[19] ( .CK(clk), .CE(w_load_cddip3_out_ia_wdata_part0), .R(n260), .D(f32_data[19]), .Q(o_cddip3_out_ia_wdata_part0[19]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[20] ( .CK(clk), .CE(w_load_cddip3_out_ia_wdata_part0), .R(n260), .D(f32_data[20]), .Q(o_cddip3_out_ia_wdata_part0[20]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[21] ( .CK(clk), .CE(w_load_cddip3_out_ia_wdata_part0), .R(n260), .D(f32_data[21]), .Q(o_cddip3_out_ia_wdata_part0[21]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[22] ( .CK(clk), .CE(w_load_cddip3_out_ia_wdata_part0), .R(n260), .D(f32_data[22]), .Q(o_cddip3_out_ia_wdata_part0[22]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[23] ( .CK(clk), .CE(w_load_cddip3_out_ia_wdata_part0), .R(n260), .D(f32_data[23]), .Q(o_cddip3_out_ia_wdata_part0[23]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[24] ( .CK(clk), .CE(w_load_cddip3_out_ia_wdata_part0), .R(n260), .D(f32_data[24]), .Q(o_cddip3_out_ia_wdata_part0[24]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[25] ( .CK(clk), .CE(w_load_cddip3_out_ia_wdata_part0), .R(n260), .D(f32_data[25]), .Q(o_cddip3_out_ia_wdata_part0[25]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[26] ( .CK(clk), .CE(w_load_cddip3_out_ia_wdata_part0), .R(n260), .D(f32_data[26]), .Q(o_cddip3_out_ia_wdata_part0[26]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[27] ( .CK(clk), .CE(w_load_cddip3_out_ia_wdata_part0), .R(n260), .D(f32_data[27]), .Q(o_cddip3_out_ia_wdata_part0[27]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[28] ( .CK(clk), .CE(w_load_cddip3_out_ia_wdata_part0), .R(n260), .D(f32_data[28]), .Q(o_cddip3_out_ia_wdata_part0[28]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[29] ( .CK(clk), .CE(w_load_cddip3_out_ia_wdata_part0), .R(n260), .D(f32_data[29]), .Q(o_cddip3_out_ia_wdata_part0[29]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[30] ( .CK(clk), .CE(w_load_cddip3_out_ia_wdata_part0), .R(n260), .D(f32_data[30]), .Q(o_cddip3_out_ia_wdata_part0[30]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[31] ( .CK(clk), .CE(w_load_cddip3_out_ia_wdata_part0), .R(n260), .D(f32_data[31]), .Q(o_cddip3_out_ia_wdata_part0[31]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[6] ( .CK(clk), .CE(w_load_cddip2_out_ia_wdata_part0), .R(n260), .D(f32_data[6]), .Q(o_cddip2_out_ia_wdata_part0[6]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[7] ( .CK(clk), .CE(w_load_cddip2_out_ia_wdata_part0), .R(n260), .D(f32_data[7]), .Q(o_cddip2_out_ia_wdata_part0[7]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[8] ( .CK(clk), .CE(w_load_cddip2_out_ia_wdata_part0), .R(n260), .D(f32_data[8]), .Q(o_cddip2_out_ia_wdata_part0[8]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[9] ( .CK(clk), .CE(w_load_cddip2_out_ia_wdata_part0), .R(n260), .D(f32_data[9]), .Q(o_cddip2_out_ia_wdata_part0[9]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[10] ( .CK(clk), .CE(w_load_cddip2_out_ia_wdata_part0), .R(n260), .D(f32_data[10]), .Q(o_cddip2_out_ia_wdata_part0[10]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[11] ( .CK(clk), .CE(w_load_cddip2_out_ia_wdata_part0), .R(n260), .D(f32_data[11]), .Q(o_cddip2_out_ia_wdata_part0[11]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[12] ( .CK(clk), .CE(w_load_cddip2_out_ia_wdata_part0), .R(n260), .D(f32_data[12]), .Q(o_cddip2_out_ia_wdata_part0[12]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[13] ( .CK(clk), .CE(w_load_cddip2_out_ia_wdata_part0), .R(n260), .D(f32_data[13]), .Q(o_cddip2_out_ia_wdata_part0[13]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[14] ( .CK(clk), .CE(w_load_cddip2_out_ia_wdata_part0), .R(n260), .D(f32_data[14]), .Q(o_cddip2_out_ia_wdata_part0[14]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[15] ( .CK(clk), .CE(w_load_cddip2_out_ia_wdata_part0), .R(n260), .D(f32_data[15]), .Q(o_cddip2_out_ia_wdata_part0[15]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[16] ( .CK(clk), .CE(w_load_cddip2_out_ia_wdata_part0), .R(n260), .D(f32_data[16]), .Q(o_cddip2_out_ia_wdata_part0[16]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[17] ( .CK(clk), .CE(w_load_cddip2_out_ia_wdata_part0), .R(n260), .D(f32_data[17]), .Q(o_cddip2_out_ia_wdata_part0[17]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[18] ( .CK(clk), .CE(w_load_cddip2_out_ia_wdata_part0), .R(n260), .D(f32_data[18]), .Q(o_cddip2_out_ia_wdata_part0[18]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[19] ( .CK(clk), .CE(w_load_cddip2_out_ia_wdata_part0), .R(n260), .D(f32_data[19]), .Q(o_cddip2_out_ia_wdata_part0[19]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[20] ( .CK(clk), .CE(w_load_cddip2_out_ia_wdata_part0), .R(n260), .D(f32_data[20]), .Q(o_cddip2_out_ia_wdata_part0[20]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[21] ( .CK(clk), .CE(w_load_cddip2_out_ia_wdata_part0), .R(n260), .D(f32_data[21]), .Q(o_cddip2_out_ia_wdata_part0[21]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[22] ( .CK(clk), .CE(w_load_cddip2_out_ia_wdata_part0), .R(n260), .D(f32_data[22]), .Q(o_cddip2_out_ia_wdata_part0[22]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[23] ( .CK(clk), .CE(w_load_cddip2_out_ia_wdata_part0), .R(n260), .D(f32_data[23]), .Q(o_cddip2_out_ia_wdata_part0[23]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[24] ( .CK(clk), .CE(w_load_cddip2_out_ia_wdata_part0), .R(n260), .D(f32_data[24]), .Q(o_cddip2_out_ia_wdata_part0[24]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[25] ( .CK(clk), .CE(w_load_cddip2_out_ia_wdata_part0), .R(n260), .D(f32_data[25]), .Q(o_cddip2_out_ia_wdata_part0[25]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[26] ( .CK(clk), .CE(w_load_cddip2_out_ia_wdata_part0), .R(n260), .D(f32_data[26]), .Q(o_cddip2_out_ia_wdata_part0[26]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[27] ( .CK(clk), .CE(w_load_cddip2_out_ia_wdata_part0), .R(n260), .D(f32_data[27]), .Q(o_cddip2_out_ia_wdata_part0[27]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[28] ( .CK(clk), .CE(w_load_cddip2_out_ia_wdata_part0), .R(n260), .D(f32_data[28]), .Q(o_cddip2_out_ia_wdata_part0[28]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[29] ( .CK(clk), .CE(w_load_cddip2_out_ia_wdata_part0), .R(n260), .D(f32_data[29]), .Q(o_cddip2_out_ia_wdata_part0[29]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[30] ( .CK(clk), .CE(w_load_cddip2_out_ia_wdata_part0), .R(n260), .D(f32_data[30]), .Q(o_cddip2_out_ia_wdata_part0[30]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[31] ( .CK(clk), .CE(w_load_cddip2_out_ia_wdata_part0), .R(n260), .D(f32_data[31]), .Q(o_cddip2_out_ia_wdata_part0[31]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[6] ( .CK(clk), .CE(w_load_cddip1_out_ia_wdata_part0), .R(n260), .D(f32_data[6]), .Q(o_cddip1_out_ia_wdata_part0[6]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[7] ( .CK(clk), .CE(w_load_cddip1_out_ia_wdata_part0), .R(n260), .D(f32_data[7]), .Q(o_cddip1_out_ia_wdata_part0[7]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[8] ( .CK(clk), .CE(w_load_cddip1_out_ia_wdata_part0), .R(n260), .D(f32_data[8]), .Q(o_cddip1_out_ia_wdata_part0[8]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[9] ( .CK(clk), .CE(w_load_cddip1_out_ia_wdata_part0), .R(n260), .D(f32_data[9]), .Q(o_cddip1_out_ia_wdata_part0[9]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[10] ( .CK(clk), .CE(w_load_cddip1_out_ia_wdata_part0), .R(n260), .D(f32_data[10]), .Q(o_cddip1_out_ia_wdata_part0[10]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[11] ( .CK(clk), .CE(w_load_cddip1_out_ia_wdata_part0), .R(n260), .D(f32_data[11]), .Q(o_cddip1_out_ia_wdata_part0[11]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[12] ( .CK(clk), .CE(w_load_cddip1_out_ia_wdata_part0), .R(n260), .D(f32_data[12]), .Q(o_cddip1_out_ia_wdata_part0[12]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[13] ( .CK(clk), .CE(w_load_cddip1_out_ia_wdata_part0), .R(n260), .D(f32_data[13]), .Q(o_cddip1_out_ia_wdata_part0[13]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[14] ( .CK(clk), .CE(w_load_cddip1_out_ia_wdata_part0), .R(n260), .D(f32_data[14]), .Q(o_cddip1_out_ia_wdata_part0[14]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[15] ( .CK(clk), .CE(w_load_cddip1_out_ia_wdata_part0), .R(n260), .D(f32_data[15]), .Q(o_cddip1_out_ia_wdata_part0[15]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[16] ( .CK(clk), .CE(w_load_cddip1_out_ia_wdata_part0), .R(n260), .D(f32_data[16]), .Q(o_cddip1_out_ia_wdata_part0[16]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[17] ( .CK(clk), .CE(w_load_cddip1_out_ia_wdata_part0), .R(n260), .D(f32_data[17]), .Q(o_cddip1_out_ia_wdata_part0[17]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[18] ( .CK(clk), .CE(w_load_cddip1_out_ia_wdata_part0), .R(n260), .D(f32_data[18]), .Q(o_cddip1_out_ia_wdata_part0[18]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[19] ( .CK(clk), .CE(w_load_cddip1_out_ia_wdata_part0), .R(n260), .D(f32_data[19]), .Q(o_cddip1_out_ia_wdata_part0[19]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[20] ( .CK(clk), .CE(w_load_cddip1_out_ia_wdata_part0), .R(n260), .D(f32_data[20]), .Q(o_cddip1_out_ia_wdata_part0[20]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[21] ( .CK(clk), .CE(w_load_cddip1_out_ia_wdata_part0), .R(n260), .D(f32_data[21]), .Q(o_cddip1_out_ia_wdata_part0[21]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[22] ( .CK(clk), .CE(w_load_cddip1_out_ia_wdata_part0), .R(n260), .D(f32_data[22]), .Q(o_cddip1_out_ia_wdata_part0[22]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[23] ( .CK(clk), .CE(w_load_cddip1_out_ia_wdata_part0), .R(n260), .D(f32_data[23]), .Q(o_cddip1_out_ia_wdata_part0[23]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[24] ( .CK(clk), .CE(w_load_cddip1_out_ia_wdata_part0), .R(n260), .D(f32_data[24]), .Q(o_cddip1_out_ia_wdata_part0[24]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[25] ( .CK(clk), .CE(w_load_cddip1_out_ia_wdata_part0), .R(n260), .D(f32_data[25]), .Q(o_cddip1_out_ia_wdata_part0[25]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[26] ( .CK(clk), .CE(w_load_cddip1_out_ia_wdata_part0), .R(n260), .D(f32_data[26]), .Q(o_cddip1_out_ia_wdata_part0[26]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[27] ( .CK(clk), .CE(w_load_cddip1_out_ia_wdata_part0), .R(n260), .D(f32_data[27]), .Q(o_cddip1_out_ia_wdata_part0[27]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[28] ( .CK(clk), .CE(w_load_cddip1_out_ia_wdata_part0), .R(n260), .D(f32_data[28]), .Q(o_cddip1_out_ia_wdata_part0[28]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[29] ( .CK(clk), .CE(w_load_cddip1_out_ia_wdata_part0), .R(n260), .D(f32_data[29]), .Q(o_cddip1_out_ia_wdata_part0[29]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[30] ( .CK(clk), .CE(w_load_cddip1_out_ia_wdata_part0), .R(n260), .D(f32_data[30]), .Q(o_cddip1_out_ia_wdata_part0[30]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[31] ( .CK(clk), .CE(w_load_cddip1_out_ia_wdata_part0), .R(n260), .D(f32_data[31]), .Q(o_cddip1_out_ia_wdata_part0[31]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[6] ( .CK(clk), .CE(w_load_cddip0_out_ia_wdata_part0), .R(n260), .D(f32_data[6]), .Q(o_cddip0_out_ia_wdata_part0[6]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[7] ( .CK(clk), .CE(w_load_cddip0_out_ia_wdata_part0), .R(n260), .D(f32_data[7]), .Q(o_cddip0_out_ia_wdata_part0[7]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[8] ( .CK(clk), .CE(w_load_cddip0_out_ia_wdata_part0), .R(n260), .D(f32_data[8]), .Q(o_cddip0_out_ia_wdata_part0[8]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[9] ( .CK(clk), .CE(w_load_cddip0_out_ia_wdata_part0), .R(n260), .D(f32_data[9]), .Q(o_cddip0_out_ia_wdata_part0[9]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[10] ( .CK(clk), .CE(w_load_cddip0_out_ia_wdata_part0), .R(n260), .D(f32_data[10]), .Q(o_cddip0_out_ia_wdata_part0[10]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[11] ( .CK(clk), .CE(w_load_cddip0_out_ia_wdata_part0), .R(n260), .D(f32_data[11]), .Q(o_cddip0_out_ia_wdata_part0[11]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[12] ( .CK(clk), .CE(w_load_cddip0_out_ia_wdata_part0), .R(n260), .D(f32_data[12]), .Q(o_cddip0_out_ia_wdata_part0[12]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[13] ( .CK(clk), .CE(w_load_cddip0_out_ia_wdata_part0), .R(n260), .D(f32_data[13]), .Q(o_cddip0_out_ia_wdata_part0[13]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[14] ( .CK(clk), .CE(w_load_cddip0_out_ia_wdata_part0), .R(n260), .D(f32_data[14]), .Q(o_cddip0_out_ia_wdata_part0[14]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[15] ( .CK(clk), .CE(w_load_cddip0_out_ia_wdata_part0), .R(n260), .D(f32_data[15]), .Q(o_cddip0_out_ia_wdata_part0[15]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[16] ( .CK(clk), .CE(w_load_cddip0_out_ia_wdata_part0), .R(n260), .D(f32_data[16]), .Q(o_cddip0_out_ia_wdata_part0[16]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[17] ( .CK(clk), .CE(w_load_cddip0_out_ia_wdata_part0), .R(n260), .D(f32_data[17]), .Q(o_cddip0_out_ia_wdata_part0[17]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[18] ( .CK(clk), .CE(w_load_cddip0_out_ia_wdata_part0), .R(n260), .D(f32_data[18]), .Q(o_cddip0_out_ia_wdata_part0[18]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[19] ( .CK(clk), .CE(w_load_cddip0_out_ia_wdata_part0), .R(n260), .D(f32_data[19]), .Q(o_cddip0_out_ia_wdata_part0[19]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[20] ( .CK(clk), .CE(w_load_cddip0_out_ia_wdata_part0), .R(n260), .D(f32_data[20]), .Q(o_cddip0_out_ia_wdata_part0[20]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[21] ( .CK(clk), .CE(w_load_cddip0_out_ia_wdata_part0), .R(n260), .D(f32_data[21]), .Q(o_cddip0_out_ia_wdata_part0[21]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[22] ( .CK(clk), .CE(w_load_cddip0_out_ia_wdata_part0), .R(n260), .D(f32_data[22]), .Q(o_cddip0_out_ia_wdata_part0[22]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[23] ( .CK(clk), .CE(w_load_cddip0_out_ia_wdata_part0), .R(n260), .D(f32_data[23]), .Q(o_cddip0_out_ia_wdata_part0[23]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[24] ( .CK(clk), .CE(w_load_cddip0_out_ia_wdata_part0), .R(n260), .D(f32_data[24]), .Q(o_cddip0_out_ia_wdata_part0[24]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[25] ( .CK(clk), .CE(w_load_cddip0_out_ia_wdata_part0), .R(n260), .D(f32_data[25]), .Q(o_cddip0_out_ia_wdata_part0[25]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[26] ( .CK(clk), .CE(w_load_cddip0_out_ia_wdata_part0), .R(n260), .D(f32_data[26]), .Q(o_cddip0_out_ia_wdata_part0[26]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[27] ( .CK(clk), .CE(w_load_cddip0_out_ia_wdata_part0), .R(n260), .D(f32_data[27]), .Q(o_cddip0_out_ia_wdata_part0[27]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[28] ( .CK(clk), .CE(w_load_cddip0_out_ia_wdata_part0), .R(n260), .D(f32_data[28]), .Q(o_cddip0_out_ia_wdata_part0[28]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[29] ( .CK(clk), .CE(w_load_cddip0_out_ia_wdata_part0), .R(n260), .D(f32_data[29]), .Q(o_cddip0_out_ia_wdata_part0[29]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[30] ( .CK(clk), .CE(w_load_cddip0_out_ia_wdata_part0), .R(n260), .D(f32_data[30]), .Q(o_cddip0_out_ia_wdata_part0[30]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[31] ( .CK(clk), .CE(w_load_cddip0_out_ia_wdata_part0), .R(n260), .D(f32_data[31]), .Q(o_cddip0_out_ia_wdata_part0[31]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[6] ( .CK(clk), .CE(w_load_cceip3_out_ia_wdata_part0), .R(n260), .D(f32_data[6]), .Q(o_cceip3_out_ia_wdata_part0[6]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[7] ( .CK(clk), .CE(w_load_cceip3_out_ia_wdata_part0), .R(n260), .D(f32_data[7]), .Q(o_cceip3_out_ia_wdata_part0[7]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[8] ( .CK(clk), .CE(w_load_cceip3_out_ia_wdata_part0), .R(n260), .D(f32_data[8]), .Q(o_cceip3_out_ia_wdata_part0[8]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[9] ( .CK(clk), .CE(w_load_cceip3_out_ia_wdata_part0), .R(n260), .D(f32_data[9]), .Q(o_cceip3_out_ia_wdata_part0[9]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[10] ( .CK(clk), .CE(w_load_cceip3_out_ia_wdata_part0), .R(n260), .D(f32_data[10]), .Q(o_cceip3_out_ia_wdata_part0[10]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[11] ( .CK(clk), .CE(w_load_cceip3_out_ia_wdata_part0), .R(n260), .D(f32_data[11]), .Q(o_cceip3_out_ia_wdata_part0[11]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[12] ( .CK(clk), .CE(w_load_cceip3_out_ia_wdata_part0), .R(n260), .D(f32_data[12]), .Q(o_cceip3_out_ia_wdata_part0[12]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[13] ( .CK(clk), .CE(w_load_cceip3_out_ia_wdata_part0), .R(n260), .D(f32_data[13]), .Q(o_cceip3_out_ia_wdata_part0[13]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[14] ( .CK(clk), .CE(w_load_cceip3_out_ia_wdata_part0), .R(n260), .D(f32_data[14]), .Q(o_cceip3_out_ia_wdata_part0[14]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[15] ( .CK(clk), .CE(w_load_cceip3_out_ia_wdata_part0), .R(n260), .D(f32_data[15]), .Q(o_cceip3_out_ia_wdata_part0[15]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[16] ( .CK(clk), .CE(w_load_cceip3_out_ia_wdata_part0), .R(n260), .D(f32_data[16]), .Q(o_cceip3_out_ia_wdata_part0[16]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[17] ( .CK(clk), .CE(w_load_cceip3_out_ia_wdata_part0), .R(n260), .D(f32_data[17]), .Q(o_cceip3_out_ia_wdata_part0[17]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[18] ( .CK(clk), .CE(w_load_cceip3_out_ia_wdata_part0), .R(n260), .D(f32_data[18]), .Q(o_cceip3_out_ia_wdata_part0[18]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[19] ( .CK(clk), .CE(w_load_cceip3_out_ia_wdata_part0), .R(n260), .D(f32_data[19]), .Q(o_cceip3_out_ia_wdata_part0[19]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[20] ( .CK(clk), .CE(w_load_cceip3_out_ia_wdata_part0), .R(n260), .D(f32_data[20]), .Q(o_cceip3_out_ia_wdata_part0[20]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[21] ( .CK(clk), .CE(w_load_cceip3_out_ia_wdata_part0), .R(n260), .D(f32_data[21]), .Q(o_cceip3_out_ia_wdata_part0[21]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[22] ( .CK(clk), .CE(w_load_cceip3_out_ia_wdata_part0), .R(n260), .D(f32_data[22]), .Q(o_cceip3_out_ia_wdata_part0[22]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[23] ( .CK(clk), .CE(w_load_cceip3_out_ia_wdata_part0), .R(n260), .D(f32_data[23]), .Q(o_cceip3_out_ia_wdata_part0[23]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[24] ( .CK(clk), .CE(w_load_cceip3_out_ia_wdata_part0), .R(n260), .D(f32_data[24]), .Q(o_cceip3_out_ia_wdata_part0[24]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[25] ( .CK(clk), .CE(w_load_cceip3_out_ia_wdata_part0), .R(n260), .D(f32_data[25]), .Q(o_cceip3_out_ia_wdata_part0[25]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[26] ( .CK(clk), .CE(w_load_cceip3_out_ia_wdata_part0), .R(n260), .D(f32_data[26]), .Q(o_cceip3_out_ia_wdata_part0[26]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[27] ( .CK(clk), .CE(w_load_cceip3_out_ia_wdata_part0), .R(n260), .D(f32_data[27]), .Q(o_cceip3_out_ia_wdata_part0[27]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[28] ( .CK(clk), .CE(w_load_cceip3_out_ia_wdata_part0), .R(n260), .D(f32_data[28]), .Q(o_cceip3_out_ia_wdata_part0[28]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[29] ( .CK(clk), .CE(w_load_cceip3_out_ia_wdata_part0), .R(n260), .D(f32_data[29]), .Q(o_cceip3_out_ia_wdata_part0[29]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[30] ( .CK(clk), .CE(w_load_cceip3_out_ia_wdata_part0), .R(n260), .D(f32_data[30]), .Q(o_cceip3_out_ia_wdata_part0[30]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[31] ( .CK(clk), .CE(w_load_cceip3_out_ia_wdata_part0), .R(n260), .D(f32_data[31]), .Q(o_cceip3_out_ia_wdata_part0[31]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[6] ( .CK(clk), .CE(w_load_cceip2_out_ia_wdata_part0), .R(n260), .D(f32_data[6]), .Q(o_cceip2_out_ia_wdata_part0[6]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[7] ( .CK(clk), .CE(w_load_cceip2_out_ia_wdata_part0), .R(n260), .D(f32_data[7]), .Q(o_cceip2_out_ia_wdata_part0[7]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[8] ( .CK(clk), .CE(w_load_cceip2_out_ia_wdata_part0), .R(n260), .D(f32_data[8]), .Q(o_cceip2_out_ia_wdata_part0[8]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[9] ( .CK(clk), .CE(w_load_cceip2_out_ia_wdata_part0), .R(n260), .D(f32_data[9]), .Q(o_cceip2_out_ia_wdata_part0[9]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[10] ( .CK(clk), .CE(w_load_cceip2_out_ia_wdata_part0), .R(n260), .D(f32_data[10]), .Q(o_cceip2_out_ia_wdata_part0[10]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[11] ( .CK(clk), .CE(w_load_cceip2_out_ia_wdata_part0), .R(n260), .D(f32_data[11]), .Q(o_cceip2_out_ia_wdata_part0[11]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[12] ( .CK(clk), .CE(w_load_cceip2_out_ia_wdata_part0), .R(n260), .D(f32_data[12]), .Q(o_cceip2_out_ia_wdata_part0[12]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[13] ( .CK(clk), .CE(w_load_cceip2_out_ia_wdata_part0), .R(n260), .D(f32_data[13]), .Q(o_cceip2_out_ia_wdata_part0[13]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[14] ( .CK(clk), .CE(w_load_cceip2_out_ia_wdata_part0), .R(n260), .D(f32_data[14]), .Q(o_cceip2_out_ia_wdata_part0[14]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[15] ( .CK(clk), .CE(w_load_cceip2_out_ia_wdata_part0), .R(n260), .D(f32_data[15]), .Q(o_cceip2_out_ia_wdata_part0[15]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[16] ( .CK(clk), .CE(w_load_cceip2_out_ia_wdata_part0), .R(n260), .D(f32_data[16]), .Q(o_cceip2_out_ia_wdata_part0[16]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[17] ( .CK(clk), .CE(w_load_cceip2_out_ia_wdata_part0), .R(n260), .D(f32_data[17]), .Q(o_cceip2_out_ia_wdata_part0[17]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[18] ( .CK(clk), .CE(w_load_cceip2_out_ia_wdata_part0), .R(n260), .D(f32_data[18]), .Q(o_cceip2_out_ia_wdata_part0[18]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[19] ( .CK(clk), .CE(w_load_cceip2_out_ia_wdata_part0), .R(n260), .D(f32_data[19]), .Q(o_cceip2_out_ia_wdata_part0[19]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[20] ( .CK(clk), .CE(w_load_cceip2_out_ia_wdata_part0), .R(n260), .D(f32_data[20]), .Q(o_cceip2_out_ia_wdata_part0[20]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[21] ( .CK(clk), .CE(w_load_cceip2_out_ia_wdata_part0), .R(n260), .D(f32_data[21]), .Q(o_cceip2_out_ia_wdata_part0[21]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[22] ( .CK(clk), .CE(w_load_cceip2_out_ia_wdata_part0), .R(n260), .D(f32_data[22]), .Q(o_cceip2_out_ia_wdata_part0[22]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[23] ( .CK(clk), .CE(w_load_cceip2_out_ia_wdata_part0), .R(n260), .D(f32_data[23]), .Q(o_cceip2_out_ia_wdata_part0[23]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[24] ( .CK(clk), .CE(w_load_cceip2_out_ia_wdata_part0), .R(n260), .D(f32_data[24]), .Q(o_cceip2_out_ia_wdata_part0[24]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[25] ( .CK(clk), .CE(w_load_cceip2_out_ia_wdata_part0), .R(n260), .D(f32_data[25]), .Q(o_cceip2_out_ia_wdata_part0[25]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[26] ( .CK(clk), .CE(w_load_cceip2_out_ia_wdata_part0), .R(n260), .D(f32_data[26]), .Q(o_cceip2_out_ia_wdata_part0[26]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[27] ( .CK(clk), .CE(w_load_cceip2_out_ia_wdata_part0), .R(n260), .D(f32_data[27]), .Q(o_cceip2_out_ia_wdata_part0[27]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[28] ( .CK(clk), .CE(w_load_cceip2_out_ia_wdata_part0), .R(n260), .D(f32_data[28]), .Q(o_cceip2_out_ia_wdata_part0[28]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[29] ( .CK(clk), .CE(w_load_cceip2_out_ia_wdata_part0), .R(n260), .D(f32_data[29]), .Q(o_cceip2_out_ia_wdata_part0[29]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[30] ( .CK(clk), .CE(w_load_cceip2_out_ia_wdata_part0), .R(n260), .D(f32_data[30]), .Q(o_cceip2_out_ia_wdata_part0[30]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[31] ( .CK(clk), .CE(w_load_cceip2_out_ia_wdata_part0), .R(n260), .D(f32_data[31]), .Q(o_cceip2_out_ia_wdata_part0[31]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[6] ( .CK(clk), .CE(w_load_cceip1_out_ia_wdata_part0), .R(n260), .D(f32_data[6]), .Q(o_cceip1_out_ia_wdata_part0[6]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[7] ( .CK(clk), .CE(w_load_cceip1_out_ia_wdata_part0), .R(n260), .D(f32_data[7]), .Q(o_cceip1_out_ia_wdata_part0[7]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[8] ( .CK(clk), .CE(w_load_cceip1_out_ia_wdata_part0), .R(n260), .D(f32_data[8]), .Q(o_cceip1_out_ia_wdata_part0[8]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[9] ( .CK(clk), .CE(w_load_cceip1_out_ia_wdata_part0), .R(n260), .D(f32_data[9]), .Q(o_cceip1_out_ia_wdata_part0[9]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[10] ( .CK(clk), .CE(w_load_cceip1_out_ia_wdata_part0), .R(n260), .D(f32_data[10]), .Q(o_cceip1_out_ia_wdata_part0[10]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[11] ( .CK(clk), .CE(w_load_cceip1_out_ia_wdata_part0), .R(n260), .D(f32_data[11]), .Q(o_cceip1_out_ia_wdata_part0[11]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[12] ( .CK(clk), .CE(w_load_cceip1_out_ia_wdata_part0), .R(n260), .D(f32_data[12]), .Q(o_cceip1_out_ia_wdata_part0[12]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[13] ( .CK(clk), .CE(w_load_cceip1_out_ia_wdata_part0), .R(n260), .D(f32_data[13]), .Q(o_cceip1_out_ia_wdata_part0[13]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[14] ( .CK(clk), .CE(w_load_cceip1_out_ia_wdata_part0), .R(n260), .D(f32_data[14]), .Q(o_cceip1_out_ia_wdata_part0[14]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[15] ( .CK(clk), .CE(w_load_cceip1_out_ia_wdata_part0), .R(n260), .D(f32_data[15]), .Q(o_cceip1_out_ia_wdata_part0[15]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[16] ( .CK(clk), .CE(w_load_cceip1_out_ia_wdata_part0), .R(n260), .D(f32_data[16]), .Q(o_cceip1_out_ia_wdata_part0[16]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[17] ( .CK(clk), .CE(w_load_cceip1_out_ia_wdata_part0), .R(n260), .D(f32_data[17]), .Q(o_cceip1_out_ia_wdata_part0[17]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[18] ( .CK(clk), .CE(w_load_cceip1_out_ia_wdata_part0), .R(n260), .D(f32_data[18]), .Q(o_cceip1_out_ia_wdata_part0[18]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[19] ( .CK(clk), .CE(w_load_cceip1_out_ia_wdata_part0), .R(n260), .D(f32_data[19]), .Q(o_cceip1_out_ia_wdata_part0[19]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[20] ( .CK(clk), .CE(w_load_cceip1_out_ia_wdata_part0), .R(n260), .D(f32_data[20]), .Q(o_cceip1_out_ia_wdata_part0[20]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[21] ( .CK(clk), .CE(w_load_cceip1_out_ia_wdata_part0), .R(n260), .D(f32_data[21]), .Q(o_cceip1_out_ia_wdata_part0[21]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[22] ( .CK(clk), .CE(w_load_cceip1_out_ia_wdata_part0), .R(n260), .D(f32_data[22]), .Q(o_cceip1_out_ia_wdata_part0[22]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[23] ( .CK(clk), .CE(w_load_cceip1_out_ia_wdata_part0), .R(n260), .D(f32_data[23]), .Q(o_cceip1_out_ia_wdata_part0[23]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[24] ( .CK(clk), .CE(w_load_cceip1_out_ia_wdata_part0), .R(n260), .D(f32_data[24]), .Q(o_cceip1_out_ia_wdata_part0[24]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[25] ( .CK(clk), .CE(w_load_cceip1_out_ia_wdata_part0), .R(n260), .D(f32_data[25]), .Q(o_cceip1_out_ia_wdata_part0[25]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[26] ( .CK(clk), .CE(w_load_cceip1_out_ia_wdata_part0), .R(n260), .D(f32_data[26]), .Q(o_cceip1_out_ia_wdata_part0[26]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[27] ( .CK(clk), .CE(w_load_cceip1_out_ia_wdata_part0), .R(n260), .D(f32_data[27]), .Q(o_cceip1_out_ia_wdata_part0[27]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[28] ( .CK(clk), .CE(w_load_cceip1_out_ia_wdata_part0), .R(n260), .D(f32_data[28]), .Q(o_cceip1_out_ia_wdata_part0[28]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[29] ( .CK(clk), .CE(w_load_cceip1_out_ia_wdata_part0), .R(n260), .D(f32_data[29]), .Q(o_cceip1_out_ia_wdata_part0[29]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[30] ( .CK(clk), .CE(w_load_cceip1_out_ia_wdata_part0), .R(n260), .D(f32_data[30]), .Q(o_cceip1_out_ia_wdata_part0[30]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[31] ( .CK(clk), .CE(w_load_cceip1_out_ia_wdata_part0), .R(n260), .D(f32_data[31]), .Q(o_cceip1_out_ia_wdata_part0[31]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[6] ( .CK(clk), .CE(w_load_cceip0_out_ia_wdata_part0), .R(n260), .D(f32_data[6]), .Q(o_cceip0_out_ia_wdata_part0[6]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[7] ( .CK(clk), .CE(w_load_cceip0_out_ia_wdata_part0), .R(n260), .D(f32_data[7]), .Q(o_cceip0_out_ia_wdata_part0[7]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[8] ( .CK(clk), .CE(w_load_cceip0_out_ia_wdata_part0), .R(n260), .D(f32_data[8]), .Q(o_cceip0_out_ia_wdata_part0[8]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[9] ( .CK(clk), .CE(w_load_cceip0_out_ia_wdata_part0), .R(n260), .D(f32_data[9]), .Q(o_cceip0_out_ia_wdata_part0[9]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[10] ( .CK(clk), .CE(w_load_cceip0_out_ia_wdata_part0), .R(n260), .D(f32_data[10]), .Q(o_cceip0_out_ia_wdata_part0[10]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[11] ( .CK(clk), .CE(w_load_cceip0_out_ia_wdata_part0), .R(n260), .D(f32_data[11]), .Q(o_cceip0_out_ia_wdata_part0[11]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[12] ( .CK(clk), .CE(w_load_cceip0_out_ia_wdata_part0), .R(n260), .D(f32_data[12]), .Q(o_cceip0_out_ia_wdata_part0[12]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[13] ( .CK(clk), .CE(w_load_cceip0_out_ia_wdata_part0), .R(n260), .D(f32_data[13]), .Q(o_cceip0_out_ia_wdata_part0[13]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[14] ( .CK(clk), .CE(w_load_cceip0_out_ia_wdata_part0), .R(n260), .D(f32_data[14]), .Q(o_cceip0_out_ia_wdata_part0[14]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[15] ( .CK(clk), .CE(w_load_cceip0_out_ia_wdata_part0), .R(n260), .D(f32_data[15]), .Q(o_cceip0_out_ia_wdata_part0[15]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[16] ( .CK(clk), .CE(w_load_cceip0_out_ia_wdata_part0), .R(n260), .D(f32_data[16]), .Q(o_cceip0_out_ia_wdata_part0[16]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[17] ( .CK(clk), .CE(w_load_cceip0_out_ia_wdata_part0), .R(n260), .D(f32_data[17]), .Q(o_cceip0_out_ia_wdata_part0[17]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[18] ( .CK(clk), .CE(w_load_cceip0_out_ia_wdata_part0), .R(n260), .D(f32_data[18]), .Q(o_cceip0_out_ia_wdata_part0[18]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[19] ( .CK(clk), .CE(w_load_cceip0_out_ia_wdata_part0), .R(n260), .D(f32_data[19]), .Q(o_cceip0_out_ia_wdata_part0[19]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[20] ( .CK(clk), .CE(w_load_cceip0_out_ia_wdata_part0), .R(n260), .D(f32_data[20]), .Q(o_cceip0_out_ia_wdata_part0[20]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[21] ( .CK(clk), .CE(w_load_cceip0_out_ia_wdata_part0), .R(n260), .D(f32_data[21]), .Q(o_cceip0_out_ia_wdata_part0[21]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[22] ( .CK(clk), .CE(w_load_cceip0_out_ia_wdata_part0), .R(n260), .D(f32_data[22]), .Q(o_cceip0_out_ia_wdata_part0[22]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[23] ( .CK(clk), .CE(w_load_cceip0_out_ia_wdata_part0), .R(n260), .D(f32_data[23]), .Q(o_cceip0_out_ia_wdata_part0[23]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[24] ( .CK(clk), .CE(w_load_cceip0_out_ia_wdata_part0), .R(n260), .D(f32_data[24]), .Q(o_cceip0_out_ia_wdata_part0[24]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[25] ( .CK(clk), .CE(w_load_cceip0_out_ia_wdata_part0), .R(n260), .D(f32_data[25]), .Q(o_cceip0_out_ia_wdata_part0[25]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[26] ( .CK(clk), .CE(w_load_cceip0_out_ia_wdata_part0), .R(n260), .D(f32_data[26]), .Q(o_cceip0_out_ia_wdata_part0[26]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[27] ( .CK(clk), .CE(w_load_cceip0_out_ia_wdata_part0), .R(n260), .D(f32_data[27]), .Q(o_cceip0_out_ia_wdata_part0[27]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[28] ( .CK(clk), .CE(w_load_cceip0_out_ia_wdata_part0), .R(n260), .D(f32_data[28]), .Q(o_cceip0_out_ia_wdata_part0[28]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[29] ( .CK(clk), .CE(w_load_cceip0_out_ia_wdata_part0), .R(n260), .D(f32_data[29]), .Q(o_cceip0_out_ia_wdata_part0[29]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[30] ( .CK(clk), .CE(w_load_cceip0_out_ia_wdata_part0), .R(n260), .D(f32_data[30]), .Q(o_cceip0_out_ia_wdata_part0[30]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[31] ( .CK(clk), .CE(w_load_cceip0_out_ia_wdata_part0), .R(n260), .D(f32_data[31]), .Q(o_cceip0_out_ia_wdata_part0[31]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[0] ( .CK(clk), .CE(n259), .R(n261), .D(n6), .Q(o_kdf_test_key_size_config[0]));
Q_INV U693 ( .A(i_reset_), .Z(n261));
Q_FDP4EP \o_kdf_test_key_size_config_REG[1] ( .CK(clk), .CE(n259), .R(n261), .D(n7), .Q(o_kdf_test_key_size_config[1]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[2] ( .CK(clk), .CE(n259), .R(n261), .D(n8), .Q(o_kdf_test_key_size_config[2]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[3] ( .CK(clk), .CE(n259), .R(n261), .D(n9), .Q(o_kdf_test_key_size_config[3]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[4] ( .CK(clk), .CE(n259), .R(n261), .D(n10), .Q(o_kdf_test_key_size_config[4]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[5] ( .CK(clk), .CE(n259), .R(n261), .D(n11), .Q(o_kdf_test_key_size_config[5]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[6] ( .CK(clk), .CE(n259), .R(n261), .D(n12), .Q(o_kdf_test_key_size_config[6]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[7] ( .CK(clk), .CE(n259), .R(n261), .D(n13), .Q(o_kdf_test_key_size_config[7]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[8] ( .CK(clk), .CE(n259), .R(n261), .D(n14), .Q(o_kdf_test_key_size_config[8]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[9] ( .CK(clk), .CE(n259), .R(n261), .D(n15), .Q(o_kdf_test_key_size_config[9]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[10] ( .CK(clk), .CE(n259), .R(n261), .D(n16), .Q(o_kdf_test_key_size_config[10]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[11] ( .CK(clk), .CE(n259), .R(n261), .D(n17), .Q(o_kdf_test_key_size_config[11]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[12] ( .CK(clk), .CE(n259), .R(n261), .D(n18), .Q(o_kdf_test_key_size_config[12]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[13] ( .CK(clk), .CE(n259), .R(n261), .D(n19), .Q(o_kdf_test_key_size_config[13]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[14] ( .CK(clk), .CE(n259), .R(n261), .D(n20), .Q(o_kdf_test_key_size_config[14]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[15] ( .CK(clk), .CE(n259), .R(n261), .D(n21), .Q(o_kdf_test_key_size_config[15]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[16] ( .CK(clk), .CE(n259), .R(n261), .D(n22), .Q(o_kdf_test_key_size_config[16]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[17] ( .CK(clk), .CE(n259), .R(n261), .D(n23), .Q(o_kdf_test_key_size_config[17]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[18] ( .CK(clk), .CE(n259), .R(n261), .D(n24), .Q(o_kdf_test_key_size_config[18]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[19] ( .CK(clk), .CE(n259), .R(n261), .D(n25), .Q(o_kdf_test_key_size_config[19]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[20] ( .CK(clk), .CE(n259), .R(n261), .D(n26), .Q(o_kdf_test_key_size_config[20]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[21] ( .CK(clk), .CE(n259), .R(n261), .D(n27), .Q(o_kdf_test_key_size_config[21]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[22] ( .CK(clk), .CE(n259), .R(n261), .D(n28), .Q(o_kdf_test_key_size_config[22]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[23] ( .CK(clk), .CE(n259), .R(n261), .D(n29), .Q(o_kdf_test_key_size_config[23]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[24] ( .CK(clk), .CE(n259), .R(n261), .D(n30), .Q(o_kdf_test_key_size_config[24]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[25] ( .CK(clk), .CE(n259), .R(n261), .D(n31), .Q(o_kdf_test_key_size_config[25]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[26] ( .CK(clk), .CE(n259), .R(n261), .D(n32), .Q(o_kdf_test_key_size_config[26]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[27] ( .CK(clk), .CE(n259), .R(n261), .D(n33), .Q(o_kdf_test_key_size_config[27]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[28] ( .CK(clk), .CE(n259), .R(n261), .D(n34), .Q(o_kdf_test_key_size_config[28]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[29] ( .CK(clk), .CE(n259), .R(n261), .D(n35), .Q(o_kdf_test_key_size_config[29]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[30] ( .CK(clk), .CE(n259), .R(n261), .D(n36), .Q(o_kdf_test_key_size_config[30]));
Q_FDP4EP \o_kdf_test_key_size_config_REG[31] ( .CK(clk), .CE(n259), .R(n261), .D(n37), .Q(o_kdf_test_key_size_config[31]));
Q_FDP4EP \o_sa_ctrl_ia_config_REG[0] ( .CK(clk), .CE(n258), .R(n261), .D(n6), .Q(o_sa_ctrl_ia_config[0]));
Q_FDP4EP \o_sa_ctrl_ia_config_REG[1] ( .CK(clk), .CE(n258), .R(n261), .D(n7), .Q(o_sa_ctrl_ia_config[1]));
Q_FDP4EP \o_sa_ctrl_ia_config_REG[2] ( .CK(clk), .CE(n258), .R(n261), .D(n8), .Q(o_sa_ctrl_ia_config[2]));
Q_FDP4EP \o_sa_ctrl_ia_config_REG[3] ( .CK(clk), .CE(n258), .R(n261), .D(n9), .Q(o_sa_ctrl_ia_config[3]));
Q_FDP4EP \o_sa_ctrl_ia_config_REG[4] ( .CK(clk), .CE(n258), .R(n261), .D(n10), .Q(o_sa_ctrl_ia_config[4]));
Q_FDP4EP \o_sa_ctrl_ia_config_REG[5] ( .CK(clk), .CE(n258), .R(n261), .D(n34), .Q(o_sa_ctrl_ia_config[5]));
Q_FDP4EP \o_sa_ctrl_ia_config_REG[6] ( .CK(clk), .CE(n258), .R(n261), .D(n35), .Q(o_sa_ctrl_ia_config[6]));
Q_FDP4EP \o_sa_ctrl_ia_config_REG[7] ( .CK(clk), .CE(n258), .R(n261), .D(n36), .Q(o_sa_ctrl_ia_config[7]));
Q_FDP4EP \o_sa_ctrl_ia_config_REG[8] ( .CK(clk), .CE(n258), .R(n261), .D(n37), .Q(o_sa_ctrl_ia_config[8]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[0] ( .CK(clk), .CE(n257), .R(n261), .D(n6), .Q(o_sa_ctrl_ia_wdata_part0[0]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[1] ( .CK(clk), .CE(n257), .R(n261), .D(n7), .Q(o_sa_ctrl_ia_wdata_part0[1]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[2] ( .CK(clk), .CE(n257), .R(n261), .D(n8), .Q(o_sa_ctrl_ia_wdata_part0[2]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[3] ( .CK(clk), .CE(n257), .R(n261), .D(n9), .Q(o_sa_ctrl_ia_wdata_part0[3]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[4] ( .CK(clk), .CE(n257), .R(n261), .D(n10), .Q(o_sa_ctrl_ia_wdata_part0[4]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[5] ( .CK(clk), .CE(n257), .R(n261), .D(n11), .Q(o_sa_ctrl_ia_wdata_part0[5]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[6] ( .CK(clk), .CE(n257), .R(n261), .D(n12), .Q(o_sa_ctrl_ia_wdata_part0[6]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[7] ( .CK(clk), .CE(n257), .R(n261), .D(n13), .Q(o_sa_ctrl_ia_wdata_part0[7]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[8] ( .CK(clk), .CE(n257), .R(n261), .D(n14), .Q(o_sa_ctrl_ia_wdata_part0[8]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[9] ( .CK(clk), .CE(n257), .R(n261), .D(n15), .Q(o_sa_ctrl_ia_wdata_part0[9]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[10] ( .CK(clk), .CE(n257), .R(n261), .D(n16), .Q(o_sa_ctrl_ia_wdata_part0[10]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[11] ( .CK(clk), .CE(n257), .R(n261), .D(n17), .Q(o_sa_ctrl_ia_wdata_part0[11]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[12] ( .CK(clk), .CE(n257), .R(n261), .D(n18), .Q(o_sa_ctrl_ia_wdata_part0[12]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[13] ( .CK(clk), .CE(n257), .R(n261), .D(n19), .Q(o_sa_ctrl_ia_wdata_part0[13]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[14] ( .CK(clk), .CE(n257), .R(n261), .D(n20), .Q(o_sa_ctrl_ia_wdata_part0[14]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[15] ( .CK(clk), .CE(n257), .R(n261), .D(n21), .Q(o_sa_ctrl_ia_wdata_part0[15]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[16] ( .CK(clk), .CE(n257), .R(n261), .D(n22), .Q(o_sa_ctrl_ia_wdata_part0[16]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[17] ( .CK(clk), .CE(n257), .R(n261), .D(n23), .Q(o_sa_ctrl_ia_wdata_part0[17]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[18] ( .CK(clk), .CE(n257), .R(n261), .D(n24), .Q(o_sa_ctrl_ia_wdata_part0[18]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[19] ( .CK(clk), .CE(n257), .R(n261), .D(n25), .Q(o_sa_ctrl_ia_wdata_part0[19]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[20] ( .CK(clk), .CE(n257), .R(n261), .D(n26), .Q(o_sa_ctrl_ia_wdata_part0[20]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[21] ( .CK(clk), .CE(n257), .R(n261), .D(n27), .Q(o_sa_ctrl_ia_wdata_part0[21]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[22] ( .CK(clk), .CE(n257), .R(n261), .D(n28), .Q(o_sa_ctrl_ia_wdata_part0[22]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[23] ( .CK(clk), .CE(n257), .R(n261), .D(n29), .Q(o_sa_ctrl_ia_wdata_part0[23]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[24] ( .CK(clk), .CE(n257), .R(n261), .D(n30), .Q(o_sa_ctrl_ia_wdata_part0[24]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[25] ( .CK(clk), .CE(n257), .R(n261), .D(n31), .Q(o_sa_ctrl_ia_wdata_part0[25]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[26] ( .CK(clk), .CE(n257), .R(n261), .D(n32), .Q(o_sa_ctrl_ia_wdata_part0[26]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[27] ( .CK(clk), .CE(n257), .R(n261), .D(n33), .Q(o_sa_ctrl_ia_wdata_part0[27]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[28] ( .CK(clk), .CE(n257), .R(n261), .D(n34), .Q(o_sa_ctrl_ia_wdata_part0[28]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[29] ( .CK(clk), .CE(n257), .R(n261), .D(n35), .Q(o_sa_ctrl_ia_wdata_part0[29]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[30] ( .CK(clk), .CE(n257), .R(n261), .D(n36), .Q(o_sa_ctrl_ia_wdata_part0[30]));
Q_FDP4EP \o_sa_ctrl_ia_wdata_part0_REG[31] ( .CK(clk), .CE(n257), .R(n261), .D(n37), .Q(o_sa_ctrl_ia_wdata_part0[31]));
Q_FDP4EP \o_sa_global_ctrl_REG[0] ( .CK(clk), .CE(n256), .R(n261), .D(n6), .Q(o_sa_global_ctrl[0]));
Q_FDP4EP \o_sa_global_ctrl_REG[1] ( .CK(clk), .CE(n256), .R(n261), .D(n7), .Q(o_sa_global_ctrl[1]));
Q_FDP4EP \o_sa_global_ctrl_REG[2] ( .CK(clk), .CE(n256), .R(n261), .D(n8), .Q(o_sa_global_ctrl[2]));
Q_FDP4EP \o_sa_global_ctrl_REG[3] ( .CK(clk), .CE(n256), .R(n261), .D(n9), .Q(o_sa_global_ctrl[3]));
Q_FDP4EP \o_sa_global_ctrl_REG[4] ( .CK(clk), .CE(n256), .R(n261), .D(n10), .Q(o_sa_global_ctrl[4]));
Q_FDP4EP \o_sa_global_ctrl_REG[5] ( .CK(clk), .CE(n256), .R(n261), .D(n11), .Q(o_sa_global_ctrl[5]));
Q_FDP4EP \o_sa_global_ctrl_REG[6] ( .CK(clk), .CE(n256), .R(n261), .D(n12), .Q(o_sa_global_ctrl[6]));
Q_FDP4EP \o_sa_global_ctrl_REG[7] ( .CK(clk), .CE(n256), .R(n261), .D(n13), .Q(o_sa_global_ctrl[7]));
Q_FDP4EP \o_sa_global_ctrl_REG[8] ( .CK(clk), .CE(n256), .R(n261), .D(n14), .Q(o_sa_global_ctrl[8]));
Q_FDP4EP \o_sa_global_ctrl_REG[9] ( .CK(clk), .CE(n256), .R(n261), .D(n15), .Q(o_sa_global_ctrl[9]));
Q_FDP4EP \o_sa_global_ctrl_REG[10] ( .CK(clk), .CE(n256), .R(n261), .D(n16), .Q(o_sa_global_ctrl[10]));
Q_FDP4EP \o_sa_global_ctrl_REG[11] ( .CK(clk), .CE(n256), .R(n261), .D(n17), .Q(o_sa_global_ctrl[11]));
Q_FDP4EP \o_sa_global_ctrl_REG[12] ( .CK(clk), .CE(n256), .R(n261), .D(n18), .Q(o_sa_global_ctrl[12]));
Q_FDP4EP \o_sa_global_ctrl_REG[13] ( .CK(clk), .CE(n256), .R(n261), .D(n19), .Q(o_sa_global_ctrl[13]));
Q_FDP4EP \o_sa_global_ctrl_REG[14] ( .CK(clk), .CE(n256), .R(n261), .D(n20), .Q(o_sa_global_ctrl[14]));
Q_FDP4EP \o_sa_global_ctrl_REG[15] ( .CK(clk), .CE(n256), .R(n261), .D(n21), .Q(o_sa_global_ctrl[15]));
Q_FDP4EP \o_sa_global_ctrl_REG[16] ( .CK(clk), .CE(n256), .R(n261), .D(n22), .Q(o_sa_global_ctrl[16]));
Q_FDP4EP \o_sa_global_ctrl_REG[17] ( .CK(clk), .CE(n256), .R(n261), .D(n23), .Q(o_sa_global_ctrl[17]));
Q_FDP4EP \o_sa_global_ctrl_REG[18] ( .CK(clk), .CE(n256), .R(n261), .D(n24), .Q(o_sa_global_ctrl[18]));
Q_FDP4EP \o_sa_global_ctrl_REG[19] ( .CK(clk), .CE(n256), .R(n261), .D(n25), .Q(o_sa_global_ctrl[19]));
Q_FDP4EP \o_sa_global_ctrl_REG[20] ( .CK(clk), .CE(n256), .R(n261), .D(n26), .Q(o_sa_global_ctrl[20]));
Q_FDP4EP \o_sa_global_ctrl_REG[21] ( .CK(clk), .CE(n256), .R(n261), .D(n27), .Q(o_sa_global_ctrl[21]));
Q_FDP4EP \o_sa_global_ctrl_REG[22] ( .CK(clk), .CE(n256), .R(n261), .D(n28), .Q(o_sa_global_ctrl[22]));
Q_FDP4EP \o_sa_global_ctrl_REG[23] ( .CK(clk), .CE(n256), .R(n261), .D(n29), .Q(o_sa_global_ctrl[23]));
Q_FDP4EP \o_sa_global_ctrl_REG[24] ( .CK(clk), .CE(n256), .R(n261), .D(n30), .Q(o_sa_global_ctrl[24]));
Q_FDP4EP \o_sa_global_ctrl_REG[25] ( .CK(clk), .CE(n256), .R(n261), .D(n31), .Q(o_sa_global_ctrl[25]));
Q_FDP4EP \o_sa_global_ctrl_REG[26] ( .CK(clk), .CE(n256), .R(n261), .D(n32), .Q(o_sa_global_ctrl[26]));
Q_FDP4EP \o_sa_global_ctrl_REG[27] ( .CK(clk), .CE(n256), .R(n261), .D(n33), .Q(o_sa_global_ctrl[27]));
Q_FDP4EP \o_sa_global_ctrl_REG[28] ( .CK(clk), .CE(n256), .R(n261), .D(n34), .Q(o_sa_global_ctrl[28]));
Q_FDP4EP \o_sa_global_ctrl_REG[29] ( .CK(clk), .CE(n256), .R(n261), .D(n35), .Q(o_sa_global_ctrl[29]));
Q_FDP4EP \o_sa_global_ctrl_REG[30] ( .CK(clk), .CE(n256), .R(n261), .D(n36), .Q(o_sa_global_ctrl[30]));
Q_FDP4EP \o_sa_global_ctrl_REG[31] ( .CK(clk), .CE(n256), .R(n261), .D(n37), .Q(o_sa_global_ctrl[31]));
Q_FDP4EP \o_cddip_decrypt_kop_fifo_override_REG[0] ( .CK(clk), .CE(n255), .R(n261), .D(n6), .Q(o_cddip_decrypt_kop_fifo_override[0]));
Q_FDP4EP \o_cddip_decrypt_kop_fifo_override_REG[1] ( .CK(clk), .CE(n255), .R(n261), .D(n7), .Q(o_cddip_decrypt_kop_fifo_override[1]));
Q_FDP4EP \o_cddip_decrypt_kop_fifo_override_REG[2] ( .CK(clk), .CE(n255), .R(n261), .D(n8), .Q(o_cddip_decrypt_kop_fifo_override[2]));
Q_FDP4EP \o_cddip_decrypt_kop_fifo_override_REG[3] ( .CK(clk), .CE(n255), .R(n261), .D(n9), .Q(o_cddip_decrypt_kop_fifo_override[3]));
Q_FDP4EP \o_cddip_decrypt_kop_fifo_override_REG[4] ( .CK(clk), .CE(n255), .R(n261), .D(n10), .Q(o_cddip_decrypt_kop_fifo_override[4]));
Q_FDP4EP \o_cddip_decrypt_kop_fifo_override_REG[5] ( .CK(clk), .CE(n255), .R(n261), .D(n11), .Q(o_cddip_decrypt_kop_fifo_override[5]));
Q_FDP4EP \o_cddip_decrypt_kop_fifo_override_REG[6] ( .CK(clk), .CE(n255), .R(n261), .D(n12), .Q(o_cddip_decrypt_kop_fifo_override[6]));
Q_FDP4EP \o_cceip_validate_kop_fifo_override_REG[0] ( .CK(clk), .CE(n254), .R(n261), .D(n6), .Q(o_cceip_validate_kop_fifo_override[0]));
Q_FDP4EP \o_cceip_validate_kop_fifo_override_REG[1] ( .CK(clk), .CE(n254), .R(n261), .D(n7), .Q(o_cceip_validate_kop_fifo_override[1]));
Q_FDP4EP \o_cceip_validate_kop_fifo_override_REG[2] ( .CK(clk), .CE(n254), .R(n261), .D(n8), .Q(o_cceip_validate_kop_fifo_override[2]));
Q_FDP4EP \o_cceip_validate_kop_fifo_override_REG[3] ( .CK(clk), .CE(n254), .R(n261), .D(n9), .Q(o_cceip_validate_kop_fifo_override[3]));
Q_FDP4EP \o_cceip_validate_kop_fifo_override_REG[4] ( .CK(clk), .CE(n254), .R(n261), .D(n10), .Q(o_cceip_validate_kop_fifo_override[4]));
Q_FDP4EP \o_cceip_validate_kop_fifo_override_REG[5] ( .CK(clk), .CE(n254), .R(n261), .D(n11), .Q(o_cceip_validate_kop_fifo_override[5]));
Q_FDP4EP \o_cceip_validate_kop_fifo_override_REG[6] ( .CK(clk), .CE(n254), .R(n261), .D(n12), .Q(o_cceip_validate_kop_fifo_override[6]));
Q_FDP4EP \o_cceip_encrypt_kop_fifo_override_REG[0] ( .CK(clk), .CE(n253), .R(n261), .D(n6), .Q(o_cceip_encrypt_kop_fifo_override[0]));
Q_FDP4EP \o_cceip_encrypt_kop_fifo_override_REG[1] ( .CK(clk), .CE(n253), .R(n261), .D(n7), .Q(o_cceip_encrypt_kop_fifo_override[1]));
Q_FDP4EP \o_cceip_encrypt_kop_fifo_override_REG[2] ( .CK(clk), .CE(n253), .R(n261), .D(n8), .Q(o_cceip_encrypt_kop_fifo_override[2]));
Q_FDP4EP \o_cceip_encrypt_kop_fifo_override_REG[3] ( .CK(clk), .CE(n253), .R(n261), .D(n9), .Q(o_cceip_encrypt_kop_fifo_override[3]));
Q_FDP4EP \o_cceip_encrypt_kop_fifo_override_REG[4] ( .CK(clk), .CE(n253), .R(n261), .D(n10), .Q(o_cceip_encrypt_kop_fifo_override[4]));
Q_FDP4EP \o_cceip_encrypt_kop_fifo_override_REG[5] ( .CK(clk), .CE(n253), .R(n261), .D(n11), .Q(o_cceip_encrypt_kop_fifo_override[5]));
Q_FDP4EP \o_cceip_encrypt_kop_fifo_override_REG[6] ( .CK(clk), .CE(n253), .R(n261), .D(n12), .Q(o_cceip_encrypt_kop_fifo_override[6]));
Q_FDP4EP \o_sa_count_ia_config_REG[0] ( .CK(clk), .CE(n252), .R(n261), .D(n6), .Q(o_sa_count_ia_config[0]));
Q_FDP4EP \o_sa_count_ia_config_REG[1] ( .CK(clk), .CE(n252), .R(n261), .D(n7), .Q(o_sa_count_ia_config[1]));
Q_FDP4EP \o_sa_count_ia_config_REG[2] ( .CK(clk), .CE(n252), .R(n261), .D(n8), .Q(o_sa_count_ia_config[2]));
Q_FDP4EP \o_sa_count_ia_config_REG[3] ( .CK(clk), .CE(n252), .R(n261), .D(n9), .Q(o_sa_count_ia_config[3]));
Q_FDP4EP \o_sa_count_ia_config_REG[4] ( .CK(clk), .CE(n252), .R(n261), .D(n10), .Q(o_sa_count_ia_config[4]));
Q_FDP4EP \o_sa_count_ia_config_REG[5] ( .CK(clk), .CE(n252), .R(n261), .D(n34), .Q(o_sa_count_ia_config[5]));
Q_FDP4EP \o_sa_count_ia_config_REG[6] ( .CK(clk), .CE(n252), .R(n261), .D(n35), .Q(o_sa_count_ia_config[6]));
Q_FDP4EP \o_sa_count_ia_config_REG[7] ( .CK(clk), .CE(n252), .R(n261), .D(n36), .Q(o_sa_count_ia_config[7]));
Q_FDP4EP \o_sa_count_ia_config_REG[8] ( .CK(clk), .CE(n252), .R(n261), .D(n37), .Q(o_sa_count_ia_config[8]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[0] ( .CK(clk), .CE(n251), .R(n261), .D(n6), .Q(o_sa_count_ia_wdata_part1[0]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[1] ( .CK(clk), .CE(n251), .R(n261), .D(n7), .Q(o_sa_count_ia_wdata_part1[1]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[2] ( .CK(clk), .CE(n251), .R(n261), .D(n8), .Q(o_sa_count_ia_wdata_part1[2]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[3] ( .CK(clk), .CE(n251), .R(n261), .D(n9), .Q(o_sa_count_ia_wdata_part1[3]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[4] ( .CK(clk), .CE(n251), .R(n261), .D(n10), .Q(o_sa_count_ia_wdata_part1[4]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[5] ( .CK(clk), .CE(n251), .R(n261), .D(n11), .Q(o_sa_count_ia_wdata_part1[5]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[6] ( .CK(clk), .CE(n251), .R(n261), .D(n12), .Q(o_sa_count_ia_wdata_part1[6]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[7] ( .CK(clk), .CE(n251), .R(n261), .D(n13), .Q(o_sa_count_ia_wdata_part1[7]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[8] ( .CK(clk), .CE(n251), .R(n261), .D(n14), .Q(o_sa_count_ia_wdata_part1[8]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[9] ( .CK(clk), .CE(n251), .R(n261), .D(n15), .Q(o_sa_count_ia_wdata_part1[9]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[10] ( .CK(clk), .CE(n251), .R(n261), .D(n16), .Q(o_sa_count_ia_wdata_part1[10]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[11] ( .CK(clk), .CE(n251), .R(n261), .D(n17), .Q(o_sa_count_ia_wdata_part1[11]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[12] ( .CK(clk), .CE(n251), .R(n261), .D(n18), .Q(o_sa_count_ia_wdata_part1[12]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[13] ( .CK(clk), .CE(n251), .R(n261), .D(n19), .Q(o_sa_count_ia_wdata_part1[13]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[14] ( .CK(clk), .CE(n251), .R(n261), .D(n20), .Q(o_sa_count_ia_wdata_part1[14]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[15] ( .CK(clk), .CE(n251), .R(n261), .D(n21), .Q(o_sa_count_ia_wdata_part1[15]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[16] ( .CK(clk), .CE(n251), .R(n261), .D(n22), .Q(o_sa_count_ia_wdata_part1[16]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[17] ( .CK(clk), .CE(n251), .R(n261), .D(n23), .Q(o_sa_count_ia_wdata_part1[17]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[18] ( .CK(clk), .CE(n251), .R(n261), .D(n24), .Q(o_sa_count_ia_wdata_part1[18]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[19] ( .CK(clk), .CE(n251), .R(n261), .D(n25), .Q(o_sa_count_ia_wdata_part1[19]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[20] ( .CK(clk), .CE(n251), .R(n261), .D(n26), .Q(o_sa_count_ia_wdata_part1[20]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[21] ( .CK(clk), .CE(n251), .R(n261), .D(n27), .Q(o_sa_count_ia_wdata_part1[21]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[22] ( .CK(clk), .CE(n251), .R(n261), .D(n28), .Q(o_sa_count_ia_wdata_part1[22]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[23] ( .CK(clk), .CE(n251), .R(n261), .D(n29), .Q(o_sa_count_ia_wdata_part1[23]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[24] ( .CK(clk), .CE(n251), .R(n261), .D(n30), .Q(o_sa_count_ia_wdata_part1[24]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[25] ( .CK(clk), .CE(n251), .R(n261), .D(n31), .Q(o_sa_count_ia_wdata_part1[25]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[26] ( .CK(clk), .CE(n251), .R(n261), .D(n32), .Q(o_sa_count_ia_wdata_part1[26]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[27] ( .CK(clk), .CE(n251), .R(n261), .D(n33), .Q(o_sa_count_ia_wdata_part1[27]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[28] ( .CK(clk), .CE(n251), .R(n261), .D(n34), .Q(o_sa_count_ia_wdata_part1[28]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[29] ( .CK(clk), .CE(n251), .R(n261), .D(n35), .Q(o_sa_count_ia_wdata_part1[29]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[30] ( .CK(clk), .CE(n251), .R(n261), .D(n36), .Q(o_sa_count_ia_wdata_part1[30]));
Q_FDP4EP \o_sa_count_ia_wdata_part1_REG[31] ( .CK(clk), .CE(n251), .R(n261), .D(n37), .Q(o_sa_count_ia_wdata_part1[31]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[0] ( .CK(clk), .CE(n250), .R(n261), .D(n6), .Q(o_sa_count_ia_wdata_part0[0]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[1] ( .CK(clk), .CE(n250), .R(n261), .D(n7), .Q(o_sa_count_ia_wdata_part0[1]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[2] ( .CK(clk), .CE(n250), .R(n261), .D(n8), .Q(o_sa_count_ia_wdata_part0[2]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[3] ( .CK(clk), .CE(n250), .R(n261), .D(n9), .Q(o_sa_count_ia_wdata_part0[3]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[4] ( .CK(clk), .CE(n250), .R(n261), .D(n10), .Q(o_sa_count_ia_wdata_part0[4]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[5] ( .CK(clk), .CE(n250), .R(n261), .D(n11), .Q(o_sa_count_ia_wdata_part0[5]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[6] ( .CK(clk), .CE(n250), .R(n261), .D(n12), .Q(o_sa_count_ia_wdata_part0[6]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[7] ( .CK(clk), .CE(n250), .R(n261), .D(n13), .Q(o_sa_count_ia_wdata_part0[7]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[8] ( .CK(clk), .CE(n250), .R(n261), .D(n14), .Q(o_sa_count_ia_wdata_part0[8]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[9] ( .CK(clk), .CE(n250), .R(n261), .D(n15), .Q(o_sa_count_ia_wdata_part0[9]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[10] ( .CK(clk), .CE(n250), .R(n261), .D(n16), .Q(o_sa_count_ia_wdata_part0[10]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[11] ( .CK(clk), .CE(n250), .R(n261), .D(n17), .Q(o_sa_count_ia_wdata_part0[11]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[12] ( .CK(clk), .CE(n250), .R(n261), .D(n18), .Q(o_sa_count_ia_wdata_part0[12]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[13] ( .CK(clk), .CE(n250), .R(n261), .D(n19), .Q(o_sa_count_ia_wdata_part0[13]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[14] ( .CK(clk), .CE(n250), .R(n261), .D(n20), .Q(o_sa_count_ia_wdata_part0[14]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[15] ( .CK(clk), .CE(n250), .R(n261), .D(n21), .Q(o_sa_count_ia_wdata_part0[15]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[16] ( .CK(clk), .CE(n250), .R(n261), .D(n22), .Q(o_sa_count_ia_wdata_part0[16]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[17] ( .CK(clk), .CE(n250), .R(n261), .D(n23), .Q(o_sa_count_ia_wdata_part0[17]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[18] ( .CK(clk), .CE(n250), .R(n261), .D(n24), .Q(o_sa_count_ia_wdata_part0[18]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[19] ( .CK(clk), .CE(n250), .R(n261), .D(n25), .Q(o_sa_count_ia_wdata_part0[19]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[20] ( .CK(clk), .CE(n250), .R(n261), .D(n26), .Q(o_sa_count_ia_wdata_part0[20]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[21] ( .CK(clk), .CE(n250), .R(n261), .D(n27), .Q(o_sa_count_ia_wdata_part0[21]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[22] ( .CK(clk), .CE(n250), .R(n261), .D(n28), .Q(o_sa_count_ia_wdata_part0[22]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[23] ( .CK(clk), .CE(n250), .R(n261), .D(n29), .Q(o_sa_count_ia_wdata_part0[23]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[24] ( .CK(clk), .CE(n250), .R(n261), .D(n30), .Q(o_sa_count_ia_wdata_part0[24]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[25] ( .CK(clk), .CE(n250), .R(n261), .D(n31), .Q(o_sa_count_ia_wdata_part0[25]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[26] ( .CK(clk), .CE(n250), .R(n261), .D(n32), .Q(o_sa_count_ia_wdata_part0[26]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[27] ( .CK(clk), .CE(n250), .R(n261), .D(n33), .Q(o_sa_count_ia_wdata_part0[27]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[28] ( .CK(clk), .CE(n250), .R(n261), .D(n34), .Q(o_sa_count_ia_wdata_part0[28]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[29] ( .CK(clk), .CE(n250), .R(n261), .D(n35), .Q(o_sa_count_ia_wdata_part0[29]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[30] ( .CK(clk), .CE(n250), .R(n261), .D(n36), .Q(o_sa_count_ia_wdata_part0[30]));
Q_FDP4EP \o_sa_count_ia_wdata_part0_REG[31] ( .CK(clk), .CE(n250), .R(n261), .D(n37), .Q(o_sa_count_ia_wdata_part0[31]));
Q_FDP4EP \o_sa_snapshot_ia_config_REG[0] ( .CK(clk), .CE(n249), .R(n261), .D(n6), .Q(o_sa_snapshot_ia_config[0]));
Q_FDP4EP \o_sa_snapshot_ia_config_REG[1] ( .CK(clk), .CE(n249), .R(n261), .D(n7), .Q(o_sa_snapshot_ia_config[1]));
Q_FDP4EP \o_sa_snapshot_ia_config_REG[2] ( .CK(clk), .CE(n249), .R(n261), .D(n8), .Q(o_sa_snapshot_ia_config[2]));
Q_FDP4EP \o_sa_snapshot_ia_config_REG[3] ( .CK(clk), .CE(n249), .R(n261), .D(n9), .Q(o_sa_snapshot_ia_config[3]));
Q_FDP4EP \o_sa_snapshot_ia_config_REG[4] ( .CK(clk), .CE(n249), .R(n261), .D(n10), .Q(o_sa_snapshot_ia_config[4]));
Q_FDP4EP \o_sa_snapshot_ia_config_REG[5] ( .CK(clk), .CE(n249), .R(n261), .D(n34), .Q(o_sa_snapshot_ia_config[5]));
Q_FDP4EP \o_sa_snapshot_ia_config_REG[6] ( .CK(clk), .CE(n249), .R(n261), .D(n35), .Q(o_sa_snapshot_ia_config[6]));
Q_FDP4EP \o_sa_snapshot_ia_config_REG[7] ( .CK(clk), .CE(n249), .R(n261), .D(n36), .Q(o_sa_snapshot_ia_config[7]));
Q_FDP4EP \o_sa_snapshot_ia_config_REG[8] ( .CK(clk), .CE(n249), .R(n261), .D(n37), .Q(o_sa_snapshot_ia_config[8]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[0] ( .CK(clk), .CE(n248), .R(n261), .D(n6), .Q(o_sa_snapshot_ia_wdata_part1[0]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[1] ( .CK(clk), .CE(n248), .R(n261), .D(n7), .Q(o_sa_snapshot_ia_wdata_part1[1]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[2] ( .CK(clk), .CE(n248), .R(n261), .D(n8), .Q(o_sa_snapshot_ia_wdata_part1[2]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[3] ( .CK(clk), .CE(n248), .R(n261), .D(n9), .Q(o_sa_snapshot_ia_wdata_part1[3]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[4] ( .CK(clk), .CE(n248), .R(n261), .D(n10), .Q(o_sa_snapshot_ia_wdata_part1[4]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[5] ( .CK(clk), .CE(n248), .R(n261), .D(n11), .Q(o_sa_snapshot_ia_wdata_part1[5]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[6] ( .CK(clk), .CE(n248), .R(n261), .D(n12), .Q(o_sa_snapshot_ia_wdata_part1[6]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[7] ( .CK(clk), .CE(n248), .R(n261), .D(n13), .Q(o_sa_snapshot_ia_wdata_part1[7]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[8] ( .CK(clk), .CE(n248), .R(n261), .D(n14), .Q(o_sa_snapshot_ia_wdata_part1[8]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[9] ( .CK(clk), .CE(n248), .R(n261), .D(n15), .Q(o_sa_snapshot_ia_wdata_part1[9]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[10] ( .CK(clk), .CE(n248), .R(n261), .D(n16), .Q(o_sa_snapshot_ia_wdata_part1[10]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[11] ( .CK(clk), .CE(n248), .R(n261), .D(n17), .Q(o_sa_snapshot_ia_wdata_part1[11]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[12] ( .CK(clk), .CE(n248), .R(n261), .D(n18), .Q(o_sa_snapshot_ia_wdata_part1[12]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[13] ( .CK(clk), .CE(n248), .R(n261), .D(n19), .Q(o_sa_snapshot_ia_wdata_part1[13]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[14] ( .CK(clk), .CE(n248), .R(n261), .D(n20), .Q(o_sa_snapshot_ia_wdata_part1[14]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[15] ( .CK(clk), .CE(n248), .R(n261), .D(n21), .Q(o_sa_snapshot_ia_wdata_part1[15]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[16] ( .CK(clk), .CE(n248), .R(n261), .D(n22), .Q(o_sa_snapshot_ia_wdata_part1[16]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[17] ( .CK(clk), .CE(n248), .R(n261), .D(n23), .Q(o_sa_snapshot_ia_wdata_part1[17]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[18] ( .CK(clk), .CE(n248), .R(n261), .D(n24), .Q(o_sa_snapshot_ia_wdata_part1[18]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[19] ( .CK(clk), .CE(n248), .R(n261), .D(n25), .Q(o_sa_snapshot_ia_wdata_part1[19]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[20] ( .CK(clk), .CE(n248), .R(n261), .D(n26), .Q(o_sa_snapshot_ia_wdata_part1[20]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[21] ( .CK(clk), .CE(n248), .R(n261), .D(n27), .Q(o_sa_snapshot_ia_wdata_part1[21]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[22] ( .CK(clk), .CE(n248), .R(n261), .D(n28), .Q(o_sa_snapshot_ia_wdata_part1[22]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[23] ( .CK(clk), .CE(n248), .R(n261), .D(n29), .Q(o_sa_snapshot_ia_wdata_part1[23]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[24] ( .CK(clk), .CE(n248), .R(n261), .D(n30), .Q(o_sa_snapshot_ia_wdata_part1[24]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[25] ( .CK(clk), .CE(n248), .R(n261), .D(n31), .Q(o_sa_snapshot_ia_wdata_part1[25]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[26] ( .CK(clk), .CE(n248), .R(n261), .D(n32), .Q(o_sa_snapshot_ia_wdata_part1[26]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[27] ( .CK(clk), .CE(n248), .R(n261), .D(n33), .Q(o_sa_snapshot_ia_wdata_part1[27]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[28] ( .CK(clk), .CE(n248), .R(n261), .D(n34), .Q(o_sa_snapshot_ia_wdata_part1[28]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[29] ( .CK(clk), .CE(n248), .R(n261), .D(n35), .Q(o_sa_snapshot_ia_wdata_part1[29]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[30] ( .CK(clk), .CE(n248), .R(n261), .D(n36), .Q(o_sa_snapshot_ia_wdata_part1[30]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part1_REG[31] ( .CK(clk), .CE(n248), .R(n261), .D(n37), .Q(o_sa_snapshot_ia_wdata_part1[31]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[0] ( .CK(clk), .CE(n247), .R(n261), .D(n6), .Q(o_sa_snapshot_ia_wdata_part0[0]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[1] ( .CK(clk), .CE(n247), .R(n261), .D(n7), .Q(o_sa_snapshot_ia_wdata_part0[1]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[2] ( .CK(clk), .CE(n247), .R(n261), .D(n8), .Q(o_sa_snapshot_ia_wdata_part0[2]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[3] ( .CK(clk), .CE(n247), .R(n261), .D(n9), .Q(o_sa_snapshot_ia_wdata_part0[3]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[4] ( .CK(clk), .CE(n247), .R(n261), .D(n10), .Q(o_sa_snapshot_ia_wdata_part0[4]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[5] ( .CK(clk), .CE(n247), .R(n261), .D(n11), .Q(o_sa_snapshot_ia_wdata_part0[5]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[6] ( .CK(clk), .CE(n247), .R(n261), .D(n12), .Q(o_sa_snapshot_ia_wdata_part0[6]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[7] ( .CK(clk), .CE(n247), .R(n261), .D(n13), .Q(o_sa_snapshot_ia_wdata_part0[7]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[8] ( .CK(clk), .CE(n247), .R(n261), .D(n14), .Q(o_sa_snapshot_ia_wdata_part0[8]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[9] ( .CK(clk), .CE(n247), .R(n261), .D(n15), .Q(o_sa_snapshot_ia_wdata_part0[9]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[10] ( .CK(clk), .CE(n247), .R(n261), .D(n16), .Q(o_sa_snapshot_ia_wdata_part0[10]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[11] ( .CK(clk), .CE(n247), .R(n261), .D(n17), .Q(o_sa_snapshot_ia_wdata_part0[11]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[12] ( .CK(clk), .CE(n247), .R(n261), .D(n18), .Q(o_sa_snapshot_ia_wdata_part0[12]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[13] ( .CK(clk), .CE(n247), .R(n261), .D(n19), .Q(o_sa_snapshot_ia_wdata_part0[13]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[14] ( .CK(clk), .CE(n247), .R(n261), .D(n20), .Q(o_sa_snapshot_ia_wdata_part0[14]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[15] ( .CK(clk), .CE(n247), .R(n261), .D(n21), .Q(o_sa_snapshot_ia_wdata_part0[15]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[16] ( .CK(clk), .CE(n247), .R(n261), .D(n22), .Q(o_sa_snapshot_ia_wdata_part0[16]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[17] ( .CK(clk), .CE(n247), .R(n261), .D(n23), .Q(o_sa_snapshot_ia_wdata_part0[17]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[18] ( .CK(clk), .CE(n247), .R(n261), .D(n24), .Q(o_sa_snapshot_ia_wdata_part0[18]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[19] ( .CK(clk), .CE(n247), .R(n261), .D(n25), .Q(o_sa_snapshot_ia_wdata_part0[19]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[20] ( .CK(clk), .CE(n247), .R(n261), .D(n26), .Q(o_sa_snapshot_ia_wdata_part0[20]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[21] ( .CK(clk), .CE(n247), .R(n261), .D(n27), .Q(o_sa_snapshot_ia_wdata_part0[21]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[22] ( .CK(clk), .CE(n247), .R(n261), .D(n28), .Q(o_sa_snapshot_ia_wdata_part0[22]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[23] ( .CK(clk), .CE(n247), .R(n261), .D(n29), .Q(o_sa_snapshot_ia_wdata_part0[23]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[24] ( .CK(clk), .CE(n247), .R(n261), .D(n30), .Q(o_sa_snapshot_ia_wdata_part0[24]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[25] ( .CK(clk), .CE(n247), .R(n261), .D(n31), .Q(o_sa_snapshot_ia_wdata_part0[25]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[26] ( .CK(clk), .CE(n247), .R(n261), .D(n32), .Q(o_sa_snapshot_ia_wdata_part0[26]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[27] ( .CK(clk), .CE(n247), .R(n261), .D(n33), .Q(o_sa_snapshot_ia_wdata_part0[27]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[28] ( .CK(clk), .CE(n247), .R(n261), .D(n34), .Q(o_sa_snapshot_ia_wdata_part0[28]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[29] ( .CK(clk), .CE(n247), .R(n261), .D(n35), .Q(o_sa_snapshot_ia_wdata_part0[29]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[30] ( .CK(clk), .CE(n247), .R(n261), .D(n36), .Q(o_sa_snapshot_ia_wdata_part0[30]));
Q_FDP4EP \o_sa_snapshot_ia_wdata_part0_REG[31] ( .CK(clk), .CE(n247), .R(n261), .D(n37), .Q(o_sa_snapshot_ia_wdata_part0[31]));
Q_FDP4EP \o_regs_sa_ctrl_REG[0] ( .CK(clk), .CE(n246), .R(n261), .D(n6), .Q(o_regs_sa_ctrl[0]));
Q_FDP4EP \o_regs_sa_ctrl_REG[1] ( .CK(clk), .CE(n246), .R(n261), .D(n7), .Q(o_regs_sa_ctrl[1]));
Q_FDP4EP \o_regs_sa_ctrl_REG[2] ( .CK(clk), .CE(n246), .R(n261), .D(n8), .Q(o_regs_sa_ctrl[2]));
Q_FDP4EP \o_regs_sa_ctrl_REG[3] ( .CK(clk), .CE(n246), .R(n261), .D(n9), .Q(o_regs_sa_ctrl[3]));
Q_FDP4EP \o_regs_sa_ctrl_REG[4] ( .CK(clk), .CE(n246), .R(n261), .D(n10), .Q(o_regs_sa_ctrl[4]));
Q_FDP4EP \o_regs_sa_ctrl_REG[5] ( .CK(clk), .CE(n246), .R(n261), .D(n11), .Q(o_regs_sa_ctrl[5]));
Q_FDP4EP \o_regs_sa_ctrl_REG[6] ( .CK(clk), .CE(n246), .R(n261), .D(n12), .Q(o_regs_sa_ctrl[6]));
Q_FDP4EP \o_regs_sa_ctrl_REG[7] ( .CK(clk), .CE(n246), .R(n261), .D(n13), .Q(o_regs_sa_ctrl[7]));
Q_FDP4EP \o_regs_sa_ctrl_REG[8] ( .CK(clk), .CE(n246), .R(n261), .D(n14), .Q(o_regs_sa_ctrl[8]));
Q_FDP4EP \o_regs_sa_ctrl_REG[9] ( .CK(clk), .CE(n246), .R(n261), .D(n15), .Q(o_regs_sa_ctrl[9]));
Q_FDP4EP \o_regs_sa_ctrl_REG[10] ( .CK(clk), .CE(n246), .R(n261), .D(n16), .Q(o_regs_sa_ctrl[10]));
Q_FDP4EP \o_regs_sa_ctrl_REG[11] ( .CK(clk), .CE(n246), .R(n261), .D(n17), .Q(o_regs_sa_ctrl[11]));
Q_FDP4EP \o_regs_sa_ctrl_REG[12] ( .CK(clk), .CE(n246), .R(n261), .D(n18), .Q(o_regs_sa_ctrl[12]));
Q_FDP4EP \o_regs_sa_ctrl_REG[13] ( .CK(clk), .CE(n246), .R(n261), .D(n19), .Q(o_regs_sa_ctrl[13]));
Q_FDP4EP \o_regs_sa_ctrl_REG[14] ( .CK(clk), .CE(n246), .R(n261), .D(n20), .Q(o_regs_sa_ctrl[14]));
Q_FDP4EP \o_regs_sa_ctrl_REG[15] ( .CK(clk), .CE(n246), .R(n261), .D(n21), .Q(o_regs_sa_ctrl[15]));
Q_FDP4EP \o_regs_sa_ctrl_REG[16] ( .CK(clk), .CE(n246), .R(n261), .D(n22), .Q(o_regs_sa_ctrl[16]));
Q_FDP4EP \o_regs_sa_ctrl_REG[17] ( .CK(clk), .CE(n246), .R(n261), .D(n23), .Q(o_regs_sa_ctrl[17]));
Q_FDP4EP \o_regs_sa_ctrl_REG[18] ( .CK(clk), .CE(n246), .R(n261), .D(n24), .Q(o_regs_sa_ctrl[18]));
Q_FDP4EP \o_regs_sa_ctrl_REG[19] ( .CK(clk), .CE(n246), .R(n261), .D(n25), .Q(o_regs_sa_ctrl[19]));
Q_FDP4EP \o_regs_sa_ctrl_REG[20] ( .CK(clk), .CE(n246), .R(n261), .D(n26), .Q(o_regs_sa_ctrl[20]));
Q_FDP4EP \o_regs_sa_ctrl_REG[21] ( .CK(clk), .CE(n246), .R(n261), .D(n27), .Q(o_regs_sa_ctrl[21]));
Q_FDP4EP \o_regs_sa_ctrl_REG[22] ( .CK(clk), .CE(n246), .R(n261), .D(n28), .Q(o_regs_sa_ctrl[22]));
Q_FDP4EP \o_regs_sa_ctrl_REG[23] ( .CK(clk), .CE(n246), .R(n261), .D(n29), .Q(o_regs_sa_ctrl[23]));
Q_FDP4EP \o_regs_sa_ctrl_REG[24] ( .CK(clk), .CE(n246), .R(n261), .D(n30), .Q(o_regs_sa_ctrl[24]));
Q_FDP4EP \o_regs_sa_ctrl_REG[25] ( .CK(clk), .CE(n246), .R(n261), .D(n31), .Q(o_regs_sa_ctrl[25]));
Q_FDP4EP \o_regs_sa_ctrl_REG[26] ( .CK(clk), .CE(n246), .R(n261), .D(n32), .Q(o_regs_sa_ctrl[26]));
Q_FDP4EP \o_regs_sa_ctrl_REG[27] ( .CK(clk), .CE(n246), .R(n261), .D(n33), .Q(o_regs_sa_ctrl[27]));
Q_FDP4EP \o_regs_sa_ctrl_REG[28] ( .CK(clk), .CE(n246), .R(n261), .D(n34), .Q(o_regs_sa_ctrl[28]));
Q_FDP4EP \o_regs_sa_ctrl_REG[29] ( .CK(clk), .CE(n246), .R(n261), .D(n35), .Q(o_regs_sa_ctrl[29]));
Q_FDP4EP \o_regs_sa_ctrl_REG[30] ( .CK(clk), .CE(n246), .R(n261), .D(n36), .Q(o_regs_sa_ctrl[30]));
Q_FDP4EP \o_regs_sa_ctrl_REG[31] ( .CK(clk), .CE(n246), .R(n261), .D(n37), .Q(o_regs_sa_ctrl[31]));
Q_FDP4EP \o_tready_override_REG[0] ( .CK(clk), .CE(n245), .R(n261), .D(n6), .Q(o_tready_override[0]));
Q_FDP4EP \o_tready_override_REG[1] ( .CK(clk), .CE(n245), .R(n261), .D(n7), .Q(o_tready_override[1]));
Q_FDP4EP \o_tready_override_REG[2] ( .CK(clk), .CE(n245), .R(n261), .D(n8), .Q(o_tready_override[2]));
Q_FDP4EP \o_tready_override_REG[3] ( .CK(clk), .CE(n245), .R(n261), .D(n9), .Q(o_tready_override[3]));
Q_FDP4EP \o_tready_override_REG[4] ( .CK(clk), .CE(n245), .R(n261), .D(n10), .Q(o_tready_override[4]));
Q_FDP4EP \o_tready_override_REG[5] ( .CK(clk), .CE(n245), .R(n261), .D(n11), .Q(o_tready_override[5]));
Q_FDP4EP \o_tready_override_REG[6] ( .CK(clk), .CE(n245), .R(n261), .D(n12), .Q(o_tready_override[6]));
Q_FDP4EP \o_tready_override_REG[7] ( .CK(clk), .CE(n245), .R(n261), .D(n13), .Q(o_tready_override[7]));
Q_FDP4EP \o_tready_override_REG[8] ( .CK(clk), .CE(n245), .R(n261), .D(n14), .Q(o_tready_override[8]));
Q_FDP4EP \o_im_consumed_REG[0] ( .CK(clk), .CE(n244), .R(n261), .D(n6), .Q(o_im_consumed[0]));
Q_FDP4EP \o_im_consumed_REG[1] ( .CK(clk), .CE(n244), .R(n261), .D(n7), .Q(o_im_consumed[1]));
Q_FDP4EP \o_im_consumed_REG[2] ( .CK(clk), .CE(n244), .R(n261), .D(n8), .Q(o_im_consumed[2]));
Q_FDP4EP \o_im_consumed_REG[3] ( .CK(clk), .CE(n244), .R(n261), .D(n9), .Q(o_im_consumed[3]));
Q_FDP4EP \o_im_consumed_REG[4] ( .CK(clk), .CE(n244), .R(n261), .D(n10), .Q(o_im_consumed[4]));
Q_FDP4EP \o_im_consumed_REG[5] ( .CK(clk), .CE(n244), .R(n261), .D(n11), .Q(o_im_consumed[5]));
Q_FDP4EP \o_im_consumed_REG[6] ( .CK(clk), .CE(n244), .R(n261), .D(n12), .Q(o_im_consumed[6]));
Q_FDP4EP \o_im_consumed_REG[7] ( .CK(clk), .CE(n244), .R(n261), .D(n13), .Q(o_im_consumed[7]));
Q_FDP4EP \o_im_consumed_REG[8] ( .CK(clk), .CE(n244), .R(n261), .D(n14), .Q(o_im_consumed[8]));
Q_FDP4EP \o_im_consumed_REG[9] ( .CK(clk), .CE(n244), .R(n261), .D(n15), .Q(o_im_consumed[9]));
Q_FDP4EP \o_im_consumed_REG[10] ( .CK(clk), .CE(n244), .R(n261), .D(n16), .Q(o_im_consumed[10]));
Q_FDP4EP \o_im_consumed_REG[11] ( .CK(clk), .CE(n244), .R(n261), .D(n17), .Q(o_im_consumed[11]));
Q_FDP4EP \o_im_consumed_REG[12] ( .CK(clk), .CE(n244), .R(n261), .D(n18), .Q(o_im_consumed[12]));
Q_FDP4EP \o_im_consumed_REG[13] ( .CK(clk), .CE(n244), .R(n261), .D(n19), .Q(o_im_consumed[13]));
Q_FDP4EP \o_im_consumed_REG[14] ( .CK(clk), .CE(n244), .R(n261), .D(n20), .Q(o_im_consumed[14]));
Q_FDP4EP \o_im_consumed_REG[15] ( .CK(clk), .CE(n244), .R(n261), .D(n21), .Q(o_im_consumed[15]));
Q_FDP4EP \o_bimc_dbgcmd2_REG[0] ( .CK(clk), .CE(n243), .R(n261), .D(n6), .Q(o_bimc_dbgcmd2[0]));
Q_FDP4EP \o_bimc_dbgcmd2_REG[1] ( .CK(clk), .CE(n243), .R(n261), .D(n7), .Q(o_bimc_dbgcmd2[1]));
Q_FDP4EP \o_bimc_dbgcmd2_REG[2] ( .CK(clk), .CE(n243), .R(n261), .D(n8), .Q(o_bimc_dbgcmd2[2]));
Q_FDP4EP \o_bimc_dbgcmd2_REG[3] ( .CK(clk), .CE(n243), .R(n261), .D(n9), .Q(o_bimc_dbgcmd2[3]));
Q_FDP4EP \o_bimc_dbgcmd2_REG[4] ( .CK(clk), .CE(n243), .R(n261), .D(n10), .Q(o_bimc_dbgcmd2[4]));
Q_FDP4EP \o_bimc_dbgcmd2_REG[5] ( .CK(clk), .CE(n243), .R(n261), .D(n11), .Q(o_bimc_dbgcmd2[5]));
Q_FDP4EP \o_bimc_dbgcmd2_REG[6] ( .CK(clk), .CE(n243), .R(n261), .D(n12), .Q(o_bimc_dbgcmd2[6]));
Q_FDP4EP \o_bimc_dbgcmd2_REG[7] ( .CK(clk), .CE(n243), .R(n261), .D(n13), .Q(o_bimc_dbgcmd2[7]));
Q_FDP4EP \o_bimc_dbgcmd2_REG[8] ( .CK(clk), .CE(n243), .R(n261), .D(n14), .Q(o_bimc_dbgcmd2[8]));
Q_FDP4EP \o_bimc_pollrsp2_REG[0] ( .CK(clk), .CE(n242), .R(n261), .D(n6), .Q(o_bimc_pollrsp2[0]));
Q_FDP4EP \o_bimc_pollrsp2_REG[1] ( .CK(clk), .CE(n242), .R(n261), .D(n7), .Q(o_bimc_pollrsp2[1]));
Q_FDP4EP \o_bimc_pollrsp2_REG[2] ( .CK(clk), .CE(n242), .R(n261), .D(n8), .Q(o_bimc_pollrsp2[2]));
Q_FDP4EP \o_bimc_pollrsp2_REG[3] ( .CK(clk), .CE(n242), .R(n261), .D(n9), .Q(o_bimc_pollrsp2[3]));
Q_FDP4EP \o_bimc_pollrsp2_REG[4] ( .CK(clk), .CE(n242), .R(n261), .D(n10), .Q(o_bimc_pollrsp2[4]));
Q_FDP4EP \o_bimc_pollrsp2_REG[5] ( .CK(clk), .CE(n242), .R(n261), .D(n11), .Q(o_bimc_pollrsp2[5]));
Q_FDP4EP \o_bimc_pollrsp2_REG[6] ( .CK(clk), .CE(n242), .R(n261), .D(n12), .Q(o_bimc_pollrsp2[6]));
Q_FDP4EP \o_bimc_pollrsp2_REG[7] ( .CK(clk), .CE(n242), .R(n261), .D(n13), .Q(o_bimc_pollrsp2[7]));
Q_FDP4EP \o_bimc_pollrsp2_REG[8] ( .CK(clk), .CE(n242), .R(n261), .D(n14), .Q(o_bimc_pollrsp2[8]));
Q_FDP4EP \o_bimc_rxrsp2_REG[0] ( .CK(clk), .CE(n241), .R(n261), .D(n6), .Q(o_bimc_rxrsp2[0]));
Q_FDP4EP \o_bimc_rxrsp2_REG[1] ( .CK(clk), .CE(n241), .R(n261), .D(n7), .Q(o_bimc_rxrsp2[1]));
Q_FDP4EP \o_bimc_rxrsp2_REG[2] ( .CK(clk), .CE(n241), .R(n261), .D(n8), .Q(o_bimc_rxrsp2[2]));
Q_FDP4EP \o_bimc_rxrsp2_REG[3] ( .CK(clk), .CE(n241), .R(n261), .D(n9), .Q(o_bimc_rxrsp2[3]));
Q_FDP4EP \o_bimc_rxrsp2_REG[4] ( .CK(clk), .CE(n241), .R(n261), .D(n10), .Q(o_bimc_rxrsp2[4]));
Q_FDP4EP \o_bimc_rxrsp2_REG[5] ( .CK(clk), .CE(n241), .R(n261), .D(n11), .Q(o_bimc_rxrsp2[5]));
Q_FDP4EP \o_bimc_rxrsp2_REG[6] ( .CK(clk), .CE(n241), .R(n261), .D(n12), .Q(o_bimc_rxrsp2[6]));
Q_FDP4EP \o_bimc_rxrsp2_REG[7] ( .CK(clk), .CE(n241), .R(n261), .D(n13), .Q(o_bimc_rxrsp2[7]));
Q_FDP4EP \o_bimc_rxrsp2_REG[8] ( .CK(clk), .CE(n241), .R(n261), .D(n14), .Q(o_bimc_rxrsp2[8]));
Q_FDP4EP \o_bimc_rxcmd2_REG[0] ( .CK(clk), .CE(n240), .R(n261), .D(n6), .Q(o_bimc_rxcmd2[0]));
Q_FDP4EP \o_bimc_rxcmd2_REG[1] ( .CK(clk), .CE(n240), .R(n261), .D(n7), .Q(o_bimc_rxcmd2[1]));
Q_FDP4EP \o_bimc_rxcmd2_REG[2] ( .CK(clk), .CE(n240), .R(n261), .D(n8), .Q(o_bimc_rxcmd2[2]));
Q_FDP4EP \o_bimc_rxcmd2_REG[3] ( .CK(clk), .CE(n240), .R(n261), .D(n9), .Q(o_bimc_rxcmd2[3]));
Q_FDP4EP \o_bimc_rxcmd2_REG[4] ( .CK(clk), .CE(n240), .R(n261), .D(n10), .Q(o_bimc_rxcmd2[4]));
Q_FDP4EP \o_bimc_rxcmd2_REG[5] ( .CK(clk), .CE(n240), .R(n261), .D(n11), .Q(o_bimc_rxcmd2[5]));
Q_FDP4EP \o_bimc_rxcmd2_REG[6] ( .CK(clk), .CE(n240), .R(n261), .D(n12), .Q(o_bimc_rxcmd2[6]));
Q_FDP4EP \o_bimc_rxcmd2_REG[7] ( .CK(clk), .CE(n240), .R(n261), .D(n13), .Q(o_bimc_rxcmd2[7]));
Q_FDP4EP \o_bimc_rxcmd2_REG[8] ( .CK(clk), .CE(n240), .R(n261), .D(n14), .Q(o_bimc_rxcmd2[8]));
Q_FDP4EP \o_bimc_cmd0_REG[0] ( .CK(clk), .CE(n239), .R(n261), .D(n6), .Q(o_bimc_cmd0[0]));
Q_FDP4EP \o_bimc_cmd0_REG[1] ( .CK(clk), .CE(n239), .R(n261), .D(n7), .Q(o_bimc_cmd0[1]));
Q_FDP4EP \o_bimc_cmd0_REG[2] ( .CK(clk), .CE(n239), .R(n261), .D(n8), .Q(o_bimc_cmd0[2]));
Q_FDP4EP \o_bimc_cmd0_REG[3] ( .CK(clk), .CE(n239), .R(n261), .D(n9), .Q(o_bimc_cmd0[3]));
Q_FDP4EP \o_bimc_cmd0_REG[4] ( .CK(clk), .CE(n239), .R(n261), .D(n10), .Q(o_bimc_cmd0[4]));
Q_FDP4EP \o_bimc_cmd0_REG[5] ( .CK(clk), .CE(n239), .R(n261), .D(n11), .Q(o_bimc_cmd0[5]));
Q_FDP4EP \o_bimc_cmd0_REG[6] ( .CK(clk), .CE(n239), .R(n261), .D(n12), .Q(o_bimc_cmd0[6]));
Q_FDP4EP \o_bimc_cmd0_REG[7] ( .CK(clk), .CE(n239), .R(n261), .D(n13), .Q(o_bimc_cmd0[7]));
Q_FDP4EP \o_bimc_cmd0_REG[8] ( .CK(clk), .CE(n239), .R(n261), .D(n14), .Q(o_bimc_cmd0[8]));
Q_FDP4EP \o_bimc_cmd0_REG[9] ( .CK(clk), .CE(n239), .R(n261), .D(n15), .Q(o_bimc_cmd0[9]));
Q_FDP4EP \o_bimc_cmd0_REG[10] ( .CK(clk), .CE(n239), .R(n261), .D(n16), .Q(o_bimc_cmd0[10]));
Q_FDP4EP \o_bimc_cmd0_REG[11] ( .CK(clk), .CE(n239), .R(n261), .D(n17), .Q(o_bimc_cmd0[11]));
Q_FDP4EP \o_bimc_cmd0_REG[12] ( .CK(clk), .CE(n239), .R(n261), .D(n18), .Q(o_bimc_cmd0[12]));
Q_FDP4EP \o_bimc_cmd0_REG[13] ( .CK(clk), .CE(n239), .R(n261), .D(n19), .Q(o_bimc_cmd0[13]));
Q_FDP4EP \o_bimc_cmd0_REG[14] ( .CK(clk), .CE(n239), .R(n261), .D(n20), .Q(o_bimc_cmd0[14]));
Q_FDP4EP \o_bimc_cmd0_REG[15] ( .CK(clk), .CE(n239), .R(n261), .D(n21), .Q(o_bimc_cmd0[15]));
Q_FDP4EP \o_bimc_cmd0_REG[16] ( .CK(clk), .CE(n239), .R(n261), .D(n22), .Q(o_bimc_cmd0[16]));
Q_FDP4EP \o_bimc_cmd0_REG[17] ( .CK(clk), .CE(n239), .R(n261), .D(n23), .Q(o_bimc_cmd0[17]));
Q_FDP4EP \o_bimc_cmd0_REG[18] ( .CK(clk), .CE(n239), .R(n261), .D(n24), .Q(o_bimc_cmd0[18]));
Q_FDP4EP \o_bimc_cmd0_REG[19] ( .CK(clk), .CE(n239), .R(n261), .D(n25), .Q(o_bimc_cmd0[19]));
Q_FDP4EP \o_bimc_cmd0_REG[20] ( .CK(clk), .CE(n239), .R(n261), .D(n26), .Q(o_bimc_cmd0[20]));
Q_FDP4EP \o_bimc_cmd0_REG[21] ( .CK(clk), .CE(n239), .R(n261), .D(n27), .Q(o_bimc_cmd0[21]));
Q_FDP4EP \o_bimc_cmd0_REG[22] ( .CK(clk), .CE(n239), .R(n261), .D(n28), .Q(o_bimc_cmd0[22]));
Q_FDP4EP \o_bimc_cmd0_REG[23] ( .CK(clk), .CE(n239), .R(n261), .D(n29), .Q(o_bimc_cmd0[23]));
Q_FDP4EP \o_bimc_cmd0_REG[24] ( .CK(clk), .CE(n239), .R(n261), .D(n30), .Q(o_bimc_cmd0[24]));
Q_FDP4EP \o_bimc_cmd0_REG[25] ( .CK(clk), .CE(n239), .R(n261), .D(n31), .Q(o_bimc_cmd0[25]));
Q_FDP4EP \o_bimc_cmd0_REG[26] ( .CK(clk), .CE(n239), .R(n261), .D(n32), .Q(o_bimc_cmd0[26]));
Q_FDP4EP \o_bimc_cmd0_REG[27] ( .CK(clk), .CE(n239), .R(n261), .D(n33), .Q(o_bimc_cmd0[27]));
Q_FDP4EP \o_bimc_cmd0_REG[28] ( .CK(clk), .CE(n239), .R(n261), .D(n34), .Q(o_bimc_cmd0[28]));
Q_FDP4EP \o_bimc_cmd0_REG[29] ( .CK(clk), .CE(n239), .R(n261), .D(n35), .Q(o_bimc_cmd0[29]));
Q_FDP4EP \o_bimc_cmd0_REG[30] ( .CK(clk), .CE(n239), .R(n261), .D(n36), .Q(o_bimc_cmd0[30]));
Q_FDP4EP \o_bimc_cmd0_REG[31] ( .CK(clk), .CE(n239), .R(n261), .D(n37), .Q(o_bimc_cmd0[31]));
Q_FDP4EP \o_bimc_cmd1_REG[0] ( .CK(clk), .CE(n238), .R(n261), .D(n6), .Q(o_bimc_cmd1[0]));
Q_FDP4EP \o_bimc_cmd1_REG[1] ( .CK(clk), .CE(n238), .R(n261), .D(n7), .Q(o_bimc_cmd1[1]));
Q_FDP4EP \o_bimc_cmd1_REG[2] ( .CK(clk), .CE(n238), .R(n261), .D(n8), .Q(o_bimc_cmd1[2]));
Q_FDP4EP \o_bimc_cmd1_REG[3] ( .CK(clk), .CE(n238), .R(n261), .D(n9), .Q(o_bimc_cmd1[3]));
Q_FDP4EP \o_bimc_cmd1_REG[4] ( .CK(clk), .CE(n238), .R(n261), .D(n10), .Q(o_bimc_cmd1[4]));
Q_FDP4EP \o_bimc_cmd1_REG[5] ( .CK(clk), .CE(n238), .R(n261), .D(n11), .Q(o_bimc_cmd1[5]));
Q_FDP4EP \o_bimc_cmd1_REG[6] ( .CK(clk), .CE(n238), .R(n261), .D(n12), .Q(o_bimc_cmd1[6]));
Q_FDP4EP \o_bimc_cmd1_REG[7] ( .CK(clk), .CE(n238), .R(n261), .D(n13), .Q(o_bimc_cmd1[7]));
Q_FDP4EP \o_bimc_cmd1_REG[8] ( .CK(clk), .CE(n238), .R(n261), .D(n14), .Q(o_bimc_cmd1[8]));
Q_FDP4EP \o_bimc_cmd1_REG[9] ( .CK(clk), .CE(n238), .R(n261), .D(n15), .Q(o_bimc_cmd1[9]));
Q_FDP4EP \o_bimc_cmd1_REG[10] ( .CK(clk), .CE(n238), .R(n261), .D(n16), .Q(o_bimc_cmd1[10]));
Q_FDP4EP \o_bimc_cmd1_REG[11] ( .CK(clk), .CE(n238), .R(n261), .D(n17), .Q(o_bimc_cmd1[11]));
Q_FDP4EP \o_bimc_cmd1_REG[12] ( .CK(clk), .CE(n238), .R(n261), .D(n18), .Q(o_bimc_cmd1[12]));
Q_FDP4EP \o_bimc_cmd1_REG[13] ( .CK(clk), .CE(n238), .R(n261), .D(n19), .Q(o_bimc_cmd1[13]));
Q_FDP4EP \o_bimc_cmd1_REG[14] ( .CK(clk), .CE(n238), .R(n261), .D(n20), .Q(o_bimc_cmd1[14]));
Q_FDP4EP \o_bimc_cmd1_REG[15] ( .CK(clk), .CE(n238), .R(n261), .D(n21), .Q(o_bimc_cmd1[15]));
Q_FDP4EP \o_bimc_cmd1_REG[16] ( .CK(clk), .CE(n238), .R(n261), .D(n22), .Q(o_bimc_cmd1[16]));
Q_FDP4EP \o_bimc_cmd1_REG[17] ( .CK(clk), .CE(n238), .R(n261), .D(n23), .Q(o_bimc_cmd1[17]));
Q_FDP4EP \o_bimc_cmd1_REG[18] ( .CK(clk), .CE(n238), .R(n261), .D(n24), .Q(o_bimc_cmd1[18]));
Q_FDP4EP \o_bimc_cmd1_REG[19] ( .CK(clk), .CE(n238), .R(n261), .D(n25), .Q(o_bimc_cmd1[19]));
Q_FDP4EP \o_bimc_cmd1_REG[20] ( .CK(clk), .CE(n238), .R(n261), .D(n26), .Q(o_bimc_cmd1[20]));
Q_FDP4EP \o_bimc_cmd1_REG[21] ( .CK(clk), .CE(n238), .R(n261), .D(n27), .Q(o_bimc_cmd1[21]));
Q_FDP4EP \o_bimc_cmd1_REG[22] ( .CK(clk), .CE(n238), .R(n261), .D(n28), .Q(o_bimc_cmd1[22]));
Q_FDP4EP \o_bimc_cmd1_REG[23] ( .CK(clk), .CE(n238), .R(n261), .D(n29), .Q(o_bimc_cmd1[23]));
Q_FDP4EP \o_bimc_cmd1_REG[24] ( .CK(clk), .CE(n238), .R(n261), .D(n30), .Q(o_bimc_cmd1[24]));
Q_FDP4EP \o_bimc_cmd1_REG[25] ( .CK(clk), .CE(n238), .R(n261), .D(n31), .Q(o_bimc_cmd1[25]));
Q_FDP4EP \o_bimc_cmd1_REG[26] ( .CK(clk), .CE(n238), .R(n261), .D(n32), .Q(o_bimc_cmd1[26]));
Q_FDP4EP \o_bimc_cmd1_REG[27] ( .CK(clk), .CE(n238), .R(n261), .D(n33), .Q(o_bimc_cmd1[27]));
Q_FDP4EP \o_bimc_cmd1_REG[28] ( .CK(clk), .CE(n238), .R(n261), .D(n34), .Q(o_bimc_cmd1[28]));
Q_FDP4EP \o_bimc_cmd1_REG[29] ( .CK(clk), .CE(n238), .R(n261), .D(n35), .Q(o_bimc_cmd1[29]));
Q_FDP4EP \o_bimc_cmd1_REG[30] ( .CK(clk), .CE(n238), .R(n261), .D(n36), .Q(o_bimc_cmd1[30]));
Q_FDP4EP \o_bimc_cmd1_REG[31] ( .CK(clk), .CE(n238), .R(n261), .D(n37), .Q(o_bimc_cmd1[31]));
Q_FDP4EP \o_bimc_cmd2_REG[0] ( .CK(clk), .CE(n237), .R(n261), .D(n6), .Q(o_bimc_cmd2[0]));
Q_FDP4EP \o_bimc_cmd2_REG[1] ( .CK(clk), .CE(n237), .R(n261), .D(n7), .Q(o_bimc_cmd2[1]));
Q_FDP4EP \o_bimc_cmd2_REG[2] ( .CK(clk), .CE(n237), .R(n261), .D(n8), .Q(o_bimc_cmd2[2]));
Q_FDP4EP \o_bimc_cmd2_REG[3] ( .CK(clk), .CE(n237), .R(n261), .D(n9), .Q(o_bimc_cmd2[3]));
Q_FDP4EP \o_bimc_cmd2_REG[4] ( .CK(clk), .CE(n237), .R(n261), .D(n10), .Q(o_bimc_cmd2[4]));
Q_FDP4EP \o_bimc_cmd2_REG[5] ( .CK(clk), .CE(n237), .R(n261), .D(n11), .Q(o_bimc_cmd2[5]));
Q_FDP4EP \o_bimc_cmd2_REG[6] ( .CK(clk), .CE(n237), .R(n261), .D(n12), .Q(o_bimc_cmd2[6]));
Q_FDP4EP \o_bimc_cmd2_REG[7] ( .CK(clk), .CE(n237), .R(n261), .D(n13), .Q(o_bimc_cmd2[7]));
Q_FDP4EP \o_bimc_cmd2_REG[8] ( .CK(clk), .CE(n237), .R(n261), .D(n14), .Q(o_bimc_cmd2[8]));
Q_FDP4EP \o_bimc_cmd2_REG[9] ( .CK(clk), .CE(n237), .R(n261), .D(n15), .Q(o_bimc_cmd2[9]));
Q_FDP4EP \o_bimc_cmd2_REG[10] ( .CK(clk), .CE(n237), .R(n261), .D(n16), .Q(o_bimc_cmd2[10]));
Q_FDP4EP \o_bimc_eccpar_debug_REG[0] ( .CK(clk), .CE(n236), .R(n261), .D(n6), .Q(o_bimc_eccpar_debug[0]));
Q_FDP4EP \o_bimc_eccpar_debug_REG[1] ( .CK(clk), .CE(n236), .R(n261), .D(n7), .Q(o_bimc_eccpar_debug[1]));
Q_FDP4EP \o_bimc_eccpar_debug_REG[2] ( .CK(clk), .CE(n236), .R(n261), .D(n8), .Q(o_bimc_eccpar_debug[2]));
Q_FDP4EP \o_bimc_eccpar_debug_REG[3] ( .CK(clk), .CE(n236), .R(n261), .D(n9), .Q(o_bimc_eccpar_debug[3]));
Q_FDP4EP \o_bimc_eccpar_debug_REG[4] ( .CK(clk), .CE(n236), .R(n261), .D(n10), .Q(o_bimc_eccpar_debug[4]));
Q_FDP4EP \o_bimc_eccpar_debug_REG[5] ( .CK(clk), .CE(n236), .R(n261), .D(n11), .Q(o_bimc_eccpar_debug[5]));
Q_FDP4EP \o_bimc_eccpar_debug_REG[6] ( .CK(clk), .CE(n236), .R(n261), .D(n12), .Q(o_bimc_eccpar_debug[6]));
Q_FDP4EP \o_bimc_eccpar_debug_REG[7] ( .CK(clk), .CE(n236), .R(n261), .D(n13), .Q(o_bimc_eccpar_debug[7]));
Q_FDP4EP \o_bimc_eccpar_debug_REG[8] ( .CK(clk), .CE(n236), .R(n261), .D(n14), .Q(o_bimc_eccpar_debug[8]));
Q_FDP4EP \o_bimc_eccpar_debug_REG[9] ( .CK(clk), .CE(n236), .R(n261), .D(n15), .Q(o_bimc_eccpar_debug[9]));
Q_FDP4EP \o_bimc_eccpar_debug_REG[10] ( .CK(clk), .CE(n236), .R(n261), .D(n16), .Q(o_bimc_eccpar_debug[10]));
Q_FDP4EP \o_bimc_eccpar_debug_REG[11] ( .CK(clk), .CE(n236), .R(n261), .D(n17), .Q(o_bimc_eccpar_debug[11]));
Q_FDP4EP \o_bimc_eccpar_debug_REG[12] ( .CK(clk), .CE(n236), .R(n261), .D(n18), .Q(o_bimc_eccpar_debug[12]));
Q_FDP4EP \o_bimc_eccpar_debug_REG[13] ( .CK(clk), .CE(n236), .R(n261), .D(n19), .Q(o_bimc_eccpar_debug[13]));
Q_FDP4EP \o_bimc_eccpar_debug_REG[14] ( .CK(clk), .CE(n236), .R(n261), .D(n20), .Q(o_bimc_eccpar_debug[14]));
Q_FDP4EP \o_bimc_eccpar_debug_REG[15] ( .CK(clk), .CE(n236), .R(n261), .D(n21), .Q(o_bimc_eccpar_debug[15]));
Q_FDP4EP \o_bimc_eccpar_debug_REG[16] ( .CK(clk), .CE(n236), .R(n261), .D(n22), .Q(o_bimc_eccpar_debug[16]));
Q_FDP4EP \o_bimc_eccpar_debug_REG[17] ( .CK(clk), .CE(n236), .R(n261), .D(n23), .Q(o_bimc_eccpar_debug[17]));
Q_FDP4EP \o_bimc_eccpar_debug_REG[18] ( .CK(clk), .CE(n236), .R(n261), .D(n24), .Q(o_bimc_eccpar_debug[18]));
Q_FDP4EP \o_bimc_eccpar_debug_REG[19] ( .CK(clk), .CE(n236), .R(n261), .D(n25), .Q(o_bimc_eccpar_debug[19]));
Q_FDP4EP \o_bimc_eccpar_debug_REG[20] ( .CK(clk), .CE(n236), .R(n261), .D(n26), .Q(o_bimc_eccpar_debug[20]));
Q_FDP4EP \o_bimc_eccpar_debug_REG[21] ( .CK(clk), .CE(n236), .R(n261), .D(n27), .Q(o_bimc_eccpar_debug[21]));
Q_FDP4EP \o_bimc_eccpar_debug_REG[22] ( .CK(clk), .CE(n236), .R(n261), .D(n28), .Q(o_bimc_eccpar_debug[22]));
Q_FDP4EP \o_bimc_eccpar_debug_REG[23] ( .CK(clk), .CE(n236), .R(n261), .D(n29), .Q(o_bimc_eccpar_debug[23]));
Q_FDP4EP \o_bimc_eccpar_debug_REG[24] ( .CK(clk), .CE(n236), .R(n261), .D(n30), .Q(o_bimc_eccpar_debug[24]));
Q_FDP4EP \o_bimc_eccpar_debug_REG[25] ( .CK(clk), .CE(n236), .R(n261), .D(n31), .Q(o_bimc_eccpar_debug[25]));
Q_FDP4EP \o_bimc_eccpar_debug_REG[26] ( .CK(clk), .CE(n236), .R(n261), .D(n32), .Q(o_bimc_eccpar_debug[26]));
Q_FDP4EP \o_bimc_eccpar_debug_REG[27] ( .CK(clk), .CE(n236), .R(n261), .D(n33), .Q(o_bimc_eccpar_debug[27]));
Q_FDP4EP \o_bimc_eccpar_debug_REG[28] ( .CK(clk), .CE(n236), .R(n261), .D(n34), .Q(o_bimc_eccpar_debug[28]));
Q_FDP4EP \o_bimc_global_config_REG[1] ( .CK(clk), .CE(n235), .R(n261), .D(n7), .Q(o_bimc_global_config[1]));
Q_FDP4EP \o_bimc_global_config_REG[2] ( .CK(clk), .CE(n235), .R(n261), .D(n8), .Q(o_bimc_global_config[2]));
Q_FDP4EP \o_bimc_global_config_REG[3] ( .CK(clk), .CE(n235), .R(n261), .D(n9), .Q(o_bimc_global_config[3]));
Q_FDP4EP \o_bimc_global_config_REG[4] ( .CK(clk), .CE(n235), .R(n261), .D(n10), .Q(o_bimc_global_config[4]));
Q_FDP4EP \o_bimc_global_config_REG[5] ( .CK(clk), .CE(n235), .R(n261), .D(n11), .Q(o_bimc_global_config[5]));
Q_FDP4EP \o_bimc_global_config_REG[6] ( .CK(clk), .CE(n235), .R(n261), .D(n12), .Q(o_bimc_global_config[6]));
Q_FDP4EP \o_bimc_global_config_REG[7] ( .CK(clk), .CE(n235), .R(n261), .D(n13), .Q(o_bimc_global_config[7]));
Q_FDP4EP \o_bimc_global_config_REG[8] ( .CK(clk), .CE(n235), .R(n261), .D(n14), .Q(o_bimc_global_config[8]));
Q_FDP4EP \o_bimc_global_config_REG[9] ( .CK(clk), .CE(n235), .R(n261), .D(n15), .Q(o_bimc_global_config[9]));
Q_FDP4EP \o_bimc_global_config_REG[10] ( .CK(clk), .CE(n235), .R(n261), .D(n16), .Q(o_bimc_global_config[10]));
Q_FDP4EP \o_bimc_global_config_REG[11] ( .CK(clk), .CE(n235), .R(n261), .D(n17), .Q(o_bimc_global_config[11]));
Q_FDP4EP \o_bimc_global_config_REG[12] ( .CK(clk), .CE(n235), .R(n261), .D(n18), .Q(o_bimc_global_config[12]));
Q_FDP4EP \o_bimc_global_config_REG[13] ( .CK(clk), .CE(n235), .R(n261), .D(n19), .Q(o_bimc_global_config[13]));
Q_FDP4EP \o_bimc_global_config_REG[14] ( .CK(clk), .CE(n235), .R(n261), .D(n20), .Q(o_bimc_global_config[14]));
Q_FDP4EP \o_bimc_global_config_REG[15] ( .CK(clk), .CE(n235), .R(n261), .D(n21), .Q(o_bimc_global_config[15]));
Q_FDP4EP \o_bimc_global_config_REG[16] ( .CK(clk), .CE(n235), .R(n261), .D(n22), .Q(o_bimc_global_config[16]));
Q_FDP4EP \o_bimc_global_config_REG[17] ( .CK(clk), .CE(n235), .R(n261), .D(n23), .Q(o_bimc_global_config[17]));
Q_FDP4EP \o_bimc_global_config_REG[18] ( .CK(clk), .CE(n235), .R(n261), .D(n24), .Q(o_bimc_global_config[18]));
Q_FDP4EP \o_bimc_global_config_REG[19] ( .CK(clk), .CE(n235), .R(n261), .D(n25), .Q(o_bimc_global_config[19]));
Q_FDP4EP \o_bimc_global_config_REG[20] ( .CK(clk), .CE(n235), .R(n261), .D(n26), .Q(o_bimc_global_config[20]));
Q_FDP4EP \o_bimc_global_config_REG[21] ( .CK(clk), .CE(n235), .R(n261), .D(n27), .Q(o_bimc_global_config[21]));
Q_FDP4EP \o_bimc_global_config_REG[22] ( .CK(clk), .CE(n235), .R(n261), .D(n28), .Q(o_bimc_global_config[22]));
Q_FDP4EP \o_bimc_global_config_REG[23] ( .CK(clk), .CE(n235), .R(n261), .D(n29), .Q(o_bimc_global_config[23]));
Q_FDP4EP \o_bimc_global_config_REG[24] ( .CK(clk), .CE(n235), .R(n261), .D(n30), .Q(o_bimc_global_config[24]));
Q_FDP4EP \o_bimc_global_config_REG[25] ( .CK(clk), .CE(n235), .R(n261), .D(n31), .Q(o_bimc_global_config[25]));
Q_FDP4EP \o_bimc_global_config_REG[26] ( .CK(clk), .CE(n235), .R(n261), .D(n32), .Q(o_bimc_global_config[26]));
Q_FDP4EP \o_bimc_global_config_REG[27] ( .CK(clk), .CE(n235), .R(n261), .D(n33), .Q(o_bimc_global_config[27]));
Q_FDP4EP \o_bimc_global_config_REG[28] ( .CK(clk), .CE(n235), .R(n261), .D(n34), .Q(o_bimc_global_config[28]));
Q_FDP4EP \o_bimc_global_config_REG[29] ( .CK(clk), .CE(n235), .R(n261), .D(n35), .Q(o_bimc_global_config[29]));
Q_FDP4EP \o_bimc_global_config_REG[30] ( .CK(clk), .CE(n235), .R(n261), .D(n36), .Q(o_bimc_global_config[30]));
Q_FDP4EP \o_bimc_global_config_REG[31] ( .CK(clk), .CE(n235), .R(n261), .D(n37), .Q(o_bimc_global_config[31]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[0] ( .CK(clk), .CE(n234), .R(n261), .D(n6), .Q(o_bimc_parity_error_cnt[0]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[1] ( .CK(clk), .CE(n234), .R(n261), .D(n7), .Q(o_bimc_parity_error_cnt[1]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[2] ( .CK(clk), .CE(n234), .R(n261), .D(n8), .Q(o_bimc_parity_error_cnt[2]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[3] ( .CK(clk), .CE(n234), .R(n261), .D(n9), .Q(o_bimc_parity_error_cnt[3]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[4] ( .CK(clk), .CE(n234), .R(n261), .D(n10), .Q(o_bimc_parity_error_cnt[4]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[5] ( .CK(clk), .CE(n234), .R(n261), .D(n11), .Q(o_bimc_parity_error_cnt[5]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[6] ( .CK(clk), .CE(n234), .R(n261), .D(n12), .Q(o_bimc_parity_error_cnt[6]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[7] ( .CK(clk), .CE(n234), .R(n261), .D(n13), .Q(o_bimc_parity_error_cnt[7]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[8] ( .CK(clk), .CE(n234), .R(n261), .D(n14), .Q(o_bimc_parity_error_cnt[8]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[9] ( .CK(clk), .CE(n234), .R(n261), .D(n15), .Q(o_bimc_parity_error_cnt[9]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[10] ( .CK(clk), .CE(n234), .R(n261), .D(n16), .Q(o_bimc_parity_error_cnt[10]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[11] ( .CK(clk), .CE(n234), .R(n261), .D(n17), .Q(o_bimc_parity_error_cnt[11]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[12] ( .CK(clk), .CE(n234), .R(n261), .D(n18), .Q(o_bimc_parity_error_cnt[12]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[13] ( .CK(clk), .CE(n234), .R(n261), .D(n19), .Q(o_bimc_parity_error_cnt[13]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[14] ( .CK(clk), .CE(n234), .R(n261), .D(n20), .Q(o_bimc_parity_error_cnt[14]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[15] ( .CK(clk), .CE(n234), .R(n261), .D(n21), .Q(o_bimc_parity_error_cnt[15]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[16] ( .CK(clk), .CE(n234), .R(n261), .D(n22), .Q(o_bimc_parity_error_cnt[16]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[17] ( .CK(clk), .CE(n234), .R(n261), .D(n23), .Q(o_bimc_parity_error_cnt[17]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[18] ( .CK(clk), .CE(n234), .R(n261), .D(n24), .Q(o_bimc_parity_error_cnt[18]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[19] ( .CK(clk), .CE(n234), .R(n261), .D(n25), .Q(o_bimc_parity_error_cnt[19]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[20] ( .CK(clk), .CE(n234), .R(n261), .D(n26), .Q(o_bimc_parity_error_cnt[20]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[21] ( .CK(clk), .CE(n234), .R(n261), .D(n27), .Q(o_bimc_parity_error_cnt[21]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[22] ( .CK(clk), .CE(n234), .R(n261), .D(n28), .Q(o_bimc_parity_error_cnt[22]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[23] ( .CK(clk), .CE(n234), .R(n261), .D(n29), .Q(o_bimc_parity_error_cnt[23]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[24] ( .CK(clk), .CE(n234), .R(n261), .D(n30), .Q(o_bimc_parity_error_cnt[24]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[25] ( .CK(clk), .CE(n234), .R(n261), .D(n31), .Q(o_bimc_parity_error_cnt[25]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[26] ( .CK(clk), .CE(n234), .R(n261), .D(n32), .Q(o_bimc_parity_error_cnt[26]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[27] ( .CK(clk), .CE(n234), .R(n261), .D(n33), .Q(o_bimc_parity_error_cnt[27]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[28] ( .CK(clk), .CE(n234), .R(n261), .D(n34), .Q(o_bimc_parity_error_cnt[28]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[29] ( .CK(clk), .CE(n234), .R(n261), .D(n35), .Q(o_bimc_parity_error_cnt[29]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[30] ( .CK(clk), .CE(n234), .R(n261), .D(n36), .Q(o_bimc_parity_error_cnt[30]));
Q_FDP4EP \o_bimc_parity_error_cnt_REG[31] ( .CK(clk), .CE(n234), .R(n261), .D(n37), .Q(o_bimc_parity_error_cnt[31]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[0] ( .CK(clk), .CE(n233), .R(n261), .D(n6), .Q(o_bimc_ecc_correctable_error_cnt[0]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[1] ( .CK(clk), .CE(n233), .R(n261), .D(n7), .Q(o_bimc_ecc_correctable_error_cnt[1]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[2] ( .CK(clk), .CE(n233), .R(n261), .D(n8), .Q(o_bimc_ecc_correctable_error_cnt[2]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[3] ( .CK(clk), .CE(n233), .R(n261), .D(n9), .Q(o_bimc_ecc_correctable_error_cnt[3]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[4] ( .CK(clk), .CE(n233), .R(n261), .D(n10), .Q(o_bimc_ecc_correctable_error_cnt[4]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[5] ( .CK(clk), .CE(n233), .R(n261), .D(n11), .Q(o_bimc_ecc_correctable_error_cnt[5]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[6] ( .CK(clk), .CE(n233), .R(n261), .D(n12), .Q(o_bimc_ecc_correctable_error_cnt[6]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[7] ( .CK(clk), .CE(n233), .R(n261), .D(n13), .Q(o_bimc_ecc_correctable_error_cnt[7]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[8] ( .CK(clk), .CE(n233), .R(n261), .D(n14), .Q(o_bimc_ecc_correctable_error_cnt[8]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[9] ( .CK(clk), .CE(n233), .R(n261), .D(n15), .Q(o_bimc_ecc_correctable_error_cnt[9]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[10] ( .CK(clk), .CE(n233), .R(n261), .D(n16), .Q(o_bimc_ecc_correctable_error_cnt[10]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[11] ( .CK(clk), .CE(n233), .R(n261), .D(n17), .Q(o_bimc_ecc_correctable_error_cnt[11]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[12] ( .CK(clk), .CE(n233), .R(n261), .D(n18), .Q(o_bimc_ecc_correctable_error_cnt[12]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[13] ( .CK(clk), .CE(n233), .R(n261), .D(n19), .Q(o_bimc_ecc_correctable_error_cnt[13]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[14] ( .CK(clk), .CE(n233), .R(n261), .D(n20), .Q(o_bimc_ecc_correctable_error_cnt[14]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[15] ( .CK(clk), .CE(n233), .R(n261), .D(n21), .Q(o_bimc_ecc_correctable_error_cnt[15]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[16] ( .CK(clk), .CE(n233), .R(n261), .D(n22), .Q(o_bimc_ecc_correctable_error_cnt[16]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[17] ( .CK(clk), .CE(n233), .R(n261), .D(n23), .Q(o_bimc_ecc_correctable_error_cnt[17]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[18] ( .CK(clk), .CE(n233), .R(n261), .D(n24), .Q(o_bimc_ecc_correctable_error_cnt[18]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[19] ( .CK(clk), .CE(n233), .R(n261), .D(n25), .Q(o_bimc_ecc_correctable_error_cnt[19]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[20] ( .CK(clk), .CE(n233), .R(n261), .D(n26), .Q(o_bimc_ecc_correctable_error_cnt[20]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[21] ( .CK(clk), .CE(n233), .R(n261), .D(n27), .Q(o_bimc_ecc_correctable_error_cnt[21]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[22] ( .CK(clk), .CE(n233), .R(n261), .D(n28), .Q(o_bimc_ecc_correctable_error_cnt[22]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[23] ( .CK(clk), .CE(n233), .R(n261), .D(n29), .Q(o_bimc_ecc_correctable_error_cnt[23]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[24] ( .CK(clk), .CE(n233), .R(n261), .D(n30), .Q(o_bimc_ecc_correctable_error_cnt[24]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[25] ( .CK(clk), .CE(n233), .R(n261), .D(n31), .Q(o_bimc_ecc_correctable_error_cnt[25]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[26] ( .CK(clk), .CE(n233), .R(n261), .D(n32), .Q(o_bimc_ecc_correctable_error_cnt[26]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[27] ( .CK(clk), .CE(n233), .R(n261), .D(n33), .Q(o_bimc_ecc_correctable_error_cnt[27]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[28] ( .CK(clk), .CE(n233), .R(n261), .D(n34), .Q(o_bimc_ecc_correctable_error_cnt[28]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[29] ( .CK(clk), .CE(n233), .R(n261), .D(n35), .Q(o_bimc_ecc_correctable_error_cnt[29]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[30] ( .CK(clk), .CE(n233), .R(n261), .D(n36), .Q(o_bimc_ecc_correctable_error_cnt[30]));
Q_FDP4EP \o_bimc_ecc_correctable_error_cnt_REG[31] ( .CK(clk), .CE(n233), .R(n261), .D(n37), .Q(o_bimc_ecc_correctable_error_cnt[31]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[0] ( .CK(clk), .CE(n232), .R(n261), .D(n6), .Q(o_bimc_ecc_uncorrectable_error_cnt[0]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[1] ( .CK(clk), .CE(n232), .R(n261), .D(n7), .Q(o_bimc_ecc_uncorrectable_error_cnt[1]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[2] ( .CK(clk), .CE(n232), .R(n261), .D(n8), .Q(o_bimc_ecc_uncorrectable_error_cnt[2]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[3] ( .CK(clk), .CE(n232), .R(n261), .D(n9), .Q(o_bimc_ecc_uncorrectable_error_cnt[3]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[4] ( .CK(clk), .CE(n232), .R(n261), .D(n10), .Q(o_bimc_ecc_uncorrectable_error_cnt[4]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[5] ( .CK(clk), .CE(n232), .R(n261), .D(n11), .Q(o_bimc_ecc_uncorrectable_error_cnt[5]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[6] ( .CK(clk), .CE(n232), .R(n261), .D(n12), .Q(o_bimc_ecc_uncorrectable_error_cnt[6]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[7] ( .CK(clk), .CE(n232), .R(n261), .D(n13), .Q(o_bimc_ecc_uncorrectable_error_cnt[7]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[8] ( .CK(clk), .CE(n232), .R(n261), .D(n14), .Q(o_bimc_ecc_uncorrectable_error_cnt[8]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[9] ( .CK(clk), .CE(n232), .R(n261), .D(n15), .Q(o_bimc_ecc_uncorrectable_error_cnt[9]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[10] ( .CK(clk), .CE(n232), .R(n261), .D(n16), .Q(o_bimc_ecc_uncorrectable_error_cnt[10]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[11] ( .CK(clk), .CE(n232), .R(n261), .D(n17), .Q(o_bimc_ecc_uncorrectable_error_cnt[11]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[12] ( .CK(clk), .CE(n232), .R(n261), .D(n18), .Q(o_bimc_ecc_uncorrectable_error_cnt[12]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[13] ( .CK(clk), .CE(n232), .R(n261), .D(n19), .Q(o_bimc_ecc_uncorrectable_error_cnt[13]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[14] ( .CK(clk), .CE(n232), .R(n261), .D(n20), .Q(o_bimc_ecc_uncorrectable_error_cnt[14]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[15] ( .CK(clk), .CE(n232), .R(n261), .D(n21), .Q(o_bimc_ecc_uncorrectable_error_cnt[15]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[16] ( .CK(clk), .CE(n232), .R(n261), .D(n22), .Q(o_bimc_ecc_uncorrectable_error_cnt[16]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[17] ( .CK(clk), .CE(n232), .R(n261), .D(n23), .Q(o_bimc_ecc_uncorrectable_error_cnt[17]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[18] ( .CK(clk), .CE(n232), .R(n261), .D(n24), .Q(o_bimc_ecc_uncorrectable_error_cnt[18]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[19] ( .CK(clk), .CE(n232), .R(n261), .D(n25), .Q(o_bimc_ecc_uncorrectable_error_cnt[19]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[20] ( .CK(clk), .CE(n232), .R(n261), .D(n26), .Q(o_bimc_ecc_uncorrectable_error_cnt[20]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[21] ( .CK(clk), .CE(n232), .R(n261), .D(n27), .Q(o_bimc_ecc_uncorrectable_error_cnt[21]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[22] ( .CK(clk), .CE(n232), .R(n261), .D(n28), .Q(o_bimc_ecc_uncorrectable_error_cnt[22]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[23] ( .CK(clk), .CE(n232), .R(n261), .D(n29), .Q(o_bimc_ecc_uncorrectable_error_cnt[23]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[24] ( .CK(clk), .CE(n232), .R(n261), .D(n30), .Q(o_bimc_ecc_uncorrectable_error_cnt[24]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[25] ( .CK(clk), .CE(n232), .R(n261), .D(n31), .Q(o_bimc_ecc_uncorrectable_error_cnt[25]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[26] ( .CK(clk), .CE(n232), .R(n261), .D(n32), .Q(o_bimc_ecc_uncorrectable_error_cnt[26]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[27] ( .CK(clk), .CE(n232), .R(n261), .D(n33), .Q(o_bimc_ecc_uncorrectable_error_cnt[27]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[28] ( .CK(clk), .CE(n232), .R(n261), .D(n34), .Q(o_bimc_ecc_uncorrectable_error_cnt[28]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[29] ( .CK(clk), .CE(n232), .R(n261), .D(n35), .Q(o_bimc_ecc_uncorrectable_error_cnt[29]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[30] ( .CK(clk), .CE(n232), .R(n261), .D(n36), .Q(o_bimc_ecc_uncorrectable_error_cnt[30]));
Q_FDP4EP \o_bimc_ecc_uncorrectable_error_cnt_REG[31] ( .CK(clk), .CE(n232), .R(n261), .D(n37), .Q(o_bimc_ecc_uncorrectable_error_cnt[31]));
Q_FDP4EP \o_bimc_monitor_mask_REG[0] ( .CK(clk), .CE(n231), .R(n261), .D(n6), .Q(o_bimc_monitor_mask[0]));
Q_FDP4EP \o_bimc_monitor_mask_REG[1] ( .CK(clk), .CE(n231), .R(n261), .D(n7), .Q(o_bimc_monitor_mask[1]));
Q_FDP4EP \o_bimc_monitor_mask_REG[2] ( .CK(clk), .CE(n231), .R(n261), .D(n8), .Q(o_bimc_monitor_mask[2]));
Q_FDP4EP \o_bimc_monitor_mask_REG[3] ( .CK(clk), .CE(n231), .R(n261), .D(n9), .Q(o_bimc_monitor_mask[3]));
Q_FDP4EP \o_bimc_monitor_mask_REG[4] ( .CK(clk), .CE(n231), .R(n261), .D(n10), .Q(o_bimc_monitor_mask[4]));
Q_FDP4EP \o_bimc_monitor_mask_REG[5] ( .CK(clk), .CE(n231), .R(n261), .D(n11), .Q(o_bimc_monitor_mask[5]));
Q_FDP4EP \o_bimc_monitor_mask_REG[6] ( .CK(clk), .CE(n231), .R(n261), .D(n12), .Q(o_bimc_monitor_mask[6]));
Q_FDP4EP \o_engine_sticky_status_REG[0] ( .CK(clk), .CE(n230), .R(n261), .D(n6), .Q(o_engine_sticky_status[0]));
Q_FDP4EP \o_engine_sticky_status_REG[1] ( .CK(clk), .CE(n230), .R(n261), .D(n7), .Q(o_engine_sticky_status[1]));
Q_FDP4EP \o_engine_sticky_status_REG[2] ( .CK(clk), .CE(n230), .R(n261), .D(n8), .Q(o_engine_sticky_status[2]));
Q_FDP4EP \o_engine_sticky_status_REG[3] ( .CK(clk), .CE(n230), .R(n261), .D(n9), .Q(o_engine_sticky_status[3]));
Q_FDP4EP \o_engine_sticky_status_REG[4] ( .CK(clk), .CE(n230), .R(n261), .D(n10), .Q(o_engine_sticky_status[4]));
Q_FDP4EP \o_engine_sticky_status_REG[5] ( .CK(clk), .CE(n230), .R(n261), .D(n11), .Q(o_engine_sticky_status[5]));
Q_FDP4EP \o_engine_sticky_status_REG[6] ( .CK(clk), .CE(n230), .R(n261), .D(n12), .Q(o_engine_sticky_status[6]));
Q_FDP4EP \o_engine_sticky_status_REG[7] ( .CK(clk), .CE(n230), .R(n261), .D(n13), .Q(o_engine_sticky_status[7]));
Q_FDP4EP \o_interrupt_mask_REG[0] ( .CK(clk), .CE(n229), .R(n261), .D(n6), .Q(o_interrupt_mask[0]));
Q_FDP4EP \o_interrupt_mask_REG[1] ( .CK(clk), .CE(n229), .R(n261), .D(n7), .Q(o_interrupt_mask[1]));
Q_FDP4EP \o_interrupt_mask_REG[2] ( .CK(clk), .CE(n229), .R(n261), .D(n8), .Q(o_interrupt_mask[2]));
Q_FDP4EP \o_interrupt_mask_REG[3] ( .CK(clk), .CE(n229), .R(n261), .D(n9), .Q(o_interrupt_mask[3]));
Q_FDP4EP \o_interrupt_mask_REG[4] ( .CK(clk), .CE(n229), .R(n261), .D(n10), .Q(o_interrupt_mask[4]));
Q_FDP4EP \o_interrupt_status_REG[0] ( .CK(clk), .CE(n228), .R(n261), .D(n6), .Q(o_interrupt_status[0]));
Q_FDP4EP \o_interrupt_status_REG[1] ( .CK(clk), .CE(n228), .R(n261), .D(n7), .Q(o_interrupt_status[1]));
Q_FDP4EP \o_interrupt_status_REG[2] ( .CK(clk), .CE(n228), .R(n261), .D(n8), .Q(o_interrupt_status[2]));
Q_FDP4EP \o_interrupt_status_REG[3] ( .CK(clk), .CE(n228), .R(n261), .D(n9), .Q(o_interrupt_status[3]));
Q_FDP4EP \o_interrupt_status_REG[4] ( .CK(clk), .CE(n228), .R(n261), .D(n10), .Q(o_interrupt_status[4]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_1_REG[0] ( .CK(clk), .CE(n227), .R(n261), .D(n6), .Q(o_kdf_drbg_seed_1_reseed_interval_1[0]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_1_REG[1] ( .CK(clk), .CE(n227), .R(n261), .D(n7), .Q(o_kdf_drbg_seed_1_reseed_interval_1[1]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_1_REG[2] ( .CK(clk), .CE(n227), .R(n261), .D(n8), .Q(o_kdf_drbg_seed_1_reseed_interval_1[2]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_1_REG[3] ( .CK(clk), .CE(n227), .R(n261), .D(n9), .Q(o_kdf_drbg_seed_1_reseed_interval_1[3]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_1_REG[4] ( .CK(clk), .CE(n227), .R(n261), .D(n10), .Q(o_kdf_drbg_seed_1_reseed_interval_1[4]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_1_REG[5] ( .CK(clk), .CE(n227), .R(n261), .D(n11), .Q(o_kdf_drbg_seed_1_reseed_interval_1[5]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_1_REG[6] ( .CK(clk), .CE(n227), .R(n261), .D(n12), .Q(o_kdf_drbg_seed_1_reseed_interval_1[6]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_1_REG[7] ( .CK(clk), .CE(n227), .R(n261), .D(n13), .Q(o_kdf_drbg_seed_1_reseed_interval_1[7]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_1_REG[8] ( .CK(clk), .CE(n227), .R(n261), .D(n14), .Q(o_kdf_drbg_seed_1_reseed_interval_1[8]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_1_REG[9] ( .CK(clk), .CE(n227), .R(n261), .D(n15), .Q(o_kdf_drbg_seed_1_reseed_interval_1[9]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_1_REG[10] ( .CK(clk), .CE(n227), .R(n261), .D(n16), .Q(o_kdf_drbg_seed_1_reseed_interval_1[10]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_1_REG[11] ( .CK(clk), .CE(n227), .R(n261), .D(n17), .Q(o_kdf_drbg_seed_1_reseed_interval_1[11]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_1_REG[12] ( .CK(clk), .CE(n227), .R(n261), .D(n18), .Q(o_kdf_drbg_seed_1_reseed_interval_1[12]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_1_REG[13] ( .CK(clk), .CE(n227), .R(n261), .D(n19), .Q(o_kdf_drbg_seed_1_reseed_interval_1[13]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_1_REG[14] ( .CK(clk), .CE(n227), .R(n261), .D(n20), .Q(o_kdf_drbg_seed_1_reseed_interval_1[14]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_1_REG[15] ( .CK(clk), .CE(n227), .R(n261), .D(n21), .Q(o_kdf_drbg_seed_1_reseed_interval_1[15]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[0] ( .CK(clk), .CE(n226), .R(n261), .D(n6), .Q(o_kdf_drbg_seed_1_reseed_interval_0[0]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[1] ( .CK(clk), .CE(n226), .R(n261), .D(n7), .Q(o_kdf_drbg_seed_1_reseed_interval_0[1]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[2] ( .CK(clk), .CE(n226), .R(n261), .D(n8), .Q(o_kdf_drbg_seed_1_reseed_interval_0[2]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[3] ( .CK(clk), .CE(n226), .R(n261), .D(n9), .Q(o_kdf_drbg_seed_1_reseed_interval_0[3]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[4] ( .CK(clk), .CE(n226), .R(n261), .D(n10), .Q(o_kdf_drbg_seed_1_reseed_interval_0[4]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[5] ( .CK(clk), .CE(n226), .R(n261), .D(n11), .Q(o_kdf_drbg_seed_1_reseed_interval_0[5]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[6] ( .CK(clk), .CE(n226), .R(n261), .D(n12), .Q(o_kdf_drbg_seed_1_reseed_interval_0[6]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[7] ( .CK(clk), .CE(n226), .R(n261), .D(n13), .Q(o_kdf_drbg_seed_1_reseed_interval_0[7]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[8] ( .CK(clk), .CE(n226), .R(n261), .D(n14), .Q(o_kdf_drbg_seed_1_reseed_interval_0[8]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[9] ( .CK(clk), .CE(n226), .R(n261), .D(n15), .Q(o_kdf_drbg_seed_1_reseed_interval_0[9]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[10] ( .CK(clk), .CE(n226), .R(n261), .D(n16), .Q(o_kdf_drbg_seed_1_reseed_interval_0[10]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[11] ( .CK(clk), .CE(n226), .R(n261), .D(n17), .Q(o_kdf_drbg_seed_1_reseed_interval_0[11]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[12] ( .CK(clk), .CE(n226), .R(n261), .D(n18), .Q(o_kdf_drbg_seed_1_reseed_interval_0[12]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[13] ( .CK(clk), .CE(n226), .R(n261), .D(n19), .Q(o_kdf_drbg_seed_1_reseed_interval_0[13]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[14] ( .CK(clk), .CE(n226), .R(n261), .D(n20), .Q(o_kdf_drbg_seed_1_reseed_interval_0[14]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[15] ( .CK(clk), .CE(n226), .R(n261), .D(n21), .Q(o_kdf_drbg_seed_1_reseed_interval_0[15]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[16] ( .CK(clk), .CE(n226), .R(n261), .D(n22), .Q(o_kdf_drbg_seed_1_reseed_interval_0[16]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[17] ( .CK(clk), .CE(n226), .R(n261), .D(n23), .Q(o_kdf_drbg_seed_1_reseed_interval_0[17]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[18] ( .CK(clk), .CE(n226), .R(n261), .D(n24), .Q(o_kdf_drbg_seed_1_reseed_interval_0[18]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[19] ( .CK(clk), .CE(n226), .R(n261), .D(n25), .Q(o_kdf_drbg_seed_1_reseed_interval_0[19]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[20] ( .CK(clk), .CE(n226), .R(n261), .D(n26), .Q(o_kdf_drbg_seed_1_reseed_interval_0[20]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[21] ( .CK(clk), .CE(n226), .R(n261), .D(n27), .Q(o_kdf_drbg_seed_1_reseed_interval_0[21]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[22] ( .CK(clk), .CE(n226), .R(n261), .D(n28), .Q(o_kdf_drbg_seed_1_reseed_interval_0[22]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[23] ( .CK(clk), .CE(n226), .R(n261), .D(n29), .Q(o_kdf_drbg_seed_1_reseed_interval_0[23]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[24] ( .CK(clk), .CE(n226), .R(n261), .D(n30), .Q(o_kdf_drbg_seed_1_reseed_interval_0[24]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[25] ( .CK(clk), .CE(n226), .R(n261), .D(n31), .Q(o_kdf_drbg_seed_1_reseed_interval_0[25]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[26] ( .CK(clk), .CE(n226), .R(n261), .D(n32), .Q(o_kdf_drbg_seed_1_reseed_interval_0[26]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[27] ( .CK(clk), .CE(n226), .R(n261), .D(n33), .Q(o_kdf_drbg_seed_1_reseed_interval_0[27]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[28] ( .CK(clk), .CE(n226), .R(n261), .D(n34), .Q(o_kdf_drbg_seed_1_reseed_interval_0[28]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[29] ( .CK(clk), .CE(n226), .R(n261), .D(n35), .Q(o_kdf_drbg_seed_1_reseed_interval_0[29]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[30] ( .CK(clk), .CE(n226), .R(n261), .D(n36), .Q(o_kdf_drbg_seed_1_reseed_interval_0[30]));
Q_FDP4EP \o_kdf_drbg_seed_1_reseed_interval_0_REG[31] ( .CK(clk), .CE(n226), .R(n261), .D(n37), .Q(o_kdf_drbg_seed_1_reseed_interval_0[31]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[0] ( .CK(clk), .CE(n225), .R(n261), .D(n6), .Q(o_kdf_drbg_seed_1_state_value_127_96[0]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[1] ( .CK(clk), .CE(n225), .R(n261), .D(n7), .Q(o_kdf_drbg_seed_1_state_value_127_96[1]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[2] ( .CK(clk), .CE(n225), .R(n261), .D(n8), .Q(o_kdf_drbg_seed_1_state_value_127_96[2]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[3] ( .CK(clk), .CE(n225), .R(n261), .D(n9), .Q(o_kdf_drbg_seed_1_state_value_127_96[3]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[4] ( .CK(clk), .CE(n225), .R(n261), .D(n10), .Q(o_kdf_drbg_seed_1_state_value_127_96[4]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[5] ( .CK(clk), .CE(n225), .R(n261), .D(n11), .Q(o_kdf_drbg_seed_1_state_value_127_96[5]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[6] ( .CK(clk), .CE(n225), .R(n261), .D(n12), .Q(o_kdf_drbg_seed_1_state_value_127_96[6]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[7] ( .CK(clk), .CE(n225), .R(n261), .D(n13), .Q(o_kdf_drbg_seed_1_state_value_127_96[7]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[8] ( .CK(clk), .CE(n225), .R(n261), .D(n14), .Q(o_kdf_drbg_seed_1_state_value_127_96[8]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[9] ( .CK(clk), .CE(n225), .R(n261), .D(n15), .Q(o_kdf_drbg_seed_1_state_value_127_96[9]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[10] ( .CK(clk), .CE(n225), .R(n261), .D(n16), .Q(o_kdf_drbg_seed_1_state_value_127_96[10]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[11] ( .CK(clk), .CE(n225), .R(n261), .D(n17), .Q(o_kdf_drbg_seed_1_state_value_127_96[11]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[12] ( .CK(clk), .CE(n225), .R(n261), .D(n18), .Q(o_kdf_drbg_seed_1_state_value_127_96[12]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[13] ( .CK(clk), .CE(n225), .R(n261), .D(n19), .Q(o_kdf_drbg_seed_1_state_value_127_96[13]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[14] ( .CK(clk), .CE(n225), .R(n261), .D(n20), .Q(o_kdf_drbg_seed_1_state_value_127_96[14]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[15] ( .CK(clk), .CE(n225), .R(n261), .D(n21), .Q(o_kdf_drbg_seed_1_state_value_127_96[15]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[16] ( .CK(clk), .CE(n225), .R(n261), .D(n22), .Q(o_kdf_drbg_seed_1_state_value_127_96[16]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[17] ( .CK(clk), .CE(n225), .R(n261), .D(n23), .Q(o_kdf_drbg_seed_1_state_value_127_96[17]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[18] ( .CK(clk), .CE(n225), .R(n261), .D(n24), .Q(o_kdf_drbg_seed_1_state_value_127_96[18]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[19] ( .CK(clk), .CE(n225), .R(n261), .D(n25), .Q(o_kdf_drbg_seed_1_state_value_127_96[19]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[20] ( .CK(clk), .CE(n225), .R(n261), .D(n26), .Q(o_kdf_drbg_seed_1_state_value_127_96[20]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[21] ( .CK(clk), .CE(n225), .R(n261), .D(n27), .Q(o_kdf_drbg_seed_1_state_value_127_96[21]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[22] ( .CK(clk), .CE(n225), .R(n261), .D(n28), .Q(o_kdf_drbg_seed_1_state_value_127_96[22]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[23] ( .CK(clk), .CE(n225), .R(n261), .D(n29), .Q(o_kdf_drbg_seed_1_state_value_127_96[23]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[24] ( .CK(clk), .CE(n225), .R(n261), .D(n30), .Q(o_kdf_drbg_seed_1_state_value_127_96[24]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[25] ( .CK(clk), .CE(n225), .R(n261), .D(n31), .Q(o_kdf_drbg_seed_1_state_value_127_96[25]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[26] ( .CK(clk), .CE(n225), .R(n261), .D(n32), .Q(o_kdf_drbg_seed_1_state_value_127_96[26]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[27] ( .CK(clk), .CE(n225), .R(n261), .D(n33), .Q(o_kdf_drbg_seed_1_state_value_127_96[27]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[28] ( .CK(clk), .CE(n225), .R(n261), .D(n34), .Q(o_kdf_drbg_seed_1_state_value_127_96[28]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[29] ( .CK(clk), .CE(n225), .R(n261), .D(n35), .Q(o_kdf_drbg_seed_1_state_value_127_96[29]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[30] ( .CK(clk), .CE(n225), .R(n261), .D(n36), .Q(o_kdf_drbg_seed_1_state_value_127_96[30]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_127_96_REG[31] ( .CK(clk), .CE(n225), .R(n261), .D(n37), .Q(o_kdf_drbg_seed_1_state_value_127_96[31]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[0] ( .CK(clk), .CE(n224), .R(n261), .D(n6), .Q(o_kdf_drbg_seed_1_state_value_95_64[0]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[1] ( .CK(clk), .CE(n224), .R(n261), .D(n7), .Q(o_kdf_drbg_seed_1_state_value_95_64[1]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[2] ( .CK(clk), .CE(n224), .R(n261), .D(n8), .Q(o_kdf_drbg_seed_1_state_value_95_64[2]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[3] ( .CK(clk), .CE(n224), .R(n261), .D(n9), .Q(o_kdf_drbg_seed_1_state_value_95_64[3]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[4] ( .CK(clk), .CE(n224), .R(n261), .D(n10), .Q(o_kdf_drbg_seed_1_state_value_95_64[4]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[5] ( .CK(clk), .CE(n224), .R(n261), .D(n11), .Q(o_kdf_drbg_seed_1_state_value_95_64[5]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[6] ( .CK(clk), .CE(n224), .R(n261), .D(n12), .Q(o_kdf_drbg_seed_1_state_value_95_64[6]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[7] ( .CK(clk), .CE(n224), .R(n261), .D(n13), .Q(o_kdf_drbg_seed_1_state_value_95_64[7]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[8] ( .CK(clk), .CE(n224), .R(n261), .D(n14), .Q(o_kdf_drbg_seed_1_state_value_95_64[8]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[9] ( .CK(clk), .CE(n224), .R(n261), .D(n15), .Q(o_kdf_drbg_seed_1_state_value_95_64[9]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[10] ( .CK(clk), .CE(n224), .R(n261), .D(n16), .Q(o_kdf_drbg_seed_1_state_value_95_64[10]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[11] ( .CK(clk), .CE(n224), .R(n261), .D(n17), .Q(o_kdf_drbg_seed_1_state_value_95_64[11]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[12] ( .CK(clk), .CE(n224), .R(n261), .D(n18), .Q(o_kdf_drbg_seed_1_state_value_95_64[12]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[13] ( .CK(clk), .CE(n224), .R(n261), .D(n19), .Q(o_kdf_drbg_seed_1_state_value_95_64[13]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[14] ( .CK(clk), .CE(n224), .R(n261), .D(n20), .Q(o_kdf_drbg_seed_1_state_value_95_64[14]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[15] ( .CK(clk), .CE(n224), .R(n261), .D(n21), .Q(o_kdf_drbg_seed_1_state_value_95_64[15]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[16] ( .CK(clk), .CE(n224), .R(n261), .D(n22), .Q(o_kdf_drbg_seed_1_state_value_95_64[16]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[17] ( .CK(clk), .CE(n224), .R(n261), .D(n23), .Q(o_kdf_drbg_seed_1_state_value_95_64[17]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[18] ( .CK(clk), .CE(n224), .R(n261), .D(n24), .Q(o_kdf_drbg_seed_1_state_value_95_64[18]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[19] ( .CK(clk), .CE(n224), .R(n261), .D(n25), .Q(o_kdf_drbg_seed_1_state_value_95_64[19]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[20] ( .CK(clk), .CE(n224), .R(n261), .D(n26), .Q(o_kdf_drbg_seed_1_state_value_95_64[20]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[21] ( .CK(clk), .CE(n224), .R(n261), .D(n27), .Q(o_kdf_drbg_seed_1_state_value_95_64[21]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[22] ( .CK(clk), .CE(n224), .R(n261), .D(n28), .Q(o_kdf_drbg_seed_1_state_value_95_64[22]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[23] ( .CK(clk), .CE(n224), .R(n261), .D(n29), .Q(o_kdf_drbg_seed_1_state_value_95_64[23]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[24] ( .CK(clk), .CE(n224), .R(n261), .D(n30), .Q(o_kdf_drbg_seed_1_state_value_95_64[24]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[25] ( .CK(clk), .CE(n224), .R(n261), .D(n31), .Q(o_kdf_drbg_seed_1_state_value_95_64[25]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[26] ( .CK(clk), .CE(n224), .R(n261), .D(n32), .Q(o_kdf_drbg_seed_1_state_value_95_64[26]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[27] ( .CK(clk), .CE(n224), .R(n261), .D(n33), .Q(o_kdf_drbg_seed_1_state_value_95_64[27]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[28] ( .CK(clk), .CE(n224), .R(n261), .D(n34), .Q(o_kdf_drbg_seed_1_state_value_95_64[28]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[29] ( .CK(clk), .CE(n224), .R(n261), .D(n35), .Q(o_kdf_drbg_seed_1_state_value_95_64[29]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[30] ( .CK(clk), .CE(n224), .R(n261), .D(n36), .Q(o_kdf_drbg_seed_1_state_value_95_64[30]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_95_64_REG[31] ( .CK(clk), .CE(n224), .R(n261), .D(n37), .Q(o_kdf_drbg_seed_1_state_value_95_64[31]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[0] ( .CK(clk), .CE(n223), .R(n261), .D(n6), .Q(o_kdf_drbg_seed_1_state_value_63_32[0]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[1] ( .CK(clk), .CE(n223), .R(n261), .D(n7), .Q(o_kdf_drbg_seed_1_state_value_63_32[1]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[2] ( .CK(clk), .CE(n223), .R(n261), .D(n8), .Q(o_kdf_drbg_seed_1_state_value_63_32[2]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[3] ( .CK(clk), .CE(n223), .R(n261), .D(n9), .Q(o_kdf_drbg_seed_1_state_value_63_32[3]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[4] ( .CK(clk), .CE(n223), .R(n261), .D(n10), .Q(o_kdf_drbg_seed_1_state_value_63_32[4]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[5] ( .CK(clk), .CE(n223), .R(n261), .D(n11), .Q(o_kdf_drbg_seed_1_state_value_63_32[5]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[6] ( .CK(clk), .CE(n223), .R(n261), .D(n12), .Q(o_kdf_drbg_seed_1_state_value_63_32[6]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[7] ( .CK(clk), .CE(n223), .R(n261), .D(n13), .Q(o_kdf_drbg_seed_1_state_value_63_32[7]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[8] ( .CK(clk), .CE(n223), .R(n261), .D(n14), .Q(o_kdf_drbg_seed_1_state_value_63_32[8]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[9] ( .CK(clk), .CE(n223), .R(n261), .D(n15), .Q(o_kdf_drbg_seed_1_state_value_63_32[9]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[10] ( .CK(clk), .CE(n223), .R(n261), .D(n16), .Q(o_kdf_drbg_seed_1_state_value_63_32[10]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[11] ( .CK(clk), .CE(n223), .R(n261), .D(n17), .Q(o_kdf_drbg_seed_1_state_value_63_32[11]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[12] ( .CK(clk), .CE(n223), .R(n261), .D(n18), .Q(o_kdf_drbg_seed_1_state_value_63_32[12]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[13] ( .CK(clk), .CE(n223), .R(n261), .D(n19), .Q(o_kdf_drbg_seed_1_state_value_63_32[13]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[14] ( .CK(clk), .CE(n223), .R(n261), .D(n20), .Q(o_kdf_drbg_seed_1_state_value_63_32[14]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[15] ( .CK(clk), .CE(n223), .R(n261), .D(n21), .Q(o_kdf_drbg_seed_1_state_value_63_32[15]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[16] ( .CK(clk), .CE(n223), .R(n261), .D(n22), .Q(o_kdf_drbg_seed_1_state_value_63_32[16]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[17] ( .CK(clk), .CE(n223), .R(n261), .D(n23), .Q(o_kdf_drbg_seed_1_state_value_63_32[17]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[18] ( .CK(clk), .CE(n223), .R(n261), .D(n24), .Q(o_kdf_drbg_seed_1_state_value_63_32[18]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[19] ( .CK(clk), .CE(n223), .R(n261), .D(n25), .Q(o_kdf_drbg_seed_1_state_value_63_32[19]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[20] ( .CK(clk), .CE(n223), .R(n261), .D(n26), .Q(o_kdf_drbg_seed_1_state_value_63_32[20]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[21] ( .CK(clk), .CE(n223), .R(n261), .D(n27), .Q(o_kdf_drbg_seed_1_state_value_63_32[21]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[22] ( .CK(clk), .CE(n223), .R(n261), .D(n28), .Q(o_kdf_drbg_seed_1_state_value_63_32[22]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[23] ( .CK(clk), .CE(n223), .R(n261), .D(n29), .Q(o_kdf_drbg_seed_1_state_value_63_32[23]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[24] ( .CK(clk), .CE(n223), .R(n261), .D(n30), .Q(o_kdf_drbg_seed_1_state_value_63_32[24]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[25] ( .CK(clk), .CE(n223), .R(n261), .D(n31), .Q(o_kdf_drbg_seed_1_state_value_63_32[25]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[26] ( .CK(clk), .CE(n223), .R(n261), .D(n32), .Q(o_kdf_drbg_seed_1_state_value_63_32[26]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[27] ( .CK(clk), .CE(n223), .R(n261), .D(n33), .Q(o_kdf_drbg_seed_1_state_value_63_32[27]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[28] ( .CK(clk), .CE(n223), .R(n261), .D(n34), .Q(o_kdf_drbg_seed_1_state_value_63_32[28]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[29] ( .CK(clk), .CE(n223), .R(n261), .D(n35), .Q(o_kdf_drbg_seed_1_state_value_63_32[29]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[30] ( .CK(clk), .CE(n223), .R(n261), .D(n36), .Q(o_kdf_drbg_seed_1_state_value_63_32[30]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_63_32_REG[31] ( .CK(clk), .CE(n223), .R(n261), .D(n37), .Q(o_kdf_drbg_seed_1_state_value_63_32[31]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[0] ( .CK(clk), .CE(n222), .R(n261), .D(n6), .Q(o_kdf_drbg_seed_1_state_value_31_0[0]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[1] ( .CK(clk), .CE(n222), .R(n261), .D(n7), .Q(o_kdf_drbg_seed_1_state_value_31_0[1]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[2] ( .CK(clk), .CE(n222), .R(n261), .D(n8), .Q(o_kdf_drbg_seed_1_state_value_31_0[2]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[3] ( .CK(clk), .CE(n222), .R(n261), .D(n9), .Q(o_kdf_drbg_seed_1_state_value_31_0[3]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[4] ( .CK(clk), .CE(n222), .R(n261), .D(n10), .Q(o_kdf_drbg_seed_1_state_value_31_0[4]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[5] ( .CK(clk), .CE(n222), .R(n261), .D(n11), .Q(o_kdf_drbg_seed_1_state_value_31_0[5]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[6] ( .CK(clk), .CE(n222), .R(n261), .D(n12), .Q(o_kdf_drbg_seed_1_state_value_31_0[6]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[7] ( .CK(clk), .CE(n222), .R(n261), .D(n13), .Q(o_kdf_drbg_seed_1_state_value_31_0[7]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[8] ( .CK(clk), .CE(n222), .R(n261), .D(n14), .Q(o_kdf_drbg_seed_1_state_value_31_0[8]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[9] ( .CK(clk), .CE(n222), .R(n261), .D(n15), .Q(o_kdf_drbg_seed_1_state_value_31_0[9]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[10] ( .CK(clk), .CE(n222), .R(n261), .D(n16), .Q(o_kdf_drbg_seed_1_state_value_31_0[10]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[11] ( .CK(clk), .CE(n222), .R(n261), .D(n17), .Q(o_kdf_drbg_seed_1_state_value_31_0[11]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[12] ( .CK(clk), .CE(n222), .R(n261), .D(n18), .Q(o_kdf_drbg_seed_1_state_value_31_0[12]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[13] ( .CK(clk), .CE(n222), .R(n261), .D(n19), .Q(o_kdf_drbg_seed_1_state_value_31_0[13]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[14] ( .CK(clk), .CE(n222), .R(n261), .D(n20), .Q(o_kdf_drbg_seed_1_state_value_31_0[14]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[15] ( .CK(clk), .CE(n222), .R(n261), .D(n21), .Q(o_kdf_drbg_seed_1_state_value_31_0[15]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[16] ( .CK(clk), .CE(n222), .R(n261), .D(n22), .Q(o_kdf_drbg_seed_1_state_value_31_0[16]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[17] ( .CK(clk), .CE(n222), .R(n261), .D(n23), .Q(o_kdf_drbg_seed_1_state_value_31_0[17]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[18] ( .CK(clk), .CE(n222), .R(n261), .D(n24), .Q(o_kdf_drbg_seed_1_state_value_31_0[18]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[19] ( .CK(clk), .CE(n222), .R(n261), .D(n25), .Q(o_kdf_drbg_seed_1_state_value_31_0[19]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[20] ( .CK(clk), .CE(n222), .R(n261), .D(n26), .Q(o_kdf_drbg_seed_1_state_value_31_0[20]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[21] ( .CK(clk), .CE(n222), .R(n261), .D(n27), .Q(o_kdf_drbg_seed_1_state_value_31_0[21]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[22] ( .CK(clk), .CE(n222), .R(n261), .D(n28), .Q(o_kdf_drbg_seed_1_state_value_31_0[22]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[23] ( .CK(clk), .CE(n222), .R(n261), .D(n29), .Q(o_kdf_drbg_seed_1_state_value_31_0[23]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[24] ( .CK(clk), .CE(n222), .R(n261), .D(n30), .Q(o_kdf_drbg_seed_1_state_value_31_0[24]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[25] ( .CK(clk), .CE(n222), .R(n261), .D(n31), .Q(o_kdf_drbg_seed_1_state_value_31_0[25]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[26] ( .CK(clk), .CE(n222), .R(n261), .D(n32), .Q(o_kdf_drbg_seed_1_state_value_31_0[26]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[27] ( .CK(clk), .CE(n222), .R(n261), .D(n33), .Q(o_kdf_drbg_seed_1_state_value_31_0[27]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[28] ( .CK(clk), .CE(n222), .R(n261), .D(n34), .Q(o_kdf_drbg_seed_1_state_value_31_0[28]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[29] ( .CK(clk), .CE(n222), .R(n261), .D(n35), .Q(o_kdf_drbg_seed_1_state_value_31_0[29]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[30] ( .CK(clk), .CE(n222), .R(n261), .D(n36), .Q(o_kdf_drbg_seed_1_state_value_31_0[30]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_value_31_0_REG[31] ( .CK(clk), .CE(n222), .R(n261), .D(n37), .Q(o_kdf_drbg_seed_1_state_value_31_0[31]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[0] ( .CK(clk), .CE(n221), .R(n261), .D(n6), .Q(o_kdf_drbg_seed_1_state_key_255_224[0]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[1] ( .CK(clk), .CE(n221), .R(n261), .D(n7), .Q(o_kdf_drbg_seed_1_state_key_255_224[1]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[2] ( .CK(clk), .CE(n221), .R(n261), .D(n8), .Q(o_kdf_drbg_seed_1_state_key_255_224[2]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[3] ( .CK(clk), .CE(n221), .R(n261), .D(n9), .Q(o_kdf_drbg_seed_1_state_key_255_224[3]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[4] ( .CK(clk), .CE(n221), .R(n261), .D(n10), .Q(o_kdf_drbg_seed_1_state_key_255_224[4]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[5] ( .CK(clk), .CE(n221), .R(n261), .D(n11), .Q(o_kdf_drbg_seed_1_state_key_255_224[5]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[6] ( .CK(clk), .CE(n221), .R(n261), .D(n12), .Q(o_kdf_drbg_seed_1_state_key_255_224[6]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[7] ( .CK(clk), .CE(n221), .R(n261), .D(n13), .Q(o_kdf_drbg_seed_1_state_key_255_224[7]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[8] ( .CK(clk), .CE(n221), .R(n261), .D(n14), .Q(o_kdf_drbg_seed_1_state_key_255_224[8]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[9] ( .CK(clk), .CE(n221), .R(n261), .D(n15), .Q(o_kdf_drbg_seed_1_state_key_255_224[9]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[10] ( .CK(clk), .CE(n221), .R(n261), .D(n16), .Q(o_kdf_drbg_seed_1_state_key_255_224[10]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[11] ( .CK(clk), .CE(n221), .R(n261), .D(n17), .Q(o_kdf_drbg_seed_1_state_key_255_224[11]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[12] ( .CK(clk), .CE(n221), .R(n261), .D(n18), .Q(o_kdf_drbg_seed_1_state_key_255_224[12]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[13] ( .CK(clk), .CE(n221), .R(n261), .D(n19), .Q(o_kdf_drbg_seed_1_state_key_255_224[13]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[14] ( .CK(clk), .CE(n221), .R(n261), .D(n20), .Q(o_kdf_drbg_seed_1_state_key_255_224[14]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[15] ( .CK(clk), .CE(n221), .R(n261), .D(n21), .Q(o_kdf_drbg_seed_1_state_key_255_224[15]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[16] ( .CK(clk), .CE(n221), .R(n261), .D(n22), .Q(o_kdf_drbg_seed_1_state_key_255_224[16]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[17] ( .CK(clk), .CE(n221), .R(n261), .D(n23), .Q(o_kdf_drbg_seed_1_state_key_255_224[17]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[18] ( .CK(clk), .CE(n221), .R(n261), .D(n24), .Q(o_kdf_drbg_seed_1_state_key_255_224[18]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[19] ( .CK(clk), .CE(n221), .R(n261), .D(n25), .Q(o_kdf_drbg_seed_1_state_key_255_224[19]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[20] ( .CK(clk), .CE(n221), .R(n261), .D(n26), .Q(o_kdf_drbg_seed_1_state_key_255_224[20]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[21] ( .CK(clk), .CE(n221), .R(n261), .D(n27), .Q(o_kdf_drbg_seed_1_state_key_255_224[21]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[22] ( .CK(clk), .CE(n221), .R(n261), .D(n28), .Q(o_kdf_drbg_seed_1_state_key_255_224[22]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[23] ( .CK(clk), .CE(n221), .R(n261), .D(n29), .Q(o_kdf_drbg_seed_1_state_key_255_224[23]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[24] ( .CK(clk), .CE(n221), .R(n261), .D(n30), .Q(o_kdf_drbg_seed_1_state_key_255_224[24]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[25] ( .CK(clk), .CE(n221), .R(n261), .D(n31), .Q(o_kdf_drbg_seed_1_state_key_255_224[25]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[26] ( .CK(clk), .CE(n221), .R(n261), .D(n32), .Q(o_kdf_drbg_seed_1_state_key_255_224[26]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[27] ( .CK(clk), .CE(n221), .R(n261), .D(n33), .Q(o_kdf_drbg_seed_1_state_key_255_224[27]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[28] ( .CK(clk), .CE(n221), .R(n261), .D(n34), .Q(o_kdf_drbg_seed_1_state_key_255_224[28]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[29] ( .CK(clk), .CE(n221), .R(n261), .D(n35), .Q(o_kdf_drbg_seed_1_state_key_255_224[29]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[30] ( .CK(clk), .CE(n221), .R(n261), .D(n36), .Q(o_kdf_drbg_seed_1_state_key_255_224[30]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_255_224_REG[31] ( .CK(clk), .CE(n221), .R(n261), .D(n37), .Q(o_kdf_drbg_seed_1_state_key_255_224[31]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[0] ( .CK(clk), .CE(n220), .R(n261), .D(n6), .Q(o_kdf_drbg_seed_1_state_key_223_192[0]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[1] ( .CK(clk), .CE(n220), .R(n261), .D(n7), .Q(o_kdf_drbg_seed_1_state_key_223_192[1]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[2] ( .CK(clk), .CE(n220), .R(n261), .D(n8), .Q(o_kdf_drbg_seed_1_state_key_223_192[2]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[3] ( .CK(clk), .CE(n220), .R(n261), .D(n9), .Q(o_kdf_drbg_seed_1_state_key_223_192[3]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[4] ( .CK(clk), .CE(n220), .R(n261), .D(n10), .Q(o_kdf_drbg_seed_1_state_key_223_192[4]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[5] ( .CK(clk), .CE(n220), .R(n261), .D(n11), .Q(o_kdf_drbg_seed_1_state_key_223_192[5]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[6] ( .CK(clk), .CE(n220), .R(n261), .D(n12), .Q(o_kdf_drbg_seed_1_state_key_223_192[6]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[7] ( .CK(clk), .CE(n220), .R(n261), .D(n13), .Q(o_kdf_drbg_seed_1_state_key_223_192[7]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[8] ( .CK(clk), .CE(n220), .R(n261), .D(n14), .Q(o_kdf_drbg_seed_1_state_key_223_192[8]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[9] ( .CK(clk), .CE(n220), .R(n261), .D(n15), .Q(o_kdf_drbg_seed_1_state_key_223_192[9]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[10] ( .CK(clk), .CE(n220), .R(n261), .D(n16), .Q(o_kdf_drbg_seed_1_state_key_223_192[10]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[11] ( .CK(clk), .CE(n220), .R(n261), .D(n17), .Q(o_kdf_drbg_seed_1_state_key_223_192[11]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[12] ( .CK(clk), .CE(n220), .R(n261), .D(n18), .Q(o_kdf_drbg_seed_1_state_key_223_192[12]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[13] ( .CK(clk), .CE(n220), .R(n261), .D(n19), .Q(o_kdf_drbg_seed_1_state_key_223_192[13]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[14] ( .CK(clk), .CE(n220), .R(n261), .D(n20), .Q(o_kdf_drbg_seed_1_state_key_223_192[14]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[15] ( .CK(clk), .CE(n220), .R(n261), .D(n21), .Q(o_kdf_drbg_seed_1_state_key_223_192[15]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[16] ( .CK(clk), .CE(n220), .R(n261), .D(n22), .Q(o_kdf_drbg_seed_1_state_key_223_192[16]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[17] ( .CK(clk), .CE(n220), .R(n261), .D(n23), .Q(o_kdf_drbg_seed_1_state_key_223_192[17]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[18] ( .CK(clk), .CE(n220), .R(n261), .D(n24), .Q(o_kdf_drbg_seed_1_state_key_223_192[18]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[19] ( .CK(clk), .CE(n220), .R(n261), .D(n25), .Q(o_kdf_drbg_seed_1_state_key_223_192[19]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[20] ( .CK(clk), .CE(n220), .R(n261), .D(n26), .Q(o_kdf_drbg_seed_1_state_key_223_192[20]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[21] ( .CK(clk), .CE(n220), .R(n261), .D(n27), .Q(o_kdf_drbg_seed_1_state_key_223_192[21]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[22] ( .CK(clk), .CE(n220), .R(n261), .D(n28), .Q(o_kdf_drbg_seed_1_state_key_223_192[22]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[23] ( .CK(clk), .CE(n220), .R(n261), .D(n29), .Q(o_kdf_drbg_seed_1_state_key_223_192[23]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[24] ( .CK(clk), .CE(n220), .R(n261), .D(n30), .Q(o_kdf_drbg_seed_1_state_key_223_192[24]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[25] ( .CK(clk), .CE(n220), .R(n261), .D(n31), .Q(o_kdf_drbg_seed_1_state_key_223_192[25]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[26] ( .CK(clk), .CE(n220), .R(n261), .D(n32), .Q(o_kdf_drbg_seed_1_state_key_223_192[26]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[27] ( .CK(clk), .CE(n220), .R(n261), .D(n33), .Q(o_kdf_drbg_seed_1_state_key_223_192[27]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[28] ( .CK(clk), .CE(n220), .R(n261), .D(n34), .Q(o_kdf_drbg_seed_1_state_key_223_192[28]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[29] ( .CK(clk), .CE(n220), .R(n261), .D(n35), .Q(o_kdf_drbg_seed_1_state_key_223_192[29]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[30] ( .CK(clk), .CE(n220), .R(n261), .D(n36), .Q(o_kdf_drbg_seed_1_state_key_223_192[30]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_223_192_REG[31] ( .CK(clk), .CE(n220), .R(n261), .D(n37), .Q(o_kdf_drbg_seed_1_state_key_223_192[31]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[0] ( .CK(clk), .CE(n219), .R(n261), .D(n6), .Q(o_kdf_drbg_seed_1_state_key_191_160[0]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[1] ( .CK(clk), .CE(n219), .R(n261), .D(n7), .Q(o_kdf_drbg_seed_1_state_key_191_160[1]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[2] ( .CK(clk), .CE(n219), .R(n261), .D(n8), .Q(o_kdf_drbg_seed_1_state_key_191_160[2]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[3] ( .CK(clk), .CE(n219), .R(n261), .D(n9), .Q(o_kdf_drbg_seed_1_state_key_191_160[3]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[4] ( .CK(clk), .CE(n219), .R(n261), .D(n10), .Q(o_kdf_drbg_seed_1_state_key_191_160[4]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[5] ( .CK(clk), .CE(n219), .R(n261), .D(n11), .Q(o_kdf_drbg_seed_1_state_key_191_160[5]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[6] ( .CK(clk), .CE(n219), .R(n261), .D(n12), .Q(o_kdf_drbg_seed_1_state_key_191_160[6]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[7] ( .CK(clk), .CE(n219), .R(n261), .D(n13), .Q(o_kdf_drbg_seed_1_state_key_191_160[7]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[8] ( .CK(clk), .CE(n219), .R(n261), .D(n14), .Q(o_kdf_drbg_seed_1_state_key_191_160[8]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[9] ( .CK(clk), .CE(n219), .R(n261), .D(n15), .Q(o_kdf_drbg_seed_1_state_key_191_160[9]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[10] ( .CK(clk), .CE(n219), .R(n261), .D(n16), .Q(o_kdf_drbg_seed_1_state_key_191_160[10]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[11] ( .CK(clk), .CE(n219), .R(n261), .D(n17), .Q(o_kdf_drbg_seed_1_state_key_191_160[11]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[12] ( .CK(clk), .CE(n219), .R(n261), .D(n18), .Q(o_kdf_drbg_seed_1_state_key_191_160[12]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[13] ( .CK(clk), .CE(n219), .R(n261), .D(n19), .Q(o_kdf_drbg_seed_1_state_key_191_160[13]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[14] ( .CK(clk), .CE(n219), .R(n261), .D(n20), .Q(o_kdf_drbg_seed_1_state_key_191_160[14]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[15] ( .CK(clk), .CE(n219), .R(n261), .D(n21), .Q(o_kdf_drbg_seed_1_state_key_191_160[15]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[16] ( .CK(clk), .CE(n219), .R(n261), .D(n22), .Q(o_kdf_drbg_seed_1_state_key_191_160[16]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[17] ( .CK(clk), .CE(n219), .R(n261), .D(n23), .Q(o_kdf_drbg_seed_1_state_key_191_160[17]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[18] ( .CK(clk), .CE(n219), .R(n261), .D(n24), .Q(o_kdf_drbg_seed_1_state_key_191_160[18]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[19] ( .CK(clk), .CE(n219), .R(n261), .D(n25), .Q(o_kdf_drbg_seed_1_state_key_191_160[19]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[20] ( .CK(clk), .CE(n219), .R(n261), .D(n26), .Q(o_kdf_drbg_seed_1_state_key_191_160[20]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[21] ( .CK(clk), .CE(n219), .R(n261), .D(n27), .Q(o_kdf_drbg_seed_1_state_key_191_160[21]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[22] ( .CK(clk), .CE(n219), .R(n261), .D(n28), .Q(o_kdf_drbg_seed_1_state_key_191_160[22]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[23] ( .CK(clk), .CE(n219), .R(n261), .D(n29), .Q(o_kdf_drbg_seed_1_state_key_191_160[23]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[24] ( .CK(clk), .CE(n219), .R(n261), .D(n30), .Q(o_kdf_drbg_seed_1_state_key_191_160[24]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[25] ( .CK(clk), .CE(n219), .R(n261), .D(n31), .Q(o_kdf_drbg_seed_1_state_key_191_160[25]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[26] ( .CK(clk), .CE(n219), .R(n261), .D(n32), .Q(o_kdf_drbg_seed_1_state_key_191_160[26]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[27] ( .CK(clk), .CE(n219), .R(n261), .D(n33), .Q(o_kdf_drbg_seed_1_state_key_191_160[27]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[28] ( .CK(clk), .CE(n219), .R(n261), .D(n34), .Q(o_kdf_drbg_seed_1_state_key_191_160[28]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[29] ( .CK(clk), .CE(n219), .R(n261), .D(n35), .Q(o_kdf_drbg_seed_1_state_key_191_160[29]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[30] ( .CK(clk), .CE(n219), .R(n261), .D(n36), .Q(o_kdf_drbg_seed_1_state_key_191_160[30]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_191_160_REG[31] ( .CK(clk), .CE(n219), .R(n261), .D(n37), .Q(o_kdf_drbg_seed_1_state_key_191_160[31]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[0] ( .CK(clk), .CE(n218), .R(n261), .D(n6), .Q(o_kdf_drbg_seed_1_state_key_159_128[0]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[1] ( .CK(clk), .CE(n218), .R(n261), .D(n7), .Q(o_kdf_drbg_seed_1_state_key_159_128[1]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[2] ( .CK(clk), .CE(n218), .R(n261), .D(n8), .Q(o_kdf_drbg_seed_1_state_key_159_128[2]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[3] ( .CK(clk), .CE(n218), .R(n261), .D(n9), .Q(o_kdf_drbg_seed_1_state_key_159_128[3]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[4] ( .CK(clk), .CE(n218), .R(n261), .D(n10), .Q(o_kdf_drbg_seed_1_state_key_159_128[4]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[5] ( .CK(clk), .CE(n218), .R(n261), .D(n11), .Q(o_kdf_drbg_seed_1_state_key_159_128[5]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[6] ( .CK(clk), .CE(n218), .R(n261), .D(n12), .Q(o_kdf_drbg_seed_1_state_key_159_128[6]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[7] ( .CK(clk), .CE(n218), .R(n261), .D(n13), .Q(o_kdf_drbg_seed_1_state_key_159_128[7]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[8] ( .CK(clk), .CE(n218), .R(n261), .D(n14), .Q(o_kdf_drbg_seed_1_state_key_159_128[8]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[9] ( .CK(clk), .CE(n218), .R(n261), .D(n15), .Q(o_kdf_drbg_seed_1_state_key_159_128[9]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[10] ( .CK(clk), .CE(n218), .R(n261), .D(n16), .Q(o_kdf_drbg_seed_1_state_key_159_128[10]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[11] ( .CK(clk), .CE(n218), .R(n261), .D(n17), .Q(o_kdf_drbg_seed_1_state_key_159_128[11]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[12] ( .CK(clk), .CE(n218), .R(n261), .D(n18), .Q(o_kdf_drbg_seed_1_state_key_159_128[12]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[13] ( .CK(clk), .CE(n218), .R(n261), .D(n19), .Q(o_kdf_drbg_seed_1_state_key_159_128[13]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[14] ( .CK(clk), .CE(n218), .R(n261), .D(n20), .Q(o_kdf_drbg_seed_1_state_key_159_128[14]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[15] ( .CK(clk), .CE(n218), .R(n261), .D(n21), .Q(o_kdf_drbg_seed_1_state_key_159_128[15]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[16] ( .CK(clk), .CE(n218), .R(n261), .D(n22), .Q(o_kdf_drbg_seed_1_state_key_159_128[16]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[17] ( .CK(clk), .CE(n218), .R(n261), .D(n23), .Q(o_kdf_drbg_seed_1_state_key_159_128[17]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[18] ( .CK(clk), .CE(n218), .R(n261), .D(n24), .Q(o_kdf_drbg_seed_1_state_key_159_128[18]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[19] ( .CK(clk), .CE(n218), .R(n261), .D(n25), .Q(o_kdf_drbg_seed_1_state_key_159_128[19]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[20] ( .CK(clk), .CE(n218), .R(n261), .D(n26), .Q(o_kdf_drbg_seed_1_state_key_159_128[20]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[21] ( .CK(clk), .CE(n218), .R(n261), .D(n27), .Q(o_kdf_drbg_seed_1_state_key_159_128[21]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[22] ( .CK(clk), .CE(n218), .R(n261), .D(n28), .Q(o_kdf_drbg_seed_1_state_key_159_128[22]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[23] ( .CK(clk), .CE(n218), .R(n261), .D(n29), .Q(o_kdf_drbg_seed_1_state_key_159_128[23]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[24] ( .CK(clk), .CE(n218), .R(n261), .D(n30), .Q(o_kdf_drbg_seed_1_state_key_159_128[24]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[25] ( .CK(clk), .CE(n218), .R(n261), .D(n31), .Q(o_kdf_drbg_seed_1_state_key_159_128[25]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[26] ( .CK(clk), .CE(n218), .R(n261), .D(n32), .Q(o_kdf_drbg_seed_1_state_key_159_128[26]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[27] ( .CK(clk), .CE(n218), .R(n261), .D(n33), .Q(o_kdf_drbg_seed_1_state_key_159_128[27]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[28] ( .CK(clk), .CE(n218), .R(n261), .D(n34), .Q(o_kdf_drbg_seed_1_state_key_159_128[28]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[29] ( .CK(clk), .CE(n218), .R(n261), .D(n35), .Q(o_kdf_drbg_seed_1_state_key_159_128[29]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[30] ( .CK(clk), .CE(n218), .R(n261), .D(n36), .Q(o_kdf_drbg_seed_1_state_key_159_128[30]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_159_128_REG[31] ( .CK(clk), .CE(n218), .R(n261), .D(n37), .Q(o_kdf_drbg_seed_1_state_key_159_128[31]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[0] ( .CK(clk), .CE(n217), .R(n261), .D(n6), .Q(o_kdf_drbg_seed_1_state_key_127_96[0]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[1] ( .CK(clk), .CE(n217), .R(n261), .D(n7), .Q(o_kdf_drbg_seed_1_state_key_127_96[1]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[2] ( .CK(clk), .CE(n217), .R(n261), .D(n8), .Q(o_kdf_drbg_seed_1_state_key_127_96[2]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[3] ( .CK(clk), .CE(n217), .R(n261), .D(n9), .Q(o_kdf_drbg_seed_1_state_key_127_96[3]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[4] ( .CK(clk), .CE(n217), .R(n261), .D(n10), .Q(o_kdf_drbg_seed_1_state_key_127_96[4]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[5] ( .CK(clk), .CE(n217), .R(n261), .D(n11), .Q(o_kdf_drbg_seed_1_state_key_127_96[5]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[6] ( .CK(clk), .CE(n217), .R(n261), .D(n12), .Q(o_kdf_drbg_seed_1_state_key_127_96[6]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[7] ( .CK(clk), .CE(n217), .R(n261), .D(n13), .Q(o_kdf_drbg_seed_1_state_key_127_96[7]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[8] ( .CK(clk), .CE(n217), .R(n261), .D(n14), .Q(o_kdf_drbg_seed_1_state_key_127_96[8]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[9] ( .CK(clk), .CE(n217), .R(n261), .D(n15), .Q(o_kdf_drbg_seed_1_state_key_127_96[9]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[10] ( .CK(clk), .CE(n217), .R(n261), .D(n16), .Q(o_kdf_drbg_seed_1_state_key_127_96[10]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[11] ( .CK(clk), .CE(n217), .R(n261), .D(n17), .Q(o_kdf_drbg_seed_1_state_key_127_96[11]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[12] ( .CK(clk), .CE(n217), .R(n261), .D(n18), .Q(o_kdf_drbg_seed_1_state_key_127_96[12]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[13] ( .CK(clk), .CE(n217), .R(n261), .D(n19), .Q(o_kdf_drbg_seed_1_state_key_127_96[13]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[14] ( .CK(clk), .CE(n217), .R(n261), .D(n20), .Q(o_kdf_drbg_seed_1_state_key_127_96[14]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[15] ( .CK(clk), .CE(n217), .R(n261), .D(n21), .Q(o_kdf_drbg_seed_1_state_key_127_96[15]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[16] ( .CK(clk), .CE(n217), .R(n261), .D(n22), .Q(o_kdf_drbg_seed_1_state_key_127_96[16]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[17] ( .CK(clk), .CE(n217), .R(n261), .D(n23), .Q(o_kdf_drbg_seed_1_state_key_127_96[17]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[18] ( .CK(clk), .CE(n217), .R(n261), .D(n24), .Q(o_kdf_drbg_seed_1_state_key_127_96[18]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[19] ( .CK(clk), .CE(n217), .R(n261), .D(n25), .Q(o_kdf_drbg_seed_1_state_key_127_96[19]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[20] ( .CK(clk), .CE(n217), .R(n261), .D(n26), .Q(o_kdf_drbg_seed_1_state_key_127_96[20]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[21] ( .CK(clk), .CE(n217), .R(n261), .D(n27), .Q(o_kdf_drbg_seed_1_state_key_127_96[21]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[22] ( .CK(clk), .CE(n217), .R(n261), .D(n28), .Q(o_kdf_drbg_seed_1_state_key_127_96[22]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[23] ( .CK(clk), .CE(n217), .R(n261), .D(n29), .Q(o_kdf_drbg_seed_1_state_key_127_96[23]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[24] ( .CK(clk), .CE(n217), .R(n261), .D(n30), .Q(o_kdf_drbg_seed_1_state_key_127_96[24]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[25] ( .CK(clk), .CE(n217), .R(n261), .D(n31), .Q(o_kdf_drbg_seed_1_state_key_127_96[25]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[26] ( .CK(clk), .CE(n217), .R(n261), .D(n32), .Q(o_kdf_drbg_seed_1_state_key_127_96[26]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[27] ( .CK(clk), .CE(n217), .R(n261), .D(n33), .Q(o_kdf_drbg_seed_1_state_key_127_96[27]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[28] ( .CK(clk), .CE(n217), .R(n261), .D(n34), .Q(o_kdf_drbg_seed_1_state_key_127_96[28]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[29] ( .CK(clk), .CE(n217), .R(n261), .D(n35), .Q(o_kdf_drbg_seed_1_state_key_127_96[29]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[30] ( .CK(clk), .CE(n217), .R(n261), .D(n36), .Q(o_kdf_drbg_seed_1_state_key_127_96[30]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_127_96_REG[31] ( .CK(clk), .CE(n217), .R(n261), .D(n37), .Q(o_kdf_drbg_seed_1_state_key_127_96[31]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[0] ( .CK(clk), .CE(n216), .R(n261), .D(n6), .Q(o_kdf_drbg_seed_1_state_key_95_64[0]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[1] ( .CK(clk), .CE(n216), .R(n261), .D(n7), .Q(o_kdf_drbg_seed_1_state_key_95_64[1]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[2] ( .CK(clk), .CE(n216), .R(n261), .D(n8), .Q(o_kdf_drbg_seed_1_state_key_95_64[2]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[3] ( .CK(clk), .CE(n216), .R(n261), .D(n9), .Q(o_kdf_drbg_seed_1_state_key_95_64[3]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[4] ( .CK(clk), .CE(n216), .R(n261), .D(n10), .Q(o_kdf_drbg_seed_1_state_key_95_64[4]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[5] ( .CK(clk), .CE(n216), .R(n261), .D(n11), .Q(o_kdf_drbg_seed_1_state_key_95_64[5]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[6] ( .CK(clk), .CE(n216), .R(n261), .D(n12), .Q(o_kdf_drbg_seed_1_state_key_95_64[6]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[7] ( .CK(clk), .CE(n216), .R(n261), .D(n13), .Q(o_kdf_drbg_seed_1_state_key_95_64[7]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[8] ( .CK(clk), .CE(n216), .R(n261), .D(n14), .Q(o_kdf_drbg_seed_1_state_key_95_64[8]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[9] ( .CK(clk), .CE(n216), .R(n261), .D(n15), .Q(o_kdf_drbg_seed_1_state_key_95_64[9]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[10] ( .CK(clk), .CE(n216), .R(n261), .D(n16), .Q(o_kdf_drbg_seed_1_state_key_95_64[10]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[11] ( .CK(clk), .CE(n216), .R(n261), .D(n17), .Q(o_kdf_drbg_seed_1_state_key_95_64[11]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[12] ( .CK(clk), .CE(n216), .R(n261), .D(n18), .Q(o_kdf_drbg_seed_1_state_key_95_64[12]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[13] ( .CK(clk), .CE(n216), .R(n261), .D(n19), .Q(o_kdf_drbg_seed_1_state_key_95_64[13]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[14] ( .CK(clk), .CE(n216), .R(n261), .D(n20), .Q(o_kdf_drbg_seed_1_state_key_95_64[14]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[15] ( .CK(clk), .CE(n216), .R(n261), .D(n21), .Q(o_kdf_drbg_seed_1_state_key_95_64[15]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[16] ( .CK(clk), .CE(n216), .R(n261), .D(n22), .Q(o_kdf_drbg_seed_1_state_key_95_64[16]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[17] ( .CK(clk), .CE(n216), .R(n261), .D(n23), .Q(o_kdf_drbg_seed_1_state_key_95_64[17]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[18] ( .CK(clk), .CE(n216), .R(n261), .D(n24), .Q(o_kdf_drbg_seed_1_state_key_95_64[18]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[19] ( .CK(clk), .CE(n216), .R(n261), .D(n25), .Q(o_kdf_drbg_seed_1_state_key_95_64[19]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[20] ( .CK(clk), .CE(n216), .R(n261), .D(n26), .Q(o_kdf_drbg_seed_1_state_key_95_64[20]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[21] ( .CK(clk), .CE(n216), .R(n261), .D(n27), .Q(o_kdf_drbg_seed_1_state_key_95_64[21]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[22] ( .CK(clk), .CE(n216), .R(n261), .D(n28), .Q(o_kdf_drbg_seed_1_state_key_95_64[22]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[23] ( .CK(clk), .CE(n216), .R(n261), .D(n29), .Q(o_kdf_drbg_seed_1_state_key_95_64[23]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[24] ( .CK(clk), .CE(n216), .R(n261), .D(n30), .Q(o_kdf_drbg_seed_1_state_key_95_64[24]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[25] ( .CK(clk), .CE(n216), .R(n261), .D(n31), .Q(o_kdf_drbg_seed_1_state_key_95_64[25]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[26] ( .CK(clk), .CE(n216), .R(n261), .D(n32), .Q(o_kdf_drbg_seed_1_state_key_95_64[26]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[27] ( .CK(clk), .CE(n216), .R(n261), .D(n33), .Q(o_kdf_drbg_seed_1_state_key_95_64[27]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[28] ( .CK(clk), .CE(n216), .R(n261), .D(n34), .Q(o_kdf_drbg_seed_1_state_key_95_64[28]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[29] ( .CK(clk), .CE(n216), .R(n261), .D(n35), .Q(o_kdf_drbg_seed_1_state_key_95_64[29]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[30] ( .CK(clk), .CE(n216), .R(n261), .D(n36), .Q(o_kdf_drbg_seed_1_state_key_95_64[30]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_95_64_REG[31] ( .CK(clk), .CE(n216), .R(n261), .D(n37), .Q(o_kdf_drbg_seed_1_state_key_95_64[31]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[0] ( .CK(clk), .CE(n215), .R(n261), .D(n6), .Q(o_kdf_drbg_seed_1_state_key_63_32[0]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[1] ( .CK(clk), .CE(n215), .R(n261), .D(n7), .Q(o_kdf_drbg_seed_1_state_key_63_32[1]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[2] ( .CK(clk), .CE(n215), .R(n261), .D(n8), .Q(o_kdf_drbg_seed_1_state_key_63_32[2]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[3] ( .CK(clk), .CE(n215), .R(n261), .D(n9), .Q(o_kdf_drbg_seed_1_state_key_63_32[3]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[4] ( .CK(clk), .CE(n215), .R(n261), .D(n10), .Q(o_kdf_drbg_seed_1_state_key_63_32[4]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[5] ( .CK(clk), .CE(n215), .R(n261), .D(n11), .Q(o_kdf_drbg_seed_1_state_key_63_32[5]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[6] ( .CK(clk), .CE(n215), .R(n261), .D(n12), .Q(o_kdf_drbg_seed_1_state_key_63_32[6]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[7] ( .CK(clk), .CE(n215), .R(n261), .D(n13), .Q(o_kdf_drbg_seed_1_state_key_63_32[7]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[8] ( .CK(clk), .CE(n215), .R(n261), .D(n14), .Q(o_kdf_drbg_seed_1_state_key_63_32[8]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[9] ( .CK(clk), .CE(n215), .R(n261), .D(n15), .Q(o_kdf_drbg_seed_1_state_key_63_32[9]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[10] ( .CK(clk), .CE(n215), .R(n261), .D(n16), .Q(o_kdf_drbg_seed_1_state_key_63_32[10]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[11] ( .CK(clk), .CE(n215), .R(n261), .D(n17), .Q(o_kdf_drbg_seed_1_state_key_63_32[11]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[12] ( .CK(clk), .CE(n215), .R(n261), .D(n18), .Q(o_kdf_drbg_seed_1_state_key_63_32[12]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[13] ( .CK(clk), .CE(n215), .R(n261), .D(n19), .Q(o_kdf_drbg_seed_1_state_key_63_32[13]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[14] ( .CK(clk), .CE(n215), .R(n261), .D(n20), .Q(o_kdf_drbg_seed_1_state_key_63_32[14]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[15] ( .CK(clk), .CE(n215), .R(n261), .D(n21), .Q(o_kdf_drbg_seed_1_state_key_63_32[15]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[16] ( .CK(clk), .CE(n215), .R(n261), .D(n22), .Q(o_kdf_drbg_seed_1_state_key_63_32[16]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[17] ( .CK(clk), .CE(n215), .R(n261), .D(n23), .Q(o_kdf_drbg_seed_1_state_key_63_32[17]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[18] ( .CK(clk), .CE(n215), .R(n261), .D(n24), .Q(o_kdf_drbg_seed_1_state_key_63_32[18]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[19] ( .CK(clk), .CE(n215), .R(n261), .D(n25), .Q(o_kdf_drbg_seed_1_state_key_63_32[19]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[20] ( .CK(clk), .CE(n215), .R(n261), .D(n26), .Q(o_kdf_drbg_seed_1_state_key_63_32[20]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[21] ( .CK(clk), .CE(n215), .R(n261), .D(n27), .Q(o_kdf_drbg_seed_1_state_key_63_32[21]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[22] ( .CK(clk), .CE(n215), .R(n261), .D(n28), .Q(o_kdf_drbg_seed_1_state_key_63_32[22]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[23] ( .CK(clk), .CE(n215), .R(n261), .D(n29), .Q(o_kdf_drbg_seed_1_state_key_63_32[23]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[24] ( .CK(clk), .CE(n215), .R(n261), .D(n30), .Q(o_kdf_drbg_seed_1_state_key_63_32[24]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[25] ( .CK(clk), .CE(n215), .R(n261), .D(n31), .Q(o_kdf_drbg_seed_1_state_key_63_32[25]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[26] ( .CK(clk), .CE(n215), .R(n261), .D(n32), .Q(o_kdf_drbg_seed_1_state_key_63_32[26]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[27] ( .CK(clk), .CE(n215), .R(n261), .D(n33), .Q(o_kdf_drbg_seed_1_state_key_63_32[27]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[28] ( .CK(clk), .CE(n215), .R(n261), .D(n34), .Q(o_kdf_drbg_seed_1_state_key_63_32[28]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[29] ( .CK(clk), .CE(n215), .R(n261), .D(n35), .Q(o_kdf_drbg_seed_1_state_key_63_32[29]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[30] ( .CK(clk), .CE(n215), .R(n261), .D(n36), .Q(o_kdf_drbg_seed_1_state_key_63_32[30]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_63_32_REG[31] ( .CK(clk), .CE(n215), .R(n261), .D(n37), .Q(o_kdf_drbg_seed_1_state_key_63_32[31]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[0] ( .CK(clk), .CE(n214), .R(n261), .D(n6), .Q(o_kdf_drbg_seed_1_state_key_31_0[0]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[1] ( .CK(clk), .CE(n214), .R(n261), .D(n7), .Q(o_kdf_drbg_seed_1_state_key_31_0[1]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[2] ( .CK(clk), .CE(n214), .R(n261), .D(n8), .Q(o_kdf_drbg_seed_1_state_key_31_0[2]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[3] ( .CK(clk), .CE(n214), .R(n261), .D(n9), .Q(o_kdf_drbg_seed_1_state_key_31_0[3]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[4] ( .CK(clk), .CE(n214), .R(n261), .D(n10), .Q(o_kdf_drbg_seed_1_state_key_31_0[4]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[5] ( .CK(clk), .CE(n214), .R(n261), .D(n11), .Q(o_kdf_drbg_seed_1_state_key_31_0[5]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[6] ( .CK(clk), .CE(n214), .R(n261), .D(n12), .Q(o_kdf_drbg_seed_1_state_key_31_0[6]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[7] ( .CK(clk), .CE(n214), .R(n261), .D(n13), .Q(o_kdf_drbg_seed_1_state_key_31_0[7]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[8] ( .CK(clk), .CE(n214), .R(n261), .D(n14), .Q(o_kdf_drbg_seed_1_state_key_31_0[8]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[9] ( .CK(clk), .CE(n214), .R(n261), .D(n15), .Q(o_kdf_drbg_seed_1_state_key_31_0[9]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[10] ( .CK(clk), .CE(n214), .R(n261), .D(n16), .Q(o_kdf_drbg_seed_1_state_key_31_0[10]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[11] ( .CK(clk), .CE(n214), .R(n261), .D(n17), .Q(o_kdf_drbg_seed_1_state_key_31_0[11]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[12] ( .CK(clk), .CE(n214), .R(n261), .D(n18), .Q(o_kdf_drbg_seed_1_state_key_31_0[12]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[13] ( .CK(clk), .CE(n214), .R(n261), .D(n19), .Q(o_kdf_drbg_seed_1_state_key_31_0[13]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[14] ( .CK(clk), .CE(n214), .R(n261), .D(n20), .Q(o_kdf_drbg_seed_1_state_key_31_0[14]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[15] ( .CK(clk), .CE(n214), .R(n261), .D(n21), .Q(o_kdf_drbg_seed_1_state_key_31_0[15]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[16] ( .CK(clk), .CE(n214), .R(n261), .D(n22), .Q(o_kdf_drbg_seed_1_state_key_31_0[16]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[17] ( .CK(clk), .CE(n214), .R(n261), .D(n23), .Q(o_kdf_drbg_seed_1_state_key_31_0[17]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[18] ( .CK(clk), .CE(n214), .R(n261), .D(n24), .Q(o_kdf_drbg_seed_1_state_key_31_0[18]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[19] ( .CK(clk), .CE(n214), .R(n261), .D(n25), .Q(o_kdf_drbg_seed_1_state_key_31_0[19]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[20] ( .CK(clk), .CE(n214), .R(n261), .D(n26), .Q(o_kdf_drbg_seed_1_state_key_31_0[20]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[21] ( .CK(clk), .CE(n214), .R(n261), .D(n27), .Q(o_kdf_drbg_seed_1_state_key_31_0[21]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[22] ( .CK(clk), .CE(n214), .R(n261), .D(n28), .Q(o_kdf_drbg_seed_1_state_key_31_0[22]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[23] ( .CK(clk), .CE(n214), .R(n261), .D(n29), .Q(o_kdf_drbg_seed_1_state_key_31_0[23]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[24] ( .CK(clk), .CE(n214), .R(n261), .D(n30), .Q(o_kdf_drbg_seed_1_state_key_31_0[24]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[25] ( .CK(clk), .CE(n214), .R(n261), .D(n31), .Q(o_kdf_drbg_seed_1_state_key_31_0[25]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[26] ( .CK(clk), .CE(n214), .R(n261), .D(n32), .Q(o_kdf_drbg_seed_1_state_key_31_0[26]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[27] ( .CK(clk), .CE(n214), .R(n261), .D(n33), .Q(o_kdf_drbg_seed_1_state_key_31_0[27]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[28] ( .CK(clk), .CE(n214), .R(n261), .D(n34), .Q(o_kdf_drbg_seed_1_state_key_31_0[28]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[29] ( .CK(clk), .CE(n214), .R(n261), .D(n35), .Q(o_kdf_drbg_seed_1_state_key_31_0[29]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[30] ( .CK(clk), .CE(n214), .R(n261), .D(n36), .Q(o_kdf_drbg_seed_1_state_key_31_0[30]));
Q_FDP4EP \o_kdf_drbg_seed_1_state_key_31_0_REG[31] ( .CK(clk), .CE(n214), .R(n261), .D(n37), .Q(o_kdf_drbg_seed_1_state_key_31_0[31]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_1_REG[0] ( .CK(clk), .CE(n213), .R(n261), .D(n6), .Q(o_kdf_drbg_seed_0_reseed_interval_1[0]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_1_REG[1] ( .CK(clk), .CE(n213), .R(n261), .D(n7), .Q(o_kdf_drbg_seed_0_reseed_interval_1[1]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_1_REG[2] ( .CK(clk), .CE(n213), .R(n261), .D(n8), .Q(o_kdf_drbg_seed_0_reseed_interval_1[2]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_1_REG[3] ( .CK(clk), .CE(n213), .R(n261), .D(n9), .Q(o_kdf_drbg_seed_0_reseed_interval_1[3]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_1_REG[4] ( .CK(clk), .CE(n213), .R(n261), .D(n10), .Q(o_kdf_drbg_seed_0_reseed_interval_1[4]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_1_REG[5] ( .CK(clk), .CE(n213), .R(n261), .D(n11), .Q(o_kdf_drbg_seed_0_reseed_interval_1[5]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_1_REG[6] ( .CK(clk), .CE(n213), .R(n261), .D(n12), .Q(o_kdf_drbg_seed_0_reseed_interval_1[6]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_1_REG[7] ( .CK(clk), .CE(n213), .R(n261), .D(n13), .Q(o_kdf_drbg_seed_0_reseed_interval_1[7]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_1_REG[8] ( .CK(clk), .CE(n213), .R(n261), .D(n14), .Q(o_kdf_drbg_seed_0_reseed_interval_1[8]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_1_REG[9] ( .CK(clk), .CE(n213), .R(n261), .D(n15), .Q(o_kdf_drbg_seed_0_reseed_interval_1[9]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_1_REG[10] ( .CK(clk), .CE(n213), .R(n261), .D(n16), .Q(o_kdf_drbg_seed_0_reseed_interval_1[10]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_1_REG[11] ( .CK(clk), .CE(n213), .R(n261), .D(n17), .Q(o_kdf_drbg_seed_0_reseed_interval_1[11]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_1_REG[12] ( .CK(clk), .CE(n213), .R(n261), .D(n18), .Q(o_kdf_drbg_seed_0_reseed_interval_1[12]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_1_REG[13] ( .CK(clk), .CE(n213), .R(n261), .D(n19), .Q(o_kdf_drbg_seed_0_reseed_interval_1[13]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_1_REG[14] ( .CK(clk), .CE(n213), .R(n261), .D(n20), .Q(o_kdf_drbg_seed_0_reseed_interval_1[14]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_1_REG[15] ( .CK(clk), .CE(n213), .R(n261), .D(n21), .Q(o_kdf_drbg_seed_0_reseed_interval_1[15]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[0] ( .CK(clk), .CE(n212), .R(n261), .D(n6), .Q(o_kdf_drbg_seed_0_reseed_interval_0[0]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[1] ( .CK(clk), .CE(n212), .R(n261), .D(n7), .Q(o_kdf_drbg_seed_0_reseed_interval_0[1]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[2] ( .CK(clk), .CE(n212), .R(n261), .D(n8), .Q(o_kdf_drbg_seed_0_reseed_interval_0[2]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[3] ( .CK(clk), .CE(n212), .R(n261), .D(n9), .Q(o_kdf_drbg_seed_0_reseed_interval_0[3]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[4] ( .CK(clk), .CE(n212), .R(n261), .D(n10), .Q(o_kdf_drbg_seed_0_reseed_interval_0[4]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[5] ( .CK(clk), .CE(n212), .R(n261), .D(n11), .Q(o_kdf_drbg_seed_0_reseed_interval_0[5]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[6] ( .CK(clk), .CE(n212), .R(n261), .D(n12), .Q(o_kdf_drbg_seed_0_reseed_interval_0[6]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[7] ( .CK(clk), .CE(n212), .R(n261), .D(n13), .Q(o_kdf_drbg_seed_0_reseed_interval_0[7]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[8] ( .CK(clk), .CE(n212), .R(n261), .D(n14), .Q(o_kdf_drbg_seed_0_reseed_interval_0[8]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[9] ( .CK(clk), .CE(n212), .R(n261), .D(n15), .Q(o_kdf_drbg_seed_0_reseed_interval_0[9]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[10] ( .CK(clk), .CE(n212), .R(n261), .D(n16), .Q(o_kdf_drbg_seed_0_reseed_interval_0[10]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[11] ( .CK(clk), .CE(n212), .R(n261), .D(n17), .Q(o_kdf_drbg_seed_0_reseed_interval_0[11]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[12] ( .CK(clk), .CE(n212), .R(n261), .D(n18), .Q(o_kdf_drbg_seed_0_reseed_interval_0[12]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[13] ( .CK(clk), .CE(n212), .R(n261), .D(n19), .Q(o_kdf_drbg_seed_0_reseed_interval_0[13]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[14] ( .CK(clk), .CE(n212), .R(n261), .D(n20), .Q(o_kdf_drbg_seed_0_reseed_interval_0[14]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[15] ( .CK(clk), .CE(n212), .R(n261), .D(n21), .Q(o_kdf_drbg_seed_0_reseed_interval_0[15]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[16] ( .CK(clk), .CE(n212), .R(n261), .D(n22), .Q(o_kdf_drbg_seed_0_reseed_interval_0[16]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[17] ( .CK(clk), .CE(n212), .R(n261), .D(n23), .Q(o_kdf_drbg_seed_0_reseed_interval_0[17]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[18] ( .CK(clk), .CE(n212), .R(n261), .D(n24), .Q(o_kdf_drbg_seed_0_reseed_interval_0[18]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[19] ( .CK(clk), .CE(n212), .R(n261), .D(n25), .Q(o_kdf_drbg_seed_0_reseed_interval_0[19]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[20] ( .CK(clk), .CE(n212), .R(n261), .D(n26), .Q(o_kdf_drbg_seed_0_reseed_interval_0[20]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[21] ( .CK(clk), .CE(n212), .R(n261), .D(n27), .Q(o_kdf_drbg_seed_0_reseed_interval_0[21]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[22] ( .CK(clk), .CE(n212), .R(n261), .D(n28), .Q(o_kdf_drbg_seed_0_reseed_interval_0[22]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[23] ( .CK(clk), .CE(n212), .R(n261), .D(n29), .Q(o_kdf_drbg_seed_0_reseed_interval_0[23]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[24] ( .CK(clk), .CE(n212), .R(n261), .D(n30), .Q(o_kdf_drbg_seed_0_reseed_interval_0[24]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[25] ( .CK(clk), .CE(n212), .R(n261), .D(n31), .Q(o_kdf_drbg_seed_0_reseed_interval_0[25]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[26] ( .CK(clk), .CE(n212), .R(n261), .D(n32), .Q(o_kdf_drbg_seed_0_reseed_interval_0[26]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[27] ( .CK(clk), .CE(n212), .R(n261), .D(n33), .Q(o_kdf_drbg_seed_0_reseed_interval_0[27]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[28] ( .CK(clk), .CE(n212), .R(n261), .D(n34), .Q(o_kdf_drbg_seed_0_reseed_interval_0[28]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[29] ( .CK(clk), .CE(n212), .R(n261), .D(n35), .Q(o_kdf_drbg_seed_0_reseed_interval_0[29]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[30] ( .CK(clk), .CE(n212), .R(n261), .D(n36), .Q(o_kdf_drbg_seed_0_reseed_interval_0[30]));
Q_FDP4EP \o_kdf_drbg_seed_0_reseed_interval_0_REG[31] ( .CK(clk), .CE(n212), .R(n261), .D(n37), .Q(o_kdf_drbg_seed_0_reseed_interval_0[31]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[0] ( .CK(clk), .CE(n211), .R(n261), .D(n6), .Q(o_kdf_drbg_seed_0_state_value_127_96[0]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[1] ( .CK(clk), .CE(n211), .R(n261), .D(n7), .Q(o_kdf_drbg_seed_0_state_value_127_96[1]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[2] ( .CK(clk), .CE(n211), .R(n261), .D(n8), .Q(o_kdf_drbg_seed_0_state_value_127_96[2]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[3] ( .CK(clk), .CE(n211), .R(n261), .D(n9), .Q(o_kdf_drbg_seed_0_state_value_127_96[3]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[4] ( .CK(clk), .CE(n211), .R(n261), .D(n10), .Q(o_kdf_drbg_seed_0_state_value_127_96[4]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[5] ( .CK(clk), .CE(n211), .R(n261), .D(n11), .Q(o_kdf_drbg_seed_0_state_value_127_96[5]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[6] ( .CK(clk), .CE(n211), .R(n261), .D(n12), .Q(o_kdf_drbg_seed_0_state_value_127_96[6]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[7] ( .CK(clk), .CE(n211), .R(n261), .D(n13), .Q(o_kdf_drbg_seed_0_state_value_127_96[7]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[8] ( .CK(clk), .CE(n211), .R(n261), .D(n14), .Q(o_kdf_drbg_seed_0_state_value_127_96[8]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[9] ( .CK(clk), .CE(n211), .R(n261), .D(n15), .Q(o_kdf_drbg_seed_0_state_value_127_96[9]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[10] ( .CK(clk), .CE(n211), .R(n261), .D(n16), .Q(o_kdf_drbg_seed_0_state_value_127_96[10]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[11] ( .CK(clk), .CE(n211), .R(n261), .D(n17), .Q(o_kdf_drbg_seed_0_state_value_127_96[11]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[12] ( .CK(clk), .CE(n211), .R(n261), .D(n18), .Q(o_kdf_drbg_seed_0_state_value_127_96[12]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[13] ( .CK(clk), .CE(n211), .R(n261), .D(n19), .Q(o_kdf_drbg_seed_0_state_value_127_96[13]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[14] ( .CK(clk), .CE(n211), .R(n261), .D(n20), .Q(o_kdf_drbg_seed_0_state_value_127_96[14]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[15] ( .CK(clk), .CE(n211), .R(n261), .D(n21), .Q(o_kdf_drbg_seed_0_state_value_127_96[15]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[16] ( .CK(clk), .CE(n211), .R(n261), .D(n22), .Q(o_kdf_drbg_seed_0_state_value_127_96[16]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[17] ( .CK(clk), .CE(n211), .R(n261), .D(n23), .Q(o_kdf_drbg_seed_0_state_value_127_96[17]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[18] ( .CK(clk), .CE(n211), .R(n261), .D(n24), .Q(o_kdf_drbg_seed_0_state_value_127_96[18]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[19] ( .CK(clk), .CE(n211), .R(n261), .D(n25), .Q(o_kdf_drbg_seed_0_state_value_127_96[19]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[20] ( .CK(clk), .CE(n211), .R(n261), .D(n26), .Q(o_kdf_drbg_seed_0_state_value_127_96[20]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[21] ( .CK(clk), .CE(n211), .R(n261), .D(n27), .Q(o_kdf_drbg_seed_0_state_value_127_96[21]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[22] ( .CK(clk), .CE(n211), .R(n261), .D(n28), .Q(o_kdf_drbg_seed_0_state_value_127_96[22]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[23] ( .CK(clk), .CE(n211), .R(n261), .D(n29), .Q(o_kdf_drbg_seed_0_state_value_127_96[23]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[24] ( .CK(clk), .CE(n211), .R(n261), .D(n30), .Q(o_kdf_drbg_seed_0_state_value_127_96[24]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[25] ( .CK(clk), .CE(n211), .R(n261), .D(n31), .Q(o_kdf_drbg_seed_0_state_value_127_96[25]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[26] ( .CK(clk), .CE(n211), .R(n261), .D(n32), .Q(o_kdf_drbg_seed_0_state_value_127_96[26]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[27] ( .CK(clk), .CE(n211), .R(n261), .D(n33), .Q(o_kdf_drbg_seed_0_state_value_127_96[27]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[28] ( .CK(clk), .CE(n211), .R(n261), .D(n34), .Q(o_kdf_drbg_seed_0_state_value_127_96[28]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[29] ( .CK(clk), .CE(n211), .R(n261), .D(n35), .Q(o_kdf_drbg_seed_0_state_value_127_96[29]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[30] ( .CK(clk), .CE(n211), .R(n261), .D(n36), .Q(o_kdf_drbg_seed_0_state_value_127_96[30]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_127_96_REG[31] ( .CK(clk), .CE(n211), .R(n261), .D(n37), .Q(o_kdf_drbg_seed_0_state_value_127_96[31]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[0] ( .CK(clk), .CE(n210), .R(n261), .D(n6), .Q(o_kdf_drbg_seed_0_state_value_95_64[0]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[1] ( .CK(clk), .CE(n210), .R(n261), .D(n7), .Q(o_kdf_drbg_seed_0_state_value_95_64[1]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[2] ( .CK(clk), .CE(n210), .R(n261), .D(n8), .Q(o_kdf_drbg_seed_0_state_value_95_64[2]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[3] ( .CK(clk), .CE(n210), .R(n261), .D(n9), .Q(o_kdf_drbg_seed_0_state_value_95_64[3]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[4] ( .CK(clk), .CE(n210), .R(n261), .D(n10), .Q(o_kdf_drbg_seed_0_state_value_95_64[4]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[5] ( .CK(clk), .CE(n210), .R(n261), .D(n11), .Q(o_kdf_drbg_seed_0_state_value_95_64[5]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[6] ( .CK(clk), .CE(n210), .R(n261), .D(n12), .Q(o_kdf_drbg_seed_0_state_value_95_64[6]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[7] ( .CK(clk), .CE(n210), .R(n261), .D(n13), .Q(o_kdf_drbg_seed_0_state_value_95_64[7]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[8] ( .CK(clk), .CE(n210), .R(n261), .D(n14), .Q(o_kdf_drbg_seed_0_state_value_95_64[8]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[9] ( .CK(clk), .CE(n210), .R(n261), .D(n15), .Q(o_kdf_drbg_seed_0_state_value_95_64[9]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[10] ( .CK(clk), .CE(n210), .R(n261), .D(n16), .Q(o_kdf_drbg_seed_0_state_value_95_64[10]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[11] ( .CK(clk), .CE(n210), .R(n261), .D(n17), .Q(o_kdf_drbg_seed_0_state_value_95_64[11]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[12] ( .CK(clk), .CE(n210), .R(n261), .D(n18), .Q(o_kdf_drbg_seed_0_state_value_95_64[12]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[13] ( .CK(clk), .CE(n210), .R(n261), .D(n19), .Q(o_kdf_drbg_seed_0_state_value_95_64[13]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[14] ( .CK(clk), .CE(n210), .R(n261), .D(n20), .Q(o_kdf_drbg_seed_0_state_value_95_64[14]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[15] ( .CK(clk), .CE(n210), .R(n261), .D(n21), .Q(o_kdf_drbg_seed_0_state_value_95_64[15]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[16] ( .CK(clk), .CE(n210), .R(n261), .D(n22), .Q(o_kdf_drbg_seed_0_state_value_95_64[16]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[17] ( .CK(clk), .CE(n210), .R(n261), .D(n23), .Q(o_kdf_drbg_seed_0_state_value_95_64[17]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[18] ( .CK(clk), .CE(n210), .R(n261), .D(n24), .Q(o_kdf_drbg_seed_0_state_value_95_64[18]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[19] ( .CK(clk), .CE(n210), .R(n261), .D(n25), .Q(o_kdf_drbg_seed_0_state_value_95_64[19]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[20] ( .CK(clk), .CE(n210), .R(n261), .D(n26), .Q(o_kdf_drbg_seed_0_state_value_95_64[20]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[21] ( .CK(clk), .CE(n210), .R(n261), .D(n27), .Q(o_kdf_drbg_seed_0_state_value_95_64[21]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[22] ( .CK(clk), .CE(n210), .R(n261), .D(n28), .Q(o_kdf_drbg_seed_0_state_value_95_64[22]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[23] ( .CK(clk), .CE(n210), .R(n261), .D(n29), .Q(o_kdf_drbg_seed_0_state_value_95_64[23]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[24] ( .CK(clk), .CE(n210), .R(n261), .D(n30), .Q(o_kdf_drbg_seed_0_state_value_95_64[24]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[25] ( .CK(clk), .CE(n210), .R(n261), .D(n31), .Q(o_kdf_drbg_seed_0_state_value_95_64[25]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[26] ( .CK(clk), .CE(n210), .R(n261), .D(n32), .Q(o_kdf_drbg_seed_0_state_value_95_64[26]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[27] ( .CK(clk), .CE(n210), .R(n261), .D(n33), .Q(o_kdf_drbg_seed_0_state_value_95_64[27]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[28] ( .CK(clk), .CE(n210), .R(n261), .D(n34), .Q(o_kdf_drbg_seed_0_state_value_95_64[28]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[29] ( .CK(clk), .CE(n210), .R(n261), .D(n35), .Q(o_kdf_drbg_seed_0_state_value_95_64[29]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[30] ( .CK(clk), .CE(n210), .R(n261), .D(n36), .Q(o_kdf_drbg_seed_0_state_value_95_64[30]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_95_64_REG[31] ( .CK(clk), .CE(n210), .R(n261), .D(n37), .Q(o_kdf_drbg_seed_0_state_value_95_64[31]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[0] ( .CK(clk), .CE(n209), .R(n261), .D(n6), .Q(o_kdf_drbg_seed_0_state_value_63_32[0]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[1] ( .CK(clk), .CE(n209), .R(n261), .D(n7), .Q(o_kdf_drbg_seed_0_state_value_63_32[1]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[2] ( .CK(clk), .CE(n209), .R(n261), .D(n8), .Q(o_kdf_drbg_seed_0_state_value_63_32[2]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[3] ( .CK(clk), .CE(n209), .R(n261), .D(n9), .Q(o_kdf_drbg_seed_0_state_value_63_32[3]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[4] ( .CK(clk), .CE(n209), .R(n261), .D(n10), .Q(o_kdf_drbg_seed_0_state_value_63_32[4]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[5] ( .CK(clk), .CE(n209), .R(n261), .D(n11), .Q(o_kdf_drbg_seed_0_state_value_63_32[5]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[6] ( .CK(clk), .CE(n209), .R(n261), .D(n12), .Q(o_kdf_drbg_seed_0_state_value_63_32[6]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[7] ( .CK(clk), .CE(n209), .R(n261), .D(n13), .Q(o_kdf_drbg_seed_0_state_value_63_32[7]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[8] ( .CK(clk), .CE(n209), .R(n261), .D(n14), .Q(o_kdf_drbg_seed_0_state_value_63_32[8]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[9] ( .CK(clk), .CE(n209), .R(n261), .D(n15), .Q(o_kdf_drbg_seed_0_state_value_63_32[9]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[10] ( .CK(clk), .CE(n209), .R(n261), .D(n16), .Q(o_kdf_drbg_seed_0_state_value_63_32[10]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[11] ( .CK(clk), .CE(n209), .R(n261), .D(n17), .Q(o_kdf_drbg_seed_0_state_value_63_32[11]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[12] ( .CK(clk), .CE(n209), .R(n261), .D(n18), .Q(o_kdf_drbg_seed_0_state_value_63_32[12]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[13] ( .CK(clk), .CE(n209), .R(n261), .D(n19), .Q(o_kdf_drbg_seed_0_state_value_63_32[13]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[14] ( .CK(clk), .CE(n209), .R(n261), .D(n20), .Q(o_kdf_drbg_seed_0_state_value_63_32[14]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[15] ( .CK(clk), .CE(n209), .R(n261), .D(n21), .Q(o_kdf_drbg_seed_0_state_value_63_32[15]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[16] ( .CK(clk), .CE(n209), .R(n261), .D(n22), .Q(o_kdf_drbg_seed_0_state_value_63_32[16]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[17] ( .CK(clk), .CE(n209), .R(n261), .D(n23), .Q(o_kdf_drbg_seed_0_state_value_63_32[17]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[18] ( .CK(clk), .CE(n209), .R(n261), .D(n24), .Q(o_kdf_drbg_seed_0_state_value_63_32[18]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[19] ( .CK(clk), .CE(n209), .R(n261), .D(n25), .Q(o_kdf_drbg_seed_0_state_value_63_32[19]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[20] ( .CK(clk), .CE(n209), .R(n261), .D(n26), .Q(o_kdf_drbg_seed_0_state_value_63_32[20]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[21] ( .CK(clk), .CE(n209), .R(n261), .D(n27), .Q(o_kdf_drbg_seed_0_state_value_63_32[21]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[22] ( .CK(clk), .CE(n209), .R(n261), .D(n28), .Q(o_kdf_drbg_seed_0_state_value_63_32[22]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[23] ( .CK(clk), .CE(n209), .R(n261), .D(n29), .Q(o_kdf_drbg_seed_0_state_value_63_32[23]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[24] ( .CK(clk), .CE(n209), .R(n261), .D(n30), .Q(o_kdf_drbg_seed_0_state_value_63_32[24]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[25] ( .CK(clk), .CE(n209), .R(n261), .D(n31), .Q(o_kdf_drbg_seed_0_state_value_63_32[25]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[26] ( .CK(clk), .CE(n209), .R(n261), .D(n32), .Q(o_kdf_drbg_seed_0_state_value_63_32[26]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[27] ( .CK(clk), .CE(n209), .R(n261), .D(n33), .Q(o_kdf_drbg_seed_0_state_value_63_32[27]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[28] ( .CK(clk), .CE(n209), .R(n261), .D(n34), .Q(o_kdf_drbg_seed_0_state_value_63_32[28]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[29] ( .CK(clk), .CE(n209), .R(n261), .D(n35), .Q(o_kdf_drbg_seed_0_state_value_63_32[29]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[30] ( .CK(clk), .CE(n209), .R(n261), .D(n36), .Q(o_kdf_drbg_seed_0_state_value_63_32[30]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_63_32_REG[31] ( .CK(clk), .CE(n209), .R(n261), .D(n37), .Q(o_kdf_drbg_seed_0_state_value_63_32[31]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[0] ( .CK(clk), .CE(n208), .R(n261), .D(n6), .Q(o_kdf_drbg_seed_0_state_value_31_0[0]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[1] ( .CK(clk), .CE(n208), .R(n261), .D(n7), .Q(o_kdf_drbg_seed_0_state_value_31_0[1]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[2] ( .CK(clk), .CE(n208), .R(n261), .D(n8), .Q(o_kdf_drbg_seed_0_state_value_31_0[2]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[3] ( .CK(clk), .CE(n208), .R(n261), .D(n9), .Q(o_kdf_drbg_seed_0_state_value_31_0[3]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[4] ( .CK(clk), .CE(n208), .R(n261), .D(n10), .Q(o_kdf_drbg_seed_0_state_value_31_0[4]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[5] ( .CK(clk), .CE(n208), .R(n261), .D(n11), .Q(o_kdf_drbg_seed_0_state_value_31_0[5]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[6] ( .CK(clk), .CE(n208), .R(n261), .D(n12), .Q(o_kdf_drbg_seed_0_state_value_31_0[6]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[7] ( .CK(clk), .CE(n208), .R(n261), .D(n13), .Q(o_kdf_drbg_seed_0_state_value_31_0[7]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[8] ( .CK(clk), .CE(n208), .R(n261), .D(n14), .Q(o_kdf_drbg_seed_0_state_value_31_0[8]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[9] ( .CK(clk), .CE(n208), .R(n261), .D(n15), .Q(o_kdf_drbg_seed_0_state_value_31_0[9]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[10] ( .CK(clk), .CE(n208), .R(n261), .D(n16), .Q(o_kdf_drbg_seed_0_state_value_31_0[10]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[11] ( .CK(clk), .CE(n208), .R(n261), .D(n17), .Q(o_kdf_drbg_seed_0_state_value_31_0[11]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[12] ( .CK(clk), .CE(n208), .R(n261), .D(n18), .Q(o_kdf_drbg_seed_0_state_value_31_0[12]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[13] ( .CK(clk), .CE(n208), .R(n261), .D(n19), .Q(o_kdf_drbg_seed_0_state_value_31_0[13]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[14] ( .CK(clk), .CE(n208), .R(n261), .D(n20), .Q(o_kdf_drbg_seed_0_state_value_31_0[14]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[15] ( .CK(clk), .CE(n208), .R(n261), .D(n21), .Q(o_kdf_drbg_seed_0_state_value_31_0[15]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[16] ( .CK(clk), .CE(n208), .R(n261), .D(n22), .Q(o_kdf_drbg_seed_0_state_value_31_0[16]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[17] ( .CK(clk), .CE(n208), .R(n261), .D(n23), .Q(o_kdf_drbg_seed_0_state_value_31_0[17]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[18] ( .CK(clk), .CE(n208), .R(n261), .D(n24), .Q(o_kdf_drbg_seed_0_state_value_31_0[18]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[19] ( .CK(clk), .CE(n208), .R(n261), .D(n25), .Q(o_kdf_drbg_seed_0_state_value_31_0[19]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[20] ( .CK(clk), .CE(n208), .R(n261), .D(n26), .Q(o_kdf_drbg_seed_0_state_value_31_0[20]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[21] ( .CK(clk), .CE(n208), .R(n261), .D(n27), .Q(o_kdf_drbg_seed_0_state_value_31_0[21]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[22] ( .CK(clk), .CE(n208), .R(n261), .D(n28), .Q(o_kdf_drbg_seed_0_state_value_31_0[22]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[23] ( .CK(clk), .CE(n208), .R(n261), .D(n29), .Q(o_kdf_drbg_seed_0_state_value_31_0[23]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[24] ( .CK(clk), .CE(n208), .R(n261), .D(n30), .Q(o_kdf_drbg_seed_0_state_value_31_0[24]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[25] ( .CK(clk), .CE(n208), .R(n261), .D(n31), .Q(o_kdf_drbg_seed_0_state_value_31_0[25]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[26] ( .CK(clk), .CE(n208), .R(n261), .D(n32), .Q(o_kdf_drbg_seed_0_state_value_31_0[26]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[27] ( .CK(clk), .CE(n208), .R(n261), .D(n33), .Q(o_kdf_drbg_seed_0_state_value_31_0[27]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[28] ( .CK(clk), .CE(n208), .R(n261), .D(n34), .Q(o_kdf_drbg_seed_0_state_value_31_0[28]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[29] ( .CK(clk), .CE(n208), .R(n261), .D(n35), .Q(o_kdf_drbg_seed_0_state_value_31_0[29]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[30] ( .CK(clk), .CE(n208), .R(n261), .D(n36), .Q(o_kdf_drbg_seed_0_state_value_31_0[30]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_value_31_0_REG[31] ( .CK(clk), .CE(n208), .R(n261), .D(n37), .Q(o_kdf_drbg_seed_0_state_value_31_0[31]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[0] ( .CK(clk), .CE(n207), .R(n261), .D(n6), .Q(o_kdf_drbg_seed_0_state_key_255_224[0]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[1] ( .CK(clk), .CE(n207), .R(n261), .D(n7), .Q(o_kdf_drbg_seed_0_state_key_255_224[1]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[2] ( .CK(clk), .CE(n207), .R(n261), .D(n8), .Q(o_kdf_drbg_seed_0_state_key_255_224[2]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[3] ( .CK(clk), .CE(n207), .R(n261), .D(n9), .Q(o_kdf_drbg_seed_0_state_key_255_224[3]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[4] ( .CK(clk), .CE(n207), .R(n261), .D(n10), .Q(o_kdf_drbg_seed_0_state_key_255_224[4]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[5] ( .CK(clk), .CE(n207), .R(n261), .D(n11), .Q(o_kdf_drbg_seed_0_state_key_255_224[5]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[6] ( .CK(clk), .CE(n207), .R(n261), .D(n12), .Q(o_kdf_drbg_seed_0_state_key_255_224[6]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[7] ( .CK(clk), .CE(n207), .R(n261), .D(n13), .Q(o_kdf_drbg_seed_0_state_key_255_224[7]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[8] ( .CK(clk), .CE(n207), .R(n261), .D(n14), .Q(o_kdf_drbg_seed_0_state_key_255_224[8]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[9] ( .CK(clk), .CE(n207), .R(n261), .D(n15), .Q(o_kdf_drbg_seed_0_state_key_255_224[9]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[10] ( .CK(clk), .CE(n207), .R(n261), .D(n16), .Q(o_kdf_drbg_seed_0_state_key_255_224[10]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[11] ( .CK(clk), .CE(n207), .R(n261), .D(n17), .Q(o_kdf_drbg_seed_0_state_key_255_224[11]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[12] ( .CK(clk), .CE(n207), .R(n261), .D(n18), .Q(o_kdf_drbg_seed_0_state_key_255_224[12]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[13] ( .CK(clk), .CE(n207), .R(n261), .D(n19), .Q(o_kdf_drbg_seed_0_state_key_255_224[13]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[14] ( .CK(clk), .CE(n207), .R(n261), .D(n20), .Q(o_kdf_drbg_seed_0_state_key_255_224[14]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[15] ( .CK(clk), .CE(n207), .R(n261), .D(n21), .Q(o_kdf_drbg_seed_0_state_key_255_224[15]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[16] ( .CK(clk), .CE(n207), .R(n261), .D(n22), .Q(o_kdf_drbg_seed_0_state_key_255_224[16]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[17] ( .CK(clk), .CE(n207), .R(n261), .D(n23), .Q(o_kdf_drbg_seed_0_state_key_255_224[17]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[18] ( .CK(clk), .CE(n207), .R(n261), .D(n24), .Q(o_kdf_drbg_seed_0_state_key_255_224[18]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[19] ( .CK(clk), .CE(n207), .R(n261), .D(n25), .Q(o_kdf_drbg_seed_0_state_key_255_224[19]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[20] ( .CK(clk), .CE(n207), .R(n261), .D(n26), .Q(o_kdf_drbg_seed_0_state_key_255_224[20]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[21] ( .CK(clk), .CE(n207), .R(n261), .D(n27), .Q(o_kdf_drbg_seed_0_state_key_255_224[21]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[22] ( .CK(clk), .CE(n207), .R(n261), .D(n28), .Q(o_kdf_drbg_seed_0_state_key_255_224[22]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[23] ( .CK(clk), .CE(n207), .R(n261), .D(n29), .Q(o_kdf_drbg_seed_0_state_key_255_224[23]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[24] ( .CK(clk), .CE(n207), .R(n261), .D(n30), .Q(o_kdf_drbg_seed_0_state_key_255_224[24]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[25] ( .CK(clk), .CE(n207), .R(n261), .D(n31), .Q(o_kdf_drbg_seed_0_state_key_255_224[25]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[26] ( .CK(clk), .CE(n207), .R(n261), .D(n32), .Q(o_kdf_drbg_seed_0_state_key_255_224[26]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[27] ( .CK(clk), .CE(n207), .R(n261), .D(n33), .Q(o_kdf_drbg_seed_0_state_key_255_224[27]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[28] ( .CK(clk), .CE(n207), .R(n261), .D(n34), .Q(o_kdf_drbg_seed_0_state_key_255_224[28]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[29] ( .CK(clk), .CE(n207), .R(n261), .D(n35), .Q(o_kdf_drbg_seed_0_state_key_255_224[29]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[30] ( .CK(clk), .CE(n207), .R(n261), .D(n36), .Q(o_kdf_drbg_seed_0_state_key_255_224[30]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_255_224_REG[31] ( .CK(clk), .CE(n207), .R(n261), .D(n37), .Q(o_kdf_drbg_seed_0_state_key_255_224[31]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[0] ( .CK(clk), .CE(n206), .R(n261), .D(n6), .Q(o_kdf_drbg_seed_0_state_key_223_192[0]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[1] ( .CK(clk), .CE(n206), .R(n261), .D(n7), .Q(o_kdf_drbg_seed_0_state_key_223_192[1]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[2] ( .CK(clk), .CE(n206), .R(n261), .D(n8), .Q(o_kdf_drbg_seed_0_state_key_223_192[2]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[3] ( .CK(clk), .CE(n206), .R(n261), .D(n9), .Q(o_kdf_drbg_seed_0_state_key_223_192[3]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[4] ( .CK(clk), .CE(n206), .R(n261), .D(n10), .Q(o_kdf_drbg_seed_0_state_key_223_192[4]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[5] ( .CK(clk), .CE(n206), .R(n261), .D(n11), .Q(o_kdf_drbg_seed_0_state_key_223_192[5]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[6] ( .CK(clk), .CE(n206), .R(n261), .D(n12), .Q(o_kdf_drbg_seed_0_state_key_223_192[6]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[7] ( .CK(clk), .CE(n206), .R(n261), .D(n13), .Q(o_kdf_drbg_seed_0_state_key_223_192[7]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[8] ( .CK(clk), .CE(n206), .R(n261), .D(n14), .Q(o_kdf_drbg_seed_0_state_key_223_192[8]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[9] ( .CK(clk), .CE(n206), .R(n261), .D(n15), .Q(o_kdf_drbg_seed_0_state_key_223_192[9]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[10] ( .CK(clk), .CE(n206), .R(n261), .D(n16), .Q(o_kdf_drbg_seed_0_state_key_223_192[10]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[11] ( .CK(clk), .CE(n206), .R(n261), .D(n17), .Q(o_kdf_drbg_seed_0_state_key_223_192[11]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[12] ( .CK(clk), .CE(n206), .R(n261), .D(n18), .Q(o_kdf_drbg_seed_0_state_key_223_192[12]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[13] ( .CK(clk), .CE(n206), .R(n261), .D(n19), .Q(o_kdf_drbg_seed_0_state_key_223_192[13]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[14] ( .CK(clk), .CE(n206), .R(n261), .D(n20), .Q(o_kdf_drbg_seed_0_state_key_223_192[14]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[15] ( .CK(clk), .CE(n206), .R(n261), .D(n21), .Q(o_kdf_drbg_seed_0_state_key_223_192[15]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[16] ( .CK(clk), .CE(n206), .R(n261), .D(n22), .Q(o_kdf_drbg_seed_0_state_key_223_192[16]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[17] ( .CK(clk), .CE(n206), .R(n261), .D(n23), .Q(o_kdf_drbg_seed_0_state_key_223_192[17]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[18] ( .CK(clk), .CE(n206), .R(n261), .D(n24), .Q(o_kdf_drbg_seed_0_state_key_223_192[18]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[19] ( .CK(clk), .CE(n206), .R(n261), .D(n25), .Q(o_kdf_drbg_seed_0_state_key_223_192[19]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[20] ( .CK(clk), .CE(n206), .R(n261), .D(n26), .Q(o_kdf_drbg_seed_0_state_key_223_192[20]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[21] ( .CK(clk), .CE(n206), .R(n261), .D(n27), .Q(o_kdf_drbg_seed_0_state_key_223_192[21]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[22] ( .CK(clk), .CE(n206), .R(n261), .D(n28), .Q(o_kdf_drbg_seed_0_state_key_223_192[22]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[23] ( .CK(clk), .CE(n206), .R(n261), .D(n29), .Q(o_kdf_drbg_seed_0_state_key_223_192[23]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[24] ( .CK(clk), .CE(n206), .R(n261), .D(n30), .Q(o_kdf_drbg_seed_0_state_key_223_192[24]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[25] ( .CK(clk), .CE(n206), .R(n261), .D(n31), .Q(o_kdf_drbg_seed_0_state_key_223_192[25]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[26] ( .CK(clk), .CE(n206), .R(n261), .D(n32), .Q(o_kdf_drbg_seed_0_state_key_223_192[26]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[27] ( .CK(clk), .CE(n206), .R(n261), .D(n33), .Q(o_kdf_drbg_seed_0_state_key_223_192[27]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[28] ( .CK(clk), .CE(n206), .R(n261), .D(n34), .Q(o_kdf_drbg_seed_0_state_key_223_192[28]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[29] ( .CK(clk), .CE(n206), .R(n261), .D(n35), .Q(o_kdf_drbg_seed_0_state_key_223_192[29]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[30] ( .CK(clk), .CE(n206), .R(n261), .D(n36), .Q(o_kdf_drbg_seed_0_state_key_223_192[30]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_223_192_REG[31] ( .CK(clk), .CE(n206), .R(n261), .D(n37), .Q(o_kdf_drbg_seed_0_state_key_223_192[31]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[0] ( .CK(clk), .CE(n205), .R(n261), .D(n6), .Q(o_kdf_drbg_seed_0_state_key_191_160[0]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[1] ( .CK(clk), .CE(n205), .R(n261), .D(n7), .Q(o_kdf_drbg_seed_0_state_key_191_160[1]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[2] ( .CK(clk), .CE(n205), .R(n261), .D(n8), .Q(o_kdf_drbg_seed_0_state_key_191_160[2]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[3] ( .CK(clk), .CE(n205), .R(n261), .D(n9), .Q(o_kdf_drbg_seed_0_state_key_191_160[3]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[4] ( .CK(clk), .CE(n205), .R(n261), .D(n10), .Q(o_kdf_drbg_seed_0_state_key_191_160[4]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[5] ( .CK(clk), .CE(n205), .R(n261), .D(n11), .Q(o_kdf_drbg_seed_0_state_key_191_160[5]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[6] ( .CK(clk), .CE(n205), .R(n261), .D(n12), .Q(o_kdf_drbg_seed_0_state_key_191_160[6]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[7] ( .CK(clk), .CE(n205), .R(n261), .D(n13), .Q(o_kdf_drbg_seed_0_state_key_191_160[7]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[8] ( .CK(clk), .CE(n205), .R(n261), .D(n14), .Q(o_kdf_drbg_seed_0_state_key_191_160[8]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[9] ( .CK(clk), .CE(n205), .R(n261), .D(n15), .Q(o_kdf_drbg_seed_0_state_key_191_160[9]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[10] ( .CK(clk), .CE(n205), .R(n261), .D(n16), .Q(o_kdf_drbg_seed_0_state_key_191_160[10]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[11] ( .CK(clk), .CE(n205), .R(n261), .D(n17), .Q(o_kdf_drbg_seed_0_state_key_191_160[11]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[12] ( .CK(clk), .CE(n205), .R(n261), .D(n18), .Q(o_kdf_drbg_seed_0_state_key_191_160[12]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[13] ( .CK(clk), .CE(n205), .R(n261), .D(n19), .Q(o_kdf_drbg_seed_0_state_key_191_160[13]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[14] ( .CK(clk), .CE(n205), .R(n261), .D(n20), .Q(o_kdf_drbg_seed_0_state_key_191_160[14]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[15] ( .CK(clk), .CE(n205), .R(n261), .D(n21), .Q(o_kdf_drbg_seed_0_state_key_191_160[15]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[16] ( .CK(clk), .CE(n205), .R(n261), .D(n22), .Q(o_kdf_drbg_seed_0_state_key_191_160[16]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[17] ( .CK(clk), .CE(n205), .R(n261), .D(n23), .Q(o_kdf_drbg_seed_0_state_key_191_160[17]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[18] ( .CK(clk), .CE(n205), .R(n261), .D(n24), .Q(o_kdf_drbg_seed_0_state_key_191_160[18]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[19] ( .CK(clk), .CE(n205), .R(n261), .D(n25), .Q(o_kdf_drbg_seed_0_state_key_191_160[19]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[20] ( .CK(clk), .CE(n205), .R(n261), .D(n26), .Q(o_kdf_drbg_seed_0_state_key_191_160[20]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[21] ( .CK(clk), .CE(n205), .R(n261), .D(n27), .Q(o_kdf_drbg_seed_0_state_key_191_160[21]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[22] ( .CK(clk), .CE(n205), .R(n261), .D(n28), .Q(o_kdf_drbg_seed_0_state_key_191_160[22]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[23] ( .CK(clk), .CE(n205), .R(n261), .D(n29), .Q(o_kdf_drbg_seed_0_state_key_191_160[23]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[24] ( .CK(clk), .CE(n205), .R(n261), .D(n30), .Q(o_kdf_drbg_seed_0_state_key_191_160[24]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[25] ( .CK(clk), .CE(n205), .R(n261), .D(n31), .Q(o_kdf_drbg_seed_0_state_key_191_160[25]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[26] ( .CK(clk), .CE(n205), .R(n261), .D(n32), .Q(o_kdf_drbg_seed_0_state_key_191_160[26]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[27] ( .CK(clk), .CE(n205), .R(n261), .D(n33), .Q(o_kdf_drbg_seed_0_state_key_191_160[27]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[28] ( .CK(clk), .CE(n205), .R(n261), .D(n34), .Q(o_kdf_drbg_seed_0_state_key_191_160[28]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[29] ( .CK(clk), .CE(n205), .R(n261), .D(n35), .Q(o_kdf_drbg_seed_0_state_key_191_160[29]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[30] ( .CK(clk), .CE(n205), .R(n261), .D(n36), .Q(o_kdf_drbg_seed_0_state_key_191_160[30]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_191_160_REG[31] ( .CK(clk), .CE(n205), .R(n261), .D(n37), .Q(o_kdf_drbg_seed_0_state_key_191_160[31]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[0] ( .CK(clk), .CE(n204), .R(n261), .D(n6), .Q(o_kdf_drbg_seed_0_state_key_159_128[0]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[1] ( .CK(clk), .CE(n204), .R(n261), .D(n7), .Q(o_kdf_drbg_seed_0_state_key_159_128[1]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[2] ( .CK(clk), .CE(n204), .R(n261), .D(n8), .Q(o_kdf_drbg_seed_0_state_key_159_128[2]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[3] ( .CK(clk), .CE(n204), .R(n261), .D(n9), .Q(o_kdf_drbg_seed_0_state_key_159_128[3]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[4] ( .CK(clk), .CE(n204), .R(n261), .D(n10), .Q(o_kdf_drbg_seed_0_state_key_159_128[4]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[5] ( .CK(clk), .CE(n204), .R(n261), .D(n11), .Q(o_kdf_drbg_seed_0_state_key_159_128[5]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[6] ( .CK(clk), .CE(n204), .R(n261), .D(n12), .Q(o_kdf_drbg_seed_0_state_key_159_128[6]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[7] ( .CK(clk), .CE(n204), .R(n261), .D(n13), .Q(o_kdf_drbg_seed_0_state_key_159_128[7]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[8] ( .CK(clk), .CE(n204), .R(n261), .D(n14), .Q(o_kdf_drbg_seed_0_state_key_159_128[8]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[9] ( .CK(clk), .CE(n204), .R(n261), .D(n15), .Q(o_kdf_drbg_seed_0_state_key_159_128[9]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[10] ( .CK(clk), .CE(n204), .R(n261), .D(n16), .Q(o_kdf_drbg_seed_0_state_key_159_128[10]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[11] ( .CK(clk), .CE(n204), .R(n261), .D(n17), .Q(o_kdf_drbg_seed_0_state_key_159_128[11]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[12] ( .CK(clk), .CE(n204), .R(n261), .D(n18), .Q(o_kdf_drbg_seed_0_state_key_159_128[12]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[13] ( .CK(clk), .CE(n204), .R(n261), .D(n19), .Q(o_kdf_drbg_seed_0_state_key_159_128[13]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[14] ( .CK(clk), .CE(n204), .R(n261), .D(n20), .Q(o_kdf_drbg_seed_0_state_key_159_128[14]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[15] ( .CK(clk), .CE(n204), .R(n261), .D(n21), .Q(o_kdf_drbg_seed_0_state_key_159_128[15]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[16] ( .CK(clk), .CE(n204), .R(n261), .D(n22), .Q(o_kdf_drbg_seed_0_state_key_159_128[16]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[17] ( .CK(clk), .CE(n204), .R(n261), .D(n23), .Q(o_kdf_drbg_seed_0_state_key_159_128[17]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[18] ( .CK(clk), .CE(n204), .R(n261), .D(n24), .Q(o_kdf_drbg_seed_0_state_key_159_128[18]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[19] ( .CK(clk), .CE(n204), .R(n261), .D(n25), .Q(o_kdf_drbg_seed_0_state_key_159_128[19]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[20] ( .CK(clk), .CE(n204), .R(n261), .D(n26), .Q(o_kdf_drbg_seed_0_state_key_159_128[20]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[21] ( .CK(clk), .CE(n204), .R(n261), .D(n27), .Q(o_kdf_drbg_seed_0_state_key_159_128[21]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[22] ( .CK(clk), .CE(n204), .R(n261), .D(n28), .Q(o_kdf_drbg_seed_0_state_key_159_128[22]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[23] ( .CK(clk), .CE(n204), .R(n261), .D(n29), .Q(o_kdf_drbg_seed_0_state_key_159_128[23]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[24] ( .CK(clk), .CE(n204), .R(n261), .D(n30), .Q(o_kdf_drbg_seed_0_state_key_159_128[24]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[25] ( .CK(clk), .CE(n204), .R(n261), .D(n31), .Q(o_kdf_drbg_seed_0_state_key_159_128[25]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[26] ( .CK(clk), .CE(n204), .R(n261), .D(n32), .Q(o_kdf_drbg_seed_0_state_key_159_128[26]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[27] ( .CK(clk), .CE(n204), .R(n261), .D(n33), .Q(o_kdf_drbg_seed_0_state_key_159_128[27]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[28] ( .CK(clk), .CE(n204), .R(n261), .D(n34), .Q(o_kdf_drbg_seed_0_state_key_159_128[28]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[29] ( .CK(clk), .CE(n204), .R(n261), .D(n35), .Q(o_kdf_drbg_seed_0_state_key_159_128[29]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[30] ( .CK(clk), .CE(n204), .R(n261), .D(n36), .Q(o_kdf_drbg_seed_0_state_key_159_128[30]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_159_128_REG[31] ( .CK(clk), .CE(n204), .R(n261), .D(n37), .Q(o_kdf_drbg_seed_0_state_key_159_128[31]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[0] ( .CK(clk), .CE(n203), .R(n261), .D(n6), .Q(o_kdf_drbg_seed_0_state_key_127_96[0]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[1] ( .CK(clk), .CE(n203), .R(n261), .D(n7), .Q(o_kdf_drbg_seed_0_state_key_127_96[1]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[2] ( .CK(clk), .CE(n203), .R(n261), .D(n8), .Q(o_kdf_drbg_seed_0_state_key_127_96[2]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[3] ( .CK(clk), .CE(n203), .R(n261), .D(n9), .Q(o_kdf_drbg_seed_0_state_key_127_96[3]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[4] ( .CK(clk), .CE(n203), .R(n261), .D(n10), .Q(o_kdf_drbg_seed_0_state_key_127_96[4]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[5] ( .CK(clk), .CE(n203), .R(n261), .D(n11), .Q(o_kdf_drbg_seed_0_state_key_127_96[5]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[6] ( .CK(clk), .CE(n203), .R(n261), .D(n12), .Q(o_kdf_drbg_seed_0_state_key_127_96[6]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[7] ( .CK(clk), .CE(n203), .R(n261), .D(n13), .Q(o_kdf_drbg_seed_0_state_key_127_96[7]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[8] ( .CK(clk), .CE(n203), .R(n261), .D(n14), .Q(o_kdf_drbg_seed_0_state_key_127_96[8]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[9] ( .CK(clk), .CE(n203), .R(n261), .D(n15), .Q(o_kdf_drbg_seed_0_state_key_127_96[9]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[10] ( .CK(clk), .CE(n203), .R(n261), .D(n16), .Q(o_kdf_drbg_seed_0_state_key_127_96[10]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[11] ( .CK(clk), .CE(n203), .R(n261), .D(n17), .Q(o_kdf_drbg_seed_0_state_key_127_96[11]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[12] ( .CK(clk), .CE(n203), .R(n261), .D(n18), .Q(o_kdf_drbg_seed_0_state_key_127_96[12]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[13] ( .CK(clk), .CE(n203), .R(n261), .D(n19), .Q(o_kdf_drbg_seed_0_state_key_127_96[13]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[14] ( .CK(clk), .CE(n203), .R(n261), .D(n20), .Q(o_kdf_drbg_seed_0_state_key_127_96[14]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[15] ( .CK(clk), .CE(n203), .R(n261), .D(n21), .Q(o_kdf_drbg_seed_0_state_key_127_96[15]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[16] ( .CK(clk), .CE(n203), .R(n261), .D(n22), .Q(o_kdf_drbg_seed_0_state_key_127_96[16]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[17] ( .CK(clk), .CE(n203), .R(n261), .D(n23), .Q(o_kdf_drbg_seed_0_state_key_127_96[17]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[18] ( .CK(clk), .CE(n203), .R(n261), .D(n24), .Q(o_kdf_drbg_seed_0_state_key_127_96[18]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[19] ( .CK(clk), .CE(n203), .R(n261), .D(n25), .Q(o_kdf_drbg_seed_0_state_key_127_96[19]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[20] ( .CK(clk), .CE(n203), .R(n261), .D(n26), .Q(o_kdf_drbg_seed_0_state_key_127_96[20]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[21] ( .CK(clk), .CE(n203), .R(n261), .D(n27), .Q(o_kdf_drbg_seed_0_state_key_127_96[21]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[22] ( .CK(clk), .CE(n203), .R(n261), .D(n28), .Q(o_kdf_drbg_seed_0_state_key_127_96[22]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[23] ( .CK(clk), .CE(n203), .R(n261), .D(n29), .Q(o_kdf_drbg_seed_0_state_key_127_96[23]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[24] ( .CK(clk), .CE(n203), .R(n261), .D(n30), .Q(o_kdf_drbg_seed_0_state_key_127_96[24]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[25] ( .CK(clk), .CE(n203), .R(n261), .D(n31), .Q(o_kdf_drbg_seed_0_state_key_127_96[25]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[26] ( .CK(clk), .CE(n203), .R(n261), .D(n32), .Q(o_kdf_drbg_seed_0_state_key_127_96[26]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[27] ( .CK(clk), .CE(n203), .R(n261), .D(n33), .Q(o_kdf_drbg_seed_0_state_key_127_96[27]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[28] ( .CK(clk), .CE(n203), .R(n261), .D(n34), .Q(o_kdf_drbg_seed_0_state_key_127_96[28]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[29] ( .CK(clk), .CE(n203), .R(n261), .D(n35), .Q(o_kdf_drbg_seed_0_state_key_127_96[29]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[30] ( .CK(clk), .CE(n203), .R(n261), .D(n36), .Q(o_kdf_drbg_seed_0_state_key_127_96[30]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_127_96_REG[31] ( .CK(clk), .CE(n203), .R(n261), .D(n37), .Q(o_kdf_drbg_seed_0_state_key_127_96[31]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[0] ( .CK(clk), .CE(n202), .R(n261), .D(n6), .Q(o_kdf_drbg_seed_0_state_key_95_64[0]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[1] ( .CK(clk), .CE(n202), .R(n261), .D(n7), .Q(o_kdf_drbg_seed_0_state_key_95_64[1]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[2] ( .CK(clk), .CE(n202), .R(n261), .D(n8), .Q(o_kdf_drbg_seed_0_state_key_95_64[2]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[3] ( .CK(clk), .CE(n202), .R(n261), .D(n9), .Q(o_kdf_drbg_seed_0_state_key_95_64[3]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[4] ( .CK(clk), .CE(n202), .R(n261), .D(n10), .Q(o_kdf_drbg_seed_0_state_key_95_64[4]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[5] ( .CK(clk), .CE(n202), .R(n261), .D(n11), .Q(o_kdf_drbg_seed_0_state_key_95_64[5]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[6] ( .CK(clk), .CE(n202), .R(n261), .D(n12), .Q(o_kdf_drbg_seed_0_state_key_95_64[6]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[7] ( .CK(clk), .CE(n202), .R(n261), .D(n13), .Q(o_kdf_drbg_seed_0_state_key_95_64[7]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[8] ( .CK(clk), .CE(n202), .R(n261), .D(n14), .Q(o_kdf_drbg_seed_0_state_key_95_64[8]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[9] ( .CK(clk), .CE(n202), .R(n261), .D(n15), .Q(o_kdf_drbg_seed_0_state_key_95_64[9]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[10] ( .CK(clk), .CE(n202), .R(n261), .D(n16), .Q(o_kdf_drbg_seed_0_state_key_95_64[10]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[11] ( .CK(clk), .CE(n202), .R(n261), .D(n17), .Q(o_kdf_drbg_seed_0_state_key_95_64[11]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[12] ( .CK(clk), .CE(n202), .R(n261), .D(n18), .Q(o_kdf_drbg_seed_0_state_key_95_64[12]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[13] ( .CK(clk), .CE(n202), .R(n261), .D(n19), .Q(o_kdf_drbg_seed_0_state_key_95_64[13]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[14] ( .CK(clk), .CE(n202), .R(n261), .D(n20), .Q(o_kdf_drbg_seed_0_state_key_95_64[14]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[15] ( .CK(clk), .CE(n202), .R(n261), .D(n21), .Q(o_kdf_drbg_seed_0_state_key_95_64[15]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[16] ( .CK(clk), .CE(n202), .R(n261), .D(n22), .Q(o_kdf_drbg_seed_0_state_key_95_64[16]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[17] ( .CK(clk), .CE(n202), .R(n261), .D(n23), .Q(o_kdf_drbg_seed_0_state_key_95_64[17]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[18] ( .CK(clk), .CE(n202), .R(n261), .D(n24), .Q(o_kdf_drbg_seed_0_state_key_95_64[18]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[19] ( .CK(clk), .CE(n202), .R(n261), .D(n25), .Q(o_kdf_drbg_seed_0_state_key_95_64[19]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[20] ( .CK(clk), .CE(n202), .R(n261), .D(n26), .Q(o_kdf_drbg_seed_0_state_key_95_64[20]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[21] ( .CK(clk), .CE(n202), .R(n261), .D(n27), .Q(o_kdf_drbg_seed_0_state_key_95_64[21]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[22] ( .CK(clk), .CE(n202), .R(n261), .D(n28), .Q(o_kdf_drbg_seed_0_state_key_95_64[22]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[23] ( .CK(clk), .CE(n202), .R(n261), .D(n29), .Q(o_kdf_drbg_seed_0_state_key_95_64[23]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[24] ( .CK(clk), .CE(n202), .R(n261), .D(n30), .Q(o_kdf_drbg_seed_0_state_key_95_64[24]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[25] ( .CK(clk), .CE(n202), .R(n261), .D(n31), .Q(o_kdf_drbg_seed_0_state_key_95_64[25]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[26] ( .CK(clk), .CE(n202), .R(n261), .D(n32), .Q(o_kdf_drbg_seed_0_state_key_95_64[26]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[27] ( .CK(clk), .CE(n202), .R(n261), .D(n33), .Q(o_kdf_drbg_seed_0_state_key_95_64[27]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[28] ( .CK(clk), .CE(n202), .R(n261), .D(n34), .Q(o_kdf_drbg_seed_0_state_key_95_64[28]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[29] ( .CK(clk), .CE(n202), .R(n261), .D(n35), .Q(o_kdf_drbg_seed_0_state_key_95_64[29]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[30] ( .CK(clk), .CE(n202), .R(n261), .D(n36), .Q(o_kdf_drbg_seed_0_state_key_95_64[30]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_95_64_REG[31] ( .CK(clk), .CE(n202), .R(n261), .D(n37), .Q(o_kdf_drbg_seed_0_state_key_95_64[31]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[0] ( .CK(clk), .CE(n201), .R(n261), .D(n6), .Q(o_kdf_drbg_seed_0_state_key_63_32[0]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[1] ( .CK(clk), .CE(n201), .R(n261), .D(n7), .Q(o_kdf_drbg_seed_0_state_key_63_32[1]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[2] ( .CK(clk), .CE(n201), .R(n261), .D(n8), .Q(o_kdf_drbg_seed_0_state_key_63_32[2]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[3] ( .CK(clk), .CE(n201), .R(n261), .D(n9), .Q(o_kdf_drbg_seed_0_state_key_63_32[3]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[4] ( .CK(clk), .CE(n201), .R(n261), .D(n10), .Q(o_kdf_drbg_seed_0_state_key_63_32[4]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[5] ( .CK(clk), .CE(n201), .R(n261), .D(n11), .Q(o_kdf_drbg_seed_0_state_key_63_32[5]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[6] ( .CK(clk), .CE(n201), .R(n261), .D(n12), .Q(o_kdf_drbg_seed_0_state_key_63_32[6]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[7] ( .CK(clk), .CE(n201), .R(n261), .D(n13), .Q(o_kdf_drbg_seed_0_state_key_63_32[7]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[8] ( .CK(clk), .CE(n201), .R(n261), .D(n14), .Q(o_kdf_drbg_seed_0_state_key_63_32[8]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[9] ( .CK(clk), .CE(n201), .R(n261), .D(n15), .Q(o_kdf_drbg_seed_0_state_key_63_32[9]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[10] ( .CK(clk), .CE(n201), .R(n261), .D(n16), .Q(o_kdf_drbg_seed_0_state_key_63_32[10]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[11] ( .CK(clk), .CE(n201), .R(n261), .D(n17), .Q(o_kdf_drbg_seed_0_state_key_63_32[11]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[12] ( .CK(clk), .CE(n201), .R(n261), .D(n18), .Q(o_kdf_drbg_seed_0_state_key_63_32[12]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[13] ( .CK(clk), .CE(n201), .R(n261), .D(n19), .Q(o_kdf_drbg_seed_0_state_key_63_32[13]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[14] ( .CK(clk), .CE(n201), .R(n261), .D(n20), .Q(o_kdf_drbg_seed_0_state_key_63_32[14]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[15] ( .CK(clk), .CE(n201), .R(n261), .D(n21), .Q(o_kdf_drbg_seed_0_state_key_63_32[15]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[16] ( .CK(clk), .CE(n201), .R(n261), .D(n22), .Q(o_kdf_drbg_seed_0_state_key_63_32[16]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[17] ( .CK(clk), .CE(n201), .R(n261), .D(n23), .Q(o_kdf_drbg_seed_0_state_key_63_32[17]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[18] ( .CK(clk), .CE(n201), .R(n261), .D(n24), .Q(o_kdf_drbg_seed_0_state_key_63_32[18]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[19] ( .CK(clk), .CE(n201), .R(n261), .D(n25), .Q(o_kdf_drbg_seed_0_state_key_63_32[19]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[20] ( .CK(clk), .CE(n201), .R(n261), .D(n26), .Q(o_kdf_drbg_seed_0_state_key_63_32[20]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[21] ( .CK(clk), .CE(n201), .R(n261), .D(n27), .Q(o_kdf_drbg_seed_0_state_key_63_32[21]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[22] ( .CK(clk), .CE(n201), .R(n261), .D(n28), .Q(o_kdf_drbg_seed_0_state_key_63_32[22]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[23] ( .CK(clk), .CE(n201), .R(n261), .D(n29), .Q(o_kdf_drbg_seed_0_state_key_63_32[23]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[24] ( .CK(clk), .CE(n201), .R(n261), .D(n30), .Q(o_kdf_drbg_seed_0_state_key_63_32[24]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[25] ( .CK(clk), .CE(n201), .R(n261), .D(n31), .Q(o_kdf_drbg_seed_0_state_key_63_32[25]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[26] ( .CK(clk), .CE(n201), .R(n261), .D(n32), .Q(o_kdf_drbg_seed_0_state_key_63_32[26]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[27] ( .CK(clk), .CE(n201), .R(n261), .D(n33), .Q(o_kdf_drbg_seed_0_state_key_63_32[27]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[28] ( .CK(clk), .CE(n201), .R(n261), .D(n34), .Q(o_kdf_drbg_seed_0_state_key_63_32[28]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[29] ( .CK(clk), .CE(n201), .R(n261), .D(n35), .Q(o_kdf_drbg_seed_0_state_key_63_32[29]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[30] ( .CK(clk), .CE(n201), .R(n261), .D(n36), .Q(o_kdf_drbg_seed_0_state_key_63_32[30]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_63_32_REG[31] ( .CK(clk), .CE(n201), .R(n261), .D(n37), .Q(o_kdf_drbg_seed_0_state_key_63_32[31]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[0] ( .CK(clk), .CE(n200), .R(n261), .D(n6), .Q(o_kdf_drbg_seed_0_state_key_31_0[0]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[1] ( .CK(clk), .CE(n200), .R(n261), .D(n7), .Q(o_kdf_drbg_seed_0_state_key_31_0[1]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[2] ( .CK(clk), .CE(n200), .R(n261), .D(n8), .Q(o_kdf_drbg_seed_0_state_key_31_0[2]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[3] ( .CK(clk), .CE(n200), .R(n261), .D(n9), .Q(o_kdf_drbg_seed_0_state_key_31_0[3]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[4] ( .CK(clk), .CE(n200), .R(n261), .D(n10), .Q(o_kdf_drbg_seed_0_state_key_31_0[4]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[5] ( .CK(clk), .CE(n200), .R(n261), .D(n11), .Q(o_kdf_drbg_seed_0_state_key_31_0[5]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[6] ( .CK(clk), .CE(n200), .R(n261), .D(n12), .Q(o_kdf_drbg_seed_0_state_key_31_0[6]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[7] ( .CK(clk), .CE(n200), .R(n261), .D(n13), .Q(o_kdf_drbg_seed_0_state_key_31_0[7]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[8] ( .CK(clk), .CE(n200), .R(n261), .D(n14), .Q(o_kdf_drbg_seed_0_state_key_31_0[8]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[9] ( .CK(clk), .CE(n200), .R(n261), .D(n15), .Q(o_kdf_drbg_seed_0_state_key_31_0[9]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[10] ( .CK(clk), .CE(n200), .R(n261), .D(n16), .Q(o_kdf_drbg_seed_0_state_key_31_0[10]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[11] ( .CK(clk), .CE(n200), .R(n261), .D(n17), .Q(o_kdf_drbg_seed_0_state_key_31_0[11]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[12] ( .CK(clk), .CE(n200), .R(n261), .D(n18), .Q(o_kdf_drbg_seed_0_state_key_31_0[12]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[13] ( .CK(clk), .CE(n200), .R(n261), .D(n19), .Q(o_kdf_drbg_seed_0_state_key_31_0[13]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[14] ( .CK(clk), .CE(n200), .R(n261), .D(n20), .Q(o_kdf_drbg_seed_0_state_key_31_0[14]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[15] ( .CK(clk), .CE(n200), .R(n261), .D(n21), .Q(o_kdf_drbg_seed_0_state_key_31_0[15]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[16] ( .CK(clk), .CE(n200), .R(n261), .D(n22), .Q(o_kdf_drbg_seed_0_state_key_31_0[16]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[17] ( .CK(clk), .CE(n200), .R(n261), .D(n23), .Q(o_kdf_drbg_seed_0_state_key_31_0[17]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[18] ( .CK(clk), .CE(n200), .R(n261), .D(n24), .Q(o_kdf_drbg_seed_0_state_key_31_0[18]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[19] ( .CK(clk), .CE(n200), .R(n261), .D(n25), .Q(o_kdf_drbg_seed_0_state_key_31_0[19]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[20] ( .CK(clk), .CE(n200), .R(n261), .D(n26), .Q(o_kdf_drbg_seed_0_state_key_31_0[20]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[21] ( .CK(clk), .CE(n200), .R(n261), .D(n27), .Q(o_kdf_drbg_seed_0_state_key_31_0[21]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[22] ( .CK(clk), .CE(n200), .R(n261), .D(n28), .Q(o_kdf_drbg_seed_0_state_key_31_0[22]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[23] ( .CK(clk), .CE(n200), .R(n261), .D(n29), .Q(o_kdf_drbg_seed_0_state_key_31_0[23]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[24] ( .CK(clk), .CE(n200), .R(n261), .D(n30), .Q(o_kdf_drbg_seed_0_state_key_31_0[24]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[25] ( .CK(clk), .CE(n200), .R(n261), .D(n31), .Q(o_kdf_drbg_seed_0_state_key_31_0[25]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[26] ( .CK(clk), .CE(n200), .R(n261), .D(n32), .Q(o_kdf_drbg_seed_0_state_key_31_0[26]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[27] ( .CK(clk), .CE(n200), .R(n261), .D(n33), .Q(o_kdf_drbg_seed_0_state_key_31_0[27]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[28] ( .CK(clk), .CE(n200), .R(n261), .D(n34), .Q(o_kdf_drbg_seed_0_state_key_31_0[28]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[29] ( .CK(clk), .CE(n200), .R(n261), .D(n35), .Q(o_kdf_drbg_seed_0_state_key_31_0[29]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[30] ( .CK(clk), .CE(n200), .R(n261), .D(n36), .Q(o_kdf_drbg_seed_0_state_key_31_0[30]));
Q_FDP4EP \o_kdf_drbg_seed_0_state_key_31_0_REG[31] ( .CK(clk), .CE(n200), .R(n261), .D(n37), .Q(o_kdf_drbg_seed_0_state_key_31_0[31]));
Q_FDP4EP \o_kdf_drbg_ctrl_REG[0] ( .CK(clk), .CE(n199), .R(n261), .D(n6), .Q(o_kdf_drbg_ctrl[0]));
Q_FDP4EP \o_kdf_drbg_ctrl_REG[1] ( .CK(clk), .CE(n199), .R(n261), .D(n7), .Q(o_kdf_drbg_ctrl[1]));
Q_FDP4EP \o_label7_data0_REG[0] ( .CK(clk), .CE(n198), .R(n261), .D(n6), .Q(o_label7_data0[0]));
Q_FDP4EP \o_label7_data0_REG[1] ( .CK(clk), .CE(n198), .R(n261), .D(n7), .Q(o_label7_data0[1]));
Q_FDP4EP \o_label7_data0_REG[2] ( .CK(clk), .CE(n198), .R(n261), .D(n8), .Q(o_label7_data0[2]));
Q_FDP4EP \o_label7_data0_REG[3] ( .CK(clk), .CE(n198), .R(n261), .D(n9), .Q(o_label7_data0[3]));
Q_FDP4EP \o_label7_data0_REG[4] ( .CK(clk), .CE(n198), .R(n261), .D(n10), .Q(o_label7_data0[4]));
Q_FDP4EP \o_label7_data0_REG[5] ( .CK(clk), .CE(n198), .R(n261), .D(n11), .Q(o_label7_data0[5]));
Q_FDP4EP \o_label7_data0_REG[6] ( .CK(clk), .CE(n198), .R(n261), .D(n12), .Q(o_label7_data0[6]));
Q_FDP4EP \o_label7_data0_REG[7] ( .CK(clk), .CE(n198), .R(n261), .D(n13), .Q(o_label7_data0[7]));
Q_FDP4EP \o_label7_data0_REG[8] ( .CK(clk), .CE(n198), .R(n261), .D(n14), .Q(o_label7_data0[8]));
Q_FDP4EP \o_label7_data0_REG[9] ( .CK(clk), .CE(n198), .R(n261), .D(n15), .Q(o_label7_data0[9]));
Q_FDP4EP \o_label7_data0_REG[10] ( .CK(clk), .CE(n198), .R(n261), .D(n16), .Q(o_label7_data0[10]));
Q_FDP4EP \o_label7_data0_REG[11] ( .CK(clk), .CE(n198), .R(n261), .D(n17), .Q(o_label7_data0[11]));
Q_FDP4EP \o_label7_data0_REG[12] ( .CK(clk), .CE(n198), .R(n261), .D(n18), .Q(o_label7_data0[12]));
Q_FDP4EP \o_label7_data0_REG[13] ( .CK(clk), .CE(n198), .R(n261), .D(n19), .Q(o_label7_data0[13]));
Q_FDP4EP \o_label7_data0_REG[14] ( .CK(clk), .CE(n198), .R(n261), .D(n20), .Q(o_label7_data0[14]));
Q_FDP4EP \o_label7_data0_REG[15] ( .CK(clk), .CE(n198), .R(n261), .D(n21), .Q(o_label7_data0[15]));
Q_FDP4EP \o_label7_data0_REG[16] ( .CK(clk), .CE(n198), .R(n261), .D(n22), .Q(o_label7_data0[16]));
Q_FDP4EP \o_label7_data0_REG[17] ( .CK(clk), .CE(n198), .R(n261), .D(n23), .Q(o_label7_data0[17]));
Q_FDP4EP \o_label7_data0_REG[18] ( .CK(clk), .CE(n198), .R(n261), .D(n24), .Q(o_label7_data0[18]));
Q_FDP4EP \o_label7_data0_REG[19] ( .CK(clk), .CE(n198), .R(n261), .D(n25), .Q(o_label7_data0[19]));
Q_FDP4EP \o_label7_data0_REG[20] ( .CK(clk), .CE(n198), .R(n261), .D(n26), .Q(o_label7_data0[20]));
Q_FDP4EP \o_label7_data0_REG[21] ( .CK(clk), .CE(n198), .R(n261), .D(n27), .Q(o_label7_data0[21]));
Q_FDP4EP \o_label7_data0_REG[22] ( .CK(clk), .CE(n198), .R(n261), .D(n28), .Q(o_label7_data0[22]));
Q_FDP4EP \o_label7_data0_REG[23] ( .CK(clk), .CE(n198), .R(n261), .D(n29), .Q(o_label7_data0[23]));
Q_FDP4EP \o_label7_data0_REG[24] ( .CK(clk), .CE(n198), .R(n261), .D(n30), .Q(o_label7_data0[24]));
Q_FDP4EP \o_label7_data0_REG[25] ( .CK(clk), .CE(n198), .R(n261), .D(n31), .Q(o_label7_data0[25]));
Q_FDP4EP \o_label7_data0_REG[26] ( .CK(clk), .CE(n198), .R(n261), .D(n32), .Q(o_label7_data0[26]));
Q_FDP4EP \o_label7_data0_REG[27] ( .CK(clk), .CE(n198), .R(n261), .D(n33), .Q(o_label7_data0[27]));
Q_FDP4EP \o_label7_data0_REG[28] ( .CK(clk), .CE(n198), .R(n261), .D(n34), .Q(o_label7_data0[28]));
Q_FDP4EP \o_label7_data0_REG[29] ( .CK(clk), .CE(n198), .R(n261), .D(n35), .Q(o_label7_data0[29]));
Q_FDP4EP \o_label7_data0_REG[30] ( .CK(clk), .CE(n198), .R(n261), .D(n36), .Q(o_label7_data0[30]));
Q_FDP4EP \o_label7_data0_REG[31] ( .CK(clk), .CE(n198), .R(n261), .D(n37), .Q(o_label7_data0[31]));
Q_FDP4EP \o_label7_data1_REG[0] ( .CK(clk), .CE(n197), .R(n261), .D(n6), .Q(o_label7_data1[0]));
Q_FDP4EP \o_label7_data1_REG[1] ( .CK(clk), .CE(n197), .R(n261), .D(n7), .Q(o_label7_data1[1]));
Q_FDP4EP \o_label7_data1_REG[2] ( .CK(clk), .CE(n197), .R(n261), .D(n8), .Q(o_label7_data1[2]));
Q_FDP4EP \o_label7_data1_REG[3] ( .CK(clk), .CE(n197), .R(n261), .D(n9), .Q(o_label7_data1[3]));
Q_FDP4EP \o_label7_data1_REG[4] ( .CK(clk), .CE(n197), .R(n261), .D(n10), .Q(o_label7_data1[4]));
Q_FDP4EP \o_label7_data1_REG[5] ( .CK(clk), .CE(n197), .R(n261), .D(n11), .Q(o_label7_data1[5]));
Q_FDP4EP \o_label7_data1_REG[6] ( .CK(clk), .CE(n197), .R(n261), .D(n12), .Q(o_label7_data1[6]));
Q_FDP4EP \o_label7_data1_REG[7] ( .CK(clk), .CE(n197), .R(n261), .D(n13), .Q(o_label7_data1[7]));
Q_FDP4EP \o_label7_data1_REG[8] ( .CK(clk), .CE(n197), .R(n261), .D(n14), .Q(o_label7_data1[8]));
Q_FDP4EP \o_label7_data1_REG[9] ( .CK(clk), .CE(n197), .R(n261), .D(n15), .Q(o_label7_data1[9]));
Q_FDP4EP \o_label7_data1_REG[10] ( .CK(clk), .CE(n197), .R(n261), .D(n16), .Q(o_label7_data1[10]));
Q_FDP4EP \o_label7_data1_REG[11] ( .CK(clk), .CE(n197), .R(n261), .D(n17), .Q(o_label7_data1[11]));
Q_FDP4EP \o_label7_data1_REG[12] ( .CK(clk), .CE(n197), .R(n261), .D(n18), .Q(o_label7_data1[12]));
Q_FDP4EP \o_label7_data1_REG[13] ( .CK(clk), .CE(n197), .R(n261), .D(n19), .Q(o_label7_data1[13]));
Q_FDP4EP \o_label7_data1_REG[14] ( .CK(clk), .CE(n197), .R(n261), .D(n20), .Q(o_label7_data1[14]));
Q_FDP4EP \o_label7_data1_REG[15] ( .CK(clk), .CE(n197), .R(n261), .D(n21), .Q(o_label7_data1[15]));
Q_FDP4EP \o_label7_data1_REG[16] ( .CK(clk), .CE(n197), .R(n261), .D(n22), .Q(o_label7_data1[16]));
Q_FDP4EP \o_label7_data1_REG[17] ( .CK(clk), .CE(n197), .R(n261), .D(n23), .Q(o_label7_data1[17]));
Q_FDP4EP \o_label7_data1_REG[18] ( .CK(clk), .CE(n197), .R(n261), .D(n24), .Q(o_label7_data1[18]));
Q_FDP4EP \o_label7_data1_REG[19] ( .CK(clk), .CE(n197), .R(n261), .D(n25), .Q(o_label7_data1[19]));
Q_FDP4EP \o_label7_data1_REG[20] ( .CK(clk), .CE(n197), .R(n261), .D(n26), .Q(o_label7_data1[20]));
Q_FDP4EP \o_label7_data1_REG[21] ( .CK(clk), .CE(n197), .R(n261), .D(n27), .Q(o_label7_data1[21]));
Q_FDP4EP \o_label7_data1_REG[22] ( .CK(clk), .CE(n197), .R(n261), .D(n28), .Q(o_label7_data1[22]));
Q_FDP4EP \o_label7_data1_REG[23] ( .CK(clk), .CE(n197), .R(n261), .D(n29), .Q(o_label7_data1[23]));
Q_FDP4EP \o_label7_data1_REG[24] ( .CK(clk), .CE(n197), .R(n261), .D(n30), .Q(o_label7_data1[24]));
Q_FDP4EP \o_label7_data1_REG[25] ( .CK(clk), .CE(n197), .R(n261), .D(n31), .Q(o_label7_data1[25]));
Q_FDP4EP \o_label7_data1_REG[26] ( .CK(clk), .CE(n197), .R(n261), .D(n32), .Q(o_label7_data1[26]));
Q_FDP4EP \o_label7_data1_REG[27] ( .CK(clk), .CE(n197), .R(n261), .D(n33), .Q(o_label7_data1[27]));
Q_FDP4EP \o_label7_data1_REG[28] ( .CK(clk), .CE(n197), .R(n261), .D(n34), .Q(o_label7_data1[28]));
Q_FDP4EP \o_label7_data1_REG[29] ( .CK(clk), .CE(n197), .R(n261), .D(n35), .Q(o_label7_data1[29]));
Q_FDP4EP \o_label7_data1_REG[30] ( .CK(clk), .CE(n197), .R(n261), .D(n36), .Q(o_label7_data1[30]));
Q_FDP4EP \o_label7_data1_REG[31] ( .CK(clk), .CE(n197), .R(n261), .D(n37), .Q(o_label7_data1[31]));
Q_FDP4EP \o_label7_data2_REG[0] ( .CK(clk), .CE(n196), .R(n261), .D(n6), .Q(o_label7_data2[0]));
Q_FDP4EP \o_label7_data2_REG[1] ( .CK(clk), .CE(n196), .R(n261), .D(n7), .Q(o_label7_data2[1]));
Q_FDP4EP \o_label7_data2_REG[2] ( .CK(clk), .CE(n196), .R(n261), .D(n8), .Q(o_label7_data2[2]));
Q_FDP4EP \o_label7_data2_REG[3] ( .CK(clk), .CE(n196), .R(n261), .D(n9), .Q(o_label7_data2[3]));
Q_FDP4EP \o_label7_data2_REG[4] ( .CK(clk), .CE(n196), .R(n261), .D(n10), .Q(o_label7_data2[4]));
Q_FDP4EP \o_label7_data2_REG[5] ( .CK(clk), .CE(n196), .R(n261), .D(n11), .Q(o_label7_data2[5]));
Q_FDP4EP \o_label7_data2_REG[6] ( .CK(clk), .CE(n196), .R(n261), .D(n12), .Q(o_label7_data2[6]));
Q_FDP4EP \o_label7_data2_REG[7] ( .CK(clk), .CE(n196), .R(n261), .D(n13), .Q(o_label7_data2[7]));
Q_FDP4EP \o_label7_data2_REG[8] ( .CK(clk), .CE(n196), .R(n261), .D(n14), .Q(o_label7_data2[8]));
Q_FDP4EP \o_label7_data2_REG[9] ( .CK(clk), .CE(n196), .R(n261), .D(n15), .Q(o_label7_data2[9]));
Q_FDP4EP \o_label7_data2_REG[10] ( .CK(clk), .CE(n196), .R(n261), .D(n16), .Q(o_label7_data2[10]));
Q_FDP4EP \o_label7_data2_REG[11] ( .CK(clk), .CE(n196), .R(n261), .D(n17), .Q(o_label7_data2[11]));
Q_FDP4EP \o_label7_data2_REG[12] ( .CK(clk), .CE(n196), .R(n261), .D(n18), .Q(o_label7_data2[12]));
Q_FDP4EP \o_label7_data2_REG[13] ( .CK(clk), .CE(n196), .R(n261), .D(n19), .Q(o_label7_data2[13]));
Q_FDP4EP \o_label7_data2_REG[14] ( .CK(clk), .CE(n196), .R(n261), .D(n20), .Q(o_label7_data2[14]));
Q_FDP4EP \o_label7_data2_REG[15] ( .CK(clk), .CE(n196), .R(n261), .D(n21), .Q(o_label7_data2[15]));
Q_FDP4EP \o_label7_data2_REG[16] ( .CK(clk), .CE(n196), .R(n261), .D(n22), .Q(o_label7_data2[16]));
Q_FDP4EP \o_label7_data2_REG[17] ( .CK(clk), .CE(n196), .R(n261), .D(n23), .Q(o_label7_data2[17]));
Q_FDP4EP \o_label7_data2_REG[18] ( .CK(clk), .CE(n196), .R(n261), .D(n24), .Q(o_label7_data2[18]));
Q_FDP4EP \o_label7_data2_REG[19] ( .CK(clk), .CE(n196), .R(n261), .D(n25), .Q(o_label7_data2[19]));
Q_FDP4EP \o_label7_data2_REG[20] ( .CK(clk), .CE(n196), .R(n261), .D(n26), .Q(o_label7_data2[20]));
Q_FDP4EP \o_label7_data2_REG[21] ( .CK(clk), .CE(n196), .R(n261), .D(n27), .Q(o_label7_data2[21]));
Q_FDP4EP \o_label7_data2_REG[22] ( .CK(clk), .CE(n196), .R(n261), .D(n28), .Q(o_label7_data2[22]));
Q_FDP4EP \o_label7_data2_REG[23] ( .CK(clk), .CE(n196), .R(n261), .D(n29), .Q(o_label7_data2[23]));
Q_FDP4EP \o_label7_data2_REG[24] ( .CK(clk), .CE(n196), .R(n261), .D(n30), .Q(o_label7_data2[24]));
Q_FDP4EP \o_label7_data2_REG[25] ( .CK(clk), .CE(n196), .R(n261), .D(n31), .Q(o_label7_data2[25]));
Q_FDP4EP \o_label7_data2_REG[26] ( .CK(clk), .CE(n196), .R(n261), .D(n32), .Q(o_label7_data2[26]));
Q_FDP4EP \o_label7_data2_REG[27] ( .CK(clk), .CE(n196), .R(n261), .D(n33), .Q(o_label7_data2[27]));
Q_FDP4EP \o_label7_data2_REG[28] ( .CK(clk), .CE(n196), .R(n261), .D(n34), .Q(o_label7_data2[28]));
Q_FDP4EP \o_label7_data2_REG[29] ( .CK(clk), .CE(n196), .R(n261), .D(n35), .Q(o_label7_data2[29]));
Q_FDP4EP \o_label7_data2_REG[30] ( .CK(clk), .CE(n196), .R(n261), .D(n36), .Q(o_label7_data2[30]));
Q_FDP4EP \o_label7_data2_REG[31] ( .CK(clk), .CE(n196), .R(n261), .D(n37), .Q(o_label7_data2[31]));
Q_FDP4EP \o_label7_data3_REG[0] ( .CK(clk), .CE(n195), .R(n261), .D(n6), .Q(o_label7_data3[0]));
Q_FDP4EP \o_label7_data3_REG[1] ( .CK(clk), .CE(n195), .R(n261), .D(n7), .Q(o_label7_data3[1]));
Q_FDP4EP \o_label7_data3_REG[2] ( .CK(clk), .CE(n195), .R(n261), .D(n8), .Q(o_label7_data3[2]));
Q_FDP4EP \o_label7_data3_REG[3] ( .CK(clk), .CE(n195), .R(n261), .D(n9), .Q(o_label7_data3[3]));
Q_FDP4EP \o_label7_data3_REG[4] ( .CK(clk), .CE(n195), .R(n261), .D(n10), .Q(o_label7_data3[4]));
Q_FDP4EP \o_label7_data3_REG[5] ( .CK(clk), .CE(n195), .R(n261), .D(n11), .Q(o_label7_data3[5]));
Q_FDP4EP \o_label7_data3_REG[6] ( .CK(clk), .CE(n195), .R(n261), .D(n12), .Q(o_label7_data3[6]));
Q_FDP4EP \o_label7_data3_REG[7] ( .CK(clk), .CE(n195), .R(n261), .D(n13), .Q(o_label7_data3[7]));
Q_FDP4EP \o_label7_data3_REG[8] ( .CK(clk), .CE(n195), .R(n261), .D(n14), .Q(o_label7_data3[8]));
Q_FDP4EP \o_label7_data3_REG[9] ( .CK(clk), .CE(n195), .R(n261), .D(n15), .Q(o_label7_data3[9]));
Q_FDP4EP \o_label7_data3_REG[10] ( .CK(clk), .CE(n195), .R(n261), .D(n16), .Q(o_label7_data3[10]));
Q_FDP4EP \o_label7_data3_REG[11] ( .CK(clk), .CE(n195), .R(n261), .D(n17), .Q(o_label7_data3[11]));
Q_FDP4EP \o_label7_data3_REG[12] ( .CK(clk), .CE(n195), .R(n261), .D(n18), .Q(o_label7_data3[12]));
Q_FDP4EP \o_label7_data3_REG[13] ( .CK(clk), .CE(n195), .R(n261), .D(n19), .Q(o_label7_data3[13]));
Q_FDP4EP \o_label7_data3_REG[14] ( .CK(clk), .CE(n195), .R(n261), .D(n20), .Q(o_label7_data3[14]));
Q_FDP4EP \o_label7_data3_REG[15] ( .CK(clk), .CE(n195), .R(n261), .D(n21), .Q(o_label7_data3[15]));
Q_FDP4EP \o_label7_data3_REG[16] ( .CK(clk), .CE(n195), .R(n261), .D(n22), .Q(o_label7_data3[16]));
Q_FDP4EP \o_label7_data3_REG[17] ( .CK(clk), .CE(n195), .R(n261), .D(n23), .Q(o_label7_data3[17]));
Q_FDP4EP \o_label7_data3_REG[18] ( .CK(clk), .CE(n195), .R(n261), .D(n24), .Q(o_label7_data3[18]));
Q_FDP4EP \o_label7_data3_REG[19] ( .CK(clk), .CE(n195), .R(n261), .D(n25), .Q(o_label7_data3[19]));
Q_FDP4EP \o_label7_data3_REG[20] ( .CK(clk), .CE(n195), .R(n261), .D(n26), .Q(o_label7_data3[20]));
Q_FDP4EP \o_label7_data3_REG[21] ( .CK(clk), .CE(n195), .R(n261), .D(n27), .Q(o_label7_data3[21]));
Q_FDP4EP \o_label7_data3_REG[22] ( .CK(clk), .CE(n195), .R(n261), .D(n28), .Q(o_label7_data3[22]));
Q_FDP4EP \o_label7_data3_REG[23] ( .CK(clk), .CE(n195), .R(n261), .D(n29), .Q(o_label7_data3[23]));
Q_FDP4EP \o_label7_data3_REG[24] ( .CK(clk), .CE(n195), .R(n261), .D(n30), .Q(o_label7_data3[24]));
Q_FDP4EP \o_label7_data3_REG[25] ( .CK(clk), .CE(n195), .R(n261), .D(n31), .Q(o_label7_data3[25]));
Q_FDP4EP \o_label7_data3_REG[26] ( .CK(clk), .CE(n195), .R(n261), .D(n32), .Q(o_label7_data3[26]));
Q_FDP4EP \o_label7_data3_REG[27] ( .CK(clk), .CE(n195), .R(n261), .D(n33), .Q(o_label7_data3[27]));
Q_FDP4EP \o_label7_data3_REG[28] ( .CK(clk), .CE(n195), .R(n261), .D(n34), .Q(o_label7_data3[28]));
Q_FDP4EP \o_label7_data3_REG[29] ( .CK(clk), .CE(n195), .R(n261), .D(n35), .Q(o_label7_data3[29]));
Q_FDP4EP \o_label7_data3_REG[30] ( .CK(clk), .CE(n195), .R(n261), .D(n36), .Q(o_label7_data3[30]));
Q_FDP4EP \o_label7_data3_REG[31] ( .CK(clk), .CE(n195), .R(n261), .D(n37), .Q(o_label7_data3[31]));
Q_FDP4EP \o_label7_data4_REG[0] ( .CK(clk), .CE(n194), .R(n261), .D(n6), .Q(o_label7_data4[0]));
Q_FDP4EP \o_label7_data4_REG[1] ( .CK(clk), .CE(n194), .R(n261), .D(n7), .Q(o_label7_data4[1]));
Q_FDP4EP \o_label7_data4_REG[2] ( .CK(clk), .CE(n194), .R(n261), .D(n8), .Q(o_label7_data4[2]));
Q_FDP4EP \o_label7_data4_REG[3] ( .CK(clk), .CE(n194), .R(n261), .D(n9), .Q(o_label7_data4[3]));
Q_FDP4EP \o_label7_data4_REG[4] ( .CK(clk), .CE(n194), .R(n261), .D(n10), .Q(o_label7_data4[4]));
Q_FDP4EP \o_label7_data4_REG[5] ( .CK(clk), .CE(n194), .R(n261), .D(n11), .Q(o_label7_data4[5]));
Q_FDP4EP \o_label7_data4_REG[6] ( .CK(clk), .CE(n194), .R(n261), .D(n12), .Q(o_label7_data4[6]));
Q_FDP4EP \o_label7_data4_REG[7] ( .CK(clk), .CE(n194), .R(n261), .D(n13), .Q(o_label7_data4[7]));
Q_FDP4EP \o_label7_data4_REG[8] ( .CK(clk), .CE(n194), .R(n261), .D(n14), .Q(o_label7_data4[8]));
Q_FDP4EP \o_label7_data4_REG[9] ( .CK(clk), .CE(n194), .R(n261), .D(n15), .Q(o_label7_data4[9]));
Q_FDP4EP \o_label7_data4_REG[10] ( .CK(clk), .CE(n194), .R(n261), .D(n16), .Q(o_label7_data4[10]));
Q_FDP4EP \o_label7_data4_REG[11] ( .CK(clk), .CE(n194), .R(n261), .D(n17), .Q(o_label7_data4[11]));
Q_FDP4EP \o_label7_data4_REG[12] ( .CK(clk), .CE(n194), .R(n261), .D(n18), .Q(o_label7_data4[12]));
Q_FDP4EP \o_label7_data4_REG[13] ( .CK(clk), .CE(n194), .R(n261), .D(n19), .Q(o_label7_data4[13]));
Q_FDP4EP \o_label7_data4_REG[14] ( .CK(clk), .CE(n194), .R(n261), .D(n20), .Q(o_label7_data4[14]));
Q_FDP4EP \o_label7_data4_REG[15] ( .CK(clk), .CE(n194), .R(n261), .D(n21), .Q(o_label7_data4[15]));
Q_FDP4EP \o_label7_data4_REG[16] ( .CK(clk), .CE(n194), .R(n261), .D(n22), .Q(o_label7_data4[16]));
Q_FDP4EP \o_label7_data4_REG[17] ( .CK(clk), .CE(n194), .R(n261), .D(n23), .Q(o_label7_data4[17]));
Q_FDP4EP \o_label7_data4_REG[18] ( .CK(clk), .CE(n194), .R(n261), .D(n24), .Q(o_label7_data4[18]));
Q_FDP4EP \o_label7_data4_REG[19] ( .CK(clk), .CE(n194), .R(n261), .D(n25), .Q(o_label7_data4[19]));
Q_FDP4EP \o_label7_data4_REG[20] ( .CK(clk), .CE(n194), .R(n261), .D(n26), .Q(o_label7_data4[20]));
Q_FDP4EP \o_label7_data4_REG[21] ( .CK(clk), .CE(n194), .R(n261), .D(n27), .Q(o_label7_data4[21]));
Q_FDP4EP \o_label7_data4_REG[22] ( .CK(clk), .CE(n194), .R(n261), .D(n28), .Q(o_label7_data4[22]));
Q_FDP4EP \o_label7_data4_REG[23] ( .CK(clk), .CE(n194), .R(n261), .D(n29), .Q(o_label7_data4[23]));
Q_FDP4EP \o_label7_data4_REG[24] ( .CK(clk), .CE(n194), .R(n261), .D(n30), .Q(o_label7_data4[24]));
Q_FDP4EP \o_label7_data4_REG[25] ( .CK(clk), .CE(n194), .R(n261), .D(n31), .Q(o_label7_data4[25]));
Q_FDP4EP \o_label7_data4_REG[26] ( .CK(clk), .CE(n194), .R(n261), .D(n32), .Q(o_label7_data4[26]));
Q_FDP4EP \o_label7_data4_REG[27] ( .CK(clk), .CE(n194), .R(n261), .D(n33), .Q(o_label7_data4[27]));
Q_FDP4EP \o_label7_data4_REG[28] ( .CK(clk), .CE(n194), .R(n261), .D(n34), .Q(o_label7_data4[28]));
Q_FDP4EP \o_label7_data4_REG[29] ( .CK(clk), .CE(n194), .R(n261), .D(n35), .Q(o_label7_data4[29]));
Q_FDP4EP \o_label7_data4_REG[30] ( .CK(clk), .CE(n194), .R(n261), .D(n36), .Q(o_label7_data4[30]));
Q_FDP4EP \o_label7_data4_REG[31] ( .CK(clk), .CE(n194), .R(n261), .D(n37), .Q(o_label7_data4[31]));
Q_FDP4EP \o_label7_data5_REG[0] ( .CK(clk), .CE(n193), .R(n261), .D(n6), .Q(o_label7_data5[0]));
Q_FDP4EP \o_label7_data5_REG[1] ( .CK(clk), .CE(n193), .R(n261), .D(n7), .Q(o_label7_data5[1]));
Q_FDP4EP \o_label7_data5_REG[2] ( .CK(clk), .CE(n193), .R(n261), .D(n8), .Q(o_label7_data5[2]));
Q_FDP4EP \o_label7_data5_REG[3] ( .CK(clk), .CE(n193), .R(n261), .D(n9), .Q(o_label7_data5[3]));
Q_FDP4EP \o_label7_data5_REG[4] ( .CK(clk), .CE(n193), .R(n261), .D(n10), .Q(o_label7_data5[4]));
Q_FDP4EP \o_label7_data5_REG[5] ( .CK(clk), .CE(n193), .R(n261), .D(n11), .Q(o_label7_data5[5]));
Q_FDP4EP \o_label7_data5_REG[6] ( .CK(clk), .CE(n193), .R(n261), .D(n12), .Q(o_label7_data5[6]));
Q_FDP4EP \o_label7_data5_REG[7] ( .CK(clk), .CE(n193), .R(n261), .D(n13), .Q(o_label7_data5[7]));
Q_FDP4EP \o_label7_data5_REG[8] ( .CK(clk), .CE(n193), .R(n261), .D(n14), .Q(o_label7_data5[8]));
Q_FDP4EP \o_label7_data5_REG[9] ( .CK(clk), .CE(n193), .R(n261), .D(n15), .Q(o_label7_data5[9]));
Q_FDP4EP \o_label7_data5_REG[10] ( .CK(clk), .CE(n193), .R(n261), .D(n16), .Q(o_label7_data5[10]));
Q_FDP4EP \o_label7_data5_REG[11] ( .CK(clk), .CE(n193), .R(n261), .D(n17), .Q(o_label7_data5[11]));
Q_FDP4EP \o_label7_data5_REG[12] ( .CK(clk), .CE(n193), .R(n261), .D(n18), .Q(o_label7_data5[12]));
Q_FDP4EP \o_label7_data5_REG[13] ( .CK(clk), .CE(n193), .R(n261), .D(n19), .Q(o_label7_data5[13]));
Q_FDP4EP \o_label7_data5_REG[14] ( .CK(clk), .CE(n193), .R(n261), .D(n20), .Q(o_label7_data5[14]));
Q_FDP4EP \o_label7_data5_REG[15] ( .CK(clk), .CE(n193), .R(n261), .D(n21), .Q(o_label7_data5[15]));
Q_FDP4EP \o_label7_data5_REG[16] ( .CK(clk), .CE(n193), .R(n261), .D(n22), .Q(o_label7_data5[16]));
Q_FDP4EP \o_label7_data5_REG[17] ( .CK(clk), .CE(n193), .R(n261), .D(n23), .Q(o_label7_data5[17]));
Q_FDP4EP \o_label7_data5_REG[18] ( .CK(clk), .CE(n193), .R(n261), .D(n24), .Q(o_label7_data5[18]));
Q_FDP4EP \o_label7_data5_REG[19] ( .CK(clk), .CE(n193), .R(n261), .D(n25), .Q(o_label7_data5[19]));
Q_FDP4EP \o_label7_data5_REG[20] ( .CK(clk), .CE(n193), .R(n261), .D(n26), .Q(o_label7_data5[20]));
Q_FDP4EP \o_label7_data5_REG[21] ( .CK(clk), .CE(n193), .R(n261), .D(n27), .Q(o_label7_data5[21]));
Q_FDP4EP \o_label7_data5_REG[22] ( .CK(clk), .CE(n193), .R(n261), .D(n28), .Q(o_label7_data5[22]));
Q_FDP4EP \o_label7_data5_REG[23] ( .CK(clk), .CE(n193), .R(n261), .D(n29), .Q(o_label7_data5[23]));
Q_FDP4EP \o_label7_data5_REG[24] ( .CK(clk), .CE(n193), .R(n261), .D(n30), .Q(o_label7_data5[24]));
Q_FDP4EP \o_label7_data5_REG[25] ( .CK(clk), .CE(n193), .R(n261), .D(n31), .Q(o_label7_data5[25]));
Q_FDP4EP \o_label7_data5_REG[26] ( .CK(clk), .CE(n193), .R(n261), .D(n32), .Q(o_label7_data5[26]));
Q_FDP4EP \o_label7_data5_REG[27] ( .CK(clk), .CE(n193), .R(n261), .D(n33), .Q(o_label7_data5[27]));
Q_FDP4EP \o_label7_data5_REG[28] ( .CK(clk), .CE(n193), .R(n261), .D(n34), .Q(o_label7_data5[28]));
Q_FDP4EP \o_label7_data5_REG[29] ( .CK(clk), .CE(n193), .R(n261), .D(n35), .Q(o_label7_data5[29]));
Q_FDP4EP \o_label7_data5_REG[30] ( .CK(clk), .CE(n193), .R(n261), .D(n36), .Q(o_label7_data5[30]));
Q_FDP4EP \o_label7_data5_REG[31] ( .CK(clk), .CE(n193), .R(n261), .D(n37), .Q(o_label7_data5[31]));
Q_FDP4EP \o_label7_data6_REG[0] ( .CK(clk), .CE(n192), .R(n261), .D(n6), .Q(o_label7_data6[0]));
Q_FDP4EP \o_label7_data6_REG[1] ( .CK(clk), .CE(n192), .R(n261), .D(n7), .Q(o_label7_data6[1]));
Q_FDP4EP \o_label7_data6_REG[2] ( .CK(clk), .CE(n192), .R(n261), .D(n8), .Q(o_label7_data6[2]));
Q_FDP4EP \o_label7_data6_REG[3] ( .CK(clk), .CE(n192), .R(n261), .D(n9), .Q(o_label7_data6[3]));
Q_FDP4EP \o_label7_data6_REG[4] ( .CK(clk), .CE(n192), .R(n261), .D(n10), .Q(o_label7_data6[4]));
Q_FDP4EP \o_label7_data6_REG[5] ( .CK(clk), .CE(n192), .R(n261), .D(n11), .Q(o_label7_data6[5]));
Q_FDP4EP \o_label7_data6_REG[6] ( .CK(clk), .CE(n192), .R(n261), .D(n12), .Q(o_label7_data6[6]));
Q_FDP4EP \o_label7_data6_REG[7] ( .CK(clk), .CE(n192), .R(n261), .D(n13), .Q(o_label7_data6[7]));
Q_FDP4EP \o_label7_data6_REG[8] ( .CK(clk), .CE(n192), .R(n261), .D(n14), .Q(o_label7_data6[8]));
Q_FDP4EP \o_label7_data6_REG[9] ( .CK(clk), .CE(n192), .R(n261), .D(n15), .Q(o_label7_data6[9]));
Q_FDP4EP \o_label7_data6_REG[10] ( .CK(clk), .CE(n192), .R(n261), .D(n16), .Q(o_label7_data6[10]));
Q_FDP4EP \o_label7_data6_REG[11] ( .CK(clk), .CE(n192), .R(n261), .D(n17), .Q(o_label7_data6[11]));
Q_FDP4EP \o_label7_data6_REG[12] ( .CK(clk), .CE(n192), .R(n261), .D(n18), .Q(o_label7_data6[12]));
Q_FDP4EP \o_label7_data6_REG[13] ( .CK(clk), .CE(n192), .R(n261), .D(n19), .Q(o_label7_data6[13]));
Q_FDP4EP \o_label7_data6_REG[14] ( .CK(clk), .CE(n192), .R(n261), .D(n20), .Q(o_label7_data6[14]));
Q_FDP4EP \o_label7_data6_REG[15] ( .CK(clk), .CE(n192), .R(n261), .D(n21), .Q(o_label7_data6[15]));
Q_FDP4EP \o_label7_data6_REG[16] ( .CK(clk), .CE(n192), .R(n261), .D(n22), .Q(o_label7_data6[16]));
Q_FDP4EP \o_label7_data6_REG[17] ( .CK(clk), .CE(n192), .R(n261), .D(n23), .Q(o_label7_data6[17]));
Q_FDP4EP \o_label7_data6_REG[18] ( .CK(clk), .CE(n192), .R(n261), .D(n24), .Q(o_label7_data6[18]));
Q_FDP4EP \o_label7_data6_REG[19] ( .CK(clk), .CE(n192), .R(n261), .D(n25), .Q(o_label7_data6[19]));
Q_FDP4EP \o_label7_data6_REG[20] ( .CK(clk), .CE(n192), .R(n261), .D(n26), .Q(o_label7_data6[20]));
Q_FDP4EP \o_label7_data6_REG[21] ( .CK(clk), .CE(n192), .R(n261), .D(n27), .Q(o_label7_data6[21]));
Q_FDP4EP \o_label7_data6_REG[22] ( .CK(clk), .CE(n192), .R(n261), .D(n28), .Q(o_label7_data6[22]));
Q_FDP4EP \o_label7_data6_REG[23] ( .CK(clk), .CE(n192), .R(n261), .D(n29), .Q(o_label7_data6[23]));
Q_FDP4EP \o_label7_data6_REG[24] ( .CK(clk), .CE(n192), .R(n261), .D(n30), .Q(o_label7_data6[24]));
Q_FDP4EP \o_label7_data6_REG[25] ( .CK(clk), .CE(n192), .R(n261), .D(n31), .Q(o_label7_data6[25]));
Q_FDP4EP \o_label7_data6_REG[26] ( .CK(clk), .CE(n192), .R(n261), .D(n32), .Q(o_label7_data6[26]));
Q_FDP4EP \o_label7_data6_REG[27] ( .CK(clk), .CE(n192), .R(n261), .D(n33), .Q(o_label7_data6[27]));
Q_FDP4EP \o_label7_data6_REG[28] ( .CK(clk), .CE(n192), .R(n261), .D(n34), .Q(o_label7_data6[28]));
Q_FDP4EP \o_label7_data6_REG[29] ( .CK(clk), .CE(n192), .R(n261), .D(n35), .Q(o_label7_data6[29]));
Q_FDP4EP \o_label7_data6_REG[30] ( .CK(clk), .CE(n192), .R(n261), .D(n36), .Q(o_label7_data6[30]));
Q_FDP4EP \o_label7_data6_REG[31] ( .CK(clk), .CE(n192), .R(n261), .D(n37), .Q(o_label7_data6[31]));
Q_FDP4EP \o_label7_data7_REG[0] ( .CK(clk), .CE(n191), .R(n261), .D(n6), .Q(o_label7_data7[0]));
Q_FDP4EP \o_label7_data7_REG[1] ( .CK(clk), .CE(n191), .R(n261), .D(n7), .Q(o_label7_data7[1]));
Q_FDP4EP \o_label7_data7_REG[2] ( .CK(clk), .CE(n191), .R(n261), .D(n8), .Q(o_label7_data7[2]));
Q_FDP4EP \o_label7_data7_REG[3] ( .CK(clk), .CE(n191), .R(n261), .D(n9), .Q(o_label7_data7[3]));
Q_FDP4EP \o_label7_data7_REG[4] ( .CK(clk), .CE(n191), .R(n261), .D(n10), .Q(o_label7_data7[4]));
Q_FDP4EP \o_label7_data7_REG[5] ( .CK(clk), .CE(n191), .R(n261), .D(n11), .Q(o_label7_data7[5]));
Q_FDP4EP \o_label7_data7_REG[6] ( .CK(clk), .CE(n191), .R(n261), .D(n12), .Q(o_label7_data7[6]));
Q_FDP4EP \o_label7_data7_REG[7] ( .CK(clk), .CE(n191), .R(n261), .D(n13), .Q(o_label7_data7[7]));
Q_FDP4EP \o_label7_data7_REG[8] ( .CK(clk), .CE(n191), .R(n261), .D(n14), .Q(o_label7_data7[8]));
Q_FDP4EP \o_label7_data7_REG[9] ( .CK(clk), .CE(n191), .R(n261), .D(n15), .Q(o_label7_data7[9]));
Q_FDP4EP \o_label7_data7_REG[10] ( .CK(clk), .CE(n191), .R(n261), .D(n16), .Q(o_label7_data7[10]));
Q_FDP4EP \o_label7_data7_REG[11] ( .CK(clk), .CE(n191), .R(n261), .D(n17), .Q(o_label7_data7[11]));
Q_FDP4EP \o_label7_data7_REG[12] ( .CK(clk), .CE(n191), .R(n261), .D(n18), .Q(o_label7_data7[12]));
Q_FDP4EP \o_label7_data7_REG[13] ( .CK(clk), .CE(n191), .R(n261), .D(n19), .Q(o_label7_data7[13]));
Q_FDP4EP \o_label7_data7_REG[14] ( .CK(clk), .CE(n191), .R(n261), .D(n20), .Q(o_label7_data7[14]));
Q_FDP4EP \o_label7_data7_REG[15] ( .CK(clk), .CE(n191), .R(n261), .D(n21), .Q(o_label7_data7[15]));
Q_FDP4EP \o_label7_data7_REG[16] ( .CK(clk), .CE(n191), .R(n261), .D(n22), .Q(o_label7_data7[16]));
Q_FDP4EP \o_label7_data7_REG[17] ( .CK(clk), .CE(n191), .R(n261), .D(n23), .Q(o_label7_data7[17]));
Q_FDP4EP \o_label7_data7_REG[18] ( .CK(clk), .CE(n191), .R(n261), .D(n24), .Q(o_label7_data7[18]));
Q_FDP4EP \o_label7_data7_REG[19] ( .CK(clk), .CE(n191), .R(n261), .D(n25), .Q(o_label7_data7[19]));
Q_FDP4EP \o_label7_data7_REG[20] ( .CK(clk), .CE(n191), .R(n261), .D(n26), .Q(o_label7_data7[20]));
Q_FDP4EP \o_label7_data7_REG[21] ( .CK(clk), .CE(n191), .R(n261), .D(n27), .Q(o_label7_data7[21]));
Q_FDP4EP \o_label7_data7_REG[22] ( .CK(clk), .CE(n191), .R(n261), .D(n28), .Q(o_label7_data7[22]));
Q_FDP4EP \o_label7_data7_REG[23] ( .CK(clk), .CE(n191), .R(n261), .D(n29), .Q(o_label7_data7[23]));
Q_FDP4EP \o_label7_data7_REG[24] ( .CK(clk), .CE(n191), .R(n261), .D(n30), .Q(o_label7_data7[24]));
Q_FDP4EP \o_label7_data7_REG[25] ( .CK(clk), .CE(n191), .R(n261), .D(n31), .Q(o_label7_data7[25]));
Q_FDP4EP \o_label7_data7_REG[26] ( .CK(clk), .CE(n191), .R(n261), .D(n32), .Q(o_label7_data7[26]));
Q_FDP4EP \o_label7_data7_REG[27] ( .CK(clk), .CE(n191), .R(n261), .D(n33), .Q(o_label7_data7[27]));
Q_FDP4EP \o_label7_data7_REG[28] ( .CK(clk), .CE(n191), .R(n261), .D(n34), .Q(o_label7_data7[28]));
Q_FDP4EP \o_label7_data7_REG[29] ( .CK(clk), .CE(n191), .R(n261), .D(n35), .Q(o_label7_data7[29]));
Q_FDP4EP \o_label7_data7_REG[30] ( .CK(clk), .CE(n191), .R(n261), .D(n36), .Q(o_label7_data7[30]));
Q_FDP4EP \o_label7_data7_REG[31] ( .CK(clk), .CE(n191), .R(n261), .D(n37), .Q(o_label7_data7[31]));
Q_FDP4EP \o_label7_config_REG[0] ( .CK(clk), .CE(n190), .R(n261), .D(n6), .Q(o_label7_config[0]));
Q_FDP4EP \o_label7_config_REG[1] ( .CK(clk), .CE(n190), .R(n261), .D(n7), .Q(o_label7_config[1]));
Q_FDP4EP \o_label7_config_REG[2] ( .CK(clk), .CE(n190), .R(n261), .D(n8), .Q(o_label7_config[2]));
Q_FDP4EP \o_label7_config_REG[3] ( .CK(clk), .CE(n190), .R(n261), .D(n9), .Q(o_label7_config[3]));
Q_FDP4EP \o_label7_config_REG[4] ( .CK(clk), .CE(n190), .R(n261), .D(n10), .Q(o_label7_config[4]));
Q_FDP4EP \o_label7_config_REG[5] ( .CK(clk), .CE(n190), .R(n261), .D(n11), .Q(o_label7_config[5]));
Q_FDP4EP \o_label7_config_REG[6] ( .CK(clk), .CE(n190), .R(n261), .D(n12), .Q(o_label7_config[6]));
Q_FDP4EP \o_label7_config_REG[7] ( .CK(clk), .CE(n190), .R(n261), .D(n13), .Q(o_label7_config[7]));
Q_FDP4EP \o_label7_config_REG[9] ( .CK(clk), .CE(n190), .R(n261), .D(n31), .Q(o_label7_config[9]));
Q_FDP4EP \o_label7_config_REG[10] ( .CK(clk), .CE(n190), .R(n261), .D(n32), .Q(o_label7_config[10]));
Q_FDP4EP \o_label7_config_REG[11] ( .CK(clk), .CE(n190), .R(n261), .D(n33), .Q(o_label7_config[11]));
Q_FDP4EP \o_label7_config_REG[12] ( .CK(clk), .CE(n190), .R(n261), .D(n34), .Q(o_label7_config[12]));
Q_FDP4EP \o_label7_config_REG[13] ( .CK(clk), .CE(n190), .R(n261), .D(n35), .Q(o_label7_config[13]));
Q_FDP4EP \o_label7_config_REG[14] ( .CK(clk), .CE(n190), .R(n261), .D(n36), .Q(o_label7_config[14]));
Q_FDP4EP \o_label7_config_REG[15] ( .CK(clk), .CE(n190), .R(n261), .D(n37), .Q(o_label7_config[15]));
Q_FDP4EP \o_label6_data0_REG[0] ( .CK(clk), .CE(n189), .R(n261), .D(n6), .Q(o_label6_data0[0]));
Q_FDP4EP \o_label6_data0_REG[1] ( .CK(clk), .CE(n189), .R(n261), .D(n7), .Q(o_label6_data0[1]));
Q_FDP4EP \o_label6_data0_REG[2] ( .CK(clk), .CE(n189), .R(n261), .D(n8), .Q(o_label6_data0[2]));
Q_FDP4EP \o_label6_data0_REG[3] ( .CK(clk), .CE(n189), .R(n261), .D(n9), .Q(o_label6_data0[3]));
Q_FDP4EP \o_label6_data0_REG[4] ( .CK(clk), .CE(n189), .R(n261), .D(n10), .Q(o_label6_data0[4]));
Q_FDP4EP \o_label6_data0_REG[5] ( .CK(clk), .CE(n189), .R(n261), .D(n11), .Q(o_label6_data0[5]));
Q_FDP4EP \o_label6_data0_REG[6] ( .CK(clk), .CE(n189), .R(n261), .D(n12), .Q(o_label6_data0[6]));
Q_FDP4EP \o_label6_data0_REG[7] ( .CK(clk), .CE(n189), .R(n261), .D(n13), .Q(o_label6_data0[7]));
Q_FDP4EP \o_label6_data0_REG[8] ( .CK(clk), .CE(n189), .R(n261), .D(n14), .Q(o_label6_data0[8]));
Q_FDP4EP \o_label6_data0_REG[9] ( .CK(clk), .CE(n189), .R(n261), .D(n15), .Q(o_label6_data0[9]));
Q_FDP4EP \o_label6_data0_REG[10] ( .CK(clk), .CE(n189), .R(n261), .D(n16), .Q(o_label6_data0[10]));
Q_FDP4EP \o_label6_data0_REG[11] ( .CK(clk), .CE(n189), .R(n261), .D(n17), .Q(o_label6_data0[11]));
Q_FDP4EP \o_label6_data0_REG[12] ( .CK(clk), .CE(n189), .R(n261), .D(n18), .Q(o_label6_data0[12]));
Q_FDP4EP \o_label6_data0_REG[13] ( .CK(clk), .CE(n189), .R(n261), .D(n19), .Q(o_label6_data0[13]));
Q_FDP4EP \o_label6_data0_REG[14] ( .CK(clk), .CE(n189), .R(n261), .D(n20), .Q(o_label6_data0[14]));
Q_FDP4EP \o_label6_data0_REG[15] ( .CK(clk), .CE(n189), .R(n261), .D(n21), .Q(o_label6_data0[15]));
Q_FDP4EP \o_label6_data0_REG[16] ( .CK(clk), .CE(n189), .R(n261), .D(n22), .Q(o_label6_data0[16]));
Q_FDP4EP \o_label6_data0_REG[17] ( .CK(clk), .CE(n189), .R(n261), .D(n23), .Q(o_label6_data0[17]));
Q_FDP4EP \o_label6_data0_REG[18] ( .CK(clk), .CE(n189), .R(n261), .D(n24), .Q(o_label6_data0[18]));
Q_FDP4EP \o_label6_data0_REG[19] ( .CK(clk), .CE(n189), .R(n261), .D(n25), .Q(o_label6_data0[19]));
Q_FDP4EP \o_label6_data0_REG[20] ( .CK(clk), .CE(n189), .R(n261), .D(n26), .Q(o_label6_data0[20]));
Q_FDP4EP \o_label6_data0_REG[21] ( .CK(clk), .CE(n189), .R(n261), .D(n27), .Q(o_label6_data0[21]));
Q_FDP4EP \o_label6_data0_REG[22] ( .CK(clk), .CE(n189), .R(n261), .D(n28), .Q(o_label6_data0[22]));
Q_FDP4EP \o_label6_data0_REG[23] ( .CK(clk), .CE(n189), .R(n261), .D(n29), .Q(o_label6_data0[23]));
Q_FDP4EP \o_label6_data0_REG[24] ( .CK(clk), .CE(n189), .R(n261), .D(n30), .Q(o_label6_data0[24]));
Q_FDP4EP \o_label6_data0_REG[25] ( .CK(clk), .CE(n189), .R(n261), .D(n31), .Q(o_label6_data0[25]));
Q_FDP4EP \o_label6_data0_REG[26] ( .CK(clk), .CE(n189), .R(n261), .D(n32), .Q(o_label6_data0[26]));
Q_FDP4EP \o_label6_data0_REG[27] ( .CK(clk), .CE(n189), .R(n261), .D(n33), .Q(o_label6_data0[27]));
Q_FDP4EP \o_label6_data0_REG[28] ( .CK(clk), .CE(n189), .R(n261), .D(n34), .Q(o_label6_data0[28]));
Q_FDP4EP \o_label6_data0_REG[29] ( .CK(clk), .CE(n189), .R(n261), .D(n35), .Q(o_label6_data0[29]));
Q_FDP4EP \o_label6_data0_REG[30] ( .CK(clk), .CE(n189), .R(n261), .D(n36), .Q(o_label6_data0[30]));
Q_FDP4EP \o_label6_data0_REG[31] ( .CK(clk), .CE(n189), .R(n261), .D(n37), .Q(o_label6_data0[31]));
Q_FDP4EP \o_label6_data1_REG[0] ( .CK(clk), .CE(n188), .R(n261), .D(n6), .Q(o_label6_data1[0]));
Q_FDP4EP \o_label6_data1_REG[1] ( .CK(clk), .CE(n188), .R(n261), .D(n7), .Q(o_label6_data1[1]));
Q_FDP4EP \o_label6_data1_REG[2] ( .CK(clk), .CE(n188), .R(n261), .D(n8), .Q(o_label6_data1[2]));
Q_FDP4EP \o_label6_data1_REG[3] ( .CK(clk), .CE(n188), .R(n261), .D(n9), .Q(o_label6_data1[3]));
Q_FDP4EP \o_label6_data1_REG[4] ( .CK(clk), .CE(n188), .R(n261), .D(n10), .Q(o_label6_data1[4]));
Q_FDP4EP \o_label6_data1_REG[5] ( .CK(clk), .CE(n188), .R(n261), .D(n11), .Q(o_label6_data1[5]));
Q_FDP4EP \o_label6_data1_REG[6] ( .CK(clk), .CE(n188), .R(n261), .D(n12), .Q(o_label6_data1[6]));
Q_FDP4EP \o_label6_data1_REG[7] ( .CK(clk), .CE(n188), .R(n261), .D(n13), .Q(o_label6_data1[7]));
Q_FDP4EP \o_label6_data1_REG[8] ( .CK(clk), .CE(n188), .R(n261), .D(n14), .Q(o_label6_data1[8]));
Q_FDP4EP \o_label6_data1_REG[9] ( .CK(clk), .CE(n188), .R(n261), .D(n15), .Q(o_label6_data1[9]));
Q_FDP4EP \o_label6_data1_REG[10] ( .CK(clk), .CE(n188), .R(n261), .D(n16), .Q(o_label6_data1[10]));
Q_FDP4EP \o_label6_data1_REG[11] ( .CK(clk), .CE(n188), .R(n261), .D(n17), .Q(o_label6_data1[11]));
Q_FDP4EP \o_label6_data1_REG[12] ( .CK(clk), .CE(n188), .R(n261), .D(n18), .Q(o_label6_data1[12]));
Q_FDP4EP \o_label6_data1_REG[13] ( .CK(clk), .CE(n188), .R(n261), .D(n19), .Q(o_label6_data1[13]));
Q_FDP4EP \o_label6_data1_REG[14] ( .CK(clk), .CE(n188), .R(n261), .D(n20), .Q(o_label6_data1[14]));
Q_FDP4EP \o_label6_data1_REG[15] ( .CK(clk), .CE(n188), .R(n261), .D(n21), .Q(o_label6_data1[15]));
Q_FDP4EP \o_label6_data1_REG[16] ( .CK(clk), .CE(n188), .R(n261), .D(n22), .Q(o_label6_data1[16]));
Q_FDP4EP \o_label6_data1_REG[17] ( .CK(clk), .CE(n188), .R(n261), .D(n23), .Q(o_label6_data1[17]));
Q_FDP4EP \o_label6_data1_REG[18] ( .CK(clk), .CE(n188), .R(n261), .D(n24), .Q(o_label6_data1[18]));
Q_FDP4EP \o_label6_data1_REG[19] ( .CK(clk), .CE(n188), .R(n261), .D(n25), .Q(o_label6_data1[19]));
Q_FDP4EP \o_label6_data1_REG[20] ( .CK(clk), .CE(n188), .R(n261), .D(n26), .Q(o_label6_data1[20]));
Q_FDP4EP \o_label6_data1_REG[21] ( .CK(clk), .CE(n188), .R(n261), .D(n27), .Q(o_label6_data1[21]));
Q_FDP4EP \o_label6_data1_REG[22] ( .CK(clk), .CE(n188), .R(n261), .D(n28), .Q(o_label6_data1[22]));
Q_FDP4EP \o_label6_data1_REG[23] ( .CK(clk), .CE(n188), .R(n261), .D(n29), .Q(o_label6_data1[23]));
Q_FDP4EP \o_label6_data1_REG[24] ( .CK(clk), .CE(n188), .R(n261), .D(n30), .Q(o_label6_data1[24]));
Q_FDP4EP \o_label6_data1_REG[25] ( .CK(clk), .CE(n188), .R(n261), .D(n31), .Q(o_label6_data1[25]));
Q_FDP4EP \o_label6_data1_REG[26] ( .CK(clk), .CE(n188), .R(n261), .D(n32), .Q(o_label6_data1[26]));
Q_FDP4EP \o_label6_data1_REG[27] ( .CK(clk), .CE(n188), .R(n261), .D(n33), .Q(o_label6_data1[27]));
Q_FDP4EP \o_label6_data1_REG[28] ( .CK(clk), .CE(n188), .R(n261), .D(n34), .Q(o_label6_data1[28]));
Q_FDP4EP \o_label6_data1_REG[29] ( .CK(clk), .CE(n188), .R(n261), .D(n35), .Q(o_label6_data1[29]));
Q_FDP4EP \o_label6_data1_REG[30] ( .CK(clk), .CE(n188), .R(n261), .D(n36), .Q(o_label6_data1[30]));
Q_FDP4EP \o_label6_data1_REG[31] ( .CK(clk), .CE(n188), .R(n261), .D(n37), .Q(o_label6_data1[31]));
Q_FDP4EP \o_label6_data2_REG[0] ( .CK(clk), .CE(n187), .R(n261), .D(n6), .Q(o_label6_data2[0]));
Q_FDP4EP \o_label6_data2_REG[1] ( .CK(clk), .CE(n187), .R(n261), .D(n7), .Q(o_label6_data2[1]));
Q_FDP4EP \o_label6_data2_REG[2] ( .CK(clk), .CE(n187), .R(n261), .D(n8), .Q(o_label6_data2[2]));
Q_FDP4EP \o_label6_data2_REG[3] ( .CK(clk), .CE(n187), .R(n261), .D(n9), .Q(o_label6_data2[3]));
Q_FDP4EP \o_label6_data2_REG[4] ( .CK(clk), .CE(n187), .R(n261), .D(n10), .Q(o_label6_data2[4]));
Q_FDP4EP \o_label6_data2_REG[5] ( .CK(clk), .CE(n187), .R(n261), .D(n11), .Q(o_label6_data2[5]));
Q_FDP4EP \o_label6_data2_REG[6] ( .CK(clk), .CE(n187), .R(n261), .D(n12), .Q(o_label6_data2[6]));
Q_FDP4EP \o_label6_data2_REG[7] ( .CK(clk), .CE(n187), .R(n261), .D(n13), .Q(o_label6_data2[7]));
Q_FDP4EP \o_label6_data2_REG[8] ( .CK(clk), .CE(n187), .R(n261), .D(n14), .Q(o_label6_data2[8]));
Q_FDP4EP \o_label6_data2_REG[9] ( .CK(clk), .CE(n187), .R(n261), .D(n15), .Q(o_label6_data2[9]));
Q_FDP4EP \o_label6_data2_REG[10] ( .CK(clk), .CE(n187), .R(n261), .D(n16), .Q(o_label6_data2[10]));
Q_FDP4EP \o_label6_data2_REG[11] ( .CK(clk), .CE(n187), .R(n261), .D(n17), .Q(o_label6_data2[11]));
Q_FDP4EP \o_label6_data2_REG[12] ( .CK(clk), .CE(n187), .R(n261), .D(n18), .Q(o_label6_data2[12]));
Q_FDP4EP \o_label6_data2_REG[13] ( .CK(clk), .CE(n187), .R(n261), .D(n19), .Q(o_label6_data2[13]));
Q_FDP4EP \o_label6_data2_REG[14] ( .CK(clk), .CE(n187), .R(n261), .D(n20), .Q(o_label6_data2[14]));
Q_FDP4EP \o_label6_data2_REG[15] ( .CK(clk), .CE(n187), .R(n261), .D(n21), .Q(o_label6_data2[15]));
Q_FDP4EP \o_label6_data2_REG[16] ( .CK(clk), .CE(n187), .R(n261), .D(n22), .Q(o_label6_data2[16]));
Q_FDP4EP \o_label6_data2_REG[17] ( .CK(clk), .CE(n187), .R(n261), .D(n23), .Q(o_label6_data2[17]));
Q_FDP4EP \o_label6_data2_REG[18] ( .CK(clk), .CE(n187), .R(n261), .D(n24), .Q(o_label6_data2[18]));
Q_FDP4EP \o_label6_data2_REG[19] ( .CK(clk), .CE(n187), .R(n261), .D(n25), .Q(o_label6_data2[19]));
Q_FDP4EP \o_label6_data2_REG[20] ( .CK(clk), .CE(n187), .R(n261), .D(n26), .Q(o_label6_data2[20]));
Q_FDP4EP \o_label6_data2_REG[21] ( .CK(clk), .CE(n187), .R(n261), .D(n27), .Q(o_label6_data2[21]));
Q_FDP4EP \o_label6_data2_REG[22] ( .CK(clk), .CE(n187), .R(n261), .D(n28), .Q(o_label6_data2[22]));
Q_FDP4EP \o_label6_data2_REG[23] ( .CK(clk), .CE(n187), .R(n261), .D(n29), .Q(o_label6_data2[23]));
Q_FDP4EP \o_label6_data2_REG[24] ( .CK(clk), .CE(n187), .R(n261), .D(n30), .Q(o_label6_data2[24]));
Q_FDP4EP \o_label6_data2_REG[25] ( .CK(clk), .CE(n187), .R(n261), .D(n31), .Q(o_label6_data2[25]));
Q_FDP4EP \o_label6_data2_REG[26] ( .CK(clk), .CE(n187), .R(n261), .D(n32), .Q(o_label6_data2[26]));
Q_FDP4EP \o_label6_data2_REG[27] ( .CK(clk), .CE(n187), .R(n261), .D(n33), .Q(o_label6_data2[27]));
Q_FDP4EP \o_label6_data2_REG[28] ( .CK(clk), .CE(n187), .R(n261), .D(n34), .Q(o_label6_data2[28]));
Q_FDP4EP \o_label6_data2_REG[29] ( .CK(clk), .CE(n187), .R(n261), .D(n35), .Q(o_label6_data2[29]));
Q_FDP4EP \o_label6_data2_REG[30] ( .CK(clk), .CE(n187), .R(n261), .D(n36), .Q(o_label6_data2[30]));
Q_FDP4EP \o_label6_data2_REG[31] ( .CK(clk), .CE(n187), .R(n261), .D(n37), .Q(o_label6_data2[31]));
Q_FDP4EP \o_label6_data3_REG[0] ( .CK(clk), .CE(n186), .R(n261), .D(n6), .Q(o_label6_data3[0]));
Q_FDP4EP \o_label6_data3_REG[1] ( .CK(clk), .CE(n186), .R(n261), .D(n7), .Q(o_label6_data3[1]));
Q_FDP4EP \o_label6_data3_REG[2] ( .CK(clk), .CE(n186), .R(n261), .D(n8), .Q(o_label6_data3[2]));
Q_FDP4EP \o_label6_data3_REG[3] ( .CK(clk), .CE(n186), .R(n261), .D(n9), .Q(o_label6_data3[3]));
Q_FDP4EP \o_label6_data3_REG[4] ( .CK(clk), .CE(n186), .R(n261), .D(n10), .Q(o_label6_data3[4]));
Q_FDP4EP \o_label6_data3_REG[5] ( .CK(clk), .CE(n186), .R(n261), .D(n11), .Q(o_label6_data3[5]));
Q_FDP4EP \o_label6_data3_REG[6] ( .CK(clk), .CE(n186), .R(n261), .D(n12), .Q(o_label6_data3[6]));
Q_FDP4EP \o_label6_data3_REG[7] ( .CK(clk), .CE(n186), .R(n261), .D(n13), .Q(o_label6_data3[7]));
Q_FDP4EP \o_label6_data3_REG[8] ( .CK(clk), .CE(n186), .R(n261), .D(n14), .Q(o_label6_data3[8]));
Q_FDP4EP \o_label6_data3_REG[9] ( .CK(clk), .CE(n186), .R(n261), .D(n15), .Q(o_label6_data3[9]));
Q_FDP4EP \o_label6_data3_REG[10] ( .CK(clk), .CE(n186), .R(n261), .D(n16), .Q(o_label6_data3[10]));
Q_FDP4EP \o_label6_data3_REG[11] ( .CK(clk), .CE(n186), .R(n261), .D(n17), .Q(o_label6_data3[11]));
Q_FDP4EP \o_label6_data3_REG[12] ( .CK(clk), .CE(n186), .R(n261), .D(n18), .Q(o_label6_data3[12]));
Q_FDP4EP \o_label6_data3_REG[13] ( .CK(clk), .CE(n186), .R(n261), .D(n19), .Q(o_label6_data3[13]));
Q_FDP4EP \o_label6_data3_REG[14] ( .CK(clk), .CE(n186), .R(n261), .D(n20), .Q(o_label6_data3[14]));
Q_FDP4EP \o_label6_data3_REG[15] ( .CK(clk), .CE(n186), .R(n261), .D(n21), .Q(o_label6_data3[15]));
Q_FDP4EP \o_label6_data3_REG[16] ( .CK(clk), .CE(n186), .R(n261), .D(n22), .Q(o_label6_data3[16]));
Q_FDP4EP \o_label6_data3_REG[17] ( .CK(clk), .CE(n186), .R(n261), .D(n23), .Q(o_label6_data3[17]));
Q_FDP4EP \o_label6_data3_REG[18] ( .CK(clk), .CE(n186), .R(n261), .D(n24), .Q(o_label6_data3[18]));
Q_FDP4EP \o_label6_data3_REG[19] ( .CK(clk), .CE(n186), .R(n261), .D(n25), .Q(o_label6_data3[19]));
Q_FDP4EP \o_label6_data3_REG[20] ( .CK(clk), .CE(n186), .R(n261), .D(n26), .Q(o_label6_data3[20]));
Q_FDP4EP \o_label6_data3_REG[21] ( .CK(clk), .CE(n186), .R(n261), .D(n27), .Q(o_label6_data3[21]));
Q_FDP4EP \o_label6_data3_REG[22] ( .CK(clk), .CE(n186), .R(n261), .D(n28), .Q(o_label6_data3[22]));
Q_FDP4EP \o_label6_data3_REG[23] ( .CK(clk), .CE(n186), .R(n261), .D(n29), .Q(o_label6_data3[23]));
Q_FDP4EP \o_label6_data3_REG[24] ( .CK(clk), .CE(n186), .R(n261), .D(n30), .Q(o_label6_data3[24]));
Q_FDP4EP \o_label6_data3_REG[25] ( .CK(clk), .CE(n186), .R(n261), .D(n31), .Q(o_label6_data3[25]));
Q_FDP4EP \o_label6_data3_REG[26] ( .CK(clk), .CE(n186), .R(n261), .D(n32), .Q(o_label6_data3[26]));
Q_FDP4EP \o_label6_data3_REG[27] ( .CK(clk), .CE(n186), .R(n261), .D(n33), .Q(o_label6_data3[27]));
Q_FDP4EP \o_label6_data3_REG[28] ( .CK(clk), .CE(n186), .R(n261), .D(n34), .Q(o_label6_data3[28]));
Q_FDP4EP \o_label6_data3_REG[29] ( .CK(clk), .CE(n186), .R(n261), .D(n35), .Q(o_label6_data3[29]));
Q_FDP4EP \o_label6_data3_REG[30] ( .CK(clk), .CE(n186), .R(n261), .D(n36), .Q(o_label6_data3[30]));
Q_FDP4EP \o_label6_data3_REG[31] ( .CK(clk), .CE(n186), .R(n261), .D(n37), .Q(o_label6_data3[31]));
Q_FDP4EP \o_label6_data4_REG[0] ( .CK(clk), .CE(n185), .R(n261), .D(n6), .Q(o_label6_data4[0]));
Q_FDP4EP \o_label6_data4_REG[1] ( .CK(clk), .CE(n185), .R(n261), .D(n7), .Q(o_label6_data4[1]));
Q_FDP4EP \o_label6_data4_REG[2] ( .CK(clk), .CE(n185), .R(n261), .D(n8), .Q(o_label6_data4[2]));
Q_FDP4EP \o_label6_data4_REG[3] ( .CK(clk), .CE(n185), .R(n261), .D(n9), .Q(o_label6_data4[3]));
Q_FDP4EP \o_label6_data4_REG[4] ( .CK(clk), .CE(n185), .R(n261), .D(n10), .Q(o_label6_data4[4]));
Q_FDP4EP \o_label6_data4_REG[5] ( .CK(clk), .CE(n185), .R(n261), .D(n11), .Q(o_label6_data4[5]));
Q_FDP4EP \o_label6_data4_REG[6] ( .CK(clk), .CE(n185), .R(n261), .D(n12), .Q(o_label6_data4[6]));
Q_FDP4EP \o_label6_data4_REG[7] ( .CK(clk), .CE(n185), .R(n261), .D(n13), .Q(o_label6_data4[7]));
Q_FDP4EP \o_label6_data4_REG[8] ( .CK(clk), .CE(n185), .R(n261), .D(n14), .Q(o_label6_data4[8]));
Q_FDP4EP \o_label6_data4_REG[9] ( .CK(clk), .CE(n185), .R(n261), .D(n15), .Q(o_label6_data4[9]));
Q_FDP4EP \o_label6_data4_REG[10] ( .CK(clk), .CE(n185), .R(n261), .D(n16), .Q(o_label6_data4[10]));
Q_FDP4EP \o_label6_data4_REG[11] ( .CK(clk), .CE(n185), .R(n261), .D(n17), .Q(o_label6_data4[11]));
Q_FDP4EP \o_label6_data4_REG[12] ( .CK(clk), .CE(n185), .R(n261), .D(n18), .Q(o_label6_data4[12]));
Q_FDP4EP \o_label6_data4_REG[13] ( .CK(clk), .CE(n185), .R(n261), .D(n19), .Q(o_label6_data4[13]));
Q_FDP4EP \o_label6_data4_REG[14] ( .CK(clk), .CE(n185), .R(n261), .D(n20), .Q(o_label6_data4[14]));
Q_FDP4EP \o_label6_data4_REG[15] ( .CK(clk), .CE(n185), .R(n261), .D(n21), .Q(o_label6_data4[15]));
Q_FDP4EP \o_label6_data4_REG[16] ( .CK(clk), .CE(n185), .R(n261), .D(n22), .Q(o_label6_data4[16]));
Q_FDP4EP \o_label6_data4_REG[17] ( .CK(clk), .CE(n185), .R(n261), .D(n23), .Q(o_label6_data4[17]));
Q_FDP4EP \o_label6_data4_REG[18] ( .CK(clk), .CE(n185), .R(n261), .D(n24), .Q(o_label6_data4[18]));
Q_FDP4EP \o_label6_data4_REG[19] ( .CK(clk), .CE(n185), .R(n261), .D(n25), .Q(o_label6_data4[19]));
Q_FDP4EP \o_label6_data4_REG[20] ( .CK(clk), .CE(n185), .R(n261), .D(n26), .Q(o_label6_data4[20]));
Q_FDP4EP \o_label6_data4_REG[21] ( .CK(clk), .CE(n185), .R(n261), .D(n27), .Q(o_label6_data4[21]));
Q_FDP4EP \o_label6_data4_REG[22] ( .CK(clk), .CE(n185), .R(n261), .D(n28), .Q(o_label6_data4[22]));
Q_FDP4EP \o_label6_data4_REG[23] ( .CK(clk), .CE(n185), .R(n261), .D(n29), .Q(o_label6_data4[23]));
Q_FDP4EP \o_label6_data4_REG[24] ( .CK(clk), .CE(n185), .R(n261), .D(n30), .Q(o_label6_data4[24]));
Q_FDP4EP \o_label6_data4_REG[25] ( .CK(clk), .CE(n185), .R(n261), .D(n31), .Q(o_label6_data4[25]));
Q_FDP4EP \o_label6_data4_REG[26] ( .CK(clk), .CE(n185), .R(n261), .D(n32), .Q(o_label6_data4[26]));
Q_FDP4EP \o_label6_data4_REG[27] ( .CK(clk), .CE(n185), .R(n261), .D(n33), .Q(o_label6_data4[27]));
Q_FDP4EP \o_label6_data4_REG[28] ( .CK(clk), .CE(n185), .R(n261), .D(n34), .Q(o_label6_data4[28]));
Q_FDP4EP \o_label6_data4_REG[29] ( .CK(clk), .CE(n185), .R(n261), .D(n35), .Q(o_label6_data4[29]));
Q_FDP4EP \o_label6_data4_REG[30] ( .CK(clk), .CE(n185), .R(n261), .D(n36), .Q(o_label6_data4[30]));
Q_FDP4EP \o_label6_data4_REG[31] ( .CK(clk), .CE(n185), .R(n261), .D(n37), .Q(o_label6_data4[31]));
Q_FDP4EP \o_label6_data5_REG[0] ( .CK(clk), .CE(n184), .R(n261), .D(n6), .Q(o_label6_data5[0]));
Q_FDP4EP \o_label6_data5_REG[1] ( .CK(clk), .CE(n184), .R(n261), .D(n7), .Q(o_label6_data5[1]));
Q_FDP4EP \o_label6_data5_REG[2] ( .CK(clk), .CE(n184), .R(n261), .D(n8), .Q(o_label6_data5[2]));
Q_FDP4EP \o_label6_data5_REG[3] ( .CK(clk), .CE(n184), .R(n261), .D(n9), .Q(o_label6_data5[3]));
Q_FDP4EP \o_label6_data5_REG[4] ( .CK(clk), .CE(n184), .R(n261), .D(n10), .Q(o_label6_data5[4]));
Q_FDP4EP \o_label6_data5_REG[5] ( .CK(clk), .CE(n184), .R(n261), .D(n11), .Q(o_label6_data5[5]));
Q_FDP4EP \o_label6_data5_REG[6] ( .CK(clk), .CE(n184), .R(n261), .D(n12), .Q(o_label6_data5[6]));
Q_FDP4EP \o_label6_data5_REG[7] ( .CK(clk), .CE(n184), .R(n261), .D(n13), .Q(o_label6_data5[7]));
Q_FDP4EP \o_label6_data5_REG[8] ( .CK(clk), .CE(n184), .R(n261), .D(n14), .Q(o_label6_data5[8]));
Q_FDP4EP \o_label6_data5_REG[9] ( .CK(clk), .CE(n184), .R(n261), .D(n15), .Q(o_label6_data5[9]));
Q_FDP4EP \o_label6_data5_REG[10] ( .CK(clk), .CE(n184), .R(n261), .D(n16), .Q(o_label6_data5[10]));
Q_FDP4EP \o_label6_data5_REG[11] ( .CK(clk), .CE(n184), .R(n261), .D(n17), .Q(o_label6_data5[11]));
Q_FDP4EP \o_label6_data5_REG[12] ( .CK(clk), .CE(n184), .R(n261), .D(n18), .Q(o_label6_data5[12]));
Q_FDP4EP \o_label6_data5_REG[13] ( .CK(clk), .CE(n184), .R(n261), .D(n19), .Q(o_label6_data5[13]));
Q_FDP4EP \o_label6_data5_REG[14] ( .CK(clk), .CE(n184), .R(n261), .D(n20), .Q(o_label6_data5[14]));
Q_FDP4EP \o_label6_data5_REG[15] ( .CK(clk), .CE(n184), .R(n261), .D(n21), .Q(o_label6_data5[15]));
Q_FDP4EP \o_label6_data5_REG[16] ( .CK(clk), .CE(n184), .R(n261), .D(n22), .Q(o_label6_data5[16]));
Q_FDP4EP \o_label6_data5_REG[17] ( .CK(clk), .CE(n184), .R(n261), .D(n23), .Q(o_label6_data5[17]));
Q_FDP4EP \o_label6_data5_REG[18] ( .CK(clk), .CE(n184), .R(n261), .D(n24), .Q(o_label6_data5[18]));
Q_FDP4EP \o_label6_data5_REG[19] ( .CK(clk), .CE(n184), .R(n261), .D(n25), .Q(o_label6_data5[19]));
Q_FDP4EP \o_label6_data5_REG[20] ( .CK(clk), .CE(n184), .R(n261), .D(n26), .Q(o_label6_data5[20]));
Q_FDP4EP \o_label6_data5_REG[21] ( .CK(clk), .CE(n184), .R(n261), .D(n27), .Q(o_label6_data5[21]));
Q_FDP4EP \o_label6_data5_REG[22] ( .CK(clk), .CE(n184), .R(n261), .D(n28), .Q(o_label6_data5[22]));
Q_FDP4EP \o_label6_data5_REG[23] ( .CK(clk), .CE(n184), .R(n261), .D(n29), .Q(o_label6_data5[23]));
Q_FDP4EP \o_label6_data5_REG[24] ( .CK(clk), .CE(n184), .R(n261), .D(n30), .Q(o_label6_data5[24]));
Q_FDP4EP \o_label6_data5_REG[25] ( .CK(clk), .CE(n184), .R(n261), .D(n31), .Q(o_label6_data5[25]));
Q_FDP4EP \o_label6_data5_REG[26] ( .CK(clk), .CE(n184), .R(n261), .D(n32), .Q(o_label6_data5[26]));
Q_FDP4EP \o_label6_data5_REG[27] ( .CK(clk), .CE(n184), .R(n261), .D(n33), .Q(o_label6_data5[27]));
Q_FDP4EP \o_label6_data5_REG[28] ( .CK(clk), .CE(n184), .R(n261), .D(n34), .Q(o_label6_data5[28]));
Q_FDP4EP \o_label6_data5_REG[29] ( .CK(clk), .CE(n184), .R(n261), .D(n35), .Q(o_label6_data5[29]));
Q_FDP4EP \o_label6_data5_REG[30] ( .CK(clk), .CE(n184), .R(n261), .D(n36), .Q(o_label6_data5[30]));
Q_FDP4EP \o_label6_data5_REG[31] ( .CK(clk), .CE(n184), .R(n261), .D(n37), .Q(o_label6_data5[31]));
Q_FDP4EP \o_label6_data6_REG[0] ( .CK(clk), .CE(n183), .R(n261), .D(n6), .Q(o_label6_data6[0]));
Q_FDP4EP \o_label6_data6_REG[1] ( .CK(clk), .CE(n183), .R(n261), .D(n7), .Q(o_label6_data6[1]));
Q_FDP4EP \o_label6_data6_REG[2] ( .CK(clk), .CE(n183), .R(n261), .D(n8), .Q(o_label6_data6[2]));
Q_FDP4EP \o_label6_data6_REG[3] ( .CK(clk), .CE(n183), .R(n261), .D(n9), .Q(o_label6_data6[3]));
Q_FDP4EP \o_label6_data6_REG[4] ( .CK(clk), .CE(n183), .R(n261), .D(n10), .Q(o_label6_data6[4]));
Q_FDP4EP \o_label6_data6_REG[5] ( .CK(clk), .CE(n183), .R(n261), .D(n11), .Q(o_label6_data6[5]));
Q_FDP4EP \o_label6_data6_REG[6] ( .CK(clk), .CE(n183), .R(n261), .D(n12), .Q(o_label6_data6[6]));
Q_FDP4EP \o_label6_data6_REG[7] ( .CK(clk), .CE(n183), .R(n261), .D(n13), .Q(o_label6_data6[7]));
Q_FDP4EP \o_label6_data6_REG[8] ( .CK(clk), .CE(n183), .R(n261), .D(n14), .Q(o_label6_data6[8]));
Q_FDP4EP \o_label6_data6_REG[9] ( .CK(clk), .CE(n183), .R(n261), .D(n15), .Q(o_label6_data6[9]));
Q_FDP4EP \o_label6_data6_REG[10] ( .CK(clk), .CE(n183), .R(n261), .D(n16), .Q(o_label6_data6[10]));
Q_FDP4EP \o_label6_data6_REG[11] ( .CK(clk), .CE(n183), .R(n261), .D(n17), .Q(o_label6_data6[11]));
Q_FDP4EP \o_label6_data6_REG[12] ( .CK(clk), .CE(n183), .R(n261), .D(n18), .Q(o_label6_data6[12]));
Q_FDP4EP \o_label6_data6_REG[13] ( .CK(clk), .CE(n183), .R(n261), .D(n19), .Q(o_label6_data6[13]));
Q_FDP4EP \o_label6_data6_REG[14] ( .CK(clk), .CE(n183), .R(n261), .D(n20), .Q(o_label6_data6[14]));
Q_FDP4EP \o_label6_data6_REG[15] ( .CK(clk), .CE(n183), .R(n261), .D(n21), .Q(o_label6_data6[15]));
Q_FDP4EP \o_label6_data6_REG[16] ( .CK(clk), .CE(n183), .R(n261), .D(n22), .Q(o_label6_data6[16]));
Q_FDP4EP \o_label6_data6_REG[17] ( .CK(clk), .CE(n183), .R(n261), .D(n23), .Q(o_label6_data6[17]));
Q_FDP4EP \o_label6_data6_REG[18] ( .CK(clk), .CE(n183), .R(n261), .D(n24), .Q(o_label6_data6[18]));
Q_FDP4EP \o_label6_data6_REG[19] ( .CK(clk), .CE(n183), .R(n261), .D(n25), .Q(o_label6_data6[19]));
Q_FDP4EP \o_label6_data6_REG[20] ( .CK(clk), .CE(n183), .R(n261), .D(n26), .Q(o_label6_data6[20]));
Q_FDP4EP \o_label6_data6_REG[21] ( .CK(clk), .CE(n183), .R(n261), .D(n27), .Q(o_label6_data6[21]));
Q_FDP4EP \o_label6_data6_REG[22] ( .CK(clk), .CE(n183), .R(n261), .D(n28), .Q(o_label6_data6[22]));
Q_FDP4EP \o_label6_data6_REG[23] ( .CK(clk), .CE(n183), .R(n261), .D(n29), .Q(o_label6_data6[23]));
Q_FDP4EP \o_label6_data6_REG[24] ( .CK(clk), .CE(n183), .R(n261), .D(n30), .Q(o_label6_data6[24]));
Q_FDP4EP \o_label6_data6_REG[25] ( .CK(clk), .CE(n183), .R(n261), .D(n31), .Q(o_label6_data6[25]));
Q_FDP4EP \o_label6_data6_REG[26] ( .CK(clk), .CE(n183), .R(n261), .D(n32), .Q(o_label6_data6[26]));
Q_FDP4EP \o_label6_data6_REG[27] ( .CK(clk), .CE(n183), .R(n261), .D(n33), .Q(o_label6_data6[27]));
Q_FDP4EP \o_label6_data6_REG[28] ( .CK(clk), .CE(n183), .R(n261), .D(n34), .Q(o_label6_data6[28]));
Q_FDP4EP \o_label6_data6_REG[29] ( .CK(clk), .CE(n183), .R(n261), .D(n35), .Q(o_label6_data6[29]));
Q_FDP4EP \o_label6_data6_REG[30] ( .CK(clk), .CE(n183), .R(n261), .D(n36), .Q(o_label6_data6[30]));
Q_FDP4EP \o_label6_data6_REG[31] ( .CK(clk), .CE(n183), .R(n261), .D(n37), .Q(o_label6_data6[31]));
Q_FDP4EP \o_label6_data7_REG[0] ( .CK(clk), .CE(n182), .R(n261), .D(n6), .Q(o_label6_data7[0]));
Q_FDP4EP \o_label6_data7_REG[1] ( .CK(clk), .CE(n182), .R(n261), .D(n7), .Q(o_label6_data7[1]));
Q_FDP4EP \o_label6_data7_REG[2] ( .CK(clk), .CE(n182), .R(n261), .D(n8), .Q(o_label6_data7[2]));
Q_FDP4EP \o_label6_data7_REG[3] ( .CK(clk), .CE(n182), .R(n261), .D(n9), .Q(o_label6_data7[3]));
Q_FDP4EP \o_label6_data7_REG[4] ( .CK(clk), .CE(n182), .R(n261), .D(n10), .Q(o_label6_data7[4]));
Q_FDP4EP \o_label6_data7_REG[5] ( .CK(clk), .CE(n182), .R(n261), .D(n11), .Q(o_label6_data7[5]));
Q_FDP4EP \o_label6_data7_REG[6] ( .CK(clk), .CE(n182), .R(n261), .D(n12), .Q(o_label6_data7[6]));
Q_FDP4EP \o_label6_data7_REG[7] ( .CK(clk), .CE(n182), .R(n261), .D(n13), .Q(o_label6_data7[7]));
Q_FDP4EP \o_label6_data7_REG[8] ( .CK(clk), .CE(n182), .R(n261), .D(n14), .Q(o_label6_data7[8]));
Q_FDP4EP \o_label6_data7_REG[9] ( .CK(clk), .CE(n182), .R(n261), .D(n15), .Q(o_label6_data7[9]));
Q_FDP4EP \o_label6_data7_REG[10] ( .CK(clk), .CE(n182), .R(n261), .D(n16), .Q(o_label6_data7[10]));
Q_FDP4EP \o_label6_data7_REG[11] ( .CK(clk), .CE(n182), .R(n261), .D(n17), .Q(o_label6_data7[11]));
Q_FDP4EP \o_label6_data7_REG[12] ( .CK(clk), .CE(n182), .R(n261), .D(n18), .Q(o_label6_data7[12]));
Q_FDP4EP \o_label6_data7_REG[13] ( .CK(clk), .CE(n182), .R(n261), .D(n19), .Q(o_label6_data7[13]));
Q_FDP4EP \o_label6_data7_REG[14] ( .CK(clk), .CE(n182), .R(n261), .D(n20), .Q(o_label6_data7[14]));
Q_FDP4EP \o_label6_data7_REG[15] ( .CK(clk), .CE(n182), .R(n261), .D(n21), .Q(o_label6_data7[15]));
Q_FDP4EP \o_label6_data7_REG[16] ( .CK(clk), .CE(n182), .R(n261), .D(n22), .Q(o_label6_data7[16]));
Q_FDP4EP \o_label6_data7_REG[17] ( .CK(clk), .CE(n182), .R(n261), .D(n23), .Q(o_label6_data7[17]));
Q_FDP4EP \o_label6_data7_REG[18] ( .CK(clk), .CE(n182), .R(n261), .D(n24), .Q(o_label6_data7[18]));
Q_FDP4EP \o_label6_data7_REG[19] ( .CK(clk), .CE(n182), .R(n261), .D(n25), .Q(o_label6_data7[19]));
Q_FDP4EP \o_label6_data7_REG[20] ( .CK(clk), .CE(n182), .R(n261), .D(n26), .Q(o_label6_data7[20]));
Q_FDP4EP \o_label6_data7_REG[21] ( .CK(clk), .CE(n182), .R(n261), .D(n27), .Q(o_label6_data7[21]));
Q_FDP4EP \o_label6_data7_REG[22] ( .CK(clk), .CE(n182), .R(n261), .D(n28), .Q(o_label6_data7[22]));
Q_FDP4EP \o_label6_data7_REG[23] ( .CK(clk), .CE(n182), .R(n261), .D(n29), .Q(o_label6_data7[23]));
Q_FDP4EP \o_label6_data7_REG[24] ( .CK(clk), .CE(n182), .R(n261), .D(n30), .Q(o_label6_data7[24]));
Q_FDP4EP \o_label6_data7_REG[25] ( .CK(clk), .CE(n182), .R(n261), .D(n31), .Q(o_label6_data7[25]));
Q_FDP4EP \o_label6_data7_REG[26] ( .CK(clk), .CE(n182), .R(n261), .D(n32), .Q(o_label6_data7[26]));
Q_FDP4EP \o_label6_data7_REG[27] ( .CK(clk), .CE(n182), .R(n261), .D(n33), .Q(o_label6_data7[27]));
Q_FDP4EP \o_label6_data7_REG[28] ( .CK(clk), .CE(n182), .R(n261), .D(n34), .Q(o_label6_data7[28]));
Q_FDP4EP \o_label6_data7_REG[29] ( .CK(clk), .CE(n182), .R(n261), .D(n35), .Q(o_label6_data7[29]));
Q_FDP4EP \o_label6_data7_REG[30] ( .CK(clk), .CE(n182), .R(n261), .D(n36), .Q(o_label6_data7[30]));
Q_FDP4EP \o_label6_data7_REG[31] ( .CK(clk), .CE(n182), .R(n261), .D(n37), .Q(o_label6_data7[31]));
Q_FDP4EP \o_label6_config_REG[0] ( .CK(clk), .CE(n181), .R(n261), .D(n6), .Q(o_label6_config[0]));
Q_FDP4EP \o_label6_config_REG[1] ( .CK(clk), .CE(n181), .R(n261), .D(n7), .Q(o_label6_config[1]));
Q_FDP4EP \o_label6_config_REG[2] ( .CK(clk), .CE(n181), .R(n261), .D(n8), .Q(o_label6_config[2]));
Q_FDP4EP \o_label6_config_REG[3] ( .CK(clk), .CE(n181), .R(n261), .D(n9), .Q(o_label6_config[3]));
Q_FDP4EP \o_label6_config_REG[4] ( .CK(clk), .CE(n181), .R(n261), .D(n10), .Q(o_label6_config[4]));
Q_FDP4EP \o_label6_config_REG[5] ( .CK(clk), .CE(n181), .R(n261), .D(n11), .Q(o_label6_config[5]));
Q_FDP4EP \o_label6_config_REG[6] ( .CK(clk), .CE(n181), .R(n261), .D(n12), .Q(o_label6_config[6]));
Q_FDP4EP \o_label6_config_REG[7] ( .CK(clk), .CE(n181), .R(n261), .D(n13), .Q(o_label6_config[7]));
Q_FDP4EP \o_label6_config_REG[9] ( .CK(clk), .CE(n181), .R(n261), .D(n31), .Q(o_label6_config[9]));
Q_FDP4EP \o_label6_config_REG[10] ( .CK(clk), .CE(n181), .R(n261), .D(n32), .Q(o_label6_config[10]));
Q_FDP4EP \o_label6_config_REG[11] ( .CK(clk), .CE(n181), .R(n261), .D(n33), .Q(o_label6_config[11]));
Q_FDP4EP \o_label6_config_REG[12] ( .CK(clk), .CE(n181), .R(n261), .D(n34), .Q(o_label6_config[12]));
Q_FDP4EP \o_label6_config_REG[13] ( .CK(clk), .CE(n181), .R(n261), .D(n35), .Q(o_label6_config[13]));
Q_FDP4EP \o_label6_config_REG[14] ( .CK(clk), .CE(n181), .R(n261), .D(n36), .Q(o_label6_config[14]));
Q_FDP4EP \o_label6_config_REG[15] ( .CK(clk), .CE(n181), .R(n261), .D(n37), .Q(o_label6_config[15]));
Q_FDP4EP \o_label5_data0_REG[0] ( .CK(clk), .CE(n180), .R(n261), .D(n6), .Q(o_label5_data0[0]));
Q_FDP4EP \o_label5_data0_REG[1] ( .CK(clk), .CE(n180), .R(n261), .D(n7), .Q(o_label5_data0[1]));
Q_FDP4EP \o_label5_data0_REG[2] ( .CK(clk), .CE(n180), .R(n261), .D(n8), .Q(o_label5_data0[2]));
Q_FDP4EP \o_label5_data0_REG[3] ( .CK(clk), .CE(n180), .R(n261), .D(n9), .Q(o_label5_data0[3]));
Q_FDP4EP \o_label5_data0_REG[4] ( .CK(clk), .CE(n180), .R(n261), .D(n10), .Q(o_label5_data0[4]));
Q_FDP4EP \o_label5_data0_REG[5] ( .CK(clk), .CE(n180), .R(n261), .D(n11), .Q(o_label5_data0[5]));
Q_FDP4EP \o_label5_data0_REG[6] ( .CK(clk), .CE(n180), .R(n261), .D(n12), .Q(o_label5_data0[6]));
Q_FDP4EP \o_label5_data0_REG[7] ( .CK(clk), .CE(n180), .R(n261), .D(n13), .Q(o_label5_data0[7]));
Q_FDP4EP \o_label5_data0_REG[8] ( .CK(clk), .CE(n180), .R(n261), .D(n14), .Q(o_label5_data0[8]));
Q_FDP4EP \o_label5_data0_REG[9] ( .CK(clk), .CE(n180), .R(n261), .D(n15), .Q(o_label5_data0[9]));
Q_FDP4EP \o_label5_data0_REG[10] ( .CK(clk), .CE(n180), .R(n261), .D(n16), .Q(o_label5_data0[10]));
Q_FDP4EP \o_label5_data0_REG[11] ( .CK(clk), .CE(n180), .R(n261), .D(n17), .Q(o_label5_data0[11]));
Q_FDP4EP \o_label5_data0_REG[12] ( .CK(clk), .CE(n180), .R(n261), .D(n18), .Q(o_label5_data0[12]));
Q_FDP4EP \o_label5_data0_REG[13] ( .CK(clk), .CE(n180), .R(n261), .D(n19), .Q(o_label5_data0[13]));
Q_FDP4EP \o_label5_data0_REG[14] ( .CK(clk), .CE(n180), .R(n261), .D(n20), .Q(o_label5_data0[14]));
Q_FDP4EP \o_label5_data0_REG[15] ( .CK(clk), .CE(n180), .R(n261), .D(n21), .Q(o_label5_data0[15]));
Q_FDP4EP \o_label5_data0_REG[16] ( .CK(clk), .CE(n180), .R(n261), .D(n22), .Q(o_label5_data0[16]));
Q_FDP4EP \o_label5_data0_REG[17] ( .CK(clk), .CE(n180), .R(n261), .D(n23), .Q(o_label5_data0[17]));
Q_FDP4EP \o_label5_data0_REG[18] ( .CK(clk), .CE(n180), .R(n261), .D(n24), .Q(o_label5_data0[18]));
Q_FDP4EP \o_label5_data0_REG[19] ( .CK(clk), .CE(n180), .R(n261), .D(n25), .Q(o_label5_data0[19]));
Q_FDP4EP \o_label5_data0_REG[20] ( .CK(clk), .CE(n180), .R(n261), .D(n26), .Q(o_label5_data0[20]));
Q_FDP4EP \o_label5_data0_REG[21] ( .CK(clk), .CE(n180), .R(n261), .D(n27), .Q(o_label5_data0[21]));
Q_FDP4EP \o_label5_data0_REG[22] ( .CK(clk), .CE(n180), .R(n261), .D(n28), .Q(o_label5_data0[22]));
Q_FDP4EP \o_label5_data0_REG[23] ( .CK(clk), .CE(n180), .R(n261), .D(n29), .Q(o_label5_data0[23]));
Q_FDP4EP \o_label5_data0_REG[24] ( .CK(clk), .CE(n180), .R(n261), .D(n30), .Q(o_label5_data0[24]));
Q_FDP4EP \o_label5_data0_REG[25] ( .CK(clk), .CE(n180), .R(n261), .D(n31), .Q(o_label5_data0[25]));
Q_FDP4EP \o_label5_data0_REG[26] ( .CK(clk), .CE(n180), .R(n261), .D(n32), .Q(o_label5_data0[26]));
Q_FDP4EP \o_label5_data0_REG[27] ( .CK(clk), .CE(n180), .R(n261), .D(n33), .Q(o_label5_data0[27]));
Q_FDP4EP \o_label5_data0_REG[28] ( .CK(clk), .CE(n180), .R(n261), .D(n34), .Q(o_label5_data0[28]));
Q_FDP4EP \o_label5_data0_REG[29] ( .CK(clk), .CE(n180), .R(n261), .D(n35), .Q(o_label5_data0[29]));
Q_FDP4EP \o_label5_data0_REG[30] ( .CK(clk), .CE(n180), .R(n261), .D(n36), .Q(o_label5_data0[30]));
Q_FDP4EP \o_label5_data0_REG[31] ( .CK(clk), .CE(n180), .R(n261), .D(n37), .Q(o_label5_data0[31]));
Q_FDP4EP \o_label5_data1_REG[0] ( .CK(clk), .CE(n179), .R(n261), .D(n6), .Q(o_label5_data1[0]));
Q_FDP4EP \o_label5_data1_REG[1] ( .CK(clk), .CE(n179), .R(n261), .D(n7), .Q(o_label5_data1[1]));
Q_FDP4EP \o_label5_data1_REG[2] ( .CK(clk), .CE(n179), .R(n261), .D(n8), .Q(o_label5_data1[2]));
Q_FDP4EP \o_label5_data1_REG[3] ( .CK(clk), .CE(n179), .R(n261), .D(n9), .Q(o_label5_data1[3]));
Q_FDP4EP \o_label5_data1_REG[4] ( .CK(clk), .CE(n179), .R(n261), .D(n10), .Q(o_label5_data1[4]));
Q_FDP4EP \o_label5_data1_REG[5] ( .CK(clk), .CE(n179), .R(n261), .D(n11), .Q(o_label5_data1[5]));
Q_FDP4EP \o_label5_data1_REG[6] ( .CK(clk), .CE(n179), .R(n261), .D(n12), .Q(o_label5_data1[6]));
Q_FDP4EP \o_label5_data1_REG[7] ( .CK(clk), .CE(n179), .R(n261), .D(n13), .Q(o_label5_data1[7]));
Q_FDP4EP \o_label5_data1_REG[8] ( .CK(clk), .CE(n179), .R(n261), .D(n14), .Q(o_label5_data1[8]));
Q_FDP4EP \o_label5_data1_REG[9] ( .CK(clk), .CE(n179), .R(n261), .D(n15), .Q(o_label5_data1[9]));
Q_FDP4EP \o_label5_data1_REG[10] ( .CK(clk), .CE(n179), .R(n261), .D(n16), .Q(o_label5_data1[10]));
Q_FDP4EP \o_label5_data1_REG[11] ( .CK(clk), .CE(n179), .R(n261), .D(n17), .Q(o_label5_data1[11]));
Q_FDP4EP \o_label5_data1_REG[12] ( .CK(clk), .CE(n179), .R(n261), .D(n18), .Q(o_label5_data1[12]));
Q_FDP4EP \o_label5_data1_REG[13] ( .CK(clk), .CE(n179), .R(n261), .D(n19), .Q(o_label5_data1[13]));
Q_FDP4EP \o_label5_data1_REG[14] ( .CK(clk), .CE(n179), .R(n261), .D(n20), .Q(o_label5_data1[14]));
Q_FDP4EP \o_label5_data1_REG[15] ( .CK(clk), .CE(n179), .R(n261), .D(n21), .Q(o_label5_data1[15]));
Q_FDP4EP \o_label5_data1_REG[16] ( .CK(clk), .CE(n179), .R(n261), .D(n22), .Q(o_label5_data1[16]));
Q_FDP4EP \o_label5_data1_REG[17] ( .CK(clk), .CE(n179), .R(n261), .D(n23), .Q(o_label5_data1[17]));
Q_FDP4EP \o_label5_data1_REG[18] ( .CK(clk), .CE(n179), .R(n261), .D(n24), .Q(o_label5_data1[18]));
Q_FDP4EP \o_label5_data1_REG[19] ( .CK(clk), .CE(n179), .R(n261), .D(n25), .Q(o_label5_data1[19]));
Q_FDP4EP \o_label5_data1_REG[20] ( .CK(clk), .CE(n179), .R(n261), .D(n26), .Q(o_label5_data1[20]));
Q_FDP4EP \o_label5_data1_REG[21] ( .CK(clk), .CE(n179), .R(n261), .D(n27), .Q(o_label5_data1[21]));
Q_FDP4EP \o_label5_data1_REG[22] ( .CK(clk), .CE(n179), .R(n261), .D(n28), .Q(o_label5_data1[22]));
Q_FDP4EP \o_label5_data1_REG[23] ( .CK(clk), .CE(n179), .R(n261), .D(n29), .Q(o_label5_data1[23]));
Q_FDP4EP \o_label5_data1_REG[24] ( .CK(clk), .CE(n179), .R(n261), .D(n30), .Q(o_label5_data1[24]));
Q_FDP4EP \o_label5_data1_REG[25] ( .CK(clk), .CE(n179), .R(n261), .D(n31), .Q(o_label5_data1[25]));
Q_FDP4EP \o_label5_data1_REG[26] ( .CK(clk), .CE(n179), .R(n261), .D(n32), .Q(o_label5_data1[26]));
Q_FDP4EP \o_label5_data1_REG[27] ( .CK(clk), .CE(n179), .R(n261), .D(n33), .Q(o_label5_data1[27]));
Q_FDP4EP \o_label5_data1_REG[28] ( .CK(clk), .CE(n179), .R(n261), .D(n34), .Q(o_label5_data1[28]));
Q_FDP4EP \o_label5_data1_REG[29] ( .CK(clk), .CE(n179), .R(n261), .D(n35), .Q(o_label5_data1[29]));
Q_FDP4EP \o_label5_data1_REG[30] ( .CK(clk), .CE(n179), .R(n261), .D(n36), .Q(o_label5_data1[30]));
Q_FDP4EP \o_label5_data1_REG[31] ( .CK(clk), .CE(n179), .R(n261), .D(n37), .Q(o_label5_data1[31]));
Q_FDP4EP \o_label5_data2_REG[0] ( .CK(clk), .CE(n178), .R(n261), .D(n6), .Q(o_label5_data2[0]));
Q_FDP4EP \o_label5_data2_REG[1] ( .CK(clk), .CE(n178), .R(n261), .D(n7), .Q(o_label5_data2[1]));
Q_FDP4EP \o_label5_data2_REG[2] ( .CK(clk), .CE(n178), .R(n261), .D(n8), .Q(o_label5_data2[2]));
Q_FDP4EP \o_label5_data2_REG[3] ( .CK(clk), .CE(n178), .R(n261), .D(n9), .Q(o_label5_data2[3]));
Q_FDP4EP \o_label5_data2_REG[4] ( .CK(clk), .CE(n178), .R(n261), .D(n10), .Q(o_label5_data2[4]));
Q_FDP4EP \o_label5_data2_REG[5] ( .CK(clk), .CE(n178), .R(n261), .D(n11), .Q(o_label5_data2[5]));
Q_FDP4EP \o_label5_data2_REG[6] ( .CK(clk), .CE(n178), .R(n261), .D(n12), .Q(o_label5_data2[6]));
Q_FDP4EP \o_label5_data2_REG[7] ( .CK(clk), .CE(n178), .R(n261), .D(n13), .Q(o_label5_data2[7]));
Q_FDP4EP \o_label5_data2_REG[8] ( .CK(clk), .CE(n178), .R(n261), .D(n14), .Q(o_label5_data2[8]));
Q_FDP4EP \o_label5_data2_REG[9] ( .CK(clk), .CE(n178), .R(n261), .D(n15), .Q(o_label5_data2[9]));
Q_FDP4EP \o_label5_data2_REG[10] ( .CK(clk), .CE(n178), .R(n261), .D(n16), .Q(o_label5_data2[10]));
Q_FDP4EP \o_label5_data2_REG[11] ( .CK(clk), .CE(n178), .R(n261), .D(n17), .Q(o_label5_data2[11]));
Q_FDP4EP \o_label5_data2_REG[12] ( .CK(clk), .CE(n178), .R(n261), .D(n18), .Q(o_label5_data2[12]));
Q_FDP4EP \o_label5_data2_REG[13] ( .CK(clk), .CE(n178), .R(n261), .D(n19), .Q(o_label5_data2[13]));
Q_FDP4EP \o_label5_data2_REG[14] ( .CK(clk), .CE(n178), .R(n261), .D(n20), .Q(o_label5_data2[14]));
Q_FDP4EP \o_label5_data2_REG[15] ( .CK(clk), .CE(n178), .R(n261), .D(n21), .Q(o_label5_data2[15]));
Q_FDP4EP \o_label5_data2_REG[16] ( .CK(clk), .CE(n178), .R(n261), .D(n22), .Q(o_label5_data2[16]));
Q_FDP4EP \o_label5_data2_REG[17] ( .CK(clk), .CE(n178), .R(n261), .D(n23), .Q(o_label5_data2[17]));
Q_FDP4EP \o_label5_data2_REG[18] ( .CK(clk), .CE(n178), .R(n261), .D(n24), .Q(o_label5_data2[18]));
Q_FDP4EP \o_label5_data2_REG[19] ( .CK(clk), .CE(n178), .R(n261), .D(n25), .Q(o_label5_data2[19]));
Q_FDP4EP \o_label5_data2_REG[20] ( .CK(clk), .CE(n178), .R(n261), .D(n26), .Q(o_label5_data2[20]));
Q_FDP4EP \o_label5_data2_REG[21] ( .CK(clk), .CE(n178), .R(n261), .D(n27), .Q(o_label5_data2[21]));
Q_FDP4EP \o_label5_data2_REG[22] ( .CK(clk), .CE(n178), .R(n261), .D(n28), .Q(o_label5_data2[22]));
Q_FDP4EP \o_label5_data2_REG[23] ( .CK(clk), .CE(n178), .R(n261), .D(n29), .Q(o_label5_data2[23]));
Q_FDP4EP \o_label5_data2_REG[24] ( .CK(clk), .CE(n178), .R(n261), .D(n30), .Q(o_label5_data2[24]));
Q_FDP4EP \o_label5_data2_REG[25] ( .CK(clk), .CE(n178), .R(n261), .D(n31), .Q(o_label5_data2[25]));
Q_FDP4EP \o_label5_data2_REG[26] ( .CK(clk), .CE(n178), .R(n261), .D(n32), .Q(o_label5_data2[26]));
Q_FDP4EP \o_label5_data2_REG[27] ( .CK(clk), .CE(n178), .R(n261), .D(n33), .Q(o_label5_data2[27]));
Q_FDP4EP \o_label5_data2_REG[28] ( .CK(clk), .CE(n178), .R(n261), .D(n34), .Q(o_label5_data2[28]));
Q_FDP4EP \o_label5_data2_REG[29] ( .CK(clk), .CE(n178), .R(n261), .D(n35), .Q(o_label5_data2[29]));
Q_FDP4EP \o_label5_data2_REG[30] ( .CK(clk), .CE(n178), .R(n261), .D(n36), .Q(o_label5_data2[30]));
Q_FDP4EP \o_label5_data2_REG[31] ( .CK(clk), .CE(n178), .R(n261), .D(n37), .Q(o_label5_data2[31]));
Q_FDP4EP \o_label5_data3_REG[0] ( .CK(clk), .CE(n177), .R(n261), .D(n6), .Q(o_label5_data3[0]));
Q_FDP4EP \o_label5_data3_REG[1] ( .CK(clk), .CE(n177), .R(n261), .D(n7), .Q(o_label5_data3[1]));
Q_FDP4EP \o_label5_data3_REG[2] ( .CK(clk), .CE(n177), .R(n261), .D(n8), .Q(o_label5_data3[2]));
Q_FDP4EP \o_label5_data3_REG[3] ( .CK(clk), .CE(n177), .R(n261), .D(n9), .Q(o_label5_data3[3]));
Q_FDP4EP \o_label5_data3_REG[4] ( .CK(clk), .CE(n177), .R(n261), .D(n10), .Q(o_label5_data3[4]));
Q_FDP4EP \o_label5_data3_REG[5] ( .CK(clk), .CE(n177), .R(n261), .D(n11), .Q(o_label5_data3[5]));
Q_FDP4EP \o_label5_data3_REG[6] ( .CK(clk), .CE(n177), .R(n261), .D(n12), .Q(o_label5_data3[6]));
Q_FDP4EP \o_label5_data3_REG[7] ( .CK(clk), .CE(n177), .R(n261), .D(n13), .Q(o_label5_data3[7]));
Q_FDP4EP \o_label5_data3_REG[8] ( .CK(clk), .CE(n177), .R(n261), .D(n14), .Q(o_label5_data3[8]));
Q_FDP4EP \o_label5_data3_REG[9] ( .CK(clk), .CE(n177), .R(n261), .D(n15), .Q(o_label5_data3[9]));
Q_FDP4EP \o_label5_data3_REG[10] ( .CK(clk), .CE(n177), .R(n261), .D(n16), .Q(o_label5_data3[10]));
Q_FDP4EP \o_label5_data3_REG[11] ( .CK(clk), .CE(n177), .R(n261), .D(n17), .Q(o_label5_data3[11]));
Q_FDP4EP \o_label5_data3_REG[12] ( .CK(clk), .CE(n177), .R(n261), .D(n18), .Q(o_label5_data3[12]));
Q_FDP4EP \o_label5_data3_REG[13] ( .CK(clk), .CE(n177), .R(n261), .D(n19), .Q(o_label5_data3[13]));
Q_FDP4EP \o_label5_data3_REG[14] ( .CK(clk), .CE(n177), .R(n261), .D(n20), .Q(o_label5_data3[14]));
Q_FDP4EP \o_label5_data3_REG[15] ( .CK(clk), .CE(n177), .R(n261), .D(n21), .Q(o_label5_data3[15]));
Q_FDP4EP \o_label5_data3_REG[16] ( .CK(clk), .CE(n177), .R(n261), .D(n22), .Q(o_label5_data3[16]));
Q_FDP4EP \o_label5_data3_REG[17] ( .CK(clk), .CE(n177), .R(n261), .D(n23), .Q(o_label5_data3[17]));
Q_FDP4EP \o_label5_data3_REG[18] ( .CK(clk), .CE(n177), .R(n261), .D(n24), .Q(o_label5_data3[18]));
Q_FDP4EP \o_label5_data3_REG[19] ( .CK(clk), .CE(n177), .R(n261), .D(n25), .Q(o_label5_data3[19]));
Q_FDP4EP \o_label5_data3_REG[20] ( .CK(clk), .CE(n177), .R(n261), .D(n26), .Q(o_label5_data3[20]));
Q_FDP4EP \o_label5_data3_REG[21] ( .CK(clk), .CE(n177), .R(n261), .D(n27), .Q(o_label5_data3[21]));
Q_FDP4EP \o_label5_data3_REG[22] ( .CK(clk), .CE(n177), .R(n261), .D(n28), .Q(o_label5_data3[22]));
Q_FDP4EP \o_label5_data3_REG[23] ( .CK(clk), .CE(n177), .R(n261), .D(n29), .Q(o_label5_data3[23]));
Q_FDP4EP \o_label5_data3_REG[24] ( .CK(clk), .CE(n177), .R(n261), .D(n30), .Q(o_label5_data3[24]));
Q_FDP4EP \o_label5_data3_REG[25] ( .CK(clk), .CE(n177), .R(n261), .D(n31), .Q(o_label5_data3[25]));
Q_FDP4EP \o_label5_data3_REG[26] ( .CK(clk), .CE(n177), .R(n261), .D(n32), .Q(o_label5_data3[26]));
Q_FDP4EP \o_label5_data3_REG[27] ( .CK(clk), .CE(n177), .R(n261), .D(n33), .Q(o_label5_data3[27]));
Q_FDP4EP \o_label5_data3_REG[28] ( .CK(clk), .CE(n177), .R(n261), .D(n34), .Q(o_label5_data3[28]));
Q_FDP4EP \o_label5_data3_REG[29] ( .CK(clk), .CE(n177), .R(n261), .D(n35), .Q(o_label5_data3[29]));
Q_FDP4EP \o_label5_data3_REG[30] ( .CK(clk), .CE(n177), .R(n261), .D(n36), .Q(o_label5_data3[30]));
Q_FDP4EP \o_label5_data3_REG[31] ( .CK(clk), .CE(n177), .R(n261), .D(n37), .Q(o_label5_data3[31]));
Q_FDP4EP \o_label5_data4_REG[0] ( .CK(clk), .CE(n176), .R(n261), .D(n6), .Q(o_label5_data4[0]));
Q_FDP4EP \o_label5_data4_REG[1] ( .CK(clk), .CE(n176), .R(n261), .D(n7), .Q(o_label5_data4[1]));
Q_FDP4EP \o_label5_data4_REG[2] ( .CK(clk), .CE(n176), .R(n261), .D(n8), .Q(o_label5_data4[2]));
Q_FDP4EP \o_label5_data4_REG[3] ( .CK(clk), .CE(n176), .R(n261), .D(n9), .Q(o_label5_data4[3]));
Q_FDP4EP \o_label5_data4_REG[4] ( .CK(clk), .CE(n176), .R(n261), .D(n10), .Q(o_label5_data4[4]));
Q_FDP4EP \o_label5_data4_REG[5] ( .CK(clk), .CE(n176), .R(n261), .D(n11), .Q(o_label5_data4[5]));
Q_FDP4EP \o_label5_data4_REG[6] ( .CK(clk), .CE(n176), .R(n261), .D(n12), .Q(o_label5_data4[6]));
Q_FDP4EP \o_label5_data4_REG[7] ( .CK(clk), .CE(n176), .R(n261), .D(n13), .Q(o_label5_data4[7]));
Q_FDP4EP \o_label5_data4_REG[8] ( .CK(clk), .CE(n176), .R(n261), .D(n14), .Q(o_label5_data4[8]));
Q_FDP4EP \o_label5_data4_REG[9] ( .CK(clk), .CE(n176), .R(n261), .D(n15), .Q(o_label5_data4[9]));
Q_FDP4EP \o_label5_data4_REG[10] ( .CK(clk), .CE(n176), .R(n261), .D(n16), .Q(o_label5_data4[10]));
Q_FDP4EP \o_label5_data4_REG[11] ( .CK(clk), .CE(n176), .R(n261), .D(n17), .Q(o_label5_data4[11]));
Q_FDP4EP \o_label5_data4_REG[12] ( .CK(clk), .CE(n176), .R(n261), .D(n18), .Q(o_label5_data4[12]));
Q_FDP4EP \o_label5_data4_REG[13] ( .CK(clk), .CE(n176), .R(n261), .D(n19), .Q(o_label5_data4[13]));
Q_FDP4EP \o_label5_data4_REG[14] ( .CK(clk), .CE(n176), .R(n261), .D(n20), .Q(o_label5_data4[14]));
Q_FDP4EP \o_label5_data4_REG[15] ( .CK(clk), .CE(n176), .R(n261), .D(n21), .Q(o_label5_data4[15]));
Q_FDP4EP \o_label5_data4_REG[16] ( .CK(clk), .CE(n176), .R(n261), .D(n22), .Q(o_label5_data4[16]));
Q_FDP4EP \o_label5_data4_REG[17] ( .CK(clk), .CE(n176), .R(n261), .D(n23), .Q(o_label5_data4[17]));
Q_FDP4EP \o_label5_data4_REG[18] ( .CK(clk), .CE(n176), .R(n261), .D(n24), .Q(o_label5_data4[18]));
Q_FDP4EP \o_label5_data4_REG[19] ( .CK(clk), .CE(n176), .R(n261), .D(n25), .Q(o_label5_data4[19]));
Q_FDP4EP \o_label5_data4_REG[20] ( .CK(clk), .CE(n176), .R(n261), .D(n26), .Q(o_label5_data4[20]));
Q_FDP4EP \o_label5_data4_REG[21] ( .CK(clk), .CE(n176), .R(n261), .D(n27), .Q(o_label5_data4[21]));
Q_FDP4EP \o_label5_data4_REG[22] ( .CK(clk), .CE(n176), .R(n261), .D(n28), .Q(o_label5_data4[22]));
Q_FDP4EP \o_label5_data4_REG[23] ( .CK(clk), .CE(n176), .R(n261), .D(n29), .Q(o_label5_data4[23]));
Q_FDP4EP \o_label5_data4_REG[24] ( .CK(clk), .CE(n176), .R(n261), .D(n30), .Q(o_label5_data4[24]));
Q_FDP4EP \o_label5_data4_REG[25] ( .CK(clk), .CE(n176), .R(n261), .D(n31), .Q(o_label5_data4[25]));
Q_FDP4EP \o_label5_data4_REG[26] ( .CK(clk), .CE(n176), .R(n261), .D(n32), .Q(o_label5_data4[26]));
Q_FDP4EP \o_label5_data4_REG[27] ( .CK(clk), .CE(n176), .R(n261), .D(n33), .Q(o_label5_data4[27]));
Q_FDP4EP \o_label5_data4_REG[28] ( .CK(clk), .CE(n176), .R(n261), .D(n34), .Q(o_label5_data4[28]));
Q_FDP4EP \o_label5_data4_REG[29] ( .CK(clk), .CE(n176), .R(n261), .D(n35), .Q(o_label5_data4[29]));
Q_FDP4EP \o_label5_data4_REG[30] ( .CK(clk), .CE(n176), .R(n261), .D(n36), .Q(o_label5_data4[30]));
Q_FDP4EP \o_label5_data4_REG[31] ( .CK(clk), .CE(n176), .R(n261), .D(n37), .Q(o_label5_data4[31]));
Q_FDP4EP \o_label5_data5_REG[0] ( .CK(clk), .CE(n175), .R(n261), .D(n6), .Q(o_label5_data5[0]));
Q_FDP4EP \o_label5_data5_REG[1] ( .CK(clk), .CE(n175), .R(n261), .D(n7), .Q(o_label5_data5[1]));
Q_FDP4EP \o_label5_data5_REG[2] ( .CK(clk), .CE(n175), .R(n261), .D(n8), .Q(o_label5_data5[2]));
Q_FDP4EP \o_label5_data5_REG[3] ( .CK(clk), .CE(n175), .R(n261), .D(n9), .Q(o_label5_data5[3]));
Q_FDP4EP \o_label5_data5_REG[4] ( .CK(clk), .CE(n175), .R(n261), .D(n10), .Q(o_label5_data5[4]));
Q_FDP4EP \o_label5_data5_REG[5] ( .CK(clk), .CE(n175), .R(n261), .D(n11), .Q(o_label5_data5[5]));
Q_FDP4EP \o_label5_data5_REG[6] ( .CK(clk), .CE(n175), .R(n261), .D(n12), .Q(o_label5_data5[6]));
Q_FDP4EP \o_label5_data5_REG[7] ( .CK(clk), .CE(n175), .R(n261), .D(n13), .Q(o_label5_data5[7]));
Q_FDP4EP \o_label5_data5_REG[8] ( .CK(clk), .CE(n175), .R(n261), .D(n14), .Q(o_label5_data5[8]));
Q_FDP4EP \o_label5_data5_REG[9] ( .CK(clk), .CE(n175), .R(n261), .D(n15), .Q(o_label5_data5[9]));
Q_FDP4EP \o_label5_data5_REG[10] ( .CK(clk), .CE(n175), .R(n261), .D(n16), .Q(o_label5_data5[10]));
Q_FDP4EP \o_label5_data5_REG[11] ( .CK(clk), .CE(n175), .R(n261), .D(n17), .Q(o_label5_data5[11]));
Q_FDP4EP \o_label5_data5_REG[12] ( .CK(clk), .CE(n175), .R(n261), .D(n18), .Q(o_label5_data5[12]));
Q_FDP4EP \o_label5_data5_REG[13] ( .CK(clk), .CE(n175), .R(n261), .D(n19), .Q(o_label5_data5[13]));
Q_FDP4EP \o_label5_data5_REG[14] ( .CK(clk), .CE(n175), .R(n261), .D(n20), .Q(o_label5_data5[14]));
Q_FDP4EP \o_label5_data5_REG[15] ( .CK(clk), .CE(n175), .R(n261), .D(n21), .Q(o_label5_data5[15]));
Q_FDP4EP \o_label5_data5_REG[16] ( .CK(clk), .CE(n175), .R(n261), .D(n22), .Q(o_label5_data5[16]));
Q_FDP4EP \o_label5_data5_REG[17] ( .CK(clk), .CE(n175), .R(n261), .D(n23), .Q(o_label5_data5[17]));
Q_FDP4EP \o_label5_data5_REG[18] ( .CK(clk), .CE(n175), .R(n261), .D(n24), .Q(o_label5_data5[18]));
Q_FDP4EP \o_label5_data5_REG[19] ( .CK(clk), .CE(n175), .R(n261), .D(n25), .Q(o_label5_data5[19]));
Q_FDP4EP \o_label5_data5_REG[20] ( .CK(clk), .CE(n175), .R(n261), .D(n26), .Q(o_label5_data5[20]));
Q_FDP4EP \o_label5_data5_REG[21] ( .CK(clk), .CE(n175), .R(n261), .D(n27), .Q(o_label5_data5[21]));
Q_FDP4EP \o_label5_data5_REG[22] ( .CK(clk), .CE(n175), .R(n261), .D(n28), .Q(o_label5_data5[22]));
Q_FDP4EP \o_label5_data5_REG[23] ( .CK(clk), .CE(n175), .R(n261), .D(n29), .Q(o_label5_data5[23]));
Q_FDP4EP \o_label5_data5_REG[24] ( .CK(clk), .CE(n175), .R(n261), .D(n30), .Q(o_label5_data5[24]));
Q_FDP4EP \o_label5_data5_REG[25] ( .CK(clk), .CE(n175), .R(n261), .D(n31), .Q(o_label5_data5[25]));
Q_FDP4EP \o_label5_data5_REG[26] ( .CK(clk), .CE(n175), .R(n261), .D(n32), .Q(o_label5_data5[26]));
Q_FDP4EP \o_label5_data5_REG[27] ( .CK(clk), .CE(n175), .R(n261), .D(n33), .Q(o_label5_data5[27]));
Q_FDP4EP \o_label5_data5_REG[28] ( .CK(clk), .CE(n175), .R(n261), .D(n34), .Q(o_label5_data5[28]));
Q_FDP4EP \o_label5_data5_REG[29] ( .CK(clk), .CE(n175), .R(n261), .D(n35), .Q(o_label5_data5[29]));
Q_FDP4EP \o_label5_data5_REG[30] ( .CK(clk), .CE(n175), .R(n261), .D(n36), .Q(o_label5_data5[30]));
Q_FDP4EP \o_label5_data5_REG[31] ( .CK(clk), .CE(n175), .R(n261), .D(n37), .Q(o_label5_data5[31]));
Q_FDP4EP \o_label5_data6_REG[0] ( .CK(clk), .CE(n174), .R(n261), .D(n6), .Q(o_label5_data6[0]));
Q_FDP4EP \o_label5_data6_REG[1] ( .CK(clk), .CE(n174), .R(n261), .D(n7), .Q(o_label5_data6[1]));
Q_FDP4EP \o_label5_data6_REG[2] ( .CK(clk), .CE(n174), .R(n261), .D(n8), .Q(o_label5_data6[2]));
Q_FDP4EP \o_label5_data6_REG[3] ( .CK(clk), .CE(n174), .R(n261), .D(n9), .Q(o_label5_data6[3]));
Q_FDP4EP \o_label5_data6_REG[4] ( .CK(clk), .CE(n174), .R(n261), .D(n10), .Q(o_label5_data6[4]));
Q_FDP4EP \o_label5_data6_REG[5] ( .CK(clk), .CE(n174), .R(n261), .D(n11), .Q(o_label5_data6[5]));
Q_FDP4EP \o_label5_data6_REG[6] ( .CK(clk), .CE(n174), .R(n261), .D(n12), .Q(o_label5_data6[6]));
Q_FDP4EP \o_label5_data6_REG[7] ( .CK(clk), .CE(n174), .R(n261), .D(n13), .Q(o_label5_data6[7]));
Q_FDP4EP \o_label5_data6_REG[8] ( .CK(clk), .CE(n174), .R(n261), .D(n14), .Q(o_label5_data6[8]));
Q_FDP4EP \o_label5_data6_REG[9] ( .CK(clk), .CE(n174), .R(n261), .D(n15), .Q(o_label5_data6[9]));
Q_FDP4EP \o_label5_data6_REG[10] ( .CK(clk), .CE(n174), .R(n261), .D(n16), .Q(o_label5_data6[10]));
Q_FDP4EP \o_label5_data6_REG[11] ( .CK(clk), .CE(n174), .R(n261), .D(n17), .Q(o_label5_data6[11]));
Q_FDP4EP \o_label5_data6_REG[12] ( .CK(clk), .CE(n174), .R(n261), .D(n18), .Q(o_label5_data6[12]));
Q_FDP4EP \o_label5_data6_REG[13] ( .CK(clk), .CE(n174), .R(n261), .D(n19), .Q(o_label5_data6[13]));
Q_FDP4EP \o_label5_data6_REG[14] ( .CK(clk), .CE(n174), .R(n261), .D(n20), .Q(o_label5_data6[14]));
Q_FDP4EP \o_label5_data6_REG[15] ( .CK(clk), .CE(n174), .R(n261), .D(n21), .Q(o_label5_data6[15]));
Q_FDP4EP \o_label5_data6_REG[16] ( .CK(clk), .CE(n174), .R(n261), .D(n22), .Q(o_label5_data6[16]));
Q_FDP4EP \o_label5_data6_REG[17] ( .CK(clk), .CE(n174), .R(n261), .D(n23), .Q(o_label5_data6[17]));
Q_FDP4EP \o_label5_data6_REG[18] ( .CK(clk), .CE(n174), .R(n261), .D(n24), .Q(o_label5_data6[18]));
Q_FDP4EP \o_label5_data6_REG[19] ( .CK(clk), .CE(n174), .R(n261), .D(n25), .Q(o_label5_data6[19]));
Q_FDP4EP \o_label5_data6_REG[20] ( .CK(clk), .CE(n174), .R(n261), .D(n26), .Q(o_label5_data6[20]));
Q_FDP4EP \o_label5_data6_REG[21] ( .CK(clk), .CE(n174), .R(n261), .D(n27), .Q(o_label5_data6[21]));
Q_FDP4EP \o_label5_data6_REG[22] ( .CK(clk), .CE(n174), .R(n261), .D(n28), .Q(o_label5_data6[22]));
Q_FDP4EP \o_label5_data6_REG[23] ( .CK(clk), .CE(n174), .R(n261), .D(n29), .Q(o_label5_data6[23]));
Q_FDP4EP \o_label5_data6_REG[24] ( .CK(clk), .CE(n174), .R(n261), .D(n30), .Q(o_label5_data6[24]));
Q_FDP4EP \o_label5_data6_REG[25] ( .CK(clk), .CE(n174), .R(n261), .D(n31), .Q(o_label5_data6[25]));
Q_FDP4EP \o_label5_data6_REG[26] ( .CK(clk), .CE(n174), .R(n261), .D(n32), .Q(o_label5_data6[26]));
Q_FDP4EP \o_label5_data6_REG[27] ( .CK(clk), .CE(n174), .R(n261), .D(n33), .Q(o_label5_data6[27]));
Q_FDP4EP \o_label5_data6_REG[28] ( .CK(clk), .CE(n174), .R(n261), .D(n34), .Q(o_label5_data6[28]));
Q_FDP4EP \o_label5_data6_REG[29] ( .CK(clk), .CE(n174), .R(n261), .D(n35), .Q(o_label5_data6[29]));
Q_FDP4EP \o_label5_data6_REG[30] ( .CK(clk), .CE(n174), .R(n261), .D(n36), .Q(o_label5_data6[30]));
Q_FDP4EP \o_label5_data6_REG[31] ( .CK(clk), .CE(n174), .R(n261), .D(n37), .Q(o_label5_data6[31]));
Q_FDP4EP \o_label5_data7_REG[0] ( .CK(clk), .CE(n173), .R(n261), .D(n6), .Q(o_label5_data7[0]));
Q_FDP4EP \o_label5_data7_REG[1] ( .CK(clk), .CE(n173), .R(n261), .D(n7), .Q(o_label5_data7[1]));
Q_FDP4EP \o_label5_data7_REG[2] ( .CK(clk), .CE(n173), .R(n261), .D(n8), .Q(o_label5_data7[2]));
Q_FDP4EP \o_label5_data7_REG[3] ( .CK(clk), .CE(n173), .R(n261), .D(n9), .Q(o_label5_data7[3]));
Q_FDP4EP \o_label5_data7_REG[4] ( .CK(clk), .CE(n173), .R(n261), .D(n10), .Q(o_label5_data7[4]));
Q_FDP4EP \o_label5_data7_REG[5] ( .CK(clk), .CE(n173), .R(n261), .D(n11), .Q(o_label5_data7[5]));
Q_FDP4EP \o_label5_data7_REG[6] ( .CK(clk), .CE(n173), .R(n261), .D(n12), .Q(o_label5_data7[6]));
Q_FDP4EP \o_label5_data7_REG[7] ( .CK(clk), .CE(n173), .R(n261), .D(n13), .Q(o_label5_data7[7]));
Q_FDP4EP \o_label5_data7_REG[8] ( .CK(clk), .CE(n173), .R(n261), .D(n14), .Q(o_label5_data7[8]));
Q_FDP4EP \o_label5_data7_REG[9] ( .CK(clk), .CE(n173), .R(n261), .D(n15), .Q(o_label5_data7[9]));
Q_FDP4EP \o_label5_data7_REG[10] ( .CK(clk), .CE(n173), .R(n261), .D(n16), .Q(o_label5_data7[10]));
Q_FDP4EP \o_label5_data7_REG[11] ( .CK(clk), .CE(n173), .R(n261), .D(n17), .Q(o_label5_data7[11]));
Q_FDP4EP \o_label5_data7_REG[12] ( .CK(clk), .CE(n173), .R(n261), .D(n18), .Q(o_label5_data7[12]));
Q_FDP4EP \o_label5_data7_REG[13] ( .CK(clk), .CE(n173), .R(n261), .D(n19), .Q(o_label5_data7[13]));
Q_FDP4EP \o_label5_data7_REG[14] ( .CK(clk), .CE(n173), .R(n261), .D(n20), .Q(o_label5_data7[14]));
Q_FDP4EP \o_label5_data7_REG[15] ( .CK(clk), .CE(n173), .R(n261), .D(n21), .Q(o_label5_data7[15]));
Q_FDP4EP \o_label5_data7_REG[16] ( .CK(clk), .CE(n173), .R(n261), .D(n22), .Q(o_label5_data7[16]));
Q_FDP4EP \o_label5_data7_REG[17] ( .CK(clk), .CE(n173), .R(n261), .D(n23), .Q(o_label5_data7[17]));
Q_FDP4EP \o_label5_data7_REG[18] ( .CK(clk), .CE(n173), .R(n261), .D(n24), .Q(o_label5_data7[18]));
Q_FDP4EP \o_label5_data7_REG[19] ( .CK(clk), .CE(n173), .R(n261), .D(n25), .Q(o_label5_data7[19]));
Q_FDP4EP \o_label5_data7_REG[20] ( .CK(clk), .CE(n173), .R(n261), .D(n26), .Q(o_label5_data7[20]));
Q_FDP4EP \o_label5_data7_REG[21] ( .CK(clk), .CE(n173), .R(n261), .D(n27), .Q(o_label5_data7[21]));
Q_FDP4EP \o_label5_data7_REG[22] ( .CK(clk), .CE(n173), .R(n261), .D(n28), .Q(o_label5_data7[22]));
Q_FDP4EP \o_label5_data7_REG[23] ( .CK(clk), .CE(n173), .R(n261), .D(n29), .Q(o_label5_data7[23]));
Q_FDP4EP \o_label5_data7_REG[24] ( .CK(clk), .CE(n173), .R(n261), .D(n30), .Q(o_label5_data7[24]));
Q_FDP4EP \o_label5_data7_REG[25] ( .CK(clk), .CE(n173), .R(n261), .D(n31), .Q(o_label5_data7[25]));
Q_FDP4EP \o_label5_data7_REG[26] ( .CK(clk), .CE(n173), .R(n261), .D(n32), .Q(o_label5_data7[26]));
Q_FDP4EP \o_label5_data7_REG[27] ( .CK(clk), .CE(n173), .R(n261), .D(n33), .Q(o_label5_data7[27]));
Q_FDP4EP \o_label5_data7_REG[28] ( .CK(clk), .CE(n173), .R(n261), .D(n34), .Q(o_label5_data7[28]));
Q_FDP4EP \o_label5_data7_REG[29] ( .CK(clk), .CE(n173), .R(n261), .D(n35), .Q(o_label5_data7[29]));
Q_FDP4EP \o_label5_data7_REG[30] ( .CK(clk), .CE(n173), .R(n261), .D(n36), .Q(o_label5_data7[30]));
Q_FDP4EP \o_label5_data7_REG[31] ( .CK(clk), .CE(n173), .R(n261), .D(n37), .Q(o_label5_data7[31]));
Q_FDP4EP \o_label5_config_REG[0] ( .CK(clk), .CE(n172), .R(n261), .D(n6), .Q(o_label5_config[0]));
Q_FDP4EP \o_label5_config_REG[1] ( .CK(clk), .CE(n172), .R(n261), .D(n7), .Q(o_label5_config[1]));
Q_FDP4EP \o_label5_config_REG[2] ( .CK(clk), .CE(n172), .R(n261), .D(n8), .Q(o_label5_config[2]));
Q_FDP4EP \o_label5_config_REG[3] ( .CK(clk), .CE(n172), .R(n261), .D(n9), .Q(o_label5_config[3]));
Q_FDP4EP \o_label5_config_REG[4] ( .CK(clk), .CE(n172), .R(n261), .D(n10), .Q(o_label5_config[4]));
Q_FDP4EP \o_label5_config_REG[5] ( .CK(clk), .CE(n172), .R(n261), .D(n11), .Q(o_label5_config[5]));
Q_FDP4EP \o_label5_config_REG[6] ( .CK(clk), .CE(n172), .R(n261), .D(n12), .Q(o_label5_config[6]));
Q_FDP4EP \o_label5_config_REG[7] ( .CK(clk), .CE(n172), .R(n261), .D(n13), .Q(o_label5_config[7]));
Q_FDP4EP \o_label5_config_REG[9] ( .CK(clk), .CE(n172), .R(n261), .D(n31), .Q(o_label5_config[9]));
Q_FDP4EP \o_label5_config_REG[10] ( .CK(clk), .CE(n172), .R(n261), .D(n32), .Q(o_label5_config[10]));
Q_FDP4EP \o_label5_config_REG[11] ( .CK(clk), .CE(n172), .R(n261), .D(n33), .Q(o_label5_config[11]));
Q_FDP4EP \o_label5_config_REG[12] ( .CK(clk), .CE(n172), .R(n261), .D(n34), .Q(o_label5_config[12]));
Q_FDP4EP \o_label5_config_REG[13] ( .CK(clk), .CE(n172), .R(n261), .D(n35), .Q(o_label5_config[13]));
Q_FDP4EP \o_label5_config_REG[14] ( .CK(clk), .CE(n172), .R(n261), .D(n36), .Q(o_label5_config[14]));
Q_FDP4EP \o_label5_config_REG[15] ( .CK(clk), .CE(n172), .R(n261), .D(n37), .Q(o_label5_config[15]));
Q_FDP4EP \o_label4_data0_REG[0] ( .CK(clk), .CE(n171), .R(n261), .D(n6), .Q(o_label4_data0[0]));
Q_FDP4EP \o_label4_data0_REG[1] ( .CK(clk), .CE(n171), .R(n261), .D(n7), .Q(o_label4_data0[1]));
Q_FDP4EP \o_label4_data0_REG[2] ( .CK(clk), .CE(n171), .R(n261), .D(n8), .Q(o_label4_data0[2]));
Q_FDP4EP \o_label4_data0_REG[3] ( .CK(clk), .CE(n171), .R(n261), .D(n9), .Q(o_label4_data0[3]));
Q_FDP4EP \o_label4_data0_REG[4] ( .CK(clk), .CE(n171), .R(n261), .D(n10), .Q(o_label4_data0[4]));
Q_FDP4EP \o_label4_data0_REG[5] ( .CK(clk), .CE(n171), .R(n261), .D(n11), .Q(o_label4_data0[5]));
Q_FDP4EP \o_label4_data0_REG[6] ( .CK(clk), .CE(n171), .R(n261), .D(n12), .Q(o_label4_data0[6]));
Q_FDP4EP \o_label4_data0_REG[7] ( .CK(clk), .CE(n171), .R(n261), .D(n13), .Q(o_label4_data0[7]));
Q_FDP4EP \o_label4_data0_REG[8] ( .CK(clk), .CE(n171), .R(n261), .D(n14), .Q(o_label4_data0[8]));
Q_FDP4EP \o_label4_data0_REG[9] ( .CK(clk), .CE(n171), .R(n261), .D(n15), .Q(o_label4_data0[9]));
Q_FDP4EP \o_label4_data0_REG[10] ( .CK(clk), .CE(n171), .R(n261), .D(n16), .Q(o_label4_data0[10]));
Q_FDP4EP \o_label4_data0_REG[11] ( .CK(clk), .CE(n171), .R(n261), .D(n17), .Q(o_label4_data0[11]));
Q_FDP4EP \o_label4_data0_REG[12] ( .CK(clk), .CE(n171), .R(n261), .D(n18), .Q(o_label4_data0[12]));
Q_FDP4EP \o_label4_data0_REG[13] ( .CK(clk), .CE(n171), .R(n261), .D(n19), .Q(o_label4_data0[13]));
Q_FDP4EP \o_label4_data0_REG[14] ( .CK(clk), .CE(n171), .R(n261), .D(n20), .Q(o_label4_data0[14]));
Q_FDP4EP \o_label4_data0_REG[15] ( .CK(clk), .CE(n171), .R(n261), .D(n21), .Q(o_label4_data0[15]));
Q_FDP4EP \o_label4_data0_REG[16] ( .CK(clk), .CE(n171), .R(n261), .D(n22), .Q(o_label4_data0[16]));
Q_FDP4EP \o_label4_data0_REG[17] ( .CK(clk), .CE(n171), .R(n261), .D(n23), .Q(o_label4_data0[17]));
Q_FDP4EP \o_label4_data0_REG[18] ( .CK(clk), .CE(n171), .R(n261), .D(n24), .Q(o_label4_data0[18]));
Q_FDP4EP \o_label4_data0_REG[19] ( .CK(clk), .CE(n171), .R(n261), .D(n25), .Q(o_label4_data0[19]));
Q_FDP4EP \o_label4_data0_REG[20] ( .CK(clk), .CE(n171), .R(n261), .D(n26), .Q(o_label4_data0[20]));
Q_FDP4EP \o_label4_data0_REG[21] ( .CK(clk), .CE(n171), .R(n261), .D(n27), .Q(o_label4_data0[21]));
Q_FDP4EP \o_label4_data0_REG[22] ( .CK(clk), .CE(n171), .R(n261), .D(n28), .Q(o_label4_data0[22]));
Q_FDP4EP \o_label4_data0_REG[23] ( .CK(clk), .CE(n171), .R(n261), .D(n29), .Q(o_label4_data0[23]));
Q_FDP4EP \o_label4_data0_REG[24] ( .CK(clk), .CE(n171), .R(n261), .D(n30), .Q(o_label4_data0[24]));
Q_FDP4EP \o_label4_data0_REG[25] ( .CK(clk), .CE(n171), .R(n261), .D(n31), .Q(o_label4_data0[25]));
Q_FDP4EP \o_label4_data0_REG[26] ( .CK(clk), .CE(n171), .R(n261), .D(n32), .Q(o_label4_data0[26]));
Q_FDP4EP \o_label4_data0_REG[27] ( .CK(clk), .CE(n171), .R(n261), .D(n33), .Q(o_label4_data0[27]));
Q_FDP4EP \o_label4_data0_REG[28] ( .CK(clk), .CE(n171), .R(n261), .D(n34), .Q(o_label4_data0[28]));
Q_FDP4EP \o_label4_data0_REG[29] ( .CK(clk), .CE(n171), .R(n261), .D(n35), .Q(o_label4_data0[29]));
Q_FDP4EP \o_label4_data0_REG[30] ( .CK(clk), .CE(n171), .R(n261), .D(n36), .Q(o_label4_data0[30]));
Q_FDP4EP \o_label4_data0_REG[31] ( .CK(clk), .CE(n171), .R(n261), .D(n37), .Q(o_label4_data0[31]));
Q_FDP4EP \o_label4_data1_REG[0] ( .CK(clk), .CE(n170), .R(n261), .D(n6), .Q(o_label4_data1[0]));
Q_FDP4EP \o_label4_data1_REG[1] ( .CK(clk), .CE(n170), .R(n261), .D(n7), .Q(o_label4_data1[1]));
Q_FDP4EP \o_label4_data1_REG[2] ( .CK(clk), .CE(n170), .R(n261), .D(n8), .Q(o_label4_data1[2]));
Q_FDP4EP \o_label4_data1_REG[3] ( .CK(clk), .CE(n170), .R(n261), .D(n9), .Q(o_label4_data1[3]));
Q_FDP4EP \o_label4_data1_REG[4] ( .CK(clk), .CE(n170), .R(n261), .D(n10), .Q(o_label4_data1[4]));
Q_FDP4EP \o_label4_data1_REG[5] ( .CK(clk), .CE(n170), .R(n261), .D(n11), .Q(o_label4_data1[5]));
Q_FDP4EP \o_label4_data1_REG[6] ( .CK(clk), .CE(n170), .R(n261), .D(n12), .Q(o_label4_data1[6]));
Q_FDP4EP \o_label4_data1_REG[7] ( .CK(clk), .CE(n170), .R(n261), .D(n13), .Q(o_label4_data1[7]));
Q_FDP4EP \o_label4_data1_REG[8] ( .CK(clk), .CE(n170), .R(n261), .D(n14), .Q(o_label4_data1[8]));
Q_FDP4EP \o_label4_data1_REG[9] ( .CK(clk), .CE(n170), .R(n261), .D(n15), .Q(o_label4_data1[9]));
Q_FDP4EP \o_label4_data1_REG[10] ( .CK(clk), .CE(n170), .R(n261), .D(n16), .Q(o_label4_data1[10]));
Q_FDP4EP \o_label4_data1_REG[11] ( .CK(clk), .CE(n170), .R(n261), .D(n17), .Q(o_label4_data1[11]));
Q_FDP4EP \o_label4_data1_REG[12] ( .CK(clk), .CE(n170), .R(n261), .D(n18), .Q(o_label4_data1[12]));
Q_FDP4EP \o_label4_data1_REG[13] ( .CK(clk), .CE(n170), .R(n261), .D(n19), .Q(o_label4_data1[13]));
Q_FDP4EP \o_label4_data1_REG[14] ( .CK(clk), .CE(n170), .R(n261), .D(n20), .Q(o_label4_data1[14]));
Q_FDP4EP \o_label4_data1_REG[15] ( .CK(clk), .CE(n170), .R(n261), .D(n21), .Q(o_label4_data1[15]));
Q_FDP4EP \o_label4_data1_REG[16] ( .CK(clk), .CE(n170), .R(n261), .D(n22), .Q(o_label4_data1[16]));
Q_FDP4EP \o_label4_data1_REG[17] ( .CK(clk), .CE(n170), .R(n261), .D(n23), .Q(o_label4_data1[17]));
Q_FDP4EP \o_label4_data1_REG[18] ( .CK(clk), .CE(n170), .R(n261), .D(n24), .Q(o_label4_data1[18]));
Q_FDP4EP \o_label4_data1_REG[19] ( .CK(clk), .CE(n170), .R(n261), .D(n25), .Q(o_label4_data1[19]));
Q_FDP4EP \o_label4_data1_REG[20] ( .CK(clk), .CE(n170), .R(n261), .D(n26), .Q(o_label4_data1[20]));
Q_FDP4EP \o_label4_data1_REG[21] ( .CK(clk), .CE(n170), .R(n261), .D(n27), .Q(o_label4_data1[21]));
Q_FDP4EP \o_label4_data1_REG[22] ( .CK(clk), .CE(n170), .R(n261), .D(n28), .Q(o_label4_data1[22]));
Q_FDP4EP \o_label4_data1_REG[23] ( .CK(clk), .CE(n170), .R(n261), .D(n29), .Q(o_label4_data1[23]));
Q_FDP4EP \o_label4_data1_REG[24] ( .CK(clk), .CE(n170), .R(n261), .D(n30), .Q(o_label4_data1[24]));
Q_FDP4EP \o_label4_data1_REG[25] ( .CK(clk), .CE(n170), .R(n261), .D(n31), .Q(o_label4_data1[25]));
Q_FDP4EP \o_label4_data1_REG[26] ( .CK(clk), .CE(n170), .R(n261), .D(n32), .Q(o_label4_data1[26]));
Q_FDP4EP \o_label4_data1_REG[27] ( .CK(clk), .CE(n170), .R(n261), .D(n33), .Q(o_label4_data1[27]));
Q_FDP4EP \o_label4_data1_REG[28] ( .CK(clk), .CE(n170), .R(n261), .D(n34), .Q(o_label4_data1[28]));
Q_FDP4EP \o_label4_data1_REG[29] ( .CK(clk), .CE(n170), .R(n261), .D(n35), .Q(o_label4_data1[29]));
Q_FDP4EP \o_label4_data1_REG[30] ( .CK(clk), .CE(n170), .R(n261), .D(n36), .Q(o_label4_data1[30]));
Q_FDP4EP \o_label4_data1_REG[31] ( .CK(clk), .CE(n170), .R(n261), .D(n37), .Q(o_label4_data1[31]));
Q_FDP4EP \o_label4_data2_REG[0] ( .CK(clk), .CE(n169), .R(n261), .D(n6), .Q(o_label4_data2[0]));
Q_FDP4EP \o_label4_data2_REG[1] ( .CK(clk), .CE(n169), .R(n261), .D(n7), .Q(o_label4_data2[1]));
Q_FDP4EP \o_label4_data2_REG[2] ( .CK(clk), .CE(n169), .R(n261), .D(n8), .Q(o_label4_data2[2]));
Q_FDP4EP \o_label4_data2_REG[3] ( .CK(clk), .CE(n169), .R(n261), .D(n9), .Q(o_label4_data2[3]));
Q_FDP4EP \o_label4_data2_REG[4] ( .CK(clk), .CE(n169), .R(n261), .D(n10), .Q(o_label4_data2[4]));
Q_FDP4EP \o_label4_data2_REG[5] ( .CK(clk), .CE(n169), .R(n261), .D(n11), .Q(o_label4_data2[5]));
Q_FDP4EP \o_label4_data2_REG[6] ( .CK(clk), .CE(n169), .R(n261), .D(n12), .Q(o_label4_data2[6]));
Q_FDP4EP \o_label4_data2_REG[7] ( .CK(clk), .CE(n169), .R(n261), .D(n13), .Q(o_label4_data2[7]));
Q_FDP4EP \o_label4_data2_REG[8] ( .CK(clk), .CE(n169), .R(n261), .D(n14), .Q(o_label4_data2[8]));
Q_FDP4EP \o_label4_data2_REG[9] ( .CK(clk), .CE(n169), .R(n261), .D(n15), .Q(o_label4_data2[9]));
Q_FDP4EP \o_label4_data2_REG[10] ( .CK(clk), .CE(n169), .R(n261), .D(n16), .Q(o_label4_data2[10]));
Q_FDP4EP \o_label4_data2_REG[11] ( .CK(clk), .CE(n169), .R(n261), .D(n17), .Q(o_label4_data2[11]));
Q_FDP4EP \o_label4_data2_REG[12] ( .CK(clk), .CE(n169), .R(n261), .D(n18), .Q(o_label4_data2[12]));
Q_FDP4EP \o_label4_data2_REG[13] ( .CK(clk), .CE(n169), .R(n261), .D(n19), .Q(o_label4_data2[13]));
Q_FDP4EP \o_label4_data2_REG[14] ( .CK(clk), .CE(n169), .R(n261), .D(n20), .Q(o_label4_data2[14]));
Q_FDP4EP \o_label4_data2_REG[15] ( .CK(clk), .CE(n169), .R(n261), .D(n21), .Q(o_label4_data2[15]));
Q_FDP4EP \o_label4_data2_REG[16] ( .CK(clk), .CE(n169), .R(n261), .D(n22), .Q(o_label4_data2[16]));
Q_FDP4EP \o_label4_data2_REG[17] ( .CK(clk), .CE(n169), .R(n261), .D(n23), .Q(o_label4_data2[17]));
Q_FDP4EP \o_label4_data2_REG[18] ( .CK(clk), .CE(n169), .R(n261), .D(n24), .Q(o_label4_data2[18]));
Q_FDP4EP \o_label4_data2_REG[19] ( .CK(clk), .CE(n169), .R(n261), .D(n25), .Q(o_label4_data2[19]));
Q_FDP4EP \o_label4_data2_REG[20] ( .CK(clk), .CE(n169), .R(n261), .D(n26), .Q(o_label4_data2[20]));
Q_FDP4EP \o_label4_data2_REG[21] ( .CK(clk), .CE(n169), .R(n261), .D(n27), .Q(o_label4_data2[21]));
Q_FDP4EP \o_label4_data2_REG[22] ( .CK(clk), .CE(n169), .R(n261), .D(n28), .Q(o_label4_data2[22]));
Q_FDP4EP \o_label4_data2_REG[23] ( .CK(clk), .CE(n169), .R(n261), .D(n29), .Q(o_label4_data2[23]));
Q_FDP4EP \o_label4_data2_REG[24] ( .CK(clk), .CE(n169), .R(n261), .D(n30), .Q(o_label4_data2[24]));
Q_FDP4EP \o_label4_data2_REG[25] ( .CK(clk), .CE(n169), .R(n261), .D(n31), .Q(o_label4_data2[25]));
Q_FDP4EP \o_label4_data2_REG[26] ( .CK(clk), .CE(n169), .R(n261), .D(n32), .Q(o_label4_data2[26]));
Q_FDP4EP \o_label4_data2_REG[27] ( .CK(clk), .CE(n169), .R(n261), .D(n33), .Q(o_label4_data2[27]));
Q_FDP4EP \o_label4_data2_REG[28] ( .CK(clk), .CE(n169), .R(n261), .D(n34), .Q(o_label4_data2[28]));
Q_FDP4EP \o_label4_data2_REG[29] ( .CK(clk), .CE(n169), .R(n261), .D(n35), .Q(o_label4_data2[29]));
Q_FDP4EP \o_label4_data2_REG[30] ( .CK(clk), .CE(n169), .R(n261), .D(n36), .Q(o_label4_data2[30]));
Q_FDP4EP \o_label4_data2_REG[31] ( .CK(clk), .CE(n169), .R(n261), .D(n37), .Q(o_label4_data2[31]));
Q_FDP4EP \o_label4_data3_REG[0] ( .CK(clk), .CE(n168), .R(n261), .D(n6), .Q(o_label4_data3[0]));
Q_FDP4EP \o_label4_data3_REG[1] ( .CK(clk), .CE(n168), .R(n261), .D(n7), .Q(o_label4_data3[1]));
Q_FDP4EP \o_label4_data3_REG[2] ( .CK(clk), .CE(n168), .R(n261), .D(n8), .Q(o_label4_data3[2]));
Q_FDP4EP \o_label4_data3_REG[3] ( .CK(clk), .CE(n168), .R(n261), .D(n9), .Q(o_label4_data3[3]));
Q_FDP4EP \o_label4_data3_REG[4] ( .CK(clk), .CE(n168), .R(n261), .D(n10), .Q(o_label4_data3[4]));
Q_FDP4EP \o_label4_data3_REG[5] ( .CK(clk), .CE(n168), .R(n261), .D(n11), .Q(o_label4_data3[5]));
Q_FDP4EP \o_label4_data3_REG[6] ( .CK(clk), .CE(n168), .R(n261), .D(n12), .Q(o_label4_data3[6]));
Q_FDP4EP \o_label4_data3_REG[7] ( .CK(clk), .CE(n168), .R(n261), .D(n13), .Q(o_label4_data3[7]));
Q_FDP4EP \o_label4_data3_REG[8] ( .CK(clk), .CE(n168), .R(n261), .D(n14), .Q(o_label4_data3[8]));
Q_FDP4EP \o_label4_data3_REG[9] ( .CK(clk), .CE(n168), .R(n261), .D(n15), .Q(o_label4_data3[9]));
Q_FDP4EP \o_label4_data3_REG[10] ( .CK(clk), .CE(n168), .R(n261), .D(n16), .Q(o_label4_data3[10]));
Q_FDP4EP \o_label4_data3_REG[11] ( .CK(clk), .CE(n168), .R(n261), .D(n17), .Q(o_label4_data3[11]));
Q_FDP4EP \o_label4_data3_REG[12] ( .CK(clk), .CE(n168), .R(n261), .D(n18), .Q(o_label4_data3[12]));
Q_FDP4EP \o_label4_data3_REG[13] ( .CK(clk), .CE(n168), .R(n261), .D(n19), .Q(o_label4_data3[13]));
Q_FDP4EP \o_label4_data3_REG[14] ( .CK(clk), .CE(n168), .R(n261), .D(n20), .Q(o_label4_data3[14]));
Q_FDP4EP \o_label4_data3_REG[15] ( .CK(clk), .CE(n168), .R(n261), .D(n21), .Q(o_label4_data3[15]));
Q_FDP4EP \o_label4_data3_REG[16] ( .CK(clk), .CE(n168), .R(n261), .D(n22), .Q(o_label4_data3[16]));
Q_FDP4EP \o_label4_data3_REG[17] ( .CK(clk), .CE(n168), .R(n261), .D(n23), .Q(o_label4_data3[17]));
Q_FDP4EP \o_label4_data3_REG[18] ( .CK(clk), .CE(n168), .R(n261), .D(n24), .Q(o_label4_data3[18]));
Q_FDP4EP \o_label4_data3_REG[19] ( .CK(clk), .CE(n168), .R(n261), .D(n25), .Q(o_label4_data3[19]));
Q_FDP4EP \o_label4_data3_REG[20] ( .CK(clk), .CE(n168), .R(n261), .D(n26), .Q(o_label4_data3[20]));
Q_FDP4EP \o_label4_data3_REG[21] ( .CK(clk), .CE(n168), .R(n261), .D(n27), .Q(o_label4_data3[21]));
Q_FDP4EP \o_label4_data3_REG[22] ( .CK(clk), .CE(n168), .R(n261), .D(n28), .Q(o_label4_data3[22]));
Q_FDP4EP \o_label4_data3_REG[23] ( .CK(clk), .CE(n168), .R(n261), .D(n29), .Q(o_label4_data3[23]));
Q_FDP4EP \o_label4_data3_REG[24] ( .CK(clk), .CE(n168), .R(n261), .D(n30), .Q(o_label4_data3[24]));
Q_FDP4EP \o_label4_data3_REG[25] ( .CK(clk), .CE(n168), .R(n261), .D(n31), .Q(o_label4_data3[25]));
Q_FDP4EP \o_label4_data3_REG[26] ( .CK(clk), .CE(n168), .R(n261), .D(n32), .Q(o_label4_data3[26]));
Q_FDP4EP \o_label4_data3_REG[27] ( .CK(clk), .CE(n168), .R(n261), .D(n33), .Q(o_label4_data3[27]));
Q_FDP4EP \o_label4_data3_REG[28] ( .CK(clk), .CE(n168), .R(n261), .D(n34), .Q(o_label4_data3[28]));
Q_FDP4EP \o_label4_data3_REG[29] ( .CK(clk), .CE(n168), .R(n261), .D(n35), .Q(o_label4_data3[29]));
Q_FDP4EP \o_label4_data3_REG[30] ( .CK(clk), .CE(n168), .R(n261), .D(n36), .Q(o_label4_data3[30]));
Q_FDP4EP \o_label4_data3_REG[31] ( .CK(clk), .CE(n168), .R(n261), .D(n37), .Q(o_label4_data3[31]));
Q_FDP4EP \o_label4_data4_REG[0] ( .CK(clk), .CE(n167), .R(n261), .D(n6), .Q(o_label4_data4[0]));
Q_FDP4EP \o_label4_data4_REG[1] ( .CK(clk), .CE(n167), .R(n261), .D(n7), .Q(o_label4_data4[1]));
Q_FDP4EP \o_label4_data4_REG[2] ( .CK(clk), .CE(n167), .R(n261), .D(n8), .Q(o_label4_data4[2]));
Q_FDP4EP \o_label4_data4_REG[3] ( .CK(clk), .CE(n167), .R(n261), .D(n9), .Q(o_label4_data4[3]));
Q_FDP4EP \o_label4_data4_REG[4] ( .CK(clk), .CE(n167), .R(n261), .D(n10), .Q(o_label4_data4[4]));
Q_FDP4EP \o_label4_data4_REG[5] ( .CK(clk), .CE(n167), .R(n261), .D(n11), .Q(o_label4_data4[5]));
Q_FDP4EP \o_label4_data4_REG[6] ( .CK(clk), .CE(n167), .R(n261), .D(n12), .Q(o_label4_data4[6]));
Q_FDP4EP \o_label4_data4_REG[7] ( .CK(clk), .CE(n167), .R(n261), .D(n13), .Q(o_label4_data4[7]));
Q_FDP4EP \o_label4_data4_REG[8] ( .CK(clk), .CE(n167), .R(n261), .D(n14), .Q(o_label4_data4[8]));
Q_FDP4EP \o_label4_data4_REG[9] ( .CK(clk), .CE(n167), .R(n261), .D(n15), .Q(o_label4_data4[9]));
Q_FDP4EP \o_label4_data4_REG[10] ( .CK(clk), .CE(n167), .R(n261), .D(n16), .Q(o_label4_data4[10]));
Q_FDP4EP \o_label4_data4_REG[11] ( .CK(clk), .CE(n167), .R(n261), .D(n17), .Q(o_label4_data4[11]));
Q_FDP4EP \o_label4_data4_REG[12] ( .CK(clk), .CE(n167), .R(n261), .D(n18), .Q(o_label4_data4[12]));
Q_FDP4EP \o_label4_data4_REG[13] ( .CK(clk), .CE(n167), .R(n261), .D(n19), .Q(o_label4_data4[13]));
Q_FDP4EP \o_label4_data4_REG[14] ( .CK(clk), .CE(n167), .R(n261), .D(n20), .Q(o_label4_data4[14]));
Q_FDP4EP \o_label4_data4_REG[15] ( .CK(clk), .CE(n167), .R(n261), .D(n21), .Q(o_label4_data4[15]));
Q_FDP4EP \o_label4_data4_REG[16] ( .CK(clk), .CE(n167), .R(n261), .D(n22), .Q(o_label4_data4[16]));
Q_FDP4EP \o_label4_data4_REG[17] ( .CK(clk), .CE(n167), .R(n261), .D(n23), .Q(o_label4_data4[17]));
Q_FDP4EP \o_label4_data4_REG[18] ( .CK(clk), .CE(n167), .R(n261), .D(n24), .Q(o_label4_data4[18]));
Q_FDP4EP \o_label4_data4_REG[19] ( .CK(clk), .CE(n167), .R(n261), .D(n25), .Q(o_label4_data4[19]));
Q_FDP4EP \o_label4_data4_REG[20] ( .CK(clk), .CE(n167), .R(n261), .D(n26), .Q(o_label4_data4[20]));
Q_FDP4EP \o_label4_data4_REG[21] ( .CK(clk), .CE(n167), .R(n261), .D(n27), .Q(o_label4_data4[21]));
Q_FDP4EP \o_label4_data4_REG[22] ( .CK(clk), .CE(n167), .R(n261), .D(n28), .Q(o_label4_data4[22]));
Q_FDP4EP \o_label4_data4_REG[23] ( .CK(clk), .CE(n167), .R(n261), .D(n29), .Q(o_label4_data4[23]));
Q_FDP4EP \o_label4_data4_REG[24] ( .CK(clk), .CE(n167), .R(n261), .D(n30), .Q(o_label4_data4[24]));
Q_FDP4EP \o_label4_data4_REG[25] ( .CK(clk), .CE(n167), .R(n261), .D(n31), .Q(o_label4_data4[25]));
Q_FDP4EP \o_label4_data4_REG[26] ( .CK(clk), .CE(n167), .R(n261), .D(n32), .Q(o_label4_data4[26]));
Q_FDP4EP \o_label4_data4_REG[27] ( .CK(clk), .CE(n167), .R(n261), .D(n33), .Q(o_label4_data4[27]));
Q_FDP4EP \o_label4_data4_REG[28] ( .CK(clk), .CE(n167), .R(n261), .D(n34), .Q(o_label4_data4[28]));
Q_FDP4EP \o_label4_data4_REG[29] ( .CK(clk), .CE(n167), .R(n261), .D(n35), .Q(o_label4_data4[29]));
Q_FDP4EP \o_label4_data4_REG[30] ( .CK(clk), .CE(n167), .R(n261), .D(n36), .Q(o_label4_data4[30]));
Q_FDP4EP \o_label4_data4_REG[31] ( .CK(clk), .CE(n167), .R(n261), .D(n37), .Q(o_label4_data4[31]));
Q_FDP4EP \o_label4_data5_REG[0] ( .CK(clk), .CE(n166), .R(n261), .D(n6), .Q(o_label4_data5[0]));
Q_FDP4EP \o_label4_data5_REG[1] ( .CK(clk), .CE(n166), .R(n261), .D(n7), .Q(o_label4_data5[1]));
Q_FDP4EP \o_label4_data5_REG[2] ( .CK(clk), .CE(n166), .R(n261), .D(n8), .Q(o_label4_data5[2]));
Q_FDP4EP \o_label4_data5_REG[3] ( .CK(clk), .CE(n166), .R(n261), .D(n9), .Q(o_label4_data5[3]));
Q_FDP4EP \o_label4_data5_REG[4] ( .CK(clk), .CE(n166), .R(n261), .D(n10), .Q(o_label4_data5[4]));
Q_FDP4EP \o_label4_data5_REG[5] ( .CK(clk), .CE(n166), .R(n261), .D(n11), .Q(o_label4_data5[5]));
Q_FDP4EP \o_label4_data5_REG[6] ( .CK(clk), .CE(n166), .R(n261), .D(n12), .Q(o_label4_data5[6]));
Q_FDP4EP \o_label4_data5_REG[7] ( .CK(clk), .CE(n166), .R(n261), .D(n13), .Q(o_label4_data5[7]));
Q_FDP4EP \o_label4_data5_REG[8] ( .CK(clk), .CE(n166), .R(n261), .D(n14), .Q(o_label4_data5[8]));
Q_FDP4EP \o_label4_data5_REG[9] ( .CK(clk), .CE(n166), .R(n261), .D(n15), .Q(o_label4_data5[9]));
Q_FDP4EP \o_label4_data5_REG[10] ( .CK(clk), .CE(n166), .R(n261), .D(n16), .Q(o_label4_data5[10]));
Q_FDP4EP \o_label4_data5_REG[11] ( .CK(clk), .CE(n166), .R(n261), .D(n17), .Q(o_label4_data5[11]));
Q_FDP4EP \o_label4_data5_REG[12] ( .CK(clk), .CE(n166), .R(n261), .D(n18), .Q(o_label4_data5[12]));
Q_FDP4EP \o_label4_data5_REG[13] ( .CK(clk), .CE(n166), .R(n261), .D(n19), .Q(o_label4_data5[13]));
Q_FDP4EP \o_label4_data5_REG[14] ( .CK(clk), .CE(n166), .R(n261), .D(n20), .Q(o_label4_data5[14]));
Q_FDP4EP \o_label4_data5_REG[15] ( .CK(clk), .CE(n166), .R(n261), .D(n21), .Q(o_label4_data5[15]));
Q_FDP4EP \o_label4_data5_REG[16] ( .CK(clk), .CE(n166), .R(n261), .D(n22), .Q(o_label4_data5[16]));
Q_FDP4EP \o_label4_data5_REG[17] ( .CK(clk), .CE(n166), .R(n261), .D(n23), .Q(o_label4_data5[17]));
Q_FDP4EP \o_label4_data5_REG[18] ( .CK(clk), .CE(n166), .R(n261), .D(n24), .Q(o_label4_data5[18]));
Q_FDP4EP \o_label4_data5_REG[19] ( .CK(clk), .CE(n166), .R(n261), .D(n25), .Q(o_label4_data5[19]));
Q_FDP4EP \o_label4_data5_REG[20] ( .CK(clk), .CE(n166), .R(n261), .D(n26), .Q(o_label4_data5[20]));
Q_FDP4EP \o_label4_data5_REG[21] ( .CK(clk), .CE(n166), .R(n261), .D(n27), .Q(o_label4_data5[21]));
Q_FDP4EP \o_label4_data5_REG[22] ( .CK(clk), .CE(n166), .R(n261), .D(n28), .Q(o_label4_data5[22]));
Q_FDP4EP \o_label4_data5_REG[23] ( .CK(clk), .CE(n166), .R(n261), .D(n29), .Q(o_label4_data5[23]));
Q_FDP4EP \o_label4_data5_REG[24] ( .CK(clk), .CE(n166), .R(n261), .D(n30), .Q(o_label4_data5[24]));
Q_FDP4EP \o_label4_data5_REG[25] ( .CK(clk), .CE(n166), .R(n261), .D(n31), .Q(o_label4_data5[25]));
Q_FDP4EP \o_label4_data5_REG[26] ( .CK(clk), .CE(n166), .R(n261), .D(n32), .Q(o_label4_data5[26]));
Q_FDP4EP \o_label4_data5_REG[27] ( .CK(clk), .CE(n166), .R(n261), .D(n33), .Q(o_label4_data5[27]));
Q_FDP4EP \o_label4_data5_REG[28] ( .CK(clk), .CE(n166), .R(n261), .D(n34), .Q(o_label4_data5[28]));
Q_FDP4EP \o_label4_data5_REG[29] ( .CK(clk), .CE(n166), .R(n261), .D(n35), .Q(o_label4_data5[29]));
Q_FDP4EP \o_label4_data5_REG[30] ( .CK(clk), .CE(n166), .R(n261), .D(n36), .Q(o_label4_data5[30]));
Q_FDP4EP \o_label4_data5_REG[31] ( .CK(clk), .CE(n166), .R(n261), .D(n37), .Q(o_label4_data5[31]));
Q_FDP4EP \o_label4_data6_REG[0] ( .CK(clk), .CE(n165), .R(n261), .D(n6), .Q(o_label4_data6[0]));
Q_FDP4EP \o_label4_data6_REG[1] ( .CK(clk), .CE(n165), .R(n261), .D(n7), .Q(o_label4_data6[1]));
Q_FDP4EP \o_label4_data6_REG[2] ( .CK(clk), .CE(n165), .R(n261), .D(n8), .Q(o_label4_data6[2]));
Q_FDP4EP \o_label4_data6_REG[3] ( .CK(clk), .CE(n165), .R(n261), .D(n9), .Q(o_label4_data6[3]));
Q_FDP4EP \o_label4_data6_REG[4] ( .CK(clk), .CE(n165), .R(n261), .D(n10), .Q(o_label4_data6[4]));
Q_FDP4EP \o_label4_data6_REG[5] ( .CK(clk), .CE(n165), .R(n261), .D(n11), .Q(o_label4_data6[5]));
Q_FDP4EP \o_label4_data6_REG[6] ( .CK(clk), .CE(n165), .R(n261), .D(n12), .Q(o_label4_data6[6]));
Q_FDP4EP \o_label4_data6_REG[7] ( .CK(clk), .CE(n165), .R(n261), .D(n13), .Q(o_label4_data6[7]));
Q_FDP4EP \o_label4_data6_REG[8] ( .CK(clk), .CE(n165), .R(n261), .D(n14), .Q(o_label4_data6[8]));
Q_FDP4EP \o_label4_data6_REG[9] ( .CK(clk), .CE(n165), .R(n261), .D(n15), .Q(o_label4_data6[9]));
Q_FDP4EP \o_label4_data6_REG[10] ( .CK(clk), .CE(n165), .R(n261), .D(n16), .Q(o_label4_data6[10]));
Q_FDP4EP \o_label4_data6_REG[11] ( .CK(clk), .CE(n165), .R(n261), .D(n17), .Q(o_label4_data6[11]));
Q_FDP4EP \o_label4_data6_REG[12] ( .CK(clk), .CE(n165), .R(n261), .D(n18), .Q(o_label4_data6[12]));
Q_FDP4EP \o_label4_data6_REG[13] ( .CK(clk), .CE(n165), .R(n261), .D(n19), .Q(o_label4_data6[13]));
Q_FDP4EP \o_label4_data6_REG[14] ( .CK(clk), .CE(n165), .R(n261), .D(n20), .Q(o_label4_data6[14]));
Q_FDP4EP \o_label4_data6_REG[15] ( .CK(clk), .CE(n165), .R(n261), .D(n21), .Q(o_label4_data6[15]));
Q_FDP4EP \o_label4_data6_REG[16] ( .CK(clk), .CE(n165), .R(n261), .D(n22), .Q(o_label4_data6[16]));
Q_FDP4EP \o_label4_data6_REG[17] ( .CK(clk), .CE(n165), .R(n261), .D(n23), .Q(o_label4_data6[17]));
Q_FDP4EP \o_label4_data6_REG[18] ( .CK(clk), .CE(n165), .R(n261), .D(n24), .Q(o_label4_data6[18]));
Q_FDP4EP \o_label4_data6_REG[19] ( .CK(clk), .CE(n165), .R(n261), .D(n25), .Q(o_label4_data6[19]));
Q_FDP4EP \o_label4_data6_REG[20] ( .CK(clk), .CE(n165), .R(n261), .D(n26), .Q(o_label4_data6[20]));
Q_FDP4EP \o_label4_data6_REG[21] ( .CK(clk), .CE(n165), .R(n261), .D(n27), .Q(o_label4_data6[21]));
Q_FDP4EP \o_label4_data6_REG[22] ( .CK(clk), .CE(n165), .R(n261), .D(n28), .Q(o_label4_data6[22]));
Q_FDP4EP \o_label4_data6_REG[23] ( .CK(clk), .CE(n165), .R(n261), .D(n29), .Q(o_label4_data6[23]));
Q_FDP4EP \o_label4_data6_REG[24] ( .CK(clk), .CE(n165), .R(n261), .D(n30), .Q(o_label4_data6[24]));
Q_FDP4EP \o_label4_data6_REG[25] ( .CK(clk), .CE(n165), .R(n261), .D(n31), .Q(o_label4_data6[25]));
Q_FDP4EP \o_label4_data6_REG[26] ( .CK(clk), .CE(n165), .R(n261), .D(n32), .Q(o_label4_data6[26]));
Q_FDP4EP \o_label4_data6_REG[27] ( .CK(clk), .CE(n165), .R(n261), .D(n33), .Q(o_label4_data6[27]));
Q_FDP4EP \o_label4_data6_REG[28] ( .CK(clk), .CE(n165), .R(n261), .D(n34), .Q(o_label4_data6[28]));
Q_FDP4EP \o_label4_data6_REG[29] ( .CK(clk), .CE(n165), .R(n261), .D(n35), .Q(o_label4_data6[29]));
Q_FDP4EP \o_label4_data6_REG[30] ( .CK(clk), .CE(n165), .R(n261), .D(n36), .Q(o_label4_data6[30]));
Q_FDP4EP \o_label4_data6_REG[31] ( .CK(clk), .CE(n165), .R(n261), .D(n37), .Q(o_label4_data6[31]));
Q_FDP4EP \o_label4_data7_REG[0] ( .CK(clk), .CE(n164), .R(n261), .D(n6), .Q(o_label4_data7[0]));
Q_FDP4EP \o_label4_data7_REG[1] ( .CK(clk), .CE(n164), .R(n261), .D(n7), .Q(o_label4_data7[1]));
Q_FDP4EP \o_label4_data7_REG[2] ( .CK(clk), .CE(n164), .R(n261), .D(n8), .Q(o_label4_data7[2]));
Q_FDP4EP \o_label4_data7_REG[3] ( .CK(clk), .CE(n164), .R(n261), .D(n9), .Q(o_label4_data7[3]));
Q_FDP4EP \o_label4_data7_REG[4] ( .CK(clk), .CE(n164), .R(n261), .D(n10), .Q(o_label4_data7[4]));
Q_FDP4EP \o_label4_data7_REG[5] ( .CK(clk), .CE(n164), .R(n261), .D(n11), .Q(o_label4_data7[5]));
Q_FDP4EP \o_label4_data7_REG[6] ( .CK(clk), .CE(n164), .R(n261), .D(n12), .Q(o_label4_data7[6]));
Q_FDP4EP \o_label4_data7_REG[7] ( .CK(clk), .CE(n164), .R(n261), .D(n13), .Q(o_label4_data7[7]));
Q_FDP4EP \o_label4_data7_REG[8] ( .CK(clk), .CE(n164), .R(n261), .D(n14), .Q(o_label4_data7[8]));
Q_FDP4EP \o_label4_data7_REG[9] ( .CK(clk), .CE(n164), .R(n261), .D(n15), .Q(o_label4_data7[9]));
Q_FDP4EP \o_label4_data7_REG[10] ( .CK(clk), .CE(n164), .R(n261), .D(n16), .Q(o_label4_data7[10]));
Q_FDP4EP \o_label4_data7_REG[11] ( .CK(clk), .CE(n164), .R(n261), .D(n17), .Q(o_label4_data7[11]));
Q_FDP4EP \o_label4_data7_REG[12] ( .CK(clk), .CE(n164), .R(n261), .D(n18), .Q(o_label4_data7[12]));
Q_FDP4EP \o_label4_data7_REG[13] ( .CK(clk), .CE(n164), .R(n261), .D(n19), .Q(o_label4_data7[13]));
Q_FDP4EP \o_label4_data7_REG[14] ( .CK(clk), .CE(n164), .R(n261), .D(n20), .Q(o_label4_data7[14]));
Q_FDP4EP \o_label4_data7_REG[15] ( .CK(clk), .CE(n164), .R(n261), .D(n21), .Q(o_label4_data7[15]));
Q_FDP4EP \o_label4_data7_REG[16] ( .CK(clk), .CE(n164), .R(n261), .D(n22), .Q(o_label4_data7[16]));
Q_FDP4EP \o_label4_data7_REG[17] ( .CK(clk), .CE(n164), .R(n261), .D(n23), .Q(o_label4_data7[17]));
Q_FDP4EP \o_label4_data7_REG[18] ( .CK(clk), .CE(n164), .R(n261), .D(n24), .Q(o_label4_data7[18]));
Q_FDP4EP \o_label4_data7_REG[19] ( .CK(clk), .CE(n164), .R(n261), .D(n25), .Q(o_label4_data7[19]));
Q_FDP4EP \o_label4_data7_REG[20] ( .CK(clk), .CE(n164), .R(n261), .D(n26), .Q(o_label4_data7[20]));
Q_FDP4EP \o_label4_data7_REG[21] ( .CK(clk), .CE(n164), .R(n261), .D(n27), .Q(o_label4_data7[21]));
Q_FDP4EP \o_label4_data7_REG[22] ( .CK(clk), .CE(n164), .R(n261), .D(n28), .Q(o_label4_data7[22]));
Q_FDP4EP \o_label4_data7_REG[23] ( .CK(clk), .CE(n164), .R(n261), .D(n29), .Q(o_label4_data7[23]));
Q_FDP4EP \o_label4_data7_REG[24] ( .CK(clk), .CE(n164), .R(n261), .D(n30), .Q(o_label4_data7[24]));
Q_FDP4EP \o_label4_data7_REG[25] ( .CK(clk), .CE(n164), .R(n261), .D(n31), .Q(o_label4_data7[25]));
Q_FDP4EP \o_label4_data7_REG[26] ( .CK(clk), .CE(n164), .R(n261), .D(n32), .Q(o_label4_data7[26]));
Q_FDP4EP \o_label4_data7_REG[27] ( .CK(clk), .CE(n164), .R(n261), .D(n33), .Q(o_label4_data7[27]));
Q_FDP4EP \o_label4_data7_REG[28] ( .CK(clk), .CE(n164), .R(n261), .D(n34), .Q(o_label4_data7[28]));
Q_FDP4EP \o_label4_data7_REG[29] ( .CK(clk), .CE(n164), .R(n261), .D(n35), .Q(o_label4_data7[29]));
Q_FDP4EP \o_label4_data7_REG[30] ( .CK(clk), .CE(n164), .R(n261), .D(n36), .Q(o_label4_data7[30]));
Q_FDP4EP \o_label4_data7_REG[31] ( .CK(clk), .CE(n164), .R(n261), .D(n37), .Q(o_label4_data7[31]));
Q_FDP4EP \o_label4_config_REG[0] ( .CK(clk), .CE(n163), .R(n261), .D(n6), .Q(o_label4_config[0]));
Q_FDP4EP \o_label4_config_REG[1] ( .CK(clk), .CE(n163), .R(n261), .D(n7), .Q(o_label4_config[1]));
Q_FDP4EP \o_label4_config_REG[2] ( .CK(clk), .CE(n163), .R(n261), .D(n8), .Q(o_label4_config[2]));
Q_FDP4EP \o_label4_config_REG[3] ( .CK(clk), .CE(n163), .R(n261), .D(n9), .Q(o_label4_config[3]));
Q_FDP4EP \o_label4_config_REG[4] ( .CK(clk), .CE(n163), .R(n261), .D(n10), .Q(o_label4_config[4]));
Q_FDP4EP \o_label4_config_REG[5] ( .CK(clk), .CE(n163), .R(n261), .D(n11), .Q(o_label4_config[5]));
Q_FDP4EP \o_label4_config_REG[6] ( .CK(clk), .CE(n163), .R(n261), .D(n12), .Q(o_label4_config[6]));
Q_FDP4EP \o_label4_config_REG[7] ( .CK(clk), .CE(n163), .R(n261), .D(n13), .Q(o_label4_config[7]));
Q_FDP4EP \o_label4_config_REG[9] ( .CK(clk), .CE(n163), .R(n261), .D(n31), .Q(o_label4_config[9]));
Q_FDP4EP \o_label4_config_REG[10] ( .CK(clk), .CE(n163), .R(n261), .D(n32), .Q(o_label4_config[10]));
Q_FDP4EP \o_label4_config_REG[11] ( .CK(clk), .CE(n163), .R(n261), .D(n33), .Q(o_label4_config[11]));
Q_FDP4EP \o_label4_config_REG[12] ( .CK(clk), .CE(n163), .R(n261), .D(n34), .Q(o_label4_config[12]));
Q_FDP4EP \o_label4_config_REG[13] ( .CK(clk), .CE(n163), .R(n261), .D(n35), .Q(o_label4_config[13]));
Q_FDP4EP \o_label4_config_REG[14] ( .CK(clk), .CE(n163), .R(n261), .D(n36), .Q(o_label4_config[14]));
Q_FDP4EP \o_label4_config_REG[15] ( .CK(clk), .CE(n163), .R(n261), .D(n37), .Q(o_label4_config[15]));
Q_FDP4EP \o_label3_data0_REG[0] ( .CK(clk), .CE(n162), .R(n261), .D(n6), .Q(o_label3_data0[0]));
Q_FDP4EP \o_label3_data0_REG[1] ( .CK(clk), .CE(n162), .R(n261), .D(n7), .Q(o_label3_data0[1]));
Q_FDP4EP \o_label3_data0_REG[2] ( .CK(clk), .CE(n162), .R(n261), .D(n8), .Q(o_label3_data0[2]));
Q_FDP4EP \o_label3_data0_REG[3] ( .CK(clk), .CE(n162), .R(n261), .D(n9), .Q(o_label3_data0[3]));
Q_FDP4EP \o_label3_data0_REG[4] ( .CK(clk), .CE(n162), .R(n261), .D(n10), .Q(o_label3_data0[4]));
Q_FDP4EP \o_label3_data0_REG[5] ( .CK(clk), .CE(n162), .R(n261), .D(n11), .Q(o_label3_data0[5]));
Q_FDP4EP \o_label3_data0_REG[6] ( .CK(clk), .CE(n162), .R(n261), .D(n12), .Q(o_label3_data0[6]));
Q_FDP4EP \o_label3_data0_REG[7] ( .CK(clk), .CE(n162), .R(n261), .D(n13), .Q(o_label3_data0[7]));
Q_FDP4EP \o_label3_data0_REG[8] ( .CK(clk), .CE(n162), .R(n261), .D(n14), .Q(o_label3_data0[8]));
Q_FDP4EP \o_label3_data0_REG[9] ( .CK(clk), .CE(n162), .R(n261), .D(n15), .Q(o_label3_data0[9]));
Q_FDP4EP \o_label3_data0_REG[10] ( .CK(clk), .CE(n162), .R(n261), .D(n16), .Q(o_label3_data0[10]));
Q_FDP4EP \o_label3_data0_REG[11] ( .CK(clk), .CE(n162), .R(n261), .D(n17), .Q(o_label3_data0[11]));
Q_FDP4EP \o_label3_data0_REG[12] ( .CK(clk), .CE(n162), .R(n261), .D(n18), .Q(o_label3_data0[12]));
Q_FDP4EP \o_label3_data0_REG[13] ( .CK(clk), .CE(n162), .R(n261), .D(n19), .Q(o_label3_data0[13]));
Q_FDP4EP \o_label3_data0_REG[14] ( .CK(clk), .CE(n162), .R(n261), .D(n20), .Q(o_label3_data0[14]));
Q_FDP4EP \o_label3_data0_REG[15] ( .CK(clk), .CE(n162), .R(n261), .D(n21), .Q(o_label3_data0[15]));
Q_FDP4EP \o_label3_data0_REG[16] ( .CK(clk), .CE(n162), .R(n261), .D(n22), .Q(o_label3_data0[16]));
Q_FDP4EP \o_label3_data0_REG[17] ( .CK(clk), .CE(n162), .R(n261), .D(n23), .Q(o_label3_data0[17]));
Q_FDP4EP \o_label3_data0_REG[18] ( .CK(clk), .CE(n162), .R(n261), .D(n24), .Q(o_label3_data0[18]));
Q_FDP4EP \o_label3_data0_REG[19] ( .CK(clk), .CE(n162), .R(n261), .D(n25), .Q(o_label3_data0[19]));
Q_FDP4EP \o_label3_data0_REG[20] ( .CK(clk), .CE(n162), .R(n261), .D(n26), .Q(o_label3_data0[20]));
Q_FDP4EP \o_label3_data0_REG[21] ( .CK(clk), .CE(n162), .R(n261), .D(n27), .Q(o_label3_data0[21]));
Q_FDP4EP \o_label3_data0_REG[22] ( .CK(clk), .CE(n162), .R(n261), .D(n28), .Q(o_label3_data0[22]));
Q_FDP4EP \o_label3_data0_REG[23] ( .CK(clk), .CE(n162), .R(n261), .D(n29), .Q(o_label3_data0[23]));
Q_FDP4EP \o_label3_data0_REG[24] ( .CK(clk), .CE(n162), .R(n261), .D(n30), .Q(o_label3_data0[24]));
Q_FDP4EP \o_label3_data0_REG[25] ( .CK(clk), .CE(n162), .R(n261), .D(n31), .Q(o_label3_data0[25]));
Q_FDP4EP \o_label3_data0_REG[26] ( .CK(clk), .CE(n162), .R(n261), .D(n32), .Q(o_label3_data0[26]));
Q_FDP4EP \o_label3_data0_REG[27] ( .CK(clk), .CE(n162), .R(n261), .D(n33), .Q(o_label3_data0[27]));
Q_FDP4EP \o_label3_data0_REG[28] ( .CK(clk), .CE(n162), .R(n261), .D(n34), .Q(o_label3_data0[28]));
Q_FDP4EP \o_label3_data0_REG[29] ( .CK(clk), .CE(n162), .R(n261), .D(n35), .Q(o_label3_data0[29]));
Q_FDP4EP \o_label3_data0_REG[30] ( .CK(clk), .CE(n162), .R(n261), .D(n36), .Q(o_label3_data0[30]));
Q_FDP4EP \o_label3_data0_REG[31] ( .CK(clk), .CE(n162), .R(n261), .D(n37), .Q(o_label3_data0[31]));
Q_FDP4EP \o_label3_data1_REG[0] ( .CK(clk), .CE(n161), .R(n261), .D(n6), .Q(o_label3_data1[0]));
Q_FDP4EP \o_label3_data1_REG[1] ( .CK(clk), .CE(n161), .R(n261), .D(n7), .Q(o_label3_data1[1]));
Q_FDP4EP \o_label3_data1_REG[2] ( .CK(clk), .CE(n161), .R(n261), .D(n8), .Q(o_label3_data1[2]));
Q_FDP4EP \o_label3_data1_REG[3] ( .CK(clk), .CE(n161), .R(n261), .D(n9), .Q(o_label3_data1[3]));
Q_FDP4EP \o_label3_data1_REG[4] ( .CK(clk), .CE(n161), .R(n261), .D(n10), .Q(o_label3_data1[4]));
Q_FDP4EP \o_label3_data1_REG[5] ( .CK(clk), .CE(n161), .R(n261), .D(n11), .Q(o_label3_data1[5]));
Q_FDP4EP \o_label3_data1_REG[6] ( .CK(clk), .CE(n161), .R(n261), .D(n12), .Q(o_label3_data1[6]));
Q_FDP4EP \o_label3_data1_REG[7] ( .CK(clk), .CE(n161), .R(n261), .D(n13), .Q(o_label3_data1[7]));
Q_FDP4EP \o_label3_data1_REG[8] ( .CK(clk), .CE(n161), .R(n261), .D(n14), .Q(o_label3_data1[8]));
Q_FDP4EP \o_label3_data1_REG[9] ( .CK(clk), .CE(n161), .R(n261), .D(n15), .Q(o_label3_data1[9]));
Q_FDP4EP \o_label3_data1_REG[10] ( .CK(clk), .CE(n161), .R(n261), .D(n16), .Q(o_label3_data1[10]));
Q_FDP4EP \o_label3_data1_REG[11] ( .CK(clk), .CE(n161), .R(n261), .D(n17), .Q(o_label3_data1[11]));
Q_FDP4EP \o_label3_data1_REG[12] ( .CK(clk), .CE(n161), .R(n261), .D(n18), .Q(o_label3_data1[12]));
Q_FDP4EP \o_label3_data1_REG[13] ( .CK(clk), .CE(n161), .R(n261), .D(n19), .Q(o_label3_data1[13]));
Q_FDP4EP \o_label3_data1_REG[14] ( .CK(clk), .CE(n161), .R(n261), .D(n20), .Q(o_label3_data1[14]));
Q_FDP4EP \o_label3_data1_REG[15] ( .CK(clk), .CE(n161), .R(n261), .D(n21), .Q(o_label3_data1[15]));
Q_FDP4EP \o_label3_data1_REG[16] ( .CK(clk), .CE(n161), .R(n261), .D(n22), .Q(o_label3_data1[16]));
Q_FDP4EP \o_label3_data1_REG[17] ( .CK(clk), .CE(n161), .R(n261), .D(n23), .Q(o_label3_data1[17]));
Q_FDP4EP \o_label3_data1_REG[18] ( .CK(clk), .CE(n161), .R(n261), .D(n24), .Q(o_label3_data1[18]));
Q_FDP4EP \o_label3_data1_REG[19] ( .CK(clk), .CE(n161), .R(n261), .D(n25), .Q(o_label3_data1[19]));
Q_FDP4EP \o_label3_data1_REG[20] ( .CK(clk), .CE(n161), .R(n261), .D(n26), .Q(o_label3_data1[20]));
Q_FDP4EP \o_label3_data1_REG[21] ( .CK(clk), .CE(n161), .R(n261), .D(n27), .Q(o_label3_data1[21]));
Q_FDP4EP \o_label3_data1_REG[22] ( .CK(clk), .CE(n161), .R(n261), .D(n28), .Q(o_label3_data1[22]));
Q_FDP4EP \o_label3_data1_REG[23] ( .CK(clk), .CE(n161), .R(n261), .D(n29), .Q(o_label3_data1[23]));
Q_FDP4EP \o_label3_data1_REG[24] ( .CK(clk), .CE(n161), .R(n261), .D(n30), .Q(o_label3_data1[24]));
Q_FDP4EP \o_label3_data1_REG[25] ( .CK(clk), .CE(n161), .R(n261), .D(n31), .Q(o_label3_data1[25]));
Q_FDP4EP \o_label3_data1_REG[26] ( .CK(clk), .CE(n161), .R(n261), .D(n32), .Q(o_label3_data1[26]));
Q_FDP4EP \o_label3_data1_REG[27] ( .CK(clk), .CE(n161), .R(n261), .D(n33), .Q(o_label3_data1[27]));
Q_FDP4EP \o_label3_data1_REG[28] ( .CK(clk), .CE(n161), .R(n261), .D(n34), .Q(o_label3_data1[28]));
Q_FDP4EP \o_label3_data1_REG[29] ( .CK(clk), .CE(n161), .R(n261), .D(n35), .Q(o_label3_data1[29]));
Q_FDP4EP \o_label3_data1_REG[30] ( .CK(clk), .CE(n161), .R(n261), .D(n36), .Q(o_label3_data1[30]));
Q_FDP4EP \o_label3_data1_REG[31] ( .CK(clk), .CE(n161), .R(n261), .D(n37), .Q(o_label3_data1[31]));
Q_FDP4EP \o_label3_data2_REG[0] ( .CK(clk), .CE(n160), .R(n261), .D(n6), .Q(o_label3_data2[0]));
Q_FDP4EP \o_label3_data2_REG[1] ( .CK(clk), .CE(n160), .R(n261), .D(n7), .Q(o_label3_data2[1]));
Q_FDP4EP \o_label3_data2_REG[2] ( .CK(clk), .CE(n160), .R(n261), .D(n8), .Q(o_label3_data2[2]));
Q_FDP4EP \o_label3_data2_REG[3] ( .CK(clk), .CE(n160), .R(n261), .D(n9), .Q(o_label3_data2[3]));
Q_FDP4EP \o_label3_data2_REG[4] ( .CK(clk), .CE(n160), .R(n261), .D(n10), .Q(o_label3_data2[4]));
Q_FDP4EP \o_label3_data2_REG[5] ( .CK(clk), .CE(n160), .R(n261), .D(n11), .Q(o_label3_data2[5]));
Q_FDP4EP \o_label3_data2_REG[6] ( .CK(clk), .CE(n160), .R(n261), .D(n12), .Q(o_label3_data2[6]));
Q_FDP4EP \o_label3_data2_REG[7] ( .CK(clk), .CE(n160), .R(n261), .D(n13), .Q(o_label3_data2[7]));
Q_FDP4EP \o_label3_data2_REG[8] ( .CK(clk), .CE(n160), .R(n261), .D(n14), .Q(o_label3_data2[8]));
Q_FDP4EP \o_label3_data2_REG[9] ( .CK(clk), .CE(n160), .R(n261), .D(n15), .Q(o_label3_data2[9]));
Q_FDP4EP \o_label3_data2_REG[10] ( .CK(clk), .CE(n160), .R(n261), .D(n16), .Q(o_label3_data2[10]));
Q_FDP4EP \o_label3_data2_REG[11] ( .CK(clk), .CE(n160), .R(n261), .D(n17), .Q(o_label3_data2[11]));
Q_FDP4EP \o_label3_data2_REG[12] ( .CK(clk), .CE(n160), .R(n261), .D(n18), .Q(o_label3_data2[12]));
Q_FDP4EP \o_label3_data2_REG[13] ( .CK(clk), .CE(n160), .R(n261), .D(n19), .Q(o_label3_data2[13]));
Q_FDP4EP \o_label3_data2_REG[14] ( .CK(clk), .CE(n160), .R(n261), .D(n20), .Q(o_label3_data2[14]));
Q_FDP4EP \o_label3_data2_REG[15] ( .CK(clk), .CE(n160), .R(n261), .D(n21), .Q(o_label3_data2[15]));
Q_FDP4EP \o_label3_data2_REG[16] ( .CK(clk), .CE(n160), .R(n261), .D(n22), .Q(o_label3_data2[16]));
Q_FDP4EP \o_label3_data2_REG[17] ( .CK(clk), .CE(n160), .R(n261), .D(n23), .Q(o_label3_data2[17]));
Q_FDP4EP \o_label3_data2_REG[18] ( .CK(clk), .CE(n160), .R(n261), .D(n24), .Q(o_label3_data2[18]));
Q_FDP4EP \o_label3_data2_REG[19] ( .CK(clk), .CE(n160), .R(n261), .D(n25), .Q(o_label3_data2[19]));
Q_FDP4EP \o_label3_data2_REG[20] ( .CK(clk), .CE(n160), .R(n261), .D(n26), .Q(o_label3_data2[20]));
Q_FDP4EP \o_label3_data2_REG[21] ( .CK(clk), .CE(n160), .R(n261), .D(n27), .Q(o_label3_data2[21]));
Q_FDP4EP \o_label3_data2_REG[22] ( .CK(clk), .CE(n160), .R(n261), .D(n28), .Q(o_label3_data2[22]));
Q_FDP4EP \o_label3_data2_REG[23] ( .CK(clk), .CE(n160), .R(n261), .D(n29), .Q(o_label3_data2[23]));
Q_FDP4EP \o_label3_data2_REG[24] ( .CK(clk), .CE(n160), .R(n261), .D(n30), .Q(o_label3_data2[24]));
Q_FDP4EP \o_label3_data2_REG[25] ( .CK(clk), .CE(n160), .R(n261), .D(n31), .Q(o_label3_data2[25]));
Q_FDP4EP \o_label3_data2_REG[26] ( .CK(clk), .CE(n160), .R(n261), .D(n32), .Q(o_label3_data2[26]));
Q_FDP4EP \o_label3_data2_REG[27] ( .CK(clk), .CE(n160), .R(n261), .D(n33), .Q(o_label3_data2[27]));
Q_FDP4EP \o_label3_data2_REG[28] ( .CK(clk), .CE(n160), .R(n261), .D(n34), .Q(o_label3_data2[28]));
Q_FDP4EP \o_label3_data2_REG[29] ( .CK(clk), .CE(n160), .R(n261), .D(n35), .Q(o_label3_data2[29]));
Q_FDP4EP \o_label3_data2_REG[30] ( .CK(clk), .CE(n160), .R(n261), .D(n36), .Q(o_label3_data2[30]));
Q_FDP4EP \o_label3_data2_REG[31] ( .CK(clk), .CE(n160), .R(n261), .D(n37), .Q(o_label3_data2[31]));
Q_FDP4EP \o_label3_data3_REG[0] ( .CK(clk), .CE(n159), .R(n261), .D(n6), .Q(o_label3_data3[0]));
Q_FDP4EP \o_label3_data3_REG[1] ( .CK(clk), .CE(n159), .R(n261), .D(n7), .Q(o_label3_data3[1]));
Q_FDP4EP \o_label3_data3_REG[2] ( .CK(clk), .CE(n159), .R(n261), .D(n8), .Q(o_label3_data3[2]));
Q_FDP4EP \o_label3_data3_REG[3] ( .CK(clk), .CE(n159), .R(n261), .D(n9), .Q(o_label3_data3[3]));
Q_FDP4EP \o_label3_data3_REG[4] ( .CK(clk), .CE(n159), .R(n261), .D(n10), .Q(o_label3_data3[4]));
Q_FDP4EP \o_label3_data3_REG[5] ( .CK(clk), .CE(n159), .R(n261), .D(n11), .Q(o_label3_data3[5]));
Q_FDP4EP \o_label3_data3_REG[6] ( .CK(clk), .CE(n159), .R(n261), .D(n12), .Q(o_label3_data3[6]));
Q_FDP4EP \o_label3_data3_REG[7] ( .CK(clk), .CE(n159), .R(n261), .D(n13), .Q(o_label3_data3[7]));
Q_FDP4EP \o_label3_data3_REG[8] ( .CK(clk), .CE(n159), .R(n261), .D(n14), .Q(o_label3_data3[8]));
Q_FDP4EP \o_label3_data3_REG[9] ( .CK(clk), .CE(n159), .R(n261), .D(n15), .Q(o_label3_data3[9]));
Q_FDP4EP \o_label3_data3_REG[10] ( .CK(clk), .CE(n159), .R(n261), .D(n16), .Q(o_label3_data3[10]));
Q_FDP4EP \o_label3_data3_REG[11] ( .CK(clk), .CE(n159), .R(n261), .D(n17), .Q(o_label3_data3[11]));
Q_FDP4EP \o_label3_data3_REG[12] ( .CK(clk), .CE(n159), .R(n261), .D(n18), .Q(o_label3_data3[12]));
Q_FDP4EP \o_label3_data3_REG[13] ( .CK(clk), .CE(n159), .R(n261), .D(n19), .Q(o_label3_data3[13]));
Q_FDP4EP \o_label3_data3_REG[14] ( .CK(clk), .CE(n159), .R(n261), .D(n20), .Q(o_label3_data3[14]));
Q_FDP4EP \o_label3_data3_REG[15] ( .CK(clk), .CE(n159), .R(n261), .D(n21), .Q(o_label3_data3[15]));
Q_FDP4EP \o_label3_data3_REG[16] ( .CK(clk), .CE(n159), .R(n261), .D(n22), .Q(o_label3_data3[16]));
Q_FDP4EP \o_label3_data3_REG[17] ( .CK(clk), .CE(n159), .R(n261), .D(n23), .Q(o_label3_data3[17]));
Q_FDP4EP \o_label3_data3_REG[18] ( .CK(clk), .CE(n159), .R(n261), .D(n24), .Q(o_label3_data3[18]));
Q_FDP4EP \o_label3_data3_REG[19] ( .CK(clk), .CE(n159), .R(n261), .D(n25), .Q(o_label3_data3[19]));
Q_FDP4EP \o_label3_data3_REG[20] ( .CK(clk), .CE(n159), .R(n261), .D(n26), .Q(o_label3_data3[20]));
Q_FDP4EP \o_label3_data3_REG[21] ( .CK(clk), .CE(n159), .R(n261), .D(n27), .Q(o_label3_data3[21]));
Q_FDP4EP \o_label3_data3_REG[22] ( .CK(clk), .CE(n159), .R(n261), .D(n28), .Q(o_label3_data3[22]));
Q_FDP4EP \o_label3_data3_REG[23] ( .CK(clk), .CE(n159), .R(n261), .D(n29), .Q(o_label3_data3[23]));
Q_FDP4EP \o_label3_data3_REG[24] ( .CK(clk), .CE(n159), .R(n261), .D(n30), .Q(o_label3_data3[24]));
Q_FDP4EP \o_label3_data3_REG[25] ( .CK(clk), .CE(n159), .R(n261), .D(n31), .Q(o_label3_data3[25]));
Q_FDP4EP \o_label3_data3_REG[26] ( .CK(clk), .CE(n159), .R(n261), .D(n32), .Q(o_label3_data3[26]));
Q_FDP4EP \o_label3_data3_REG[27] ( .CK(clk), .CE(n159), .R(n261), .D(n33), .Q(o_label3_data3[27]));
Q_FDP4EP \o_label3_data3_REG[28] ( .CK(clk), .CE(n159), .R(n261), .D(n34), .Q(o_label3_data3[28]));
Q_FDP4EP \o_label3_data3_REG[29] ( .CK(clk), .CE(n159), .R(n261), .D(n35), .Q(o_label3_data3[29]));
Q_FDP4EP \o_label3_data3_REG[30] ( .CK(clk), .CE(n159), .R(n261), .D(n36), .Q(o_label3_data3[30]));
Q_FDP4EP \o_label3_data3_REG[31] ( .CK(clk), .CE(n159), .R(n261), .D(n37), .Q(o_label3_data3[31]));
Q_FDP4EP \o_label3_data4_REG[0] ( .CK(clk), .CE(n158), .R(n261), .D(n6), .Q(o_label3_data4[0]));
Q_FDP4EP \o_label3_data4_REG[1] ( .CK(clk), .CE(n158), .R(n261), .D(n7), .Q(o_label3_data4[1]));
Q_FDP4EP \o_label3_data4_REG[2] ( .CK(clk), .CE(n158), .R(n261), .D(n8), .Q(o_label3_data4[2]));
Q_FDP4EP \o_label3_data4_REG[3] ( .CK(clk), .CE(n158), .R(n261), .D(n9), .Q(o_label3_data4[3]));
Q_FDP4EP \o_label3_data4_REG[4] ( .CK(clk), .CE(n158), .R(n261), .D(n10), .Q(o_label3_data4[4]));
Q_FDP4EP \o_label3_data4_REG[5] ( .CK(clk), .CE(n158), .R(n261), .D(n11), .Q(o_label3_data4[5]));
Q_FDP4EP \o_label3_data4_REG[6] ( .CK(clk), .CE(n158), .R(n261), .D(n12), .Q(o_label3_data4[6]));
Q_FDP4EP \o_label3_data4_REG[7] ( .CK(clk), .CE(n158), .R(n261), .D(n13), .Q(o_label3_data4[7]));
Q_FDP4EP \o_label3_data4_REG[8] ( .CK(clk), .CE(n158), .R(n261), .D(n14), .Q(o_label3_data4[8]));
Q_FDP4EP \o_label3_data4_REG[9] ( .CK(clk), .CE(n158), .R(n261), .D(n15), .Q(o_label3_data4[9]));
Q_FDP4EP \o_label3_data4_REG[10] ( .CK(clk), .CE(n158), .R(n261), .D(n16), .Q(o_label3_data4[10]));
Q_FDP4EP \o_label3_data4_REG[11] ( .CK(clk), .CE(n158), .R(n261), .D(n17), .Q(o_label3_data4[11]));
Q_FDP4EP \o_label3_data4_REG[12] ( .CK(clk), .CE(n158), .R(n261), .D(n18), .Q(o_label3_data4[12]));
Q_FDP4EP \o_label3_data4_REG[13] ( .CK(clk), .CE(n158), .R(n261), .D(n19), .Q(o_label3_data4[13]));
Q_FDP4EP \o_label3_data4_REG[14] ( .CK(clk), .CE(n158), .R(n261), .D(n20), .Q(o_label3_data4[14]));
Q_FDP4EP \o_label3_data4_REG[15] ( .CK(clk), .CE(n158), .R(n261), .D(n21), .Q(o_label3_data4[15]));
Q_FDP4EP \o_label3_data4_REG[16] ( .CK(clk), .CE(n158), .R(n261), .D(n22), .Q(o_label3_data4[16]));
Q_FDP4EP \o_label3_data4_REG[17] ( .CK(clk), .CE(n158), .R(n261), .D(n23), .Q(o_label3_data4[17]));
Q_FDP4EP \o_label3_data4_REG[18] ( .CK(clk), .CE(n158), .R(n261), .D(n24), .Q(o_label3_data4[18]));
Q_FDP4EP \o_label3_data4_REG[19] ( .CK(clk), .CE(n158), .R(n261), .D(n25), .Q(o_label3_data4[19]));
Q_FDP4EP \o_label3_data4_REG[20] ( .CK(clk), .CE(n158), .R(n261), .D(n26), .Q(o_label3_data4[20]));
Q_FDP4EP \o_label3_data4_REG[21] ( .CK(clk), .CE(n158), .R(n261), .D(n27), .Q(o_label3_data4[21]));
Q_FDP4EP \o_label3_data4_REG[22] ( .CK(clk), .CE(n158), .R(n261), .D(n28), .Q(o_label3_data4[22]));
Q_FDP4EP \o_label3_data4_REG[23] ( .CK(clk), .CE(n158), .R(n261), .D(n29), .Q(o_label3_data4[23]));
Q_FDP4EP \o_label3_data4_REG[24] ( .CK(clk), .CE(n158), .R(n261), .D(n30), .Q(o_label3_data4[24]));
Q_FDP4EP \o_label3_data4_REG[25] ( .CK(clk), .CE(n158), .R(n261), .D(n31), .Q(o_label3_data4[25]));
Q_FDP4EP \o_label3_data4_REG[26] ( .CK(clk), .CE(n158), .R(n261), .D(n32), .Q(o_label3_data4[26]));
Q_FDP4EP \o_label3_data4_REG[27] ( .CK(clk), .CE(n158), .R(n261), .D(n33), .Q(o_label3_data4[27]));
Q_FDP4EP \o_label3_data4_REG[28] ( .CK(clk), .CE(n158), .R(n261), .D(n34), .Q(o_label3_data4[28]));
Q_FDP4EP \o_label3_data4_REG[29] ( .CK(clk), .CE(n158), .R(n261), .D(n35), .Q(o_label3_data4[29]));
Q_FDP4EP \o_label3_data4_REG[30] ( .CK(clk), .CE(n158), .R(n261), .D(n36), .Q(o_label3_data4[30]));
Q_FDP4EP \o_label3_data4_REG[31] ( .CK(clk), .CE(n158), .R(n261), .D(n37), .Q(o_label3_data4[31]));
Q_FDP4EP \o_label3_data5_REG[0] ( .CK(clk), .CE(n157), .R(n261), .D(n6), .Q(o_label3_data5[0]));
Q_FDP4EP \o_label3_data5_REG[1] ( .CK(clk), .CE(n157), .R(n261), .D(n7), .Q(o_label3_data5[1]));
Q_FDP4EP \o_label3_data5_REG[2] ( .CK(clk), .CE(n157), .R(n261), .D(n8), .Q(o_label3_data5[2]));
Q_FDP4EP \o_label3_data5_REG[3] ( .CK(clk), .CE(n157), .R(n261), .D(n9), .Q(o_label3_data5[3]));
Q_FDP4EP \o_label3_data5_REG[4] ( .CK(clk), .CE(n157), .R(n261), .D(n10), .Q(o_label3_data5[4]));
Q_FDP4EP \o_label3_data5_REG[5] ( .CK(clk), .CE(n157), .R(n261), .D(n11), .Q(o_label3_data5[5]));
Q_FDP4EP \o_label3_data5_REG[6] ( .CK(clk), .CE(n157), .R(n261), .D(n12), .Q(o_label3_data5[6]));
Q_FDP4EP \o_label3_data5_REG[7] ( .CK(clk), .CE(n157), .R(n261), .D(n13), .Q(o_label3_data5[7]));
Q_FDP4EP \o_label3_data5_REG[8] ( .CK(clk), .CE(n157), .R(n261), .D(n14), .Q(o_label3_data5[8]));
Q_FDP4EP \o_label3_data5_REG[9] ( .CK(clk), .CE(n157), .R(n261), .D(n15), .Q(o_label3_data5[9]));
Q_FDP4EP \o_label3_data5_REG[10] ( .CK(clk), .CE(n157), .R(n261), .D(n16), .Q(o_label3_data5[10]));
Q_FDP4EP \o_label3_data5_REG[11] ( .CK(clk), .CE(n157), .R(n261), .D(n17), .Q(o_label3_data5[11]));
Q_FDP4EP \o_label3_data5_REG[12] ( .CK(clk), .CE(n157), .R(n261), .D(n18), .Q(o_label3_data5[12]));
Q_FDP4EP \o_label3_data5_REG[13] ( .CK(clk), .CE(n157), .R(n261), .D(n19), .Q(o_label3_data5[13]));
Q_FDP4EP \o_label3_data5_REG[14] ( .CK(clk), .CE(n157), .R(n261), .D(n20), .Q(o_label3_data5[14]));
Q_FDP4EP \o_label3_data5_REG[15] ( .CK(clk), .CE(n157), .R(n261), .D(n21), .Q(o_label3_data5[15]));
Q_FDP4EP \o_label3_data5_REG[16] ( .CK(clk), .CE(n157), .R(n261), .D(n22), .Q(o_label3_data5[16]));
Q_FDP4EP \o_label3_data5_REG[17] ( .CK(clk), .CE(n157), .R(n261), .D(n23), .Q(o_label3_data5[17]));
Q_FDP4EP \o_label3_data5_REG[18] ( .CK(clk), .CE(n157), .R(n261), .D(n24), .Q(o_label3_data5[18]));
Q_FDP4EP \o_label3_data5_REG[19] ( .CK(clk), .CE(n157), .R(n261), .D(n25), .Q(o_label3_data5[19]));
Q_FDP4EP \o_label3_data5_REG[20] ( .CK(clk), .CE(n157), .R(n261), .D(n26), .Q(o_label3_data5[20]));
Q_FDP4EP \o_label3_data5_REG[21] ( .CK(clk), .CE(n157), .R(n261), .D(n27), .Q(o_label3_data5[21]));
Q_FDP4EP \o_label3_data5_REG[22] ( .CK(clk), .CE(n157), .R(n261), .D(n28), .Q(o_label3_data5[22]));
Q_FDP4EP \o_label3_data5_REG[23] ( .CK(clk), .CE(n157), .R(n261), .D(n29), .Q(o_label3_data5[23]));
Q_FDP4EP \o_label3_data5_REG[24] ( .CK(clk), .CE(n157), .R(n261), .D(n30), .Q(o_label3_data5[24]));
Q_FDP4EP \o_label3_data5_REG[25] ( .CK(clk), .CE(n157), .R(n261), .D(n31), .Q(o_label3_data5[25]));
Q_FDP4EP \o_label3_data5_REG[26] ( .CK(clk), .CE(n157), .R(n261), .D(n32), .Q(o_label3_data5[26]));
Q_FDP4EP \o_label3_data5_REG[27] ( .CK(clk), .CE(n157), .R(n261), .D(n33), .Q(o_label3_data5[27]));
Q_FDP4EP \o_label3_data5_REG[28] ( .CK(clk), .CE(n157), .R(n261), .D(n34), .Q(o_label3_data5[28]));
Q_FDP4EP \o_label3_data5_REG[29] ( .CK(clk), .CE(n157), .R(n261), .D(n35), .Q(o_label3_data5[29]));
Q_FDP4EP \o_label3_data5_REG[30] ( .CK(clk), .CE(n157), .R(n261), .D(n36), .Q(o_label3_data5[30]));
Q_FDP4EP \o_label3_data5_REG[31] ( .CK(clk), .CE(n157), .R(n261), .D(n37), .Q(o_label3_data5[31]));
Q_FDP4EP \o_label3_data6_REG[0] ( .CK(clk), .CE(n156), .R(n261), .D(n6), .Q(o_label3_data6[0]));
Q_FDP4EP \o_label3_data6_REG[1] ( .CK(clk), .CE(n156), .R(n261), .D(n7), .Q(o_label3_data6[1]));
Q_FDP4EP \o_label3_data6_REG[2] ( .CK(clk), .CE(n156), .R(n261), .D(n8), .Q(o_label3_data6[2]));
Q_FDP4EP \o_label3_data6_REG[3] ( .CK(clk), .CE(n156), .R(n261), .D(n9), .Q(o_label3_data6[3]));
Q_FDP4EP \o_label3_data6_REG[4] ( .CK(clk), .CE(n156), .R(n261), .D(n10), .Q(o_label3_data6[4]));
Q_FDP4EP \o_label3_data6_REG[5] ( .CK(clk), .CE(n156), .R(n261), .D(n11), .Q(o_label3_data6[5]));
Q_FDP4EP \o_label3_data6_REG[6] ( .CK(clk), .CE(n156), .R(n261), .D(n12), .Q(o_label3_data6[6]));
Q_FDP4EP \o_label3_data6_REG[7] ( .CK(clk), .CE(n156), .R(n261), .D(n13), .Q(o_label3_data6[7]));
Q_FDP4EP \o_label3_data6_REG[8] ( .CK(clk), .CE(n156), .R(n261), .D(n14), .Q(o_label3_data6[8]));
Q_FDP4EP \o_label3_data6_REG[9] ( .CK(clk), .CE(n156), .R(n261), .D(n15), .Q(o_label3_data6[9]));
Q_FDP4EP \o_label3_data6_REG[10] ( .CK(clk), .CE(n156), .R(n261), .D(n16), .Q(o_label3_data6[10]));
Q_FDP4EP \o_label3_data6_REG[11] ( .CK(clk), .CE(n156), .R(n261), .D(n17), .Q(o_label3_data6[11]));
Q_FDP4EP \o_label3_data6_REG[12] ( .CK(clk), .CE(n156), .R(n261), .D(n18), .Q(o_label3_data6[12]));
Q_FDP4EP \o_label3_data6_REG[13] ( .CK(clk), .CE(n156), .R(n261), .D(n19), .Q(o_label3_data6[13]));
Q_FDP4EP \o_label3_data6_REG[14] ( .CK(clk), .CE(n156), .R(n261), .D(n20), .Q(o_label3_data6[14]));
Q_FDP4EP \o_label3_data6_REG[15] ( .CK(clk), .CE(n156), .R(n261), .D(n21), .Q(o_label3_data6[15]));
Q_FDP4EP \o_label3_data6_REG[16] ( .CK(clk), .CE(n156), .R(n261), .D(n22), .Q(o_label3_data6[16]));
Q_FDP4EP \o_label3_data6_REG[17] ( .CK(clk), .CE(n156), .R(n261), .D(n23), .Q(o_label3_data6[17]));
Q_FDP4EP \o_label3_data6_REG[18] ( .CK(clk), .CE(n156), .R(n261), .D(n24), .Q(o_label3_data6[18]));
Q_FDP4EP \o_label3_data6_REG[19] ( .CK(clk), .CE(n156), .R(n261), .D(n25), .Q(o_label3_data6[19]));
Q_FDP4EP \o_label3_data6_REG[20] ( .CK(clk), .CE(n156), .R(n261), .D(n26), .Q(o_label3_data6[20]));
Q_FDP4EP \o_label3_data6_REG[21] ( .CK(clk), .CE(n156), .R(n261), .D(n27), .Q(o_label3_data6[21]));
Q_FDP4EP \o_label3_data6_REG[22] ( .CK(clk), .CE(n156), .R(n261), .D(n28), .Q(o_label3_data6[22]));
Q_FDP4EP \o_label3_data6_REG[23] ( .CK(clk), .CE(n156), .R(n261), .D(n29), .Q(o_label3_data6[23]));
Q_FDP4EP \o_label3_data6_REG[24] ( .CK(clk), .CE(n156), .R(n261), .D(n30), .Q(o_label3_data6[24]));
Q_FDP4EP \o_label3_data6_REG[25] ( .CK(clk), .CE(n156), .R(n261), .D(n31), .Q(o_label3_data6[25]));
Q_FDP4EP \o_label3_data6_REG[26] ( .CK(clk), .CE(n156), .R(n261), .D(n32), .Q(o_label3_data6[26]));
Q_FDP4EP \o_label3_data6_REG[27] ( .CK(clk), .CE(n156), .R(n261), .D(n33), .Q(o_label3_data6[27]));
Q_FDP4EP \o_label3_data6_REG[28] ( .CK(clk), .CE(n156), .R(n261), .D(n34), .Q(o_label3_data6[28]));
Q_FDP4EP \o_label3_data6_REG[29] ( .CK(clk), .CE(n156), .R(n261), .D(n35), .Q(o_label3_data6[29]));
Q_FDP4EP \o_label3_data6_REG[30] ( .CK(clk), .CE(n156), .R(n261), .D(n36), .Q(o_label3_data6[30]));
Q_FDP4EP \o_label3_data6_REG[31] ( .CK(clk), .CE(n156), .R(n261), .D(n37), .Q(o_label3_data6[31]));
Q_FDP4EP \o_label3_data7_REG[0] ( .CK(clk), .CE(n155), .R(n261), .D(n6), .Q(o_label3_data7[0]));
Q_FDP4EP \o_label3_data7_REG[1] ( .CK(clk), .CE(n155), .R(n261), .D(n7), .Q(o_label3_data7[1]));
Q_FDP4EP \o_label3_data7_REG[2] ( .CK(clk), .CE(n155), .R(n261), .D(n8), .Q(o_label3_data7[2]));
Q_FDP4EP \o_label3_data7_REG[3] ( .CK(clk), .CE(n155), .R(n261), .D(n9), .Q(o_label3_data7[3]));
Q_FDP4EP \o_label3_data7_REG[4] ( .CK(clk), .CE(n155), .R(n261), .D(n10), .Q(o_label3_data7[4]));
Q_FDP4EP \o_label3_data7_REG[5] ( .CK(clk), .CE(n155), .R(n261), .D(n11), .Q(o_label3_data7[5]));
Q_FDP4EP \o_label3_data7_REG[6] ( .CK(clk), .CE(n155), .R(n261), .D(n12), .Q(o_label3_data7[6]));
Q_FDP4EP \o_label3_data7_REG[7] ( .CK(clk), .CE(n155), .R(n261), .D(n13), .Q(o_label3_data7[7]));
Q_FDP4EP \o_label3_data7_REG[8] ( .CK(clk), .CE(n155), .R(n261), .D(n14), .Q(o_label3_data7[8]));
Q_FDP4EP \o_label3_data7_REG[9] ( .CK(clk), .CE(n155), .R(n261), .D(n15), .Q(o_label3_data7[9]));
Q_FDP4EP \o_label3_data7_REG[10] ( .CK(clk), .CE(n155), .R(n261), .D(n16), .Q(o_label3_data7[10]));
Q_FDP4EP \o_label3_data7_REG[11] ( .CK(clk), .CE(n155), .R(n261), .D(n17), .Q(o_label3_data7[11]));
Q_FDP4EP \o_label3_data7_REG[12] ( .CK(clk), .CE(n155), .R(n261), .D(n18), .Q(o_label3_data7[12]));
Q_FDP4EP \o_label3_data7_REG[13] ( .CK(clk), .CE(n155), .R(n261), .D(n19), .Q(o_label3_data7[13]));
Q_FDP4EP \o_label3_data7_REG[14] ( .CK(clk), .CE(n155), .R(n261), .D(n20), .Q(o_label3_data7[14]));
Q_FDP4EP \o_label3_data7_REG[15] ( .CK(clk), .CE(n155), .R(n261), .D(n21), .Q(o_label3_data7[15]));
Q_FDP4EP \o_label3_data7_REG[16] ( .CK(clk), .CE(n155), .R(n261), .D(n22), .Q(o_label3_data7[16]));
Q_FDP4EP \o_label3_data7_REG[17] ( .CK(clk), .CE(n155), .R(n261), .D(n23), .Q(o_label3_data7[17]));
Q_FDP4EP \o_label3_data7_REG[18] ( .CK(clk), .CE(n155), .R(n261), .D(n24), .Q(o_label3_data7[18]));
Q_FDP4EP \o_label3_data7_REG[19] ( .CK(clk), .CE(n155), .R(n261), .D(n25), .Q(o_label3_data7[19]));
Q_FDP4EP \o_label3_data7_REG[20] ( .CK(clk), .CE(n155), .R(n261), .D(n26), .Q(o_label3_data7[20]));
Q_FDP4EP \o_label3_data7_REG[21] ( .CK(clk), .CE(n155), .R(n261), .D(n27), .Q(o_label3_data7[21]));
Q_FDP4EP \o_label3_data7_REG[22] ( .CK(clk), .CE(n155), .R(n261), .D(n28), .Q(o_label3_data7[22]));
Q_FDP4EP \o_label3_data7_REG[23] ( .CK(clk), .CE(n155), .R(n261), .D(n29), .Q(o_label3_data7[23]));
Q_FDP4EP \o_label3_data7_REG[24] ( .CK(clk), .CE(n155), .R(n261), .D(n30), .Q(o_label3_data7[24]));
Q_FDP4EP \o_label3_data7_REG[25] ( .CK(clk), .CE(n155), .R(n261), .D(n31), .Q(o_label3_data7[25]));
Q_FDP4EP \o_label3_data7_REG[26] ( .CK(clk), .CE(n155), .R(n261), .D(n32), .Q(o_label3_data7[26]));
Q_FDP4EP \o_label3_data7_REG[27] ( .CK(clk), .CE(n155), .R(n261), .D(n33), .Q(o_label3_data7[27]));
Q_FDP4EP \o_label3_data7_REG[28] ( .CK(clk), .CE(n155), .R(n261), .D(n34), .Q(o_label3_data7[28]));
Q_FDP4EP \o_label3_data7_REG[29] ( .CK(clk), .CE(n155), .R(n261), .D(n35), .Q(o_label3_data7[29]));
Q_FDP4EP \o_label3_data7_REG[30] ( .CK(clk), .CE(n155), .R(n261), .D(n36), .Q(o_label3_data7[30]));
Q_FDP4EP \o_label3_data7_REG[31] ( .CK(clk), .CE(n155), .R(n261), .D(n37), .Q(o_label3_data7[31]));
Q_FDP4EP \o_label3_config_REG[0] ( .CK(clk), .CE(n154), .R(n261), .D(n6), .Q(o_label3_config[0]));
Q_FDP4EP \o_label3_config_REG[1] ( .CK(clk), .CE(n154), .R(n261), .D(n7), .Q(o_label3_config[1]));
Q_FDP4EP \o_label3_config_REG[2] ( .CK(clk), .CE(n154), .R(n261), .D(n8), .Q(o_label3_config[2]));
Q_FDP4EP \o_label3_config_REG[3] ( .CK(clk), .CE(n154), .R(n261), .D(n9), .Q(o_label3_config[3]));
Q_FDP4EP \o_label3_config_REG[4] ( .CK(clk), .CE(n154), .R(n261), .D(n10), .Q(o_label3_config[4]));
Q_FDP4EP \o_label3_config_REG[5] ( .CK(clk), .CE(n154), .R(n261), .D(n11), .Q(o_label3_config[5]));
Q_FDP4EP \o_label3_config_REG[6] ( .CK(clk), .CE(n154), .R(n261), .D(n12), .Q(o_label3_config[6]));
Q_FDP4EP \o_label3_config_REG[7] ( .CK(clk), .CE(n154), .R(n261), .D(n13), .Q(o_label3_config[7]));
Q_FDP4EP \o_label3_config_REG[9] ( .CK(clk), .CE(n154), .R(n261), .D(n31), .Q(o_label3_config[9]));
Q_FDP4EP \o_label3_config_REG[10] ( .CK(clk), .CE(n154), .R(n261), .D(n32), .Q(o_label3_config[10]));
Q_FDP4EP \o_label3_config_REG[11] ( .CK(clk), .CE(n154), .R(n261), .D(n33), .Q(o_label3_config[11]));
Q_FDP4EP \o_label3_config_REG[12] ( .CK(clk), .CE(n154), .R(n261), .D(n34), .Q(o_label3_config[12]));
Q_FDP4EP \o_label3_config_REG[13] ( .CK(clk), .CE(n154), .R(n261), .D(n35), .Q(o_label3_config[13]));
Q_FDP4EP \o_label3_config_REG[14] ( .CK(clk), .CE(n154), .R(n261), .D(n36), .Q(o_label3_config[14]));
Q_FDP4EP \o_label3_config_REG[15] ( .CK(clk), .CE(n154), .R(n261), .D(n37), .Q(o_label3_config[15]));
Q_FDP4EP \o_label2_data0_REG[0] ( .CK(clk), .CE(n153), .R(n261), .D(n6), .Q(o_label2_data0[0]));
Q_FDP4EP \o_label2_data0_REG[1] ( .CK(clk), .CE(n153), .R(n261), .D(n7), .Q(o_label2_data0[1]));
Q_FDP4EP \o_label2_data0_REG[2] ( .CK(clk), .CE(n153), .R(n261), .D(n8), .Q(o_label2_data0[2]));
Q_FDP4EP \o_label2_data0_REG[3] ( .CK(clk), .CE(n153), .R(n261), .D(n9), .Q(o_label2_data0[3]));
Q_FDP4EP \o_label2_data0_REG[4] ( .CK(clk), .CE(n153), .R(n261), .D(n10), .Q(o_label2_data0[4]));
Q_FDP4EP \o_label2_data0_REG[5] ( .CK(clk), .CE(n153), .R(n261), .D(n11), .Q(o_label2_data0[5]));
Q_FDP4EP \o_label2_data0_REG[6] ( .CK(clk), .CE(n153), .R(n261), .D(n12), .Q(o_label2_data0[6]));
Q_FDP4EP \o_label2_data0_REG[7] ( .CK(clk), .CE(n153), .R(n261), .D(n13), .Q(o_label2_data0[7]));
Q_FDP4EP \o_label2_data0_REG[8] ( .CK(clk), .CE(n153), .R(n261), .D(n14), .Q(o_label2_data0[8]));
Q_FDP4EP \o_label2_data0_REG[9] ( .CK(clk), .CE(n153), .R(n261), .D(n15), .Q(o_label2_data0[9]));
Q_FDP4EP \o_label2_data0_REG[10] ( .CK(clk), .CE(n153), .R(n261), .D(n16), .Q(o_label2_data0[10]));
Q_FDP4EP \o_label2_data0_REG[11] ( .CK(clk), .CE(n153), .R(n261), .D(n17), .Q(o_label2_data0[11]));
Q_FDP4EP \o_label2_data0_REG[12] ( .CK(clk), .CE(n153), .R(n261), .D(n18), .Q(o_label2_data0[12]));
Q_FDP4EP \o_label2_data0_REG[13] ( .CK(clk), .CE(n153), .R(n261), .D(n19), .Q(o_label2_data0[13]));
Q_FDP4EP \o_label2_data0_REG[14] ( .CK(clk), .CE(n153), .R(n261), .D(n20), .Q(o_label2_data0[14]));
Q_FDP4EP \o_label2_data0_REG[15] ( .CK(clk), .CE(n153), .R(n261), .D(n21), .Q(o_label2_data0[15]));
Q_FDP4EP \o_label2_data0_REG[16] ( .CK(clk), .CE(n153), .R(n261), .D(n22), .Q(o_label2_data0[16]));
Q_FDP4EP \o_label2_data0_REG[17] ( .CK(clk), .CE(n153), .R(n261), .D(n23), .Q(o_label2_data0[17]));
Q_FDP4EP \o_label2_data0_REG[18] ( .CK(clk), .CE(n153), .R(n261), .D(n24), .Q(o_label2_data0[18]));
Q_FDP4EP \o_label2_data0_REG[19] ( .CK(clk), .CE(n153), .R(n261), .D(n25), .Q(o_label2_data0[19]));
Q_FDP4EP \o_label2_data0_REG[20] ( .CK(clk), .CE(n153), .R(n261), .D(n26), .Q(o_label2_data0[20]));
Q_FDP4EP \o_label2_data0_REG[21] ( .CK(clk), .CE(n153), .R(n261), .D(n27), .Q(o_label2_data0[21]));
Q_FDP4EP \o_label2_data0_REG[22] ( .CK(clk), .CE(n153), .R(n261), .D(n28), .Q(o_label2_data0[22]));
Q_FDP4EP \o_label2_data0_REG[23] ( .CK(clk), .CE(n153), .R(n261), .D(n29), .Q(o_label2_data0[23]));
Q_FDP4EP \o_label2_data0_REG[24] ( .CK(clk), .CE(n153), .R(n261), .D(n30), .Q(o_label2_data0[24]));
Q_FDP4EP \o_label2_data0_REG[25] ( .CK(clk), .CE(n153), .R(n261), .D(n31), .Q(o_label2_data0[25]));
Q_FDP4EP \o_label2_data0_REG[26] ( .CK(clk), .CE(n153), .R(n261), .D(n32), .Q(o_label2_data0[26]));
Q_FDP4EP \o_label2_data0_REG[27] ( .CK(clk), .CE(n153), .R(n261), .D(n33), .Q(o_label2_data0[27]));
Q_FDP4EP \o_label2_data0_REG[28] ( .CK(clk), .CE(n153), .R(n261), .D(n34), .Q(o_label2_data0[28]));
Q_FDP4EP \o_label2_data0_REG[29] ( .CK(clk), .CE(n153), .R(n261), .D(n35), .Q(o_label2_data0[29]));
Q_FDP4EP \o_label2_data0_REG[30] ( .CK(clk), .CE(n153), .R(n261), .D(n36), .Q(o_label2_data0[30]));
Q_FDP4EP \o_label2_data0_REG[31] ( .CK(clk), .CE(n153), .R(n261), .D(n37), .Q(o_label2_data0[31]));
Q_FDP4EP \o_label2_data1_REG[0] ( .CK(clk), .CE(n152), .R(n261), .D(n6), .Q(o_label2_data1[0]));
Q_FDP4EP \o_label2_data1_REG[1] ( .CK(clk), .CE(n152), .R(n261), .D(n7), .Q(o_label2_data1[1]));
Q_FDP4EP \o_label2_data1_REG[2] ( .CK(clk), .CE(n152), .R(n261), .D(n8), .Q(o_label2_data1[2]));
Q_FDP4EP \o_label2_data1_REG[3] ( .CK(clk), .CE(n152), .R(n261), .D(n9), .Q(o_label2_data1[3]));
Q_FDP4EP \o_label2_data1_REG[4] ( .CK(clk), .CE(n152), .R(n261), .D(n10), .Q(o_label2_data1[4]));
Q_FDP4EP \o_label2_data1_REG[5] ( .CK(clk), .CE(n152), .R(n261), .D(n11), .Q(o_label2_data1[5]));
Q_FDP4EP \o_label2_data1_REG[6] ( .CK(clk), .CE(n152), .R(n261), .D(n12), .Q(o_label2_data1[6]));
Q_FDP4EP \o_label2_data1_REG[7] ( .CK(clk), .CE(n152), .R(n261), .D(n13), .Q(o_label2_data1[7]));
Q_FDP4EP \o_label2_data1_REG[8] ( .CK(clk), .CE(n152), .R(n261), .D(n14), .Q(o_label2_data1[8]));
Q_FDP4EP \o_label2_data1_REG[9] ( .CK(clk), .CE(n152), .R(n261), .D(n15), .Q(o_label2_data1[9]));
Q_FDP4EP \o_label2_data1_REG[10] ( .CK(clk), .CE(n152), .R(n261), .D(n16), .Q(o_label2_data1[10]));
Q_FDP4EP \o_label2_data1_REG[11] ( .CK(clk), .CE(n152), .R(n261), .D(n17), .Q(o_label2_data1[11]));
Q_FDP4EP \o_label2_data1_REG[12] ( .CK(clk), .CE(n152), .R(n261), .D(n18), .Q(o_label2_data1[12]));
Q_FDP4EP \o_label2_data1_REG[13] ( .CK(clk), .CE(n152), .R(n261), .D(n19), .Q(o_label2_data1[13]));
Q_FDP4EP \o_label2_data1_REG[14] ( .CK(clk), .CE(n152), .R(n261), .D(n20), .Q(o_label2_data1[14]));
Q_FDP4EP \o_label2_data1_REG[15] ( .CK(clk), .CE(n152), .R(n261), .D(n21), .Q(o_label2_data1[15]));
Q_FDP4EP \o_label2_data1_REG[16] ( .CK(clk), .CE(n152), .R(n261), .D(n22), .Q(o_label2_data1[16]));
Q_FDP4EP \o_label2_data1_REG[17] ( .CK(clk), .CE(n152), .R(n261), .D(n23), .Q(o_label2_data1[17]));
Q_FDP4EP \o_label2_data1_REG[18] ( .CK(clk), .CE(n152), .R(n261), .D(n24), .Q(o_label2_data1[18]));
Q_FDP4EP \o_label2_data1_REG[19] ( .CK(clk), .CE(n152), .R(n261), .D(n25), .Q(o_label2_data1[19]));
Q_FDP4EP \o_label2_data1_REG[20] ( .CK(clk), .CE(n152), .R(n261), .D(n26), .Q(o_label2_data1[20]));
Q_FDP4EP \o_label2_data1_REG[21] ( .CK(clk), .CE(n152), .R(n261), .D(n27), .Q(o_label2_data1[21]));
Q_FDP4EP \o_label2_data1_REG[22] ( .CK(clk), .CE(n152), .R(n261), .D(n28), .Q(o_label2_data1[22]));
Q_FDP4EP \o_label2_data1_REG[23] ( .CK(clk), .CE(n152), .R(n261), .D(n29), .Q(o_label2_data1[23]));
Q_FDP4EP \o_label2_data1_REG[24] ( .CK(clk), .CE(n152), .R(n261), .D(n30), .Q(o_label2_data1[24]));
Q_FDP4EP \o_label2_data1_REG[25] ( .CK(clk), .CE(n152), .R(n261), .D(n31), .Q(o_label2_data1[25]));
Q_FDP4EP \o_label2_data1_REG[26] ( .CK(clk), .CE(n152), .R(n261), .D(n32), .Q(o_label2_data1[26]));
Q_FDP4EP \o_label2_data1_REG[27] ( .CK(clk), .CE(n152), .R(n261), .D(n33), .Q(o_label2_data1[27]));
Q_FDP4EP \o_label2_data1_REG[28] ( .CK(clk), .CE(n152), .R(n261), .D(n34), .Q(o_label2_data1[28]));
Q_FDP4EP \o_label2_data1_REG[29] ( .CK(clk), .CE(n152), .R(n261), .D(n35), .Q(o_label2_data1[29]));
Q_FDP4EP \o_label2_data1_REG[30] ( .CK(clk), .CE(n152), .R(n261), .D(n36), .Q(o_label2_data1[30]));
Q_FDP4EP \o_label2_data1_REG[31] ( .CK(clk), .CE(n152), .R(n261), .D(n37), .Q(o_label2_data1[31]));
Q_FDP4EP \o_label2_data2_REG[0] ( .CK(clk), .CE(n151), .R(n261), .D(n6), .Q(o_label2_data2[0]));
Q_FDP4EP \o_label2_data2_REG[1] ( .CK(clk), .CE(n151), .R(n261), .D(n7), .Q(o_label2_data2[1]));
Q_FDP4EP \o_label2_data2_REG[2] ( .CK(clk), .CE(n151), .R(n261), .D(n8), .Q(o_label2_data2[2]));
Q_FDP4EP \o_label2_data2_REG[3] ( .CK(clk), .CE(n151), .R(n261), .D(n9), .Q(o_label2_data2[3]));
Q_FDP4EP \o_label2_data2_REG[4] ( .CK(clk), .CE(n151), .R(n261), .D(n10), .Q(o_label2_data2[4]));
Q_FDP4EP \o_label2_data2_REG[5] ( .CK(clk), .CE(n151), .R(n261), .D(n11), .Q(o_label2_data2[5]));
Q_FDP4EP \o_label2_data2_REG[6] ( .CK(clk), .CE(n151), .R(n261), .D(n12), .Q(o_label2_data2[6]));
Q_FDP4EP \o_label2_data2_REG[7] ( .CK(clk), .CE(n151), .R(n261), .D(n13), .Q(o_label2_data2[7]));
Q_FDP4EP \o_label2_data2_REG[8] ( .CK(clk), .CE(n151), .R(n261), .D(n14), .Q(o_label2_data2[8]));
Q_FDP4EP \o_label2_data2_REG[9] ( .CK(clk), .CE(n151), .R(n261), .D(n15), .Q(o_label2_data2[9]));
Q_FDP4EP \o_label2_data2_REG[10] ( .CK(clk), .CE(n151), .R(n261), .D(n16), .Q(o_label2_data2[10]));
Q_FDP4EP \o_label2_data2_REG[11] ( .CK(clk), .CE(n151), .R(n261), .D(n17), .Q(o_label2_data2[11]));
Q_FDP4EP \o_label2_data2_REG[12] ( .CK(clk), .CE(n151), .R(n261), .D(n18), .Q(o_label2_data2[12]));
Q_FDP4EP \o_label2_data2_REG[13] ( .CK(clk), .CE(n151), .R(n261), .D(n19), .Q(o_label2_data2[13]));
Q_FDP4EP \o_label2_data2_REG[14] ( .CK(clk), .CE(n151), .R(n261), .D(n20), .Q(o_label2_data2[14]));
Q_FDP4EP \o_label2_data2_REG[15] ( .CK(clk), .CE(n151), .R(n261), .D(n21), .Q(o_label2_data2[15]));
Q_FDP4EP \o_label2_data2_REG[16] ( .CK(clk), .CE(n151), .R(n261), .D(n22), .Q(o_label2_data2[16]));
Q_FDP4EP \o_label2_data2_REG[17] ( .CK(clk), .CE(n151), .R(n261), .D(n23), .Q(o_label2_data2[17]));
Q_FDP4EP \o_label2_data2_REG[18] ( .CK(clk), .CE(n151), .R(n261), .D(n24), .Q(o_label2_data2[18]));
Q_FDP4EP \o_label2_data2_REG[19] ( .CK(clk), .CE(n151), .R(n261), .D(n25), .Q(o_label2_data2[19]));
Q_FDP4EP \o_label2_data2_REG[20] ( .CK(clk), .CE(n151), .R(n261), .D(n26), .Q(o_label2_data2[20]));
Q_FDP4EP \o_label2_data2_REG[21] ( .CK(clk), .CE(n151), .R(n261), .D(n27), .Q(o_label2_data2[21]));
Q_FDP4EP \o_label2_data2_REG[22] ( .CK(clk), .CE(n151), .R(n261), .D(n28), .Q(o_label2_data2[22]));
Q_FDP4EP \o_label2_data2_REG[23] ( .CK(clk), .CE(n151), .R(n261), .D(n29), .Q(o_label2_data2[23]));
Q_FDP4EP \o_label2_data2_REG[24] ( .CK(clk), .CE(n151), .R(n261), .D(n30), .Q(o_label2_data2[24]));
Q_FDP4EP \o_label2_data2_REG[25] ( .CK(clk), .CE(n151), .R(n261), .D(n31), .Q(o_label2_data2[25]));
Q_FDP4EP \o_label2_data2_REG[26] ( .CK(clk), .CE(n151), .R(n261), .D(n32), .Q(o_label2_data2[26]));
Q_FDP4EP \o_label2_data2_REG[27] ( .CK(clk), .CE(n151), .R(n261), .D(n33), .Q(o_label2_data2[27]));
Q_FDP4EP \o_label2_data2_REG[28] ( .CK(clk), .CE(n151), .R(n261), .D(n34), .Q(o_label2_data2[28]));
Q_FDP4EP \o_label2_data2_REG[29] ( .CK(clk), .CE(n151), .R(n261), .D(n35), .Q(o_label2_data2[29]));
Q_FDP4EP \o_label2_data2_REG[30] ( .CK(clk), .CE(n151), .R(n261), .D(n36), .Q(o_label2_data2[30]));
Q_FDP4EP \o_label2_data2_REG[31] ( .CK(clk), .CE(n151), .R(n261), .D(n37), .Q(o_label2_data2[31]));
Q_FDP4EP \o_label2_data3_REG[0] ( .CK(clk), .CE(n150), .R(n261), .D(n6), .Q(o_label2_data3[0]));
Q_FDP4EP \o_label2_data3_REG[1] ( .CK(clk), .CE(n150), .R(n261), .D(n7), .Q(o_label2_data3[1]));
Q_FDP4EP \o_label2_data3_REG[2] ( .CK(clk), .CE(n150), .R(n261), .D(n8), .Q(o_label2_data3[2]));
Q_FDP4EP \o_label2_data3_REG[3] ( .CK(clk), .CE(n150), .R(n261), .D(n9), .Q(o_label2_data3[3]));
Q_FDP4EP \o_label2_data3_REG[4] ( .CK(clk), .CE(n150), .R(n261), .D(n10), .Q(o_label2_data3[4]));
Q_FDP4EP \o_label2_data3_REG[5] ( .CK(clk), .CE(n150), .R(n261), .D(n11), .Q(o_label2_data3[5]));
Q_FDP4EP \o_label2_data3_REG[6] ( .CK(clk), .CE(n150), .R(n261), .D(n12), .Q(o_label2_data3[6]));
Q_FDP4EP \o_label2_data3_REG[7] ( .CK(clk), .CE(n150), .R(n261), .D(n13), .Q(o_label2_data3[7]));
Q_FDP4EP \o_label2_data3_REG[8] ( .CK(clk), .CE(n150), .R(n261), .D(n14), .Q(o_label2_data3[8]));
Q_FDP4EP \o_label2_data3_REG[9] ( .CK(clk), .CE(n150), .R(n261), .D(n15), .Q(o_label2_data3[9]));
Q_FDP4EP \o_label2_data3_REG[10] ( .CK(clk), .CE(n150), .R(n261), .D(n16), .Q(o_label2_data3[10]));
Q_FDP4EP \o_label2_data3_REG[11] ( .CK(clk), .CE(n150), .R(n261), .D(n17), .Q(o_label2_data3[11]));
Q_FDP4EP \o_label2_data3_REG[12] ( .CK(clk), .CE(n150), .R(n261), .D(n18), .Q(o_label2_data3[12]));
Q_FDP4EP \o_label2_data3_REG[13] ( .CK(clk), .CE(n150), .R(n261), .D(n19), .Q(o_label2_data3[13]));
Q_FDP4EP \o_label2_data3_REG[14] ( .CK(clk), .CE(n150), .R(n261), .D(n20), .Q(o_label2_data3[14]));
Q_FDP4EP \o_label2_data3_REG[15] ( .CK(clk), .CE(n150), .R(n261), .D(n21), .Q(o_label2_data3[15]));
Q_FDP4EP \o_label2_data3_REG[16] ( .CK(clk), .CE(n150), .R(n261), .D(n22), .Q(o_label2_data3[16]));
Q_FDP4EP \o_label2_data3_REG[17] ( .CK(clk), .CE(n150), .R(n261), .D(n23), .Q(o_label2_data3[17]));
Q_FDP4EP \o_label2_data3_REG[18] ( .CK(clk), .CE(n150), .R(n261), .D(n24), .Q(o_label2_data3[18]));
Q_FDP4EP \o_label2_data3_REG[19] ( .CK(clk), .CE(n150), .R(n261), .D(n25), .Q(o_label2_data3[19]));
Q_FDP4EP \o_label2_data3_REG[20] ( .CK(clk), .CE(n150), .R(n261), .D(n26), .Q(o_label2_data3[20]));
Q_FDP4EP \o_label2_data3_REG[21] ( .CK(clk), .CE(n150), .R(n261), .D(n27), .Q(o_label2_data3[21]));
Q_FDP4EP \o_label2_data3_REG[22] ( .CK(clk), .CE(n150), .R(n261), .D(n28), .Q(o_label2_data3[22]));
Q_FDP4EP \o_label2_data3_REG[23] ( .CK(clk), .CE(n150), .R(n261), .D(n29), .Q(o_label2_data3[23]));
Q_FDP4EP \o_label2_data3_REG[24] ( .CK(clk), .CE(n150), .R(n261), .D(n30), .Q(o_label2_data3[24]));
Q_FDP4EP \o_label2_data3_REG[25] ( .CK(clk), .CE(n150), .R(n261), .D(n31), .Q(o_label2_data3[25]));
Q_FDP4EP \o_label2_data3_REG[26] ( .CK(clk), .CE(n150), .R(n261), .D(n32), .Q(o_label2_data3[26]));
Q_FDP4EP \o_label2_data3_REG[27] ( .CK(clk), .CE(n150), .R(n261), .D(n33), .Q(o_label2_data3[27]));
Q_FDP4EP \o_label2_data3_REG[28] ( .CK(clk), .CE(n150), .R(n261), .D(n34), .Q(o_label2_data3[28]));
Q_FDP4EP \o_label2_data3_REG[29] ( .CK(clk), .CE(n150), .R(n261), .D(n35), .Q(o_label2_data3[29]));
Q_FDP4EP \o_label2_data3_REG[30] ( .CK(clk), .CE(n150), .R(n261), .D(n36), .Q(o_label2_data3[30]));
Q_FDP4EP \o_label2_data3_REG[31] ( .CK(clk), .CE(n150), .R(n261), .D(n37), .Q(o_label2_data3[31]));
Q_FDP4EP \o_label2_data4_REG[0] ( .CK(clk), .CE(n149), .R(n261), .D(n6), .Q(o_label2_data4[0]));
Q_FDP4EP \o_label2_data4_REG[1] ( .CK(clk), .CE(n149), .R(n261), .D(n7), .Q(o_label2_data4[1]));
Q_FDP4EP \o_label2_data4_REG[2] ( .CK(clk), .CE(n149), .R(n261), .D(n8), .Q(o_label2_data4[2]));
Q_FDP4EP \o_label2_data4_REG[3] ( .CK(clk), .CE(n149), .R(n261), .D(n9), .Q(o_label2_data4[3]));
Q_FDP4EP \o_label2_data4_REG[4] ( .CK(clk), .CE(n149), .R(n261), .D(n10), .Q(o_label2_data4[4]));
Q_FDP4EP \o_label2_data4_REG[5] ( .CK(clk), .CE(n149), .R(n261), .D(n11), .Q(o_label2_data4[5]));
Q_FDP4EP \o_label2_data4_REG[6] ( .CK(clk), .CE(n149), .R(n261), .D(n12), .Q(o_label2_data4[6]));
Q_FDP4EP \o_label2_data4_REG[7] ( .CK(clk), .CE(n149), .R(n261), .D(n13), .Q(o_label2_data4[7]));
Q_FDP4EP \o_label2_data4_REG[8] ( .CK(clk), .CE(n149), .R(n261), .D(n14), .Q(o_label2_data4[8]));
Q_FDP4EP \o_label2_data4_REG[9] ( .CK(clk), .CE(n149), .R(n261), .D(n15), .Q(o_label2_data4[9]));
Q_FDP4EP \o_label2_data4_REG[10] ( .CK(clk), .CE(n149), .R(n261), .D(n16), .Q(o_label2_data4[10]));
Q_FDP4EP \o_label2_data4_REG[11] ( .CK(clk), .CE(n149), .R(n261), .D(n17), .Q(o_label2_data4[11]));
Q_FDP4EP \o_label2_data4_REG[12] ( .CK(clk), .CE(n149), .R(n261), .D(n18), .Q(o_label2_data4[12]));
Q_FDP4EP \o_label2_data4_REG[13] ( .CK(clk), .CE(n149), .R(n261), .D(n19), .Q(o_label2_data4[13]));
Q_FDP4EP \o_label2_data4_REG[14] ( .CK(clk), .CE(n149), .R(n261), .D(n20), .Q(o_label2_data4[14]));
Q_FDP4EP \o_label2_data4_REG[15] ( .CK(clk), .CE(n149), .R(n261), .D(n21), .Q(o_label2_data4[15]));
Q_FDP4EP \o_label2_data4_REG[16] ( .CK(clk), .CE(n149), .R(n261), .D(n22), .Q(o_label2_data4[16]));
Q_FDP4EP \o_label2_data4_REG[17] ( .CK(clk), .CE(n149), .R(n261), .D(n23), .Q(o_label2_data4[17]));
Q_FDP4EP \o_label2_data4_REG[18] ( .CK(clk), .CE(n149), .R(n261), .D(n24), .Q(o_label2_data4[18]));
Q_FDP4EP \o_label2_data4_REG[19] ( .CK(clk), .CE(n149), .R(n261), .D(n25), .Q(o_label2_data4[19]));
Q_FDP4EP \o_label2_data4_REG[20] ( .CK(clk), .CE(n149), .R(n261), .D(n26), .Q(o_label2_data4[20]));
Q_FDP4EP \o_label2_data4_REG[21] ( .CK(clk), .CE(n149), .R(n261), .D(n27), .Q(o_label2_data4[21]));
Q_FDP4EP \o_label2_data4_REG[22] ( .CK(clk), .CE(n149), .R(n261), .D(n28), .Q(o_label2_data4[22]));
Q_FDP4EP \o_label2_data4_REG[23] ( .CK(clk), .CE(n149), .R(n261), .D(n29), .Q(o_label2_data4[23]));
Q_FDP4EP \o_label2_data4_REG[24] ( .CK(clk), .CE(n149), .R(n261), .D(n30), .Q(o_label2_data4[24]));
Q_FDP4EP \o_label2_data4_REG[25] ( .CK(clk), .CE(n149), .R(n261), .D(n31), .Q(o_label2_data4[25]));
Q_FDP4EP \o_label2_data4_REG[26] ( .CK(clk), .CE(n149), .R(n261), .D(n32), .Q(o_label2_data4[26]));
Q_FDP4EP \o_label2_data4_REG[27] ( .CK(clk), .CE(n149), .R(n261), .D(n33), .Q(o_label2_data4[27]));
Q_FDP4EP \o_label2_data4_REG[28] ( .CK(clk), .CE(n149), .R(n261), .D(n34), .Q(o_label2_data4[28]));
Q_FDP4EP \o_label2_data4_REG[29] ( .CK(clk), .CE(n149), .R(n261), .D(n35), .Q(o_label2_data4[29]));
Q_FDP4EP \o_label2_data4_REG[30] ( .CK(clk), .CE(n149), .R(n261), .D(n36), .Q(o_label2_data4[30]));
Q_FDP4EP \o_label2_data4_REG[31] ( .CK(clk), .CE(n149), .R(n261), .D(n37), .Q(o_label2_data4[31]));
Q_FDP4EP \o_label2_data5_REG[0] ( .CK(clk), .CE(n148), .R(n261), .D(n6), .Q(o_label2_data5[0]));
Q_FDP4EP \o_label2_data5_REG[1] ( .CK(clk), .CE(n148), .R(n261), .D(n7), .Q(o_label2_data5[1]));
Q_FDP4EP \o_label2_data5_REG[2] ( .CK(clk), .CE(n148), .R(n261), .D(n8), .Q(o_label2_data5[2]));
Q_FDP4EP \o_label2_data5_REG[3] ( .CK(clk), .CE(n148), .R(n261), .D(n9), .Q(o_label2_data5[3]));
Q_FDP4EP \o_label2_data5_REG[4] ( .CK(clk), .CE(n148), .R(n261), .D(n10), .Q(o_label2_data5[4]));
Q_FDP4EP \o_label2_data5_REG[5] ( .CK(clk), .CE(n148), .R(n261), .D(n11), .Q(o_label2_data5[5]));
Q_FDP4EP \o_label2_data5_REG[6] ( .CK(clk), .CE(n148), .R(n261), .D(n12), .Q(o_label2_data5[6]));
Q_FDP4EP \o_label2_data5_REG[7] ( .CK(clk), .CE(n148), .R(n261), .D(n13), .Q(o_label2_data5[7]));
Q_FDP4EP \o_label2_data5_REG[8] ( .CK(clk), .CE(n148), .R(n261), .D(n14), .Q(o_label2_data5[8]));
Q_FDP4EP \o_label2_data5_REG[9] ( .CK(clk), .CE(n148), .R(n261), .D(n15), .Q(o_label2_data5[9]));
Q_FDP4EP \o_label2_data5_REG[10] ( .CK(clk), .CE(n148), .R(n261), .D(n16), .Q(o_label2_data5[10]));
Q_FDP4EP \o_label2_data5_REG[11] ( .CK(clk), .CE(n148), .R(n261), .D(n17), .Q(o_label2_data5[11]));
Q_FDP4EP \o_label2_data5_REG[12] ( .CK(clk), .CE(n148), .R(n261), .D(n18), .Q(o_label2_data5[12]));
Q_FDP4EP \o_label2_data5_REG[13] ( .CK(clk), .CE(n148), .R(n261), .D(n19), .Q(o_label2_data5[13]));
Q_FDP4EP \o_label2_data5_REG[14] ( .CK(clk), .CE(n148), .R(n261), .D(n20), .Q(o_label2_data5[14]));
Q_FDP4EP \o_label2_data5_REG[15] ( .CK(clk), .CE(n148), .R(n261), .D(n21), .Q(o_label2_data5[15]));
Q_FDP4EP \o_label2_data5_REG[16] ( .CK(clk), .CE(n148), .R(n261), .D(n22), .Q(o_label2_data5[16]));
Q_FDP4EP \o_label2_data5_REG[17] ( .CK(clk), .CE(n148), .R(n261), .D(n23), .Q(o_label2_data5[17]));
Q_FDP4EP \o_label2_data5_REG[18] ( .CK(clk), .CE(n148), .R(n261), .D(n24), .Q(o_label2_data5[18]));
Q_FDP4EP \o_label2_data5_REG[19] ( .CK(clk), .CE(n148), .R(n261), .D(n25), .Q(o_label2_data5[19]));
Q_FDP4EP \o_label2_data5_REG[20] ( .CK(clk), .CE(n148), .R(n261), .D(n26), .Q(o_label2_data5[20]));
Q_FDP4EP \o_label2_data5_REG[21] ( .CK(clk), .CE(n148), .R(n261), .D(n27), .Q(o_label2_data5[21]));
Q_FDP4EP \o_label2_data5_REG[22] ( .CK(clk), .CE(n148), .R(n261), .D(n28), .Q(o_label2_data5[22]));
Q_FDP4EP \o_label2_data5_REG[23] ( .CK(clk), .CE(n148), .R(n261), .D(n29), .Q(o_label2_data5[23]));
Q_FDP4EP \o_label2_data5_REG[24] ( .CK(clk), .CE(n148), .R(n261), .D(n30), .Q(o_label2_data5[24]));
Q_FDP4EP \o_label2_data5_REG[25] ( .CK(clk), .CE(n148), .R(n261), .D(n31), .Q(o_label2_data5[25]));
Q_FDP4EP \o_label2_data5_REG[26] ( .CK(clk), .CE(n148), .R(n261), .D(n32), .Q(o_label2_data5[26]));
Q_FDP4EP \o_label2_data5_REG[27] ( .CK(clk), .CE(n148), .R(n261), .D(n33), .Q(o_label2_data5[27]));
Q_FDP4EP \o_label2_data5_REG[28] ( .CK(clk), .CE(n148), .R(n261), .D(n34), .Q(o_label2_data5[28]));
Q_FDP4EP \o_label2_data5_REG[29] ( .CK(clk), .CE(n148), .R(n261), .D(n35), .Q(o_label2_data5[29]));
Q_FDP4EP \o_label2_data5_REG[30] ( .CK(clk), .CE(n148), .R(n261), .D(n36), .Q(o_label2_data5[30]));
Q_FDP4EP \o_label2_data5_REG[31] ( .CK(clk), .CE(n148), .R(n261), .D(n37), .Q(o_label2_data5[31]));
Q_FDP4EP \o_label2_data6_REG[0] ( .CK(clk), .CE(n147), .R(n261), .D(n6), .Q(o_label2_data6[0]));
Q_FDP4EP \o_label2_data6_REG[1] ( .CK(clk), .CE(n147), .R(n261), .D(n7), .Q(o_label2_data6[1]));
Q_FDP4EP \o_label2_data6_REG[2] ( .CK(clk), .CE(n147), .R(n261), .D(n8), .Q(o_label2_data6[2]));
Q_FDP4EP \o_label2_data6_REG[3] ( .CK(clk), .CE(n147), .R(n261), .D(n9), .Q(o_label2_data6[3]));
Q_FDP4EP \o_label2_data6_REG[4] ( .CK(clk), .CE(n147), .R(n261), .D(n10), .Q(o_label2_data6[4]));
Q_FDP4EP \o_label2_data6_REG[5] ( .CK(clk), .CE(n147), .R(n261), .D(n11), .Q(o_label2_data6[5]));
Q_FDP4EP \o_label2_data6_REG[6] ( .CK(clk), .CE(n147), .R(n261), .D(n12), .Q(o_label2_data6[6]));
Q_FDP4EP \o_label2_data6_REG[7] ( .CK(clk), .CE(n147), .R(n261), .D(n13), .Q(o_label2_data6[7]));
Q_FDP4EP \o_label2_data6_REG[8] ( .CK(clk), .CE(n147), .R(n261), .D(n14), .Q(o_label2_data6[8]));
Q_FDP4EP \o_label2_data6_REG[9] ( .CK(clk), .CE(n147), .R(n261), .D(n15), .Q(o_label2_data6[9]));
Q_FDP4EP \o_label2_data6_REG[10] ( .CK(clk), .CE(n147), .R(n261), .D(n16), .Q(o_label2_data6[10]));
Q_FDP4EP \o_label2_data6_REG[11] ( .CK(clk), .CE(n147), .R(n261), .D(n17), .Q(o_label2_data6[11]));
Q_FDP4EP \o_label2_data6_REG[12] ( .CK(clk), .CE(n147), .R(n261), .D(n18), .Q(o_label2_data6[12]));
Q_FDP4EP \o_label2_data6_REG[13] ( .CK(clk), .CE(n147), .R(n261), .D(n19), .Q(o_label2_data6[13]));
Q_FDP4EP \o_label2_data6_REG[14] ( .CK(clk), .CE(n147), .R(n261), .D(n20), .Q(o_label2_data6[14]));
Q_FDP4EP \o_label2_data6_REG[15] ( .CK(clk), .CE(n147), .R(n261), .D(n21), .Q(o_label2_data6[15]));
Q_FDP4EP \o_label2_data6_REG[16] ( .CK(clk), .CE(n147), .R(n261), .D(n22), .Q(o_label2_data6[16]));
Q_FDP4EP \o_label2_data6_REG[17] ( .CK(clk), .CE(n147), .R(n261), .D(n23), .Q(o_label2_data6[17]));
Q_FDP4EP \o_label2_data6_REG[18] ( .CK(clk), .CE(n147), .R(n261), .D(n24), .Q(o_label2_data6[18]));
Q_FDP4EP \o_label2_data6_REG[19] ( .CK(clk), .CE(n147), .R(n261), .D(n25), .Q(o_label2_data6[19]));
Q_FDP4EP \o_label2_data6_REG[20] ( .CK(clk), .CE(n147), .R(n261), .D(n26), .Q(o_label2_data6[20]));
Q_FDP4EP \o_label2_data6_REG[21] ( .CK(clk), .CE(n147), .R(n261), .D(n27), .Q(o_label2_data6[21]));
Q_FDP4EP \o_label2_data6_REG[22] ( .CK(clk), .CE(n147), .R(n261), .D(n28), .Q(o_label2_data6[22]));
Q_FDP4EP \o_label2_data6_REG[23] ( .CK(clk), .CE(n147), .R(n261), .D(n29), .Q(o_label2_data6[23]));
Q_FDP4EP \o_label2_data6_REG[24] ( .CK(clk), .CE(n147), .R(n261), .D(n30), .Q(o_label2_data6[24]));
Q_FDP4EP \o_label2_data6_REG[25] ( .CK(clk), .CE(n147), .R(n261), .D(n31), .Q(o_label2_data6[25]));
Q_FDP4EP \o_label2_data6_REG[26] ( .CK(clk), .CE(n147), .R(n261), .D(n32), .Q(o_label2_data6[26]));
Q_FDP4EP \o_label2_data6_REG[27] ( .CK(clk), .CE(n147), .R(n261), .D(n33), .Q(o_label2_data6[27]));
Q_FDP4EP \o_label2_data6_REG[28] ( .CK(clk), .CE(n147), .R(n261), .D(n34), .Q(o_label2_data6[28]));
Q_FDP4EP \o_label2_data6_REG[29] ( .CK(clk), .CE(n147), .R(n261), .D(n35), .Q(o_label2_data6[29]));
Q_FDP4EP \o_label2_data6_REG[30] ( .CK(clk), .CE(n147), .R(n261), .D(n36), .Q(o_label2_data6[30]));
Q_FDP4EP \o_label2_data6_REG[31] ( .CK(clk), .CE(n147), .R(n261), .D(n37), .Q(o_label2_data6[31]));
Q_FDP4EP \o_label2_data7_REG[0] ( .CK(clk), .CE(n146), .R(n261), .D(n6), .Q(o_label2_data7[0]));
Q_FDP4EP \o_label2_data7_REG[1] ( .CK(clk), .CE(n146), .R(n261), .D(n7), .Q(o_label2_data7[1]));
Q_FDP4EP \o_label2_data7_REG[2] ( .CK(clk), .CE(n146), .R(n261), .D(n8), .Q(o_label2_data7[2]));
Q_FDP4EP \o_label2_data7_REG[3] ( .CK(clk), .CE(n146), .R(n261), .D(n9), .Q(o_label2_data7[3]));
Q_FDP4EP \o_label2_data7_REG[4] ( .CK(clk), .CE(n146), .R(n261), .D(n10), .Q(o_label2_data7[4]));
Q_FDP4EP \o_label2_data7_REG[5] ( .CK(clk), .CE(n146), .R(n261), .D(n11), .Q(o_label2_data7[5]));
Q_FDP4EP \o_label2_data7_REG[6] ( .CK(clk), .CE(n146), .R(n261), .D(n12), .Q(o_label2_data7[6]));
Q_FDP4EP \o_label2_data7_REG[7] ( .CK(clk), .CE(n146), .R(n261), .D(n13), .Q(o_label2_data7[7]));
Q_FDP4EP \o_label2_data7_REG[8] ( .CK(clk), .CE(n146), .R(n261), .D(n14), .Q(o_label2_data7[8]));
Q_FDP4EP \o_label2_data7_REG[9] ( .CK(clk), .CE(n146), .R(n261), .D(n15), .Q(o_label2_data7[9]));
Q_FDP4EP \o_label2_data7_REG[10] ( .CK(clk), .CE(n146), .R(n261), .D(n16), .Q(o_label2_data7[10]));
Q_FDP4EP \o_label2_data7_REG[11] ( .CK(clk), .CE(n146), .R(n261), .D(n17), .Q(o_label2_data7[11]));
Q_FDP4EP \o_label2_data7_REG[12] ( .CK(clk), .CE(n146), .R(n261), .D(n18), .Q(o_label2_data7[12]));
Q_FDP4EP \o_label2_data7_REG[13] ( .CK(clk), .CE(n146), .R(n261), .D(n19), .Q(o_label2_data7[13]));
Q_FDP4EP \o_label2_data7_REG[14] ( .CK(clk), .CE(n146), .R(n261), .D(n20), .Q(o_label2_data7[14]));
Q_FDP4EP \o_label2_data7_REG[15] ( .CK(clk), .CE(n146), .R(n261), .D(n21), .Q(o_label2_data7[15]));
Q_FDP4EP \o_label2_data7_REG[16] ( .CK(clk), .CE(n146), .R(n261), .D(n22), .Q(o_label2_data7[16]));
Q_FDP4EP \o_label2_data7_REG[17] ( .CK(clk), .CE(n146), .R(n261), .D(n23), .Q(o_label2_data7[17]));
Q_FDP4EP \o_label2_data7_REG[18] ( .CK(clk), .CE(n146), .R(n261), .D(n24), .Q(o_label2_data7[18]));
Q_FDP4EP \o_label2_data7_REG[19] ( .CK(clk), .CE(n146), .R(n261), .D(n25), .Q(o_label2_data7[19]));
Q_FDP4EP \o_label2_data7_REG[20] ( .CK(clk), .CE(n146), .R(n261), .D(n26), .Q(o_label2_data7[20]));
Q_FDP4EP \o_label2_data7_REG[21] ( .CK(clk), .CE(n146), .R(n261), .D(n27), .Q(o_label2_data7[21]));
Q_FDP4EP \o_label2_data7_REG[22] ( .CK(clk), .CE(n146), .R(n261), .D(n28), .Q(o_label2_data7[22]));
Q_FDP4EP \o_label2_data7_REG[23] ( .CK(clk), .CE(n146), .R(n261), .D(n29), .Q(o_label2_data7[23]));
Q_FDP4EP \o_label2_data7_REG[24] ( .CK(clk), .CE(n146), .R(n261), .D(n30), .Q(o_label2_data7[24]));
Q_FDP4EP \o_label2_data7_REG[25] ( .CK(clk), .CE(n146), .R(n261), .D(n31), .Q(o_label2_data7[25]));
Q_FDP4EP \o_label2_data7_REG[26] ( .CK(clk), .CE(n146), .R(n261), .D(n32), .Q(o_label2_data7[26]));
Q_FDP4EP \o_label2_data7_REG[27] ( .CK(clk), .CE(n146), .R(n261), .D(n33), .Q(o_label2_data7[27]));
Q_FDP4EP \o_label2_data7_REG[28] ( .CK(clk), .CE(n146), .R(n261), .D(n34), .Q(o_label2_data7[28]));
Q_FDP4EP \o_label2_data7_REG[29] ( .CK(clk), .CE(n146), .R(n261), .D(n35), .Q(o_label2_data7[29]));
Q_FDP4EP \o_label2_data7_REG[30] ( .CK(clk), .CE(n146), .R(n261), .D(n36), .Q(o_label2_data7[30]));
Q_FDP4EP \o_label2_data7_REG[31] ( .CK(clk), .CE(n146), .R(n261), .D(n37), .Q(o_label2_data7[31]));
Q_FDP4EP \o_label2_config_REG[0] ( .CK(clk), .CE(n145), .R(n261), .D(n6), .Q(o_label2_config[0]));
Q_FDP4EP \o_label2_config_REG[1] ( .CK(clk), .CE(n145), .R(n261), .D(n7), .Q(o_label2_config[1]));
Q_FDP4EP \o_label2_config_REG[2] ( .CK(clk), .CE(n145), .R(n261), .D(n8), .Q(o_label2_config[2]));
Q_FDP4EP \o_label2_config_REG[3] ( .CK(clk), .CE(n145), .R(n261), .D(n9), .Q(o_label2_config[3]));
Q_FDP4EP \o_label2_config_REG[4] ( .CK(clk), .CE(n145), .R(n261), .D(n10), .Q(o_label2_config[4]));
Q_FDP4EP \o_label2_config_REG[5] ( .CK(clk), .CE(n145), .R(n261), .D(n11), .Q(o_label2_config[5]));
Q_FDP4EP \o_label2_config_REG[6] ( .CK(clk), .CE(n145), .R(n261), .D(n12), .Q(o_label2_config[6]));
Q_FDP4EP \o_label2_config_REG[7] ( .CK(clk), .CE(n145), .R(n261), .D(n13), .Q(o_label2_config[7]));
Q_FDP4EP \o_label2_config_REG[9] ( .CK(clk), .CE(n145), .R(n261), .D(n31), .Q(o_label2_config[9]));
Q_FDP4EP \o_label2_config_REG[10] ( .CK(clk), .CE(n145), .R(n261), .D(n32), .Q(o_label2_config[10]));
Q_FDP4EP \o_label2_config_REG[11] ( .CK(clk), .CE(n145), .R(n261), .D(n33), .Q(o_label2_config[11]));
Q_FDP4EP \o_label2_config_REG[12] ( .CK(clk), .CE(n145), .R(n261), .D(n34), .Q(o_label2_config[12]));
Q_FDP4EP \o_label2_config_REG[13] ( .CK(clk), .CE(n145), .R(n261), .D(n35), .Q(o_label2_config[13]));
Q_FDP4EP \o_label2_config_REG[14] ( .CK(clk), .CE(n145), .R(n261), .D(n36), .Q(o_label2_config[14]));
Q_FDP4EP \o_label2_config_REG[15] ( .CK(clk), .CE(n145), .R(n261), .D(n37), .Q(o_label2_config[15]));
Q_FDP4EP \o_label1_data0_REG[0] ( .CK(clk), .CE(n144), .R(n261), .D(n6), .Q(o_label1_data0[0]));
Q_FDP4EP \o_label1_data0_REG[1] ( .CK(clk), .CE(n144), .R(n261), .D(n7), .Q(o_label1_data0[1]));
Q_FDP4EP \o_label1_data0_REG[2] ( .CK(clk), .CE(n144), .R(n261), .D(n8), .Q(o_label1_data0[2]));
Q_FDP4EP \o_label1_data0_REG[3] ( .CK(clk), .CE(n144), .R(n261), .D(n9), .Q(o_label1_data0[3]));
Q_FDP4EP \o_label1_data0_REG[4] ( .CK(clk), .CE(n144), .R(n261), .D(n10), .Q(o_label1_data0[4]));
Q_FDP4EP \o_label1_data0_REG[5] ( .CK(clk), .CE(n144), .R(n261), .D(n11), .Q(o_label1_data0[5]));
Q_FDP4EP \o_label1_data0_REG[6] ( .CK(clk), .CE(n144), .R(n261), .D(n12), .Q(o_label1_data0[6]));
Q_FDP4EP \o_label1_data0_REG[7] ( .CK(clk), .CE(n144), .R(n261), .D(n13), .Q(o_label1_data0[7]));
Q_FDP4EP \o_label1_data0_REG[8] ( .CK(clk), .CE(n144), .R(n261), .D(n14), .Q(o_label1_data0[8]));
Q_FDP4EP \o_label1_data0_REG[9] ( .CK(clk), .CE(n144), .R(n261), .D(n15), .Q(o_label1_data0[9]));
Q_FDP4EP \o_label1_data0_REG[10] ( .CK(clk), .CE(n144), .R(n261), .D(n16), .Q(o_label1_data0[10]));
Q_FDP4EP \o_label1_data0_REG[11] ( .CK(clk), .CE(n144), .R(n261), .D(n17), .Q(o_label1_data0[11]));
Q_FDP4EP \o_label1_data0_REG[12] ( .CK(clk), .CE(n144), .R(n261), .D(n18), .Q(o_label1_data0[12]));
Q_FDP4EP \o_label1_data0_REG[13] ( .CK(clk), .CE(n144), .R(n261), .D(n19), .Q(o_label1_data0[13]));
Q_FDP4EP \o_label1_data0_REG[14] ( .CK(clk), .CE(n144), .R(n261), .D(n20), .Q(o_label1_data0[14]));
Q_FDP4EP \o_label1_data0_REG[15] ( .CK(clk), .CE(n144), .R(n261), .D(n21), .Q(o_label1_data0[15]));
Q_FDP4EP \o_label1_data0_REG[16] ( .CK(clk), .CE(n144), .R(n261), .D(n22), .Q(o_label1_data0[16]));
Q_FDP4EP \o_label1_data0_REG[17] ( .CK(clk), .CE(n144), .R(n261), .D(n23), .Q(o_label1_data0[17]));
Q_FDP4EP \o_label1_data0_REG[18] ( .CK(clk), .CE(n144), .R(n261), .D(n24), .Q(o_label1_data0[18]));
Q_FDP4EP \o_label1_data0_REG[19] ( .CK(clk), .CE(n144), .R(n261), .D(n25), .Q(o_label1_data0[19]));
Q_FDP4EP \o_label1_data0_REG[20] ( .CK(clk), .CE(n144), .R(n261), .D(n26), .Q(o_label1_data0[20]));
Q_FDP4EP \o_label1_data0_REG[21] ( .CK(clk), .CE(n144), .R(n261), .D(n27), .Q(o_label1_data0[21]));
Q_FDP4EP \o_label1_data0_REG[22] ( .CK(clk), .CE(n144), .R(n261), .D(n28), .Q(o_label1_data0[22]));
Q_FDP4EP \o_label1_data0_REG[23] ( .CK(clk), .CE(n144), .R(n261), .D(n29), .Q(o_label1_data0[23]));
Q_FDP4EP \o_label1_data0_REG[24] ( .CK(clk), .CE(n144), .R(n261), .D(n30), .Q(o_label1_data0[24]));
Q_FDP4EP \o_label1_data0_REG[25] ( .CK(clk), .CE(n144), .R(n261), .D(n31), .Q(o_label1_data0[25]));
Q_FDP4EP \o_label1_data0_REG[26] ( .CK(clk), .CE(n144), .R(n261), .D(n32), .Q(o_label1_data0[26]));
Q_FDP4EP \o_label1_data0_REG[27] ( .CK(clk), .CE(n144), .R(n261), .D(n33), .Q(o_label1_data0[27]));
Q_FDP4EP \o_label1_data0_REG[28] ( .CK(clk), .CE(n144), .R(n261), .D(n34), .Q(o_label1_data0[28]));
Q_FDP4EP \o_label1_data0_REG[29] ( .CK(clk), .CE(n144), .R(n261), .D(n35), .Q(o_label1_data0[29]));
Q_FDP4EP \o_label1_data0_REG[30] ( .CK(clk), .CE(n144), .R(n261), .D(n36), .Q(o_label1_data0[30]));
Q_FDP4EP \o_label1_data0_REG[31] ( .CK(clk), .CE(n144), .R(n261), .D(n37), .Q(o_label1_data0[31]));
Q_FDP4EP \o_label1_data1_REG[0] ( .CK(clk), .CE(n143), .R(n261), .D(n6), .Q(o_label1_data1[0]));
Q_FDP4EP \o_label1_data1_REG[1] ( .CK(clk), .CE(n143), .R(n261), .D(n7), .Q(o_label1_data1[1]));
Q_FDP4EP \o_label1_data1_REG[2] ( .CK(clk), .CE(n143), .R(n261), .D(n8), .Q(o_label1_data1[2]));
Q_FDP4EP \o_label1_data1_REG[3] ( .CK(clk), .CE(n143), .R(n261), .D(n9), .Q(o_label1_data1[3]));
Q_FDP4EP \o_label1_data1_REG[4] ( .CK(clk), .CE(n143), .R(n261), .D(n10), .Q(o_label1_data1[4]));
Q_FDP4EP \o_label1_data1_REG[5] ( .CK(clk), .CE(n143), .R(n261), .D(n11), .Q(o_label1_data1[5]));
Q_FDP4EP \o_label1_data1_REG[6] ( .CK(clk), .CE(n143), .R(n261), .D(n12), .Q(o_label1_data1[6]));
Q_FDP4EP \o_label1_data1_REG[7] ( .CK(clk), .CE(n143), .R(n261), .D(n13), .Q(o_label1_data1[7]));
Q_FDP4EP \o_label1_data1_REG[8] ( .CK(clk), .CE(n143), .R(n261), .D(n14), .Q(o_label1_data1[8]));
Q_FDP4EP \o_label1_data1_REG[9] ( .CK(clk), .CE(n143), .R(n261), .D(n15), .Q(o_label1_data1[9]));
Q_FDP4EP \o_label1_data1_REG[10] ( .CK(clk), .CE(n143), .R(n261), .D(n16), .Q(o_label1_data1[10]));
Q_FDP4EP \o_label1_data1_REG[11] ( .CK(clk), .CE(n143), .R(n261), .D(n17), .Q(o_label1_data1[11]));
Q_FDP4EP \o_label1_data1_REG[12] ( .CK(clk), .CE(n143), .R(n261), .D(n18), .Q(o_label1_data1[12]));
Q_FDP4EP \o_label1_data1_REG[13] ( .CK(clk), .CE(n143), .R(n261), .D(n19), .Q(o_label1_data1[13]));
Q_FDP4EP \o_label1_data1_REG[14] ( .CK(clk), .CE(n143), .R(n261), .D(n20), .Q(o_label1_data1[14]));
Q_FDP4EP \o_label1_data1_REG[15] ( .CK(clk), .CE(n143), .R(n261), .D(n21), .Q(o_label1_data1[15]));
Q_FDP4EP \o_label1_data1_REG[16] ( .CK(clk), .CE(n143), .R(n261), .D(n22), .Q(o_label1_data1[16]));
Q_FDP4EP \o_label1_data1_REG[17] ( .CK(clk), .CE(n143), .R(n261), .D(n23), .Q(o_label1_data1[17]));
Q_FDP4EP \o_label1_data1_REG[18] ( .CK(clk), .CE(n143), .R(n261), .D(n24), .Q(o_label1_data1[18]));
Q_FDP4EP \o_label1_data1_REG[19] ( .CK(clk), .CE(n143), .R(n261), .D(n25), .Q(o_label1_data1[19]));
Q_FDP4EP \o_label1_data1_REG[20] ( .CK(clk), .CE(n143), .R(n261), .D(n26), .Q(o_label1_data1[20]));
Q_FDP4EP \o_label1_data1_REG[21] ( .CK(clk), .CE(n143), .R(n261), .D(n27), .Q(o_label1_data1[21]));
Q_FDP4EP \o_label1_data1_REG[22] ( .CK(clk), .CE(n143), .R(n261), .D(n28), .Q(o_label1_data1[22]));
Q_FDP4EP \o_label1_data1_REG[23] ( .CK(clk), .CE(n143), .R(n261), .D(n29), .Q(o_label1_data1[23]));
Q_FDP4EP \o_label1_data1_REG[24] ( .CK(clk), .CE(n143), .R(n261), .D(n30), .Q(o_label1_data1[24]));
Q_FDP4EP \o_label1_data1_REG[25] ( .CK(clk), .CE(n143), .R(n261), .D(n31), .Q(o_label1_data1[25]));
Q_FDP4EP \o_label1_data1_REG[26] ( .CK(clk), .CE(n143), .R(n261), .D(n32), .Q(o_label1_data1[26]));
Q_FDP4EP \o_label1_data1_REG[27] ( .CK(clk), .CE(n143), .R(n261), .D(n33), .Q(o_label1_data1[27]));
Q_FDP4EP \o_label1_data1_REG[28] ( .CK(clk), .CE(n143), .R(n261), .D(n34), .Q(o_label1_data1[28]));
Q_FDP4EP \o_label1_data1_REG[29] ( .CK(clk), .CE(n143), .R(n261), .D(n35), .Q(o_label1_data1[29]));
Q_FDP4EP \o_label1_data1_REG[30] ( .CK(clk), .CE(n143), .R(n261), .D(n36), .Q(o_label1_data1[30]));
Q_FDP4EP \o_label1_data1_REG[31] ( .CK(clk), .CE(n143), .R(n261), .D(n37), .Q(o_label1_data1[31]));
Q_FDP4EP \o_label1_data2_REG[0] ( .CK(clk), .CE(n142), .R(n261), .D(n6), .Q(o_label1_data2[0]));
Q_FDP4EP \o_label1_data2_REG[1] ( .CK(clk), .CE(n142), .R(n261), .D(n7), .Q(o_label1_data2[1]));
Q_FDP4EP \o_label1_data2_REG[2] ( .CK(clk), .CE(n142), .R(n261), .D(n8), .Q(o_label1_data2[2]));
Q_FDP4EP \o_label1_data2_REG[3] ( .CK(clk), .CE(n142), .R(n261), .D(n9), .Q(o_label1_data2[3]));
Q_FDP4EP \o_label1_data2_REG[4] ( .CK(clk), .CE(n142), .R(n261), .D(n10), .Q(o_label1_data2[4]));
Q_FDP4EP \o_label1_data2_REG[5] ( .CK(clk), .CE(n142), .R(n261), .D(n11), .Q(o_label1_data2[5]));
Q_FDP4EP \o_label1_data2_REG[6] ( .CK(clk), .CE(n142), .R(n261), .D(n12), .Q(o_label1_data2[6]));
Q_FDP4EP \o_label1_data2_REG[7] ( .CK(clk), .CE(n142), .R(n261), .D(n13), .Q(o_label1_data2[7]));
Q_FDP4EP \o_label1_data2_REG[8] ( .CK(clk), .CE(n142), .R(n261), .D(n14), .Q(o_label1_data2[8]));
Q_FDP4EP \o_label1_data2_REG[9] ( .CK(clk), .CE(n142), .R(n261), .D(n15), .Q(o_label1_data2[9]));
Q_FDP4EP \o_label1_data2_REG[10] ( .CK(clk), .CE(n142), .R(n261), .D(n16), .Q(o_label1_data2[10]));
Q_FDP4EP \o_label1_data2_REG[11] ( .CK(clk), .CE(n142), .R(n261), .D(n17), .Q(o_label1_data2[11]));
Q_FDP4EP \o_label1_data2_REG[12] ( .CK(clk), .CE(n142), .R(n261), .D(n18), .Q(o_label1_data2[12]));
Q_FDP4EP \o_label1_data2_REG[13] ( .CK(clk), .CE(n142), .R(n261), .D(n19), .Q(o_label1_data2[13]));
Q_FDP4EP \o_label1_data2_REG[14] ( .CK(clk), .CE(n142), .R(n261), .D(n20), .Q(o_label1_data2[14]));
Q_FDP4EP \o_label1_data2_REG[15] ( .CK(clk), .CE(n142), .R(n261), .D(n21), .Q(o_label1_data2[15]));
Q_FDP4EP \o_label1_data2_REG[16] ( .CK(clk), .CE(n142), .R(n261), .D(n22), .Q(o_label1_data2[16]));
Q_FDP4EP \o_label1_data2_REG[17] ( .CK(clk), .CE(n142), .R(n261), .D(n23), .Q(o_label1_data2[17]));
Q_FDP4EP \o_label1_data2_REG[18] ( .CK(clk), .CE(n142), .R(n261), .D(n24), .Q(o_label1_data2[18]));
Q_FDP4EP \o_label1_data2_REG[19] ( .CK(clk), .CE(n142), .R(n261), .D(n25), .Q(o_label1_data2[19]));
Q_FDP4EP \o_label1_data2_REG[20] ( .CK(clk), .CE(n142), .R(n261), .D(n26), .Q(o_label1_data2[20]));
Q_FDP4EP \o_label1_data2_REG[21] ( .CK(clk), .CE(n142), .R(n261), .D(n27), .Q(o_label1_data2[21]));
Q_FDP4EP \o_label1_data2_REG[22] ( .CK(clk), .CE(n142), .R(n261), .D(n28), .Q(o_label1_data2[22]));
Q_FDP4EP \o_label1_data2_REG[23] ( .CK(clk), .CE(n142), .R(n261), .D(n29), .Q(o_label1_data2[23]));
Q_FDP4EP \o_label1_data2_REG[24] ( .CK(clk), .CE(n142), .R(n261), .D(n30), .Q(o_label1_data2[24]));
Q_FDP4EP \o_label1_data2_REG[25] ( .CK(clk), .CE(n142), .R(n261), .D(n31), .Q(o_label1_data2[25]));
Q_FDP4EP \o_label1_data2_REG[26] ( .CK(clk), .CE(n142), .R(n261), .D(n32), .Q(o_label1_data2[26]));
Q_FDP4EP \o_label1_data2_REG[27] ( .CK(clk), .CE(n142), .R(n261), .D(n33), .Q(o_label1_data2[27]));
Q_FDP4EP \o_label1_data2_REG[28] ( .CK(clk), .CE(n142), .R(n261), .D(n34), .Q(o_label1_data2[28]));
Q_FDP4EP \o_label1_data2_REG[29] ( .CK(clk), .CE(n142), .R(n261), .D(n35), .Q(o_label1_data2[29]));
Q_FDP4EP \o_label1_data2_REG[30] ( .CK(clk), .CE(n142), .R(n261), .D(n36), .Q(o_label1_data2[30]));
Q_FDP4EP \o_label1_data2_REG[31] ( .CK(clk), .CE(n142), .R(n261), .D(n37), .Q(o_label1_data2[31]));
Q_FDP4EP \o_label1_data3_REG[0] ( .CK(clk), .CE(n141), .R(n261), .D(n6), .Q(o_label1_data3[0]));
Q_FDP4EP \o_label1_data3_REG[1] ( .CK(clk), .CE(n141), .R(n261), .D(n7), .Q(o_label1_data3[1]));
Q_FDP4EP \o_label1_data3_REG[2] ( .CK(clk), .CE(n141), .R(n261), .D(n8), .Q(o_label1_data3[2]));
Q_FDP4EP \o_label1_data3_REG[3] ( .CK(clk), .CE(n141), .R(n261), .D(n9), .Q(o_label1_data3[3]));
Q_FDP4EP \o_label1_data3_REG[4] ( .CK(clk), .CE(n141), .R(n261), .D(n10), .Q(o_label1_data3[4]));
Q_FDP4EP \o_label1_data3_REG[5] ( .CK(clk), .CE(n141), .R(n261), .D(n11), .Q(o_label1_data3[5]));
Q_FDP4EP \o_label1_data3_REG[6] ( .CK(clk), .CE(n141), .R(n261), .D(n12), .Q(o_label1_data3[6]));
Q_FDP4EP \o_label1_data3_REG[7] ( .CK(clk), .CE(n141), .R(n261), .D(n13), .Q(o_label1_data3[7]));
Q_FDP4EP \o_label1_data3_REG[8] ( .CK(clk), .CE(n141), .R(n261), .D(n14), .Q(o_label1_data3[8]));
Q_FDP4EP \o_label1_data3_REG[9] ( .CK(clk), .CE(n141), .R(n261), .D(n15), .Q(o_label1_data3[9]));
Q_FDP4EP \o_label1_data3_REG[10] ( .CK(clk), .CE(n141), .R(n261), .D(n16), .Q(o_label1_data3[10]));
Q_FDP4EP \o_label1_data3_REG[11] ( .CK(clk), .CE(n141), .R(n261), .D(n17), .Q(o_label1_data3[11]));
Q_FDP4EP \o_label1_data3_REG[12] ( .CK(clk), .CE(n141), .R(n261), .D(n18), .Q(o_label1_data3[12]));
Q_FDP4EP \o_label1_data3_REG[13] ( .CK(clk), .CE(n141), .R(n261), .D(n19), .Q(o_label1_data3[13]));
Q_FDP4EP \o_label1_data3_REG[14] ( .CK(clk), .CE(n141), .R(n261), .D(n20), .Q(o_label1_data3[14]));
Q_FDP4EP \o_label1_data3_REG[15] ( .CK(clk), .CE(n141), .R(n261), .D(n21), .Q(o_label1_data3[15]));
Q_FDP4EP \o_label1_data3_REG[16] ( .CK(clk), .CE(n141), .R(n261), .D(n22), .Q(o_label1_data3[16]));
Q_FDP4EP \o_label1_data3_REG[17] ( .CK(clk), .CE(n141), .R(n261), .D(n23), .Q(o_label1_data3[17]));
Q_FDP4EP \o_label1_data3_REG[18] ( .CK(clk), .CE(n141), .R(n261), .D(n24), .Q(o_label1_data3[18]));
Q_FDP4EP \o_label1_data3_REG[19] ( .CK(clk), .CE(n141), .R(n261), .D(n25), .Q(o_label1_data3[19]));
Q_FDP4EP \o_label1_data3_REG[20] ( .CK(clk), .CE(n141), .R(n261), .D(n26), .Q(o_label1_data3[20]));
Q_FDP4EP \o_label1_data3_REG[21] ( .CK(clk), .CE(n141), .R(n261), .D(n27), .Q(o_label1_data3[21]));
Q_FDP4EP \o_label1_data3_REG[22] ( .CK(clk), .CE(n141), .R(n261), .D(n28), .Q(o_label1_data3[22]));
Q_FDP4EP \o_label1_data3_REG[23] ( .CK(clk), .CE(n141), .R(n261), .D(n29), .Q(o_label1_data3[23]));
Q_FDP4EP \o_label1_data3_REG[24] ( .CK(clk), .CE(n141), .R(n261), .D(n30), .Q(o_label1_data3[24]));
Q_FDP4EP \o_label1_data3_REG[25] ( .CK(clk), .CE(n141), .R(n261), .D(n31), .Q(o_label1_data3[25]));
Q_FDP4EP \o_label1_data3_REG[26] ( .CK(clk), .CE(n141), .R(n261), .D(n32), .Q(o_label1_data3[26]));
Q_FDP4EP \o_label1_data3_REG[27] ( .CK(clk), .CE(n141), .R(n261), .D(n33), .Q(o_label1_data3[27]));
Q_FDP4EP \o_label1_data3_REG[28] ( .CK(clk), .CE(n141), .R(n261), .D(n34), .Q(o_label1_data3[28]));
Q_FDP4EP \o_label1_data3_REG[29] ( .CK(clk), .CE(n141), .R(n261), .D(n35), .Q(o_label1_data3[29]));
Q_FDP4EP \o_label1_data3_REG[30] ( .CK(clk), .CE(n141), .R(n261), .D(n36), .Q(o_label1_data3[30]));
Q_FDP4EP \o_label1_data3_REG[31] ( .CK(clk), .CE(n141), .R(n261), .D(n37), .Q(o_label1_data3[31]));
Q_FDP4EP \o_label1_data4_REG[0] ( .CK(clk), .CE(n140), .R(n261), .D(n6), .Q(o_label1_data4[0]));
Q_FDP4EP \o_label1_data4_REG[1] ( .CK(clk), .CE(n140), .R(n261), .D(n7), .Q(o_label1_data4[1]));
Q_FDP4EP \o_label1_data4_REG[2] ( .CK(clk), .CE(n140), .R(n261), .D(n8), .Q(o_label1_data4[2]));
Q_FDP4EP \o_label1_data4_REG[3] ( .CK(clk), .CE(n140), .R(n261), .D(n9), .Q(o_label1_data4[3]));
Q_FDP4EP \o_label1_data4_REG[4] ( .CK(clk), .CE(n140), .R(n261), .D(n10), .Q(o_label1_data4[4]));
Q_FDP4EP \o_label1_data4_REG[5] ( .CK(clk), .CE(n140), .R(n261), .D(n11), .Q(o_label1_data4[5]));
Q_FDP4EP \o_label1_data4_REG[6] ( .CK(clk), .CE(n140), .R(n261), .D(n12), .Q(o_label1_data4[6]));
Q_FDP4EP \o_label1_data4_REG[7] ( .CK(clk), .CE(n140), .R(n261), .D(n13), .Q(o_label1_data4[7]));
Q_FDP4EP \o_label1_data4_REG[8] ( .CK(clk), .CE(n140), .R(n261), .D(n14), .Q(o_label1_data4[8]));
Q_FDP4EP \o_label1_data4_REG[9] ( .CK(clk), .CE(n140), .R(n261), .D(n15), .Q(o_label1_data4[9]));
Q_FDP4EP \o_label1_data4_REG[10] ( .CK(clk), .CE(n140), .R(n261), .D(n16), .Q(o_label1_data4[10]));
Q_FDP4EP \o_label1_data4_REG[11] ( .CK(clk), .CE(n140), .R(n261), .D(n17), .Q(o_label1_data4[11]));
Q_FDP4EP \o_label1_data4_REG[12] ( .CK(clk), .CE(n140), .R(n261), .D(n18), .Q(o_label1_data4[12]));
Q_FDP4EP \o_label1_data4_REG[13] ( .CK(clk), .CE(n140), .R(n261), .D(n19), .Q(o_label1_data4[13]));
Q_FDP4EP \o_label1_data4_REG[14] ( .CK(clk), .CE(n140), .R(n261), .D(n20), .Q(o_label1_data4[14]));
Q_FDP4EP \o_label1_data4_REG[15] ( .CK(clk), .CE(n140), .R(n261), .D(n21), .Q(o_label1_data4[15]));
Q_FDP4EP \o_label1_data4_REG[16] ( .CK(clk), .CE(n140), .R(n261), .D(n22), .Q(o_label1_data4[16]));
Q_FDP4EP \o_label1_data4_REG[17] ( .CK(clk), .CE(n140), .R(n261), .D(n23), .Q(o_label1_data4[17]));
Q_FDP4EP \o_label1_data4_REG[18] ( .CK(clk), .CE(n140), .R(n261), .D(n24), .Q(o_label1_data4[18]));
Q_FDP4EP \o_label1_data4_REG[19] ( .CK(clk), .CE(n140), .R(n261), .D(n25), .Q(o_label1_data4[19]));
Q_FDP4EP \o_label1_data4_REG[20] ( .CK(clk), .CE(n140), .R(n261), .D(n26), .Q(o_label1_data4[20]));
Q_FDP4EP \o_label1_data4_REG[21] ( .CK(clk), .CE(n140), .R(n261), .D(n27), .Q(o_label1_data4[21]));
Q_FDP4EP \o_label1_data4_REG[22] ( .CK(clk), .CE(n140), .R(n261), .D(n28), .Q(o_label1_data4[22]));
Q_FDP4EP \o_label1_data4_REG[23] ( .CK(clk), .CE(n140), .R(n261), .D(n29), .Q(o_label1_data4[23]));
Q_FDP4EP \o_label1_data4_REG[24] ( .CK(clk), .CE(n140), .R(n261), .D(n30), .Q(o_label1_data4[24]));
Q_FDP4EP \o_label1_data4_REG[25] ( .CK(clk), .CE(n140), .R(n261), .D(n31), .Q(o_label1_data4[25]));
Q_FDP4EP \o_label1_data4_REG[26] ( .CK(clk), .CE(n140), .R(n261), .D(n32), .Q(o_label1_data4[26]));
Q_FDP4EP \o_label1_data4_REG[27] ( .CK(clk), .CE(n140), .R(n261), .D(n33), .Q(o_label1_data4[27]));
Q_FDP4EP \o_label1_data4_REG[28] ( .CK(clk), .CE(n140), .R(n261), .D(n34), .Q(o_label1_data4[28]));
Q_FDP4EP \o_label1_data4_REG[29] ( .CK(clk), .CE(n140), .R(n261), .D(n35), .Q(o_label1_data4[29]));
Q_FDP4EP \o_label1_data4_REG[30] ( .CK(clk), .CE(n140), .R(n261), .D(n36), .Q(o_label1_data4[30]));
Q_FDP4EP \o_label1_data4_REG[31] ( .CK(clk), .CE(n140), .R(n261), .D(n37), .Q(o_label1_data4[31]));
Q_FDP4EP \o_label1_data5_REG[0] ( .CK(clk), .CE(n139), .R(n261), .D(n6), .Q(o_label1_data5[0]));
Q_FDP4EP \o_label1_data5_REG[1] ( .CK(clk), .CE(n139), .R(n261), .D(n7), .Q(o_label1_data5[1]));
Q_FDP4EP \o_label1_data5_REG[2] ( .CK(clk), .CE(n139), .R(n261), .D(n8), .Q(o_label1_data5[2]));
Q_FDP4EP \o_label1_data5_REG[3] ( .CK(clk), .CE(n139), .R(n261), .D(n9), .Q(o_label1_data5[3]));
Q_FDP4EP \o_label1_data5_REG[4] ( .CK(clk), .CE(n139), .R(n261), .D(n10), .Q(o_label1_data5[4]));
Q_FDP4EP \o_label1_data5_REG[5] ( .CK(clk), .CE(n139), .R(n261), .D(n11), .Q(o_label1_data5[5]));
Q_FDP4EP \o_label1_data5_REG[6] ( .CK(clk), .CE(n139), .R(n261), .D(n12), .Q(o_label1_data5[6]));
Q_FDP4EP \o_label1_data5_REG[7] ( .CK(clk), .CE(n139), .R(n261), .D(n13), .Q(o_label1_data5[7]));
Q_FDP4EP \o_label1_data5_REG[8] ( .CK(clk), .CE(n139), .R(n261), .D(n14), .Q(o_label1_data5[8]));
Q_FDP4EP \o_label1_data5_REG[9] ( .CK(clk), .CE(n139), .R(n261), .D(n15), .Q(o_label1_data5[9]));
Q_FDP4EP \o_label1_data5_REG[10] ( .CK(clk), .CE(n139), .R(n261), .D(n16), .Q(o_label1_data5[10]));
Q_FDP4EP \o_label1_data5_REG[11] ( .CK(clk), .CE(n139), .R(n261), .D(n17), .Q(o_label1_data5[11]));
Q_FDP4EP \o_label1_data5_REG[12] ( .CK(clk), .CE(n139), .R(n261), .D(n18), .Q(o_label1_data5[12]));
Q_FDP4EP \o_label1_data5_REG[13] ( .CK(clk), .CE(n139), .R(n261), .D(n19), .Q(o_label1_data5[13]));
Q_FDP4EP \o_label1_data5_REG[14] ( .CK(clk), .CE(n139), .R(n261), .D(n20), .Q(o_label1_data5[14]));
Q_FDP4EP \o_label1_data5_REG[15] ( .CK(clk), .CE(n139), .R(n261), .D(n21), .Q(o_label1_data5[15]));
Q_FDP4EP \o_label1_data5_REG[16] ( .CK(clk), .CE(n139), .R(n261), .D(n22), .Q(o_label1_data5[16]));
Q_FDP4EP \o_label1_data5_REG[17] ( .CK(clk), .CE(n139), .R(n261), .D(n23), .Q(o_label1_data5[17]));
Q_FDP4EP \o_label1_data5_REG[18] ( .CK(clk), .CE(n139), .R(n261), .D(n24), .Q(o_label1_data5[18]));
Q_FDP4EP \o_label1_data5_REG[19] ( .CK(clk), .CE(n139), .R(n261), .D(n25), .Q(o_label1_data5[19]));
Q_FDP4EP \o_label1_data5_REG[20] ( .CK(clk), .CE(n139), .R(n261), .D(n26), .Q(o_label1_data5[20]));
Q_FDP4EP \o_label1_data5_REG[21] ( .CK(clk), .CE(n139), .R(n261), .D(n27), .Q(o_label1_data5[21]));
Q_FDP4EP \o_label1_data5_REG[22] ( .CK(clk), .CE(n139), .R(n261), .D(n28), .Q(o_label1_data5[22]));
Q_FDP4EP \o_label1_data5_REG[23] ( .CK(clk), .CE(n139), .R(n261), .D(n29), .Q(o_label1_data5[23]));
Q_FDP4EP \o_label1_data5_REG[24] ( .CK(clk), .CE(n139), .R(n261), .D(n30), .Q(o_label1_data5[24]));
Q_FDP4EP \o_label1_data5_REG[25] ( .CK(clk), .CE(n139), .R(n261), .D(n31), .Q(o_label1_data5[25]));
Q_FDP4EP \o_label1_data5_REG[26] ( .CK(clk), .CE(n139), .R(n261), .D(n32), .Q(o_label1_data5[26]));
Q_FDP4EP \o_label1_data5_REG[27] ( .CK(clk), .CE(n139), .R(n261), .D(n33), .Q(o_label1_data5[27]));
Q_FDP4EP \o_label1_data5_REG[28] ( .CK(clk), .CE(n139), .R(n261), .D(n34), .Q(o_label1_data5[28]));
Q_FDP4EP \o_label1_data5_REG[29] ( .CK(clk), .CE(n139), .R(n261), .D(n35), .Q(o_label1_data5[29]));
Q_FDP4EP \o_label1_data5_REG[30] ( .CK(clk), .CE(n139), .R(n261), .D(n36), .Q(o_label1_data5[30]));
Q_FDP4EP \o_label1_data5_REG[31] ( .CK(clk), .CE(n139), .R(n261), .D(n37), .Q(o_label1_data5[31]));
Q_FDP4EP \o_label1_data6_REG[0] ( .CK(clk), .CE(n138), .R(n261), .D(n6), .Q(o_label1_data6[0]));
Q_FDP4EP \o_label1_data6_REG[1] ( .CK(clk), .CE(n138), .R(n261), .D(n7), .Q(o_label1_data6[1]));
Q_FDP4EP \o_label1_data6_REG[2] ( .CK(clk), .CE(n138), .R(n261), .D(n8), .Q(o_label1_data6[2]));
Q_FDP4EP \o_label1_data6_REG[3] ( .CK(clk), .CE(n138), .R(n261), .D(n9), .Q(o_label1_data6[3]));
Q_FDP4EP \o_label1_data6_REG[4] ( .CK(clk), .CE(n138), .R(n261), .D(n10), .Q(o_label1_data6[4]));
Q_FDP4EP \o_label1_data6_REG[5] ( .CK(clk), .CE(n138), .R(n261), .D(n11), .Q(o_label1_data6[5]));
Q_FDP4EP \o_label1_data6_REG[6] ( .CK(clk), .CE(n138), .R(n261), .D(n12), .Q(o_label1_data6[6]));
Q_FDP4EP \o_label1_data6_REG[7] ( .CK(clk), .CE(n138), .R(n261), .D(n13), .Q(o_label1_data6[7]));
Q_FDP4EP \o_label1_data6_REG[8] ( .CK(clk), .CE(n138), .R(n261), .D(n14), .Q(o_label1_data6[8]));
Q_FDP4EP \o_label1_data6_REG[9] ( .CK(clk), .CE(n138), .R(n261), .D(n15), .Q(o_label1_data6[9]));
Q_FDP4EP \o_label1_data6_REG[10] ( .CK(clk), .CE(n138), .R(n261), .D(n16), .Q(o_label1_data6[10]));
Q_FDP4EP \o_label1_data6_REG[11] ( .CK(clk), .CE(n138), .R(n261), .D(n17), .Q(o_label1_data6[11]));
Q_FDP4EP \o_label1_data6_REG[12] ( .CK(clk), .CE(n138), .R(n261), .D(n18), .Q(o_label1_data6[12]));
Q_FDP4EP \o_label1_data6_REG[13] ( .CK(clk), .CE(n138), .R(n261), .D(n19), .Q(o_label1_data6[13]));
Q_FDP4EP \o_label1_data6_REG[14] ( .CK(clk), .CE(n138), .R(n261), .D(n20), .Q(o_label1_data6[14]));
Q_FDP4EP \o_label1_data6_REG[15] ( .CK(clk), .CE(n138), .R(n261), .D(n21), .Q(o_label1_data6[15]));
Q_FDP4EP \o_label1_data6_REG[16] ( .CK(clk), .CE(n138), .R(n261), .D(n22), .Q(o_label1_data6[16]));
Q_FDP4EP \o_label1_data6_REG[17] ( .CK(clk), .CE(n138), .R(n261), .D(n23), .Q(o_label1_data6[17]));
Q_FDP4EP \o_label1_data6_REG[18] ( .CK(clk), .CE(n138), .R(n261), .D(n24), .Q(o_label1_data6[18]));
Q_FDP4EP \o_label1_data6_REG[19] ( .CK(clk), .CE(n138), .R(n261), .D(n25), .Q(o_label1_data6[19]));
Q_FDP4EP \o_label1_data6_REG[20] ( .CK(clk), .CE(n138), .R(n261), .D(n26), .Q(o_label1_data6[20]));
Q_FDP4EP \o_label1_data6_REG[21] ( .CK(clk), .CE(n138), .R(n261), .D(n27), .Q(o_label1_data6[21]));
Q_FDP4EP \o_label1_data6_REG[22] ( .CK(clk), .CE(n138), .R(n261), .D(n28), .Q(o_label1_data6[22]));
Q_FDP4EP \o_label1_data6_REG[23] ( .CK(clk), .CE(n138), .R(n261), .D(n29), .Q(o_label1_data6[23]));
Q_FDP4EP \o_label1_data6_REG[24] ( .CK(clk), .CE(n138), .R(n261), .D(n30), .Q(o_label1_data6[24]));
Q_FDP4EP \o_label1_data6_REG[25] ( .CK(clk), .CE(n138), .R(n261), .D(n31), .Q(o_label1_data6[25]));
Q_FDP4EP \o_label1_data6_REG[26] ( .CK(clk), .CE(n138), .R(n261), .D(n32), .Q(o_label1_data6[26]));
Q_FDP4EP \o_label1_data6_REG[27] ( .CK(clk), .CE(n138), .R(n261), .D(n33), .Q(o_label1_data6[27]));
Q_FDP4EP \o_label1_data6_REG[28] ( .CK(clk), .CE(n138), .R(n261), .D(n34), .Q(o_label1_data6[28]));
Q_FDP4EP \o_label1_data6_REG[29] ( .CK(clk), .CE(n138), .R(n261), .D(n35), .Q(o_label1_data6[29]));
Q_FDP4EP \o_label1_data6_REG[30] ( .CK(clk), .CE(n138), .R(n261), .D(n36), .Q(o_label1_data6[30]));
Q_FDP4EP \o_label1_data6_REG[31] ( .CK(clk), .CE(n138), .R(n261), .D(n37), .Q(o_label1_data6[31]));
Q_FDP4EP \o_label1_data7_REG[0] ( .CK(clk), .CE(n137), .R(n261), .D(n6), .Q(o_label1_data7[0]));
Q_FDP4EP \o_label1_data7_REG[1] ( .CK(clk), .CE(n137), .R(n261), .D(n7), .Q(o_label1_data7[1]));
Q_FDP4EP \o_label1_data7_REG[2] ( .CK(clk), .CE(n137), .R(n261), .D(n8), .Q(o_label1_data7[2]));
Q_FDP4EP \o_label1_data7_REG[3] ( .CK(clk), .CE(n137), .R(n261), .D(n9), .Q(o_label1_data7[3]));
Q_FDP4EP \o_label1_data7_REG[4] ( .CK(clk), .CE(n137), .R(n261), .D(n10), .Q(o_label1_data7[4]));
Q_FDP4EP \o_label1_data7_REG[5] ( .CK(clk), .CE(n137), .R(n261), .D(n11), .Q(o_label1_data7[5]));
Q_FDP4EP \o_label1_data7_REG[6] ( .CK(clk), .CE(n137), .R(n261), .D(n12), .Q(o_label1_data7[6]));
Q_FDP4EP \o_label1_data7_REG[7] ( .CK(clk), .CE(n137), .R(n261), .D(n13), .Q(o_label1_data7[7]));
Q_FDP4EP \o_label1_data7_REG[8] ( .CK(clk), .CE(n137), .R(n261), .D(n14), .Q(o_label1_data7[8]));
Q_FDP4EP \o_label1_data7_REG[9] ( .CK(clk), .CE(n137), .R(n261), .D(n15), .Q(o_label1_data7[9]));
Q_FDP4EP \o_label1_data7_REG[10] ( .CK(clk), .CE(n137), .R(n261), .D(n16), .Q(o_label1_data7[10]));
Q_FDP4EP \o_label1_data7_REG[11] ( .CK(clk), .CE(n137), .R(n261), .D(n17), .Q(o_label1_data7[11]));
Q_FDP4EP \o_label1_data7_REG[12] ( .CK(clk), .CE(n137), .R(n261), .D(n18), .Q(o_label1_data7[12]));
Q_FDP4EP \o_label1_data7_REG[13] ( .CK(clk), .CE(n137), .R(n261), .D(n19), .Q(o_label1_data7[13]));
Q_FDP4EP \o_label1_data7_REG[14] ( .CK(clk), .CE(n137), .R(n261), .D(n20), .Q(o_label1_data7[14]));
Q_FDP4EP \o_label1_data7_REG[15] ( .CK(clk), .CE(n137), .R(n261), .D(n21), .Q(o_label1_data7[15]));
Q_FDP4EP \o_label1_data7_REG[16] ( .CK(clk), .CE(n137), .R(n261), .D(n22), .Q(o_label1_data7[16]));
Q_FDP4EP \o_label1_data7_REG[17] ( .CK(clk), .CE(n137), .R(n261), .D(n23), .Q(o_label1_data7[17]));
Q_FDP4EP \o_label1_data7_REG[18] ( .CK(clk), .CE(n137), .R(n261), .D(n24), .Q(o_label1_data7[18]));
Q_FDP4EP \o_label1_data7_REG[19] ( .CK(clk), .CE(n137), .R(n261), .D(n25), .Q(o_label1_data7[19]));
Q_FDP4EP \o_label1_data7_REG[20] ( .CK(clk), .CE(n137), .R(n261), .D(n26), .Q(o_label1_data7[20]));
Q_FDP4EP \o_label1_data7_REG[21] ( .CK(clk), .CE(n137), .R(n261), .D(n27), .Q(o_label1_data7[21]));
Q_FDP4EP \o_label1_data7_REG[22] ( .CK(clk), .CE(n137), .R(n261), .D(n28), .Q(o_label1_data7[22]));
Q_FDP4EP \o_label1_data7_REG[23] ( .CK(clk), .CE(n137), .R(n261), .D(n29), .Q(o_label1_data7[23]));
Q_FDP4EP \o_label1_data7_REG[24] ( .CK(clk), .CE(n137), .R(n261), .D(n30), .Q(o_label1_data7[24]));
Q_FDP4EP \o_label1_data7_REG[25] ( .CK(clk), .CE(n137), .R(n261), .D(n31), .Q(o_label1_data7[25]));
Q_FDP4EP \o_label1_data7_REG[26] ( .CK(clk), .CE(n137), .R(n261), .D(n32), .Q(o_label1_data7[26]));
Q_FDP4EP \o_label1_data7_REG[27] ( .CK(clk), .CE(n137), .R(n261), .D(n33), .Q(o_label1_data7[27]));
Q_FDP4EP \o_label1_data7_REG[28] ( .CK(clk), .CE(n137), .R(n261), .D(n34), .Q(o_label1_data7[28]));
Q_FDP4EP \o_label1_data7_REG[29] ( .CK(clk), .CE(n137), .R(n261), .D(n35), .Q(o_label1_data7[29]));
Q_FDP4EP \o_label1_data7_REG[30] ( .CK(clk), .CE(n137), .R(n261), .D(n36), .Q(o_label1_data7[30]));
Q_FDP4EP \o_label1_data7_REG[31] ( .CK(clk), .CE(n137), .R(n261), .D(n37), .Q(o_label1_data7[31]));
Q_FDP4EP \o_label1_config_REG[0] ( .CK(clk), .CE(n136), .R(n261), .D(n6), .Q(o_label1_config[0]));
Q_FDP4EP \o_label1_config_REG[1] ( .CK(clk), .CE(n136), .R(n261), .D(n7), .Q(o_label1_config[1]));
Q_FDP4EP \o_label1_config_REG[2] ( .CK(clk), .CE(n136), .R(n261), .D(n8), .Q(o_label1_config[2]));
Q_FDP4EP \o_label1_config_REG[3] ( .CK(clk), .CE(n136), .R(n261), .D(n9), .Q(o_label1_config[3]));
Q_FDP4EP \o_label1_config_REG[4] ( .CK(clk), .CE(n136), .R(n261), .D(n10), .Q(o_label1_config[4]));
Q_FDP4EP \o_label1_config_REG[5] ( .CK(clk), .CE(n136), .R(n261), .D(n11), .Q(o_label1_config[5]));
Q_FDP4EP \o_label1_config_REG[6] ( .CK(clk), .CE(n136), .R(n261), .D(n12), .Q(o_label1_config[6]));
Q_FDP4EP \o_label1_config_REG[7] ( .CK(clk), .CE(n136), .R(n261), .D(n13), .Q(o_label1_config[7]));
Q_FDP4EP \o_label1_config_REG[9] ( .CK(clk), .CE(n136), .R(n261), .D(n31), .Q(o_label1_config[9]));
Q_FDP4EP \o_label1_config_REG[10] ( .CK(clk), .CE(n136), .R(n261), .D(n32), .Q(o_label1_config[10]));
Q_FDP4EP \o_label1_config_REG[11] ( .CK(clk), .CE(n136), .R(n261), .D(n33), .Q(o_label1_config[11]));
Q_FDP4EP \o_label1_config_REG[12] ( .CK(clk), .CE(n136), .R(n261), .D(n34), .Q(o_label1_config[12]));
Q_FDP4EP \o_label1_config_REG[13] ( .CK(clk), .CE(n136), .R(n261), .D(n35), .Q(o_label1_config[13]));
Q_FDP4EP \o_label1_config_REG[14] ( .CK(clk), .CE(n136), .R(n261), .D(n36), .Q(o_label1_config[14]));
Q_FDP4EP \o_label1_config_REG[15] ( .CK(clk), .CE(n136), .R(n261), .D(n37), .Q(o_label1_config[15]));
Q_FDP4EP \o_label0_data0_REG[0] ( .CK(clk), .CE(n135), .R(n261), .D(n6), .Q(o_label0_data0[0]));
Q_FDP4EP \o_label0_data0_REG[1] ( .CK(clk), .CE(n135), .R(n261), .D(n7), .Q(o_label0_data0[1]));
Q_FDP4EP \o_label0_data0_REG[2] ( .CK(clk), .CE(n135), .R(n261), .D(n8), .Q(o_label0_data0[2]));
Q_FDP4EP \o_label0_data0_REG[3] ( .CK(clk), .CE(n135), .R(n261), .D(n9), .Q(o_label0_data0[3]));
Q_FDP4EP \o_label0_data0_REG[4] ( .CK(clk), .CE(n135), .R(n261), .D(n10), .Q(o_label0_data0[4]));
Q_FDP4EP \o_label0_data0_REG[5] ( .CK(clk), .CE(n135), .R(n261), .D(n11), .Q(o_label0_data0[5]));
Q_FDP4EP \o_label0_data0_REG[6] ( .CK(clk), .CE(n135), .R(n261), .D(n12), .Q(o_label0_data0[6]));
Q_FDP4EP \o_label0_data0_REG[7] ( .CK(clk), .CE(n135), .R(n261), .D(n13), .Q(o_label0_data0[7]));
Q_FDP4EP \o_label0_data0_REG[8] ( .CK(clk), .CE(n135), .R(n261), .D(n14), .Q(o_label0_data0[8]));
Q_FDP4EP \o_label0_data0_REG[9] ( .CK(clk), .CE(n135), .R(n261), .D(n15), .Q(o_label0_data0[9]));
Q_FDP4EP \o_label0_data0_REG[10] ( .CK(clk), .CE(n135), .R(n261), .D(n16), .Q(o_label0_data0[10]));
Q_FDP4EP \o_label0_data0_REG[11] ( .CK(clk), .CE(n135), .R(n261), .D(n17), .Q(o_label0_data0[11]));
Q_FDP4EP \o_label0_data0_REG[12] ( .CK(clk), .CE(n135), .R(n261), .D(n18), .Q(o_label0_data0[12]));
Q_FDP4EP \o_label0_data0_REG[13] ( .CK(clk), .CE(n135), .R(n261), .D(n19), .Q(o_label0_data0[13]));
Q_FDP4EP \o_label0_data0_REG[14] ( .CK(clk), .CE(n135), .R(n261), .D(n20), .Q(o_label0_data0[14]));
Q_FDP4EP \o_label0_data0_REG[15] ( .CK(clk), .CE(n135), .R(n261), .D(n21), .Q(o_label0_data0[15]));
Q_FDP4EP \o_label0_data0_REG[16] ( .CK(clk), .CE(n135), .R(n261), .D(n22), .Q(o_label0_data0[16]));
Q_FDP4EP \o_label0_data0_REG[17] ( .CK(clk), .CE(n135), .R(n261), .D(n23), .Q(o_label0_data0[17]));
Q_FDP4EP \o_label0_data0_REG[18] ( .CK(clk), .CE(n135), .R(n261), .D(n24), .Q(o_label0_data0[18]));
Q_FDP4EP \o_label0_data0_REG[19] ( .CK(clk), .CE(n135), .R(n261), .D(n25), .Q(o_label0_data0[19]));
Q_FDP4EP \o_label0_data0_REG[20] ( .CK(clk), .CE(n135), .R(n261), .D(n26), .Q(o_label0_data0[20]));
Q_FDP4EP \o_label0_data0_REG[21] ( .CK(clk), .CE(n135), .R(n261), .D(n27), .Q(o_label0_data0[21]));
Q_FDP4EP \o_label0_data0_REG[22] ( .CK(clk), .CE(n135), .R(n261), .D(n28), .Q(o_label0_data0[22]));
Q_FDP4EP \o_label0_data0_REG[23] ( .CK(clk), .CE(n135), .R(n261), .D(n29), .Q(o_label0_data0[23]));
Q_FDP4EP \o_label0_data0_REG[24] ( .CK(clk), .CE(n135), .R(n261), .D(n30), .Q(o_label0_data0[24]));
Q_FDP4EP \o_label0_data0_REG[25] ( .CK(clk), .CE(n135), .R(n261), .D(n31), .Q(o_label0_data0[25]));
Q_FDP4EP \o_label0_data0_REG[26] ( .CK(clk), .CE(n135), .R(n261), .D(n32), .Q(o_label0_data0[26]));
Q_FDP4EP \o_label0_data0_REG[27] ( .CK(clk), .CE(n135), .R(n261), .D(n33), .Q(o_label0_data0[27]));
Q_FDP4EP \o_label0_data0_REG[28] ( .CK(clk), .CE(n135), .R(n261), .D(n34), .Q(o_label0_data0[28]));
Q_FDP4EP \o_label0_data0_REG[29] ( .CK(clk), .CE(n135), .R(n261), .D(n35), .Q(o_label0_data0[29]));
Q_FDP4EP \o_label0_data0_REG[30] ( .CK(clk), .CE(n135), .R(n261), .D(n36), .Q(o_label0_data0[30]));
Q_FDP4EP \o_label0_data0_REG[31] ( .CK(clk), .CE(n135), .R(n261), .D(n37), .Q(o_label0_data0[31]));
Q_FDP4EP \o_label0_data1_REG[0] ( .CK(clk), .CE(n134), .R(n261), .D(n6), .Q(o_label0_data1[0]));
Q_FDP4EP \o_label0_data1_REG[1] ( .CK(clk), .CE(n134), .R(n261), .D(n7), .Q(o_label0_data1[1]));
Q_FDP4EP \o_label0_data1_REG[2] ( .CK(clk), .CE(n134), .R(n261), .D(n8), .Q(o_label0_data1[2]));
Q_FDP4EP \o_label0_data1_REG[3] ( .CK(clk), .CE(n134), .R(n261), .D(n9), .Q(o_label0_data1[3]));
Q_FDP4EP \o_label0_data1_REG[4] ( .CK(clk), .CE(n134), .R(n261), .D(n10), .Q(o_label0_data1[4]));
Q_FDP4EP \o_label0_data1_REG[5] ( .CK(clk), .CE(n134), .R(n261), .D(n11), .Q(o_label0_data1[5]));
Q_FDP4EP \o_label0_data1_REG[6] ( .CK(clk), .CE(n134), .R(n261), .D(n12), .Q(o_label0_data1[6]));
Q_FDP4EP \o_label0_data1_REG[7] ( .CK(clk), .CE(n134), .R(n261), .D(n13), .Q(o_label0_data1[7]));
Q_FDP4EP \o_label0_data1_REG[8] ( .CK(clk), .CE(n134), .R(n261), .D(n14), .Q(o_label0_data1[8]));
Q_FDP4EP \o_label0_data1_REG[9] ( .CK(clk), .CE(n134), .R(n261), .D(n15), .Q(o_label0_data1[9]));
Q_FDP4EP \o_label0_data1_REG[10] ( .CK(clk), .CE(n134), .R(n261), .D(n16), .Q(o_label0_data1[10]));
Q_FDP4EP \o_label0_data1_REG[11] ( .CK(clk), .CE(n134), .R(n261), .D(n17), .Q(o_label0_data1[11]));
Q_FDP4EP \o_label0_data1_REG[12] ( .CK(clk), .CE(n134), .R(n261), .D(n18), .Q(o_label0_data1[12]));
Q_FDP4EP \o_label0_data1_REG[13] ( .CK(clk), .CE(n134), .R(n261), .D(n19), .Q(o_label0_data1[13]));
Q_FDP4EP \o_label0_data1_REG[14] ( .CK(clk), .CE(n134), .R(n261), .D(n20), .Q(o_label0_data1[14]));
Q_FDP4EP \o_label0_data1_REG[15] ( .CK(clk), .CE(n134), .R(n261), .D(n21), .Q(o_label0_data1[15]));
Q_FDP4EP \o_label0_data1_REG[16] ( .CK(clk), .CE(n134), .R(n261), .D(n22), .Q(o_label0_data1[16]));
Q_FDP4EP \o_label0_data1_REG[17] ( .CK(clk), .CE(n134), .R(n261), .D(n23), .Q(o_label0_data1[17]));
Q_FDP4EP \o_label0_data1_REG[18] ( .CK(clk), .CE(n134), .R(n261), .D(n24), .Q(o_label0_data1[18]));
Q_FDP4EP \o_label0_data1_REG[19] ( .CK(clk), .CE(n134), .R(n261), .D(n25), .Q(o_label0_data1[19]));
Q_FDP4EP \o_label0_data1_REG[20] ( .CK(clk), .CE(n134), .R(n261), .D(n26), .Q(o_label0_data1[20]));
Q_FDP4EP \o_label0_data1_REG[21] ( .CK(clk), .CE(n134), .R(n261), .D(n27), .Q(o_label0_data1[21]));
Q_FDP4EP \o_label0_data1_REG[22] ( .CK(clk), .CE(n134), .R(n261), .D(n28), .Q(o_label0_data1[22]));
Q_FDP4EP \o_label0_data1_REG[23] ( .CK(clk), .CE(n134), .R(n261), .D(n29), .Q(o_label0_data1[23]));
Q_FDP4EP \o_label0_data1_REG[24] ( .CK(clk), .CE(n134), .R(n261), .D(n30), .Q(o_label0_data1[24]));
Q_FDP4EP \o_label0_data1_REG[25] ( .CK(clk), .CE(n134), .R(n261), .D(n31), .Q(o_label0_data1[25]));
Q_FDP4EP \o_label0_data1_REG[26] ( .CK(clk), .CE(n134), .R(n261), .D(n32), .Q(o_label0_data1[26]));
Q_FDP4EP \o_label0_data1_REG[27] ( .CK(clk), .CE(n134), .R(n261), .D(n33), .Q(o_label0_data1[27]));
Q_FDP4EP \o_label0_data1_REG[28] ( .CK(clk), .CE(n134), .R(n261), .D(n34), .Q(o_label0_data1[28]));
Q_FDP4EP \o_label0_data1_REG[29] ( .CK(clk), .CE(n134), .R(n261), .D(n35), .Q(o_label0_data1[29]));
Q_FDP4EP \o_label0_data1_REG[30] ( .CK(clk), .CE(n134), .R(n261), .D(n36), .Q(o_label0_data1[30]));
Q_FDP4EP \o_label0_data1_REG[31] ( .CK(clk), .CE(n134), .R(n261), .D(n37), .Q(o_label0_data1[31]));
Q_FDP4EP \o_label0_data2_REG[0] ( .CK(clk), .CE(n133), .R(n261), .D(n6), .Q(o_label0_data2[0]));
Q_FDP4EP \o_label0_data2_REG[1] ( .CK(clk), .CE(n133), .R(n261), .D(n7), .Q(o_label0_data2[1]));
Q_FDP4EP \o_label0_data2_REG[2] ( .CK(clk), .CE(n133), .R(n261), .D(n8), .Q(o_label0_data2[2]));
Q_FDP4EP \o_label0_data2_REG[3] ( .CK(clk), .CE(n133), .R(n261), .D(n9), .Q(o_label0_data2[3]));
Q_FDP4EP \o_label0_data2_REG[4] ( .CK(clk), .CE(n133), .R(n261), .D(n10), .Q(o_label0_data2[4]));
Q_FDP4EP \o_label0_data2_REG[5] ( .CK(clk), .CE(n133), .R(n261), .D(n11), .Q(o_label0_data2[5]));
Q_FDP4EP \o_label0_data2_REG[6] ( .CK(clk), .CE(n133), .R(n261), .D(n12), .Q(o_label0_data2[6]));
Q_FDP4EP \o_label0_data2_REG[7] ( .CK(clk), .CE(n133), .R(n261), .D(n13), .Q(o_label0_data2[7]));
Q_FDP4EP \o_label0_data2_REG[8] ( .CK(clk), .CE(n133), .R(n261), .D(n14), .Q(o_label0_data2[8]));
Q_FDP4EP \o_label0_data2_REG[9] ( .CK(clk), .CE(n133), .R(n261), .D(n15), .Q(o_label0_data2[9]));
Q_FDP4EP \o_label0_data2_REG[10] ( .CK(clk), .CE(n133), .R(n261), .D(n16), .Q(o_label0_data2[10]));
Q_FDP4EP \o_label0_data2_REG[11] ( .CK(clk), .CE(n133), .R(n261), .D(n17), .Q(o_label0_data2[11]));
Q_FDP4EP \o_label0_data2_REG[12] ( .CK(clk), .CE(n133), .R(n261), .D(n18), .Q(o_label0_data2[12]));
Q_FDP4EP \o_label0_data2_REG[13] ( .CK(clk), .CE(n133), .R(n261), .D(n19), .Q(o_label0_data2[13]));
Q_FDP4EP \o_label0_data2_REG[14] ( .CK(clk), .CE(n133), .R(n261), .D(n20), .Q(o_label0_data2[14]));
Q_FDP4EP \o_label0_data2_REG[15] ( .CK(clk), .CE(n133), .R(n261), .D(n21), .Q(o_label0_data2[15]));
Q_FDP4EP \o_label0_data2_REG[16] ( .CK(clk), .CE(n133), .R(n261), .D(n22), .Q(o_label0_data2[16]));
Q_FDP4EP \o_label0_data2_REG[17] ( .CK(clk), .CE(n133), .R(n261), .D(n23), .Q(o_label0_data2[17]));
Q_FDP4EP \o_label0_data2_REG[18] ( .CK(clk), .CE(n133), .R(n261), .D(n24), .Q(o_label0_data2[18]));
Q_FDP4EP \o_label0_data2_REG[19] ( .CK(clk), .CE(n133), .R(n261), .D(n25), .Q(o_label0_data2[19]));
Q_FDP4EP \o_label0_data2_REG[20] ( .CK(clk), .CE(n133), .R(n261), .D(n26), .Q(o_label0_data2[20]));
Q_FDP4EP \o_label0_data2_REG[21] ( .CK(clk), .CE(n133), .R(n261), .D(n27), .Q(o_label0_data2[21]));
Q_FDP4EP \o_label0_data2_REG[22] ( .CK(clk), .CE(n133), .R(n261), .D(n28), .Q(o_label0_data2[22]));
Q_FDP4EP \o_label0_data2_REG[23] ( .CK(clk), .CE(n133), .R(n261), .D(n29), .Q(o_label0_data2[23]));
Q_FDP4EP \o_label0_data2_REG[24] ( .CK(clk), .CE(n133), .R(n261), .D(n30), .Q(o_label0_data2[24]));
Q_FDP4EP \o_label0_data2_REG[25] ( .CK(clk), .CE(n133), .R(n261), .D(n31), .Q(o_label0_data2[25]));
Q_FDP4EP \o_label0_data2_REG[26] ( .CK(clk), .CE(n133), .R(n261), .D(n32), .Q(o_label0_data2[26]));
Q_FDP4EP \o_label0_data2_REG[27] ( .CK(clk), .CE(n133), .R(n261), .D(n33), .Q(o_label0_data2[27]));
Q_FDP4EP \o_label0_data2_REG[28] ( .CK(clk), .CE(n133), .R(n261), .D(n34), .Q(o_label0_data2[28]));
Q_FDP4EP \o_label0_data2_REG[29] ( .CK(clk), .CE(n133), .R(n261), .D(n35), .Q(o_label0_data2[29]));
Q_FDP4EP \o_label0_data2_REG[30] ( .CK(clk), .CE(n133), .R(n261), .D(n36), .Q(o_label0_data2[30]));
Q_FDP4EP \o_label0_data2_REG[31] ( .CK(clk), .CE(n133), .R(n261), .D(n37), .Q(o_label0_data2[31]));
Q_FDP4EP \o_label0_data3_REG[0] ( .CK(clk), .CE(n132), .R(n261), .D(n6), .Q(o_label0_data3[0]));
Q_FDP4EP \o_label0_data3_REG[1] ( .CK(clk), .CE(n132), .R(n261), .D(n7), .Q(o_label0_data3[1]));
Q_FDP4EP \o_label0_data3_REG[2] ( .CK(clk), .CE(n132), .R(n261), .D(n8), .Q(o_label0_data3[2]));
Q_FDP4EP \o_label0_data3_REG[3] ( .CK(clk), .CE(n132), .R(n261), .D(n9), .Q(o_label0_data3[3]));
Q_FDP4EP \o_label0_data3_REG[4] ( .CK(clk), .CE(n132), .R(n261), .D(n10), .Q(o_label0_data3[4]));
Q_FDP4EP \o_label0_data3_REG[5] ( .CK(clk), .CE(n132), .R(n261), .D(n11), .Q(o_label0_data3[5]));
Q_FDP4EP \o_label0_data3_REG[6] ( .CK(clk), .CE(n132), .R(n261), .D(n12), .Q(o_label0_data3[6]));
Q_FDP4EP \o_label0_data3_REG[7] ( .CK(clk), .CE(n132), .R(n261), .D(n13), .Q(o_label0_data3[7]));
Q_FDP4EP \o_label0_data3_REG[8] ( .CK(clk), .CE(n132), .R(n261), .D(n14), .Q(o_label0_data3[8]));
Q_FDP4EP \o_label0_data3_REG[9] ( .CK(clk), .CE(n132), .R(n261), .D(n15), .Q(o_label0_data3[9]));
Q_FDP4EP \o_label0_data3_REG[10] ( .CK(clk), .CE(n132), .R(n261), .D(n16), .Q(o_label0_data3[10]));
Q_FDP4EP \o_label0_data3_REG[11] ( .CK(clk), .CE(n132), .R(n261), .D(n17), .Q(o_label0_data3[11]));
Q_FDP4EP \o_label0_data3_REG[12] ( .CK(clk), .CE(n132), .R(n261), .D(n18), .Q(o_label0_data3[12]));
Q_FDP4EP \o_label0_data3_REG[13] ( .CK(clk), .CE(n132), .R(n261), .D(n19), .Q(o_label0_data3[13]));
Q_FDP4EP \o_label0_data3_REG[14] ( .CK(clk), .CE(n132), .R(n261), .D(n20), .Q(o_label0_data3[14]));
Q_FDP4EP \o_label0_data3_REG[15] ( .CK(clk), .CE(n132), .R(n261), .D(n21), .Q(o_label0_data3[15]));
Q_FDP4EP \o_label0_data3_REG[16] ( .CK(clk), .CE(n132), .R(n261), .D(n22), .Q(o_label0_data3[16]));
Q_FDP4EP \o_label0_data3_REG[17] ( .CK(clk), .CE(n132), .R(n261), .D(n23), .Q(o_label0_data3[17]));
Q_FDP4EP \o_label0_data3_REG[18] ( .CK(clk), .CE(n132), .R(n261), .D(n24), .Q(o_label0_data3[18]));
Q_FDP4EP \o_label0_data3_REG[19] ( .CK(clk), .CE(n132), .R(n261), .D(n25), .Q(o_label0_data3[19]));
Q_FDP4EP \o_label0_data3_REG[20] ( .CK(clk), .CE(n132), .R(n261), .D(n26), .Q(o_label0_data3[20]));
Q_FDP4EP \o_label0_data3_REG[21] ( .CK(clk), .CE(n132), .R(n261), .D(n27), .Q(o_label0_data3[21]));
Q_FDP4EP \o_label0_data3_REG[22] ( .CK(clk), .CE(n132), .R(n261), .D(n28), .Q(o_label0_data3[22]));
Q_FDP4EP \o_label0_data3_REG[23] ( .CK(clk), .CE(n132), .R(n261), .D(n29), .Q(o_label0_data3[23]));
Q_FDP4EP \o_label0_data3_REG[24] ( .CK(clk), .CE(n132), .R(n261), .D(n30), .Q(o_label0_data3[24]));
Q_FDP4EP \o_label0_data3_REG[25] ( .CK(clk), .CE(n132), .R(n261), .D(n31), .Q(o_label0_data3[25]));
Q_FDP4EP \o_label0_data3_REG[26] ( .CK(clk), .CE(n132), .R(n261), .D(n32), .Q(o_label0_data3[26]));
Q_FDP4EP \o_label0_data3_REG[27] ( .CK(clk), .CE(n132), .R(n261), .D(n33), .Q(o_label0_data3[27]));
Q_FDP4EP \o_label0_data3_REG[28] ( .CK(clk), .CE(n132), .R(n261), .D(n34), .Q(o_label0_data3[28]));
Q_FDP4EP \o_label0_data3_REG[29] ( .CK(clk), .CE(n132), .R(n261), .D(n35), .Q(o_label0_data3[29]));
Q_FDP4EP \o_label0_data3_REG[30] ( .CK(clk), .CE(n132), .R(n261), .D(n36), .Q(o_label0_data3[30]));
Q_FDP4EP \o_label0_data3_REG[31] ( .CK(clk), .CE(n132), .R(n261), .D(n37), .Q(o_label0_data3[31]));
Q_FDP4EP \o_label0_data4_REG[0] ( .CK(clk), .CE(n131), .R(n261), .D(n6), .Q(o_label0_data4[0]));
Q_FDP4EP \o_label0_data4_REG[1] ( .CK(clk), .CE(n131), .R(n261), .D(n7), .Q(o_label0_data4[1]));
Q_FDP4EP \o_label0_data4_REG[2] ( .CK(clk), .CE(n131), .R(n261), .D(n8), .Q(o_label0_data4[2]));
Q_FDP4EP \o_label0_data4_REG[3] ( .CK(clk), .CE(n131), .R(n261), .D(n9), .Q(o_label0_data4[3]));
Q_FDP4EP \o_label0_data4_REG[4] ( .CK(clk), .CE(n131), .R(n261), .D(n10), .Q(o_label0_data4[4]));
Q_FDP4EP \o_label0_data4_REG[5] ( .CK(clk), .CE(n131), .R(n261), .D(n11), .Q(o_label0_data4[5]));
Q_FDP4EP \o_label0_data4_REG[6] ( .CK(clk), .CE(n131), .R(n261), .D(n12), .Q(o_label0_data4[6]));
Q_FDP4EP \o_label0_data4_REG[7] ( .CK(clk), .CE(n131), .R(n261), .D(n13), .Q(o_label0_data4[7]));
Q_FDP4EP \o_label0_data4_REG[8] ( .CK(clk), .CE(n131), .R(n261), .D(n14), .Q(o_label0_data4[8]));
Q_FDP4EP \o_label0_data4_REG[9] ( .CK(clk), .CE(n131), .R(n261), .D(n15), .Q(o_label0_data4[9]));
Q_FDP4EP \o_label0_data4_REG[10] ( .CK(clk), .CE(n131), .R(n261), .D(n16), .Q(o_label0_data4[10]));
Q_FDP4EP \o_label0_data4_REG[11] ( .CK(clk), .CE(n131), .R(n261), .D(n17), .Q(o_label0_data4[11]));
Q_FDP4EP \o_label0_data4_REG[12] ( .CK(clk), .CE(n131), .R(n261), .D(n18), .Q(o_label0_data4[12]));
Q_FDP4EP \o_label0_data4_REG[13] ( .CK(clk), .CE(n131), .R(n261), .D(n19), .Q(o_label0_data4[13]));
Q_FDP4EP \o_label0_data4_REG[14] ( .CK(clk), .CE(n131), .R(n261), .D(n20), .Q(o_label0_data4[14]));
Q_FDP4EP \o_label0_data4_REG[15] ( .CK(clk), .CE(n131), .R(n261), .D(n21), .Q(o_label0_data4[15]));
Q_FDP4EP \o_label0_data4_REG[16] ( .CK(clk), .CE(n131), .R(n261), .D(n22), .Q(o_label0_data4[16]));
Q_FDP4EP \o_label0_data4_REG[17] ( .CK(clk), .CE(n131), .R(n261), .D(n23), .Q(o_label0_data4[17]));
Q_FDP4EP \o_label0_data4_REG[18] ( .CK(clk), .CE(n131), .R(n261), .D(n24), .Q(o_label0_data4[18]));
Q_FDP4EP \o_label0_data4_REG[19] ( .CK(clk), .CE(n131), .R(n261), .D(n25), .Q(o_label0_data4[19]));
Q_FDP4EP \o_label0_data4_REG[20] ( .CK(clk), .CE(n131), .R(n261), .D(n26), .Q(o_label0_data4[20]));
Q_FDP4EP \o_label0_data4_REG[21] ( .CK(clk), .CE(n131), .R(n261), .D(n27), .Q(o_label0_data4[21]));
Q_FDP4EP \o_label0_data4_REG[22] ( .CK(clk), .CE(n131), .R(n261), .D(n28), .Q(o_label0_data4[22]));
Q_FDP4EP \o_label0_data4_REG[23] ( .CK(clk), .CE(n131), .R(n261), .D(n29), .Q(o_label0_data4[23]));
Q_FDP4EP \o_label0_data4_REG[24] ( .CK(clk), .CE(n131), .R(n261), .D(n30), .Q(o_label0_data4[24]));
Q_FDP4EP \o_label0_data4_REG[25] ( .CK(clk), .CE(n131), .R(n261), .D(n31), .Q(o_label0_data4[25]));
Q_FDP4EP \o_label0_data4_REG[26] ( .CK(clk), .CE(n131), .R(n261), .D(n32), .Q(o_label0_data4[26]));
Q_FDP4EP \o_label0_data4_REG[27] ( .CK(clk), .CE(n131), .R(n261), .D(n33), .Q(o_label0_data4[27]));
Q_FDP4EP \o_label0_data4_REG[28] ( .CK(clk), .CE(n131), .R(n261), .D(n34), .Q(o_label0_data4[28]));
Q_FDP4EP \o_label0_data4_REG[29] ( .CK(clk), .CE(n131), .R(n261), .D(n35), .Q(o_label0_data4[29]));
Q_FDP4EP \o_label0_data4_REG[30] ( .CK(clk), .CE(n131), .R(n261), .D(n36), .Q(o_label0_data4[30]));
Q_FDP4EP \o_label0_data4_REG[31] ( .CK(clk), .CE(n131), .R(n261), .D(n37), .Q(o_label0_data4[31]));
Q_FDP4EP \o_label0_data5_REG[0] ( .CK(clk), .CE(n130), .R(n261), .D(n6), .Q(o_label0_data5[0]));
Q_FDP4EP \o_label0_data5_REG[1] ( .CK(clk), .CE(n130), .R(n261), .D(n7), .Q(o_label0_data5[1]));
Q_FDP4EP \o_label0_data5_REG[2] ( .CK(clk), .CE(n130), .R(n261), .D(n8), .Q(o_label0_data5[2]));
Q_FDP4EP \o_label0_data5_REG[3] ( .CK(clk), .CE(n130), .R(n261), .D(n9), .Q(o_label0_data5[3]));
Q_FDP4EP \o_label0_data5_REG[4] ( .CK(clk), .CE(n130), .R(n261), .D(n10), .Q(o_label0_data5[4]));
Q_FDP4EP \o_label0_data5_REG[5] ( .CK(clk), .CE(n130), .R(n261), .D(n11), .Q(o_label0_data5[5]));
Q_FDP4EP \o_label0_data5_REG[6] ( .CK(clk), .CE(n130), .R(n261), .D(n12), .Q(o_label0_data5[6]));
Q_FDP4EP \o_label0_data5_REG[7] ( .CK(clk), .CE(n130), .R(n261), .D(n13), .Q(o_label0_data5[7]));
Q_FDP4EP \o_label0_data5_REG[8] ( .CK(clk), .CE(n130), .R(n261), .D(n14), .Q(o_label0_data5[8]));
Q_FDP4EP \o_label0_data5_REG[9] ( .CK(clk), .CE(n130), .R(n261), .D(n15), .Q(o_label0_data5[9]));
Q_FDP4EP \o_label0_data5_REG[10] ( .CK(clk), .CE(n130), .R(n261), .D(n16), .Q(o_label0_data5[10]));
Q_FDP4EP \o_label0_data5_REG[11] ( .CK(clk), .CE(n130), .R(n261), .D(n17), .Q(o_label0_data5[11]));
Q_FDP4EP \o_label0_data5_REG[12] ( .CK(clk), .CE(n130), .R(n261), .D(n18), .Q(o_label0_data5[12]));
Q_FDP4EP \o_label0_data5_REG[13] ( .CK(clk), .CE(n130), .R(n261), .D(n19), .Q(o_label0_data5[13]));
Q_FDP4EP \o_label0_data5_REG[14] ( .CK(clk), .CE(n130), .R(n261), .D(n20), .Q(o_label0_data5[14]));
Q_FDP4EP \o_label0_data5_REG[15] ( .CK(clk), .CE(n130), .R(n261), .D(n21), .Q(o_label0_data5[15]));
Q_FDP4EP \o_label0_data5_REG[16] ( .CK(clk), .CE(n130), .R(n261), .D(n22), .Q(o_label0_data5[16]));
Q_FDP4EP \o_label0_data5_REG[17] ( .CK(clk), .CE(n130), .R(n261), .D(n23), .Q(o_label0_data5[17]));
Q_FDP4EP \o_label0_data5_REG[18] ( .CK(clk), .CE(n130), .R(n261), .D(n24), .Q(o_label0_data5[18]));
Q_FDP4EP \o_label0_data5_REG[19] ( .CK(clk), .CE(n130), .R(n261), .D(n25), .Q(o_label0_data5[19]));
Q_FDP4EP \o_label0_data5_REG[20] ( .CK(clk), .CE(n130), .R(n261), .D(n26), .Q(o_label0_data5[20]));
Q_FDP4EP \o_label0_data5_REG[21] ( .CK(clk), .CE(n130), .R(n261), .D(n27), .Q(o_label0_data5[21]));
Q_FDP4EP \o_label0_data5_REG[22] ( .CK(clk), .CE(n130), .R(n261), .D(n28), .Q(o_label0_data5[22]));
Q_FDP4EP \o_label0_data5_REG[23] ( .CK(clk), .CE(n130), .R(n261), .D(n29), .Q(o_label0_data5[23]));
Q_FDP4EP \o_label0_data5_REG[24] ( .CK(clk), .CE(n130), .R(n261), .D(n30), .Q(o_label0_data5[24]));
Q_FDP4EP \o_label0_data5_REG[25] ( .CK(clk), .CE(n130), .R(n261), .D(n31), .Q(o_label0_data5[25]));
Q_FDP4EP \o_label0_data5_REG[26] ( .CK(clk), .CE(n130), .R(n261), .D(n32), .Q(o_label0_data5[26]));
Q_FDP4EP \o_label0_data5_REG[27] ( .CK(clk), .CE(n130), .R(n261), .D(n33), .Q(o_label0_data5[27]));
Q_FDP4EP \o_label0_data5_REG[28] ( .CK(clk), .CE(n130), .R(n261), .D(n34), .Q(o_label0_data5[28]));
Q_FDP4EP \o_label0_data5_REG[29] ( .CK(clk), .CE(n130), .R(n261), .D(n35), .Q(o_label0_data5[29]));
Q_FDP4EP \o_label0_data5_REG[30] ( .CK(clk), .CE(n130), .R(n261), .D(n36), .Q(o_label0_data5[30]));
Q_FDP4EP \o_label0_data5_REG[31] ( .CK(clk), .CE(n130), .R(n261), .D(n37), .Q(o_label0_data5[31]));
Q_FDP4EP \o_label0_data6_REG[0] ( .CK(clk), .CE(n129), .R(n261), .D(n6), .Q(o_label0_data6[0]));
Q_FDP4EP \o_label0_data6_REG[1] ( .CK(clk), .CE(n129), .R(n261), .D(n7), .Q(o_label0_data6[1]));
Q_FDP4EP \o_label0_data6_REG[2] ( .CK(clk), .CE(n129), .R(n261), .D(n8), .Q(o_label0_data6[2]));
Q_FDP4EP \o_label0_data6_REG[3] ( .CK(clk), .CE(n129), .R(n261), .D(n9), .Q(o_label0_data6[3]));
Q_FDP4EP \o_label0_data6_REG[4] ( .CK(clk), .CE(n129), .R(n261), .D(n10), .Q(o_label0_data6[4]));
Q_FDP4EP \o_label0_data6_REG[5] ( .CK(clk), .CE(n129), .R(n261), .D(n11), .Q(o_label0_data6[5]));
Q_FDP4EP \o_label0_data6_REG[6] ( .CK(clk), .CE(n129), .R(n261), .D(n12), .Q(o_label0_data6[6]));
Q_FDP4EP \o_label0_data6_REG[7] ( .CK(clk), .CE(n129), .R(n261), .D(n13), .Q(o_label0_data6[7]));
Q_FDP4EP \o_label0_data6_REG[8] ( .CK(clk), .CE(n129), .R(n261), .D(n14), .Q(o_label0_data6[8]));
Q_FDP4EP \o_label0_data6_REG[9] ( .CK(clk), .CE(n129), .R(n261), .D(n15), .Q(o_label0_data6[9]));
Q_FDP4EP \o_label0_data6_REG[10] ( .CK(clk), .CE(n129), .R(n261), .D(n16), .Q(o_label0_data6[10]));
Q_FDP4EP \o_label0_data6_REG[11] ( .CK(clk), .CE(n129), .R(n261), .D(n17), .Q(o_label0_data6[11]));
Q_FDP4EP \o_label0_data6_REG[12] ( .CK(clk), .CE(n129), .R(n261), .D(n18), .Q(o_label0_data6[12]));
Q_FDP4EP \o_label0_data6_REG[13] ( .CK(clk), .CE(n129), .R(n261), .D(n19), .Q(o_label0_data6[13]));
Q_FDP4EP \o_label0_data6_REG[14] ( .CK(clk), .CE(n129), .R(n261), .D(n20), .Q(o_label0_data6[14]));
Q_FDP4EP \o_label0_data6_REG[15] ( .CK(clk), .CE(n129), .R(n261), .D(n21), .Q(o_label0_data6[15]));
Q_FDP4EP \o_label0_data6_REG[16] ( .CK(clk), .CE(n129), .R(n261), .D(n22), .Q(o_label0_data6[16]));
Q_FDP4EP \o_label0_data6_REG[17] ( .CK(clk), .CE(n129), .R(n261), .D(n23), .Q(o_label0_data6[17]));
Q_FDP4EP \o_label0_data6_REG[18] ( .CK(clk), .CE(n129), .R(n261), .D(n24), .Q(o_label0_data6[18]));
Q_FDP4EP \o_label0_data6_REG[19] ( .CK(clk), .CE(n129), .R(n261), .D(n25), .Q(o_label0_data6[19]));
Q_FDP4EP \o_label0_data6_REG[20] ( .CK(clk), .CE(n129), .R(n261), .D(n26), .Q(o_label0_data6[20]));
Q_FDP4EP \o_label0_data6_REG[21] ( .CK(clk), .CE(n129), .R(n261), .D(n27), .Q(o_label0_data6[21]));
Q_FDP4EP \o_label0_data6_REG[22] ( .CK(clk), .CE(n129), .R(n261), .D(n28), .Q(o_label0_data6[22]));
Q_FDP4EP \o_label0_data6_REG[23] ( .CK(clk), .CE(n129), .R(n261), .D(n29), .Q(o_label0_data6[23]));
Q_FDP4EP \o_label0_data6_REG[24] ( .CK(clk), .CE(n129), .R(n261), .D(n30), .Q(o_label0_data6[24]));
Q_FDP4EP \o_label0_data6_REG[25] ( .CK(clk), .CE(n129), .R(n261), .D(n31), .Q(o_label0_data6[25]));
Q_FDP4EP \o_label0_data6_REG[26] ( .CK(clk), .CE(n129), .R(n261), .D(n32), .Q(o_label0_data6[26]));
Q_FDP4EP \o_label0_data6_REG[27] ( .CK(clk), .CE(n129), .R(n261), .D(n33), .Q(o_label0_data6[27]));
Q_FDP4EP \o_label0_data6_REG[28] ( .CK(clk), .CE(n129), .R(n261), .D(n34), .Q(o_label0_data6[28]));
Q_FDP4EP \o_label0_data6_REG[29] ( .CK(clk), .CE(n129), .R(n261), .D(n35), .Q(o_label0_data6[29]));
Q_FDP4EP \o_label0_data6_REG[30] ( .CK(clk), .CE(n129), .R(n261), .D(n36), .Q(o_label0_data6[30]));
Q_FDP4EP \o_label0_data6_REG[31] ( .CK(clk), .CE(n129), .R(n261), .D(n37), .Q(o_label0_data6[31]));
Q_FDP4EP \o_label0_data7_REG[0] ( .CK(clk), .CE(n128), .R(n261), .D(n6), .Q(o_label0_data7[0]));
Q_FDP4EP \o_label0_data7_REG[1] ( .CK(clk), .CE(n128), .R(n261), .D(n7), .Q(o_label0_data7[1]));
Q_FDP4EP \o_label0_data7_REG[2] ( .CK(clk), .CE(n128), .R(n261), .D(n8), .Q(o_label0_data7[2]));
Q_FDP4EP \o_label0_data7_REG[3] ( .CK(clk), .CE(n128), .R(n261), .D(n9), .Q(o_label0_data7[3]));
Q_FDP4EP \o_label0_data7_REG[4] ( .CK(clk), .CE(n128), .R(n261), .D(n10), .Q(o_label0_data7[4]));
Q_FDP4EP \o_label0_data7_REG[5] ( .CK(clk), .CE(n128), .R(n261), .D(n11), .Q(o_label0_data7[5]));
Q_FDP4EP \o_label0_data7_REG[6] ( .CK(clk), .CE(n128), .R(n261), .D(n12), .Q(o_label0_data7[6]));
Q_FDP4EP \o_label0_data7_REG[7] ( .CK(clk), .CE(n128), .R(n261), .D(n13), .Q(o_label0_data7[7]));
Q_FDP4EP \o_label0_data7_REG[8] ( .CK(clk), .CE(n128), .R(n261), .D(n14), .Q(o_label0_data7[8]));
Q_FDP4EP \o_label0_data7_REG[9] ( .CK(clk), .CE(n128), .R(n261), .D(n15), .Q(o_label0_data7[9]));
Q_FDP4EP \o_label0_data7_REG[10] ( .CK(clk), .CE(n128), .R(n261), .D(n16), .Q(o_label0_data7[10]));
Q_FDP4EP \o_label0_data7_REG[11] ( .CK(clk), .CE(n128), .R(n261), .D(n17), .Q(o_label0_data7[11]));
Q_FDP4EP \o_label0_data7_REG[12] ( .CK(clk), .CE(n128), .R(n261), .D(n18), .Q(o_label0_data7[12]));
Q_FDP4EP \o_label0_data7_REG[13] ( .CK(clk), .CE(n128), .R(n261), .D(n19), .Q(o_label0_data7[13]));
Q_FDP4EP \o_label0_data7_REG[14] ( .CK(clk), .CE(n128), .R(n261), .D(n20), .Q(o_label0_data7[14]));
Q_FDP4EP \o_label0_data7_REG[15] ( .CK(clk), .CE(n128), .R(n261), .D(n21), .Q(o_label0_data7[15]));
Q_FDP4EP \o_label0_data7_REG[16] ( .CK(clk), .CE(n128), .R(n261), .D(n22), .Q(o_label0_data7[16]));
Q_FDP4EP \o_label0_data7_REG[17] ( .CK(clk), .CE(n128), .R(n261), .D(n23), .Q(o_label0_data7[17]));
Q_FDP4EP \o_label0_data7_REG[18] ( .CK(clk), .CE(n128), .R(n261), .D(n24), .Q(o_label0_data7[18]));
Q_FDP4EP \o_label0_data7_REG[19] ( .CK(clk), .CE(n128), .R(n261), .D(n25), .Q(o_label0_data7[19]));
Q_FDP4EP \o_label0_data7_REG[20] ( .CK(clk), .CE(n128), .R(n261), .D(n26), .Q(o_label0_data7[20]));
Q_FDP4EP \o_label0_data7_REG[21] ( .CK(clk), .CE(n128), .R(n261), .D(n27), .Q(o_label0_data7[21]));
Q_FDP4EP \o_label0_data7_REG[22] ( .CK(clk), .CE(n128), .R(n261), .D(n28), .Q(o_label0_data7[22]));
Q_FDP4EP \o_label0_data7_REG[23] ( .CK(clk), .CE(n128), .R(n261), .D(n29), .Q(o_label0_data7[23]));
Q_FDP4EP \o_label0_data7_REG[24] ( .CK(clk), .CE(n128), .R(n261), .D(n30), .Q(o_label0_data7[24]));
Q_FDP4EP \o_label0_data7_REG[25] ( .CK(clk), .CE(n128), .R(n261), .D(n31), .Q(o_label0_data7[25]));
Q_FDP4EP \o_label0_data7_REG[26] ( .CK(clk), .CE(n128), .R(n261), .D(n32), .Q(o_label0_data7[26]));
Q_FDP4EP \o_label0_data7_REG[27] ( .CK(clk), .CE(n128), .R(n261), .D(n33), .Q(o_label0_data7[27]));
Q_FDP4EP \o_label0_data7_REG[28] ( .CK(clk), .CE(n128), .R(n261), .D(n34), .Q(o_label0_data7[28]));
Q_FDP4EP \o_label0_data7_REG[29] ( .CK(clk), .CE(n128), .R(n261), .D(n35), .Q(o_label0_data7[29]));
Q_FDP4EP \o_label0_data7_REG[30] ( .CK(clk), .CE(n128), .R(n261), .D(n36), .Q(o_label0_data7[30]));
Q_FDP4EP \o_label0_data7_REG[31] ( .CK(clk), .CE(n128), .R(n261), .D(n37), .Q(o_label0_data7[31]));
Q_FDP4EP \o_label0_config_REG[0] ( .CK(clk), .CE(n127), .R(n261), .D(n6), .Q(o_label0_config[0]));
Q_FDP4EP \o_label0_config_REG[1] ( .CK(clk), .CE(n127), .R(n261), .D(n7), .Q(o_label0_config[1]));
Q_FDP4EP \o_label0_config_REG[2] ( .CK(clk), .CE(n127), .R(n261), .D(n8), .Q(o_label0_config[2]));
Q_FDP4EP \o_label0_config_REG[3] ( .CK(clk), .CE(n127), .R(n261), .D(n9), .Q(o_label0_config[3]));
Q_FDP4EP \o_label0_config_REG[4] ( .CK(clk), .CE(n127), .R(n261), .D(n10), .Q(o_label0_config[4]));
Q_FDP4EP \o_label0_config_REG[5] ( .CK(clk), .CE(n127), .R(n261), .D(n11), .Q(o_label0_config[5]));
Q_FDP4EP \o_label0_config_REG[6] ( .CK(clk), .CE(n127), .R(n261), .D(n12), .Q(o_label0_config[6]));
Q_FDP4EP \o_label0_config_REG[7] ( .CK(clk), .CE(n127), .R(n261), .D(n13), .Q(o_label0_config[7]));
Q_FDP4EP \o_label0_config_REG[9] ( .CK(clk), .CE(n127), .R(n261), .D(n31), .Q(o_label0_config[9]));
Q_FDP4EP \o_label0_config_REG[10] ( .CK(clk), .CE(n127), .R(n261), .D(n32), .Q(o_label0_config[10]));
Q_FDP4EP \o_label0_config_REG[11] ( .CK(clk), .CE(n127), .R(n261), .D(n33), .Q(o_label0_config[11]));
Q_FDP4EP \o_label0_config_REG[12] ( .CK(clk), .CE(n127), .R(n261), .D(n34), .Q(o_label0_config[12]));
Q_FDP4EP \o_label0_config_REG[13] ( .CK(clk), .CE(n127), .R(n261), .D(n35), .Q(o_label0_config[13]));
Q_FDP4EP \o_label0_config_REG[14] ( .CK(clk), .CE(n127), .R(n261), .D(n36), .Q(o_label0_config[14]));
Q_FDP4EP \o_label0_config_REG[15] ( .CK(clk), .CE(n127), .R(n261), .D(n37), .Q(o_label0_config[15]));
Q_FDP4EP \o_kim_ia_config_REG[0] ( .CK(clk), .CE(n126), .R(n261), .D(n6), .Q(o_kim_ia_config[0]));
Q_FDP4EP \o_kim_ia_config_REG[1] ( .CK(clk), .CE(n126), .R(n261), .D(n7), .Q(o_kim_ia_config[1]));
Q_FDP4EP \o_kim_ia_config_REG[2] ( .CK(clk), .CE(n126), .R(n261), .D(n8), .Q(o_kim_ia_config[2]));
Q_FDP4EP \o_kim_ia_config_REG[3] ( .CK(clk), .CE(n126), .R(n261), .D(n9), .Q(o_kim_ia_config[3]));
Q_FDP4EP \o_kim_ia_config_REG[4] ( .CK(clk), .CE(n126), .R(n261), .D(n10), .Q(o_kim_ia_config[4]));
Q_FDP4EP \o_kim_ia_config_REG[5] ( .CK(clk), .CE(n126), .R(n261), .D(n11), .Q(o_kim_ia_config[5]));
Q_FDP4EP \o_kim_ia_config_REG[6] ( .CK(clk), .CE(n126), .R(n261), .D(n12), .Q(o_kim_ia_config[6]));
Q_FDP4EP \o_kim_ia_config_REG[7] ( .CK(clk), .CE(n126), .R(n261), .D(n13), .Q(o_kim_ia_config[7]));
Q_FDP4EP \o_kim_ia_config_REG[8] ( .CK(clk), .CE(n126), .R(n261), .D(n14), .Q(o_kim_ia_config[8]));
Q_FDP4EP \o_kim_ia_config_REG[9] ( .CK(clk), .CE(n126), .R(n261), .D(n15), .Q(o_kim_ia_config[9]));
Q_FDP4EP \o_kim_ia_config_REG[10] ( .CK(clk), .CE(n126), .R(n261), .D(n16), .Q(o_kim_ia_config[10]));
Q_FDP4EP \o_kim_ia_config_REG[11] ( .CK(clk), .CE(n126), .R(n261), .D(n17), .Q(o_kim_ia_config[11]));
Q_FDP4EP \o_kim_ia_config_REG[12] ( .CK(clk), .CE(n126), .R(n261), .D(n18), .Q(o_kim_ia_config[12]));
Q_FDP4EP \o_kim_ia_config_REG[13] ( .CK(clk), .CE(n126), .R(n261), .D(n19), .Q(o_kim_ia_config[13]));
Q_FDP4EP \o_kim_ia_config_REG[14] ( .CK(clk), .CE(n126), .R(n261), .D(n34), .Q(o_kim_ia_config[14]));
Q_FDP4EP \o_kim_ia_config_REG[15] ( .CK(clk), .CE(n126), .R(n261), .D(n35), .Q(o_kim_ia_config[15]));
Q_FDP4EP \o_kim_ia_config_REG[16] ( .CK(clk), .CE(n126), .R(n261), .D(n36), .Q(o_kim_ia_config[16]));
Q_FDP4EP \o_kim_ia_config_REG[17] ( .CK(clk), .CE(n126), .R(n261), .D(n37), .Q(o_kim_ia_config[17]));
Q_FDP4EP \o_kim_ia_wdata_part1_REG[0] ( .CK(clk), .CE(n125), .R(n261), .D(n6), .Q(o_kim_ia_wdata_part1[0]));
Q_FDP4EP \o_kim_ia_wdata_part1_REG[1] ( .CK(clk), .CE(n125), .R(n261), .D(n7), .Q(o_kim_ia_wdata_part1[1]));
Q_FDP4EP \o_kim_ia_wdata_part1_REG[2] ( .CK(clk), .CE(n125), .R(n261), .D(n8), .Q(o_kim_ia_wdata_part1[2]));
Q_FDP4EP \o_kim_ia_wdata_part1_REG[3] ( .CK(clk), .CE(n125), .R(n261), .D(n9), .Q(o_kim_ia_wdata_part1[3]));
Q_FDP4EP \o_kim_ia_wdata_part1_REG[4] ( .CK(clk), .CE(n125), .R(n261), .D(n10), .Q(o_kim_ia_wdata_part1[4]));
Q_FDP4EP \o_kim_ia_wdata_part1_REG[5] ( .CK(clk), .CE(n125), .R(n261), .D(n11), .Q(o_kim_ia_wdata_part1[5]));
Q_FDP4EP \o_kim_ia_wdata_part1_REG[6] ( .CK(clk), .CE(n125), .R(n261), .D(n12), .Q(o_kim_ia_wdata_part1[6]));
Q_FDP4EP \o_kim_ia_wdata_part1_REG[7] ( .CK(clk), .CE(n125), .R(n261), .D(n13), .Q(o_kim_ia_wdata_part1[7]));
Q_FDP4EP \o_kim_ia_wdata_part1_REG[8] ( .CK(clk), .CE(n125), .R(n261), .D(n14), .Q(o_kim_ia_wdata_part1[8]));
Q_FDP4EP \o_kim_ia_wdata_part1_REG[9] ( .CK(clk), .CE(n125), .R(n261), .D(n15), .Q(o_kim_ia_wdata_part1[9]));
Q_FDP4EP \o_kim_ia_wdata_part1_REG[10] ( .CK(clk), .CE(n125), .R(n261), .D(n16), .Q(o_kim_ia_wdata_part1[10]));
Q_FDP4EP \o_kim_ia_wdata_part1_REG[11] ( .CK(clk), .CE(n125), .R(n261), .D(n17), .Q(o_kim_ia_wdata_part1[11]));
Q_FDP4EP \o_kim_ia_wdata_part1_REG[12] ( .CK(clk), .CE(n125), .R(n261), .D(n18), .Q(o_kim_ia_wdata_part1[12]));
Q_FDP4EP \o_kim_ia_wdata_part1_REG[13] ( .CK(clk), .CE(n125), .R(n261), .D(n34), .Q(o_kim_ia_wdata_part1[13]));
Q_FDP4EP \o_kim_ia_wdata_part1_REG[14] ( .CK(clk), .CE(n125), .R(n261), .D(n35), .Q(o_kim_ia_wdata_part1[14]));
Q_FDP4EP \o_kim_ia_wdata_part1_REG[15] ( .CK(clk), .CE(n125), .R(n261), .D(n36), .Q(o_kim_ia_wdata_part1[15]));
Q_FDP4EP \o_kim_ia_wdata_part1_REG[16] ( .CK(clk), .CE(n125), .R(n261), .D(n37), .Q(o_kim_ia_wdata_part1[16]));
Q_FDP4EP \o_kim_ia_wdata_part0_REG[0] ( .CK(clk), .CE(n124), .R(n261), .D(n6), .Q(o_kim_ia_wdata_part0[0]));
Q_FDP4EP \o_kim_ia_wdata_part0_REG[1] ( .CK(clk), .CE(n124), .R(n261), .D(n7), .Q(o_kim_ia_wdata_part0[1]));
Q_FDP4EP \o_kim_ia_wdata_part0_REG[2] ( .CK(clk), .CE(n124), .R(n261), .D(n8), .Q(o_kim_ia_wdata_part0[2]));
Q_FDP4EP \o_kim_ia_wdata_part0_REG[3] ( .CK(clk), .CE(n124), .R(n261), .D(n9), .Q(o_kim_ia_wdata_part0[3]));
Q_FDP4EP \o_kim_ia_wdata_part0_REG[4] ( .CK(clk), .CE(n124), .R(n261), .D(n10), .Q(o_kim_ia_wdata_part0[4]));
Q_FDP4EP \o_kim_ia_wdata_part0_REG[5] ( .CK(clk), .CE(n124), .R(n261), .D(n11), .Q(o_kim_ia_wdata_part0[5]));
Q_FDP4EP \o_kim_ia_wdata_part0_REG[6] ( .CK(clk), .CE(n124), .R(n261), .D(n12), .Q(o_kim_ia_wdata_part0[6]));
Q_FDP4EP \o_kim_ia_wdata_part0_REG[7] ( .CK(clk), .CE(n124), .R(n261), .D(n13), .Q(o_kim_ia_wdata_part0[7]));
Q_FDP4EP \o_kim_ia_wdata_part0_REG[8] ( .CK(clk), .CE(n124), .R(n261), .D(n14), .Q(o_kim_ia_wdata_part0[8]));
Q_FDP4EP \o_kim_ia_wdata_part0_REG[9] ( .CK(clk), .CE(n124), .R(n261), .D(n15), .Q(o_kim_ia_wdata_part0[9]));
Q_FDP4EP \o_kim_ia_wdata_part0_REG[10] ( .CK(clk), .CE(n124), .R(n261), .D(n16), .Q(o_kim_ia_wdata_part0[10]));
Q_FDP4EP \o_kim_ia_wdata_part0_REG[11] ( .CK(clk), .CE(n124), .R(n261), .D(n17), .Q(o_kim_ia_wdata_part0[11]));
Q_FDP4EP \o_kim_ia_wdata_part0_REG[12] ( .CK(clk), .CE(n124), .R(n261), .D(n18), .Q(o_kim_ia_wdata_part0[12]));
Q_FDP4EP \o_kim_ia_wdata_part0_REG[13] ( .CK(clk), .CE(n124), .R(n261), .D(n19), .Q(o_kim_ia_wdata_part0[13]));
Q_FDP4EP \o_kim_ia_wdata_part0_REG[14] ( .CK(clk), .CE(n124), .R(n261), .D(n20), .Q(o_kim_ia_wdata_part0[14]));
Q_FDP4EP \o_kim_ia_wdata_part0_REG[15] ( .CK(clk), .CE(n124), .R(n261), .D(n32), .Q(o_kim_ia_wdata_part0[15]));
Q_FDP4EP \o_kim_ia_wdata_part0_REG[16] ( .CK(clk), .CE(n124), .R(n261), .D(n33), .Q(o_kim_ia_wdata_part0[16]));
Q_FDP4EP \o_kim_ia_wdata_part0_REG[17] ( .CK(clk), .CE(n124), .R(n261), .D(n34), .Q(o_kim_ia_wdata_part0[17]));
Q_FDP4EP \o_kim_ia_wdata_part0_REG[18] ( .CK(clk), .CE(n124), .R(n261), .D(n35), .Q(o_kim_ia_wdata_part0[18]));
Q_FDP4EP \o_kim_ia_wdata_part0_REG[19] ( .CK(clk), .CE(n124), .R(n261), .D(n36), .Q(o_kim_ia_wdata_part0[19]));
Q_FDP4EP \o_kim_ia_wdata_part0_REG[20] ( .CK(clk), .CE(n124), .R(n261), .D(n37), .Q(o_kim_ia_wdata_part0[20]));
Q_FDP4EP \o_ckv_ia_config_REG[0] ( .CK(clk), .CE(n123), .R(n261), .D(n6), .Q(o_ckv_ia_config[0]));
Q_FDP4EP \o_ckv_ia_config_REG[1] ( .CK(clk), .CE(n123), .R(n261), .D(n7), .Q(o_ckv_ia_config[1]));
Q_FDP4EP \o_ckv_ia_config_REG[2] ( .CK(clk), .CE(n123), .R(n261), .D(n8), .Q(o_ckv_ia_config[2]));
Q_FDP4EP \o_ckv_ia_config_REG[3] ( .CK(clk), .CE(n123), .R(n261), .D(n9), .Q(o_ckv_ia_config[3]));
Q_FDP4EP \o_ckv_ia_config_REG[4] ( .CK(clk), .CE(n123), .R(n261), .D(n10), .Q(o_ckv_ia_config[4]));
Q_FDP4EP \o_ckv_ia_config_REG[5] ( .CK(clk), .CE(n123), .R(n261), .D(n11), .Q(o_ckv_ia_config[5]));
Q_FDP4EP \o_ckv_ia_config_REG[6] ( .CK(clk), .CE(n123), .R(n261), .D(n12), .Q(o_ckv_ia_config[6]));
Q_FDP4EP \o_ckv_ia_config_REG[7] ( .CK(clk), .CE(n123), .R(n261), .D(n13), .Q(o_ckv_ia_config[7]));
Q_FDP4EP \o_ckv_ia_config_REG[8] ( .CK(clk), .CE(n123), .R(n261), .D(n14), .Q(o_ckv_ia_config[8]));
Q_FDP4EP \o_ckv_ia_config_REG[9] ( .CK(clk), .CE(n123), .R(n261), .D(n15), .Q(o_ckv_ia_config[9]));
Q_FDP4EP \o_ckv_ia_config_REG[10] ( .CK(clk), .CE(n123), .R(n261), .D(n16), .Q(o_ckv_ia_config[10]));
Q_FDP4EP \o_ckv_ia_config_REG[11] ( .CK(clk), .CE(n123), .R(n261), .D(n17), .Q(o_ckv_ia_config[11]));
Q_FDP4EP \o_ckv_ia_config_REG[12] ( .CK(clk), .CE(n123), .R(n261), .D(n18), .Q(o_ckv_ia_config[12]));
Q_FDP4EP \o_ckv_ia_config_REG[13] ( .CK(clk), .CE(n123), .R(n261), .D(n19), .Q(o_ckv_ia_config[13]));
Q_FDP4EP \o_ckv_ia_config_REG[14] ( .CK(clk), .CE(n123), .R(n261), .D(n20), .Q(o_ckv_ia_config[14]));
Q_FDP4EP \o_ckv_ia_config_REG[15] ( .CK(clk), .CE(n123), .R(n261), .D(n34), .Q(o_ckv_ia_config[15]));
Q_FDP4EP \o_ckv_ia_config_REG[16] ( .CK(clk), .CE(n123), .R(n261), .D(n35), .Q(o_ckv_ia_config[16]));
Q_FDP4EP \o_ckv_ia_config_REG[17] ( .CK(clk), .CE(n123), .R(n261), .D(n36), .Q(o_ckv_ia_config[17]));
Q_FDP4EP \o_ckv_ia_config_REG[18] ( .CK(clk), .CE(n123), .R(n261), .D(n37), .Q(o_ckv_ia_config[18]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[0] ( .CK(clk), .CE(n122), .R(n261), .D(n6), .Q(o_ckv_ia_wdata_part1[0]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[1] ( .CK(clk), .CE(n122), .R(n261), .D(n7), .Q(o_ckv_ia_wdata_part1[1]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[2] ( .CK(clk), .CE(n122), .R(n261), .D(n8), .Q(o_ckv_ia_wdata_part1[2]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[3] ( .CK(clk), .CE(n122), .R(n261), .D(n9), .Q(o_ckv_ia_wdata_part1[3]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[4] ( .CK(clk), .CE(n122), .R(n261), .D(n10), .Q(o_ckv_ia_wdata_part1[4]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[5] ( .CK(clk), .CE(n122), .R(n261), .D(n11), .Q(o_ckv_ia_wdata_part1[5]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[6] ( .CK(clk), .CE(n122), .R(n261), .D(n12), .Q(o_ckv_ia_wdata_part1[6]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[7] ( .CK(clk), .CE(n122), .R(n261), .D(n13), .Q(o_ckv_ia_wdata_part1[7]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[8] ( .CK(clk), .CE(n122), .R(n261), .D(n14), .Q(o_ckv_ia_wdata_part1[8]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[9] ( .CK(clk), .CE(n122), .R(n261), .D(n15), .Q(o_ckv_ia_wdata_part1[9]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[10] ( .CK(clk), .CE(n122), .R(n261), .D(n16), .Q(o_ckv_ia_wdata_part1[10]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[11] ( .CK(clk), .CE(n122), .R(n261), .D(n17), .Q(o_ckv_ia_wdata_part1[11]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[12] ( .CK(clk), .CE(n122), .R(n261), .D(n18), .Q(o_ckv_ia_wdata_part1[12]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[13] ( .CK(clk), .CE(n122), .R(n261), .D(n19), .Q(o_ckv_ia_wdata_part1[13]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[14] ( .CK(clk), .CE(n122), .R(n261), .D(n20), .Q(o_ckv_ia_wdata_part1[14]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[15] ( .CK(clk), .CE(n122), .R(n261), .D(n21), .Q(o_ckv_ia_wdata_part1[15]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[16] ( .CK(clk), .CE(n122), .R(n261), .D(n22), .Q(o_ckv_ia_wdata_part1[16]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[17] ( .CK(clk), .CE(n122), .R(n261), .D(n23), .Q(o_ckv_ia_wdata_part1[17]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[18] ( .CK(clk), .CE(n122), .R(n261), .D(n24), .Q(o_ckv_ia_wdata_part1[18]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[19] ( .CK(clk), .CE(n122), .R(n261), .D(n25), .Q(o_ckv_ia_wdata_part1[19]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[20] ( .CK(clk), .CE(n122), .R(n261), .D(n26), .Q(o_ckv_ia_wdata_part1[20]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[21] ( .CK(clk), .CE(n122), .R(n261), .D(n27), .Q(o_ckv_ia_wdata_part1[21]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[22] ( .CK(clk), .CE(n122), .R(n261), .D(n28), .Q(o_ckv_ia_wdata_part1[22]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[23] ( .CK(clk), .CE(n122), .R(n261), .D(n29), .Q(o_ckv_ia_wdata_part1[23]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[24] ( .CK(clk), .CE(n122), .R(n261), .D(n30), .Q(o_ckv_ia_wdata_part1[24]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[25] ( .CK(clk), .CE(n122), .R(n261), .D(n31), .Q(o_ckv_ia_wdata_part1[25]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[26] ( .CK(clk), .CE(n122), .R(n261), .D(n32), .Q(o_ckv_ia_wdata_part1[26]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[27] ( .CK(clk), .CE(n122), .R(n261), .D(n33), .Q(o_ckv_ia_wdata_part1[27]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[28] ( .CK(clk), .CE(n122), .R(n261), .D(n34), .Q(o_ckv_ia_wdata_part1[28]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[29] ( .CK(clk), .CE(n122), .R(n261), .D(n35), .Q(o_ckv_ia_wdata_part1[29]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[30] ( .CK(clk), .CE(n122), .R(n261), .D(n36), .Q(o_ckv_ia_wdata_part1[30]));
Q_FDP4EP \o_ckv_ia_wdata_part1_REG[31] ( .CK(clk), .CE(n122), .R(n261), .D(n37), .Q(o_ckv_ia_wdata_part1[31]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[0] ( .CK(clk), .CE(n121), .R(n261), .D(n6), .Q(o_ckv_ia_wdata_part0[0]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[1] ( .CK(clk), .CE(n121), .R(n261), .D(n7), .Q(o_ckv_ia_wdata_part0[1]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[2] ( .CK(clk), .CE(n121), .R(n261), .D(n8), .Q(o_ckv_ia_wdata_part0[2]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[3] ( .CK(clk), .CE(n121), .R(n261), .D(n9), .Q(o_ckv_ia_wdata_part0[3]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[4] ( .CK(clk), .CE(n121), .R(n261), .D(n10), .Q(o_ckv_ia_wdata_part0[4]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[5] ( .CK(clk), .CE(n121), .R(n261), .D(n11), .Q(o_ckv_ia_wdata_part0[5]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[6] ( .CK(clk), .CE(n121), .R(n261), .D(n12), .Q(o_ckv_ia_wdata_part0[6]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[7] ( .CK(clk), .CE(n121), .R(n261), .D(n13), .Q(o_ckv_ia_wdata_part0[7]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[8] ( .CK(clk), .CE(n121), .R(n261), .D(n14), .Q(o_ckv_ia_wdata_part0[8]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[9] ( .CK(clk), .CE(n121), .R(n261), .D(n15), .Q(o_ckv_ia_wdata_part0[9]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[10] ( .CK(clk), .CE(n121), .R(n261), .D(n16), .Q(o_ckv_ia_wdata_part0[10]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[11] ( .CK(clk), .CE(n121), .R(n261), .D(n17), .Q(o_ckv_ia_wdata_part0[11]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[12] ( .CK(clk), .CE(n121), .R(n261), .D(n18), .Q(o_ckv_ia_wdata_part0[12]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[13] ( .CK(clk), .CE(n121), .R(n261), .D(n19), .Q(o_ckv_ia_wdata_part0[13]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[14] ( .CK(clk), .CE(n121), .R(n261), .D(n20), .Q(o_ckv_ia_wdata_part0[14]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[15] ( .CK(clk), .CE(n121), .R(n261), .D(n21), .Q(o_ckv_ia_wdata_part0[15]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[16] ( .CK(clk), .CE(n121), .R(n261), .D(n22), .Q(o_ckv_ia_wdata_part0[16]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[17] ( .CK(clk), .CE(n121), .R(n261), .D(n23), .Q(o_ckv_ia_wdata_part0[17]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[18] ( .CK(clk), .CE(n121), .R(n261), .D(n24), .Q(o_ckv_ia_wdata_part0[18]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[19] ( .CK(clk), .CE(n121), .R(n261), .D(n25), .Q(o_ckv_ia_wdata_part0[19]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[20] ( .CK(clk), .CE(n121), .R(n261), .D(n26), .Q(o_ckv_ia_wdata_part0[20]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[21] ( .CK(clk), .CE(n121), .R(n261), .D(n27), .Q(o_ckv_ia_wdata_part0[21]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[22] ( .CK(clk), .CE(n121), .R(n261), .D(n28), .Q(o_ckv_ia_wdata_part0[22]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[23] ( .CK(clk), .CE(n121), .R(n261), .D(n29), .Q(o_ckv_ia_wdata_part0[23]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[24] ( .CK(clk), .CE(n121), .R(n261), .D(n30), .Q(o_ckv_ia_wdata_part0[24]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[25] ( .CK(clk), .CE(n121), .R(n261), .D(n31), .Q(o_ckv_ia_wdata_part0[25]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[26] ( .CK(clk), .CE(n121), .R(n261), .D(n32), .Q(o_ckv_ia_wdata_part0[26]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[27] ( .CK(clk), .CE(n121), .R(n261), .D(n33), .Q(o_ckv_ia_wdata_part0[27]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[28] ( .CK(clk), .CE(n121), .R(n261), .D(n34), .Q(o_ckv_ia_wdata_part0[28]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[29] ( .CK(clk), .CE(n121), .R(n261), .D(n35), .Q(o_ckv_ia_wdata_part0[29]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[30] ( .CK(clk), .CE(n121), .R(n261), .D(n36), .Q(o_ckv_ia_wdata_part0[30]));
Q_FDP4EP \o_ckv_ia_wdata_part0_REG[31] ( .CK(clk), .CE(n121), .R(n261), .D(n37), .Q(o_ckv_ia_wdata_part0[31]));
Q_FDP4EP \o_cddip3_out_im_read_done_REG[0] ( .CK(clk), .CE(n120), .R(n261), .D(n36), .Q(o_cddip3_out_im_read_done[0]));
Q_FDP4EP \o_cddip3_out_im_read_done_REG[1] ( .CK(clk), .CE(n120), .R(n261), .D(n37), .Q(o_cddip3_out_im_read_done[1]));
Q_FDP4EP \o_cddip3_out_im_config_REG[0] ( .CK(clk), .CE(n119), .R(n261), .D(n6), .Q(o_cddip3_out_im_config[0]));
Q_FDP4EP \o_cddip3_out_im_config_REG[1] ( .CK(clk), .CE(n119), .R(n261), .D(n7), .Q(o_cddip3_out_im_config[1]));
Q_FDP4EP \o_cddip3_out_im_config_REG[2] ( .CK(clk), .CE(n119), .R(n261), .D(n8), .Q(o_cddip3_out_im_config[2]));
Q_FDP4EP \o_cddip3_out_im_config_REG[3] ( .CK(clk), .CE(n119), .R(n261), .D(n9), .Q(o_cddip3_out_im_config[3]));
Q_FDP4EP \o_cddip3_out_im_config_REG[4] ( .CK(clk), .CE(n119), .R(n261), .D(n10), .Q(o_cddip3_out_im_config[4]));
Q_FDP4EP \o_cddip3_out_im_config_REG[5] ( .CK(clk), .CE(n119), .R(n261), .D(n11), .Q(o_cddip3_out_im_config[5]));
Q_FDP4EP \o_cddip3_out_im_config_REG[6] ( .CK(clk), .CE(n119), .R(n261), .D(n12), .Q(o_cddip3_out_im_config[6]));
Q_FDP4EP \o_cddip3_out_im_config_REG[7] ( .CK(clk), .CE(n119), .R(n261), .D(n13), .Q(o_cddip3_out_im_config[7]));
Q_FDP4EP \o_cddip3_out_im_config_REG[8] ( .CK(clk), .CE(n119), .R(n261), .D(n14), .Q(o_cddip3_out_im_config[8]));
Q_FDP4EP \o_cddip3_out_ia_config_REG[0] ( .CK(clk), .CE(n118), .R(n261), .D(n6), .Q(o_cddip3_out_ia_config[0]));
Q_FDP4EP \o_cddip3_out_ia_config_REG[1] ( .CK(clk), .CE(n118), .R(n261), .D(n7), .Q(o_cddip3_out_ia_config[1]));
Q_FDP4EP \o_cddip3_out_ia_config_REG[2] ( .CK(clk), .CE(n118), .R(n261), .D(n8), .Q(o_cddip3_out_ia_config[2]));
Q_FDP4EP \o_cddip3_out_ia_config_REG[3] ( .CK(clk), .CE(n118), .R(n261), .D(n9), .Q(o_cddip3_out_ia_config[3]));
Q_FDP4EP \o_cddip3_out_ia_config_REG[4] ( .CK(clk), .CE(n118), .R(n261), .D(n10), .Q(o_cddip3_out_ia_config[4]));
Q_FDP4EP \o_cddip3_out_ia_config_REG[5] ( .CK(clk), .CE(n118), .R(n261), .D(n11), .Q(o_cddip3_out_ia_config[5]));
Q_FDP4EP \o_cddip3_out_ia_config_REG[6] ( .CK(clk), .CE(n118), .R(n261), .D(n12), .Q(o_cddip3_out_ia_config[6]));
Q_FDP4EP \o_cddip3_out_ia_config_REG[7] ( .CK(clk), .CE(n118), .R(n261), .D(n13), .Q(o_cddip3_out_ia_config[7]));
Q_FDP4EP \o_cddip3_out_ia_config_REG[8] ( .CK(clk), .CE(n118), .R(n261), .D(n14), .Q(o_cddip3_out_ia_config[8]));
Q_FDP4EP \o_cddip3_out_ia_config_REG[9] ( .CK(clk), .CE(n118), .R(n261), .D(n34), .Q(o_cddip3_out_ia_config[9]));
Q_FDP4EP \o_cddip3_out_ia_config_REG[10] ( .CK(clk), .CE(n118), .R(n261), .D(n35), .Q(o_cddip3_out_ia_config[10]));
Q_FDP4EP \o_cddip3_out_ia_config_REG[11] ( .CK(clk), .CE(n118), .R(n261), .D(n36), .Q(o_cddip3_out_ia_config[11]));
Q_FDP4EP \o_cddip3_out_ia_config_REG[12] ( .CK(clk), .CE(n118), .R(n261), .D(n37), .Q(o_cddip3_out_ia_config[12]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[0] ( .CK(clk), .CE(n117), .R(n261), .D(n6), .Q(o_cddip3_out_ia_wdata_part2[0]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[1] ( .CK(clk), .CE(n117), .R(n261), .D(n7), .Q(o_cddip3_out_ia_wdata_part2[1]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[2] ( .CK(clk), .CE(n117), .R(n261), .D(n8), .Q(o_cddip3_out_ia_wdata_part2[2]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[3] ( .CK(clk), .CE(n117), .R(n261), .D(n9), .Q(o_cddip3_out_ia_wdata_part2[3]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[4] ( .CK(clk), .CE(n117), .R(n261), .D(n10), .Q(o_cddip3_out_ia_wdata_part2[4]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[5] ( .CK(clk), .CE(n117), .R(n261), .D(n11), .Q(o_cddip3_out_ia_wdata_part2[5]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[6] ( .CK(clk), .CE(n117), .R(n261), .D(n12), .Q(o_cddip3_out_ia_wdata_part2[6]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[7] ( .CK(clk), .CE(n117), .R(n261), .D(n13), .Q(o_cddip3_out_ia_wdata_part2[7]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[8] ( .CK(clk), .CE(n117), .R(n261), .D(n14), .Q(o_cddip3_out_ia_wdata_part2[8]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[9] ( .CK(clk), .CE(n117), .R(n261), .D(n15), .Q(o_cddip3_out_ia_wdata_part2[9]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[10] ( .CK(clk), .CE(n117), .R(n261), .D(n16), .Q(o_cddip3_out_ia_wdata_part2[10]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[11] ( .CK(clk), .CE(n117), .R(n261), .D(n17), .Q(o_cddip3_out_ia_wdata_part2[11]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[12] ( .CK(clk), .CE(n117), .R(n261), .D(n18), .Q(o_cddip3_out_ia_wdata_part2[12]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[13] ( .CK(clk), .CE(n117), .R(n261), .D(n19), .Q(o_cddip3_out_ia_wdata_part2[13]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[14] ( .CK(clk), .CE(n117), .R(n261), .D(n20), .Q(o_cddip3_out_ia_wdata_part2[14]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[15] ( .CK(clk), .CE(n117), .R(n261), .D(n21), .Q(o_cddip3_out_ia_wdata_part2[15]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[16] ( .CK(clk), .CE(n117), .R(n261), .D(n22), .Q(o_cddip3_out_ia_wdata_part2[16]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[17] ( .CK(clk), .CE(n117), .R(n261), .D(n23), .Q(o_cddip3_out_ia_wdata_part2[17]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[18] ( .CK(clk), .CE(n117), .R(n261), .D(n24), .Q(o_cddip3_out_ia_wdata_part2[18]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[19] ( .CK(clk), .CE(n117), .R(n261), .D(n25), .Q(o_cddip3_out_ia_wdata_part2[19]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[20] ( .CK(clk), .CE(n117), .R(n261), .D(n26), .Q(o_cddip3_out_ia_wdata_part2[20]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[21] ( .CK(clk), .CE(n117), .R(n261), .D(n27), .Q(o_cddip3_out_ia_wdata_part2[21]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[22] ( .CK(clk), .CE(n117), .R(n261), .D(n28), .Q(o_cddip3_out_ia_wdata_part2[22]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[23] ( .CK(clk), .CE(n117), .R(n261), .D(n29), .Q(o_cddip3_out_ia_wdata_part2[23]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[24] ( .CK(clk), .CE(n117), .R(n261), .D(n30), .Q(o_cddip3_out_ia_wdata_part2[24]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[25] ( .CK(clk), .CE(n117), .R(n261), .D(n31), .Q(o_cddip3_out_ia_wdata_part2[25]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[26] ( .CK(clk), .CE(n117), .R(n261), .D(n32), .Q(o_cddip3_out_ia_wdata_part2[26]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[27] ( .CK(clk), .CE(n117), .R(n261), .D(n33), .Q(o_cddip3_out_ia_wdata_part2[27]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[28] ( .CK(clk), .CE(n117), .R(n261), .D(n34), .Q(o_cddip3_out_ia_wdata_part2[28]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[29] ( .CK(clk), .CE(n117), .R(n261), .D(n35), .Q(o_cddip3_out_ia_wdata_part2[29]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[30] ( .CK(clk), .CE(n117), .R(n261), .D(n36), .Q(o_cddip3_out_ia_wdata_part2[30]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part2_REG[31] ( .CK(clk), .CE(n117), .R(n261), .D(n37), .Q(o_cddip3_out_ia_wdata_part2[31]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[0] ( .CK(clk), .CE(n116), .R(n261), .D(n6), .Q(o_cddip3_out_ia_wdata_part1[0]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[1] ( .CK(clk), .CE(n116), .R(n261), .D(n7), .Q(o_cddip3_out_ia_wdata_part1[1]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[2] ( .CK(clk), .CE(n116), .R(n261), .D(n8), .Q(o_cddip3_out_ia_wdata_part1[2]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[3] ( .CK(clk), .CE(n116), .R(n261), .D(n9), .Q(o_cddip3_out_ia_wdata_part1[3]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[4] ( .CK(clk), .CE(n116), .R(n261), .D(n10), .Q(o_cddip3_out_ia_wdata_part1[4]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[5] ( .CK(clk), .CE(n116), .R(n261), .D(n11), .Q(o_cddip3_out_ia_wdata_part1[5]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[6] ( .CK(clk), .CE(n116), .R(n261), .D(n12), .Q(o_cddip3_out_ia_wdata_part1[6]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[7] ( .CK(clk), .CE(n116), .R(n261), .D(n13), .Q(o_cddip3_out_ia_wdata_part1[7]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[8] ( .CK(clk), .CE(n116), .R(n261), .D(n14), .Q(o_cddip3_out_ia_wdata_part1[8]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[9] ( .CK(clk), .CE(n116), .R(n261), .D(n15), .Q(o_cddip3_out_ia_wdata_part1[9]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[10] ( .CK(clk), .CE(n116), .R(n261), .D(n16), .Q(o_cddip3_out_ia_wdata_part1[10]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[11] ( .CK(clk), .CE(n116), .R(n261), .D(n17), .Q(o_cddip3_out_ia_wdata_part1[11]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[12] ( .CK(clk), .CE(n116), .R(n261), .D(n18), .Q(o_cddip3_out_ia_wdata_part1[12]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[13] ( .CK(clk), .CE(n116), .R(n261), .D(n19), .Q(o_cddip3_out_ia_wdata_part1[13]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[14] ( .CK(clk), .CE(n116), .R(n261), .D(n20), .Q(o_cddip3_out_ia_wdata_part1[14]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[15] ( .CK(clk), .CE(n116), .R(n261), .D(n21), .Q(o_cddip3_out_ia_wdata_part1[15]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[16] ( .CK(clk), .CE(n116), .R(n261), .D(n22), .Q(o_cddip3_out_ia_wdata_part1[16]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[17] ( .CK(clk), .CE(n116), .R(n261), .D(n23), .Q(o_cddip3_out_ia_wdata_part1[17]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[18] ( .CK(clk), .CE(n116), .R(n261), .D(n24), .Q(o_cddip3_out_ia_wdata_part1[18]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[19] ( .CK(clk), .CE(n116), .R(n261), .D(n25), .Q(o_cddip3_out_ia_wdata_part1[19]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[20] ( .CK(clk), .CE(n116), .R(n261), .D(n26), .Q(o_cddip3_out_ia_wdata_part1[20]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[21] ( .CK(clk), .CE(n116), .R(n261), .D(n27), .Q(o_cddip3_out_ia_wdata_part1[21]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[22] ( .CK(clk), .CE(n116), .R(n261), .D(n28), .Q(o_cddip3_out_ia_wdata_part1[22]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[23] ( .CK(clk), .CE(n116), .R(n261), .D(n29), .Q(o_cddip3_out_ia_wdata_part1[23]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[24] ( .CK(clk), .CE(n116), .R(n261), .D(n30), .Q(o_cddip3_out_ia_wdata_part1[24]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[25] ( .CK(clk), .CE(n116), .R(n261), .D(n31), .Q(o_cddip3_out_ia_wdata_part1[25]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[26] ( .CK(clk), .CE(n116), .R(n261), .D(n32), .Q(o_cddip3_out_ia_wdata_part1[26]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[27] ( .CK(clk), .CE(n116), .R(n261), .D(n33), .Q(o_cddip3_out_ia_wdata_part1[27]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[28] ( .CK(clk), .CE(n116), .R(n261), .D(n34), .Q(o_cddip3_out_ia_wdata_part1[28]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[29] ( .CK(clk), .CE(n116), .R(n261), .D(n35), .Q(o_cddip3_out_ia_wdata_part1[29]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[30] ( .CK(clk), .CE(n116), .R(n261), .D(n36), .Q(o_cddip3_out_ia_wdata_part1[30]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part1_REG[31] ( .CK(clk), .CE(n116), .R(n261), .D(n37), .Q(o_cddip3_out_ia_wdata_part1[31]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[0] ( .CK(clk), .CE(n115), .R(n261), .D(n6), .Q(o_cddip3_out_ia_wdata_part0[0]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[1] ( .CK(clk), .CE(n115), .R(n261), .D(n7), .Q(o_cddip3_out_ia_wdata_part0[1]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[2] ( .CK(clk), .CE(n115), .R(n261), .D(n8), .Q(o_cddip3_out_ia_wdata_part0[2]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[3] ( .CK(clk), .CE(n115), .R(n261), .D(n9), .Q(o_cddip3_out_ia_wdata_part0[3]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[4] ( .CK(clk), .CE(n115), .R(n261), .D(n10), .Q(o_cddip3_out_ia_wdata_part0[4]));
Q_FDP4EP \o_cddip3_out_ia_wdata_part0_REG[5] ( .CK(clk), .CE(n115), .R(n261), .D(n11), .Q(o_cddip3_out_ia_wdata_part0[5]));
Q_FDP4EP \o_cddip2_out_im_read_done_REG[0] ( .CK(clk), .CE(n114), .R(n261), .D(n36), .Q(o_cddip2_out_im_read_done[0]));
Q_FDP4EP \o_cddip2_out_im_read_done_REG[1] ( .CK(clk), .CE(n114), .R(n261), .D(n37), .Q(o_cddip2_out_im_read_done[1]));
Q_FDP4EP \o_cddip2_out_im_config_REG[0] ( .CK(clk), .CE(n113), .R(n261), .D(n6), .Q(o_cddip2_out_im_config[0]));
Q_FDP4EP \o_cddip2_out_im_config_REG[1] ( .CK(clk), .CE(n113), .R(n261), .D(n7), .Q(o_cddip2_out_im_config[1]));
Q_FDP4EP \o_cddip2_out_im_config_REG[2] ( .CK(clk), .CE(n113), .R(n261), .D(n8), .Q(o_cddip2_out_im_config[2]));
Q_FDP4EP \o_cddip2_out_im_config_REG[3] ( .CK(clk), .CE(n113), .R(n261), .D(n9), .Q(o_cddip2_out_im_config[3]));
Q_FDP4EP \o_cddip2_out_im_config_REG[4] ( .CK(clk), .CE(n113), .R(n261), .D(n10), .Q(o_cddip2_out_im_config[4]));
Q_FDP4EP \o_cddip2_out_im_config_REG[5] ( .CK(clk), .CE(n113), .R(n261), .D(n11), .Q(o_cddip2_out_im_config[5]));
Q_FDP4EP \o_cddip2_out_im_config_REG[6] ( .CK(clk), .CE(n113), .R(n261), .D(n12), .Q(o_cddip2_out_im_config[6]));
Q_FDP4EP \o_cddip2_out_im_config_REG[7] ( .CK(clk), .CE(n113), .R(n261), .D(n13), .Q(o_cddip2_out_im_config[7]));
Q_FDP4EP \o_cddip2_out_im_config_REG[8] ( .CK(clk), .CE(n113), .R(n261), .D(n14), .Q(o_cddip2_out_im_config[8]));
Q_FDP4EP \o_cddip2_out_ia_config_REG[0] ( .CK(clk), .CE(n112), .R(n261), .D(n6), .Q(o_cddip2_out_ia_config[0]));
Q_FDP4EP \o_cddip2_out_ia_config_REG[1] ( .CK(clk), .CE(n112), .R(n261), .D(n7), .Q(o_cddip2_out_ia_config[1]));
Q_FDP4EP \o_cddip2_out_ia_config_REG[2] ( .CK(clk), .CE(n112), .R(n261), .D(n8), .Q(o_cddip2_out_ia_config[2]));
Q_FDP4EP \o_cddip2_out_ia_config_REG[3] ( .CK(clk), .CE(n112), .R(n261), .D(n9), .Q(o_cddip2_out_ia_config[3]));
Q_FDP4EP \o_cddip2_out_ia_config_REG[4] ( .CK(clk), .CE(n112), .R(n261), .D(n10), .Q(o_cddip2_out_ia_config[4]));
Q_FDP4EP \o_cddip2_out_ia_config_REG[5] ( .CK(clk), .CE(n112), .R(n261), .D(n11), .Q(o_cddip2_out_ia_config[5]));
Q_FDP4EP \o_cddip2_out_ia_config_REG[6] ( .CK(clk), .CE(n112), .R(n261), .D(n12), .Q(o_cddip2_out_ia_config[6]));
Q_FDP4EP \o_cddip2_out_ia_config_REG[7] ( .CK(clk), .CE(n112), .R(n261), .D(n13), .Q(o_cddip2_out_ia_config[7]));
Q_FDP4EP \o_cddip2_out_ia_config_REG[8] ( .CK(clk), .CE(n112), .R(n261), .D(n14), .Q(o_cddip2_out_ia_config[8]));
Q_FDP4EP \o_cddip2_out_ia_config_REG[9] ( .CK(clk), .CE(n112), .R(n261), .D(n34), .Q(o_cddip2_out_ia_config[9]));
Q_FDP4EP \o_cddip2_out_ia_config_REG[10] ( .CK(clk), .CE(n112), .R(n261), .D(n35), .Q(o_cddip2_out_ia_config[10]));
Q_FDP4EP \o_cddip2_out_ia_config_REG[11] ( .CK(clk), .CE(n112), .R(n261), .D(n36), .Q(o_cddip2_out_ia_config[11]));
Q_FDP4EP \o_cddip2_out_ia_config_REG[12] ( .CK(clk), .CE(n112), .R(n261), .D(n37), .Q(o_cddip2_out_ia_config[12]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[0] ( .CK(clk), .CE(n111), .R(n261), .D(n6), .Q(o_cddip2_out_ia_wdata_part2[0]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[1] ( .CK(clk), .CE(n111), .R(n261), .D(n7), .Q(o_cddip2_out_ia_wdata_part2[1]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[2] ( .CK(clk), .CE(n111), .R(n261), .D(n8), .Q(o_cddip2_out_ia_wdata_part2[2]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[3] ( .CK(clk), .CE(n111), .R(n261), .D(n9), .Q(o_cddip2_out_ia_wdata_part2[3]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[4] ( .CK(clk), .CE(n111), .R(n261), .D(n10), .Q(o_cddip2_out_ia_wdata_part2[4]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[5] ( .CK(clk), .CE(n111), .R(n261), .D(n11), .Q(o_cddip2_out_ia_wdata_part2[5]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[6] ( .CK(clk), .CE(n111), .R(n261), .D(n12), .Q(o_cddip2_out_ia_wdata_part2[6]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[7] ( .CK(clk), .CE(n111), .R(n261), .D(n13), .Q(o_cddip2_out_ia_wdata_part2[7]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[8] ( .CK(clk), .CE(n111), .R(n261), .D(n14), .Q(o_cddip2_out_ia_wdata_part2[8]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[9] ( .CK(clk), .CE(n111), .R(n261), .D(n15), .Q(o_cddip2_out_ia_wdata_part2[9]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[10] ( .CK(clk), .CE(n111), .R(n261), .D(n16), .Q(o_cddip2_out_ia_wdata_part2[10]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[11] ( .CK(clk), .CE(n111), .R(n261), .D(n17), .Q(o_cddip2_out_ia_wdata_part2[11]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[12] ( .CK(clk), .CE(n111), .R(n261), .D(n18), .Q(o_cddip2_out_ia_wdata_part2[12]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[13] ( .CK(clk), .CE(n111), .R(n261), .D(n19), .Q(o_cddip2_out_ia_wdata_part2[13]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[14] ( .CK(clk), .CE(n111), .R(n261), .D(n20), .Q(o_cddip2_out_ia_wdata_part2[14]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[15] ( .CK(clk), .CE(n111), .R(n261), .D(n21), .Q(o_cddip2_out_ia_wdata_part2[15]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[16] ( .CK(clk), .CE(n111), .R(n261), .D(n22), .Q(o_cddip2_out_ia_wdata_part2[16]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[17] ( .CK(clk), .CE(n111), .R(n261), .D(n23), .Q(o_cddip2_out_ia_wdata_part2[17]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[18] ( .CK(clk), .CE(n111), .R(n261), .D(n24), .Q(o_cddip2_out_ia_wdata_part2[18]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[19] ( .CK(clk), .CE(n111), .R(n261), .D(n25), .Q(o_cddip2_out_ia_wdata_part2[19]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[20] ( .CK(clk), .CE(n111), .R(n261), .D(n26), .Q(o_cddip2_out_ia_wdata_part2[20]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[21] ( .CK(clk), .CE(n111), .R(n261), .D(n27), .Q(o_cddip2_out_ia_wdata_part2[21]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[22] ( .CK(clk), .CE(n111), .R(n261), .D(n28), .Q(o_cddip2_out_ia_wdata_part2[22]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[23] ( .CK(clk), .CE(n111), .R(n261), .D(n29), .Q(o_cddip2_out_ia_wdata_part2[23]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[24] ( .CK(clk), .CE(n111), .R(n261), .D(n30), .Q(o_cddip2_out_ia_wdata_part2[24]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[25] ( .CK(clk), .CE(n111), .R(n261), .D(n31), .Q(o_cddip2_out_ia_wdata_part2[25]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[26] ( .CK(clk), .CE(n111), .R(n261), .D(n32), .Q(o_cddip2_out_ia_wdata_part2[26]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[27] ( .CK(clk), .CE(n111), .R(n261), .D(n33), .Q(o_cddip2_out_ia_wdata_part2[27]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[28] ( .CK(clk), .CE(n111), .R(n261), .D(n34), .Q(o_cddip2_out_ia_wdata_part2[28]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[29] ( .CK(clk), .CE(n111), .R(n261), .D(n35), .Q(o_cddip2_out_ia_wdata_part2[29]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[30] ( .CK(clk), .CE(n111), .R(n261), .D(n36), .Q(o_cddip2_out_ia_wdata_part2[30]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part2_REG[31] ( .CK(clk), .CE(n111), .R(n261), .D(n37), .Q(o_cddip2_out_ia_wdata_part2[31]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[0] ( .CK(clk), .CE(n110), .R(n261), .D(n6), .Q(o_cddip2_out_ia_wdata_part1[0]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[1] ( .CK(clk), .CE(n110), .R(n261), .D(n7), .Q(o_cddip2_out_ia_wdata_part1[1]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[2] ( .CK(clk), .CE(n110), .R(n261), .D(n8), .Q(o_cddip2_out_ia_wdata_part1[2]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[3] ( .CK(clk), .CE(n110), .R(n261), .D(n9), .Q(o_cddip2_out_ia_wdata_part1[3]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[4] ( .CK(clk), .CE(n110), .R(n261), .D(n10), .Q(o_cddip2_out_ia_wdata_part1[4]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[5] ( .CK(clk), .CE(n110), .R(n261), .D(n11), .Q(o_cddip2_out_ia_wdata_part1[5]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[6] ( .CK(clk), .CE(n110), .R(n261), .D(n12), .Q(o_cddip2_out_ia_wdata_part1[6]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[7] ( .CK(clk), .CE(n110), .R(n261), .D(n13), .Q(o_cddip2_out_ia_wdata_part1[7]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[8] ( .CK(clk), .CE(n110), .R(n261), .D(n14), .Q(o_cddip2_out_ia_wdata_part1[8]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[9] ( .CK(clk), .CE(n110), .R(n261), .D(n15), .Q(o_cddip2_out_ia_wdata_part1[9]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[10] ( .CK(clk), .CE(n110), .R(n261), .D(n16), .Q(o_cddip2_out_ia_wdata_part1[10]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[11] ( .CK(clk), .CE(n110), .R(n261), .D(n17), .Q(o_cddip2_out_ia_wdata_part1[11]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[12] ( .CK(clk), .CE(n110), .R(n261), .D(n18), .Q(o_cddip2_out_ia_wdata_part1[12]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[13] ( .CK(clk), .CE(n110), .R(n261), .D(n19), .Q(o_cddip2_out_ia_wdata_part1[13]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[14] ( .CK(clk), .CE(n110), .R(n261), .D(n20), .Q(o_cddip2_out_ia_wdata_part1[14]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[15] ( .CK(clk), .CE(n110), .R(n261), .D(n21), .Q(o_cddip2_out_ia_wdata_part1[15]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[16] ( .CK(clk), .CE(n110), .R(n261), .D(n22), .Q(o_cddip2_out_ia_wdata_part1[16]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[17] ( .CK(clk), .CE(n110), .R(n261), .D(n23), .Q(o_cddip2_out_ia_wdata_part1[17]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[18] ( .CK(clk), .CE(n110), .R(n261), .D(n24), .Q(o_cddip2_out_ia_wdata_part1[18]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[19] ( .CK(clk), .CE(n110), .R(n261), .D(n25), .Q(o_cddip2_out_ia_wdata_part1[19]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[20] ( .CK(clk), .CE(n110), .R(n261), .D(n26), .Q(o_cddip2_out_ia_wdata_part1[20]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[21] ( .CK(clk), .CE(n110), .R(n261), .D(n27), .Q(o_cddip2_out_ia_wdata_part1[21]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[22] ( .CK(clk), .CE(n110), .R(n261), .D(n28), .Q(o_cddip2_out_ia_wdata_part1[22]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[23] ( .CK(clk), .CE(n110), .R(n261), .D(n29), .Q(o_cddip2_out_ia_wdata_part1[23]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[24] ( .CK(clk), .CE(n110), .R(n261), .D(n30), .Q(o_cddip2_out_ia_wdata_part1[24]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[25] ( .CK(clk), .CE(n110), .R(n261), .D(n31), .Q(o_cddip2_out_ia_wdata_part1[25]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[26] ( .CK(clk), .CE(n110), .R(n261), .D(n32), .Q(o_cddip2_out_ia_wdata_part1[26]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[27] ( .CK(clk), .CE(n110), .R(n261), .D(n33), .Q(o_cddip2_out_ia_wdata_part1[27]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[28] ( .CK(clk), .CE(n110), .R(n261), .D(n34), .Q(o_cddip2_out_ia_wdata_part1[28]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[29] ( .CK(clk), .CE(n110), .R(n261), .D(n35), .Q(o_cddip2_out_ia_wdata_part1[29]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[30] ( .CK(clk), .CE(n110), .R(n261), .D(n36), .Q(o_cddip2_out_ia_wdata_part1[30]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part1_REG[31] ( .CK(clk), .CE(n110), .R(n261), .D(n37), .Q(o_cddip2_out_ia_wdata_part1[31]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[0] ( .CK(clk), .CE(n109), .R(n261), .D(n6), .Q(o_cddip2_out_ia_wdata_part0[0]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[1] ( .CK(clk), .CE(n109), .R(n261), .D(n7), .Q(o_cddip2_out_ia_wdata_part0[1]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[2] ( .CK(clk), .CE(n109), .R(n261), .D(n8), .Q(o_cddip2_out_ia_wdata_part0[2]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[3] ( .CK(clk), .CE(n109), .R(n261), .D(n9), .Q(o_cddip2_out_ia_wdata_part0[3]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[4] ( .CK(clk), .CE(n109), .R(n261), .D(n10), .Q(o_cddip2_out_ia_wdata_part0[4]));
Q_FDP4EP \o_cddip2_out_ia_wdata_part0_REG[5] ( .CK(clk), .CE(n109), .R(n261), .D(n11), .Q(o_cddip2_out_ia_wdata_part0[5]));
Q_FDP4EP \o_cddip1_out_im_read_done_REG[0] ( .CK(clk), .CE(n108), .R(n261), .D(n36), .Q(o_cddip1_out_im_read_done[0]));
Q_FDP4EP \o_cddip1_out_im_read_done_REG[1] ( .CK(clk), .CE(n108), .R(n261), .D(n37), .Q(o_cddip1_out_im_read_done[1]));
Q_FDP4EP \o_cddip1_out_im_config_REG[0] ( .CK(clk), .CE(n107), .R(n261), .D(n6), .Q(o_cddip1_out_im_config[0]));
Q_FDP4EP \o_cddip1_out_im_config_REG[1] ( .CK(clk), .CE(n107), .R(n261), .D(n7), .Q(o_cddip1_out_im_config[1]));
Q_FDP4EP \o_cddip1_out_im_config_REG[2] ( .CK(clk), .CE(n107), .R(n261), .D(n8), .Q(o_cddip1_out_im_config[2]));
Q_FDP4EP \o_cddip1_out_im_config_REG[3] ( .CK(clk), .CE(n107), .R(n261), .D(n9), .Q(o_cddip1_out_im_config[3]));
Q_FDP4EP \o_cddip1_out_im_config_REG[4] ( .CK(clk), .CE(n107), .R(n261), .D(n10), .Q(o_cddip1_out_im_config[4]));
Q_FDP4EP \o_cddip1_out_im_config_REG[5] ( .CK(clk), .CE(n107), .R(n261), .D(n11), .Q(o_cddip1_out_im_config[5]));
Q_FDP4EP \o_cddip1_out_im_config_REG[6] ( .CK(clk), .CE(n107), .R(n261), .D(n12), .Q(o_cddip1_out_im_config[6]));
Q_FDP4EP \o_cddip1_out_im_config_REG[7] ( .CK(clk), .CE(n107), .R(n261), .D(n13), .Q(o_cddip1_out_im_config[7]));
Q_FDP4EP \o_cddip1_out_im_config_REG[8] ( .CK(clk), .CE(n107), .R(n261), .D(n14), .Q(o_cddip1_out_im_config[8]));
Q_FDP4EP \o_cddip1_out_ia_config_REG[0] ( .CK(clk), .CE(n106), .R(n261), .D(n6), .Q(o_cddip1_out_ia_config[0]));
Q_FDP4EP \o_cddip1_out_ia_config_REG[1] ( .CK(clk), .CE(n106), .R(n261), .D(n7), .Q(o_cddip1_out_ia_config[1]));
Q_FDP4EP \o_cddip1_out_ia_config_REG[2] ( .CK(clk), .CE(n106), .R(n261), .D(n8), .Q(o_cddip1_out_ia_config[2]));
Q_FDP4EP \o_cddip1_out_ia_config_REG[3] ( .CK(clk), .CE(n106), .R(n261), .D(n9), .Q(o_cddip1_out_ia_config[3]));
Q_FDP4EP \o_cddip1_out_ia_config_REG[4] ( .CK(clk), .CE(n106), .R(n261), .D(n10), .Q(o_cddip1_out_ia_config[4]));
Q_FDP4EP \o_cddip1_out_ia_config_REG[5] ( .CK(clk), .CE(n106), .R(n261), .D(n11), .Q(o_cddip1_out_ia_config[5]));
Q_FDP4EP \o_cddip1_out_ia_config_REG[6] ( .CK(clk), .CE(n106), .R(n261), .D(n12), .Q(o_cddip1_out_ia_config[6]));
Q_FDP4EP \o_cddip1_out_ia_config_REG[7] ( .CK(clk), .CE(n106), .R(n261), .D(n13), .Q(o_cddip1_out_ia_config[7]));
Q_FDP4EP \o_cddip1_out_ia_config_REG[8] ( .CK(clk), .CE(n106), .R(n261), .D(n14), .Q(o_cddip1_out_ia_config[8]));
Q_FDP4EP \o_cddip1_out_ia_config_REG[9] ( .CK(clk), .CE(n106), .R(n261), .D(n34), .Q(o_cddip1_out_ia_config[9]));
Q_FDP4EP \o_cddip1_out_ia_config_REG[10] ( .CK(clk), .CE(n106), .R(n261), .D(n35), .Q(o_cddip1_out_ia_config[10]));
Q_FDP4EP \o_cddip1_out_ia_config_REG[11] ( .CK(clk), .CE(n106), .R(n261), .D(n36), .Q(o_cddip1_out_ia_config[11]));
Q_FDP4EP \o_cddip1_out_ia_config_REG[12] ( .CK(clk), .CE(n106), .R(n261), .D(n37), .Q(o_cddip1_out_ia_config[12]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[0] ( .CK(clk), .CE(n105), .R(n261), .D(n6), .Q(o_cddip1_out_ia_wdata_part2[0]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[1] ( .CK(clk), .CE(n105), .R(n261), .D(n7), .Q(o_cddip1_out_ia_wdata_part2[1]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[2] ( .CK(clk), .CE(n105), .R(n261), .D(n8), .Q(o_cddip1_out_ia_wdata_part2[2]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[3] ( .CK(clk), .CE(n105), .R(n261), .D(n9), .Q(o_cddip1_out_ia_wdata_part2[3]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[4] ( .CK(clk), .CE(n105), .R(n261), .D(n10), .Q(o_cddip1_out_ia_wdata_part2[4]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[5] ( .CK(clk), .CE(n105), .R(n261), .D(n11), .Q(o_cddip1_out_ia_wdata_part2[5]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[6] ( .CK(clk), .CE(n105), .R(n261), .D(n12), .Q(o_cddip1_out_ia_wdata_part2[6]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[7] ( .CK(clk), .CE(n105), .R(n261), .D(n13), .Q(o_cddip1_out_ia_wdata_part2[7]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[8] ( .CK(clk), .CE(n105), .R(n261), .D(n14), .Q(o_cddip1_out_ia_wdata_part2[8]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[9] ( .CK(clk), .CE(n105), .R(n261), .D(n15), .Q(o_cddip1_out_ia_wdata_part2[9]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[10] ( .CK(clk), .CE(n105), .R(n261), .D(n16), .Q(o_cddip1_out_ia_wdata_part2[10]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[11] ( .CK(clk), .CE(n105), .R(n261), .D(n17), .Q(o_cddip1_out_ia_wdata_part2[11]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[12] ( .CK(clk), .CE(n105), .R(n261), .D(n18), .Q(o_cddip1_out_ia_wdata_part2[12]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[13] ( .CK(clk), .CE(n105), .R(n261), .D(n19), .Q(o_cddip1_out_ia_wdata_part2[13]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[14] ( .CK(clk), .CE(n105), .R(n261), .D(n20), .Q(o_cddip1_out_ia_wdata_part2[14]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[15] ( .CK(clk), .CE(n105), .R(n261), .D(n21), .Q(o_cddip1_out_ia_wdata_part2[15]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[16] ( .CK(clk), .CE(n105), .R(n261), .D(n22), .Q(o_cddip1_out_ia_wdata_part2[16]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[17] ( .CK(clk), .CE(n105), .R(n261), .D(n23), .Q(o_cddip1_out_ia_wdata_part2[17]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[18] ( .CK(clk), .CE(n105), .R(n261), .D(n24), .Q(o_cddip1_out_ia_wdata_part2[18]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[19] ( .CK(clk), .CE(n105), .R(n261), .D(n25), .Q(o_cddip1_out_ia_wdata_part2[19]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[20] ( .CK(clk), .CE(n105), .R(n261), .D(n26), .Q(o_cddip1_out_ia_wdata_part2[20]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[21] ( .CK(clk), .CE(n105), .R(n261), .D(n27), .Q(o_cddip1_out_ia_wdata_part2[21]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[22] ( .CK(clk), .CE(n105), .R(n261), .D(n28), .Q(o_cddip1_out_ia_wdata_part2[22]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[23] ( .CK(clk), .CE(n105), .R(n261), .D(n29), .Q(o_cddip1_out_ia_wdata_part2[23]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[24] ( .CK(clk), .CE(n105), .R(n261), .D(n30), .Q(o_cddip1_out_ia_wdata_part2[24]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[25] ( .CK(clk), .CE(n105), .R(n261), .D(n31), .Q(o_cddip1_out_ia_wdata_part2[25]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[26] ( .CK(clk), .CE(n105), .R(n261), .D(n32), .Q(o_cddip1_out_ia_wdata_part2[26]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[27] ( .CK(clk), .CE(n105), .R(n261), .D(n33), .Q(o_cddip1_out_ia_wdata_part2[27]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[28] ( .CK(clk), .CE(n105), .R(n261), .D(n34), .Q(o_cddip1_out_ia_wdata_part2[28]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[29] ( .CK(clk), .CE(n105), .R(n261), .D(n35), .Q(o_cddip1_out_ia_wdata_part2[29]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[30] ( .CK(clk), .CE(n105), .R(n261), .D(n36), .Q(o_cddip1_out_ia_wdata_part2[30]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part2_REG[31] ( .CK(clk), .CE(n105), .R(n261), .D(n37), .Q(o_cddip1_out_ia_wdata_part2[31]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[0] ( .CK(clk), .CE(n104), .R(n261), .D(n6), .Q(o_cddip1_out_ia_wdata_part1[0]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[1] ( .CK(clk), .CE(n104), .R(n261), .D(n7), .Q(o_cddip1_out_ia_wdata_part1[1]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[2] ( .CK(clk), .CE(n104), .R(n261), .D(n8), .Q(o_cddip1_out_ia_wdata_part1[2]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[3] ( .CK(clk), .CE(n104), .R(n261), .D(n9), .Q(o_cddip1_out_ia_wdata_part1[3]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[4] ( .CK(clk), .CE(n104), .R(n261), .D(n10), .Q(o_cddip1_out_ia_wdata_part1[4]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[5] ( .CK(clk), .CE(n104), .R(n261), .D(n11), .Q(o_cddip1_out_ia_wdata_part1[5]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[6] ( .CK(clk), .CE(n104), .R(n261), .D(n12), .Q(o_cddip1_out_ia_wdata_part1[6]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[7] ( .CK(clk), .CE(n104), .R(n261), .D(n13), .Q(o_cddip1_out_ia_wdata_part1[7]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[8] ( .CK(clk), .CE(n104), .R(n261), .D(n14), .Q(o_cddip1_out_ia_wdata_part1[8]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[9] ( .CK(clk), .CE(n104), .R(n261), .D(n15), .Q(o_cddip1_out_ia_wdata_part1[9]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[10] ( .CK(clk), .CE(n104), .R(n261), .D(n16), .Q(o_cddip1_out_ia_wdata_part1[10]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[11] ( .CK(clk), .CE(n104), .R(n261), .D(n17), .Q(o_cddip1_out_ia_wdata_part1[11]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[12] ( .CK(clk), .CE(n104), .R(n261), .D(n18), .Q(o_cddip1_out_ia_wdata_part1[12]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[13] ( .CK(clk), .CE(n104), .R(n261), .D(n19), .Q(o_cddip1_out_ia_wdata_part1[13]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[14] ( .CK(clk), .CE(n104), .R(n261), .D(n20), .Q(o_cddip1_out_ia_wdata_part1[14]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[15] ( .CK(clk), .CE(n104), .R(n261), .D(n21), .Q(o_cddip1_out_ia_wdata_part1[15]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[16] ( .CK(clk), .CE(n104), .R(n261), .D(n22), .Q(o_cddip1_out_ia_wdata_part1[16]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[17] ( .CK(clk), .CE(n104), .R(n261), .D(n23), .Q(o_cddip1_out_ia_wdata_part1[17]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[18] ( .CK(clk), .CE(n104), .R(n261), .D(n24), .Q(o_cddip1_out_ia_wdata_part1[18]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[19] ( .CK(clk), .CE(n104), .R(n261), .D(n25), .Q(o_cddip1_out_ia_wdata_part1[19]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[20] ( .CK(clk), .CE(n104), .R(n261), .D(n26), .Q(o_cddip1_out_ia_wdata_part1[20]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[21] ( .CK(clk), .CE(n104), .R(n261), .D(n27), .Q(o_cddip1_out_ia_wdata_part1[21]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[22] ( .CK(clk), .CE(n104), .R(n261), .D(n28), .Q(o_cddip1_out_ia_wdata_part1[22]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[23] ( .CK(clk), .CE(n104), .R(n261), .D(n29), .Q(o_cddip1_out_ia_wdata_part1[23]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[24] ( .CK(clk), .CE(n104), .R(n261), .D(n30), .Q(o_cddip1_out_ia_wdata_part1[24]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[25] ( .CK(clk), .CE(n104), .R(n261), .D(n31), .Q(o_cddip1_out_ia_wdata_part1[25]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[26] ( .CK(clk), .CE(n104), .R(n261), .D(n32), .Q(o_cddip1_out_ia_wdata_part1[26]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[27] ( .CK(clk), .CE(n104), .R(n261), .D(n33), .Q(o_cddip1_out_ia_wdata_part1[27]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[28] ( .CK(clk), .CE(n104), .R(n261), .D(n34), .Q(o_cddip1_out_ia_wdata_part1[28]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[29] ( .CK(clk), .CE(n104), .R(n261), .D(n35), .Q(o_cddip1_out_ia_wdata_part1[29]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[30] ( .CK(clk), .CE(n104), .R(n261), .D(n36), .Q(o_cddip1_out_ia_wdata_part1[30]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part1_REG[31] ( .CK(clk), .CE(n104), .R(n261), .D(n37), .Q(o_cddip1_out_ia_wdata_part1[31]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[0] ( .CK(clk), .CE(n103), .R(n261), .D(n6), .Q(o_cddip1_out_ia_wdata_part0[0]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[1] ( .CK(clk), .CE(n103), .R(n261), .D(n7), .Q(o_cddip1_out_ia_wdata_part0[1]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[2] ( .CK(clk), .CE(n103), .R(n261), .D(n8), .Q(o_cddip1_out_ia_wdata_part0[2]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[3] ( .CK(clk), .CE(n103), .R(n261), .D(n9), .Q(o_cddip1_out_ia_wdata_part0[3]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[4] ( .CK(clk), .CE(n103), .R(n261), .D(n10), .Q(o_cddip1_out_ia_wdata_part0[4]));
Q_FDP4EP \o_cddip1_out_ia_wdata_part0_REG[5] ( .CK(clk), .CE(n103), .R(n261), .D(n11), .Q(o_cddip1_out_ia_wdata_part0[5]));
Q_FDP4EP \o_cddip0_out_im_read_done_REG[0] ( .CK(clk), .CE(n102), .R(n261), .D(n36), .Q(o_cddip0_out_im_read_done[0]));
Q_FDP4EP \o_cddip0_out_im_read_done_REG[1] ( .CK(clk), .CE(n102), .R(n261), .D(n37), .Q(o_cddip0_out_im_read_done[1]));
Q_FDP4EP \o_cddip0_out_im_config_REG[0] ( .CK(clk), .CE(n101), .R(n261), .D(n6), .Q(o_cddip0_out_im_config[0]));
Q_FDP4EP \o_cddip0_out_im_config_REG[1] ( .CK(clk), .CE(n101), .R(n261), .D(n7), .Q(o_cddip0_out_im_config[1]));
Q_FDP4EP \o_cddip0_out_im_config_REG[2] ( .CK(clk), .CE(n101), .R(n261), .D(n8), .Q(o_cddip0_out_im_config[2]));
Q_FDP4EP \o_cddip0_out_im_config_REG[3] ( .CK(clk), .CE(n101), .R(n261), .D(n9), .Q(o_cddip0_out_im_config[3]));
Q_FDP4EP \o_cddip0_out_im_config_REG[4] ( .CK(clk), .CE(n101), .R(n261), .D(n10), .Q(o_cddip0_out_im_config[4]));
Q_FDP4EP \o_cddip0_out_im_config_REG[5] ( .CK(clk), .CE(n101), .R(n261), .D(n11), .Q(o_cddip0_out_im_config[5]));
Q_FDP4EP \o_cddip0_out_im_config_REG[6] ( .CK(clk), .CE(n101), .R(n261), .D(n12), .Q(o_cddip0_out_im_config[6]));
Q_FDP4EP \o_cddip0_out_im_config_REG[7] ( .CK(clk), .CE(n101), .R(n261), .D(n13), .Q(o_cddip0_out_im_config[7]));
Q_FDP4EP \o_cddip0_out_im_config_REG[8] ( .CK(clk), .CE(n101), .R(n261), .D(n14), .Q(o_cddip0_out_im_config[8]));
Q_FDP4EP \o_cddip0_out_ia_config_REG[0] ( .CK(clk), .CE(n100), .R(n261), .D(n6), .Q(o_cddip0_out_ia_config[0]));
Q_FDP4EP \o_cddip0_out_ia_config_REG[1] ( .CK(clk), .CE(n100), .R(n261), .D(n7), .Q(o_cddip0_out_ia_config[1]));
Q_FDP4EP \o_cddip0_out_ia_config_REG[2] ( .CK(clk), .CE(n100), .R(n261), .D(n8), .Q(o_cddip0_out_ia_config[2]));
Q_FDP4EP \o_cddip0_out_ia_config_REG[3] ( .CK(clk), .CE(n100), .R(n261), .D(n9), .Q(o_cddip0_out_ia_config[3]));
Q_FDP4EP \o_cddip0_out_ia_config_REG[4] ( .CK(clk), .CE(n100), .R(n261), .D(n10), .Q(o_cddip0_out_ia_config[4]));
Q_FDP4EP \o_cddip0_out_ia_config_REG[5] ( .CK(clk), .CE(n100), .R(n261), .D(n11), .Q(o_cddip0_out_ia_config[5]));
Q_FDP4EP \o_cddip0_out_ia_config_REG[6] ( .CK(clk), .CE(n100), .R(n261), .D(n12), .Q(o_cddip0_out_ia_config[6]));
Q_FDP4EP \o_cddip0_out_ia_config_REG[7] ( .CK(clk), .CE(n100), .R(n261), .D(n13), .Q(o_cddip0_out_ia_config[7]));
Q_FDP4EP \o_cddip0_out_ia_config_REG[8] ( .CK(clk), .CE(n100), .R(n261), .D(n14), .Q(o_cddip0_out_ia_config[8]));
Q_FDP4EP \o_cddip0_out_ia_config_REG[9] ( .CK(clk), .CE(n100), .R(n261), .D(n34), .Q(o_cddip0_out_ia_config[9]));
Q_FDP4EP \o_cddip0_out_ia_config_REG[10] ( .CK(clk), .CE(n100), .R(n261), .D(n35), .Q(o_cddip0_out_ia_config[10]));
Q_FDP4EP \o_cddip0_out_ia_config_REG[11] ( .CK(clk), .CE(n100), .R(n261), .D(n36), .Q(o_cddip0_out_ia_config[11]));
Q_FDP4EP \o_cddip0_out_ia_config_REG[12] ( .CK(clk), .CE(n100), .R(n261), .D(n37), .Q(o_cddip0_out_ia_config[12]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[0] ( .CK(clk), .CE(n99), .R(n261), .D(n6), .Q(o_cddip0_out_ia_wdata_part2[0]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[1] ( .CK(clk), .CE(n99), .R(n261), .D(n7), .Q(o_cddip0_out_ia_wdata_part2[1]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[2] ( .CK(clk), .CE(n99), .R(n261), .D(n8), .Q(o_cddip0_out_ia_wdata_part2[2]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[3] ( .CK(clk), .CE(n99), .R(n261), .D(n9), .Q(o_cddip0_out_ia_wdata_part2[3]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[4] ( .CK(clk), .CE(n99), .R(n261), .D(n10), .Q(o_cddip0_out_ia_wdata_part2[4]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[5] ( .CK(clk), .CE(n99), .R(n261), .D(n11), .Q(o_cddip0_out_ia_wdata_part2[5]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[6] ( .CK(clk), .CE(n99), .R(n261), .D(n12), .Q(o_cddip0_out_ia_wdata_part2[6]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[7] ( .CK(clk), .CE(n99), .R(n261), .D(n13), .Q(o_cddip0_out_ia_wdata_part2[7]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[8] ( .CK(clk), .CE(n99), .R(n261), .D(n14), .Q(o_cddip0_out_ia_wdata_part2[8]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[9] ( .CK(clk), .CE(n99), .R(n261), .D(n15), .Q(o_cddip0_out_ia_wdata_part2[9]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[10] ( .CK(clk), .CE(n99), .R(n261), .D(n16), .Q(o_cddip0_out_ia_wdata_part2[10]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[11] ( .CK(clk), .CE(n99), .R(n261), .D(n17), .Q(o_cddip0_out_ia_wdata_part2[11]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[12] ( .CK(clk), .CE(n99), .R(n261), .D(n18), .Q(o_cddip0_out_ia_wdata_part2[12]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[13] ( .CK(clk), .CE(n99), .R(n261), .D(n19), .Q(o_cddip0_out_ia_wdata_part2[13]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[14] ( .CK(clk), .CE(n99), .R(n261), .D(n20), .Q(o_cddip0_out_ia_wdata_part2[14]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[15] ( .CK(clk), .CE(n99), .R(n261), .D(n21), .Q(o_cddip0_out_ia_wdata_part2[15]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[16] ( .CK(clk), .CE(n99), .R(n261), .D(n22), .Q(o_cddip0_out_ia_wdata_part2[16]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[17] ( .CK(clk), .CE(n99), .R(n261), .D(n23), .Q(o_cddip0_out_ia_wdata_part2[17]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[18] ( .CK(clk), .CE(n99), .R(n261), .D(n24), .Q(o_cddip0_out_ia_wdata_part2[18]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[19] ( .CK(clk), .CE(n99), .R(n261), .D(n25), .Q(o_cddip0_out_ia_wdata_part2[19]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[20] ( .CK(clk), .CE(n99), .R(n261), .D(n26), .Q(o_cddip0_out_ia_wdata_part2[20]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[21] ( .CK(clk), .CE(n99), .R(n261), .D(n27), .Q(o_cddip0_out_ia_wdata_part2[21]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[22] ( .CK(clk), .CE(n99), .R(n261), .D(n28), .Q(o_cddip0_out_ia_wdata_part2[22]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[23] ( .CK(clk), .CE(n99), .R(n261), .D(n29), .Q(o_cddip0_out_ia_wdata_part2[23]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[24] ( .CK(clk), .CE(n99), .R(n261), .D(n30), .Q(o_cddip0_out_ia_wdata_part2[24]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[25] ( .CK(clk), .CE(n99), .R(n261), .D(n31), .Q(o_cddip0_out_ia_wdata_part2[25]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[26] ( .CK(clk), .CE(n99), .R(n261), .D(n32), .Q(o_cddip0_out_ia_wdata_part2[26]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[27] ( .CK(clk), .CE(n99), .R(n261), .D(n33), .Q(o_cddip0_out_ia_wdata_part2[27]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[28] ( .CK(clk), .CE(n99), .R(n261), .D(n34), .Q(o_cddip0_out_ia_wdata_part2[28]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[29] ( .CK(clk), .CE(n99), .R(n261), .D(n35), .Q(o_cddip0_out_ia_wdata_part2[29]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[30] ( .CK(clk), .CE(n99), .R(n261), .D(n36), .Q(o_cddip0_out_ia_wdata_part2[30]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part2_REG[31] ( .CK(clk), .CE(n99), .R(n261), .D(n37), .Q(o_cddip0_out_ia_wdata_part2[31]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[0] ( .CK(clk), .CE(n98), .R(n261), .D(n6), .Q(o_cddip0_out_ia_wdata_part1[0]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[1] ( .CK(clk), .CE(n98), .R(n261), .D(n7), .Q(o_cddip0_out_ia_wdata_part1[1]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[2] ( .CK(clk), .CE(n98), .R(n261), .D(n8), .Q(o_cddip0_out_ia_wdata_part1[2]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[3] ( .CK(clk), .CE(n98), .R(n261), .D(n9), .Q(o_cddip0_out_ia_wdata_part1[3]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[4] ( .CK(clk), .CE(n98), .R(n261), .D(n10), .Q(o_cddip0_out_ia_wdata_part1[4]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[5] ( .CK(clk), .CE(n98), .R(n261), .D(n11), .Q(o_cddip0_out_ia_wdata_part1[5]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[6] ( .CK(clk), .CE(n98), .R(n261), .D(n12), .Q(o_cddip0_out_ia_wdata_part1[6]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[7] ( .CK(clk), .CE(n98), .R(n261), .D(n13), .Q(o_cddip0_out_ia_wdata_part1[7]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[8] ( .CK(clk), .CE(n98), .R(n261), .D(n14), .Q(o_cddip0_out_ia_wdata_part1[8]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[9] ( .CK(clk), .CE(n98), .R(n261), .D(n15), .Q(o_cddip0_out_ia_wdata_part1[9]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[10] ( .CK(clk), .CE(n98), .R(n261), .D(n16), .Q(o_cddip0_out_ia_wdata_part1[10]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[11] ( .CK(clk), .CE(n98), .R(n261), .D(n17), .Q(o_cddip0_out_ia_wdata_part1[11]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[12] ( .CK(clk), .CE(n98), .R(n261), .D(n18), .Q(o_cddip0_out_ia_wdata_part1[12]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[13] ( .CK(clk), .CE(n98), .R(n261), .D(n19), .Q(o_cddip0_out_ia_wdata_part1[13]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[14] ( .CK(clk), .CE(n98), .R(n261), .D(n20), .Q(o_cddip0_out_ia_wdata_part1[14]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[15] ( .CK(clk), .CE(n98), .R(n261), .D(n21), .Q(o_cddip0_out_ia_wdata_part1[15]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[16] ( .CK(clk), .CE(n98), .R(n261), .D(n22), .Q(o_cddip0_out_ia_wdata_part1[16]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[17] ( .CK(clk), .CE(n98), .R(n261), .D(n23), .Q(o_cddip0_out_ia_wdata_part1[17]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[18] ( .CK(clk), .CE(n98), .R(n261), .D(n24), .Q(o_cddip0_out_ia_wdata_part1[18]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[19] ( .CK(clk), .CE(n98), .R(n261), .D(n25), .Q(o_cddip0_out_ia_wdata_part1[19]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[20] ( .CK(clk), .CE(n98), .R(n261), .D(n26), .Q(o_cddip0_out_ia_wdata_part1[20]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[21] ( .CK(clk), .CE(n98), .R(n261), .D(n27), .Q(o_cddip0_out_ia_wdata_part1[21]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[22] ( .CK(clk), .CE(n98), .R(n261), .D(n28), .Q(o_cddip0_out_ia_wdata_part1[22]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[23] ( .CK(clk), .CE(n98), .R(n261), .D(n29), .Q(o_cddip0_out_ia_wdata_part1[23]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[24] ( .CK(clk), .CE(n98), .R(n261), .D(n30), .Q(o_cddip0_out_ia_wdata_part1[24]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[25] ( .CK(clk), .CE(n98), .R(n261), .D(n31), .Q(o_cddip0_out_ia_wdata_part1[25]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[26] ( .CK(clk), .CE(n98), .R(n261), .D(n32), .Q(o_cddip0_out_ia_wdata_part1[26]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[27] ( .CK(clk), .CE(n98), .R(n261), .D(n33), .Q(o_cddip0_out_ia_wdata_part1[27]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[28] ( .CK(clk), .CE(n98), .R(n261), .D(n34), .Q(o_cddip0_out_ia_wdata_part1[28]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[29] ( .CK(clk), .CE(n98), .R(n261), .D(n35), .Q(o_cddip0_out_ia_wdata_part1[29]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[30] ( .CK(clk), .CE(n98), .R(n261), .D(n36), .Q(o_cddip0_out_ia_wdata_part1[30]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part1_REG[31] ( .CK(clk), .CE(n98), .R(n261), .D(n37), .Q(o_cddip0_out_ia_wdata_part1[31]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[0] ( .CK(clk), .CE(n97), .R(n261), .D(n6), .Q(o_cddip0_out_ia_wdata_part0[0]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[1] ( .CK(clk), .CE(n97), .R(n261), .D(n7), .Q(o_cddip0_out_ia_wdata_part0[1]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[2] ( .CK(clk), .CE(n97), .R(n261), .D(n8), .Q(o_cddip0_out_ia_wdata_part0[2]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[3] ( .CK(clk), .CE(n97), .R(n261), .D(n9), .Q(o_cddip0_out_ia_wdata_part0[3]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[4] ( .CK(clk), .CE(n97), .R(n261), .D(n10), .Q(o_cddip0_out_ia_wdata_part0[4]));
Q_FDP4EP \o_cddip0_out_ia_wdata_part0_REG[5] ( .CK(clk), .CE(n97), .R(n261), .D(n11), .Q(o_cddip0_out_ia_wdata_part0[5]));
Q_FDP4EP \o_cceip3_out_im_read_done_REG[0] ( .CK(clk), .CE(n96), .R(n261), .D(n36), .Q(o_cceip3_out_im_read_done[0]));
Q_FDP4EP \o_cceip3_out_im_read_done_REG[1] ( .CK(clk), .CE(n96), .R(n261), .D(n37), .Q(o_cceip3_out_im_read_done[1]));
Q_FDP4EP \o_cceip3_out_im_config_REG[0] ( .CK(clk), .CE(n95), .R(n261), .D(n6), .Q(o_cceip3_out_im_config[0]));
Q_FDP4EP \o_cceip3_out_im_config_REG[1] ( .CK(clk), .CE(n95), .R(n261), .D(n7), .Q(o_cceip3_out_im_config[1]));
Q_FDP4EP \o_cceip3_out_im_config_REG[2] ( .CK(clk), .CE(n95), .R(n261), .D(n8), .Q(o_cceip3_out_im_config[2]));
Q_FDP4EP \o_cceip3_out_im_config_REG[3] ( .CK(clk), .CE(n95), .R(n261), .D(n9), .Q(o_cceip3_out_im_config[3]));
Q_FDP4EP \o_cceip3_out_im_config_REG[4] ( .CK(clk), .CE(n95), .R(n261), .D(n10), .Q(o_cceip3_out_im_config[4]));
Q_FDP4EP \o_cceip3_out_im_config_REG[5] ( .CK(clk), .CE(n95), .R(n261), .D(n11), .Q(o_cceip3_out_im_config[5]));
Q_FDP4EP \o_cceip3_out_im_config_REG[6] ( .CK(clk), .CE(n95), .R(n261), .D(n12), .Q(o_cceip3_out_im_config[6]));
Q_FDP4EP \o_cceip3_out_im_config_REG[7] ( .CK(clk), .CE(n95), .R(n261), .D(n13), .Q(o_cceip3_out_im_config[7]));
Q_FDP4EP \o_cceip3_out_im_config_REG[8] ( .CK(clk), .CE(n95), .R(n261), .D(n14), .Q(o_cceip3_out_im_config[8]));
Q_FDP4EP \o_cceip3_out_ia_config_REG[0] ( .CK(clk), .CE(n94), .R(n261), .D(n6), .Q(o_cceip3_out_ia_config[0]));
Q_FDP4EP \o_cceip3_out_ia_config_REG[1] ( .CK(clk), .CE(n94), .R(n261), .D(n7), .Q(o_cceip3_out_ia_config[1]));
Q_FDP4EP \o_cceip3_out_ia_config_REG[2] ( .CK(clk), .CE(n94), .R(n261), .D(n8), .Q(o_cceip3_out_ia_config[2]));
Q_FDP4EP \o_cceip3_out_ia_config_REG[3] ( .CK(clk), .CE(n94), .R(n261), .D(n9), .Q(o_cceip3_out_ia_config[3]));
Q_FDP4EP \o_cceip3_out_ia_config_REG[4] ( .CK(clk), .CE(n94), .R(n261), .D(n10), .Q(o_cceip3_out_ia_config[4]));
Q_FDP4EP \o_cceip3_out_ia_config_REG[5] ( .CK(clk), .CE(n94), .R(n261), .D(n11), .Q(o_cceip3_out_ia_config[5]));
Q_FDP4EP \o_cceip3_out_ia_config_REG[6] ( .CK(clk), .CE(n94), .R(n261), .D(n12), .Q(o_cceip3_out_ia_config[6]));
Q_FDP4EP \o_cceip3_out_ia_config_REG[7] ( .CK(clk), .CE(n94), .R(n261), .D(n13), .Q(o_cceip3_out_ia_config[7]));
Q_FDP4EP \o_cceip3_out_ia_config_REG[8] ( .CK(clk), .CE(n94), .R(n261), .D(n14), .Q(o_cceip3_out_ia_config[8]));
Q_FDP4EP \o_cceip3_out_ia_config_REG[9] ( .CK(clk), .CE(n94), .R(n261), .D(n34), .Q(o_cceip3_out_ia_config[9]));
Q_FDP4EP \o_cceip3_out_ia_config_REG[10] ( .CK(clk), .CE(n94), .R(n261), .D(n35), .Q(o_cceip3_out_ia_config[10]));
Q_FDP4EP \o_cceip3_out_ia_config_REG[11] ( .CK(clk), .CE(n94), .R(n261), .D(n36), .Q(o_cceip3_out_ia_config[11]));
Q_FDP4EP \o_cceip3_out_ia_config_REG[12] ( .CK(clk), .CE(n94), .R(n261), .D(n37), .Q(o_cceip3_out_ia_config[12]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[0] ( .CK(clk), .CE(n93), .R(n261), .D(n6), .Q(o_cceip3_out_ia_wdata_part2[0]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[1] ( .CK(clk), .CE(n93), .R(n261), .D(n7), .Q(o_cceip3_out_ia_wdata_part2[1]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[2] ( .CK(clk), .CE(n93), .R(n261), .D(n8), .Q(o_cceip3_out_ia_wdata_part2[2]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[3] ( .CK(clk), .CE(n93), .R(n261), .D(n9), .Q(o_cceip3_out_ia_wdata_part2[3]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[4] ( .CK(clk), .CE(n93), .R(n261), .D(n10), .Q(o_cceip3_out_ia_wdata_part2[4]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[5] ( .CK(clk), .CE(n93), .R(n261), .D(n11), .Q(o_cceip3_out_ia_wdata_part2[5]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[6] ( .CK(clk), .CE(n93), .R(n261), .D(n12), .Q(o_cceip3_out_ia_wdata_part2[6]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[7] ( .CK(clk), .CE(n93), .R(n261), .D(n13), .Q(o_cceip3_out_ia_wdata_part2[7]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[8] ( .CK(clk), .CE(n93), .R(n261), .D(n14), .Q(o_cceip3_out_ia_wdata_part2[8]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[9] ( .CK(clk), .CE(n93), .R(n261), .D(n15), .Q(o_cceip3_out_ia_wdata_part2[9]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[10] ( .CK(clk), .CE(n93), .R(n261), .D(n16), .Q(o_cceip3_out_ia_wdata_part2[10]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[11] ( .CK(clk), .CE(n93), .R(n261), .D(n17), .Q(o_cceip3_out_ia_wdata_part2[11]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[12] ( .CK(clk), .CE(n93), .R(n261), .D(n18), .Q(o_cceip3_out_ia_wdata_part2[12]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[13] ( .CK(clk), .CE(n93), .R(n261), .D(n19), .Q(o_cceip3_out_ia_wdata_part2[13]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[14] ( .CK(clk), .CE(n93), .R(n261), .D(n20), .Q(o_cceip3_out_ia_wdata_part2[14]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[15] ( .CK(clk), .CE(n93), .R(n261), .D(n21), .Q(o_cceip3_out_ia_wdata_part2[15]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[16] ( .CK(clk), .CE(n93), .R(n261), .D(n22), .Q(o_cceip3_out_ia_wdata_part2[16]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[17] ( .CK(clk), .CE(n93), .R(n261), .D(n23), .Q(o_cceip3_out_ia_wdata_part2[17]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[18] ( .CK(clk), .CE(n93), .R(n261), .D(n24), .Q(o_cceip3_out_ia_wdata_part2[18]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[19] ( .CK(clk), .CE(n93), .R(n261), .D(n25), .Q(o_cceip3_out_ia_wdata_part2[19]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[20] ( .CK(clk), .CE(n93), .R(n261), .D(n26), .Q(o_cceip3_out_ia_wdata_part2[20]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[21] ( .CK(clk), .CE(n93), .R(n261), .D(n27), .Q(o_cceip3_out_ia_wdata_part2[21]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[22] ( .CK(clk), .CE(n93), .R(n261), .D(n28), .Q(o_cceip3_out_ia_wdata_part2[22]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[23] ( .CK(clk), .CE(n93), .R(n261), .D(n29), .Q(o_cceip3_out_ia_wdata_part2[23]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[24] ( .CK(clk), .CE(n93), .R(n261), .D(n30), .Q(o_cceip3_out_ia_wdata_part2[24]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[25] ( .CK(clk), .CE(n93), .R(n261), .D(n31), .Q(o_cceip3_out_ia_wdata_part2[25]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[26] ( .CK(clk), .CE(n93), .R(n261), .D(n32), .Q(o_cceip3_out_ia_wdata_part2[26]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[27] ( .CK(clk), .CE(n93), .R(n261), .D(n33), .Q(o_cceip3_out_ia_wdata_part2[27]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[28] ( .CK(clk), .CE(n93), .R(n261), .D(n34), .Q(o_cceip3_out_ia_wdata_part2[28]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[29] ( .CK(clk), .CE(n93), .R(n261), .D(n35), .Q(o_cceip3_out_ia_wdata_part2[29]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[30] ( .CK(clk), .CE(n93), .R(n261), .D(n36), .Q(o_cceip3_out_ia_wdata_part2[30]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part2_REG[31] ( .CK(clk), .CE(n93), .R(n261), .D(n37), .Q(o_cceip3_out_ia_wdata_part2[31]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[0] ( .CK(clk), .CE(n92), .R(n261), .D(n6), .Q(o_cceip3_out_ia_wdata_part1[0]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[1] ( .CK(clk), .CE(n92), .R(n261), .D(n7), .Q(o_cceip3_out_ia_wdata_part1[1]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[2] ( .CK(clk), .CE(n92), .R(n261), .D(n8), .Q(o_cceip3_out_ia_wdata_part1[2]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[3] ( .CK(clk), .CE(n92), .R(n261), .D(n9), .Q(o_cceip3_out_ia_wdata_part1[3]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[4] ( .CK(clk), .CE(n92), .R(n261), .D(n10), .Q(o_cceip3_out_ia_wdata_part1[4]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[5] ( .CK(clk), .CE(n92), .R(n261), .D(n11), .Q(o_cceip3_out_ia_wdata_part1[5]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[6] ( .CK(clk), .CE(n92), .R(n261), .D(n12), .Q(o_cceip3_out_ia_wdata_part1[6]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[7] ( .CK(clk), .CE(n92), .R(n261), .D(n13), .Q(o_cceip3_out_ia_wdata_part1[7]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[8] ( .CK(clk), .CE(n92), .R(n261), .D(n14), .Q(o_cceip3_out_ia_wdata_part1[8]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[9] ( .CK(clk), .CE(n92), .R(n261), .D(n15), .Q(o_cceip3_out_ia_wdata_part1[9]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[10] ( .CK(clk), .CE(n92), .R(n261), .D(n16), .Q(o_cceip3_out_ia_wdata_part1[10]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[11] ( .CK(clk), .CE(n92), .R(n261), .D(n17), .Q(o_cceip3_out_ia_wdata_part1[11]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[12] ( .CK(clk), .CE(n92), .R(n261), .D(n18), .Q(o_cceip3_out_ia_wdata_part1[12]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[13] ( .CK(clk), .CE(n92), .R(n261), .D(n19), .Q(o_cceip3_out_ia_wdata_part1[13]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[14] ( .CK(clk), .CE(n92), .R(n261), .D(n20), .Q(o_cceip3_out_ia_wdata_part1[14]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[15] ( .CK(clk), .CE(n92), .R(n261), .D(n21), .Q(o_cceip3_out_ia_wdata_part1[15]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[16] ( .CK(clk), .CE(n92), .R(n261), .D(n22), .Q(o_cceip3_out_ia_wdata_part1[16]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[17] ( .CK(clk), .CE(n92), .R(n261), .D(n23), .Q(o_cceip3_out_ia_wdata_part1[17]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[18] ( .CK(clk), .CE(n92), .R(n261), .D(n24), .Q(o_cceip3_out_ia_wdata_part1[18]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[19] ( .CK(clk), .CE(n92), .R(n261), .D(n25), .Q(o_cceip3_out_ia_wdata_part1[19]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[20] ( .CK(clk), .CE(n92), .R(n261), .D(n26), .Q(o_cceip3_out_ia_wdata_part1[20]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[21] ( .CK(clk), .CE(n92), .R(n261), .D(n27), .Q(o_cceip3_out_ia_wdata_part1[21]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[22] ( .CK(clk), .CE(n92), .R(n261), .D(n28), .Q(o_cceip3_out_ia_wdata_part1[22]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[23] ( .CK(clk), .CE(n92), .R(n261), .D(n29), .Q(o_cceip3_out_ia_wdata_part1[23]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[24] ( .CK(clk), .CE(n92), .R(n261), .D(n30), .Q(o_cceip3_out_ia_wdata_part1[24]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[25] ( .CK(clk), .CE(n92), .R(n261), .D(n31), .Q(o_cceip3_out_ia_wdata_part1[25]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[26] ( .CK(clk), .CE(n92), .R(n261), .D(n32), .Q(o_cceip3_out_ia_wdata_part1[26]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[27] ( .CK(clk), .CE(n92), .R(n261), .D(n33), .Q(o_cceip3_out_ia_wdata_part1[27]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[28] ( .CK(clk), .CE(n92), .R(n261), .D(n34), .Q(o_cceip3_out_ia_wdata_part1[28]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[29] ( .CK(clk), .CE(n92), .R(n261), .D(n35), .Q(o_cceip3_out_ia_wdata_part1[29]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[30] ( .CK(clk), .CE(n92), .R(n261), .D(n36), .Q(o_cceip3_out_ia_wdata_part1[30]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part1_REG[31] ( .CK(clk), .CE(n92), .R(n261), .D(n37), .Q(o_cceip3_out_ia_wdata_part1[31]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[0] ( .CK(clk), .CE(n91), .R(n261), .D(n6), .Q(o_cceip3_out_ia_wdata_part0[0]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[1] ( .CK(clk), .CE(n91), .R(n261), .D(n7), .Q(o_cceip3_out_ia_wdata_part0[1]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[2] ( .CK(clk), .CE(n91), .R(n261), .D(n8), .Q(o_cceip3_out_ia_wdata_part0[2]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[3] ( .CK(clk), .CE(n91), .R(n261), .D(n9), .Q(o_cceip3_out_ia_wdata_part0[3]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[4] ( .CK(clk), .CE(n91), .R(n261), .D(n10), .Q(o_cceip3_out_ia_wdata_part0[4]));
Q_FDP4EP \o_cceip3_out_ia_wdata_part0_REG[5] ( .CK(clk), .CE(n91), .R(n261), .D(n11), .Q(o_cceip3_out_ia_wdata_part0[5]));
Q_FDP4EP \o_cceip2_out_im_read_done_REG[0] ( .CK(clk), .CE(n90), .R(n261), .D(n36), .Q(o_cceip2_out_im_read_done[0]));
Q_FDP4EP \o_cceip2_out_im_read_done_REG[1] ( .CK(clk), .CE(n90), .R(n261), .D(n37), .Q(o_cceip2_out_im_read_done[1]));
Q_FDP4EP \o_cceip2_out_im_config_REG[0] ( .CK(clk), .CE(n89), .R(n261), .D(n6), .Q(o_cceip2_out_im_config[0]));
Q_FDP4EP \o_cceip2_out_im_config_REG[1] ( .CK(clk), .CE(n89), .R(n261), .D(n7), .Q(o_cceip2_out_im_config[1]));
Q_FDP4EP \o_cceip2_out_im_config_REG[2] ( .CK(clk), .CE(n89), .R(n261), .D(n8), .Q(o_cceip2_out_im_config[2]));
Q_FDP4EP \o_cceip2_out_im_config_REG[3] ( .CK(clk), .CE(n89), .R(n261), .D(n9), .Q(o_cceip2_out_im_config[3]));
Q_FDP4EP \o_cceip2_out_im_config_REG[4] ( .CK(clk), .CE(n89), .R(n261), .D(n10), .Q(o_cceip2_out_im_config[4]));
Q_FDP4EP \o_cceip2_out_im_config_REG[5] ( .CK(clk), .CE(n89), .R(n261), .D(n11), .Q(o_cceip2_out_im_config[5]));
Q_FDP4EP \o_cceip2_out_im_config_REG[6] ( .CK(clk), .CE(n89), .R(n261), .D(n12), .Q(o_cceip2_out_im_config[6]));
Q_FDP4EP \o_cceip2_out_im_config_REG[7] ( .CK(clk), .CE(n89), .R(n261), .D(n13), .Q(o_cceip2_out_im_config[7]));
Q_FDP4EP \o_cceip2_out_im_config_REG[8] ( .CK(clk), .CE(n89), .R(n261), .D(n14), .Q(o_cceip2_out_im_config[8]));
Q_FDP4EP \o_cceip2_out_ia_config_REG[0] ( .CK(clk), .CE(n88), .R(n261), .D(n6), .Q(o_cceip2_out_ia_config[0]));
Q_FDP4EP \o_cceip2_out_ia_config_REG[1] ( .CK(clk), .CE(n88), .R(n261), .D(n7), .Q(o_cceip2_out_ia_config[1]));
Q_FDP4EP \o_cceip2_out_ia_config_REG[2] ( .CK(clk), .CE(n88), .R(n261), .D(n8), .Q(o_cceip2_out_ia_config[2]));
Q_FDP4EP \o_cceip2_out_ia_config_REG[3] ( .CK(clk), .CE(n88), .R(n261), .D(n9), .Q(o_cceip2_out_ia_config[3]));
Q_FDP4EP \o_cceip2_out_ia_config_REG[4] ( .CK(clk), .CE(n88), .R(n261), .D(n10), .Q(o_cceip2_out_ia_config[4]));
Q_FDP4EP \o_cceip2_out_ia_config_REG[5] ( .CK(clk), .CE(n88), .R(n261), .D(n11), .Q(o_cceip2_out_ia_config[5]));
Q_FDP4EP \o_cceip2_out_ia_config_REG[6] ( .CK(clk), .CE(n88), .R(n261), .D(n12), .Q(o_cceip2_out_ia_config[6]));
Q_FDP4EP \o_cceip2_out_ia_config_REG[7] ( .CK(clk), .CE(n88), .R(n261), .D(n13), .Q(o_cceip2_out_ia_config[7]));
Q_FDP4EP \o_cceip2_out_ia_config_REG[8] ( .CK(clk), .CE(n88), .R(n261), .D(n14), .Q(o_cceip2_out_ia_config[8]));
Q_FDP4EP \o_cceip2_out_ia_config_REG[9] ( .CK(clk), .CE(n88), .R(n261), .D(n34), .Q(o_cceip2_out_ia_config[9]));
Q_FDP4EP \o_cceip2_out_ia_config_REG[10] ( .CK(clk), .CE(n88), .R(n261), .D(n35), .Q(o_cceip2_out_ia_config[10]));
Q_FDP4EP \o_cceip2_out_ia_config_REG[11] ( .CK(clk), .CE(n88), .R(n261), .D(n36), .Q(o_cceip2_out_ia_config[11]));
Q_FDP4EP \o_cceip2_out_ia_config_REG[12] ( .CK(clk), .CE(n88), .R(n261), .D(n37), .Q(o_cceip2_out_ia_config[12]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[0] ( .CK(clk), .CE(n87), .R(n261), .D(n6), .Q(o_cceip2_out_ia_wdata_part2[0]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[1] ( .CK(clk), .CE(n87), .R(n261), .D(n7), .Q(o_cceip2_out_ia_wdata_part2[1]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[2] ( .CK(clk), .CE(n87), .R(n261), .D(n8), .Q(o_cceip2_out_ia_wdata_part2[2]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[3] ( .CK(clk), .CE(n87), .R(n261), .D(n9), .Q(o_cceip2_out_ia_wdata_part2[3]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[4] ( .CK(clk), .CE(n87), .R(n261), .D(n10), .Q(o_cceip2_out_ia_wdata_part2[4]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[5] ( .CK(clk), .CE(n87), .R(n261), .D(n11), .Q(o_cceip2_out_ia_wdata_part2[5]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[6] ( .CK(clk), .CE(n87), .R(n261), .D(n12), .Q(o_cceip2_out_ia_wdata_part2[6]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[7] ( .CK(clk), .CE(n87), .R(n261), .D(n13), .Q(o_cceip2_out_ia_wdata_part2[7]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[8] ( .CK(clk), .CE(n87), .R(n261), .D(n14), .Q(o_cceip2_out_ia_wdata_part2[8]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[9] ( .CK(clk), .CE(n87), .R(n261), .D(n15), .Q(o_cceip2_out_ia_wdata_part2[9]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[10] ( .CK(clk), .CE(n87), .R(n261), .D(n16), .Q(o_cceip2_out_ia_wdata_part2[10]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[11] ( .CK(clk), .CE(n87), .R(n261), .D(n17), .Q(o_cceip2_out_ia_wdata_part2[11]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[12] ( .CK(clk), .CE(n87), .R(n261), .D(n18), .Q(o_cceip2_out_ia_wdata_part2[12]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[13] ( .CK(clk), .CE(n87), .R(n261), .D(n19), .Q(o_cceip2_out_ia_wdata_part2[13]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[14] ( .CK(clk), .CE(n87), .R(n261), .D(n20), .Q(o_cceip2_out_ia_wdata_part2[14]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[15] ( .CK(clk), .CE(n87), .R(n261), .D(n21), .Q(o_cceip2_out_ia_wdata_part2[15]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[16] ( .CK(clk), .CE(n87), .R(n261), .D(n22), .Q(o_cceip2_out_ia_wdata_part2[16]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[17] ( .CK(clk), .CE(n87), .R(n261), .D(n23), .Q(o_cceip2_out_ia_wdata_part2[17]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[18] ( .CK(clk), .CE(n87), .R(n261), .D(n24), .Q(o_cceip2_out_ia_wdata_part2[18]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[19] ( .CK(clk), .CE(n87), .R(n261), .D(n25), .Q(o_cceip2_out_ia_wdata_part2[19]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[20] ( .CK(clk), .CE(n87), .R(n261), .D(n26), .Q(o_cceip2_out_ia_wdata_part2[20]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[21] ( .CK(clk), .CE(n87), .R(n261), .D(n27), .Q(o_cceip2_out_ia_wdata_part2[21]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[22] ( .CK(clk), .CE(n87), .R(n261), .D(n28), .Q(o_cceip2_out_ia_wdata_part2[22]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[23] ( .CK(clk), .CE(n87), .R(n261), .D(n29), .Q(o_cceip2_out_ia_wdata_part2[23]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[24] ( .CK(clk), .CE(n87), .R(n261), .D(n30), .Q(o_cceip2_out_ia_wdata_part2[24]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[25] ( .CK(clk), .CE(n87), .R(n261), .D(n31), .Q(o_cceip2_out_ia_wdata_part2[25]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[26] ( .CK(clk), .CE(n87), .R(n261), .D(n32), .Q(o_cceip2_out_ia_wdata_part2[26]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[27] ( .CK(clk), .CE(n87), .R(n261), .D(n33), .Q(o_cceip2_out_ia_wdata_part2[27]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[28] ( .CK(clk), .CE(n87), .R(n261), .D(n34), .Q(o_cceip2_out_ia_wdata_part2[28]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[29] ( .CK(clk), .CE(n87), .R(n261), .D(n35), .Q(o_cceip2_out_ia_wdata_part2[29]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[30] ( .CK(clk), .CE(n87), .R(n261), .D(n36), .Q(o_cceip2_out_ia_wdata_part2[30]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part2_REG[31] ( .CK(clk), .CE(n87), .R(n261), .D(n37), .Q(o_cceip2_out_ia_wdata_part2[31]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[0] ( .CK(clk), .CE(n86), .R(n261), .D(n6), .Q(o_cceip2_out_ia_wdata_part1[0]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[1] ( .CK(clk), .CE(n86), .R(n261), .D(n7), .Q(o_cceip2_out_ia_wdata_part1[1]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[2] ( .CK(clk), .CE(n86), .R(n261), .D(n8), .Q(o_cceip2_out_ia_wdata_part1[2]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[3] ( .CK(clk), .CE(n86), .R(n261), .D(n9), .Q(o_cceip2_out_ia_wdata_part1[3]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[4] ( .CK(clk), .CE(n86), .R(n261), .D(n10), .Q(o_cceip2_out_ia_wdata_part1[4]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[5] ( .CK(clk), .CE(n86), .R(n261), .D(n11), .Q(o_cceip2_out_ia_wdata_part1[5]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[6] ( .CK(clk), .CE(n86), .R(n261), .D(n12), .Q(o_cceip2_out_ia_wdata_part1[6]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[7] ( .CK(clk), .CE(n86), .R(n261), .D(n13), .Q(o_cceip2_out_ia_wdata_part1[7]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[8] ( .CK(clk), .CE(n86), .R(n261), .D(n14), .Q(o_cceip2_out_ia_wdata_part1[8]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[9] ( .CK(clk), .CE(n86), .R(n261), .D(n15), .Q(o_cceip2_out_ia_wdata_part1[9]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[10] ( .CK(clk), .CE(n86), .R(n261), .D(n16), .Q(o_cceip2_out_ia_wdata_part1[10]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[11] ( .CK(clk), .CE(n86), .R(n261), .D(n17), .Q(o_cceip2_out_ia_wdata_part1[11]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[12] ( .CK(clk), .CE(n86), .R(n261), .D(n18), .Q(o_cceip2_out_ia_wdata_part1[12]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[13] ( .CK(clk), .CE(n86), .R(n261), .D(n19), .Q(o_cceip2_out_ia_wdata_part1[13]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[14] ( .CK(clk), .CE(n86), .R(n261), .D(n20), .Q(o_cceip2_out_ia_wdata_part1[14]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[15] ( .CK(clk), .CE(n86), .R(n261), .D(n21), .Q(o_cceip2_out_ia_wdata_part1[15]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[16] ( .CK(clk), .CE(n86), .R(n261), .D(n22), .Q(o_cceip2_out_ia_wdata_part1[16]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[17] ( .CK(clk), .CE(n86), .R(n261), .D(n23), .Q(o_cceip2_out_ia_wdata_part1[17]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[18] ( .CK(clk), .CE(n86), .R(n261), .D(n24), .Q(o_cceip2_out_ia_wdata_part1[18]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[19] ( .CK(clk), .CE(n86), .R(n261), .D(n25), .Q(o_cceip2_out_ia_wdata_part1[19]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[20] ( .CK(clk), .CE(n86), .R(n261), .D(n26), .Q(o_cceip2_out_ia_wdata_part1[20]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[21] ( .CK(clk), .CE(n86), .R(n261), .D(n27), .Q(o_cceip2_out_ia_wdata_part1[21]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[22] ( .CK(clk), .CE(n86), .R(n261), .D(n28), .Q(o_cceip2_out_ia_wdata_part1[22]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[23] ( .CK(clk), .CE(n86), .R(n261), .D(n29), .Q(o_cceip2_out_ia_wdata_part1[23]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[24] ( .CK(clk), .CE(n86), .R(n261), .D(n30), .Q(o_cceip2_out_ia_wdata_part1[24]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[25] ( .CK(clk), .CE(n86), .R(n261), .D(n31), .Q(o_cceip2_out_ia_wdata_part1[25]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[26] ( .CK(clk), .CE(n86), .R(n261), .D(n32), .Q(o_cceip2_out_ia_wdata_part1[26]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[27] ( .CK(clk), .CE(n86), .R(n261), .D(n33), .Q(o_cceip2_out_ia_wdata_part1[27]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[28] ( .CK(clk), .CE(n86), .R(n261), .D(n34), .Q(o_cceip2_out_ia_wdata_part1[28]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[29] ( .CK(clk), .CE(n86), .R(n261), .D(n35), .Q(o_cceip2_out_ia_wdata_part1[29]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[30] ( .CK(clk), .CE(n86), .R(n261), .D(n36), .Q(o_cceip2_out_ia_wdata_part1[30]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part1_REG[31] ( .CK(clk), .CE(n86), .R(n261), .D(n37), .Q(o_cceip2_out_ia_wdata_part1[31]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[0] ( .CK(clk), .CE(n85), .R(n261), .D(n6), .Q(o_cceip2_out_ia_wdata_part0[0]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[1] ( .CK(clk), .CE(n85), .R(n261), .D(n7), .Q(o_cceip2_out_ia_wdata_part0[1]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[2] ( .CK(clk), .CE(n85), .R(n261), .D(n8), .Q(o_cceip2_out_ia_wdata_part0[2]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[3] ( .CK(clk), .CE(n85), .R(n261), .D(n9), .Q(o_cceip2_out_ia_wdata_part0[3]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[4] ( .CK(clk), .CE(n85), .R(n261), .D(n10), .Q(o_cceip2_out_ia_wdata_part0[4]));
Q_FDP4EP \o_cceip2_out_ia_wdata_part0_REG[5] ( .CK(clk), .CE(n85), .R(n261), .D(n11), .Q(o_cceip2_out_ia_wdata_part0[5]));
Q_FDP4EP \o_cceip1_out_im_read_done_REG[0] ( .CK(clk), .CE(n84), .R(n261), .D(n36), .Q(o_cceip1_out_im_read_done[0]));
Q_FDP4EP \o_cceip1_out_im_read_done_REG[1] ( .CK(clk), .CE(n84), .R(n261), .D(n37), .Q(o_cceip1_out_im_read_done[1]));
Q_FDP4EP \o_cceip1_out_im_config_REG[0] ( .CK(clk), .CE(n83), .R(n261), .D(n6), .Q(o_cceip1_out_im_config[0]));
Q_FDP4EP \o_cceip1_out_im_config_REG[1] ( .CK(clk), .CE(n83), .R(n261), .D(n7), .Q(o_cceip1_out_im_config[1]));
Q_FDP4EP \o_cceip1_out_im_config_REG[2] ( .CK(clk), .CE(n83), .R(n261), .D(n8), .Q(o_cceip1_out_im_config[2]));
Q_FDP4EP \o_cceip1_out_im_config_REG[3] ( .CK(clk), .CE(n83), .R(n261), .D(n9), .Q(o_cceip1_out_im_config[3]));
Q_FDP4EP \o_cceip1_out_im_config_REG[4] ( .CK(clk), .CE(n83), .R(n261), .D(n10), .Q(o_cceip1_out_im_config[4]));
Q_FDP4EP \o_cceip1_out_im_config_REG[5] ( .CK(clk), .CE(n83), .R(n261), .D(n11), .Q(o_cceip1_out_im_config[5]));
Q_FDP4EP \o_cceip1_out_im_config_REG[6] ( .CK(clk), .CE(n83), .R(n261), .D(n12), .Q(o_cceip1_out_im_config[6]));
Q_FDP4EP \o_cceip1_out_im_config_REG[7] ( .CK(clk), .CE(n83), .R(n261), .D(n13), .Q(o_cceip1_out_im_config[7]));
Q_FDP4EP \o_cceip1_out_im_config_REG[8] ( .CK(clk), .CE(n83), .R(n261), .D(n14), .Q(o_cceip1_out_im_config[8]));
Q_FDP4EP \o_cceip1_out_ia_config_REG[0] ( .CK(clk), .CE(n82), .R(n261), .D(n6), .Q(o_cceip1_out_ia_config[0]));
Q_FDP4EP \o_cceip1_out_ia_config_REG[1] ( .CK(clk), .CE(n82), .R(n261), .D(n7), .Q(o_cceip1_out_ia_config[1]));
Q_FDP4EP \o_cceip1_out_ia_config_REG[2] ( .CK(clk), .CE(n82), .R(n261), .D(n8), .Q(o_cceip1_out_ia_config[2]));
Q_FDP4EP \o_cceip1_out_ia_config_REG[3] ( .CK(clk), .CE(n82), .R(n261), .D(n9), .Q(o_cceip1_out_ia_config[3]));
Q_FDP4EP \o_cceip1_out_ia_config_REG[4] ( .CK(clk), .CE(n82), .R(n261), .D(n10), .Q(o_cceip1_out_ia_config[4]));
Q_FDP4EP \o_cceip1_out_ia_config_REG[5] ( .CK(clk), .CE(n82), .R(n261), .D(n11), .Q(o_cceip1_out_ia_config[5]));
Q_FDP4EP \o_cceip1_out_ia_config_REG[6] ( .CK(clk), .CE(n82), .R(n261), .D(n12), .Q(o_cceip1_out_ia_config[6]));
Q_FDP4EP \o_cceip1_out_ia_config_REG[7] ( .CK(clk), .CE(n82), .R(n261), .D(n13), .Q(o_cceip1_out_ia_config[7]));
Q_FDP4EP \o_cceip1_out_ia_config_REG[8] ( .CK(clk), .CE(n82), .R(n261), .D(n14), .Q(o_cceip1_out_ia_config[8]));
Q_FDP4EP \o_cceip1_out_ia_config_REG[9] ( .CK(clk), .CE(n82), .R(n261), .D(n34), .Q(o_cceip1_out_ia_config[9]));
Q_FDP4EP \o_cceip1_out_ia_config_REG[10] ( .CK(clk), .CE(n82), .R(n261), .D(n35), .Q(o_cceip1_out_ia_config[10]));
Q_FDP4EP \o_cceip1_out_ia_config_REG[11] ( .CK(clk), .CE(n82), .R(n261), .D(n36), .Q(o_cceip1_out_ia_config[11]));
Q_FDP4EP \o_cceip1_out_ia_config_REG[12] ( .CK(clk), .CE(n82), .R(n261), .D(n37), .Q(o_cceip1_out_ia_config[12]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[0] ( .CK(clk), .CE(n81), .R(n261), .D(n6), .Q(o_cceip1_out_ia_wdata_part2[0]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[1] ( .CK(clk), .CE(n81), .R(n261), .D(n7), .Q(o_cceip1_out_ia_wdata_part2[1]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[2] ( .CK(clk), .CE(n81), .R(n261), .D(n8), .Q(o_cceip1_out_ia_wdata_part2[2]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[3] ( .CK(clk), .CE(n81), .R(n261), .D(n9), .Q(o_cceip1_out_ia_wdata_part2[3]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[4] ( .CK(clk), .CE(n81), .R(n261), .D(n10), .Q(o_cceip1_out_ia_wdata_part2[4]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[5] ( .CK(clk), .CE(n81), .R(n261), .D(n11), .Q(o_cceip1_out_ia_wdata_part2[5]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[6] ( .CK(clk), .CE(n81), .R(n261), .D(n12), .Q(o_cceip1_out_ia_wdata_part2[6]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[7] ( .CK(clk), .CE(n81), .R(n261), .D(n13), .Q(o_cceip1_out_ia_wdata_part2[7]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[8] ( .CK(clk), .CE(n81), .R(n261), .D(n14), .Q(o_cceip1_out_ia_wdata_part2[8]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[9] ( .CK(clk), .CE(n81), .R(n261), .D(n15), .Q(o_cceip1_out_ia_wdata_part2[9]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[10] ( .CK(clk), .CE(n81), .R(n261), .D(n16), .Q(o_cceip1_out_ia_wdata_part2[10]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[11] ( .CK(clk), .CE(n81), .R(n261), .D(n17), .Q(o_cceip1_out_ia_wdata_part2[11]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[12] ( .CK(clk), .CE(n81), .R(n261), .D(n18), .Q(o_cceip1_out_ia_wdata_part2[12]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[13] ( .CK(clk), .CE(n81), .R(n261), .D(n19), .Q(o_cceip1_out_ia_wdata_part2[13]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[14] ( .CK(clk), .CE(n81), .R(n261), .D(n20), .Q(o_cceip1_out_ia_wdata_part2[14]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[15] ( .CK(clk), .CE(n81), .R(n261), .D(n21), .Q(o_cceip1_out_ia_wdata_part2[15]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[16] ( .CK(clk), .CE(n81), .R(n261), .D(n22), .Q(o_cceip1_out_ia_wdata_part2[16]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[17] ( .CK(clk), .CE(n81), .R(n261), .D(n23), .Q(o_cceip1_out_ia_wdata_part2[17]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[18] ( .CK(clk), .CE(n81), .R(n261), .D(n24), .Q(o_cceip1_out_ia_wdata_part2[18]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[19] ( .CK(clk), .CE(n81), .R(n261), .D(n25), .Q(o_cceip1_out_ia_wdata_part2[19]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[20] ( .CK(clk), .CE(n81), .R(n261), .D(n26), .Q(o_cceip1_out_ia_wdata_part2[20]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[21] ( .CK(clk), .CE(n81), .R(n261), .D(n27), .Q(o_cceip1_out_ia_wdata_part2[21]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[22] ( .CK(clk), .CE(n81), .R(n261), .D(n28), .Q(o_cceip1_out_ia_wdata_part2[22]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[23] ( .CK(clk), .CE(n81), .R(n261), .D(n29), .Q(o_cceip1_out_ia_wdata_part2[23]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[24] ( .CK(clk), .CE(n81), .R(n261), .D(n30), .Q(o_cceip1_out_ia_wdata_part2[24]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[25] ( .CK(clk), .CE(n81), .R(n261), .D(n31), .Q(o_cceip1_out_ia_wdata_part2[25]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[26] ( .CK(clk), .CE(n81), .R(n261), .D(n32), .Q(o_cceip1_out_ia_wdata_part2[26]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[27] ( .CK(clk), .CE(n81), .R(n261), .D(n33), .Q(o_cceip1_out_ia_wdata_part2[27]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[28] ( .CK(clk), .CE(n81), .R(n261), .D(n34), .Q(o_cceip1_out_ia_wdata_part2[28]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[29] ( .CK(clk), .CE(n81), .R(n261), .D(n35), .Q(o_cceip1_out_ia_wdata_part2[29]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[30] ( .CK(clk), .CE(n81), .R(n261), .D(n36), .Q(o_cceip1_out_ia_wdata_part2[30]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part2_REG[31] ( .CK(clk), .CE(n81), .R(n261), .D(n37), .Q(o_cceip1_out_ia_wdata_part2[31]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[0] ( .CK(clk), .CE(n80), .R(n261), .D(n6), .Q(o_cceip1_out_ia_wdata_part1[0]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[1] ( .CK(clk), .CE(n80), .R(n261), .D(n7), .Q(o_cceip1_out_ia_wdata_part1[1]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[2] ( .CK(clk), .CE(n80), .R(n261), .D(n8), .Q(o_cceip1_out_ia_wdata_part1[2]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[3] ( .CK(clk), .CE(n80), .R(n261), .D(n9), .Q(o_cceip1_out_ia_wdata_part1[3]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[4] ( .CK(clk), .CE(n80), .R(n261), .D(n10), .Q(o_cceip1_out_ia_wdata_part1[4]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[5] ( .CK(clk), .CE(n80), .R(n261), .D(n11), .Q(o_cceip1_out_ia_wdata_part1[5]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[6] ( .CK(clk), .CE(n80), .R(n261), .D(n12), .Q(o_cceip1_out_ia_wdata_part1[6]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[7] ( .CK(clk), .CE(n80), .R(n261), .D(n13), .Q(o_cceip1_out_ia_wdata_part1[7]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[8] ( .CK(clk), .CE(n80), .R(n261), .D(n14), .Q(o_cceip1_out_ia_wdata_part1[8]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[9] ( .CK(clk), .CE(n80), .R(n261), .D(n15), .Q(o_cceip1_out_ia_wdata_part1[9]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[10] ( .CK(clk), .CE(n80), .R(n261), .D(n16), .Q(o_cceip1_out_ia_wdata_part1[10]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[11] ( .CK(clk), .CE(n80), .R(n261), .D(n17), .Q(o_cceip1_out_ia_wdata_part1[11]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[12] ( .CK(clk), .CE(n80), .R(n261), .D(n18), .Q(o_cceip1_out_ia_wdata_part1[12]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[13] ( .CK(clk), .CE(n80), .R(n261), .D(n19), .Q(o_cceip1_out_ia_wdata_part1[13]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[14] ( .CK(clk), .CE(n80), .R(n261), .D(n20), .Q(o_cceip1_out_ia_wdata_part1[14]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[15] ( .CK(clk), .CE(n80), .R(n261), .D(n21), .Q(o_cceip1_out_ia_wdata_part1[15]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[16] ( .CK(clk), .CE(n80), .R(n261), .D(n22), .Q(o_cceip1_out_ia_wdata_part1[16]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[17] ( .CK(clk), .CE(n80), .R(n261), .D(n23), .Q(o_cceip1_out_ia_wdata_part1[17]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[18] ( .CK(clk), .CE(n80), .R(n261), .D(n24), .Q(o_cceip1_out_ia_wdata_part1[18]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[19] ( .CK(clk), .CE(n80), .R(n261), .D(n25), .Q(o_cceip1_out_ia_wdata_part1[19]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[20] ( .CK(clk), .CE(n80), .R(n261), .D(n26), .Q(o_cceip1_out_ia_wdata_part1[20]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[21] ( .CK(clk), .CE(n80), .R(n261), .D(n27), .Q(o_cceip1_out_ia_wdata_part1[21]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[22] ( .CK(clk), .CE(n80), .R(n261), .D(n28), .Q(o_cceip1_out_ia_wdata_part1[22]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[23] ( .CK(clk), .CE(n80), .R(n261), .D(n29), .Q(o_cceip1_out_ia_wdata_part1[23]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[24] ( .CK(clk), .CE(n80), .R(n261), .D(n30), .Q(o_cceip1_out_ia_wdata_part1[24]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[25] ( .CK(clk), .CE(n80), .R(n261), .D(n31), .Q(o_cceip1_out_ia_wdata_part1[25]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[26] ( .CK(clk), .CE(n80), .R(n261), .D(n32), .Q(o_cceip1_out_ia_wdata_part1[26]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[27] ( .CK(clk), .CE(n80), .R(n261), .D(n33), .Q(o_cceip1_out_ia_wdata_part1[27]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[28] ( .CK(clk), .CE(n80), .R(n261), .D(n34), .Q(o_cceip1_out_ia_wdata_part1[28]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[29] ( .CK(clk), .CE(n80), .R(n261), .D(n35), .Q(o_cceip1_out_ia_wdata_part1[29]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[30] ( .CK(clk), .CE(n80), .R(n261), .D(n36), .Q(o_cceip1_out_ia_wdata_part1[30]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part1_REG[31] ( .CK(clk), .CE(n80), .R(n261), .D(n37), .Q(o_cceip1_out_ia_wdata_part1[31]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[0] ( .CK(clk), .CE(n79), .R(n261), .D(n6), .Q(o_cceip1_out_ia_wdata_part0[0]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[1] ( .CK(clk), .CE(n79), .R(n261), .D(n7), .Q(o_cceip1_out_ia_wdata_part0[1]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[2] ( .CK(clk), .CE(n79), .R(n261), .D(n8), .Q(o_cceip1_out_ia_wdata_part0[2]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[3] ( .CK(clk), .CE(n79), .R(n261), .D(n9), .Q(o_cceip1_out_ia_wdata_part0[3]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[4] ( .CK(clk), .CE(n79), .R(n261), .D(n10), .Q(o_cceip1_out_ia_wdata_part0[4]));
Q_FDP4EP \o_cceip1_out_ia_wdata_part0_REG[5] ( .CK(clk), .CE(n79), .R(n261), .D(n11), .Q(o_cceip1_out_ia_wdata_part0[5]));
Q_FDP4EP \o_cceip0_out_im_read_done_REG[0] ( .CK(clk), .CE(n78), .R(n261), .D(n36), .Q(o_cceip0_out_im_read_done[0]));
Q_FDP4EP \o_cceip0_out_im_read_done_REG[1] ( .CK(clk), .CE(n78), .R(n261), .D(n37), .Q(o_cceip0_out_im_read_done[1]));
Q_FDP4EP \o_cceip0_out_im_config_REG[0] ( .CK(clk), .CE(n77), .R(n261), .D(n6), .Q(o_cceip0_out_im_config[0]));
Q_FDP4EP \o_cceip0_out_im_config_REG[1] ( .CK(clk), .CE(n77), .R(n261), .D(n7), .Q(o_cceip0_out_im_config[1]));
Q_FDP4EP \o_cceip0_out_im_config_REG[2] ( .CK(clk), .CE(n77), .R(n261), .D(n8), .Q(o_cceip0_out_im_config[2]));
Q_FDP4EP \o_cceip0_out_im_config_REG[3] ( .CK(clk), .CE(n77), .R(n261), .D(n9), .Q(o_cceip0_out_im_config[3]));
Q_FDP4EP \o_cceip0_out_im_config_REG[4] ( .CK(clk), .CE(n77), .R(n261), .D(n10), .Q(o_cceip0_out_im_config[4]));
Q_FDP4EP \o_cceip0_out_im_config_REG[5] ( .CK(clk), .CE(n77), .R(n261), .D(n11), .Q(o_cceip0_out_im_config[5]));
Q_FDP4EP \o_cceip0_out_im_config_REG[6] ( .CK(clk), .CE(n77), .R(n261), .D(n12), .Q(o_cceip0_out_im_config[6]));
Q_FDP4EP \o_cceip0_out_im_config_REG[7] ( .CK(clk), .CE(n77), .R(n261), .D(n13), .Q(o_cceip0_out_im_config[7]));
Q_FDP4EP \o_cceip0_out_im_config_REG[8] ( .CK(clk), .CE(n77), .R(n261), .D(n14), .Q(o_cceip0_out_im_config[8]));
Q_FDP4EP \o_cceip0_out_ia_config_REG[0] ( .CK(clk), .CE(n76), .R(n261), .D(n6), .Q(o_cceip0_out_ia_config[0]));
Q_FDP4EP \o_cceip0_out_ia_config_REG[1] ( .CK(clk), .CE(n76), .R(n261), .D(n7), .Q(o_cceip0_out_ia_config[1]));
Q_FDP4EP \o_cceip0_out_ia_config_REG[2] ( .CK(clk), .CE(n76), .R(n261), .D(n8), .Q(o_cceip0_out_ia_config[2]));
Q_FDP4EP \o_cceip0_out_ia_config_REG[3] ( .CK(clk), .CE(n76), .R(n261), .D(n9), .Q(o_cceip0_out_ia_config[3]));
Q_FDP4EP \o_cceip0_out_ia_config_REG[4] ( .CK(clk), .CE(n76), .R(n261), .D(n10), .Q(o_cceip0_out_ia_config[4]));
Q_FDP4EP \o_cceip0_out_ia_config_REG[5] ( .CK(clk), .CE(n76), .R(n261), .D(n11), .Q(o_cceip0_out_ia_config[5]));
Q_FDP4EP \o_cceip0_out_ia_config_REG[6] ( .CK(clk), .CE(n76), .R(n261), .D(n12), .Q(o_cceip0_out_ia_config[6]));
Q_FDP4EP \o_cceip0_out_ia_config_REG[7] ( .CK(clk), .CE(n76), .R(n261), .D(n13), .Q(o_cceip0_out_ia_config[7]));
Q_FDP4EP \o_cceip0_out_ia_config_REG[8] ( .CK(clk), .CE(n76), .R(n261), .D(n14), .Q(o_cceip0_out_ia_config[8]));
Q_FDP4EP \o_cceip0_out_ia_config_REG[9] ( .CK(clk), .CE(n76), .R(n261), .D(n34), .Q(o_cceip0_out_ia_config[9]));
Q_FDP4EP \o_cceip0_out_ia_config_REG[10] ( .CK(clk), .CE(n76), .R(n261), .D(n35), .Q(o_cceip0_out_ia_config[10]));
Q_FDP4EP \o_cceip0_out_ia_config_REG[11] ( .CK(clk), .CE(n76), .R(n261), .D(n36), .Q(o_cceip0_out_ia_config[11]));
Q_FDP4EP \o_cceip0_out_ia_config_REG[12] ( .CK(clk), .CE(n76), .R(n261), .D(n37), .Q(o_cceip0_out_ia_config[12]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[0] ( .CK(clk), .CE(n75), .R(n261), .D(n6), .Q(o_cceip0_out_ia_wdata_part2[0]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[1] ( .CK(clk), .CE(n75), .R(n261), .D(n7), .Q(o_cceip0_out_ia_wdata_part2[1]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[2] ( .CK(clk), .CE(n75), .R(n261), .D(n8), .Q(o_cceip0_out_ia_wdata_part2[2]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[3] ( .CK(clk), .CE(n75), .R(n261), .D(n9), .Q(o_cceip0_out_ia_wdata_part2[3]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[4] ( .CK(clk), .CE(n75), .R(n261), .D(n10), .Q(o_cceip0_out_ia_wdata_part2[4]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[5] ( .CK(clk), .CE(n75), .R(n261), .D(n11), .Q(o_cceip0_out_ia_wdata_part2[5]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[6] ( .CK(clk), .CE(n75), .R(n261), .D(n12), .Q(o_cceip0_out_ia_wdata_part2[6]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[7] ( .CK(clk), .CE(n75), .R(n261), .D(n13), .Q(o_cceip0_out_ia_wdata_part2[7]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[8] ( .CK(clk), .CE(n75), .R(n261), .D(n14), .Q(o_cceip0_out_ia_wdata_part2[8]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[9] ( .CK(clk), .CE(n75), .R(n261), .D(n15), .Q(o_cceip0_out_ia_wdata_part2[9]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[10] ( .CK(clk), .CE(n75), .R(n261), .D(n16), .Q(o_cceip0_out_ia_wdata_part2[10]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[11] ( .CK(clk), .CE(n75), .R(n261), .D(n17), .Q(o_cceip0_out_ia_wdata_part2[11]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[12] ( .CK(clk), .CE(n75), .R(n261), .D(n18), .Q(o_cceip0_out_ia_wdata_part2[12]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[13] ( .CK(clk), .CE(n75), .R(n261), .D(n19), .Q(o_cceip0_out_ia_wdata_part2[13]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[14] ( .CK(clk), .CE(n75), .R(n261), .D(n20), .Q(o_cceip0_out_ia_wdata_part2[14]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[15] ( .CK(clk), .CE(n75), .R(n261), .D(n21), .Q(o_cceip0_out_ia_wdata_part2[15]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[16] ( .CK(clk), .CE(n75), .R(n261), .D(n22), .Q(o_cceip0_out_ia_wdata_part2[16]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[17] ( .CK(clk), .CE(n75), .R(n261), .D(n23), .Q(o_cceip0_out_ia_wdata_part2[17]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[18] ( .CK(clk), .CE(n75), .R(n261), .D(n24), .Q(o_cceip0_out_ia_wdata_part2[18]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[19] ( .CK(clk), .CE(n75), .R(n261), .D(n25), .Q(o_cceip0_out_ia_wdata_part2[19]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[20] ( .CK(clk), .CE(n75), .R(n261), .D(n26), .Q(o_cceip0_out_ia_wdata_part2[20]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[21] ( .CK(clk), .CE(n75), .R(n261), .D(n27), .Q(o_cceip0_out_ia_wdata_part2[21]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[22] ( .CK(clk), .CE(n75), .R(n261), .D(n28), .Q(o_cceip0_out_ia_wdata_part2[22]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[23] ( .CK(clk), .CE(n75), .R(n261), .D(n29), .Q(o_cceip0_out_ia_wdata_part2[23]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[24] ( .CK(clk), .CE(n75), .R(n261), .D(n30), .Q(o_cceip0_out_ia_wdata_part2[24]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[25] ( .CK(clk), .CE(n75), .R(n261), .D(n31), .Q(o_cceip0_out_ia_wdata_part2[25]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[26] ( .CK(clk), .CE(n75), .R(n261), .D(n32), .Q(o_cceip0_out_ia_wdata_part2[26]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[27] ( .CK(clk), .CE(n75), .R(n261), .D(n33), .Q(o_cceip0_out_ia_wdata_part2[27]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[28] ( .CK(clk), .CE(n75), .R(n261), .D(n34), .Q(o_cceip0_out_ia_wdata_part2[28]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[29] ( .CK(clk), .CE(n75), .R(n261), .D(n35), .Q(o_cceip0_out_ia_wdata_part2[29]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[30] ( .CK(clk), .CE(n75), .R(n261), .D(n36), .Q(o_cceip0_out_ia_wdata_part2[30]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part2_REG[31] ( .CK(clk), .CE(n75), .R(n261), .D(n37), .Q(o_cceip0_out_ia_wdata_part2[31]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[0] ( .CK(clk), .CE(n74), .R(n261), .D(n6), .Q(o_cceip0_out_ia_wdata_part1[0]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[1] ( .CK(clk), .CE(n74), .R(n261), .D(n7), .Q(o_cceip0_out_ia_wdata_part1[1]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[2] ( .CK(clk), .CE(n74), .R(n261), .D(n8), .Q(o_cceip0_out_ia_wdata_part1[2]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[3] ( .CK(clk), .CE(n74), .R(n261), .D(n9), .Q(o_cceip0_out_ia_wdata_part1[3]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[4] ( .CK(clk), .CE(n74), .R(n261), .D(n10), .Q(o_cceip0_out_ia_wdata_part1[4]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[5] ( .CK(clk), .CE(n74), .R(n261), .D(n11), .Q(o_cceip0_out_ia_wdata_part1[5]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[6] ( .CK(clk), .CE(n74), .R(n261), .D(n12), .Q(o_cceip0_out_ia_wdata_part1[6]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[7] ( .CK(clk), .CE(n74), .R(n261), .D(n13), .Q(o_cceip0_out_ia_wdata_part1[7]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[8] ( .CK(clk), .CE(n74), .R(n261), .D(n14), .Q(o_cceip0_out_ia_wdata_part1[8]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[9] ( .CK(clk), .CE(n74), .R(n261), .D(n15), .Q(o_cceip0_out_ia_wdata_part1[9]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[10] ( .CK(clk), .CE(n74), .R(n261), .D(n16), .Q(o_cceip0_out_ia_wdata_part1[10]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[11] ( .CK(clk), .CE(n74), .R(n261), .D(n17), .Q(o_cceip0_out_ia_wdata_part1[11]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[12] ( .CK(clk), .CE(n74), .R(n261), .D(n18), .Q(o_cceip0_out_ia_wdata_part1[12]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[13] ( .CK(clk), .CE(n74), .R(n261), .D(n19), .Q(o_cceip0_out_ia_wdata_part1[13]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[14] ( .CK(clk), .CE(n74), .R(n261), .D(n20), .Q(o_cceip0_out_ia_wdata_part1[14]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[15] ( .CK(clk), .CE(n74), .R(n261), .D(n21), .Q(o_cceip0_out_ia_wdata_part1[15]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[16] ( .CK(clk), .CE(n74), .R(n261), .D(n22), .Q(o_cceip0_out_ia_wdata_part1[16]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[17] ( .CK(clk), .CE(n74), .R(n261), .D(n23), .Q(o_cceip0_out_ia_wdata_part1[17]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[18] ( .CK(clk), .CE(n74), .R(n261), .D(n24), .Q(o_cceip0_out_ia_wdata_part1[18]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[19] ( .CK(clk), .CE(n74), .R(n261), .D(n25), .Q(o_cceip0_out_ia_wdata_part1[19]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[20] ( .CK(clk), .CE(n74), .R(n261), .D(n26), .Q(o_cceip0_out_ia_wdata_part1[20]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[21] ( .CK(clk), .CE(n74), .R(n261), .D(n27), .Q(o_cceip0_out_ia_wdata_part1[21]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[22] ( .CK(clk), .CE(n74), .R(n261), .D(n28), .Q(o_cceip0_out_ia_wdata_part1[22]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[23] ( .CK(clk), .CE(n74), .R(n261), .D(n29), .Q(o_cceip0_out_ia_wdata_part1[23]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[24] ( .CK(clk), .CE(n74), .R(n261), .D(n30), .Q(o_cceip0_out_ia_wdata_part1[24]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[25] ( .CK(clk), .CE(n74), .R(n261), .D(n31), .Q(o_cceip0_out_ia_wdata_part1[25]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[26] ( .CK(clk), .CE(n74), .R(n261), .D(n32), .Q(o_cceip0_out_ia_wdata_part1[26]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[27] ( .CK(clk), .CE(n74), .R(n261), .D(n33), .Q(o_cceip0_out_ia_wdata_part1[27]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[28] ( .CK(clk), .CE(n74), .R(n261), .D(n34), .Q(o_cceip0_out_ia_wdata_part1[28]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[29] ( .CK(clk), .CE(n74), .R(n261), .D(n35), .Q(o_cceip0_out_ia_wdata_part1[29]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[30] ( .CK(clk), .CE(n74), .R(n261), .D(n36), .Q(o_cceip0_out_ia_wdata_part1[30]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part1_REG[31] ( .CK(clk), .CE(n74), .R(n261), .D(n37), .Q(o_cceip0_out_ia_wdata_part1[31]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[0] ( .CK(clk), .CE(n73), .R(n261), .D(n6), .Q(o_cceip0_out_ia_wdata_part0[0]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[1] ( .CK(clk), .CE(n73), .R(n261), .D(n7), .Q(o_cceip0_out_ia_wdata_part0[1]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[2] ( .CK(clk), .CE(n73), .R(n261), .D(n8), .Q(o_cceip0_out_ia_wdata_part0[2]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[3] ( .CK(clk), .CE(n73), .R(n261), .D(n9), .Q(o_cceip0_out_ia_wdata_part0[3]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[4] ( .CK(clk), .CE(n73), .R(n261), .D(n10), .Q(o_cceip0_out_ia_wdata_part0[4]));
Q_FDP4EP \o_cceip0_out_ia_wdata_part0_REG[5] ( .CK(clk), .CE(n73), .R(n261), .D(n11), .Q(o_cceip0_out_ia_wdata_part0[5]));
Q_FDP4EP \o_spare_config_REG[0] ( .CK(clk), .CE(n72), .R(n261), .D(n6), .Q(o_spare_config[0]));
Q_FDP4EP \o_spare_config_REG[1] ( .CK(clk), .CE(n72), .R(n261), .D(n7), .Q(o_spare_config[1]));
Q_FDP4EP \o_spare_config_REG[2] ( .CK(clk), .CE(n72), .R(n261), .D(n8), .Q(o_spare_config[2]));
Q_FDP4EP \o_spare_config_REG[3] ( .CK(clk), .CE(n72), .R(n261), .D(n9), .Q(o_spare_config[3]));
Q_FDP4EP \o_spare_config_REG[4] ( .CK(clk), .CE(n72), .R(n261), .D(n10), .Q(o_spare_config[4]));
Q_FDP4EP \o_spare_config_REG[5] ( .CK(clk), .CE(n72), .R(n261), .D(n11), .Q(o_spare_config[5]));
Q_FDP4EP \o_spare_config_REG[6] ( .CK(clk), .CE(n72), .R(n261), .D(n12), .Q(o_spare_config[6]));
Q_FDP4EP \o_spare_config_REG[7] ( .CK(clk), .CE(n72), .R(n261), .D(n13), .Q(o_spare_config[7]));
Q_FDP4EP \o_spare_config_REG[8] ( .CK(clk), .CE(n72), .R(n261), .D(n14), .Q(o_spare_config[8]));
Q_FDP4EP \o_spare_config_REG[9] ( .CK(clk), .CE(n72), .R(n261), .D(n15), .Q(o_spare_config[9]));
Q_FDP4EP \o_spare_config_REG[10] ( .CK(clk), .CE(n72), .R(n261), .D(n16), .Q(o_spare_config[10]));
Q_FDP4EP \o_spare_config_REG[11] ( .CK(clk), .CE(n72), .R(n261), .D(n17), .Q(o_spare_config[11]));
Q_FDP4EP \o_spare_config_REG[12] ( .CK(clk), .CE(n72), .R(n261), .D(n18), .Q(o_spare_config[12]));
Q_FDP4EP \o_spare_config_REG[13] ( .CK(clk), .CE(n72), .R(n261), .D(n19), .Q(o_spare_config[13]));
Q_FDP4EP \o_spare_config_REG[14] ( .CK(clk), .CE(n72), .R(n261), .D(n20), .Q(o_spare_config[14]));
Q_FDP4EP \o_spare_config_REG[15] ( .CK(clk), .CE(n72), .R(n261), .D(n21), .Q(o_spare_config[15]));
Q_FDP4EP \o_spare_config_REG[16] ( .CK(clk), .CE(n72), .R(n261), .D(n22), .Q(o_spare_config[16]));
Q_FDP4EP \o_spare_config_REG[17] ( .CK(clk), .CE(n72), .R(n261), .D(n23), .Q(o_spare_config[17]));
Q_FDP4EP \o_spare_config_REG[18] ( .CK(clk), .CE(n72), .R(n261), .D(n24), .Q(o_spare_config[18]));
Q_FDP4EP \o_spare_config_REG[19] ( .CK(clk), .CE(n72), .R(n261), .D(n25), .Q(o_spare_config[19]));
Q_FDP4EP \o_spare_config_REG[20] ( .CK(clk), .CE(n72), .R(n261), .D(n26), .Q(o_spare_config[20]));
Q_FDP4EP \o_spare_config_REG[21] ( .CK(clk), .CE(n72), .R(n261), .D(n27), .Q(o_spare_config[21]));
Q_FDP4EP \o_spare_config_REG[22] ( .CK(clk), .CE(n72), .R(n261), .D(n28), .Q(o_spare_config[22]));
Q_FDP4EP \o_spare_config_REG[23] ( .CK(clk), .CE(n72), .R(n261), .D(n29), .Q(o_spare_config[23]));
Q_FDP4EP \o_spare_config_REG[24] ( .CK(clk), .CE(n72), .R(n261), .D(n30), .Q(o_spare_config[24]));
Q_FDP4EP \o_spare_config_REG[25] ( .CK(clk), .CE(n72), .R(n261), .D(n31), .Q(o_spare_config[25]));
Q_FDP4EP \o_spare_config_REG[26] ( .CK(clk), .CE(n72), .R(n261), .D(n32), .Q(o_spare_config[26]));
Q_FDP4EP \o_spare_config_REG[27] ( .CK(clk), .CE(n72), .R(n261), .D(n33), .Q(o_spare_config[27]));
Q_FDP4EP \o_spare_config_REG[28] ( .CK(clk), .CE(n72), .R(n261), .D(n34), .Q(o_spare_config[28]));
Q_FDP4EP \o_spare_config_REG[29] ( .CK(clk), .CE(n72), .R(n261), .D(n35), .Q(o_spare_config[29]));
Q_FDP4EP \o_spare_config_REG[30] ( .CK(clk), .CE(n72), .R(n261), .D(n36), .Q(o_spare_config[30]));
Q_FDP4EP \o_spare_config_REG[31] ( .CK(clk), .CE(n72), .R(n261), .D(n37), .Q(o_spare_config[31]));
endmodule
