architecture module of ixc_uClkGen is
  -- quickturn CVASTRPROP MODULE HDLICE PROP_IXCOM_MOD TRUE
  signal DUMMY0 : std_logic ;

begin
  uclk <= DUMMY0 ;
end module;
