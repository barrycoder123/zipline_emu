
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
(* celldefine = 1 *) 
module sync_fifo ( dout, full, empty, clk, rst_n, din, wr_en, rd_en, 
	space_avail);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output [95:0] dout;
output full;
output empty;
input clk;
input rst_n;
input [95:0] din;
input wr_en;
input rd_en;
output [3:0] space_avail;
wire [3:0] wr_ptr_nxt;
wire [3:0] rd_ptr_nxt;
wire full_i;
wire empty_i;
wire [95:0] default_data;
wire [3:0] wr_ptr_r;
wire [3:0] rd_ptr_r;
wire [31:0] i;
wire [95:0] dout_i;
wire [95:0] dout_r;
wire hit_flag;
supply1 n1;
Q_BUF U0 ( .A(n1), .Z(hit_flag));
Q_BUF U1 ( .A(dout_i[0]), .Z(dout_r[0]));
Q_BUF U2 ( .A(dout_i[1]), .Z(dout_r[1]));
Q_BUF U3 ( .A(dout_i[2]), .Z(dout_r[2]));
Q_BUF U4 ( .A(dout_i[3]), .Z(dout_r[3]));
Q_BUF U5 ( .A(dout_i[4]), .Z(dout_r[4]));
Q_BUF U6 ( .A(dout_i[5]), .Z(dout_r[5]));
Q_BUF U7 ( .A(dout_i[6]), .Z(dout_r[6]));
Q_BUF U8 ( .A(dout_i[7]), .Z(dout_r[7]));
Q_BUF U9 ( .A(dout_i[8]), .Z(dout_r[8]));
Q_BUF U10 ( .A(dout_i[9]), .Z(dout_r[9]));
Q_BUF U11 ( .A(dout_i[10]), .Z(dout_r[10]));
Q_BUF U12 ( .A(dout_i[11]), .Z(dout_r[11]));
Q_BUF U13 ( .A(dout_i[12]), .Z(dout_r[12]));
Q_BUF U14 ( .A(dout_i[13]), .Z(dout_r[13]));
Q_BUF U15 ( .A(dout_i[14]), .Z(dout_r[14]));
Q_BUF U16 ( .A(dout_i[15]), .Z(dout_r[15]));
Q_BUF U17 ( .A(dout_i[16]), .Z(dout_r[16]));
Q_BUF U18 ( .A(dout_i[17]), .Z(dout_r[17]));
Q_BUF U19 ( .A(dout_i[18]), .Z(dout_r[18]));
Q_BUF U20 ( .A(dout_i[19]), .Z(dout_r[19]));
Q_BUF U21 ( .A(dout_i[20]), .Z(dout_r[20]));
Q_BUF U22 ( .A(dout_i[21]), .Z(dout_r[21]));
Q_BUF U23 ( .A(dout_i[22]), .Z(dout_r[22]));
Q_BUF U24 ( .A(dout_i[23]), .Z(dout_r[23]));
Q_BUF U25 ( .A(dout_i[24]), .Z(dout_r[24]));
Q_BUF U26 ( .A(dout_i[25]), .Z(dout_r[25]));
Q_BUF U27 ( .A(dout_i[26]), .Z(dout_r[26]));
Q_BUF U28 ( .A(dout_i[27]), .Z(dout_r[27]));
Q_BUF U29 ( .A(dout_i[28]), .Z(dout_r[28]));
Q_BUF U30 ( .A(dout_i[29]), .Z(dout_r[29]));
Q_BUF U31 ( .A(dout_i[30]), .Z(dout_r[30]));
Q_BUF U32 ( .A(dout_i[31]), .Z(dout_r[31]));
Q_BUF U33 ( .A(dout_i[32]), .Z(dout_r[32]));
Q_BUF U34 ( .A(dout_i[33]), .Z(dout_r[33]));
Q_BUF U35 ( .A(dout_i[34]), .Z(dout_r[34]));
Q_BUF U36 ( .A(dout_i[35]), .Z(dout_r[35]));
Q_BUF U37 ( .A(dout_i[36]), .Z(dout_r[36]));
Q_BUF U38 ( .A(dout_i[37]), .Z(dout_r[37]));
Q_BUF U39 ( .A(dout_i[38]), .Z(dout_r[38]));
Q_BUF U40 ( .A(dout_i[39]), .Z(dout_r[39]));
Q_BUF U41 ( .A(dout_i[40]), .Z(dout_r[40]));
Q_BUF U42 ( .A(dout_i[41]), .Z(dout_r[41]));
Q_BUF U43 ( .A(dout_i[42]), .Z(dout_r[42]));
Q_BUF U44 ( .A(dout_i[43]), .Z(dout_r[43]));
Q_BUF U45 ( .A(dout_i[44]), .Z(dout_r[44]));
Q_BUF U46 ( .A(dout_i[45]), .Z(dout_r[45]));
Q_BUF U47 ( .A(dout_i[46]), .Z(dout_r[46]));
Q_BUF U48 ( .A(dout_i[47]), .Z(dout_r[47]));
Q_BUF U49 ( .A(dout_i[48]), .Z(dout_r[48]));
Q_BUF U50 ( .A(dout_i[49]), .Z(dout_r[49]));
Q_BUF U51 ( .A(dout_i[50]), .Z(dout_r[50]));
Q_BUF U52 ( .A(dout_i[51]), .Z(dout_r[51]));
Q_BUF U53 ( .A(dout_i[52]), .Z(dout_r[52]));
Q_BUF U54 ( .A(dout_i[53]), .Z(dout_r[53]));
Q_BUF U55 ( .A(dout_i[54]), .Z(dout_r[54]));
Q_BUF U56 ( .A(dout_i[55]), .Z(dout_r[55]));
Q_BUF U57 ( .A(dout_i[56]), .Z(dout_r[56]));
Q_BUF U58 ( .A(dout_i[57]), .Z(dout_r[57]));
Q_BUF U59 ( .A(dout_i[58]), .Z(dout_r[58]));
Q_BUF U60 ( .A(dout_i[59]), .Z(dout_r[59]));
Q_BUF U61 ( .A(dout_i[60]), .Z(dout_r[60]));
Q_BUF U62 ( .A(dout_i[61]), .Z(dout_r[61]));
Q_BUF U63 ( .A(dout_i[62]), .Z(dout_r[62]));
Q_BUF U64 ( .A(dout_i[63]), .Z(dout_r[63]));
Q_BUF U65 ( .A(dout_i[64]), .Z(dout_r[64]));
Q_BUF U66 ( .A(dout_i[65]), .Z(dout_r[65]));
Q_BUF U67 ( .A(dout_i[66]), .Z(dout_r[66]));
Q_BUF U68 ( .A(dout_i[67]), .Z(dout_r[67]));
Q_BUF U69 ( .A(dout_i[68]), .Z(dout_r[68]));
Q_BUF U70 ( .A(dout_i[69]), .Z(dout_r[69]));
Q_BUF U71 ( .A(dout_i[70]), .Z(dout_r[70]));
Q_BUF U72 ( .A(dout_i[71]), .Z(dout_r[71]));
Q_BUF U73 ( .A(dout_i[72]), .Z(dout_r[72]));
Q_BUF U74 ( .A(dout_i[73]), .Z(dout_r[73]));
Q_BUF U75 ( .A(dout_i[74]), .Z(dout_r[74]));
Q_BUF U76 ( .A(dout_i[75]), .Z(dout_r[75]));
Q_BUF U77 ( .A(dout_i[76]), .Z(dout_r[76]));
Q_BUF U78 ( .A(dout_i[77]), .Z(dout_r[77]));
Q_BUF U79 ( .A(dout_i[78]), .Z(dout_r[78]));
Q_BUF U80 ( .A(dout_i[79]), .Z(dout_r[79]));
Q_BUF U81 ( .A(dout_i[80]), .Z(dout_r[80]));
Q_BUF U82 ( .A(dout_i[81]), .Z(dout_r[81]));
Q_BUF U83 ( .A(dout_i[82]), .Z(dout_r[82]));
Q_BUF U84 ( .A(dout_i[83]), .Z(dout_r[83]));
Q_BUF U85 ( .A(dout_i[84]), .Z(dout_r[84]));
Q_BUF U86 ( .A(dout_i[85]), .Z(dout_r[85]));
Q_BUF U87 ( .A(dout_i[86]), .Z(dout_r[86]));
Q_BUF U88 ( .A(dout_i[87]), .Z(dout_r[87]));
Q_BUF U89 ( .A(dout_i[88]), .Z(dout_r[88]));
Q_BUF U90 ( .A(dout_i[89]), .Z(dout_r[89]));
Q_BUF U91 ( .A(dout_i[90]), .Z(dout_r[90]));
Q_BUF U92 ( .A(dout_i[91]), .Z(dout_r[91]));
Q_BUF U93 ( .A(dout_i[92]), .Z(dout_r[92]));
Q_BUF U94 ( .A(dout_i[93]), .Z(dout_r[93]));
Q_BUF U95 ( .A(dout_i[94]), .Z(dout_r[94]));
Q_BUF U96 ( .A(dout_i[95]), .Z(dout_r[95]));
ixc_assign_96 \genblk1._zz_strnp_0 ( default_data[95:0], { \mem_r[0][95] , 
	\mem_r[0][94] , \mem_r[0][93] , \mem_r[0][92] , \mem_r[0][91] , 
	\mem_r[0][90] , \mem_r[0][89] , \mem_r[0][88] , \mem_r[0][87] , 
	\mem_r[0][86] , \mem_r[0][85] , \mem_r[0][84] , \mem_r[0][83] , 
	\mem_r[0][82] , \mem_r[0][81] , \mem_r[0][80] , \mem_r[0][79] , 
	\mem_r[0][78] , \mem_r[0][77] , \mem_r[0][76] , \mem_r[0][75] , 
	\mem_r[0][74] , \mem_r[0][73] , \mem_r[0][72] , \mem_r[0][71] , 
	\mem_r[0][70] , \mem_r[0][69] , \mem_r[0][68] , \mem_r[0][67] , 
	\mem_r[0][66] , \mem_r[0][65] , \mem_r[0][64] , \mem_r[0][63] , 
	\mem_r[0][62] , \mem_r[0][61] , \mem_r[0][60] , \mem_r[0][59] , 
	\mem_r[0][58] , \mem_r[0][57] , \mem_r[0][56] , \mem_r[0][55] , 
	\mem_r[0][54] , \mem_r[0][53] , \mem_r[0][52] , \mem_r[0][51] , 
	\mem_r[0][50] , \mem_r[0][49] , \mem_r[0][48] , \mem_r[0][47] , 
	\mem_r[0][46] , \mem_r[0][45] , \mem_r[0][44] , \mem_r[0][43] , 
	\mem_r[0][42] , \mem_r[0][41] , \mem_r[0][40] , \mem_r[0][39] , 
	\mem_r[0][38] , \mem_r[0][37] , \mem_r[0][36] , \mem_r[0][35] , 
	\mem_r[0][34] , \mem_r[0][33] , \mem_r[0][32] , \mem_r[0][31] , 
	\mem_r[0][30] , \mem_r[0][29] , \mem_r[0][28] , \mem_r[0][27] , 
	\mem_r[0][26] , \mem_r[0][25] , \mem_r[0][24] , \mem_r[0][23] , 
	\mem_r[0][22] , \mem_r[0][21] , \mem_r[0][20] , \mem_r[0][19] , 
	\mem_r[0][18] , \mem_r[0][17] , \mem_r[0][16] , \mem_r[0][15] , 
	\mem_r[0][14] , \mem_r[0][13] , \mem_r[0][12] , \mem_r[0][11] , 
	\mem_r[0][10] , \mem_r[0][9] , \mem_r[0][8] , \mem_r[0][7] , 
	\mem_r[0][6] , \mem_r[0][5] , \mem_r[0][4] , \mem_r[0][3] , 
	\mem_r[0][2] , \mem_r[0][1] , \mem_r[0][0] });
ixc_assign_4 _zz_strnp_4 ( space_avail[3:0], { n2, n3, n4, n5});
ixc_assign_96 _zz_strnp_3 ( dout[95:0], dout_r[95:0]);
ixc_assign _zz_strnp_2 ( empty, empty_i);
ixc_assign _zz_strnp_1 ( full, full_i);
Q_AN02 U102 ( .A0(n6), .A1(n12), .Z(empty_i));
Q_AN03 U103 ( .A0(n10), .A1(n8), .A2(n7), .Z(n12));
Q_AN02 U104 ( .A0(n9), .A1(n11), .Z(full_i));
Q_INV U105 ( .A(n10), .Z(n11));
Q_XNR2 U106 ( .A0(rd_ptr_r[3]), .A1(wr_ptr_r[3]), .Z(n10));
Q_AN03 U107 ( .A0(n6), .A1(n7), .A2(n8), .Z(n9));
Q_XNR2 U108 ( .A0(rd_ptr_r[2]), .A1(wr_ptr_r[2]), .Z(n8));
Q_XNR2 U109 ( .A0(rd_ptr_r[1]), .A1(wr_ptr_r[1]), .Z(n7));
Q_XNR2 U110 ( .A0(rd_ptr_r[0]), .A1(wr_ptr_r[0]), .Z(n6));
Q_MX02 U111 ( .S(n10), .A0(rd_ptr_r[0]), .A1(wr_ptr_r[0]), .Z(n13));
Q_MX02 U112 ( .S(n10), .A0(rd_ptr_r[1]), .A1(wr_ptr_r[1]), .Z(n14));
Q_MX02 U113 ( .S(n10), .A0(rd_ptr_r[2]), .A1(wr_ptr_r[2]), .Z(n15));
Q_MX02 U114 ( .S(n10), .A0(wr_ptr_r[0]), .A1(rd_ptr_r[0]), .Z(n16));
Q_MX02 U115 ( .S(n10), .A0(wr_ptr_r[1]), .A1(rd_ptr_r[1]), .Z(n17));
Q_MX02 U116 ( .S(n10), .A0(wr_ptr_r[2]), .A1(rd_ptr_r[2]), .Z(n18));
Q_INV U117 ( .A(n16), .Z(n19));
Q_INV U118 ( .A(n17), .Z(n20));
Q_INV U119 ( .A(n18), .Z(n21));
Q_XNR2 U120 ( .A0(n13), .A1(n19), .Z(n5));
Q_OR02 U121 ( .A0(n13), .A1(n19), .Z(n22));
Q_AD02 U122 ( .CI(n22), .A0(n14), .A1(n15), .B0(n20), .B1(n21), .S0(n23), .S1(n24), .CO(n25));
Q_INV U123 ( .A(n25), .Z(n26));
Q_INV U124 ( .A(n5), .Z(n27));
Q_INV U125 ( .A(n23), .Z(n28));
Q_INV U126 ( .A(n24), .Z(n29));
Q_AD01HF U127 ( .A0(n27), .B0(n28), .S(n30), .CO(n31));
Q_AD01HF U128 ( .A0(n31), .B0(n29), .S(n32), .CO(n33));
Q_XNR2 U129 ( .A0(n33), .A1(n25), .Z(n34));
Q_MX02 U130 ( .S(n10), .A0(n23), .A1(n30), .Z(n4));
Q_MX02 U131 ( .S(n10), .A0(n24), .A1(n32), .Z(n3));
Q_MX02 U132 ( .S(n10), .A0(n26), .A1(n34), .Z(n2));
Q_FDP1 \rd_ptr_r_REG[0] ( .CK(clk), .R(rst_n), .D(rd_ptr_nxt[0]), .Q(rd_ptr_r[0]), .QN(n86));
Q_FDP1 \rd_ptr_r_REG[1] ( .CK(clk), .R(rst_n), .D(rd_ptr_nxt[1]), .Q(rd_ptr_r[1]), .QN( ));
Q_FDP1 \rd_ptr_r_REG[2] ( .CK(clk), .R(rst_n), .D(rd_ptr_nxt[2]), .Q(rd_ptr_r[2]), .QN( ));
Q_FDP1 \rd_ptr_r_REG[3] ( .CK(clk), .R(rst_n), .D(rd_ptr_nxt[3]), .Q(rd_ptr_r[3]), .QN( ));
Q_FDP1 \wr_ptr_r_REG[0] ( .CK(clk), .R(rst_n), .D(wr_ptr_nxt[0]), .Q(wr_ptr_r[0]), .QN(n40));
Q_FDP1 \wr_ptr_r_REG[1] ( .CK(clk), .R(rst_n), .D(wr_ptr_nxt[1]), .Q(wr_ptr_r[1]), .QN(n48));
Q_FDP1 \wr_ptr_r_REG[2] ( .CK(clk), .R(rst_n), .D(wr_ptr_nxt[2]), .Q(wr_ptr_r[2]), .QN( ));
Q_FDP1 \wr_ptr_r_REG[3] ( .CK(clk), .R(rst_n), .D(wr_ptr_nxt[3]), .Q(wr_ptr_r[3]), .QN( ));
Q_MX02 U141 ( .S(n56), .A0(\mem_r[7][0] ), .A1(din[0]), .Z(\mem_nxt[7][0] ));
Q_MX02 U142 ( .S(n56), .A0(\mem_r[7][1] ), .A1(din[1]), .Z(\mem_nxt[7][1] ));
Q_MX02 U143 ( .S(n56), .A0(\mem_r[7][2] ), .A1(din[2]), .Z(\mem_nxt[7][2] ));
Q_MX02 U144 ( .S(n56), .A0(\mem_r[7][3] ), .A1(din[3]), .Z(\mem_nxt[7][3] ));
Q_MX02 U145 ( .S(n56), .A0(\mem_r[7][4] ), .A1(din[4]), .Z(\mem_nxt[7][4] ));
Q_MX02 U146 ( .S(n56), .A0(\mem_r[7][5] ), .A1(din[5]), .Z(\mem_nxt[7][5] ));
Q_MX02 U147 ( .S(n56), .A0(\mem_r[7][6] ), .A1(din[6]), .Z(\mem_nxt[7][6] ));
Q_MX02 U148 ( .S(n56), .A0(\mem_r[7][7] ), .A1(din[7]), .Z(\mem_nxt[7][7] ));
Q_MX02 U149 ( .S(n56), .A0(\mem_r[7][8] ), .A1(din[8]), .Z(\mem_nxt[7][8] ));
Q_MX02 U150 ( .S(n56), .A0(\mem_r[7][9] ), .A1(din[9]), .Z(\mem_nxt[7][9] ));
Q_MX02 U151 ( .S(n56), .A0(\mem_r[7][10] ), .A1(din[10]), .Z(\mem_nxt[7][10] ));
Q_MX02 U152 ( .S(n56), .A0(\mem_r[7][11] ), .A1(din[11]), .Z(\mem_nxt[7][11] ));
Q_MX02 U153 ( .S(n56), .A0(\mem_r[7][12] ), .A1(din[12]), .Z(\mem_nxt[7][12] ));
Q_MX02 U154 ( .S(n56), .A0(\mem_r[7][13] ), .A1(din[13]), .Z(\mem_nxt[7][13] ));
Q_MX02 U155 ( .S(n56), .A0(\mem_r[7][14] ), .A1(din[14]), .Z(\mem_nxt[7][14] ));
Q_MX02 U156 ( .S(n56), .A0(\mem_r[7][15] ), .A1(din[15]), .Z(\mem_nxt[7][15] ));
Q_MX02 U157 ( .S(n56), .A0(\mem_r[7][16] ), .A1(din[16]), .Z(\mem_nxt[7][16] ));
Q_MX02 U158 ( .S(n56), .A0(\mem_r[7][17] ), .A1(din[17]), .Z(\mem_nxt[7][17] ));
Q_MX02 U159 ( .S(n56), .A0(\mem_r[7][18] ), .A1(din[18]), .Z(\mem_nxt[7][18] ));
Q_MX02 U160 ( .S(n56), .A0(\mem_r[7][19] ), .A1(din[19]), .Z(\mem_nxt[7][19] ));
Q_MX02 U161 ( .S(n56), .A0(\mem_r[7][20] ), .A1(din[20]), .Z(\mem_nxt[7][20] ));
Q_MX02 U162 ( .S(n56), .A0(\mem_r[7][21] ), .A1(din[21]), .Z(\mem_nxt[7][21] ));
Q_MX02 U163 ( .S(n56), .A0(\mem_r[7][22] ), .A1(din[22]), .Z(\mem_nxt[7][22] ));
Q_MX02 U164 ( .S(n56), .A0(\mem_r[7][23] ), .A1(din[23]), .Z(\mem_nxt[7][23] ));
Q_MX02 U165 ( .S(n56), .A0(\mem_r[7][24] ), .A1(din[24]), .Z(\mem_nxt[7][24] ));
Q_MX02 U166 ( .S(n56), .A0(\mem_r[7][25] ), .A1(din[25]), .Z(\mem_nxt[7][25] ));
Q_MX02 U167 ( .S(n56), .A0(\mem_r[7][26] ), .A1(din[26]), .Z(\mem_nxt[7][26] ));
Q_MX02 U168 ( .S(n56), .A0(\mem_r[7][27] ), .A1(din[27]), .Z(\mem_nxt[7][27] ));
Q_MX02 U169 ( .S(n56), .A0(\mem_r[7][28] ), .A1(din[28]), .Z(\mem_nxt[7][28] ));
Q_MX02 U170 ( .S(n56), .A0(\mem_r[7][29] ), .A1(din[29]), .Z(\mem_nxt[7][29] ));
Q_MX02 U171 ( .S(n56), .A0(\mem_r[7][30] ), .A1(din[30]), .Z(\mem_nxt[7][30] ));
Q_MX02 U172 ( .S(n56), .A0(\mem_r[7][31] ), .A1(din[31]), .Z(\mem_nxt[7][31] ));
Q_MX02 U173 ( .S(n56), .A0(\mem_r[7][32] ), .A1(din[32]), .Z(\mem_nxt[7][32] ));
Q_MX02 U174 ( .S(n56), .A0(\mem_r[7][33] ), .A1(din[33]), .Z(\mem_nxt[7][33] ));
Q_MX02 U175 ( .S(n56), .A0(\mem_r[7][34] ), .A1(din[34]), .Z(\mem_nxt[7][34] ));
Q_MX02 U176 ( .S(n56), .A0(\mem_r[7][35] ), .A1(din[35]), .Z(\mem_nxt[7][35] ));
Q_MX02 U177 ( .S(n56), .A0(\mem_r[7][36] ), .A1(din[36]), .Z(\mem_nxt[7][36] ));
Q_MX02 U178 ( .S(n56), .A0(\mem_r[7][37] ), .A1(din[37]), .Z(\mem_nxt[7][37] ));
Q_MX02 U179 ( .S(n56), .A0(\mem_r[7][38] ), .A1(din[38]), .Z(\mem_nxt[7][38] ));
Q_MX02 U180 ( .S(n56), .A0(\mem_r[7][39] ), .A1(din[39]), .Z(\mem_nxt[7][39] ));
Q_MX02 U181 ( .S(n56), .A0(\mem_r[7][40] ), .A1(din[40]), .Z(\mem_nxt[7][40] ));
Q_MX02 U182 ( .S(n56), .A0(\mem_r[7][41] ), .A1(din[41]), .Z(\mem_nxt[7][41] ));
Q_MX02 U183 ( .S(n56), .A0(\mem_r[7][42] ), .A1(din[42]), .Z(\mem_nxt[7][42] ));
Q_MX02 U184 ( .S(n56), .A0(\mem_r[7][43] ), .A1(din[43]), .Z(\mem_nxt[7][43] ));
Q_MX02 U185 ( .S(n56), .A0(\mem_r[7][44] ), .A1(din[44]), .Z(\mem_nxt[7][44] ));
Q_MX02 U186 ( .S(n56), .A0(\mem_r[7][45] ), .A1(din[45]), .Z(\mem_nxt[7][45] ));
Q_MX02 U187 ( .S(n56), .A0(\mem_r[7][46] ), .A1(din[46]), .Z(\mem_nxt[7][46] ));
Q_MX02 U188 ( .S(n56), .A0(\mem_r[7][47] ), .A1(din[47]), .Z(\mem_nxt[7][47] ));
Q_MX02 U189 ( .S(n56), .A0(\mem_r[7][48] ), .A1(din[48]), .Z(\mem_nxt[7][48] ));
Q_MX02 U190 ( .S(n56), .A0(\mem_r[7][49] ), .A1(din[49]), .Z(\mem_nxt[7][49] ));
Q_MX02 U191 ( .S(n56), .A0(\mem_r[7][50] ), .A1(din[50]), .Z(\mem_nxt[7][50] ));
Q_MX02 U192 ( .S(n56), .A0(\mem_r[7][51] ), .A1(din[51]), .Z(\mem_nxt[7][51] ));
Q_MX02 U193 ( .S(n56), .A0(\mem_r[7][52] ), .A1(din[52]), .Z(\mem_nxt[7][52] ));
Q_MX02 U194 ( .S(n56), .A0(\mem_r[7][53] ), .A1(din[53]), .Z(\mem_nxt[7][53] ));
Q_MX02 U195 ( .S(n56), .A0(\mem_r[7][54] ), .A1(din[54]), .Z(\mem_nxt[7][54] ));
Q_MX02 U196 ( .S(n56), .A0(\mem_r[7][55] ), .A1(din[55]), .Z(\mem_nxt[7][55] ));
Q_MX02 U197 ( .S(n56), .A0(\mem_r[7][56] ), .A1(din[56]), .Z(\mem_nxt[7][56] ));
Q_MX02 U198 ( .S(n56), .A0(\mem_r[7][57] ), .A1(din[57]), .Z(\mem_nxt[7][57] ));
Q_MX02 U199 ( .S(n56), .A0(\mem_r[7][58] ), .A1(din[58]), .Z(\mem_nxt[7][58] ));
Q_MX02 U200 ( .S(n56), .A0(\mem_r[7][59] ), .A1(din[59]), .Z(\mem_nxt[7][59] ));
Q_MX02 U201 ( .S(n56), .A0(\mem_r[7][60] ), .A1(din[60]), .Z(\mem_nxt[7][60] ));
Q_MX02 U202 ( .S(n56), .A0(\mem_r[7][61] ), .A1(din[61]), .Z(\mem_nxt[7][61] ));
Q_MX02 U203 ( .S(n56), .A0(\mem_r[7][62] ), .A1(din[62]), .Z(\mem_nxt[7][62] ));
Q_MX02 U204 ( .S(n56), .A0(\mem_r[7][63] ), .A1(din[63]), .Z(\mem_nxt[7][63] ));
Q_MX02 U205 ( .S(n56), .A0(\mem_r[7][64] ), .A1(din[64]), .Z(\mem_nxt[7][64] ));
Q_MX02 U206 ( .S(n56), .A0(\mem_r[7][65] ), .A1(din[65]), .Z(\mem_nxt[7][65] ));
Q_MX02 U207 ( .S(n56), .A0(\mem_r[7][66] ), .A1(din[66]), .Z(\mem_nxt[7][66] ));
Q_MX02 U208 ( .S(n56), .A0(\mem_r[7][67] ), .A1(din[67]), .Z(\mem_nxt[7][67] ));
Q_MX02 U209 ( .S(n56), .A0(\mem_r[7][68] ), .A1(din[68]), .Z(\mem_nxt[7][68] ));
Q_MX02 U210 ( .S(n56), .A0(\mem_r[7][69] ), .A1(din[69]), .Z(\mem_nxt[7][69] ));
Q_MX02 U211 ( .S(n56), .A0(\mem_r[7][70] ), .A1(din[70]), .Z(\mem_nxt[7][70] ));
Q_MX02 U212 ( .S(n56), .A0(\mem_r[7][71] ), .A1(din[71]), .Z(\mem_nxt[7][71] ));
Q_MX02 U213 ( .S(n56), .A0(\mem_r[7][72] ), .A1(din[72]), .Z(\mem_nxt[7][72] ));
Q_MX02 U214 ( .S(n56), .A0(\mem_r[7][73] ), .A1(din[73]), .Z(\mem_nxt[7][73] ));
Q_MX02 U215 ( .S(n56), .A0(\mem_r[7][74] ), .A1(din[74]), .Z(\mem_nxt[7][74] ));
Q_MX02 U216 ( .S(n56), .A0(\mem_r[7][75] ), .A1(din[75]), .Z(\mem_nxt[7][75] ));
Q_MX02 U217 ( .S(n56), .A0(\mem_r[7][76] ), .A1(din[76]), .Z(\mem_nxt[7][76] ));
Q_MX02 U218 ( .S(n56), .A0(\mem_r[7][77] ), .A1(din[77]), .Z(\mem_nxt[7][77] ));
Q_MX02 U219 ( .S(n56), .A0(\mem_r[7][78] ), .A1(din[78]), .Z(\mem_nxt[7][78] ));
Q_MX02 U220 ( .S(n56), .A0(\mem_r[7][79] ), .A1(din[79]), .Z(\mem_nxt[7][79] ));
Q_MX02 U221 ( .S(n56), .A0(\mem_r[7][80] ), .A1(din[80]), .Z(\mem_nxt[7][80] ));
Q_MX02 U222 ( .S(n56), .A0(\mem_r[7][81] ), .A1(din[81]), .Z(\mem_nxt[7][81] ));
Q_MX02 U223 ( .S(n56), .A0(\mem_r[7][82] ), .A1(din[82]), .Z(\mem_nxt[7][82] ));
Q_MX02 U224 ( .S(n56), .A0(\mem_r[7][83] ), .A1(din[83]), .Z(\mem_nxt[7][83] ));
Q_MX02 U225 ( .S(n56), .A0(\mem_r[7][84] ), .A1(din[84]), .Z(\mem_nxt[7][84] ));
Q_MX02 U226 ( .S(n56), .A0(\mem_r[7][85] ), .A1(din[85]), .Z(\mem_nxt[7][85] ));
Q_MX02 U227 ( .S(n56), .A0(\mem_r[7][86] ), .A1(din[86]), .Z(\mem_nxt[7][86] ));
Q_MX02 U228 ( .S(n56), .A0(\mem_r[7][87] ), .A1(din[87]), .Z(\mem_nxt[7][87] ));
Q_MX02 U229 ( .S(n56), .A0(\mem_r[7][88] ), .A1(din[88]), .Z(\mem_nxt[7][88] ));
Q_MX02 U230 ( .S(n56), .A0(\mem_r[7][89] ), .A1(din[89]), .Z(\mem_nxt[7][89] ));
Q_MX02 U231 ( .S(n56), .A0(\mem_r[7][90] ), .A1(din[90]), .Z(\mem_nxt[7][90] ));
Q_MX02 U232 ( .S(n56), .A0(\mem_r[7][91] ), .A1(din[91]), .Z(\mem_nxt[7][91] ));
Q_MX02 U233 ( .S(n56), .A0(\mem_r[7][92] ), .A1(din[92]), .Z(\mem_nxt[7][92] ));
Q_MX02 U234 ( .S(n56), .A0(\mem_r[7][93] ), .A1(din[93]), .Z(\mem_nxt[7][93] ));
Q_MX02 U235 ( .S(n56), .A0(\mem_r[7][94] ), .A1(din[94]), .Z(\mem_nxt[7][94] ));
Q_MX02 U236 ( .S(n56), .A0(\mem_r[7][95] ), .A1(din[95]), .Z(\mem_nxt[7][95] ));
Q_MX02 U237 ( .S(n36), .A0(\mem_r[6][0] ), .A1(din[0]), .Z(\mem_nxt[6][0] ));
Q_MX02 U238 ( .S(n36), .A0(\mem_r[6][1] ), .A1(din[1]), .Z(\mem_nxt[6][1] ));
Q_MX02 U239 ( .S(n36), .A0(\mem_r[6][2] ), .A1(din[2]), .Z(\mem_nxt[6][2] ));
Q_MX02 U240 ( .S(n36), .A0(\mem_r[6][3] ), .A1(din[3]), .Z(\mem_nxt[6][3] ));
Q_MX02 U241 ( .S(n36), .A0(\mem_r[6][4] ), .A1(din[4]), .Z(\mem_nxt[6][4] ));
Q_MX02 U242 ( .S(n36), .A0(\mem_r[6][5] ), .A1(din[5]), .Z(\mem_nxt[6][5] ));
Q_MX02 U243 ( .S(n36), .A0(\mem_r[6][6] ), .A1(din[6]), .Z(\mem_nxt[6][6] ));
Q_MX02 U244 ( .S(n36), .A0(\mem_r[6][7] ), .A1(din[7]), .Z(\mem_nxt[6][7] ));
Q_MX02 U245 ( .S(n36), .A0(\mem_r[6][8] ), .A1(din[8]), .Z(\mem_nxt[6][8] ));
Q_MX02 U246 ( .S(n36), .A0(\mem_r[6][9] ), .A1(din[9]), .Z(\mem_nxt[6][9] ));
Q_MX02 U247 ( .S(n36), .A0(\mem_r[6][10] ), .A1(din[10]), .Z(\mem_nxt[6][10] ));
Q_MX02 U248 ( .S(n36), .A0(\mem_r[6][11] ), .A1(din[11]), .Z(\mem_nxt[6][11] ));
Q_MX02 U249 ( .S(n36), .A0(\mem_r[6][12] ), .A1(din[12]), .Z(\mem_nxt[6][12] ));
Q_MX02 U250 ( .S(n36), .A0(\mem_r[6][13] ), .A1(din[13]), .Z(\mem_nxt[6][13] ));
Q_MX02 U251 ( .S(n36), .A0(\mem_r[6][14] ), .A1(din[14]), .Z(\mem_nxt[6][14] ));
Q_MX02 U252 ( .S(n36), .A0(\mem_r[6][15] ), .A1(din[15]), .Z(\mem_nxt[6][15] ));
Q_MX02 U253 ( .S(n36), .A0(\mem_r[6][16] ), .A1(din[16]), .Z(\mem_nxt[6][16] ));
Q_MX02 U254 ( .S(n36), .A0(\mem_r[6][17] ), .A1(din[17]), .Z(\mem_nxt[6][17] ));
Q_MX02 U255 ( .S(n36), .A0(\mem_r[6][18] ), .A1(din[18]), .Z(\mem_nxt[6][18] ));
Q_MX02 U256 ( .S(n36), .A0(\mem_r[6][19] ), .A1(din[19]), .Z(\mem_nxt[6][19] ));
Q_MX02 U257 ( .S(n36), .A0(\mem_r[6][20] ), .A1(din[20]), .Z(\mem_nxt[6][20] ));
Q_MX02 U258 ( .S(n36), .A0(\mem_r[6][21] ), .A1(din[21]), .Z(\mem_nxt[6][21] ));
Q_MX02 U259 ( .S(n36), .A0(\mem_r[6][22] ), .A1(din[22]), .Z(\mem_nxt[6][22] ));
Q_MX02 U260 ( .S(n36), .A0(\mem_r[6][23] ), .A1(din[23]), .Z(\mem_nxt[6][23] ));
Q_MX02 U261 ( .S(n36), .A0(\mem_r[6][24] ), .A1(din[24]), .Z(\mem_nxt[6][24] ));
Q_MX02 U262 ( .S(n36), .A0(\mem_r[6][25] ), .A1(din[25]), .Z(\mem_nxt[6][25] ));
Q_MX02 U263 ( .S(n36), .A0(\mem_r[6][26] ), .A1(din[26]), .Z(\mem_nxt[6][26] ));
Q_MX02 U264 ( .S(n36), .A0(\mem_r[6][27] ), .A1(din[27]), .Z(\mem_nxt[6][27] ));
Q_MX02 U265 ( .S(n36), .A0(\mem_r[6][28] ), .A1(din[28]), .Z(\mem_nxt[6][28] ));
Q_MX02 U266 ( .S(n36), .A0(\mem_r[6][29] ), .A1(din[29]), .Z(\mem_nxt[6][29] ));
Q_MX02 U267 ( .S(n36), .A0(\mem_r[6][30] ), .A1(din[30]), .Z(\mem_nxt[6][30] ));
Q_MX02 U268 ( .S(n36), .A0(\mem_r[6][31] ), .A1(din[31]), .Z(\mem_nxt[6][31] ));
Q_MX02 U269 ( .S(n36), .A0(\mem_r[6][32] ), .A1(din[32]), .Z(\mem_nxt[6][32] ));
Q_MX02 U270 ( .S(n36), .A0(\mem_r[6][33] ), .A1(din[33]), .Z(\mem_nxt[6][33] ));
Q_MX02 U271 ( .S(n36), .A0(\mem_r[6][34] ), .A1(din[34]), .Z(\mem_nxt[6][34] ));
Q_MX02 U272 ( .S(n36), .A0(\mem_r[6][35] ), .A1(din[35]), .Z(\mem_nxt[6][35] ));
Q_MX02 U273 ( .S(n36), .A0(\mem_r[6][36] ), .A1(din[36]), .Z(\mem_nxt[6][36] ));
Q_MX02 U274 ( .S(n36), .A0(\mem_r[6][37] ), .A1(din[37]), .Z(\mem_nxt[6][37] ));
Q_MX02 U275 ( .S(n36), .A0(\mem_r[6][38] ), .A1(din[38]), .Z(\mem_nxt[6][38] ));
Q_MX02 U276 ( .S(n36), .A0(\mem_r[6][39] ), .A1(din[39]), .Z(\mem_nxt[6][39] ));
Q_MX02 U277 ( .S(n36), .A0(\mem_r[6][40] ), .A1(din[40]), .Z(\mem_nxt[6][40] ));
Q_MX02 U278 ( .S(n36), .A0(\mem_r[6][41] ), .A1(din[41]), .Z(\mem_nxt[6][41] ));
Q_MX02 U279 ( .S(n36), .A0(\mem_r[6][42] ), .A1(din[42]), .Z(\mem_nxt[6][42] ));
Q_MX02 U280 ( .S(n36), .A0(\mem_r[6][43] ), .A1(din[43]), .Z(\mem_nxt[6][43] ));
Q_MX02 U281 ( .S(n36), .A0(\mem_r[6][44] ), .A1(din[44]), .Z(\mem_nxt[6][44] ));
Q_MX02 U282 ( .S(n36), .A0(\mem_r[6][45] ), .A1(din[45]), .Z(\mem_nxt[6][45] ));
Q_MX02 U283 ( .S(n36), .A0(\mem_r[6][46] ), .A1(din[46]), .Z(\mem_nxt[6][46] ));
Q_MX02 U284 ( .S(n36), .A0(\mem_r[6][47] ), .A1(din[47]), .Z(\mem_nxt[6][47] ));
Q_MX02 U285 ( .S(n36), .A0(\mem_r[6][48] ), .A1(din[48]), .Z(\mem_nxt[6][48] ));
Q_MX02 U286 ( .S(n36), .A0(\mem_r[6][49] ), .A1(din[49]), .Z(\mem_nxt[6][49] ));
Q_MX02 U287 ( .S(n36), .A0(\mem_r[6][50] ), .A1(din[50]), .Z(\mem_nxt[6][50] ));
Q_MX02 U288 ( .S(n36), .A0(\mem_r[6][51] ), .A1(din[51]), .Z(\mem_nxt[6][51] ));
Q_MX02 U289 ( .S(n36), .A0(\mem_r[6][52] ), .A1(din[52]), .Z(\mem_nxt[6][52] ));
Q_MX02 U290 ( .S(n36), .A0(\mem_r[6][53] ), .A1(din[53]), .Z(\mem_nxt[6][53] ));
Q_MX02 U291 ( .S(n36), .A0(\mem_r[6][54] ), .A1(din[54]), .Z(\mem_nxt[6][54] ));
Q_MX02 U292 ( .S(n36), .A0(\mem_r[6][55] ), .A1(din[55]), .Z(\mem_nxt[6][55] ));
Q_MX02 U293 ( .S(n36), .A0(\mem_r[6][56] ), .A1(din[56]), .Z(\mem_nxt[6][56] ));
Q_MX02 U294 ( .S(n36), .A0(\mem_r[6][57] ), .A1(din[57]), .Z(\mem_nxt[6][57] ));
Q_MX02 U295 ( .S(n36), .A0(\mem_r[6][58] ), .A1(din[58]), .Z(\mem_nxt[6][58] ));
Q_MX02 U296 ( .S(n36), .A0(\mem_r[6][59] ), .A1(din[59]), .Z(\mem_nxt[6][59] ));
Q_MX02 U297 ( .S(n36), .A0(\mem_r[6][60] ), .A1(din[60]), .Z(\mem_nxt[6][60] ));
Q_MX02 U298 ( .S(n36), .A0(\mem_r[6][61] ), .A1(din[61]), .Z(\mem_nxt[6][61] ));
Q_MX02 U299 ( .S(n36), .A0(\mem_r[6][62] ), .A1(din[62]), .Z(\mem_nxt[6][62] ));
Q_MX02 U300 ( .S(n36), .A0(\mem_r[6][63] ), .A1(din[63]), .Z(\mem_nxt[6][63] ));
Q_MX02 U301 ( .S(n36), .A0(\mem_r[6][64] ), .A1(din[64]), .Z(\mem_nxt[6][64] ));
Q_MX02 U302 ( .S(n36), .A0(\mem_r[6][65] ), .A1(din[65]), .Z(\mem_nxt[6][65] ));
Q_MX02 U303 ( .S(n36), .A0(\mem_r[6][66] ), .A1(din[66]), .Z(\mem_nxt[6][66] ));
Q_MX02 U304 ( .S(n36), .A0(\mem_r[6][67] ), .A1(din[67]), .Z(\mem_nxt[6][67] ));
Q_MX02 U305 ( .S(n36), .A0(\mem_r[6][68] ), .A1(din[68]), .Z(\mem_nxt[6][68] ));
Q_MX02 U306 ( .S(n36), .A0(\mem_r[6][69] ), .A1(din[69]), .Z(\mem_nxt[6][69] ));
Q_MX02 U307 ( .S(n36), .A0(\mem_r[6][70] ), .A1(din[70]), .Z(\mem_nxt[6][70] ));
Q_MX02 U308 ( .S(n36), .A0(\mem_r[6][71] ), .A1(din[71]), .Z(\mem_nxt[6][71] ));
Q_MX02 U309 ( .S(n36), .A0(\mem_r[6][72] ), .A1(din[72]), .Z(\mem_nxt[6][72] ));
Q_MX02 U310 ( .S(n36), .A0(\mem_r[6][73] ), .A1(din[73]), .Z(\mem_nxt[6][73] ));
Q_MX02 U311 ( .S(n36), .A0(\mem_r[6][74] ), .A1(din[74]), .Z(\mem_nxt[6][74] ));
Q_MX02 U312 ( .S(n36), .A0(\mem_r[6][75] ), .A1(din[75]), .Z(\mem_nxt[6][75] ));
Q_MX02 U313 ( .S(n36), .A0(\mem_r[6][76] ), .A1(din[76]), .Z(\mem_nxt[6][76] ));
Q_MX02 U314 ( .S(n36), .A0(\mem_r[6][77] ), .A1(din[77]), .Z(\mem_nxt[6][77] ));
Q_MX02 U315 ( .S(n36), .A0(\mem_r[6][78] ), .A1(din[78]), .Z(\mem_nxt[6][78] ));
Q_MX02 U316 ( .S(n36), .A0(\mem_r[6][79] ), .A1(din[79]), .Z(\mem_nxt[6][79] ));
Q_MX02 U317 ( .S(n36), .A0(\mem_r[6][80] ), .A1(din[80]), .Z(\mem_nxt[6][80] ));
Q_MX02 U318 ( .S(n36), .A0(\mem_r[6][81] ), .A1(din[81]), .Z(\mem_nxt[6][81] ));
Q_MX02 U319 ( .S(n36), .A0(\mem_r[6][82] ), .A1(din[82]), .Z(\mem_nxt[6][82] ));
Q_MX02 U320 ( .S(n36), .A0(\mem_r[6][83] ), .A1(din[83]), .Z(\mem_nxt[6][83] ));
Q_MX02 U321 ( .S(n36), .A0(\mem_r[6][84] ), .A1(din[84]), .Z(\mem_nxt[6][84] ));
Q_MX02 U322 ( .S(n36), .A0(\mem_r[6][85] ), .A1(din[85]), .Z(\mem_nxt[6][85] ));
Q_MX02 U323 ( .S(n36), .A0(\mem_r[6][86] ), .A1(din[86]), .Z(\mem_nxt[6][86] ));
Q_MX02 U324 ( .S(n36), .A0(\mem_r[6][87] ), .A1(din[87]), .Z(\mem_nxt[6][87] ));
Q_MX02 U325 ( .S(n36), .A0(\mem_r[6][88] ), .A1(din[88]), .Z(\mem_nxt[6][88] ));
Q_MX02 U326 ( .S(n36), .A0(\mem_r[6][89] ), .A1(din[89]), .Z(\mem_nxt[6][89] ));
Q_MX02 U327 ( .S(n36), .A0(\mem_r[6][90] ), .A1(din[90]), .Z(\mem_nxt[6][90] ));
Q_MX02 U328 ( .S(n36), .A0(\mem_r[6][91] ), .A1(din[91]), .Z(\mem_nxt[6][91] ));
Q_MX02 U329 ( .S(n36), .A0(\mem_r[6][92] ), .A1(din[92]), .Z(\mem_nxt[6][92] ));
Q_MX02 U330 ( .S(n36), .A0(\mem_r[6][93] ), .A1(din[93]), .Z(\mem_nxt[6][93] ));
Q_MX02 U331 ( .S(n36), .A0(\mem_r[6][94] ), .A1(din[94]), .Z(\mem_nxt[6][94] ));
Q_MX02 U332 ( .S(n36), .A0(\mem_r[6][95] ), .A1(din[95]), .Z(\mem_nxt[6][95] ));
Q_MX02 U333 ( .S(n39), .A0(\mem_r[5][0] ), .A1(din[0]), .Z(\mem_nxt[5][0] ));
Q_MX02 U334 ( .S(n39), .A0(\mem_r[5][1] ), .A1(din[1]), .Z(\mem_nxt[5][1] ));
Q_MX02 U335 ( .S(n39), .A0(\mem_r[5][2] ), .A1(din[2]), .Z(\mem_nxt[5][2] ));
Q_MX02 U336 ( .S(n39), .A0(\mem_r[5][3] ), .A1(din[3]), .Z(\mem_nxt[5][3] ));
Q_MX02 U337 ( .S(n39), .A0(\mem_r[5][4] ), .A1(din[4]), .Z(\mem_nxt[5][4] ));
Q_MX02 U338 ( .S(n39), .A0(\mem_r[5][5] ), .A1(din[5]), .Z(\mem_nxt[5][5] ));
Q_MX02 U339 ( .S(n39), .A0(\mem_r[5][6] ), .A1(din[6]), .Z(\mem_nxt[5][6] ));
Q_MX02 U340 ( .S(n39), .A0(\mem_r[5][7] ), .A1(din[7]), .Z(\mem_nxt[5][7] ));
Q_MX02 U341 ( .S(n39), .A0(\mem_r[5][8] ), .A1(din[8]), .Z(\mem_nxt[5][8] ));
Q_MX02 U342 ( .S(n39), .A0(\mem_r[5][9] ), .A1(din[9]), .Z(\mem_nxt[5][9] ));
Q_MX02 U343 ( .S(n39), .A0(\mem_r[5][10] ), .A1(din[10]), .Z(\mem_nxt[5][10] ));
Q_MX02 U344 ( .S(n39), .A0(\mem_r[5][11] ), .A1(din[11]), .Z(\mem_nxt[5][11] ));
Q_MX02 U345 ( .S(n39), .A0(\mem_r[5][12] ), .A1(din[12]), .Z(\mem_nxt[5][12] ));
Q_MX02 U346 ( .S(n39), .A0(\mem_r[5][13] ), .A1(din[13]), .Z(\mem_nxt[5][13] ));
Q_MX02 U347 ( .S(n39), .A0(\mem_r[5][14] ), .A1(din[14]), .Z(\mem_nxt[5][14] ));
Q_MX02 U348 ( .S(n39), .A0(\mem_r[5][15] ), .A1(din[15]), .Z(\mem_nxt[5][15] ));
Q_MX02 U349 ( .S(n39), .A0(\mem_r[5][16] ), .A1(din[16]), .Z(\mem_nxt[5][16] ));
Q_MX02 U350 ( .S(n39), .A0(\mem_r[5][17] ), .A1(din[17]), .Z(\mem_nxt[5][17] ));
Q_MX02 U351 ( .S(n39), .A0(\mem_r[5][18] ), .A1(din[18]), .Z(\mem_nxt[5][18] ));
Q_MX02 U352 ( .S(n39), .A0(\mem_r[5][19] ), .A1(din[19]), .Z(\mem_nxt[5][19] ));
Q_MX02 U353 ( .S(n39), .A0(\mem_r[5][20] ), .A1(din[20]), .Z(\mem_nxt[5][20] ));
Q_MX02 U354 ( .S(n39), .A0(\mem_r[5][21] ), .A1(din[21]), .Z(\mem_nxt[5][21] ));
Q_MX02 U355 ( .S(n39), .A0(\mem_r[5][22] ), .A1(din[22]), .Z(\mem_nxt[5][22] ));
Q_MX02 U356 ( .S(n39), .A0(\mem_r[5][23] ), .A1(din[23]), .Z(\mem_nxt[5][23] ));
Q_MX02 U357 ( .S(n39), .A0(\mem_r[5][24] ), .A1(din[24]), .Z(\mem_nxt[5][24] ));
Q_MX02 U358 ( .S(n39), .A0(\mem_r[5][25] ), .A1(din[25]), .Z(\mem_nxt[5][25] ));
Q_MX02 U359 ( .S(n39), .A0(\mem_r[5][26] ), .A1(din[26]), .Z(\mem_nxt[5][26] ));
Q_MX02 U360 ( .S(n39), .A0(\mem_r[5][27] ), .A1(din[27]), .Z(\mem_nxt[5][27] ));
Q_MX02 U361 ( .S(n39), .A0(\mem_r[5][28] ), .A1(din[28]), .Z(\mem_nxt[5][28] ));
Q_MX02 U362 ( .S(n39), .A0(\mem_r[5][29] ), .A1(din[29]), .Z(\mem_nxt[5][29] ));
Q_MX02 U363 ( .S(n39), .A0(\mem_r[5][30] ), .A1(din[30]), .Z(\mem_nxt[5][30] ));
Q_MX02 U364 ( .S(n39), .A0(\mem_r[5][31] ), .A1(din[31]), .Z(\mem_nxt[5][31] ));
Q_MX02 U365 ( .S(n39), .A0(\mem_r[5][32] ), .A1(din[32]), .Z(\mem_nxt[5][32] ));
Q_MX02 U366 ( .S(n39), .A0(\mem_r[5][33] ), .A1(din[33]), .Z(\mem_nxt[5][33] ));
Q_MX02 U367 ( .S(n39), .A0(\mem_r[5][34] ), .A1(din[34]), .Z(\mem_nxt[5][34] ));
Q_MX02 U368 ( .S(n39), .A0(\mem_r[5][35] ), .A1(din[35]), .Z(\mem_nxt[5][35] ));
Q_MX02 U369 ( .S(n39), .A0(\mem_r[5][36] ), .A1(din[36]), .Z(\mem_nxt[5][36] ));
Q_MX02 U370 ( .S(n39), .A0(\mem_r[5][37] ), .A1(din[37]), .Z(\mem_nxt[5][37] ));
Q_MX02 U371 ( .S(n39), .A0(\mem_r[5][38] ), .A1(din[38]), .Z(\mem_nxt[5][38] ));
Q_MX02 U372 ( .S(n39), .A0(\mem_r[5][39] ), .A1(din[39]), .Z(\mem_nxt[5][39] ));
Q_MX02 U373 ( .S(n39), .A0(\mem_r[5][40] ), .A1(din[40]), .Z(\mem_nxt[5][40] ));
Q_MX02 U374 ( .S(n39), .A0(\mem_r[5][41] ), .A1(din[41]), .Z(\mem_nxt[5][41] ));
Q_MX02 U375 ( .S(n39), .A0(\mem_r[5][42] ), .A1(din[42]), .Z(\mem_nxt[5][42] ));
Q_MX02 U376 ( .S(n39), .A0(\mem_r[5][43] ), .A1(din[43]), .Z(\mem_nxt[5][43] ));
Q_MX02 U377 ( .S(n39), .A0(\mem_r[5][44] ), .A1(din[44]), .Z(\mem_nxt[5][44] ));
Q_MX02 U378 ( .S(n39), .A0(\mem_r[5][45] ), .A1(din[45]), .Z(\mem_nxt[5][45] ));
Q_MX02 U379 ( .S(n39), .A0(\mem_r[5][46] ), .A1(din[46]), .Z(\mem_nxt[5][46] ));
Q_MX02 U380 ( .S(n39), .A0(\mem_r[5][47] ), .A1(din[47]), .Z(\mem_nxt[5][47] ));
Q_MX02 U381 ( .S(n39), .A0(\mem_r[5][48] ), .A1(din[48]), .Z(\mem_nxt[5][48] ));
Q_MX02 U382 ( .S(n39), .A0(\mem_r[5][49] ), .A1(din[49]), .Z(\mem_nxt[5][49] ));
Q_MX02 U383 ( .S(n39), .A0(\mem_r[5][50] ), .A1(din[50]), .Z(\mem_nxt[5][50] ));
Q_MX02 U384 ( .S(n39), .A0(\mem_r[5][51] ), .A1(din[51]), .Z(\mem_nxt[5][51] ));
Q_MX02 U385 ( .S(n39), .A0(\mem_r[5][52] ), .A1(din[52]), .Z(\mem_nxt[5][52] ));
Q_MX02 U386 ( .S(n39), .A0(\mem_r[5][53] ), .A1(din[53]), .Z(\mem_nxt[5][53] ));
Q_MX02 U387 ( .S(n39), .A0(\mem_r[5][54] ), .A1(din[54]), .Z(\mem_nxt[5][54] ));
Q_MX02 U388 ( .S(n39), .A0(\mem_r[5][55] ), .A1(din[55]), .Z(\mem_nxt[5][55] ));
Q_MX02 U389 ( .S(n39), .A0(\mem_r[5][56] ), .A1(din[56]), .Z(\mem_nxt[5][56] ));
Q_MX02 U390 ( .S(n39), .A0(\mem_r[5][57] ), .A1(din[57]), .Z(\mem_nxt[5][57] ));
Q_MX02 U391 ( .S(n39), .A0(\mem_r[5][58] ), .A1(din[58]), .Z(\mem_nxt[5][58] ));
Q_MX02 U392 ( .S(n39), .A0(\mem_r[5][59] ), .A1(din[59]), .Z(\mem_nxt[5][59] ));
Q_MX02 U393 ( .S(n39), .A0(\mem_r[5][60] ), .A1(din[60]), .Z(\mem_nxt[5][60] ));
Q_MX02 U394 ( .S(n39), .A0(\mem_r[5][61] ), .A1(din[61]), .Z(\mem_nxt[5][61] ));
Q_MX02 U395 ( .S(n39), .A0(\mem_r[5][62] ), .A1(din[62]), .Z(\mem_nxt[5][62] ));
Q_MX02 U396 ( .S(n39), .A0(\mem_r[5][63] ), .A1(din[63]), .Z(\mem_nxt[5][63] ));
Q_MX02 U397 ( .S(n39), .A0(\mem_r[5][64] ), .A1(din[64]), .Z(\mem_nxt[5][64] ));
Q_MX02 U398 ( .S(n39), .A0(\mem_r[5][65] ), .A1(din[65]), .Z(\mem_nxt[5][65] ));
Q_MX02 U399 ( .S(n39), .A0(\mem_r[5][66] ), .A1(din[66]), .Z(\mem_nxt[5][66] ));
Q_MX02 U400 ( .S(n39), .A0(\mem_r[5][67] ), .A1(din[67]), .Z(\mem_nxt[5][67] ));
Q_MX02 U401 ( .S(n39), .A0(\mem_r[5][68] ), .A1(din[68]), .Z(\mem_nxt[5][68] ));
Q_MX02 U402 ( .S(n39), .A0(\mem_r[5][69] ), .A1(din[69]), .Z(\mem_nxt[5][69] ));
Q_MX02 U403 ( .S(n39), .A0(\mem_r[5][70] ), .A1(din[70]), .Z(\mem_nxt[5][70] ));
Q_MX02 U404 ( .S(n39), .A0(\mem_r[5][71] ), .A1(din[71]), .Z(\mem_nxt[5][71] ));
Q_MX02 U405 ( .S(n39), .A0(\mem_r[5][72] ), .A1(din[72]), .Z(\mem_nxt[5][72] ));
Q_MX02 U406 ( .S(n39), .A0(\mem_r[5][73] ), .A1(din[73]), .Z(\mem_nxt[5][73] ));
Q_MX02 U407 ( .S(n39), .A0(\mem_r[5][74] ), .A1(din[74]), .Z(\mem_nxt[5][74] ));
Q_MX02 U408 ( .S(n39), .A0(\mem_r[5][75] ), .A1(din[75]), .Z(\mem_nxt[5][75] ));
Q_MX02 U409 ( .S(n39), .A0(\mem_r[5][76] ), .A1(din[76]), .Z(\mem_nxt[5][76] ));
Q_MX02 U410 ( .S(n39), .A0(\mem_r[5][77] ), .A1(din[77]), .Z(\mem_nxt[5][77] ));
Q_MX02 U411 ( .S(n39), .A0(\mem_r[5][78] ), .A1(din[78]), .Z(\mem_nxt[5][78] ));
Q_MX02 U412 ( .S(n39), .A0(\mem_r[5][79] ), .A1(din[79]), .Z(\mem_nxt[5][79] ));
Q_MX02 U413 ( .S(n39), .A0(\mem_r[5][80] ), .A1(din[80]), .Z(\mem_nxt[5][80] ));
Q_MX02 U414 ( .S(n39), .A0(\mem_r[5][81] ), .A1(din[81]), .Z(\mem_nxt[5][81] ));
Q_MX02 U415 ( .S(n39), .A0(\mem_r[5][82] ), .A1(din[82]), .Z(\mem_nxt[5][82] ));
Q_MX02 U416 ( .S(n39), .A0(\mem_r[5][83] ), .A1(din[83]), .Z(\mem_nxt[5][83] ));
Q_MX02 U417 ( .S(n39), .A0(\mem_r[5][84] ), .A1(din[84]), .Z(\mem_nxt[5][84] ));
Q_MX02 U418 ( .S(n39), .A0(\mem_r[5][85] ), .A1(din[85]), .Z(\mem_nxt[5][85] ));
Q_MX02 U419 ( .S(n39), .A0(\mem_r[5][86] ), .A1(din[86]), .Z(\mem_nxt[5][86] ));
Q_MX02 U420 ( .S(n39), .A0(\mem_r[5][87] ), .A1(din[87]), .Z(\mem_nxt[5][87] ));
Q_MX02 U421 ( .S(n39), .A0(\mem_r[5][88] ), .A1(din[88]), .Z(\mem_nxt[5][88] ));
Q_MX02 U422 ( .S(n39), .A0(\mem_r[5][89] ), .A1(din[89]), .Z(\mem_nxt[5][89] ));
Q_MX02 U423 ( .S(n39), .A0(\mem_r[5][90] ), .A1(din[90]), .Z(\mem_nxt[5][90] ));
Q_MX02 U424 ( .S(n39), .A0(\mem_r[5][91] ), .A1(din[91]), .Z(\mem_nxt[5][91] ));
Q_MX02 U425 ( .S(n39), .A0(\mem_r[5][92] ), .A1(din[92]), .Z(\mem_nxt[5][92] ));
Q_MX02 U426 ( .S(n39), .A0(\mem_r[5][93] ), .A1(din[93]), .Z(\mem_nxt[5][93] ));
Q_MX02 U427 ( .S(n39), .A0(\mem_r[5][94] ), .A1(din[94]), .Z(\mem_nxt[5][94] ));
Q_MX02 U428 ( .S(n39), .A0(\mem_r[5][95] ), .A1(din[95]), .Z(\mem_nxt[5][95] ));
Q_MX02 U429 ( .S(n42), .A0(\mem_r[4][0] ), .A1(din[0]), .Z(\mem_nxt[4][0] ));
Q_MX02 U430 ( .S(n42), .A0(\mem_r[4][1] ), .A1(din[1]), .Z(\mem_nxt[4][1] ));
Q_MX02 U431 ( .S(n42), .A0(\mem_r[4][2] ), .A1(din[2]), .Z(\mem_nxt[4][2] ));
Q_MX02 U432 ( .S(n42), .A0(\mem_r[4][3] ), .A1(din[3]), .Z(\mem_nxt[4][3] ));
Q_MX02 U433 ( .S(n42), .A0(\mem_r[4][4] ), .A1(din[4]), .Z(\mem_nxt[4][4] ));
Q_MX02 U434 ( .S(n42), .A0(\mem_r[4][5] ), .A1(din[5]), .Z(\mem_nxt[4][5] ));
Q_MX02 U435 ( .S(n42), .A0(\mem_r[4][6] ), .A1(din[6]), .Z(\mem_nxt[4][6] ));
Q_MX02 U436 ( .S(n42), .A0(\mem_r[4][7] ), .A1(din[7]), .Z(\mem_nxt[4][7] ));
Q_MX02 U437 ( .S(n42), .A0(\mem_r[4][8] ), .A1(din[8]), .Z(\mem_nxt[4][8] ));
Q_MX02 U438 ( .S(n42), .A0(\mem_r[4][9] ), .A1(din[9]), .Z(\mem_nxt[4][9] ));
Q_MX02 U439 ( .S(n42), .A0(\mem_r[4][10] ), .A1(din[10]), .Z(\mem_nxt[4][10] ));
Q_MX02 U440 ( .S(n42), .A0(\mem_r[4][11] ), .A1(din[11]), .Z(\mem_nxt[4][11] ));
Q_MX02 U441 ( .S(n42), .A0(\mem_r[4][12] ), .A1(din[12]), .Z(\mem_nxt[4][12] ));
Q_MX02 U442 ( .S(n42), .A0(\mem_r[4][13] ), .A1(din[13]), .Z(\mem_nxt[4][13] ));
Q_MX02 U443 ( .S(n42), .A0(\mem_r[4][14] ), .A1(din[14]), .Z(\mem_nxt[4][14] ));
Q_MX02 U444 ( .S(n42), .A0(\mem_r[4][15] ), .A1(din[15]), .Z(\mem_nxt[4][15] ));
Q_MX02 U445 ( .S(n42), .A0(\mem_r[4][16] ), .A1(din[16]), .Z(\mem_nxt[4][16] ));
Q_MX02 U446 ( .S(n42), .A0(\mem_r[4][17] ), .A1(din[17]), .Z(\mem_nxt[4][17] ));
Q_MX02 U447 ( .S(n42), .A0(\mem_r[4][18] ), .A1(din[18]), .Z(\mem_nxt[4][18] ));
Q_MX02 U448 ( .S(n42), .A0(\mem_r[4][19] ), .A1(din[19]), .Z(\mem_nxt[4][19] ));
Q_MX02 U449 ( .S(n42), .A0(\mem_r[4][20] ), .A1(din[20]), .Z(\mem_nxt[4][20] ));
Q_MX02 U450 ( .S(n42), .A0(\mem_r[4][21] ), .A1(din[21]), .Z(\mem_nxt[4][21] ));
Q_MX02 U451 ( .S(n42), .A0(\mem_r[4][22] ), .A1(din[22]), .Z(\mem_nxt[4][22] ));
Q_MX02 U452 ( .S(n42), .A0(\mem_r[4][23] ), .A1(din[23]), .Z(\mem_nxt[4][23] ));
Q_MX02 U453 ( .S(n42), .A0(\mem_r[4][24] ), .A1(din[24]), .Z(\mem_nxt[4][24] ));
Q_MX02 U454 ( .S(n42), .A0(\mem_r[4][25] ), .A1(din[25]), .Z(\mem_nxt[4][25] ));
Q_MX02 U455 ( .S(n42), .A0(\mem_r[4][26] ), .A1(din[26]), .Z(\mem_nxt[4][26] ));
Q_MX02 U456 ( .S(n42), .A0(\mem_r[4][27] ), .A1(din[27]), .Z(\mem_nxt[4][27] ));
Q_MX02 U457 ( .S(n42), .A0(\mem_r[4][28] ), .A1(din[28]), .Z(\mem_nxt[4][28] ));
Q_MX02 U458 ( .S(n42), .A0(\mem_r[4][29] ), .A1(din[29]), .Z(\mem_nxt[4][29] ));
Q_MX02 U459 ( .S(n42), .A0(\mem_r[4][30] ), .A1(din[30]), .Z(\mem_nxt[4][30] ));
Q_MX02 U460 ( .S(n42), .A0(\mem_r[4][31] ), .A1(din[31]), .Z(\mem_nxt[4][31] ));
Q_MX02 U461 ( .S(n42), .A0(\mem_r[4][32] ), .A1(din[32]), .Z(\mem_nxt[4][32] ));
Q_MX02 U462 ( .S(n42), .A0(\mem_r[4][33] ), .A1(din[33]), .Z(\mem_nxt[4][33] ));
Q_MX02 U463 ( .S(n42), .A0(\mem_r[4][34] ), .A1(din[34]), .Z(\mem_nxt[4][34] ));
Q_MX02 U464 ( .S(n42), .A0(\mem_r[4][35] ), .A1(din[35]), .Z(\mem_nxt[4][35] ));
Q_MX02 U465 ( .S(n42), .A0(\mem_r[4][36] ), .A1(din[36]), .Z(\mem_nxt[4][36] ));
Q_MX02 U466 ( .S(n42), .A0(\mem_r[4][37] ), .A1(din[37]), .Z(\mem_nxt[4][37] ));
Q_MX02 U467 ( .S(n42), .A0(\mem_r[4][38] ), .A1(din[38]), .Z(\mem_nxt[4][38] ));
Q_MX02 U468 ( .S(n42), .A0(\mem_r[4][39] ), .A1(din[39]), .Z(\mem_nxt[4][39] ));
Q_MX02 U469 ( .S(n42), .A0(\mem_r[4][40] ), .A1(din[40]), .Z(\mem_nxt[4][40] ));
Q_MX02 U470 ( .S(n42), .A0(\mem_r[4][41] ), .A1(din[41]), .Z(\mem_nxt[4][41] ));
Q_MX02 U471 ( .S(n42), .A0(\mem_r[4][42] ), .A1(din[42]), .Z(\mem_nxt[4][42] ));
Q_MX02 U472 ( .S(n42), .A0(\mem_r[4][43] ), .A1(din[43]), .Z(\mem_nxt[4][43] ));
Q_MX02 U473 ( .S(n42), .A0(\mem_r[4][44] ), .A1(din[44]), .Z(\mem_nxt[4][44] ));
Q_MX02 U474 ( .S(n42), .A0(\mem_r[4][45] ), .A1(din[45]), .Z(\mem_nxt[4][45] ));
Q_MX02 U475 ( .S(n42), .A0(\mem_r[4][46] ), .A1(din[46]), .Z(\mem_nxt[4][46] ));
Q_MX02 U476 ( .S(n42), .A0(\mem_r[4][47] ), .A1(din[47]), .Z(\mem_nxt[4][47] ));
Q_MX02 U477 ( .S(n42), .A0(\mem_r[4][48] ), .A1(din[48]), .Z(\mem_nxt[4][48] ));
Q_MX02 U478 ( .S(n42), .A0(\mem_r[4][49] ), .A1(din[49]), .Z(\mem_nxt[4][49] ));
Q_MX02 U479 ( .S(n42), .A0(\mem_r[4][50] ), .A1(din[50]), .Z(\mem_nxt[4][50] ));
Q_MX02 U480 ( .S(n42), .A0(\mem_r[4][51] ), .A1(din[51]), .Z(\mem_nxt[4][51] ));
Q_MX02 U481 ( .S(n42), .A0(\mem_r[4][52] ), .A1(din[52]), .Z(\mem_nxt[4][52] ));
Q_MX02 U482 ( .S(n42), .A0(\mem_r[4][53] ), .A1(din[53]), .Z(\mem_nxt[4][53] ));
Q_MX02 U483 ( .S(n42), .A0(\mem_r[4][54] ), .A1(din[54]), .Z(\mem_nxt[4][54] ));
Q_MX02 U484 ( .S(n42), .A0(\mem_r[4][55] ), .A1(din[55]), .Z(\mem_nxt[4][55] ));
Q_MX02 U485 ( .S(n42), .A0(\mem_r[4][56] ), .A1(din[56]), .Z(\mem_nxt[4][56] ));
Q_MX02 U486 ( .S(n42), .A0(\mem_r[4][57] ), .A1(din[57]), .Z(\mem_nxt[4][57] ));
Q_MX02 U487 ( .S(n42), .A0(\mem_r[4][58] ), .A1(din[58]), .Z(\mem_nxt[4][58] ));
Q_MX02 U488 ( .S(n42), .A0(\mem_r[4][59] ), .A1(din[59]), .Z(\mem_nxt[4][59] ));
Q_MX02 U489 ( .S(n42), .A0(\mem_r[4][60] ), .A1(din[60]), .Z(\mem_nxt[4][60] ));
Q_MX02 U490 ( .S(n42), .A0(\mem_r[4][61] ), .A1(din[61]), .Z(\mem_nxt[4][61] ));
Q_MX02 U491 ( .S(n42), .A0(\mem_r[4][62] ), .A1(din[62]), .Z(\mem_nxt[4][62] ));
Q_MX02 U492 ( .S(n42), .A0(\mem_r[4][63] ), .A1(din[63]), .Z(\mem_nxt[4][63] ));
Q_MX02 U493 ( .S(n42), .A0(\mem_r[4][64] ), .A1(din[64]), .Z(\mem_nxt[4][64] ));
Q_MX02 U494 ( .S(n42), .A0(\mem_r[4][65] ), .A1(din[65]), .Z(\mem_nxt[4][65] ));
Q_MX02 U495 ( .S(n42), .A0(\mem_r[4][66] ), .A1(din[66]), .Z(\mem_nxt[4][66] ));
Q_MX02 U496 ( .S(n42), .A0(\mem_r[4][67] ), .A1(din[67]), .Z(\mem_nxt[4][67] ));
Q_MX02 U497 ( .S(n42), .A0(\mem_r[4][68] ), .A1(din[68]), .Z(\mem_nxt[4][68] ));
Q_MX02 U498 ( .S(n42), .A0(\mem_r[4][69] ), .A1(din[69]), .Z(\mem_nxt[4][69] ));
Q_MX02 U499 ( .S(n42), .A0(\mem_r[4][70] ), .A1(din[70]), .Z(\mem_nxt[4][70] ));
Q_MX02 U500 ( .S(n42), .A0(\mem_r[4][71] ), .A1(din[71]), .Z(\mem_nxt[4][71] ));
Q_MX02 U501 ( .S(n42), .A0(\mem_r[4][72] ), .A1(din[72]), .Z(\mem_nxt[4][72] ));
Q_MX02 U502 ( .S(n42), .A0(\mem_r[4][73] ), .A1(din[73]), .Z(\mem_nxt[4][73] ));
Q_MX02 U503 ( .S(n42), .A0(\mem_r[4][74] ), .A1(din[74]), .Z(\mem_nxt[4][74] ));
Q_MX02 U504 ( .S(n42), .A0(\mem_r[4][75] ), .A1(din[75]), .Z(\mem_nxt[4][75] ));
Q_MX02 U505 ( .S(n42), .A0(\mem_r[4][76] ), .A1(din[76]), .Z(\mem_nxt[4][76] ));
Q_MX02 U506 ( .S(n42), .A0(\mem_r[4][77] ), .A1(din[77]), .Z(\mem_nxt[4][77] ));
Q_MX02 U507 ( .S(n42), .A0(\mem_r[4][78] ), .A1(din[78]), .Z(\mem_nxt[4][78] ));
Q_MX02 U508 ( .S(n42), .A0(\mem_r[4][79] ), .A1(din[79]), .Z(\mem_nxt[4][79] ));
Q_MX02 U509 ( .S(n42), .A0(\mem_r[4][80] ), .A1(din[80]), .Z(\mem_nxt[4][80] ));
Q_MX02 U510 ( .S(n42), .A0(\mem_r[4][81] ), .A1(din[81]), .Z(\mem_nxt[4][81] ));
Q_MX02 U511 ( .S(n42), .A0(\mem_r[4][82] ), .A1(din[82]), .Z(\mem_nxt[4][82] ));
Q_MX02 U512 ( .S(n42), .A0(\mem_r[4][83] ), .A1(din[83]), .Z(\mem_nxt[4][83] ));
Q_MX02 U513 ( .S(n42), .A0(\mem_r[4][84] ), .A1(din[84]), .Z(\mem_nxt[4][84] ));
Q_MX02 U514 ( .S(n42), .A0(\mem_r[4][85] ), .A1(din[85]), .Z(\mem_nxt[4][85] ));
Q_MX02 U515 ( .S(n42), .A0(\mem_r[4][86] ), .A1(din[86]), .Z(\mem_nxt[4][86] ));
Q_MX02 U516 ( .S(n42), .A0(\mem_r[4][87] ), .A1(din[87]), .Z(\mem_nxt[4][87] ));
Q_MX02 U517 ( .S(n42), .A0(\mem_r[4][88] ), .A1(din[88]), .Z(\mem_nxt[4][88] ));
Q_MX02 U518 ( .S(n42), .A0(\mem_r[4][89] ), .A1(din[89]), .Z(\mem_nxt[4][89] ));
Q_MX02 U519 ( .S(n42), .A0(\mem_r[4][90] ), .A1(din[90]), .Z(\mem_nxt[4][90] ));
Q_MX02 U520 ( .S(n42), .A0(\mem_r[4][91] ), .A1(din[91]), .Z(\mem_nxt[4][91] ));
Q_MX02 U521 ( .S(n42), .A0(\mem_r[4][92] ), .A1(din[92]), .Z(\mem_nxt[4][92] ));
Q_MX02 U522 ( .S(n42), .A0(\mem_r[4][93] ), .A1(din[93]), .Z(\mem_nxt[4][93] ));
Q_MX02 U523 ( .S(n42), .A0(\mem_r[4][94] ), .A1(din[94]), .Z(\mem_nxt[4][94] ));
Q_MX02 U524 ( .S(n42), .A0(\mem_r[4][95] ), .A1(din[95]), .Z(\mem_nxt[4][95] ));
Q_MX02 U525 ( .S(n45), .A0(\mem_r[3][0] ), .A1(din[0]), .Z(\mem_nxt[3][0] ));
Q_MX02 U526 ( .S(n45), .A0(\mem_r[3][1] ), .A1(din[1]), .Z(\mem_nxt[3][1] ));
Q_MX02 U527 ( .S(n45), .A0(\mem_r[3][2] ), .A1(din[2]), .Z(\mem_nxt[3][2] ));
Q_MX02 U528 ( .S(n45), .A0(\mem_r[3][3] ), .A1(din[3]), .Z(\mem_nxt[3][3] ));
Q_MX02 U529 ( .S(n45), .A0(\mem_r[3][4] ), .A1(din[4]), .Z(\mem_nxt[3][4] ));
Q_MX02 U530 ( .S(n45), .A0(\mem_r[3][5] ), .A1(din[5]), .Z(\mem_nxt[3][5] ));
Q_MX02 U531 ( .S(n45), .A0(\mem_r[3][6] ), .A1(din[6]), .Z(\mem_nxt[3][6] ));
Q_MX02 U532 ( .S(n45), .A0(\mem_r[3][7] ), .A1(din[7]), .Z(\mem_nxt[3][7] ));
Q_MX02 U533 ( .S(n45), .A0(\mem_r[3][8] ), .A1(din[8]), .Z(\mem_nxt[3][8] ));
Q_MX02 U534 ( .S(n45), .A0(\mem_r[3][9] ), .A1(din[9]), .Z(\mem_nxt[3][9] ));
Q_MX02 U535 ( .S(n45), .A0(\mem_r[3][10] ), .A1(din[10]), .Z(\mem_nxt[3][10] ));
Q_MX02 U536 ( .S(n45), .A0(\mem_r[3][11] ), .A1(din[11]), .Z(\mem_nxt[3][11] ));
Q_MX02 U537 ( .S(n45), .A0(\mem_r[3][12] ), .A1(din[12]), .Z(\mem_nxt[3][12] ));
Q_MX02 U538 ( .S(n45), .A0(\mem_r[3][13] ), .A1(din[13]), .Z(\mem_nxt[3][13] ));
Q_MX02 U539 ( .S(n45), .A0(\mem_r[3][14] ), .A1(din[14]), .Z(\mem_nxt[3][14] ));
Q_MX02 U540 ( .S(n45), .A0(\mem_r[3][15] ), .A1(din[15]), .Z(\mem_nxt[3][15] ));
Q_MX02 U541 ( .S(n45), .A0(\mem_r[3][16] ), .A1(din[16]), .Z(\mem_nxt[3][16] ));
Q_MX02 U542 ( .S(n45), .A0(\mem_r[3][17] ), .A1(din[17]), .Z(\mem_nxt[3][17] ));
Q_MX02 U543 ( .S(n45), .A0(\mem_r[3][18] ), .A1(din[18]), .Z(\mem_nxt[3][18] ));
Q_MX02 U544 ( .S(n45), .A0(\mem_r[3][19] ), .A1(din[19]), .Z(\mem_nxt[3][19] ));
Q_MX02 U545 ( .S(n45), .A0(\mem_r[3][20] ), .A1(din[20]), .Z(\mem_nxt[3][20] ));
Q_MX02 U546 ( .S(n45), .A0(\mem_r[3][21] ), .A1(din[21]), .Z(\mem_nxt[3][21] ));
Q_MX02 U547 ( .S(n45), .A0(\mem_r[3][22] ), .A1(din[22]), .Z(\mem_nxt[3][22] ));
Q_MX02 U548 ( .S(n45), .A0(\mem_r[3][23] ), .A1(din[23]), .Z(\mem_nxt[3][23] ));
Q_MX02 U549 ( .S(n45), .A0(\mem_r[3][24] ), .A1(din[24]), .Z(\mem_nxt[3][24] ));
Q_MX02 U550 ( .S(n45), .A0(\mem_r[3][25] ), .A1(din[25]), .Z(\mem_nxt[3][25] ));
Q_MX02 U551 ( .S(n45), .A0(\mem_r[3][26] ), .A1(din[26]), .Z(\mem_nxt[3][26] ));
Q_MX02 U552 ( .S(n45), .A0(\mem_r[3][27] ), .A1(din[27]), .Z(\mem_nxt[3][27] ));
Q_MX02 U553 ( .S(n45), .A0(\mem_r[3][28] ), .A1(din[28]), .Z(\mem_nxt[3][28] ));
Q_MX02 U554 ( .S(n45), .A0(\mem_r[3][29] ), .A1(din[29]), .Z(\mem_nxt[3][29] ));
Q_MX02 U555 ( .S(n45), .A0(\mem_r[3][30] ), .A1(din[30]), .Z(\mem_nxt[3][30] ));
Q_MX02 U556 ( .S(n45), .A0(\mem_r[3][31] ), .A1(din[31]), .Z(\mem_nxt[3][31] ));
Q_MX02 U557 ( .S(n45), .A0(\mem_r[3][32] ), .A1(din[32]), .Z(\mem_nxt[3][32] ));
Q_MX02 U558 ( .S(n45), .A0(\mem_r[3][33] ), .A1(din[33]), .Z(\mem_nxt[3][33] ));
Q_MX02 U559 ( .S(n45), .A0(\mem_r[3][34] ), .A1(din[34]), .Z(\mem_nxt[3][34] ));
Q_MX02 U560 ( .S(n45), .A0(\mem_r[3][35] ), .A1(din[35]), .Z(\mem_nxt[3][35] ));
Q_MX02 U561 ( .S(n45), .A0(\mem_r[3][36] ), .A1(din[36]), .Z(\mem_nxt[3][36] ));
Q_MX02 U562 ( .S(n45), .A0(\mem_r[3][37] ), .A1(din[37]), .Z(\mem_nxt[3][37] ));
Q_MX02 U563 ( .S(n45), .A0(\mem_r[3][38] ), .A1(din[38]), .Z(\mem_nxt[3][38] ));
Q_MX02 U564 ( .S(n45), .A0(\mem_r[3][39] ), .A1(din[39]), .Z(\mem_nxt[3][39] ));
Q_MX02 U565 ( .S(n45), .A0(\mem_r[3][40] ), .A1(din[40]), .Z(\mem_nxt[3][40] ));
Q_MX02 U566 ( .S(n45), .A0(\mem_r[3][41] ), .A1(din[41]), .Z(\mem_nxt[3][41] ));
Q_MX02 U567 ( .S(n45), .A0(\mem_r[3][42] ), .A1(din[42]), .Z(\mem_nxt[3][42] ));
Q_MX02 U568 ( .S(n45), .A0(\mem_r[3][43] ), .A1(din[43]), .Z(\mem_nxt[3][43] ));
Q_MX02 U569 ( .S(n45), .A0(\mem_r[3][44] ), .A1(din[44]), .Z(\mem_nxt[3][44] ));
Q_MX02 U570 ( .S(n45), .A0(\mem_r[3][45] ), .A1(din[45]), .Z(\mem_nxt[3][45] ));
Q_MX02 U571 ( .S(n45), .A0(\mem_r[3][46] ), .A1(din[46]), .Z(\mem_nxt[3][46] ));
Q_MX02 U572 ( .S(n45), .A0(\mem_r[3][47] ), .A1(din[47]), .Z(\mem_nxt[3][47] ));
Q_MX02 U573 ( .S(n45), .A0(\mem_r[3][48] ), .A1(din[48]), .Z(\mem_nxt[3][48] ));
Q_MX02 U574 ( .S(n45), .A0(\mem_r[3][49] ), .A1(din[49]), .Z(\mem_nxt[3][49] ));
Q_MX02 U575 ( .S(n45), .A0(\mem_r[3][50] ), .A1(din[50]), .Z(\mem_nxt[3][50] ));
Q_MX02 U576 ( .S(n45), .A0(\mem_r[3][51] ), .A1(din[51]), .Z(\mem_nxt[3][51] ));
Q_MX02 U577 ( .S(n45), .A0(\mem_r[3][52] ), .A1(din[52]), .Z(\mem_nxt[3][52] ));
Q_MX02 U578 ( .S(n45), .A0(\mem_r[3][53] ), .A1(din[53]), .Z(\mem_nxt[3][53] ));
Q_MX02 U579 ( .S(n45), .A0(\mem_r[3][54] ), .A1(din[54]), .Z(\mem_nxt[3][54] ));
Q_MX02 U580 ( .S(n45), .A0(\mem_r[3][55] ), .A1(din[55]), .Z(\mem_nxt[3][55] ));
Q_MX02 U581 ( .S(n45), .A0(\mem_r[3][56] ), .A1(din[56]), .Z(\mem_nxt[3][56] ));
Q_MX02 U582 ( .S(n45), .A0(\mem_r[3][57] ), .A1(din[57]), .Z(\mem_nxt[3][57] ));
Q_MX02 U583 ( .S(n45), .A0(\mem_r[3][58] ), .A1(din[58]), .Z(\mem_nxt[3][58] ));
Q_MX02 U584 ( .S(n45), .A0(\mem_r[3][59] ), .A1(din[59]), .Z(\mem_nxt[3][59] ));
Q_MX02 U585 ( .S(n45), .A0(\mem_r[3][60] ), .A1(din[60]), .Z(\mem_nxt[3][60] ));
Q_MX02 U586 ( .S(n45), .A0(\mem_r[3][61] ), .A1(din[61]), .Z(\mem_nxt[3][61] ));
Q_MX02 U587 ( .S(n45), .A0(\mem_r[3][62] ), .A1(din[62]), .Z(\mem_nxt[3][62] ));
Q_MX02 U588 ( .S(n45), .A0(\mem_r[3][63] ), .A1(din[63]), .Z(\mem_nxt[3][63] ));
Q_MX02 U589 ( .S(n45), .A0(\mem_r[3][64] ), .A1(din[64]), .Z(\mem_nxt[3][64] ));
Q_MX02 U590 ( .S(n45), .A0(\mem_r[3][65] ), .A1(din[65]), .Z(\mem_nxt[3][65] ));
Q_MX02 U591 ( .S(n45), .A0(\mem_r[3][66] ), .A1(din[66]), .Z(\mem_nxt[3][66] ));
Q_MX02 U592 ( .S(n45), .A0(\mem_r[3][67] ), .A1(din[67]), .Z(\mem_nxt[3][67] ));
Q_MX02 U593 ( .S(n45), .A0(\mem_r[3][68] ), .A1(din[68]), .Z(\mem_nxt[3][68] ));
Q_MX02 U594 ( .S(n45), .A0(\mem_r[3][69] ), .A1(din[69]), .Z(\mem_nxt[3][69] ));
Q_MX02 U595 ( .S(n45), .A0(\mem_r[3][70] ), .A1(din[70]), .Z(\mem_nxt[3][70] ));
Q_MX02 U596 ( .S(n45), .A0(\mem_r[3][71] ), .A1(din[71]), .Z(\mem_nxt[3][71] ));
Q_MX02 U597 ( .S(n45), .A0(\mem_r[3][72] ), .A1(din[72]), .Z(\mem_nxt[3][72] ));
Q_MX02 U598 ( .S(n45), .A0(\mem_r[3][73] ), .A1(din[73]), .Z(\mem_nxt[3][73] ));
Q_MX02 U599 ( .S(n45), .A0(\mem_r[3][74] ), .A1(din[74]), .Z(\mem_nxt[3][74] ));
Q_MX02 U600 ( .S(n45), .A0(\mem_r[3][75] ), .A1(din[75]), .Z(\mem_nxt[3][75] ));
Q_MX02 U601 ( .S(n45), .A0(\mem_r[3][76] ), .A1(din[76]), .Z(\mem_nxt[3][76] ));
Q_MX02 U602 ( .S(n45), .A0(\mem_r[3][77] ), .A1(din[77]), .Z(\mem_nxt[3][77] ));
Q_MX02 U603 ( .S(n45), .A0(\mem_r[3][78] ), .A1(din[78]), .Z(\mem_nxt[3][78] ));
Q_MX02 U604 ( .S(n45), .A0(\mem_r[3][79] ), .A1(din[79]), .Z(\mem_nxt[3][79] ));
Q_MX02 U605 ( .S(n45), .A0(\mem_r[3][80] ), .A1(din[80]), .Z(\mem_nxt[3][80] ));
Q_MX02 U606 ( .S(n45), .A0(\mem_r[3][81] ), .A1(din[81]), .Z(\mem_nxt[3][81] ));
Q_MX02 U607 ( .S(n45), .A0(\mem_r[3][82] ), .A1(din[82]), .Z(\mem_nxt[3][82] ));
Q_MX02 U608 ( .S(n45), .A0(\mem_r[3][83] ), .A1(din[83]), .Z(\mem_nxt[3][83] ));
Q_MX02 U609 ( .S(n45), .A0(\mem_r[3][84] ), .A1(din[84]), .Z(\mem_nxt[3][84] ));
Q_MX02 U610 ( .S(n45), .A0(\mem_r[3][85] ), .A1(din[85]), .Z(\mem_nxt[3][85] ));
Q_MX02 U611 ( .S(n45), .A0(\mem_r[3][86] ), .A1(din[86]), .Z(\mem_nxt[3][86] ));
Q_MX02 U612 ( .S(n45), .A0(\mem_r[3][87] ), .A1(din[87]), .Z(\mem_nxt[3][87] ));
Q_MX02 U613 ( .S(n45), .A0(\mem_r[3][88] ), .A1(din[88]), .Z(\mem_nxt[3][88] ));
Q_MX02 U614 ( .S(n45), .A0(\mem_r[3][89] ), .A1(din[89]), .Z(\mem_nxt[3][89] ));
Q_MX02 U615 ( .S(n45), .A0(\mem_r[3][90] ), .A1(din[90]), .Z(\mem_nxt[3][90] ));
Q_MX02 U616 ( .S(n45), .A0(\mem_r[3][91] ), .A1(din[91]), .Z(\mem_nxt[3][91] ));
Q_MX02 U617 ( .S(n45), .A0(\mem_r[3][92] ), .A1(din[92]), .Z(\mem_nxt[3][92] ));
Q_MX02 U618 ( .S(n45), .A0(\mem_r[3][93] ), .A1(din[93]), .Z(\mem_nxt[3][93] ));
Q_MX02 U619 ( .S(n45), .A0(\mem_r[3][94] ), .A1(din[94]), .Z(\mem_nxt[3][94] ));
Q_MX02 U620 ( .S(n45), .A0(\mem_r[3][95] ), .A1(din[95]), .Z(\mem_nxt[3][95] ));
Q_MX02 U621 ( .S(n47), .A0(\mem_r[2][0] ), .A1(din[0]), .Z(\mem_nxt[2][0] ));
Q_MX02 U622 ( .S(n47), .A0(\mem_r[2][1] ), .A1(din[1]), .Z(\mem_nxt[2][1] ));
Q_MX02 U623 ( .S(n47), .A0(\mem_r[2][2] ), .A1(din[2]), .Z(\mem_nxt[2][2] ));
Q_MX02 U624 ( .S(n47), .A0(\mem_r[2][3] ), .A1(din[3]), .Z(\mem_nxt[2][3] ));
Q_MX02 U625 ( .S(n47), .A0(\mem_r[2][4] ), .A1(din[4]), .Z(\mem_nxt[2][4] ));
Q_MX02 U626 ( .S(n47), .A0(\mem_r[2][5] ), .A1(din[5]), .Z(\mem_nxt[2][5] ));
Q_MX02 U627 ( .S(n47), .A0(\mem_r[2][6] ), .A1(din[6]), .Z(\mem_nxt[2][6] ));
Q_MX02 U628 ( .S(n47), .A0(\mem_r[2][7] ), .A1(din[7]), .Z(\mem_nxt[2][7] ));
Q_MX02 U629 ( .S(n47), .A0(\mem_r[2][8] ), .A1(din[8]), .Z(\mem_nxt[2][8] ));
Q_MX02 U630 ( .S(n47), .A0(\mem_r[2][9] ), .A1(din[9]), .Z(\mem_nxt[2][9] ));
Q_MX02 U631 ( .S(n47), .A0(\mem_r[2][10] ), .A1(din[10]), .Z(\mem_nxt[2][10] ));
Q_MX02 U632 ( .S(n47), .A0(\mem_r[2][11] ), .A1(din[11]), .Z(\mem_nxt[2][11] ));
Q_MX02 U633 ( .S(n47), .A0(\mem_r[2][12] ), .A1(din[12]), .Z(\mem_nxt[2][12] ));
Q_MX02 U634 ( .S(n47), .A0(\mem_r[2][13] ), .A1(din[13]), .Z(\mem_nxt[2][13] ));
Q_MX02 U635 ( .S(n47), .A0(\mem_r[2][14] ), .A1(din[14]), .Z(\mem_nxt[2][14] ));
Q_MX02 U636 ( .S(n47), .A0(\mem_r[2][15] ), .A1(din[15]), .Z(\mem_nxt[2][15] ));
Q_MX02 U637 ( .S(n47), .A0(\mem_r[2][16] ), .A1(din[16]), .Z(\mem_nxt[2][16] ));
Q_MX02 U638 ( .S(n47), .A0(\mem_r[2][17] ), .A1(din[17]), .Z(\mem_nxt[2][17] ));
Q_MX02 U639 ( .S(n47), .A0(\mem_r[2][18] ), .A1(din[18]), .Z(\mem_nxt[2][18] ));
Q_MX02 U640 ( .S(n47), .A0(\mem_r[2][19] ), .A1(din[19]), .Z(\mem_nxt[2][19] ));
Q_MX02 U641 ( .S(n47), .A0(\mem_r[2][20] ), .A1(din[20]), .Z(\mem_nxt[2][20] ));
Q_MX02 U642 ( .S(n47), .A0(\mem_r[2][21] ), .A1(din[21]), .Z(\mem_nxt[2][21] ));
Q_MX02 U643 ( .S(n47), .A0(\mem_r[2][22] ), .A1(din[22]), .Z(\mem_nxt[2][22] ));
Q_MX02 U644 ( .S(n47), .A0(\mem_r[2][23] ), .A1(din[23]), .Z(\mem_nxt[2][23] ));
Q_MX02 U645 ( .S(n47), .A0(\mem_r[2][24] ), .A1(din[24]), .Z(\mem_nxt[2][24] ));
Q_MX02 U646 ( .S(n47), .A0(\mem_r[2][25] ), .A1(din[25]), .Z(\mem_nxt[2][25] ));
Q_MX02 U647 ( .S(n47), .A0(\mem_r[2][26] ), .A1(din[26]), .Z(\mem_nxt[2][26] ));
Q_MX02 U648 ( .S(n47), .A0(\mem_r[2][27] ), .A1(din[27]), .Z(\mem_nxt[2][27] ));
Q_MX02 U649 ( .S(n47), .A0(\mem_r[2][28] ), .A1(din[28]), .Z(\mem_nxt[2][28] ));
Q_MX02 U650 ( .S(n47), .A0(\mem_r[2][29] ), .A1(din[29]), .Z(\mem_nxt[2][29] ));
Q_MX02 U651 ( .S(n47), .A0(\mem_r[2][30] ), .A1(din[30]), .Z(\mem_nxt[2][30] ));
Q_MX02 U652 ( .S(n47), .A0(\mem_r[2][31] ), .A1(din[31]), .Z(\mem_nxt[2][31] ));
Q_MX02 U653 ( .S(n47), .A0(\mem_r[2][32] ), .A1(din[32]), .Z(\mem_nxt[2][32] ));
Q_MX02 U654 ( .S(n47), .A0(\mem_r[2][33] ), .A1(din[33]), .Z(\mem_nxt[2][33] ));
Q_MX02 U655 ( .S(n47), .A0(\mem_r[2][34] ), .A1(din[34]), .Z(\mem_nxt[2][34] ));
Q_MX02 U656 ( .S(n47), .A0(\mem_r[2][35] ), .A1(din[35]), .Z(\mem_nxt[2][35] ));
Q_MX02 U657 ( .S(n47), .A0(\mem_r[2][36] ), .A1(din[36]), .Z(\mem_nxt[2][36] ));
Q_MX02 U658 ( .S(n47), .A0(\mem_r[2][37] ), .A1(din[37]), .Z(\mem_nxt[2][37] ));
Q_MX02 U659 ( .S(n47), .A0(\mem_r[2][38] ), .A1(din[38]), .Z(\mem_nxt[2][38] ));
Q_MX02 U660 ( .S(n47), .A0(\mem_r[2][39] ), .A1(din[39]), .Z(\mem_nxt[2][39] ));
Q_MX02 U661 ( .S(n47), .A0(\mem_r[2][40] ), .A1(din[40]), .Z(\mem_nxt[2][40] ));
Q_MX02 U662 ( .S(n47), .A0(\mem_r[2][41] ), .A1(din[41]), .Z(\mem_nxt[2][41] ));
Q_MX02 U663 ( .S(n47), .A0(\mem_r[2][42] ), .A1(din[42]), .Z(\mem_nxt[2][42] ));
Q_MX02 U664 ( .S(n47), .A0(\mem_r[2][43] ), .A1(din[43]), .Z(\mem_nxt[2][43] ));
Q_MX02 U665 ( .S(n47), .A0(\mem_r[2][44] ), .A1(din[44]), .Z(\mem_nxt[2][44] ));
Q_MX02 U666 ( .S(n47), .A0(\mem_r[2][45] ), .A1(din[45]), .Z(\mem_nxt[2][45] ));
Q_MX02 U667 ( .S(n47), .A0(\mem_r[2][46] ), .A1(din[46]), .Z(\mem_nxt[2][46] ));
Q_MX02 U668 ( .S(n47), .A0(\mem_r[2][47] ), .A1(din[47]), .Z(\mem_nxt[2][47] ));
Q_MX02 U669 ( .S(n47), .A0(\mem_r[2][48] ), .A1(din[48]), .Z(\mem_nxt[2][48] ));
Q_MX02 U670 ( .S(n47), .A0(\mem_r[2][49] ), .A1(din[49]), .Z(\mem_nxt[2][49] ));
Q_MX02 U671 ( .S(n47), .A0(\mem_r[2][50] ), .A1(din[50]), .Z(\mem_nxt[2][50] ));
Q_MX02 U672 ( .S(n47), .A0(\mem_r[2][51] ), .A1(din[51]), .Z(\mem_nxt[2][51] ));
Q_MX02 U673 ( .S(n47), .A0(\mem_r[2][52] ), .A1(din[52]), .Z(\mem_nxt[2][52] ));
Q_MX02 U674 ( .S(n47), .A0(\mem_r[2][53] ), .A1(din[53]), .Z(\mem_nxt[2][53] ));
Q_MX02 U675 ( .S(n47), .A0(\mem_r[2][54] ), .A1(din[54]), .Z(\mem_nxt[2][54] ));
Q_MX02 U676 ( .S(n47), .A0(\mem_r[2][55] ), .A1(din[55]), .Z(\mem_nxt[2][55] ));
Q_MX02 U677 ( .S(n47), .A0(\mem_r[2][56] ), .A1(din[56]), .Z(\mem_nxt[2][56] ));
Q_MX02 U678 ( .S(n47), .A0(\mem_r[2][57] ), .A1(din[57]), .Z(\mem_nxt[2][57] ));
Q_MX02 U679 ( .S(n47), .A0(\mem_r[2][58] ), .A1(din[58]), .Z(\mem_nxt[2][58] ));
Q_MX02 U680 ( .S(n47), .A0(\mem_r[2][59] ), .A1(din[59]), .Z(\mem_nxt[2][59] ));
Q_MX02 U681 ( .S(n47), .A0(\mem_r[2][60] ), .A1(din[60]), .Z(\mem_nxt[2][60] ));
Q_MX02 U682 ( .S(n47), .A0(\mem_r[2][61] ), .A1(din[61]), .Z(\mem_nxt[2][61] ));
Q_MX02 U683 ( .S(n47), .A0(\mem_r[2][62] ), .A1(din[62]), .Z(\mem_nxt[2][62] ));
Q_MX02 U684 ( .S(n47), .A0(\mem_r[2][63] ), .A1(din[63]), .Z(\mem_nxt[2][63] ));
Q_MX02 U685 ( .S(n47), .A0(\mem_r[2][64] ), .A1(din[64]), .Z(\mem_nxt[2][64] ));
Q_MX02 U686 ( .S(n47), .A0(\mem_r[2][65] ), .A1(din[65]), .Z(\mem_nxt[2][65] ));
Q_MX02 U687 ( .S(n47), .A0(\mem_r[2][66] ), .A1(din[66]), .Z(\mem_nxt[2][66] ));
Q_MX02 U688 ( .S(n47), .A0(\mem_r[2][67] ), .A1(din[67]), .Z(\mem_nxt[2][67] ));
Q_MX02 U689 ( .S(n47), .A0(\mem_r[2][68] ), .A1(din[68]), .Z(\mem_nxt[2][68] ));
Q_MX02 U690 ( .S(n47), .A0(\mem_r[2][69] ), .A1(din[69]), .Z(\mem_nxt[2][69] ));
Q_MX02 U691 ( .S(n47), .A0(\mem_r[2][70] ), .A1(din[70]), .Z(\mem_nxt[2][70] ));
Q_MX02 U692 ( .S(n47), .A0(\mem_r[2][71] ), .A1(din[71]), .Z(\mem_nxt[2][71] ));
Q_MX02 U693 ( .S(n47), .A0(\mem_r[2][72] ), .A1(din[72]), .Z(\mem_nxt[2][72] ));
Q_MX02 U694 ( .S(n47), .A0(\mem_r[2][73] ), .A1(din[73]), .Z(\mem_nxt[2][73] ));
Q_MX02 U695 ( .S(n47), .A0(\mem_r[2][74] ), .A1(din[74]), .Z(\mem_nxt[2][74] ));
Q_MX02 U696 ( .S(n47), .A0(\mem_r[2][75] ), .A1(din[75]), .Z(\mem_nxt[2][75] ));
Q_MX02 U697 ( .S(n47), .A0(\mem_r[2][76] ), .A1(din[76]), .Z(\mem_nxt[2][76] ));
Q_MX02 U698 ( .S(n47), .A0(\mem_r[2][77] ), .A1(din[77]), .Z(\mem_nxt[2][77] ));
Q_MX02 U699 ( .S(n47), .A0(\mem_r[2][78] ), .A1(din[78]), .Z(\mem_nxt[2][78] ));
Q_MX02 U700 ( .S(n47), .A0(\mem_r[2][79] ), .A1(din[79]), .Z(\mem_nxt[2][79] ));
Q_MX02 U701 ( .S(n47), .A0(\mem_r[2][80] ), .A1(din[80]), .Z(\mem_nxt[2][80] ));
Q_MX02 U702 ( .S(n47), .A0(\mem_r[2][81] ), .A1(din[81]), .Z(\mem_nxt[2][81] ));
Q_MX02 U703 ( .S(n47), .A0(\mem_r[2][82] ), .A1(din[82]), .Z(\mem_nxt[2][82] ));
Q_MX02 U704 ( .S(n47), .A0(\mem_r[2][83] ), .A1(din[83]), .Z(\mem_nxt[2][83] ));
Q_MX02 U705 ( .S(n47), .A0(\mem_r[2][84] ), .A1(din[84]), .Z(\mem_nxt[2][84] ));
Q_MX02 U706 ( .S(n47), .A0(\mem_r[2][85] ), .A1(din[85]), .Z(\mem_nxt[2][85] ));
Q_MX02 U707 ( .S(n47), .A0(\mem_r[2][86] ), .A1(din[86]), .Z(\mem_nxt[2][86] ));
Q_MX02 U708 ( .S(n47), .A0(\mem_r[2][87] ), .A1(din[87]), .Z(\mem_nxt[2][87] ));
Q_MX02 U709 ( .S(n47), .A0(\mem_r[2][88] ), .A1(din[88]), .Z(\mem_nxt[2][88] ));
Q_MX02 U710 ( .S(n47), .A0(\mem_r[2][89] ), .A1(din[89]), .Z(\mem_nxt[2][89] ));
Q_MX02 U711 ( .S(n47), .A0(\mem_r[2][90] ), .A1(din[90]), .Z(\mem_nxt[2][90] ));
Q_MX02 U712 ( .S(n47), .A0(\mem_r[2][91] ), .A1(din[91]), .Z(\mem_nxt[2][91] ));
Q_MX02 U713 ( .S(n47), .A0(\mem_r[2][92] ), .A1(din[92]), .Z(\mem_nxt[2][92] ));
Q_MX02 U714 ( .S(n47), .A0(\mem_r[2][93] ), .A1(din[93]), .Z(\mem_nxt[2][93] ));
Q_MX02 U715 ( .S(n47), .A0(\mem_r[2][94] ), .A1(din[94]), .Z(\mem_nxt[2][94] ));
Q_MX02 U716 ( .S(n47), .A0(\mem_r[2][95] ), .A1(din[95]), .Z(\mem_nxt[2][95] ));
Q_MX02 U717 ( .S(n50), .A0(\mem_r[1][0] ), .A1(din[0]), .Z(\mem_nxt[1][0] ));
Q_MX02 U718 ( .S(n50), .A0(\mem_r[1][1] ), .A1(din[1]), .Z(\mem_nxt[1][1] ));
Q_MX02 U719 ( .S(n50), .A0(\mem_r[1][2] ), .A1(din[2]), .Z(\mem_nxt[1][2] ));
Q_MX02 U720 ( .S(n50), .A0(\mem_r[1][3] ), .A1(din[3]), .Z(\mem_nxt[1][3] ));
Q_MX02 U721 ( .S(n50), .A0(\mem_r[1][4] ), .A1(din[4]), .Z(\mem_nxt[1][4] ));
Q_MX02 U722 ( .S(n50), .A0(\mem_r[1][5] ), .A1(din[5]), .Z(\mem_nxt[1][5] ));
Q_MX02 U723 ( .S(n50), .A0(\mem_r[1][6] ), .A1(din[6]), .Z(\mem_nxt[1][6] ));
Q_MX02 U724 ( .S(n50), .A0(\mem_r[1][7] ), .A1(din[7]), .Z(\mem_nxt[1][7] ));
Q_MX02 U725 ( .S(n50), .A0(\mem_r[1][8] ), .A1(din[8]), .Z(\mem_nxt[1][8] ));
Q_MX02 U726 ( .S(n50), .A0(\mem_r[1][9] ), .A1(din[9]), .Z(\mem_nxt[1][9] ));
Q_MX02 U727 ( .S(n50), .A0(\mem_r[1][10] ), .A1(din[10]), .Z(\mem_nxt[1][10] ));
Q_MX02 U728 ( .S(n50), .A0(\mem_r[1][11] ), .A1(din[11]), .Z(\mem_nxt[1][11] ));
Q_MX02 U729 ( .S(n50), .A0(\mem_r[1][12] ), .A1(din[12]), .Z(\mem_nxt[1][12] ));
Q_MX02 U730 ( .S(n50), .A0(\mem_r[1][13] ), .A1(din[13]), .Z(\mem_nxt[1][13] ));
Q_MX02 U731 ( .S(n50), .A0(\mem_r[1][14] ), .A1(din[14]), .Z(\mem_nxt[1][14] ));
Q_MX02 U732 ( .S(n50), .A0(\mem_r[1][15] ), .A1(din[15]), .Z(\mem_nxt[1][15] ));
Q_MX02 U733 ( .S(n50), .A0(\mem_r[1][16] ), .A1(din[16]), .Z(\mem_nxt[1][16] ));
Q_MX02 U734 ( .S(n50), .A0(\mem_r[1][17] ), .A1(din[17]), .Z(\mem_nxt[1][17] ));
Q_MX02 U735 ( .S(n50), .A0(\mem_r[1][18] ), .A1(din[18]), .Z(\mem_nxt[1][18] ));
Q_MX02 U736 ( .S(n50), .A0(\mem_r[1][19] ), .A1(din[19]), .Z(\mem_nxt[1][19] ));
Q_MX02 U737 ( .S(n50), .A0(\mem_r[1][20] ), .A1(din[20]), .Z(\mem_nxt[1][20] ));
Q_MX02 U738 ( .S(n50), .A0(\mem_r[1][21] ), .A1(din[21]), .Z(\mem_nxt[1][21] ));
Q_MX02 U739 ( .S(n50), .A0(\mem_r[1][22] ), .A1(din[22]), .Z(\mem_nxt[1][22] ));
Q_MX02 U740 ( .S(n50), .A0(\mem_r[1][23] ), .A1(din[23]), .Z(\mem_nxt[1][23] ));
Q_MX02 U741 ( .S(n50), .A0(\mem_r[1][24] ), .A1(din[24]), .Z(\mem_nxt[1][24] ));
Q_MX02 U742 ( .S(n50), .A0(\mem_r[1][25] ), .A1(din[25]), .Z(\mem_nxt[1][25] ));
Q_MX02 U743 ( .S(n50), .A0(\mem_r[1][26] ), .A1(din[26]), .Z(\mem_nxt[1][26] ));
Q_MX02 U744 ( .S(n50), .A0(\mem_r[1][27] ), .A1(din[27]), .Z(\mem_nxt[1][27] ));
Q_MX02 U745 ( .S(n50), .A0(\mem_r[1][28] ), .A1(din[28]), .Z(\mem_nxt[1][28] ));
Q_MX02 U746 ( .S(n50), .A0(\mem_r[1][29] ), .A1(din[29]), .Z(\mem_nxt[1][29] ));
Q_MX02 U747 ( .S(n50), .A0(\mem_r[1][30] ), .A1(din[30]), .Z(\mem_nxt[1][30] ));
Q_MX02 U748 ( .S(n50), .A0(\mem_r[1][31] ), .A1(din[31]), .Z(\mem_nxt[1][31] ));
Q_MX02 U749 ( .S(n50), .A0(\mem_r[1][32] ), .A1(din[32]), .Z(\mem_nxt[1][32] ));
Q_MX02 U750 ( .S(n50), .A0(\mem_r[1][33] ), .A1(din[33]), .Z(\mem_nxt[1][33] ));
Q_MX02 U751 ( .S(n50), .A0(\mem_r[1][34] ), .A1(din[34]), .Z(\mem_nxt[1][34] ));
Q_MX02 U752 ( .S(n50), .A0(\mem_r[1][35] ), .A1(din[35]), .Z(\mem_nxt[1][35] ));
Q_MX02 U753 ( .S(n50), .A0(\mem_r[1][36] ), .A1(din[36]), .Z(\mem_nxt[1][36] ));
Q_MX02 U754 ( .S(n50), .A0(\mem_r[1][37] ), .A1(din[37]), .Z(\mem_nxt[1][37] ));
Q_MX02 U755 ( .S(n50), .A0(\mem_r[1][38] ), .A1(din[38]), .Z(\mem_nxt[1][38] ));
Q_MX02 U756 ( .S(n50), .A0(\mem_r[1][39] ), .A1(din[39]), .Z(\mem_nxt[1][39] ));
Q_MX02 U757 ( .S(n50), .A0(\mem_r[1][40] ), .A1(din[40]), .Z(\mem_nxt[1][40] ));
Q_MX02 U758 ( .S(n50), .A0(\mem_r[1][41] ), .A1(din[41]), .Z(\mem_nxt[1][41] ));
Q_MX02 U759 ( .S(n50), .A0(\mem_r[1][42] ), .A1(din[42]), .Z(\mem_nxt[1][42] ));
Q_MX02 U760 ( .S(n50), .A0(\mem_r[1][43] ), .A1(din[43]), .Z(\mem_nxt[1][43] ));
Q_MX02 U761 ( .S(n50), .A0(\mem_r[1][44] ), .A1(din[44]), .Z(\mem_nxt[1][44] ));
Q_MX02 U762 ( .S(n50), .A0(\mem_r[1][45] ), .A1(din[45]), .Z(\mem_nxt[1][45] ));
Q_MX02 U763 ( .S(n50), .A0(\mem_r[1][46] ), .A1(din[46]), .Z(\mem_nxt[1][46] ));
Q_MX02 U764 ( .S(n50), .A0(\mem_r[1][47] ), .A1(din[47]), .Z(\mem_nxt[1][47] ));
Q_MX02 U765 ( .S(n50), .A0(\mem_r[1][48] ), .A1(din[48]), .Z(\mem_nxt[1][48] ));
Q_MX02 U766 ( .S(n50), .A0(\mem_r[1][49] ), .A1(din[49]), .Z(\mem_nxt[1][49] ));
Q_MX02 U767 ( .S(n50), .A0(\mem_r[1][50] ), .A1(din[50]), .Z(\mem_nxt[1][50] ));
Q_MX02 U768 ( .S(n50), .A0(\mem_r[1][51] ), .A1(din[51]), .Z(\mem_nxt[1][51] ));
Q_MX02 U769 ( .S(n50), .A0(\mem_r[1][52] ), .A1(din[52]), .Z(\mem_nxt[1][52] ));
Q_MX02 U770 ( .S(n50), .A0(\mem_r[1][53] ), .A1(din[53]), .Z(\mem_nxt[1][53] ));
Q_MX02 U771 ( .S(n50), .A0(\mem_r[1][54] ), .A1(din[54]), .Z(\mem_nxt[1][54] ));
Q_MX02 U772 ( .S(n50), .A0(\mem_r[1][55] ), .A1(din[55]), .Z(\mem_nxt[1][55] ));
Q_MX02 U773 ( .S(n50), .A0(\mem_r[1][56] ), .A1(din[56]), .Z(\mem_nxt[1][56] ));
Q_MX02 U774 ( .S(n50), .A0(\mem_r[1][57] ), .A1(din[57]), .Z(\mem_nxt[1][57] ));
Q_MX02 U775 ( .S(n50), .A0(\mem_r[1][58] ), .A1(din[58]), .Z(\mem_nxt[1][58] ));
Q_MX02 U776 ( .S(n50), .A0(\mem_r[1][59] ), .A1(din[59]), .Z(\mem_nxt[1][59] ));
Q_MX02 U777 ( .S(n50), .A0(\mem_r[1][60] ), .A1(din[60]), .Z(\mem_nxt[1][60] ));
Q_MX02 U778 ( .S(n50), .A0(\mem_r[1][61] ), .A1(din[61]), .Z(\mem_nxt[1][61] ));
Q_MX02 U779 ( .S(n50), .A0(\mem_r[1][62] ), .A1(din[62]), .Z(\mem_nxt[1][62] ));
Q_MX02 U780 ( .S(n50), .A0(\mem_r[1][63] ), .A1(din[63]), .Z(\mem_nxt[1][63] ));
Q_MX02 U781 ( .S(n50), .A0(\mem_r[1][64] ), .A1(din[64]), .Z(\mem_nxt[1][64] ));
Q_MX02 U782 ( .S(n50), .A0(\mem_r[1][65] ), .A1(din[65]), .Z(\mem_nxt[1][65] ));
Q_MX02 U783 ( .S(n50), .A0(\mem_r[1][66] ), .A1(din[66]), .Z(\mem_nxt[1][66] ));
Q_MX02 U784 ( .S(n50), .A0(\mem_r[1][67] ), .A1(din[67]), .Z(\mem_nxt[1][67] ));
Q_MX02 U785 ( .S(n50), .A0(\mem_r[1][68] ), .A1(din[68]), .Z(\mem_nxt[1][68] ));
Q_MX02 U786 ( .S(n50), .A0(\mem_r[1][69] ), .A1(din[69]), .Z(\mem_nxt[1][69] ));
Q_MX02 U787 ( .S(n50), .A0(\mem_r[1][70] ), .A1(din[70]), .Z(\mem_nxt[1][70] ));
Q_MX02 U788 ( .S(n50), .A0(\mem_r[1][71] ), .A1(din[71]), .Z(\mem_nxt[1][71] ));
Q_MX02 U789 ( .S(n50), .A0(\mem_r[1][72] ), .A1(din[72]), .Z(\mem_nxt[1][72] ));
Q_MX02 U790 ( .S(n50), .A0(\mem_r[1][73] ), .A1(din[73]), .Z(\mem_nxt[1][73] ));
Q_MX02 U791 ( .S(n50), .A0(\mem_r[1][74] ), .A1(din[74]), .Z(\mem_nxt[1][74] ));
Q_MX02 U792 ( .S(n50), .A0(\mem_r[1][75] ), .A1(din[75]), .Z(\mem_nxt[1][75] ));
Q_MX02 U793 ( .S(n50), .A0(\mem_r[1][76] ), .A1(din[76]), .Z(\mem_nxt[1][76] ));
Q_MX02 U794 ( .S(n50), .A0(\mem_r[1][77] ), .A1(din[77]), .Z(\mem_nxt[1][77] ));
Q_MX02 U795 ( .S(n50), .A0(\mem_r[1][78] ), .A1(din[78]), .Z(\mem_nxt[1][78] ));
Q_MX02 U796 ( .S(n50), .A0(\mem_r[1][79] ), .A1(din[79]), .Z(\mem_nxt[1][79] ));
Q_MX02 U797 ( .S(n50), .A0(\mem_r[1][80] ), .A1(din[80]), .Z(\mem_nxt[1][80] ));
Q_MX02 U798 ( .S(n50), .A0(\mem_r[1][81] ), .A1(din[81]), .Z(\mem_nxt[1][81] ));
Q_MX02 U799 ( .S(n50), .A0(\mem_r[1][82] ), .A1(din[82]), .Z(\mem_nxt[1][82] ));
Q_MX02 U800 ( .S(n50), .A0(\mem_r[1][83] ), .A1(din[83]), .Z(\mem_nxt[1][83] ));
Q_MX02 U801 ( .S(n50), .A0(\mem_r[1][84] ), .A1(din[84]), .Z(\mem_nxt[1][84] ));
Q_MX02 U802 ( .S(n50), .A0(\mem_r[1][85] ), .A1(din[85]), .Z(\mem_nxt[1][85] ));
Q_MX02 U803 ( .S(n50), .A0(\mem_r[1][86] ), .A1(din[86]), .Z(\mem_nxt[1][86] ));
Q_MX02 U804 ( .S(n50), .A0(\mem_r[1][87] ), .A1(din[87]), .Z(\mem_nxt[1][87] ));
Q_MX02 U805 ( .S(n50), .A0(\mem_r[1][88] ), .A1(din[88]), .Z(\mem_nxt[1][88] ));
Q_MX02 U806 ( .S(n50), .A0(\mem_r[1][89] ), .A1(din[89]), .Z(\mem_nxt[1][89] ));
Q_MX02 U807 ( .S(n50), .A0(\mem_r[1][90] ), .A1(din[90]), .Z(\mem_nxt[1][90] ));
Q_MX02 U808 ( .S(n50), .A0(\mem_r[1][91] ), .A1(din[91]), .Z(\mem_nxt[1][91] ));
Q_MX02 U809 ( .S(n50), .A0(\mem_r[1][92] ), .A1(din[92]), .Z(\mem_nxt[1][92] ));
Q_MX02 U810 ( .S(n50), .A0(\mem_r[1][93] ), .A1(din[93]), .Z(\mem_nxt[1][93] ));
Q_MX02 U811 ( .S(n50), .A0(\mem_r[1][94] ), .A1(din[94]), .Z(\mem_nxt[1][94] ));
Q_MX02 U812 ( .S(n50), .A0(\mem_r[1][95] ), .A1(din[95]), .Z(\mem_nxt[1][95] ));
Q_MX02 U813 ( .S(n52), .A0(\mem_r[0][0] ), .A1(din[0]), .Z(\mem_nxt[0][0] ));
Q_MX02 U814 ( .S(n52), .A0(\mem_r[0][1] ), .A1(din[1]), .Z(\mem_nxt[0][1] ));
Q_MX02 U815 ( .S(n52), .A0(\mem_r[0][2] ), .A1(din[2]), .Z(\mem_nxt[0][2] ));
Q_MX02 U816 ( .S(n52), .A0(\mem_r[0][3] ), .A1(din[3]), .Z(\mem_nxt[0][3] ));
Q_MX02 U817 ( .S(n52), .A0(\mem_r[0][4] ), .A1(din[4]), .Z(\mem_nxt[0][4] ));
Q_MX02 U818 ( .S(n52), .A0(\mem_r[0][5] ), .A1(din[5]), .Z(\mem_nxt[0][5] ));
Q_MX02 U819 ( .S(n52), .A0(\mem_r[0][6] ), .A1(din[6]), .Z(\mem_nxt[0][6] ));
Q_MX02 U820 ( .S(n52), .A0(\mem_r[0][7] ), .A1(din[7]), .Z(\mem_nxt[0][7] ));
Q_MX02 U821 ( .S(n52), .A0(\mem_r[0][8] ), .A1(din[8]), .Z(\mem_nxt[0][8] ));
Q_MX02 U822 ( .S(n52), .A0(\mem_r[0][9] ), .A1(din[9]), .Z(\mem_nxt[0][9] ));
Q_MX02 U823 ( .S(n52), .A0(\mem_r[0][10] ), .A1(din[10]), .Z(\mem_nxt[0][10] ));
Q_MX02 U824 ( .S(n52), .A0(\mem_r[0][11] ), .A1(din[11]), .Z(\mem_nxt[0][11] ));
Q_MX02 U825 ( .S(n52), .A0(\mem_r[0][12] ), .A1(din[12]), .Z(\mem_nxt[0][12] ));
Q_MX02 U826 ( .S(n52), .A0(\mem_r[0][13] ), .A1(din[13]), .Z(\mem_nxt[0][13] ));
Q_MX02 U827 ( .S(n52), .A0(\mem_r[0][14] ), .A1(din[14]), .Z(\mem_nxt[0][14] ));
Q_MX02 U828 ( .S(n52), .A0(\mem_r[0][15] ), .A1(din[15]), .Z(\mem_nxt[0][15] ));
Q_MX02 U829 ( .S(n52), .A0(\mem_r[0][16] ), .A1(din[16]), .Z(\mem_nxt[0][16] ));
Q_MX02 U830 ( .S(n52), .A0(\mem_r[0][17] ), .A1(din[17]), .Z(\mem_nxt[0][17] ));
Q_MX02 U831 ( .S(n52), .A0(\mem_r[0][18] ), .A1(din[18]), .Z(\mem_nxt[0][18] ));
Q_MX02 U832 ( .S(n52), .A0(\mem_r[0][19] ), .A1(din[19]), .Z(\mem_nxt[0][19] ));
Q_MX02 U833 ( .S(n52), .A0(\mem_r[0][20] ), .A1(din[20]), .Z(\mem_nxt[0][20] ));
Q_MX02 U834 ( .S(n52), .A0(\mem_r[0][21] ), .A1(din[21]), .Z(\mem_nxt[0][21] ));
Q_MX02 U835 ( .S(n52), .A0(\mem_r[0][22] ), .A1(din[22]), .Z(\mem_nxt[0][22] ));
Q_MX02 U836 ( .S(n52), .A0(\mem_r[0][23] ), .A1(din[23]), .Z(\mem_nxt[0][23] ));
Q_MX02 U837 ( .S(n52), .A0(\mem_r[0][24] ), .A1(din[24]), .Z(\mem_nxt[0][24] ));
Q_MX02 U838 ( .S(n52), .A0(\mem_r[0][25] ), .A1(din[25]), .Z(\mem_nxt[0][25] ));
Q_MX02 U839 ( .S(n52), .A0(\mem_r[0][26] ), .A1(din[26]), .Z(\mem_nxt[0][26] ));
Q_MX02 U840 ( .S(n52), .A0(\mem_r[0][27] ), .A1(din[27]), .Z(\mem_nxt[0][27] ));
Q_MX02 U841 ( .S(n52), .A0(\mem_r[0][28] ), .A1(din[28]), .Z(\mem_nxt[0][28] ));
Q_MX02 U842 ( .S(n52), .A0(\mem_r[0][29] ), .A1(din[29]), .Z(\mem_nxt[0][29] ));
Q_MX02 U843 ( .S(n52), .A0(\mem_r[0][30] ), .A1(din[30]), .Z(\mem_nxt[0][30] ));
Q_MX02 U844 ( .S(n52), .A0(\mem_r[0][31] ), .A1(din[31]), .Z(\mem_nxt[0][31] ));
Q_MX02 U845 ( .S(n52), .A0(\mem_r[0][32] ), .A1(din[32]), .Z(\mem_nxt[0][32] ));
Q_MX02 U846 ( .S(n52), .A0(\mem_r[0][33] ), .A1(din[33]), .Z(\mem_nxt[0][33] ));
Q_MX02 U847 ( .S(n52), .A0(\mem_r[0][34] ), .A1(din[34]), .Z(\mem_nxt[0][34] ));
Q_MX02 U848 ( .S(n52), .A0(\mem_r[0][35] ), .A1(din[35]), .Z(\mem_nxt[0][35] ));
Q_MX02 U849 ( .S(n52), .A0(\mem_r[0][36] ), .A1(din[36]), .Z(\mem_nxt[0][36] ));
Q_MX02 U850 ( .S(n52), .A0(\mem_r[0][37] ), .A1(din[37]), .Z(\mem_nxt[0][37] ));
Q_MX02 U851 ( .S(n52), .A0(\mem_r[0][38] ), .A1(din[38]), .Z(\mem_nxt[0][38] ));
Q_MX02 U852 ( .S(n52), .A0(\mem_r[0][39] ), .A1(din[39]), .Z(\mem_nxt[0][39] ));
Q_MX02 U853 ( .S(n52), .A0(\mem_r[0][40] ), .A1(din[40]), .Z(\mem_nxt[0][40] ));
Q_MX02 U854 ( .S(n52), .A0(\mem_r[0][41] ), .A1(din[41]), .Z(\mem_nxt[0][41] ));
Q_MX02 U855 ( .S(n52), .A0(\mem_r[0][42] ), .A1(din[42]), .Z(\mem_nxt[0][42] ));
Q_MX02 U856 ( .S(n52), .A0(\mem_r[0][43] ), .A1(din[43]), .Z(\mem_nxt[0][43] ));
Q_MX02 U857 ( .S(n52), .A0(\mem_r[0][44] ), .A1(din[44]), .Z(\mem_nxt[0][44] ));
Q_MX02 U858 ( .S(n52), .A0(\mem_r[0][45] ), .A1(din[45]), .Z(\mem_nxt[0][45] ));
Q_MX02 U859 ( .S(n52), .A0(\mem_r[0][46] ), .A1(din[46]), .Z(\mem_nxt[0][46] ));
Q_MX02 U860 ( .S(n52), .A0(\mem_r[0][47] ), .A1(din[47]), .Z(\mem_nxt[0][47] ));
Q_MX02 U861 ( .S(n52), .A0(\mem_r[0][48] ), .A1(din[48]), .Z(\mem_nxt[0][48] ));
Q_MX02 U862 ( .S(n52), .A0(\mem_r[0][49] ), .A1(din[49]), .Z(\mem_nxt[0][49] ));
Q_MX02 U863 ( .S(n52), .A0(\mem_r[0][50] ), .A1(din[50]), .Z(\mem_nxt[0][50] ));
Q_MX02 U864 ( .S(n52), .A0(\mem_r[0][51] ), .A1(din[51]), .Z(\mem_nxt[0][51] ));
Q_MX02 U865 ( .S(n52), .A0(\mem_r[0][52] ), .A1(din[52]), .Z(\mem_nxt[0][52] ));
Q_MX02 U866 ( .S(n52), .A0(\mem_r[0][53] ), .A1(din[53]), .Z(\mem_nxt[0][53] ));
Q_MX02 U867 ( .S(n52), .A0(\mem_r[0][54] ), .A1(din[54]), .Z(\mem_nxt[0][54] ));
Q_MX02 U868 ( .S(n52), .A0(\mem_r[0][55] ), .A1(din[55]), .Z(\mem_nxt[0][55] ));
Q_MX02 U869 ( .S(n52), .A0(\mem_r[0][56] ), .A1(din[56]), .Z(\mem_nxt[0][56] ));
Q_MX02 U870 ( .S(n52), .A0(\mem_r[0][57] ), .A1(din[57]), .Z(\mem_nxt[0][57] ));
Q_MX02 U871 ( .S(n52), .A0(\mem_r[0][58] ), .A1(din[58]), .Z(\mem_nxt[0][58] ));
Q_MX02 U872 ( .S(n52), .A0(\mem_r[0][59] ), .A1(din[59]), .Z(\mem_nxt[0][59] ));
Q_MX02 U873 ( .S(n52), .A0(\mem_r[0][60] ), .A1(din[60]), .Z(\mem_nxt[0][60] ));
Q_MX02 U874 ( .S(n52), .A0(\mem_r[0][61] ), .A1(din[61]), .Z(\mem_nxt[0][61] ));
Q_MX02 U875 ( .S(n52), .A0(\mem_r[0][62] ), .A1(din[62]), .Z(\mem_nxt[0][62] ));
Q_MX02 U876 ( .S(n52), .A0(\mem_r[0][63] ), .A1(din[63]), .Z(\mem_nxt[0][63] ));
Q_MX02 U877 ( .S(n52), .A0(\mem_r[0][64] ), .A1(din[64]), .Z(\mem_nxt[0][64] ));
Q_MX02 U878 ( .S(n52), .A0(\mem_r[0][65] ), .A1(din[65]), .Z(\mem_nxt[0][65] ));
Q_MX02 U879 ( .S(n52), .A0(\mem_r[0][66] ), .A1(din[66]), .Z(\mem_nxt[0][66] ));
Q_MX02 U880 ( .S(n52), .A0(\mem_r[0][67] ), .A1(din[67]), .Z(\mem_nxt[0][67] ));
Q_MX02 U881 ( .S(n52), .A0(\mem_r[0][68] ), .A1(din[68]), .Z(\mem_nxt[0][68] ));
Q_MX02 U882 ( .S(n52), .A0(\mem_r[0][69] ), .A1(din[69]), .Z(\mem_nxt[0][69] ));
Q_MX02 U883 ( .S(n52), .A0(\mem_r[0][70] ), .A1(din[70]), .Z(\mem_nxt[0][70] ));
Q_MX02 U884 ( .S(n52), .A0(\mem_r[0][71] ), .A1(din[71]), .Z(\mem_nxt[0][71] ));
Q_MX02 U885 ( .S(n52), .A0(\mem_r[0][72] ), .A1(din[72]), .Z(\mem_nxt[0][72] ));
Q_MX02 U886 ( .S(n52), .A0(\mem_r[0][73] ), .A1(din[73]), .Z(\mem_nxt[0][73] ));
Q_MX02 U887 ( .S(n52), .A0(\mem_r[0][74] ), .A1(din[74]), .Z(\mem_nxt[0][74] ));
Q_MX02 U888 ( .S(n52), .A0(\mem_r[0][75] ), .A1(din[75]), .Z(\mem_nxt[0][75] ));
Q_MX02 U889 ( .S(n52), .A0(\mem_r[0][76] ), .A1(din[76]), .Z(\mem_nxt[0][76] ));
Q_MX02 U890 ( .S(n52), .A0(\mem_r[0][77] ), .A1(din[77]), .Z(\mem_nxt[0][77] ));
Q_MX02 U891 ( .S(n52), .A0(\mem_r[0][78] ), .A1(din[78]), .Z(\mem_nxt[0][78] ));
Q_MX02 U892 ( .S(n52), .A0(\mem_r[0][79] ), .A1(din[79]), .Z(\mem_nxt[0][79] ));
Q_MX02 U893 ( .S(n52), .A0(\mem_r[0][80] ), .A1(din[80]), .Z(\mem_nxt[0][80] ));
Q_MX02 U894 ( .S(n52), .A0(\mem_r[0][81] ), .A1(din[81]), .Z(\mem_nxt[0][81] ));
Q_MX02 U895 ( .S(n52), .A0(\mem_r[0][82] ), .A1(din[82]), .Z(\mem_nxt[0][82] ));
Q_MX02 U896 ( .S(n52), .A0(\mem_r[0][83] ), .A1(din[83]), .Z(\mem_nxt[0][83] ));
Q_MX02 U897 ( .S(n52), .A0(\mem_r[0][84] ), .A1(din[84]), .Z(\mem_nxt[0][84] ));
Q_MX02 U898 ( .S(n52), .A0(\mem_r[0][85] ), .A1(din[85]), .Z(\mem_nxt[0][85] ));
Q_MX02 U899 ( .S(n52), .A0(\mem_r[0][86] ), .A1(din[86]), .Z(\mem_nxt[0][86] ));
Q_MX02 U900 ( .S(n52), .A0(\mem_r[0][87] ), .A1(din[87]), .Z(\mem_nxt[0][87] ));
Q_MX02 U901 ( .S(n52), .A0(\mem_r[0][88] ), .A1(din[88]), .Z(\mem_nxt[0][88] ));
Q_MX02 U902 ( .S(n52), .A0(\mem_r[0][89] ), .A1(din[89]), .Z(\mem_nxt[0][89] ));
Q_MX02 U903 ( .S(n52), .A0(\mem_r[0][90] ), .A1(din[90]), .Z(\mem_nxt[0][90] ));
Q_MX02 U904 ( .S(n52), .A0(\mem_r[0][91] ), .A1(din[91]), .Z(\mem_nxt[0][91] ));
Q_MX02 U905 ( .S(n52), .A0(\mem_r[0][92] ), .A1(din[92]), .Z(\mem_nxt[0][92] ));
Q_MX02 U906 ( .S(n52), .A0(\mem_r[0][93] ), .A1(din[93]), .Z(\mem_nxt[0][93] ));
Q_MX02 U907 ( .S(n52), .A0(\mem_r[0][94] ), .A1(din[94]), .Z(\mem_nxt[0][94] ));
Q_MX02 U908 ( .S(n52), .A0(\mem_r[0][95] ), .A1(din[95]), .Z(\mem_nxt[0][95] ));
Q_AN02 U909 ( .A0(wr_ptr_r[0]), .A1(n35), .Z(n56));
Q_NR02 U910 ( .A0(wr_ptr_r[0]), .A1(n37), .Z(n36));
Q_INV U911 ( .A(n35), .Z(n37));
Q_AN02 U912 ( .A0(wr_ptr_r[1]), .A1(n38), .Z(n35));
Q_NR02 U913 ( .A0(n40), .A1(n41), .Z(n39));
Q_NR02 U914 ( .A0(wr_ptr_r[0]), .A1(n41), .Z(n42));
Q_OR02 U915 ( .A0(wr_ptr_r[1]), .A1(n43), .Z(n41));
Q_INV U916 ( .A(n38), .Z(n43));
Q_AN02 U917 ( .A0(wr_ptr_r[2]), .A1(n44), .Z(n38));
Q_NR02 U918 ( .A0(n40), .A1(n46), .Z(n45));
Q_NR02 U919 ( .A0(wr_ptr_r[0]), .A1(n46), .Z(n47));
Q_OR02 U920 ( .A0(n48), .A1(n49), .Z(n46));
Q_NR02 U921 ( .A0(n40), .A1(n51), .Z(n50));
Q_NR02 U922 ( .A0(wr_ptr_r[0]), .A1(n51), .Z(n52));
Q_OR02 U923 ( .A0(wr_ptr_r[1]), .A1(n49), .Z(n51));
Q_OR02 U924 ( .A0(wr_ptr_r[2]), .A1(n53), .Z(n49));
Q_INV U925 ( .A(n44), .Z(n53));
Q_AN02 U926 ( .A0(wr_en), .A1(n54), .Z(n44));
Q_OR02 U927 ( .A0(rd_en), .A1(n55), .Z(n54));
Q_INV U928 ( .A(full_i), .Z(n55));
Q_FDP1 \mem_r_REG[7][0] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][0] ), .Q(\mem_r[7][0] ), .QN( ));
Q_FDP1 \mem_r_REG[7][1] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][1] ), .Q(\mem_r[7][1] ), .QN( ));
Q_FDP1 \mem_r_REG[7][2] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][2] ), .Q(\mem_r[7][2] ), .QN( ));
Q_FDP1 \mem_r_REG[7][3] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][3] ), .Q(\mem_r[7][3] ), .QN( ));
Q_FDP1 \mem_r_REG[7][4] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][4] ), .Q(\mem_r[7][4] ), .QN( ));
Q_FDP1 \mem_r_REG[7][5] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][5] ), .Q(\mem_r[7][5] ), .QN( ));
Q_FDP1 \mem_r_REG[7][6] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][6] ), .Q(\mem_r[7][6] ), .QN( ));
Q_FDP1 \mem_r_REG[7][7] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][7] ), .Q(\mem_r[7][7] ), .QN( ));
Q_FDP1 \mem_r_REG[7][8] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][8] ), .Q(\mem_r[7][8] ), .QN( ));
Q_FDP1 \mem_r_REG[7][9] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][9] ), .Q(\mem_r[7][9] ), .QN( ));
Q_FDP1 \mem_r_REG[7][10] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][10] ), .Q(\mem_r[7][10] ), .QN( ));
Q_FDP1 \mem_r_REG[7][11] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][11] ), .Q(\mem_r[7][11] ), .QN( ));
Q_FDP1 \mem_r_REG[7][12] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][12] ), .Q(\mem_r[7][12] ), .QN( ));
Q_FDP1 \mem_r_REG[7][13] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][13] ), .Q(\mem_r[7][13] ), .QN( ));
Q_FDP1 \mem_r_REG[7][14] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][14] ), .Q(\mem_r[7][14] ), .QN( ));
Q_FDP1 \mem_r_REG[7][15] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][15] ), .Q(\mem_r[7][15] ), .QN( ));
Q_FDP1 \mem_r_REG[7][16] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][16] ), .Q(\mem_r[7][16] ), .QN( ));
Q_FDP1 \mem_r_REG[7][17] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][17] ), .Q(\mem_r[7][17] ), .QN( ));
Q_FDP1 \mem_r_REG[7][18] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][18] ), .Q(\mem_r[7][18] ), .QN( ));
Q_FDP1 \mem_r_REG[7][19] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][19] ), .Q(\mem_r[7][19] ), .QN( ));
Q_FDP1 \mem_r_REG[7][20] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][20] ), .Q(\mem_r[7][20] ), .QN( ));
Q_FDP1 \mem_r_REG[7][21] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][21] ), .Q(\mem_r[7][21] ), .QN( ));
Q_FDP1 \mem_r_REG[7][22] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][22] ), .Q(\mem_r[7][22] ), .QN( ));
Q_FDP1 \mem_r_REG[7][23] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][23] ), .Q(\mem_r[7][23] ), .QN( ));
Q_FDP1 \mem_r_REG[7][24] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][24] ), .Q(\mem_r[7][24] ), .QN( ));
Q_FDP1 \mem_r_REG[7][25] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][25] ), .Q(\mem_r[7][25] ), .QN( ));
Q_FDP1 \mem_r_REG[7][26] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][26] ), .Q(\mem_r[7][26] ), .QN( ));
Q_FDP1 \mem_r_REG[7][27] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][27] ), .Q(\mem_r[7][27] ), .QN( ));
Q_FDP1 \mem_r_REG[7][28] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][28] ), .Q(\mem_r[7][28] ), .QN( ));
Q_FDP1 \mem_r_REG[7][29] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][29] ), .Q(\mem_r[7][29] ), .QN( ));
Q_FDP1 \mem_r_REG[7][30] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][30] ), .Q(\mem_r[7][30] ), .QN( ));
Q_FDP1 \mem_r_REG[7][31] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][31] ), .Q(\mem_r[7][31] ), .QN( ));
Q_FDP1 \mem_r_REG[7][32] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][32] ), .Q(\mem_r[7][32] ), .QN( ));
Q_FDP1 \mem_r_REG[7][33] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][33] ), .Q(\mem_r[7][33] ), .QN( ));
Q_FDP1 \mem_r_REG[7][34] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][34] ), .Q(\mem_r[7][34] ), .QN( ));
Q_FDP1 \mem_r_REG[7][35] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][35] ), .Q(\mem_r[7][35] ), .QN( ));
Q_FDP1 \mem_r_REG[7][36] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][36] ), .Q(\mem_r[7][36] ), .QN( ));
Q_FDP1 \mem_r_REG[7][37] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][37] ), .Q(\mem_r[7][37] ), .QN( ));
Q_FDP1 \mem_r_REG[7][38] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][38] ), .Q(\mem_r[7][38] ), .QN( ));
Q_FDP1 \mem_r_REG[7][39] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][39] ), .Q(\mem_r[7][39] ), .QN( ));
Q_FDP1 \mem_r_REG[7][40] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][40] ), .Q(\mem_r[7][40] ), .QN( ));
Q_FDP1 \mem_r_REG[7][41] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][41] ), .Q(\mem_r[7][41] ), .QN( ));
Q_FDP1 \mem_r_REG[7][42] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][42] ), .Q(\mem_r[7][42] ), .QN( ));
Q_FDP1 \mem_r_REG[7][43] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][43] ), .Q(\mem_r[7][43] ), .QN( ));
Q_FDP1 \mem_r_REG[7][44] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][44] ), .Q(\mem_r[7][44] ), .QN( ));
Q_FDP1 \mem_r_REG[7][45] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][45] ), .Q(\mem_r[7][45] ), .QN( ));
Q_FDP1 \mem_r_REG[7][46] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][46] ), .Q(\mem_r[7][46] ), .QN( ));
Q_FDP1 \mem_r_REG[7][47] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][47] ), .Q(\mem_r[7][47] ), .QN( ));
Q_FDP1 \mem_r_REG[7][48] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][48] ), .Q(\mem_r[7][48] ), .QN( ));
Q_FDP1 \mem_r_REG[7][49] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][49] ), .Q(\mem_r[7][49] ), .QN( ));
Q_FDP1 \mem_r_REG[7][50] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][50] ), .Q(\mem_r[7][50] ), .QN( ));
Q_FDP1 \mem_r_REG[7][51] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][51] ), .Q(\mem_r[7][51] ), .QN( ));
Q_FDP1 \mem_r_REG[7][52] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][52] ), .Q(\mem_r[7][52] ), .QN( ));
Q_FDP1 \mem_r_REG[7][53] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][53] ), .Q(\mem_r[7][53] ), .QN( ));
Q_FDP1 \mem_r_REG[7][54] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][54] ), .Q(\mem_r[7][54] ), .QN( ));
Q_FDP1 \mem_r_REG[7][55] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][55] ), .Q(\mem_r[7][55] ), .QN( ));
Q_FDP1 \mem_r_REG[7][56] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][56] ), .Q(\mem_r[7][56] ), .QN( ));
Q_FDP1 \mem_r_REG[7][57] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][57] ), .Q(\mem_r[7][57] ), .QN( ));
Q_FDP1 \mem_r_REG[7][58] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][58] ), .Q(\mem_r[7][58] ), .QN( ));
Q_FDP1 \mem_r_REG[7][59] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][59] ), .Q(\mem_r[7][59] ), .QN( ));
Q_FDP1 \mem_r_REG[7][60] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][60] ), .Q(\mem_r[7][60] ), .QN( ));
Q_FDP1 \mem_r_REG[7][61] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][61] ), .Q(\mem_r[7][61] ), .QN( ));
Q_FDP1 \mem_r_REG[7][62] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][62] ), .Q(\mem_r[7][62] ), .QN( ));
Q_FDP1 \mem_r_REG[7][63] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][63] ), .Q(\mem_r[7][63] ), .QN( ));
Q_FDP1 \mem_r_REG[7][64] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][64] ), .Q(\mem_r[7][64] ), .QN( ));
Q_FDP1 \mem_r_REG[7][65] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][65] ), .Q(\mem_r[7][65] ), .QN( ));
Q_FDP1 \mem_r_REG[7][66] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][66] ), .Q(\mem_r[7][66] ), .QN( ));
Q_FDP1 \mem_r_REG[7][67] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][67] ), .Q(\mem_r[7][67] ), .QN( ));
Q_FDP1 \mem_r_REG[7][68] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][68] ), .Q(\mem_r[7][68] ), .QN( ));
Q_FDP1 \mem_r_REG[7][69] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][69] ), .Q(\mem_r[7][69] ), .QN( ));
Q_FDP1 \mem_r_REG[7][70] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][70] ), .Q(\mem_r[7][70] ), .QN( ));
Q_FDP1 \mem_r_REG[7][71] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][71] ), .Q(\mem_r[7][71] ), .QN( ));
Q_FDP1 \mem_r_REG[7][72] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][72] ), .Q(\mem_r[7][72] ), .QN( ));
Q_FDP1 \mem_r_REG[7][73] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][73] ), .Q(\mem_r[7][73] ), .QN( ));
Q_FDP1 \mem_r_REG[7][74] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][74] ), .Q(\mem_r[7][74] ), .QN( ));
Q_FDP1 \mem_r_REG[7][75] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][75] ), .Q(\mem_r[7][75] ), .QN( ));
Q_FDP1 \mem_r_REG[7][76] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][76] ), .Q(\mem_r[7][76] ), .QN( ));
Q_FDP1 \mem_r_REG[7][77] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][77] ), .Q(\mem_r[7][77] ), .QN( ));
Q_FDP1 \mem_r_REG[7][78] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][78] ), .Q(\mem_r[7][78] ), .QN( ));
Q_FDP1 \mem_r_REG[7][79] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][79] ), .Q(\mem_r[7][79] ), .QN( ));
Q_FDP1 \mem_r_REG[7][80] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][80] ), .Q(\mem_r[7][80] ), .QN( ));
Q_FDP1 \mem_r_REG[7][81] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][81] ), .Q(\mem_r[7][81] ), .QN( ));
Q_FDP1 \mem_r_REG[7][82] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][82] ), .Q(\mem_r[7][82] ), .QN( ));
Q_FDP1 \mem_r_REG[7][83] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][83] ), .Q(\mem_r[7][83] ), .QN( ));
Q_FDP1 \mem_r_REG[7][84] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][84] ), .Q(\mem_r[7][84] ), .QN( ));
Q_FDP1 \mem_r_REG[7][85] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][85] ), .Q(\mem_r[7][85] ), .QN( ));
Q_FDP1 \mem_r_REG[7][86] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][86] ), .Q(\mem_r[7][86] ), .QN( ));
Q_FDP1 \mem_r_REG[7][87] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][87] ), .Q(\mem_r[7][87] ), .QN( ));
Q_FDP1 \mem_r_REG[7][88] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][88] ), .Q(\mem_r[7][88] ), .QN( ));
Q_FDP1 \mem_r_REG[7][89] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][89] ), .Q(\mem_r[7][89] ), .QN( ));
Q_FDP1 \mem_r_REG[7][90] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][90] ), .Q(\mem_r[7][90] ), .QN( ));
Q_FDP1 \mem_r_REG[7][91] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][91] ), .Q(\mem_r[7][91] ), .QN( ));
Q_FDP1 \mem_r_REG[7][92] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][92] ), .Q(\mem_r[7][92] ), .QN( ));
Q_FDP1 \mem_r_REG[7][93] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][93] ), .Q(\mem_r[7][93] ), .QN( ));
Q_FDP1 \mem_r_REG[7][94] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][94] ), .Q(\mem_r[7][94] ), .QN( ));
Q_FDP1 \mem_r_REG[7][95] ( .CK(clk), .R(rst_n), .D(\mem_nxt[7][95] ), .Q(\mem_r[7][95] ), .QN( ));
Q_FDP1 \mem_r_REG[6][0] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][0] ), .Q(\mem_r[6][0] ), .QN( ));
Q_FDP1 \mem_r_REG[6][1] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][1] ), .Q(\mem_r[6][1] ), .QN( ));
Q_FDP1 \mem_r_REG[6][2] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][2] ), .Q(\mem_r[6][2] ), .QN( ));
Q_FDP1 \mem_r_REG[6][3] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][3] ), .Q(\mem_r[6][3] ), .QN( ));
Q_FDP1 \mem_r_REG[6][4] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][4] ), .Q(\mem_r[6][4] ), .QN( ));
Q_FDP1 \mem_r_REG[6][5] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][5] ), .Q(\mem_r[6][5] ), .QN( ));
Q_FDP1 \mem_r_REG[6][6] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][6] ), .Q(\mem_r[6][6] ), .QN( ));
Q_FDP1 \mem_r_REG[6][7] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][7] ), .Q(\mem_r[6][7] ), .QN( ));
Q_FDP1 \mem_r_REG[6][8] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][8] ), .Q(\mem_r[6][8] ), .QN( ));
Q_FDP1 \mem_r_REG[6][9] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][9] ), .Q(\mem_r[6][9] ), .QN( ));
Q_FDP1 \mem_r_REG[6][10] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][10] ), .Q(\mem_r[6][10] ), .QN( ));
Q_FDP1 \mem_r_REG[6][11] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][11] ), .Q(\mem_r[6][11] ), .QN( ));
Q_FDP1 \mem_r_REG[6][12] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][12] ), .Q(\mem_r[6][12] ), .QN( ));
Q_FDP1 \mem_r_REG[6][13] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][13] ), .Q(\mem_r[6][13] ), .QN( ));
Q_FDP1 \mem_r_REG[6][14] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][14] ), .Q(\mem_r[6][14] ), .QN( ));
Q_FDP1 \mem_r_REG[6][15] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][15] ), .Q(\mem_r[6][15] ), .QN( ));
Q_FDP1 \mem_r_REG[6][16] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][16] ), .Q(\mem_r[6][16] ), .QN( ));
Q_FDP1 \mem_r_REG[6][17] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][17] ), .Q(\mem_r[6][17] ), .QN( ));
Q_FDP1 \mem_r_REG[6][18] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][18] ), .Q(\mem_r[6][18] ), .QN( ));
Q_FDP1 \mem_r_REG[6][19] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][19] ), .Q(\mem_r[6][19] ), .QN( ));
Q_FDP1 \mem_r_REG[6][20] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][20] ), .Q(\mem_r[6][20] ), .QN( ));
Q_FDP1 \mem_r_REG[6][21] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][21] ), .Q(\mem_r[6][21] ), .QN( ));
Q_FDP1 \mem_r_REG[6][22] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][22] ), .Q(\mem_r[6][22] ), .QN( ));
Q_FDP1 \mem_r_REG[6][23] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][23] ), .Q(\mem_r[6][23] ), .QN( ));
Q_FDP1 \mem_r_REG[6][24] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][24] ), .Q(\mem_r[6][24] ), .QN( ));
Q_FDP1 \mem_r_REG[6][25] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][25] ), .Q(\mem_r[6][25] ), .QN( ));
Q_FDP1 \mem_r_REG[6][26] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][26] ), .Q(\mem_r[6][26] ), .QN( ));
Q_FDP1 \mem_r_REG[6][27] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][27] ), .Q(\mem_r[6][27] ), .QN( ));
Q_FDP1 \mem_r_REG[6][28] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][28] ), .Q(\mem_r[6][28] ), .QN( ));
Q_FDP1 \mem_r_REG[6][29] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][29] ), .Q(\mem_r[6][29] ), .QN( ));
Q_FDP1 \mem_r_REG[6][30] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][30] ), .Q(\mem_r[6][30] ), .QN( ));
Q_FDP1 \mem_r_REG[6][31] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][31] ), .Q(\mem_r[6][31] ), .QN( ));
Q_FDP1 \mem_r_REG[6][32] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][32] ), .Q(\mem_r[6][32] ), .QN( ));
Q_FDP1 \mem_r_REG[6][33] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][33] ), .Q(\mem_r[6][33] ), .QN( ));
Q_FDP1 \mem_r_REG[6][34] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][34] ), .Q(\mem_r[6][34] ), .QN( ));
Q_FDP1 \mem_r_REG[6][35] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][35] ), .Q(\mem_r[6][35] ), .QN( ));
Q_FDP1 \mem_r_REG[6][36] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][36] ), .Q(\mem_r[6][36] ), .QN( ));
Q_FDP1 \mem_r_REG[6][37] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][37] ), .Q(\mem_r[6][37] ), .QN( ));
Q_FDP1 \mem_r_REG[6][38] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][38] ), .Q(\mem_r[6][38] ), .QN( ));
Q_FDP1 \mem_r_REG[6][39] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][39] ), .Q(\mem_r[6][39] ), .QN( ));
Q_FDP1 \mem_r_REG[6][40] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][40] ), .Q(\mem_r[6][40] ), .QN( ));
Q_FDP1 \mem_r_REG[6][41] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][41] ), .Q(\mem_r[6][41] ), .QN( ));
Q_FDP1 \mem_r_REG[6][42] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][42] ), .Q(\mem_r[6][42] ), .QN( ));
Q_FDP1 \mem_r_REG[6][43] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][43] ), .Q(\mem_r[6][43] ), .QN( ));
Q_FDP1 \mem_r_REG[6][44] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][44] ), .Q(\mem_r[6][44] ), .QN( ));
Q_FDP1 \mem_r_REG[6][45] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][45] ), .Q(\mem_r[6][45] ), .QN( ));
Q_FDP1 \mem_r_REG[6][46] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][46] ), .Q(\mem_r[6][46] ), .QN( ));
Q_FDP1 \mem_r_REG[6][47] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][47] ), .Q(\mem_r[6][47] ), .QN( ));
Q_FDP1 \mem_r_REG[6][48] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][48] ), .Q(\mem_r[6][48] ), .QN( ));
Q_FDP1 \mem_r_REG[6][49] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][49] ), .Q(\mem_r[6][49] ), .QN( ));
Q_FDP1 \mem_r_REG[6][50] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][50] ), .Q(\mem_r[6][50] ), .QN( ));
Q_FDP1 \mem_r_REG[6][51] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][51] ), .Q(\mem_r[6][51] ), .QN( ));
Q_FDP1 \mem_r_REG[6][52] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][52] ), .Q(\mem_r[6][52] ), .QN( ));
Q_FDP1 \mem_r_REG[6][53] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][53] ), .Q(\mem_r[6][53] ), .QN( ));
Q_FDP1 \mem_r_REG[6][54] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][54] ), .Q(\mem_r[6][54] ), .QN( ));
Q_FDP1 \mem_r_REG[6][55] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][55] ), .Q(\mem_r[6][55] ), .QN( ));
Q_FDP1 \mem_r_REG[6][56] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][56] ), .Q(\mem_r[6][56] ), .QN( ));
Q_FDP1 \mem_r_REG[6][57] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][57] ), .Q(\mem_r[6][57] ), .QN( ));
Q_FDP1 \mem_r_REG[6][58] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][58] ), .Q(\mem_r[6][58] ), .QN( ));
Q_FDP1 \mem_r_REG[6][59] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][59] ), .Q(\mem_r[6][59] ), .QN( ));
Q_FDP1 \mem_r_REG[6][60] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][60] ), .Q(\mem_r[6][60] ), .QN( ));
Q_FDP1 \mem_r_REG[6][61] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][61] ), .Q(\mem_r[6][61] ), .QN( ));
Q_FDP1 \mem_r_REG[6][62] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][62] ), .Q(\mem_r[6][62] ), .QN( ));
Q_FDP1 \mem_r_REG[6][63] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][63] ), .Q(\mem_r[6][63] ), .QN( ));
Q_FDP1 \mem_r_REG[6][64] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][64] ), .Q(\mem_r[6][64] ), .QN( ));
Q_FDP1 \mem_r_REG[6][65] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][65] ), .Q(\mem_r[6][65] ), .QN( ));
Q_FDP1 \mem_r_REG[6][66] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][66] ), .Q(\mem_r[6][66] ), .QN( ));
Q_FDP1 \mem_r_REG[6][67] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][67] ), .Q(\mem_r[6][67] ), .QN( ));
Q_FDP1 \mem_r_REG[6][68] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][68] ), .Q(\mem_r[6][68] ), .QN( ));
Q_FDP1 \mem_r_REG[6][69] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][69] ), .Q(\mem_r[6][69] ), .QN( ));
Q_FDP1 \mem_r_REG[6][70] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][70] ), .Q(\mem_r[6][70] ), .QN( ));
Q_FDP1 \mem_r_REG[6][71] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][71] ), .Q(\mem_r[6][71] ), .QN( ));
Q_FDP1 \mem_r_REG[6][72] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][72] ), .Q(\mem_r[6][72] ), .QN( ));
Q_FDP1 \mem_r_REG[6][73] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][73] ), .Q(\mem_r[6][73] ), .QN( ));
Q_FDP1 \mem_r_REG[6][74] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][74] ), .Q(\mem_r[6][74] ), .QN( ));
Q_FDP1 \mem_r_REG[6][75] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][75] ), .Q(\mem_r[6][75] ), .QN( ));
Q_FDP1 \mem_r_REG[6][76] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][76] ), .Q(\mem_r[6][76] ), .QN( ));
Q_FDP1 \mem_r_REG[6][77] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][77] ), .Q(\mem_r[6][77] ), .QN( ));
Q_FDP1 \mem_r_REG[6][78] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][78] ), .Q(\mem_r[6][78] ), .QN( ));
Q_FDP1 \mem_r_REG[6][79] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][79] ), .Q(\mem_r[6][79] ), .QN( ));
Q_FDP1 \mem_r_REG[6][80] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][80] ), .Q(\mem_r[6][80] ), .QN( ));
Q_FDP1 \mem_r_REG[6][81] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][81] ), .Q(\mem_r[6][81] ), .QN( ));
Q_FDP1 \mem_r_REG[6][82] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][82] ), .Q(\mem_r[6][82] ), .QN( ));
Q_FDP1 \mem_r_REG[6][83] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][83] ), .Q(\mem_r[6][83] ), .QN( ));
Q_FDP1 \mem_r_REG[6][84] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][84] ), .Q(\mem_r[6][84] ), .QN( ));
Q_FDP1 \mem_r_REG[6][85] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][85] ), .Q(\mem_r[6][85] ), .QN( ));
Q_FDP1 \mem_r_REG[6][86] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][86] ), .Q(\mem_r[6][86] ), .QN( ));
Q_FDP1 \mem_r_REG[6][87] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][87] ), .Q(\mem_r[6][87] ), .QN( ));
Q_FDP1 \mem_r_REG[6][88] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][88] ), .Q(\mem_r[6][88] ), .QN( ));
Q_FDP1 \mem_r_REG[6][89] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][89] ), .Q(\mem_r[6][89] ), .QN( ));
Q_FDP1 \mem_r_REG[6][90] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][90] ), .Q(\mem_r[6][90] ), .QN( ));
Q_FDP1 \mem_r_REG[6][91] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][91] ), .Q(\mem_r[6][91] ), .QN( ));
Q_FDP1 \mem_r_REG[6][92] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][92] ), .Q(\mem_r[6][92] ), .QN( ));
Q_FDP1 \mem_r_REG[6][93] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][93] ), .Q(\mem_r[6][93] ), .QN( ));
Q_FDP1 \mem_r_REG[6][94] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][94] ), .Q(\mem_r[6][94] ), .QN( ));
Q_FDP1 \mem_r_REG[6][95] ( .CK(clk), .R(rst_n), .D(\mem_nxt[6][95] ), .Q(\mem_r[6][95] ), .QN( ));
Q_FDP1 \mem_r_REG[5][0] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][0] ), .Q(\mem_r[5][0] ), .QN( ));
Q_FDP1 \mem_r_REG[5][1] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][1] ), .Q(\mem_r[5][1] ), .QN( ));
Q_FDP1 \mem_r_REG[5][2] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][2] ), .Q(\mem_r[5][2] ), .QN( ));
Q_FDP1 \mem_r_REG[5][3] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][3] ), .Q(\mem_r[5][3] ), .QN( ));
Q_FDP1 \mem_r_REG[5][4] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][4] ), .Q(\mem_r[5][4] ), .QN( ));
Q_FDP1 \mem_r_REG[5][5] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][5] ), .Q(\mem_r[5][5] ), .QN( ));
Q_FDP1 \mem_r_REG[5][6] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][6] ), .Q(\mem_r[5][6] ), .QN( ));
Q_FDP1 \mem_r_REG[5][7] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][7] ), .Q(\mem_r[5][7] ), .QN( ));
Q_FDP1 \mem_r_REG[5][8] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][8] ), .Q(\mem_r[5][8] ), .QN( ));
Q_FDP1 \mem_r_REG[5][9] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][9] ), .Q(\mem_r[5][9] ), .QN( ));
Q_FDP1 \mem_r_REG[5][10] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][10] ), .Q(\mem_r[5][10] ), .QN( ));
Q_FDP1 \mem_r_REG[5][11] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][11] ), .Q(\mem_r[5][11] ), .QN( ));
Q_FDP1 \mem_r_REG[5][12] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][12] ), .Q(\mem_r[5][12] ), .QN( ));
Q_FDP1 \mem_r_REG[5][13] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][13] ), .Q(\mem_r[5][13] ), .QN( ));
Q_FDP1 \mem_r_REG[5][14] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][14] ), .Q(\mem_r[5][14] ), .QN( ));
Q_FDP1 \mem_r_REG[5][15] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][15] ), .Q(\mem_r[5][15] ), .QN( ));
Q_FDP1 \mem_r_REG[5][16] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][16] ), .Q(\mem_r[5][16] ), .QN( ));
Q_FDP1 \mem_r_REG[5][17] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][17] ), .Q(\mem_r[5][17] ), .QN( ));
Q_FDP1 \mem_r_REG[5][18] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][18] ), .Q(\mem_r[5][18] ), .QN( ));
Q_FDP1 \mem_r_REG[5][19] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][19] ), .Q(\mem_r[5][19] ), .QN( ));
Q_FDP1 \mem_r_REG[5][20] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][20] ), .Q(\mem_r[5][20] ), .QN( ));
Q_FDP1 \mem_r_REG[5][21] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][21] ), .Q(\mem_r[5][21] ), .QN( ));
Q_FDP1 \mem_r_REG[5][22] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][22] ), .Q(\mem_r[5][22] ), .QN( ));
Q_FDP1 \mem_r_REG[5][23] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][23] ), .Q(\mem_r[5][23] ), .QN( ));
Q_FDP1 \mem_r_REG[5][24] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][24] ), .Q(\mem_r[5][24] ), .QN( ));
Q_FDP1 \mem_r_REG[5][25] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][25] ), .Q(\mem_r[5][25] ), .QN( ));
Q_FDP1 \mem_r_REG[5][26] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][26] ), .Q(\mem_r[5][26] ), .QN( ));
Q_FDP1 \mem_r_REG[5][27] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][27] ), .Q(\mem_r[5][27] ), .QN( ));
Q_FDP1 \mem_r_REG[5][28] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][28] ), .Q(\mem_r[5][28] ), .QN( ));
Q_FDP1 \mem_r_REG[5][29] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][29] ), .Q(\mem_r[5][29] ), .QN( ));
Q_FDP1 \mem_r_REG[5][30] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][30] ), .Q(\mem_r[5][30] ), .QN( ));
Q_FDP1 \mem_r_REG[5][31] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][31] ), .Q(\mem_r[5][31] ), .QN( ));
Q_FDP1 \mem_r_REG[5][32] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][32] ), .Q(\mem_r[5][32] ), .QN( ));
Q_FDP1 \mem_r_REG[5][33] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][33] ), .Q(\mem_r[5][33] ), .QN( ));
Q_FDP1 \mem_r_REG[5][34] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][34] ), .Q(\mem_r[5][34] ), .QN( ));
Q_FDP1 \mem_r_REG[5][35] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][35] ), .Q(\mem_r[5][35] ), .QN( ));
Q_FDP1 \mem_r_REG[5][36] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][36] ), .Q(\mem_r[5][36] ), .QN( ));
Q_FDP1 \mem_r_REG[5][37] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][37] ), .Q(\mem_r[5][37] ), .QN( ));
Q_FDP1 \mem_r_REG[5][38] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][38] ), .Q(\mem_r[5][38] ), .QN( ));
Q_FDP1 \mem_r_REG[5][39] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][39] ), .Q(\mem_r[5][39] ), .QN( ));
Q_FDP1 \mem_r_REG[5][40] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][40] ), .Q(\mem_r[5][40] ), .QN( ));
Q_FDP1 \mem_r_REG[5][41] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][41] ), .Q(\mem_r[5][41] ), .QN( ));
Q_FDP1 \mem_r_REG[5][42] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][42] ), .Q(\mem_r[5][42] ), .QN( ));
Q_FDP1 \mem_r_REG[5][43] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][43] ), .Q(\mem_r[5][43] ), .QN( ));
Q_FDP1 \mem_r_REG[5][44] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][44] ), .Q(\mem_r[5][44] ), .QN( ));
Q_FDP1 \mem_r_REG[5][45] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][45] ), .Q(\mem_r[5][45] ), .QN( ));
Q_FDP1 \mem_r_REG[5][46] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][46] ), .Q(\mem_r[5][46] ), .QN( ));
Q_FDP1 \mem_r_REG[5][47] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][47] ), .Q(\mem_r[5][47] ), .QN( ));
Q_FDP1 \mem_r_REG[5][48] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][48] ), .Q(\mem_r[5][48] ), .QN( ));
Q_FDP1 \mem_r_REG[5][49] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][49] ), .Q(\mem_r[5][49] ), .QN( ));
Q_FDP1 \mem_r_REG[5][50] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][50] ), .Q(\mem_r[5][50] ), .QN( ));
Q_FDP1 \mem_r_REG[5][51] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][51] ), .Q(\mem_r[5][51] ), .QN( ));
Q_FDP1 \mem_r_REG[5][52] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][52] ), .Q(\mem_r[5][52] ), .QN( ));
Q_FDP1 \mem_r_REG[5][53] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][53] ), .Q(\mem_r[5][53] ), .QN( ));
Q_FDP1 \mem_r_REG[5][54] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][54] ), .Q(\mem_r[5][54] ), .QN( ));
Q_FDP1 \mem_r_REG[5][55] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][55] ), .Q(\mem_r[5][55] ), .QN( ));
Q_FDP1 \mem_r_REG[5][56] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][56] ), .Q(\mem_r[5][56] ), .QN( ));
Q_FDP1 \mem_r_REG[5][57] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][57] ), .Q(\mem_r[5][57] ), .QN( ));
Q_FDP1 \mem_r_REG[5][58] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][58] ), .Q(\mem_r[5][58] ), .QN( ));
Q_FDP1 \mem_r_REG[5][59] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][59] ), .Q(\mem_r[5][59] ), .QN( ));
Q_FDP1 \mem_r_REG[5][60] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][60] ), .Q(\mem_r[5][60] ), .QN( ));
Q_FDP1 \mem_r_REG[5][61] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][61] ), .Q(\mem_r[5][61] ), .QN( ));
Q_FDP1 \mem_r_REG[5][62] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][62] ), .Q(\mem_r[5][62] ), .QN( ));
Q_FDP1 \mem_r_REG[5][63] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][63] ), .Q(\mem_r[5][63] ), .QN( ));
Q_FDP1 \mem_r_REG[5][64] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][64] ), .Q(\mem_r[5][64] ), .QN( ));
Q_FDP1 \mem_r_REG[5][65] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][65] ), .Q(\mem_r[5][65] ), .QN( ));
Q_FDP1 \mem_r_REG[5][66] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][66] ), .Q(\mem_r[5][66] ), .QN( ));
Q_FDP1 \mem_r_REG[5][67] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][67] ), .Q(\mem_r[5][67] ), .QN( ));
Q_FDP1 \mem_r_REG[5][68] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][68] ), .Q(\mem_r[5][68] ), .QN( ));
Q_FDP1 \mem_r_REG[5][69] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][69] ), .Q(\mem_r[5][69] ), .QN( ));
Q_FDP1 \mem_r_REG[5][70] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][70] ), .Q(\mem_r[5][70] ), .QN( ));
Q_FDP1 \mem_r_REG[5][71] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][71] ), .Q(\mem_r[5][71] ), .QN( ));
Q_FDP1 \mem_r_REG[5][72] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][72] ), .Q(\mem_r[5][72] ), .QN( ));
Q_FDP1 \mem_r_REG[5][73] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][73] ), .Q(\mem_r[5][73] ), .QN( ));
Q_FDP1 \mem_r_REG[5][74] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][74] ), .Q(\mem_r[5][74] ), .QN( ));
Q_FDP1 \mem_r_REG[5][75] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][75] ), .Q(\mem_r[5][75] ), .QN( ));
Q_FDP1 \mem_r_REG[5][76] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][76] ), .Q(\mem_r[5][76] ), .QN( ));
Q_FDP1 \mem_r_REG[5][77] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][77] ), .Q(\mem_r[5][77] ), .QN( ));
Q_FDP1 \mem_r_REG[5][78] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][78] ), .Q(\mem_r[5][78] ), .QN( ));
Q_FDP1 \mem_r_REG[5][79] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][79] ), .Q(\mem_r[5][79] ), .QN( ));
Q_FDP1 \mem_r_REG[5][80] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][80] ), .Q(\mem_r[5][80] ), .QN( ));
Q_FDP1 \mem_r_REG[5][81] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][81] ), .Q(\mem_r[5][81] ), .QN( ));
Q_FDP1 \mem_r_REG[5][82] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][82] ), .Q(\mem_r[5][82] ), .QN( ));
Q_FDP1 \mem_r_REG[5][83] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][83] ), .Q(\mem_r[5][83] ), .QN( ));
Q_FDP1 \mem_r_REG[5][84] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][84] ), .Q(\mem_r[5][84] ), .QN( ));
Q_FDP1 \mem_r_REG[5][85] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][85] ), .Q(\mem_r[5][85] ), .QN( ));
Q_FDP1 \mem_r_REG[5][86] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][86] ), .Q(\mem_r[5][86] ), .QN( ));
Q_FDP1 \mem_r_REG[5][87] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][87] ), .Q(\mem_r[5][87] ), .QN( ));
Q_FDP1 \mem_r_REG[5][88] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][88] ), .Q(\mem_r[5][88] ), .QN( ));
Q_FDP1 \mem_r_REG[5][89] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][89] ), .Q(\mem_r[5][89] ), .QN( ));
Q_FDP1 \mem_r_REG[5][90] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][90] ), .Q(\mem_r[5][90] ), .QN( ));
Q_FDP1 \mem_r_REG[5][91] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][91] ), .Q(\mem_r[5][91] ), .QN( ));
Q_FDP1 \mem_r_REG[5][92] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][92] ), .Q(\mem_r[5][92] ), .QN( ));
Q_FDP1 \mem_r_REG[5][93] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][93] ), .Q(\mem_r[5][93] ), .QN( ));
Q_FDP1 \mem_r_REG[5][94] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][94] ), .Q(\mem_r[5][94] ), .QN( ));
Q_FDP1 \mem_r_REG[5][95] ( .CK(clk), .R(rst_n), .D(\mem_nxt[5][95] ), .Q(\mem_r[5][95] ), .QN( ));
Q_FDP1 \mem_r_REG[4][0] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][0] ), .Q(\mem_r[4][0] ), .QN( ));
Q_FDP1 \mem_r_REG[4][1] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][1] ), .Q(\mem_r[4][1] ), .QN( ));
Q_FDP1 \mem_r_REG[4][2] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][2] ), .Q(\mem_r[4][2] ), .QN( ));
Q_FDP1 \mem_r_REG[4][3] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][3] ), .Q(\mem_r[4][3] ), .QN( ));
Q_FDP1 \mem_r_REG[4][4] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][4] ), .Q(\mem_r[4][4] ), .QN( ));
Q_FDP1 \mem_r_REG[4][5] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][5] ), .Q(\mem_r[4][5] ), .QN( ));
Q_FDP1 \mem_r_REG[4][6] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][6] ), .Q(\mem_r[4][6] ), .QN( ));
Q_FDP1 \mem_r_REG[4][7] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][7] ), .Q(\mem_r[4][7] ), .QN( ));
Q_FDP1 \mem_r_REG[4][8] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][8] ), .Q(\mem_r[4][8] ), .QN( ));
Q_FDP1 \mem_r_REG[4][9] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][9] ), .Q(\mem_r[4][9] ), .QN( ));
Q_FDP1 \mem_r_REG[4][10] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][10] ), .Q(\mem_r[4][10] ), .QN( ));
Q_FDP1 \mem_r_REG[4][11] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][11] ), .Q(\mem_r[4][11] ), .QN( ));
Q_FDP1 \mem_r_REG[4][12] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][12] ), .Q(\mem_r[4][12] ), .QN( ));
Q_FDP1 \mem_r_REG[4][13] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][13] ), .Q(\mem_r[4][13] ), .QN( ));
Q_FDP1 \mem_r_REG[4][14] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][14] ), .Q(\mem_r[4][14] ), .QN( ));
Q_FDP1 \mem_r_REG[4][15] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][15] ), .Q(\mem_r[4][15] ), .QN( ));
Q_FDP1 \mem_r_REG[4][16] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][16] ), .Q(\mem_r[4][16] ), .QN( ));
Q_FDP1 \mem_r_REG[4][17] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][17] ), .Q(\mem_r[4][17] ), .QN( ));
Q_FDP1 \mem_r_REG[4][18] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][18] ), .Q(\mem_r[4][18] ), .QN( ));
Q_FDP1 \mem_r_REG[4][19] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][19] ), .Q(\mem_r[4][19] ), .QN( ));
Q_FDP1 \mem_r_REG[4][20] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][20] ), .Q(\mem_r[4][20] ), .QN( ));
Q_FDP1 \mem_r_REG[4][21] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][21] ), .Q(\mem_r[4][21] ), .QN( ));
Q_FDP1 \mem_r_REG[4][22] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][22] ), .Q(\mem_r[4][22] ), .QN( ));
Q_FDP1 \mem_r_REG[4][23] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][23] ), .Q(\mem_r[4][23] ), .QN( ));
Q_FDP1 \mem_r_REG[4][24] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][24] ), .Q(\mem_r[4][24] ), .QN( ));
Q_FDP1 \mem_r_REG[4][25] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][25] ), .Q(\mem_r[4][25] ), .QN( ));
Q_FDP1 \mem_r_REG[4][26] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][26] ), .Q(\mem_r[4][26] ), .QN( ));
Q_FDP1 \mem_r_REG[4][27] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][27] ), .Q(\mem_r[4][27] ), .QN( ));
Q_FDP1 \mem_r_REG[4][28] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][28] ), .Q(\mem_r[4][28] ), .QN( ));
Q_FDP1 \mem_r_REG[4][29] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][29] ), .Q(\mem_r[4][29] ), .QN( ));
Q_FDP1 \mem_r_REG[4][30] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][30] ), .Q(\mem_r[4][30] ), .QN( ));
Q_FDP1 \mem_r_REG[4][31] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][31] ), .Q(\mem_r[4][31] ), .QN( ));
Q_FDP1 \mem_r_REG[4][32] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][32] ), .Q(\mem_r[4][32] ), .QN( ));
Q_FDP1 \mem_r_REG[4][33] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][33] ), .Q(\mem_r[4][33] ), .QN( ));
Q_FDP1 \mem_r_REG[4][34] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][34] ), .Q(\mem_r[4][34] ), .QN( ));
Q_FDP1 \mem_r_REG[4][35] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][35] ), .Q(\mem_r[4][35] ), .QN( ));
Q_FDP1 \mem_r_REG[4][36] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][36] ), .Q(\mem_r[4][36] ), .QN( ));
Q_FDP1 \mem_r_REG[4][37] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][37] ), .Q(\mem_r[4][37] ), .QN( ));
Q_FDP1 \mem_r_REG[4][38] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][38] ), .Q(\mem_r[4][38] ), .QN( ));
Q_FDP1 \mem_r_REG[4][39] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][39] ), .Q(\mem_r[4][39] ), .QN( ));
Q_FDP1 \mem_r_REG[4][40] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][40] ), .Q(\mem_r[4][40] ), .QN( ));
Q_FDP1 \mem_r_REG[4][41] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][41] ), .Q(\mem_r[4][41] ), .QN( ));
Q_FDP1 \mem_r_REG[4][42] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][42] ), .Q(\mem_r[4][42] ), .QN( ));
Q_FDP1 \mem_r_REG[4][43] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][43] ), .Q(\mem_r[4][43] ), .QN( ));
Q_FDP1 \mem_r_REG[4][44] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][44] ), .Q(\mem_r[4][44] ), .QN( ));
Q_FDP1 \mem_r_REG[4][45] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][45] ), .Q(\mem_r[4][45] ), .QN( ));
Q_FDP1 \mem_r_REG[4][46] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][46] ), .Q(\mem_r[4][46] ), .QN( ));
Q_FDP1 \mem_r_REG[4][47] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][47] ), .Q(\mem_r[4][47] ), .QN( ));
Q_FDP1 \mem_r_REG[4][48] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][48] ), .Q(\mem_r[4][48] ), .QN( ));
Q_FDP1 \mem_r_REG[4][49] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][49] ), .Q(\mem_r[4][49] ), .QN( ));
Q_FDP1 \mem_r_REG[4][50] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][50] ), .Q(\mem_r[4][50] ), .QN( ));
Q_FDP1 \mem_r_REG[4][51] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][51] ), .Q(\mem_r[4][51] ), .QN( ));
Q_FDP1 \mem_r_REG[4][52] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][52] ), .Q(\mem_r[4][52] ), .QN( ));
Q_FDP1 \mem_r_REG[4][53] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][53] ), .Q(\mem_r[4][53] ), .QN( ));
Q_FDP1 \mem_r_REG[4][54] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][54] ), .Q(\mem_r[4][54] ), .QN( ));
Q_FDP1 \mem_r_REG[4][55] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][55] ), .Q(\mem_r[4][55] ), .QN( ));
Q_FDP1 \mem_r_REG[4][56] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][56] ), .Q(\mem_r[4][56] ), .QN( ));
Q_FDP1 \mem_r_REG[4][57] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][57] ), .Q(\mem_r[4][57] ), .QN( ));
Q_FDP1 \mem_r_REG[4][58] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][58] ), .Q(\mem_r[4][58] ), .QN( ));
Q_FDP1 \mem_r_REG[4][59] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][59] ), .Q(\mem_r[4][59] ), .QN( ));
Q_FDP1 \mem_r_REG[4][60] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][60] ), .Q(\mem_r[4][60] ), .QN( ));
Q_FDP1 \mem_r_REG[4][61] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][61] ), .Q(\mem_r[4][61] ), .QN( ));
Q_FDP1 \mem_r_REG[4][62] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][62] ), .Q(\mem_r[4][62] ), .QN( ));
Q_FDP1 \mem_r_REG[4][63] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][63] ), .Q(\mem_r[4][63] ), .QN( ));
Q_FDP1 \mem_r_REG[4][64] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][64] ), .Q(\mem_r[4][64] ), .QN( ));
Q_FDP1 \mem_r_REG[4][65] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][65] ), .Q(\mem_r[4][65] ), .QN( ));
Q_FDP1 \mem_r_REG[4][66] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][66] ), .Q(\mem_r[4][66] ), .QN( ));
Q_FDP1 \mem_r_REG[4][67] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][67] ), .Q(\mem_r[4][67] ), .QN( ));
Q_FDP1 \mem_r_REG[4][68] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][68] ), .Q(\mem_r[4][68] ), .QN( ));
Q_FDP1 \mem_r_REG[4][69] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][69] ), .Q(\mem_r[4][69] ), .QN( ));
Q_FDP1 \mem_r_REG[4][70] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][70] ), .Q(\mem_r[4][70] ), .QN( ));
Q_FDP1 \mem_r_REG[4][71] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][71] ), .Q(\mem_r[4][71] ), .QN( ));
Q_FDP1 \mem_r_REG[4][72] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][72] ), .Q(\mem_r[4][72] ), .QN( ));
Q_FDP1 \mem_r_REG[4][73] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][73] ), .Q(\mem_r[4][73] ), .QN( ));
Q_FDP1 \mem_r_REG[4][74] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][74] ), .Q(\mem_r[4][74] ), .QN( ));
Q_FDP1 \mem_r_REG[4][75] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][75] ), .Q(\mem_r[4][75] ), .QN( ));
Q_FDP1 \mem_r_REG[4][76] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][76] ), .Q(\mem_r[4][76] ), .QN( ));
Q_FDP1 \mem_r_REG[4][77] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][77] ), .Q(\mem_r[4][77] ), .QN( ));
Q_FDP1 \mem_r_REG[4][78] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][78] ), .Q(\mem_r[4][78] ), .QN( ));
Q_FDP1 \mem_r_REG[4][79] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][79] ), .Q(\mem_r[4][79] ), .QN( ));
Q_FDP1 \mem_r_REG[4][80] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][80] ), .Q(\mem_r[4][80] ), .QN( ));
Q_FDP1 \mem_r_REG[4][81] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][81] ), .Q(\mem_r[4][81] ), .QN( ));
Q_FDP1 \mem_r_REG[4][82] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][82] ), .Q(\mem_r[4][82] ), .QN( ));
Q_FDP1 \mem_r_REG[4][83] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][83] ), .Q(\mem_r[4][83] ), .QN( ));
Q_FDP1 \mem_r_REG[4][84] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][84] ), .Q(\mem_r[4][84] ), .QN( ));
Q_FDP1 \mem_r_REG[4][85] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][85] ), .Q(\mem_r[4][85] ), .QN( ));
Q_FDP1 \mem_r_REG[4][86] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][86] ), .Q(\mem_r[4][86] ), .QN( ));
Q_FDP1 \mem_r_REG[4][87] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][87] ), .Q(\mem_r[4][87] ), .QN( ));
Q_FDP1 \mem_r_REG[4][88] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][88] ), .Q(\mem_r[4][88] ), .QN( ));
Q_FDP1 \mem_r_REG[4][89] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][89] ), .Q(\mem_r[4][89] ), .QN( ));
Q_FDP1 \mem_r_REG[4][90] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][90] ), .Q(\mem_r[4][90] ), .QN( ));
Q_FDP1 \mem_r_REG[4][91] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][91] ), .Q(\mem_r[4][91] ), .QN( ));
Q_FDP1 \mem_r_REG[4][92] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][92] ), .Q(\mem_r[4][92] ), .QN( ));
Q_FDP1 \mem_r_REG[4][93] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][93] ), .Q(\mem_r[4][93] ), .QN( ));
Q_FDP1 \mem_r_REG[4][94] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][94] ), .Q(\mem_r[4][94] ), .QN( ));
Q_FDP1 \mem_r_REG[4][95] ( .CK(clk), .R(rst_n), .D(\mem_nxt[4][95] ), .Q(\mem_r[4][95] ), .QN( ));
Q_FDP1 \mem_r_REG[3][0] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][0] ), .Q(\mem_r[3][0] ), .QN( ));
Q_FDP1 \mem_r_REG[3][1] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][1] ), .Q(\mem_r[3][1] ), .QN( ));
Q_FDP1 \mem_r_REG[3][2] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][2] ), .Q(\mem_r[3][2] ), .QN( ));
Q_FDP1 \mem_r_REG[3][3] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][3] ), .Q(\mem_r[3][3] ), .QN( ));
Q_FDP1 \mem_r_REG[3][4] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][4] ), .Q(\mem_r[3][4] ), .QN( ));
Q_FDP1 \mem_r_REG[3][5] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][5] ), .Q(\mem_r[3][5] ), .QN( ));
Q_FDP1 \mem_r_REG[3][6] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][6] ), .Q(\mem_r[3][6] ), .QN( ));
Q_FDP1 \mem_r_REG[3][7] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][7] ), .Q(\mem_r[3][7] ), .QN( ));
Q_FDP1 \mem_r_REG[3][8] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][8] ), .Q(\mem_r[3][8] ), .QN( ));
Q_FDP1 \mem_r_REG[3][9] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][9] ), .Q(\mem_r[3][9] ), .QN( ));
Q_FDP1 \mem_r_REG[3][10] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][10] ), .Q(\mem_r[3][10] ), .QN( ));
Q_FDP1 \mem_r_REG[3][11] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][11] ), .Q(\mem_r[3][11] ), .QN( ));
Q_FDP1 \mem_r_REG[3][12] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][12] ), .Q(\mem_r[3][12] ), .QN( ));
Q_FDP1 \mem_r_REG[3][13] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][13] ), .Q(\mem_r[3][13] ), .QN( ));
Q_FDP1 \mem_r_REG[3][14] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][14] ), .Q(\mem_r[3][14] ), .QN( ));
Q_FDP1 \mem_r_REG[3][15] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][15] ), .Q(\mem_r[3][15] ), .QN( ));
Q_FDP1 \mem_r_REG[3][16] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][16] ), .Q(\mem_r[3][16] ), .QN( ));
Q_FDP1 \mem_r_REG[3][17] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][17] ), .Q(\mem_r[3][17] ), .QN( ));
Q_FDP1 \mem_r_REG[3][18] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][18] ), .Q(\mem_r[3][18] ), .QN( ));
Q_FDP1 \mem_r_REG[3][19] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][19] ), .Q(\mem_r[3][19] ), .QN( ));
Q_FDP1 \mem_r_REG[3][20] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][20] ), .Q(\mem_r[3][20] ), .QN( ));
Q_FDP1 \mem_r_REG[3][21] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][21] ), .Q(\mem_r[3][21] ), .QN( ));
Q_FDP1 \mem_r_REG[3][22] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][22] ), .Q(\mem_r[3][22] ), .QN( ));
Q_FDP1 \mem_r_REG[3][23] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][23] ), .Q(\mem_r[3][23] ), .QN( ));
Q_FDP1 \mem_r_REG[3][24] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][24] ), .Q(\mem_r[3][24] ), .QN( ));
Q_FDP1 \mem_r_REG[3][25] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][25] ), .Q(\mem_r[3][25] ), .QN( ));
Q_FDP1 \mem_r_REG[3][26] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][26] ), .Q(\mem_r[3][26] ), .QN( ));
Q_FDP1 \mem_r_REG[3][27] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][27] ), .Q(\mem_r[3][27] ), .QN( ));
Q_FDP1 \mem_r_REG[3][28] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][28] ), .Q(\mem_r[3][28] ), .QN( ));
Q_FDP1 \mem_r_REG[3][29] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][29] ), .Q(\mem_r[3][29] ), .QN( ));
Q_FDP1 \mem_r_REG[3][30] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][30] ), .Q(\mem_r[3][30] ), .QN( ));
Q_FDP1 \mem_r_REG[3][31] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][31] ), .Q(\mem_r[3][31] ), .QN( ));
Q_FDP1 \mem_r_REG[3][32] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][32] ), .Q(\mem_r[3][32] ), .QN( ));
Q_FDP1 \mem_r_REG[3][33] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][33] ), .Q(\mem_r[3][33] ), .QN( ));
Q_FDP1 \mem_r_REG[3][34] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][34] ), .Q(\mem_r[3][34] ), .QN( ));
Q_FDP1 \mem_r_REG[3][35] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][35] ), .Q(\mem_r[3][35] ), .QN( ));
Q_FDP1 \mem_r_REG[3][36] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][36] ), .Q(\mem_r[3][36] ), .QN( ));
Q_FDP1 \mem_r_REG[3][37] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][37] ), .Q(\mem_r[3][37] ), .QN( ));
Q_FDP1 \mem_r_REG[3][38] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][38] ), .Q(\mem_r[3][38] ), .QN( ));
Q_FDP1 \mem_r_REG[3][39] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][39] ), .Q(\mem_r[3][39] ), .QN( ));
Q_FDP1 \mem_r_REG[3][40] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][40] ), .Q(\mem_r[3][40] ), .QN( ));
Q_FDP1 \mem_r_REG[3][41] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][41] ), .Q(\mem_r[3][41] ), .QN( ));
Q_FDP1 \mem_r_REG[3][42] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][42] ), .Q(\mem_r[3][42] ), .QN( ));
Q_FDP1 \mem_r_REG[3][43] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][43] ), .Q(\mem_r[3][43] ), .QN( ));
Q_FDP1 \mem_r_REG[3][44] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][44] ), .Q(\mem_r[3][44] ), .QN( ));
Q_FDP1 \mem_r_REG[3][45] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][45] ), .Q(\mem_r[3][45] ), .QN( ));
Q_FDP1 \mem_r_REG[3][46] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][46] ), .Q(\mem_r[3][46] ), .QN( ));
Q_FDP1 \mem_r_REG[3][47] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][47] ), .Q(\mem_r[3][47] ), .QN( ));
Q_FDP1 \mem_r_REG[3][48] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][48] ), .Q(\mem_r[3][48] ), .QN( ));
Q_FDP1 \mem_r_REG[3][49] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][49] ), .Q(\mem_r[3][49] ), .QN( ));
Q_FDP1 \mem_r_REG[3][50] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][50] ), .Q(\mem_r[3][50] ), .QN( ));
Q_FDP1 \mem_r_REG[3][51] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][51] ), .Q(\mem_r[3][51] ), .QN( ));
Q_FDP1 \mem_r_REG[3][52] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][52] ), .Q(\mem_r[3][52] ), .QN( ));
Q_FDP1 \mem_r_REG[3][53] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][53] ), .Q(\mem_r[3][53] ), .QN( ));
Q_FDP1 \mem_r_REG[3][54] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][54] ), .Q(\mem_r[3][54] ), .QN( ));
Q_FDP1 \mem_r_REG[3][55] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][55] ), .Q(\mem_r[3][55] ), .QN( ));
Q_FDP1 \mem_r_REG[3][56] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][56] ), .Q(\mem_r[3][56] ), .QN( ));
Q_FDP1 \mem_r_REG[3][57] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][57] ), .Q(\mem_r[3][57] ), .QN( ));
Q_FDP1 \mem_r_REG[3][58] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][58] ), .Q(\mem_r[3][58] ), .QN( ));
Q_FDP1 \mem_r_REG[3][59] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][59] ), .Q(\mem_r[3][59] ), .QN( ));
Q_FDP1 \mem_r_REG[3][60] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][60] ), .Q(\mem_r[3][60] ), .QN( ));
Q_FDP1 \mem_r_REG[3][61] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][61] ), .Q(\mem_r[3][61] ), .QN( ));
Q_FDP1 \mem_r_REG[3][62] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][62] ), .Q(\mem_r[3][62] ), .QN( ));
Q_FDP1 \mem_r_REG[3][63] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][63] ), .Q(\mem_r[3][63] ), .QN( ));
Q_FDP1 \mem_r_REG[3][64] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][64] ), .Q(\mem_r[3][64] ), .QN( ));
Q_FDP1 \mem_r_REG[3][65] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][65] ), .Q(\mem_r[3][65] ), .QN( ));
Q_FDP1 \mem_r_REG[3][66] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][66] ), .Q(\mem_r[3][66] ), .QN( ));
Q_FDP1 \mem_r_REG[3][67] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][67] ), .Q(\mem_r[3][67] ), .QN( ));
Q_FDP1 \mem_r_REG[3][68] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][68] ), .Q(\mem_r[3][68] ), .QN( ));
Q_FDP1 \mem_r_REG[3][69] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][69] ), .Q(\mem_r[3][69] ), .QN( ));
Q_FDP1 \mem_r_REG[3][70] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][70] ), .Q(\mem_r[3][70] ), .QN( ));
Q_FDP1 \mem_r_REG[3][71] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][71] ), .Q(\mem_r[3][71] ), .QN( ));
Q_FDP1 \mem_r_REG[3][72] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][72] ), .Q(\mem_r[3][72] ), .QN( ));
Q_FDP1 \mem_r_REG[3][73] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][73] ), .Q(\mem_r[3][73] ), .QN( ));
Q_FDP1 \mem_r_REG[3][74] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][74] ), .Q(\mem_r[3][74] ), .QN( ));
Q_FDP1 \mem_r_REG[3][75] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][75] ), .Q(\mem_r[3][75] ), .QN( ));
Q_FDP1 \mem_r_REG[3][76] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][76] ), .Q(\mem_r[3][76] ), .QN( ));
Q_FDP1 \mem_r_REG[3][77] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][77] ), .Q(\mem_r[3][77] ), .QN( ));
Q_FDP1 \mem_r_REG[3][78] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][78] ), .Q(\mem_r[3][78] ), .QN( ));
Q_FDP1 \mem_r_REG[3][79] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][79] ), .Q(\mem_r[3][79] ), .QN( ));
Q_FDP1 \mem_r_REG[3][80] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][80] ), .Q(\mem_r[3][80] ), .QN( ));
Q_FDP1 \mem_r_REG[3][81] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][81] ), .Q(\mem_r[3][81] ), .QN( ));
Q_FDP1 \mem_r_REG[3][82] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][82] ), .Q(\mem_r[3][82] ), .QN( ));
Q_FDP1 \mem_r_REG[3][83] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][83] ), .Q(\mem_r[3][83] ), .QN( ));
Q_FDP1 \mem_r_REG[3][84] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][84] ), .Q(\mem_r[3][84] ), .QN( ));
Q_FDP1 \mem_r_REG[3][85] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][85] ), .Q(\mem_r[3][85] ), .QN( ));
Q_FDP1 \mem_r_REG[3][86] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][86] ), .Q(\mem_r[3][86] ), .QN( ));
Q_FDP1 \mem_r_REG[3][87] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][87] ), .Q(\mem_r[3][87] ), .QN( ));
Q_FDP1 \mem_r_REG[3][88] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][88] ), .Q(\mem_r[3][88] ), .QN( ));
Q_FDP1 \mem_r_REG[3][89] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][89] ), .Q(\mem_r[3][89] ), .QN( ));
Q_FDP1 \mem_r_REG[3][90] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][90] ), .Q(\mem_r[3][90] ), .QN( ));
Q_FDP1 \mem_r_REG[3][91] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][91] ), .Q(\mem_r[3][91] ), .QN( ));
Q_FDP1 \mem_r_REG[3][92] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][92] ), .Q(\mem_r[3][92] ), .QN( ));
Q_FDP1 \mem_r_REG[3][93] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][93] ), .Q(\mem_r[3][93] ), .QN( ));
Q_FDP1 \mem_r_REG[3][94] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][94] ), .Q(\mem_r[3][94] ), .QN( ));
Q_FDP1 \mem_r_REG[3][95] ( .CK(clk), .R(rst_n), .D(\mem_nxt[3][95] ), .Q(\mem_r[3][95] ), .QN( ));
Q_FDP1 \mem_r_REG[2][0] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][0] ), .Q(\mem_r[2][0] ), .QN( ));
Q_FDP1 \mem_r_REG[2][1] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][1] ), .Q(\mem_r[2][1] ), .QN( ));
Q_FDP1 \mem_r_REG[2][2] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][2] ), .Q(\mem_r[2][2] ), .QN( ));
Q_FDP1 \mem_r_REG[2][3] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][3] ), .Q(\mem_r[2][3] ), .QN( ));
Q_FDP1 \mem_r_REG[2][4] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][4] ), .Q(\mem_r[2][4] ), .QN( ));
Q_FDP1 \mem_r_REG[2][5] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][5] ), .Q(\mem_r[2][5] ), .QN( ));
Q_FDP1 \mem_r_REG[2][6] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][6] ), .Q(\mem_r[2][6] ), .QN( ));
Q_FDP1 \mem_r_REG[2][7] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][7] ), .Q(\mem_r[2][7] ), .QN( ));
Q_FDP1 \mem_r_REG[2][8] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][8] ), .Q(\mem_r[2][8] ), .QN( ));
Q_FDP1 \mem_r_REG[2][9] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][9] ), .Q(\mem_r[2][9] ), .QN( ));
Q_FDP1 \mem_r_REG[2][10] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][10] ), .Q(\mem_r[2][10] ), .QN( ));
Q_FDP1 \mem_r_REG[2][11] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][11] ), .Q(\mem_r[2][11] ), .QN( ));
Q_FDP1 \mem_r_REG[2][12] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][12] ), .Q(\mem_r[2][12] ), .QN( ));
Q_FDP1 \mem_r_REG[2][13] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][13] ), .Q(\mem_r[2][13] ), .QN( ));
Q_FDP1 \mem_r_REG[2][14] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][14] ), .Q(\mem_r[2][14] ), .QN( ));
Q_FDP1 \mem_r_REG[2][15] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][15] ), .Q(\mem_r[2][15] ), .QN( ));
Q_FDP1 \mem_r_REG[2][16] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][16] ), .Q(\mem_r[2][16] ), .QN( ));
Q_FDP1 \mem_r_REG[2][17] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][17] ), .Q(\mem_r[2][17] ), .QN( ));
Q_FDP1 \mem_r_REG[2][18] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][18] ), .Q(\mem_r[2][18] ), .QN( ));
Q_FDP1 \mem_r_REG[2][19] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][19] ), .Q(\mem_r[2][19] ), .QN( ));
Q_FDP1 \mem_r_REG[2][20] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][20] ), .Q(\mem_r[2][20] ), .QN( ));
Q_FDP1 \mem_r_REG[2][21] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][21] ), .Q(\mem_r[2][21] ), .QN( ));
Q_FDP1 \mem_r_REG[2][22] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][22] ), .Q(\mem_r[2][22] ), .QN( ));
Q_FDP1 \mem_r_REG[2][23] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][23] ), .Q(\mem_r[2][23] ), .QN( ));
Q_FDP1 \mem_r_REG[2][24] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][24] ), .Q(\mem_r[2][24] ), .QN( ));
Q_FDP1 \mem_r_REG[2][25] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][25] ), .Q(\mem_r[2][25] ), .QN( ));
Q_FDP1 \mem_r_REG[2][26] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][26] ), .Q(\mem_r[2][26] ), .QN( ));
Q_FDP1 \mem_r_REG[2][27] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][27] ), .Q(\mem_r[2][27] ), .QN( ));
Q_FDP1 \mem_r_REG[2][28] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][28] ), .Q(\mem_r[2][28] ), .QN( ));
Q_FDP1 \mem_r_REG[2][29] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][29] ), .Q(\mem_r[2][29] ), .QN( ));
Q_FDP1 \mem_r_REG[2][30] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][30] ), .Q(\mem_r[2][30] ), .QN( ));
Q_FDP1 \mem_r_REG[2][31] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][31] ), .Q(\mem_r[2][31] ), .QN( ));
Q_FDP1 \mem_r_REG[2][32] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][32] ), .Q(\mem_r[2][32] ), .QN( ));
Q_FDP1 \mem_r_REG[2][33] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][33] ), .Q(\mem_r[2][33] ), .QN( ));
Q_FDP1 \mem_r_REG[2][34] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][34] ), .Q(\mem_r[2][34] ), .QN( ));
Q_FDP1 \mem_r_REG[2][35] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][35] ), .Q(\mem_r[2][35] ), .QN( ));
Q_FDP1 \mem_r_REG[2][36] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][36] ), .Q(\mem_r[2][36] ), .QN( ));
Q_FDP1 \mem_r_REG[2][37] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][37] ), .Q(\mem_r[2][37] ), .QN( ));
Q_FDP1 \mem_r_REG[2][38] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][38] ), .Q(\mem_r[2][38] ), .QN( ));
Q_FDP1 \mem_r_REG[2][39] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][39] ), .Q(\mem_r[2][39] ), .QN( ));
Q_FDP1 \mem_r_REG[2][40] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][40] ), .Q(\mem_r[2][40] ), .QN( ));
Q_FDP1 \mem_r_REG[2][41] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][41] ), .Q(\mem_r[2][41] ), .QN( ));
Q_FDP1 \mem_r_REG[2][42] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][42] ), .Q(\mem_r[2][42] ), .QN( ));
Q_FDP1 \mem_r_REG[2][43] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][43] ), .Q(\mem_r[2][43] ), .QN( ));
Q_FDP1 \mem_r_REG[2][44] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][44] ), .Q(\mem_r[2][44] ), .QN( ));
Q_FDP1 \mem_r_REG[2][45] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][45] ), .Q(\mem_r[2][45] ), .QN( ));
Q_FDP1 \mem_r_REG[2][46] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][46] ), .Q(\mem_r[2][46] ), .QN( ));
Q_FDP1 \mem_r_REG[2][47] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][47] ), .Q(\mem_r[2][47] ), .QN( ));
Q_FDP1 \mem_r_REG[2][48] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][48] ), .Q(\mem_r[2][48] ), .QN( ));
Q_FDP1 \mem_r_REG[2][49] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][49] ), .Q(\mem_r[2][49] ), .QN( ));
Q_FDP1 \mem_r_REG[2][50] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][50] ), .Q(\mem_r[2][50] ), .QN( ));
Q_FDP1 \mem_r_REG[2][51] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][51] ), .Q(\mem_r[2][51] ), .QN( ));
Q_FDP1 \mem_r_REG[2][52] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][52] ), .Q(\mem_r[2][52] ), .QN( ));
Q_FDP1 \mem_r_REG[2][53] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][53] ), .Q(\mem_r[2][53] ), .QN( ));
Q_FDP1 \mem_r_REG[2][54] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][54] ), .Q(\mem_r[2][54] ), .QN( ));
Q_FDP1 \mem_r_REG[2][55] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][55] ), .Q(\mem_r[2][55] ), .QN( ));
Q_FDP1 \mem_r_REG[2][56] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][56] ), .Q(\mem_r[2][56] ), .QN( ));
Q_FDP1 \mem_r_REG[2][57] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][57] ), .Q(\mem_r[2][57] ), .QN( ));
Q_FDP1 \mem_r_REG[2][58] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][58] ), .Q(\mem_r[2][58] ), .QN( ));
Q_FDP1 \mem_r_REG[2][59] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][59] ), .Q(\mem_r[2][59] ), .QN( ));
Q_FDP1 \mem_r_REG[2][60] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][60] ), .Q(\mem_r[2][60] ), .QN( ));
Q_FDP1 \mem_r_REG[2][61] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][61] ), .Q(\mem_r[2][61] ), .QN( ));
Q_FDP1 \mem_r_REG[2][62] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][62] ), .Q(\mem_r[2][62] ), .QN( ));
Q_FDP1 \mem_r_REG[2][63] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][63] ), .Q(\mem_r[2][63] ), .QN( ));
Q_FDP1 \mem_r_REG[2][64] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][64] ), .Q(\mem_r[2][64] ), .QN( ));
Q_FDP1 \mem_r_REG[2][65] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][65] ), .Q(\mem_r[2][65] ), .QN( ));
Q_FDP1 \mem_r_REG[2][66] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][66] ), .Q(\mem_r[2][66] ), .QN( ));
Q_FDP1 \mem_r_REG[2][67] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][67] ), .Q(\mem_r[2][67] ), .QN( ));
Q_FDP1 \mem_r_REG[2][68] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][68] ), .Q(\mem_r[2][68] ), .QN( ));
Q_FDP1 \mem_r_REG[2][69] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][69] ), .Q(\mem_r[2][69] ), .QN( ));
Q_FDP1 \mem_r_REG[2][70] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][70] ), .Q(\mem_r[2][70] ), .QN( ));
Q_FDP1 \mem_r_REG[2][71] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][71] ), .Q(\mem_r[2][71] ), .QN( ));
Q_FDP1 \mem_r_REG[2][72] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][72] ), .Q(\mem_r[2][72] ), .QN( ));
Q_FDP1 \mem_r_REG[2][73] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][73] ), .Q(\mem_r[2][73] ), .QN( ));
Q_FDP1 \mem_r_REG[2][74] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][74] ), .Q(\mem_r[2][74] ), .QN( ));
Q_FDP1 \mem_r_REG[2][75] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][75] ), .Q(\mem_r[2][75] ), .QN( ));
Q_FDP1 \mem_r_REG[2][76] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][76] ), .Q(\mem_r[2][76] ), .QN( ));
Q_FDP1 \mem_r_REG[2][77] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][77] ), .Q(\mem_r[2][77] ), .QN( ));
Q_FDP1 \mem_r_REG[2][78] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][78] ), .Q(\mem_r[2][78] ), .QN( ));
Q_FDP1 \mem_r_REG[2][79] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][79] ), .Q(\mem_r[2][79] ), .QN( ));
Q_FDP1 \mem_r_REG[2][80] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][80] ), .Q(\mem_r[2][80] ), .QN( ));
Q_FDP1 \mem_r_REG[2][81] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][81] ), .Q(\mem_r[2][81] ), .QN( ));
Q_FDP1 \mem_r_REG[2][82] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][82] ), .Q(\mem_r[2][82] ), .QN( ));
Q_FDP1 \mem_r_REG[2][83] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][83] ), .Q(\mem_r[2][83] ), .QN( ));
Q_FDP1 \mem_r_REG[2][84] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][84] ), .Q(\mem_r[2][84] ), .QN( ));
Q_FDP1 \mem_r_REG[2][85] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][85] ), .Q(\mem_r[2][85] ), .QN( ));
Q_FDP1 \mem_r_REG[2][86] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][86] ), .Q(\mem_r[2][86] ), .QN( ));
Q_FDP1 \mem_r_REG[2][87] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][87] ), .Q(\mem_r[2][87] ), .QN( ));
Q_FDP1 \mem_r_REG[2][88] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][88] ), .Q(\mem_r[2][88] ), .QN( ));
Q_FDP1 \mem_r_REG[2][89] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][89] ), .Q(\mem_r[2][89] ), .QN( ));
Q_FDP1 \mem_r_REG[2][90] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][90] ), .Q(\mem_r[2][90] ), .QN( ));
Q_FDP1 \mem_r_REG[2][91] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][91] ), .Q(\mem_r[2][91] ), .QN( ));
Q_FDP1 \mem_r_REG[2][92] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][92] ), .Q(\mem_r[2][92] ), .QN( ));
Q_FDP1 \mem_r_REG[2][93] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][93] ), .Q(\mem_r[2][93] ), .QN( ));
Q_FDP1 \mem_r_REG[2][94] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][94] ), .Q(\mem_r[2][94] ), .QN( ));
Q_FDP1 \mem_r_REG[2][95] ( .CK(clk), .R(rst_n), .D(\mem_nxt[2][95] ), .Q(\mem_r[2][95] ), .QN( ));
Q_FDP1 \mem_r_REG[1][0] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][0] ), .Q(\mem_r[1][0] ), .QN( ));
Q_FDP1 \mem_r_REG[1][1] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][1] ), .Q(\mem_r[1][1] ), .QN( ));
Q_FDP1 \mem_r_REG[1][2] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][2] ), .Q(\mem_r[1][2] ), .QN( ));
Q_FDP1 \mem_r_REG[1][3] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][3] ), .Q(\mem_r[1][3] ), .QN( ));
Q_FDP1 \mem_r_REG[1][4] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][4] ), .Q(\mem_r[1][4] ), .QN( ));
Q_FDP1 \mem_r_REG[1][5] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][5] ), .Q(\mem_r[1][5] ), .QN( ));
Q_FDP1 \mem_r_REG[1][6] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][6] ), .Q(\mem_r[1][6] ), .QN( ));
Q_FDP1 \mem_r_REG[1][7] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][7] ), .Q(\mem_r[1][7] ), .QN( ));
Q_FDP1 \mem_r_REG[1][8] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][8] ), .Q(\mem_r[1][8] ), .QN( ));
Q_FDP1 \mem_r_REG[1][9] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][9] ), .Q(\mem_r[1][9] ), .QN( ));
Q_FDP1 \mem_r_REG[1][10] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][10] ), .Q(\mem_r[1][10] ), .QN( ));
Q_FDP1 \mem_r_REG[1][11] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][11] ), .Q(\mem_r[1][11] ), .QN( ));
Q_FDP1 \mem_r_REG[1][12] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][12] ), .Q(\mem_r[1][12] ), .QN( ));
Q_FDP1 \mem_r_REG[1][13] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][13] ), .Q(\mem_r[1][13] ), .QN( ));
Q_FDP1 \mem_r_REG[1][14] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][14] ), .Q(\mem_r[1][14] ), .QN( ));
Q_FDP1 \mem_r_REG[1][15] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][15] ), .Q(\mem_r[1][15] ), .QN( ));
Q_FDP1 \mem_r_REG[1][16] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][16] ), .Q(\mem_r[1][16] ), .QN( ));
Q_FDP1 \mem_r_REG[1][17] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][17] ), .Q(\mem_r[1][17] ), .QN( ));
Q_FDP1 \mem_r_REG[1][18] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][18] ), .Q(\mem_r[1][18] ), .QN( ));
Q_FDP1 \mem_r_REG[1][19] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][19] ), .Q(\mem_r[1][19] ), .QN( ));
Q_FDP1 \mem_r_REG[1][20] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][20] ), .Q(\mem_r[1][20] ), .QN( ));
Q_FDP1 \mem_r_REG[1][21] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][21] ), .Q(\mem_r[1][21] ), .QN( ));
Q_FDP1 \mem_r_REG[1][22] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][22] ), .Q(\mem_r[1][22] ), .QN( ));
Q_FDP1 \mem_r_REG[1][23] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][23] ), .Q(\mem_r[1][23] ), .QN( ));
Q_FDP1 \mem_r_REG[1][24] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][24] ), .Q(\mem_r[1][24] ), .QN( ));
Q_FDP1 \mem_r_REG[1][25] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][25] ), .Q(\mem_r[1][25] ), .QN( ));
Q_FDP1 \mem_r_REG[1][26] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][26] ), .Q(\mem_r[1][26] ), .QN( ));
Q_FDP1 \mem_r_REG[1][27] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][27] ), .Q(\mem_r[1][27] ), .QN( ));
Q_FDP1 \mem_r_REG[1][28] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][28] ), .Q(\mem_r[1][28] ), .QN( ));
Q_FDP1 \mem_r_REG[1][29] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][29] ), .Q(\mem_r[1][29] ), .QN( ));
Q_FDP1 \mem_r_REG[1][30] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][30] ), .Q(\mem_r[1][30] ), .QN( ));
Q_FDP1 \mem_r_REG[1][31] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][31] ), .Q(\mem_r[1][31] ), .QN( ));
Q_FDP1 \mem_r_REG[1][32] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][32] ), .Q(\mem_r[1][32] ), .QN( ));
Q_FDP1 \mem_r_REG[1][33] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][33] ), .Q(\mem_r[1][33] ), .QN( ));
Q_FDP1 \mem_r_REG[1][34] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][34] ), .Q(\mem_r[1][34] ), .QN( ));
Q_FDP1 \mem_r_REG[1][35] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][35] ), .Q(\mem_r[1][35] ), .QN( ));
Q_FDP1 \mem_r_REG[1][36] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][36] ), .Q(\mem_r[1][36] ), .QN( ));
Q_FDP1 \mem_r_REG[1][37] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][37] ), .Q(\mem_r[1][37] ), .QN( ));
Q_FDP1 \mem_r_REG[1][38] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][38] ), .Q(\mem_r[1][38] ), .QN( ));
Q_FDP1 \mem_r_REG[1][39] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][39] ), .Q(\mem_r[1][39] ), .QN( ));
Q_FDP1 \mem_r_REG[1][40] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][40] ), .Q(\mem_r[1][40] ), .QN( ));
Q_FDP1 \mem_r_REG[1][41] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][41] ), .Q(\mem_r[1][41] ), .QN( ));
Q_FDP1 \mem_r_REG[1][42] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][42] ), .Q(\mem_r[1][42] ), .QN( ));
Q_FDP1 \mem_r_REG[1][43] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][43] ), .Q(\mem_r[1][43] ), .QN( ));
Q_FDP1 \mem_r_REG[1][44] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][44] ), .Q(\mem_r[1][44] ), .QN( ));
Q_FDP1 \mem_r_REG[1][45] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][45] ), .Q(\mem_r[1][45] ), .QN( ));
Q_FDP1 \mem_r_REG[1][46] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][46] ), .Q(\mem_r[1][46] ), .QN( ));
Q_FDP1 \mem_r_REG[1][47] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][47] ), .Q(\mem_r[1][47] ), .QN( ));
Q_FDP1 \mem_r_REG[1][48] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][48] ), .Q(\mem_r[1][48] ), .QN( ));
Q_FDP1 \mem_r_REG[1][49] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][49] ), .Q(\mem_r[1][49] ), .QN( ));
Q_FDP1 \mem_r_REG[1][50] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][50] ), .Q(\mem_r[1][50] ), .QN( ));
Q_FDP1 \mem_r_REG[1][51] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][51] ), .Q(\mem_r[1][51] ), .QN( ));
Q_FDP1 \mem_r_REG[1][52] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][52] ), .Q(\mem_r[1][52] ), .QN( ));
Q_FDP1 \mem_r_REG[1][53] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][53] ), .Q(\mem_r[1][53] ), .QN( ));
Q_FDP1 \mem_r_REG[1][54] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][54] ), .Q(\mem_r[1][54] ), .QN( ));
Q_FDP1 \mem_r_REG[1][55] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][55] ), .Q(\mem_r[1][55] ), .QN( ));
Q_FDP1 \mem_r_REG[1][56] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][56] ), .Q(\mem_r[1][56] ), .QN( ));
Q_FDP1 \mem_r_REG[1][57] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][57] ), .Q(\mem_r[1][57] ), .QN( ));
Q_FDP1 \mem_r_REG[1][58] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][58] ), .Q(\mem_r[1][58] ), .QN( ));
Q_FDP1 \mem_r_REG[1][59] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][59] ), .Q(\mem_r[1][59] ), .QN( ));
Q_FDP1 \mem_r_REG[1][60] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][60] ), .Q(\mem_r[1][60] ), .QN( ));
Q_FDP1 \mem_r_REG[1][61] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][61] ), .Q(\mem_r[1][61] ), .QN( ));
Q_FDP1 \mem_r_REG[1][62] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][62] ), .Q(\mem_r[1][62] ), .QN( ));
Q_FDP1 \mem_r_REG[1][63] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][63] ), .Q(\mem_r[1][63] ), .QN( ));
Q_FDP1 \mem_r_REG[1][64] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][64] ), .Q(\mem_r[1][64] ), .QN( ));
Q_FDP1 \mem_r_REG[1][65] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][65] ), .Q(\mem_r[1][65] ), .QN( ));
Q_FDP1 \mem_r_REG[1][66] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][66] ), .Q(\mem_r[1][66] ), .QN( ));
Q_FDP1 \mem_r_REG[1][67] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][67] ), .Q(\mem_r[1][67] ), .QN( ));
Q_FDP1 \mem_r_REG[1][68] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][68] ), .Q(\mem_r[1][68] ), .QN( ));
Q_FDP1 \mem_r_REG[1][69] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][69] ), .Q(\mem_r[1][69] ), .QN( ));
Q_FDP1 \mem_r_REG[1][70] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][70] ), .Q(\mem_r[1][70] ), .QN( ));
Q_FDP1 \mem_r_REG[1][71] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][71] ), .Q(\mem_r[1][71] ), .QN( ));
Q_FDP1 \mem_r_REG[1][72] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][72] ), .Q(\mem_r[1][72] ), .QN( ));
Q_FDP1 \mem_r_REG[1][73] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][73] ), .Q(\mem_r[1][73] ), .QN( ));
Q_FDP1 \mem_r_REG[1][74] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][74] ), .Q(\mem_r[1][74] ), .QN( ));
Q_FDP1 \mem_r_REG[1][75] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][75] ), .Q(\mem_r[1][75] ), .QN( ));
Q_FDP1 \mem_r_REG[1][76] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][76] ), .Q(\mem_r[1][76] ), .QN( ));
Q_FDP1 \mem_r_REG[1][77] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][77] ), .Q(\mem_r[1][77] ), .QN( ));
Q_FDP1 \mem_r_REG[1][78] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][78] ), .Q(\mem_r[1][78] ), .QN( ));
Q_FDP1 \mem_r_REG[1][79] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][79] ), .Q(\mem_r[1][79] ), .QN( ));
Q_FDP1 \mem_r_REG[1][80] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][80] ), .Q(\mem_r[1][80] ), .QN( ));
Q_FDP1 \mem_r_REG[1][81] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][81] ), .Q(\mem_r[1][81] ), .QN( ));
Q_FDP1 \mem_r_REG[1][82] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][82] ), .Q(\mem_r[1][82] ), .QN( ));
Q_FDP1 \mem_r_REG[1][83] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][83] ), .Q(\mem_r[1][83] ), .QN( ));
Q_FDP1 \mem_r_REG[1][84] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][84] ), .Q(\mem_r[1][84] ), .QN( ));
Q_FDP1 \mem_r_REG[1][85] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][85] ), .Q(\mem_r[1][85] ), .QN( ));
Q_FDP1 \mem_r_REG[1][86] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][86] ), .Q(\mem_r[1][86] ), .QN( ));
Q_FDP1 \mem_r_REG[1][87] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][87] ), .Q(\mem_r[1][87] ), .QN( ));
Q_FDP1 \mem_r_REG[1][88] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][88] ), .Q(\mem_r[1][88] ), .QN( ));
Q_FDP1 \mem_r_REG[1][89] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][89] ), .Q(\mem_r[1][89] ), .QN( ));
Q_FDP1 \mem_r_REG[1][90] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][90] ), .Q(\mem_r[1][90] ), .QN( ));
Q_FDP1 \mem_r_REG[1][91] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][91] ), .Q(\mem_r[1][91] ), .QN( ));
Q_FDP1 \mem_r_REG[1][92] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][92] ), .Q(\mem_r[1][92] ), .QN( ));
Q_FDP1 \mem_r_REG[1][93] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][93] ), .Q(\mem_r[1][93] ), .QN( ));
Q_FDP1 \mem_r_REG[1][94] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][94] ), .Q(\mem_r[1][94] ), .QN( ));
Q_FDP1 \mem_r_REG[1][95] ( .CK(clk), .R(rst_n), .D(\mem_nxt[1][95] ), .Q(\mem_r[1][95] ), .QN( ));
Q_FDP1 \mem_r_REG[0][0] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][0] ), .Q(\mem_r[0][0] ), .QN( ));
Q_FDP1 \mem_r_REG[0][1] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][1] ), .Q(\mem_r[0][1] ), .QN( ));
Q_FDP1 \mem_r_REG[0][2] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][2] ), .Q(\mem_r[0][2] ), .QN( ));
Q_FDP1 \mem_r_REG[0][3] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][3] ), .Q(\mem_r[0][3] ), .QN( ));
Q_FDP1 \mem_r_REG[0][4] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][4] ), .Q(\mem_r[0][4] ), .QN( ));
Q_FDP1 \mem_r_REG[0][5] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][5] ), .Q(\mem_r[0][5] ), .QN( ));
Q_FDP1 \mem_r_REG[0][6] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][6] ), .Q(\mem_r[0][6] ), .QN( ));
Q_FDP1 \mem_r_REG[0][7] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][7] ), .Q(\mem_r[0][7] ), .QN( ));
Q_FDP1 \mem_r_REG[0][8] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][8] ), .Q(\mem_r[0][8] ), .QN( ));
Q_FDP1 \mem_r_REG[0][9] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][9] ), .Q(\mem_r[0][9] ), .QN( ));
Q_FDP1 \mem_r_REG[0][10] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][10] ), .Q(\mem_r[0][10] ), .QN( ));
Q_FDP1 \mem_r_REG[0][11] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][11] ), .Q(\mem_r[0][11] ), .QN( ));
Q_FDP1 \mem_r_REG[0][12] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][12] ), .Q(\mem_r[0][12] ), .QN( ));
Q_FDP1 \mem_r_REG[0][13] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][13] ), .Q(\mem_r[0][13] ), .QN( ));
Q_FDP1 \mem_r_REG[0][14] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][14] ), .Q(\mem_r[0][14] ), .QN( ));
Q_FDP1 \mem_r_REG[0][15] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][15] ), .Q(\mem_r[0][15] ), .QN( ));
Q_FDP1 \mem_r_REG[0][16] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][16] ), .Q(\mem_r[0][16] ), .QN( ));
Q_FDP1 \mem_r_REG[0][17] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][17] ), .Q(\mem_r[0][17] ), .QN( ));
Q_FDP1 \mem_r_REG[0][18] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][18] ), .Q(\mem_r[0][18] ), .QN( ));
Q_FDP1 \mem_r_REG[0][19] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][19] ), .Q(\mem_r[0][19] ), .QN( ));
Q_FDP1 \mem_r_REG[0][20] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][20] ), .Q(\mem_r[0][20] ), .QN( ));
Q_FDP1 \mem_r_REG[0][21] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][21] ), .Q(\mem_r[0][21] ), .QN( ));
Q_FDP1 \mem_r_REG[0][22] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][22] ), .Q(\mem_r[0][22] ), .QN( ));
Q_FDP1 \mem_r_REG[0][23] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][23] ), .Q(\mem_r[0][23] ), .QN( ));
Q_FDP1 \mem_r_REG[0][24] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][24] ), .Q(\mem_r[0][24] ), .QN( ));
Q_FDP1 \mem_r_REG[0][25] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][25] ), .Q(\mem_r[0][25] ), .QN( ));
Q_FDP1 \mem_r_REG[0][26] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][26] ), .Q(\mem_r[0][26] ), .QN( ));
Q_FDP1 \mem_r_REG[0][27] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][27] ), .Q(\mem_r[0][27] ), .QN( ));
Q_FDP1 \mem_r_REG[0][28] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][28] ), .Q(\mem_r[0][28] ), .QN( ));
Q_FDP1 \mem_r_REG[0][29] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][29] ), .Q(\mem_r[0][29] ), .QN( ));
Q_FDP1 \mem_r_REG[0][30] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][30] ), .Q(\mem_r[0][30] ), .QN( ));
Q_FDP1 \mem_r_REG[0][31] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][31] ), .Q(\mem_r[0][31] ), .QN( ));
Q_FDP1 \mem_r_REG[0][32] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][32] ), .Q(\mem_r[0][32] ), .QN( ));
Q_FDP1 \mem_r_REG[0][33] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][33] ), .Q(\mem_r[0][33] ), .QN( ));
Q_FDP1 \mem_r_REG[0][34] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][34] ), .Q(\mem_r[0][34] ), .QN( ));
Q_FDP1 \mem_r_REG[0][35] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][35] ), .Q(\mem_r[0][35] ), .QN( ));
Q_FDP1 \mem_r_REG[0][36] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][36] ), .Q(\mem_r[0][36] ), .QN( ));
Q_FDP1 \mem_r_REG[0][37] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][37] ), .Q(\mem_r[0][37] ), .QN( ));
Q_FDP1 \mem_r_REG[0][38] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][38] ), .Q(\mem_r[0][38] ), .QN( ));
Q_FDP1 \mem_r_REG[0][39] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][39] ), .Q(\mem_r[0][39] ), .QN( ));
Q_FDP1 \mem_r_REG[0][40] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][40] ), .Q(\mem_r[0][40] ), .QN( ));
Q_FDP1 \mem_r_REG[0][41] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][41] ), .Q(\mem_r[0][41] ), .QN( ));
Q_FDP1 \mem_r_REG[0][42] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][42] ), .Q(\mem_r[0][42] ), .QN( ));
Q_FDP1 \mem_r_REG[0][43] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][43] ), .Q(\mem_r[0][43] ), .QN( ));
Q_FDP1 \mem_r_REG[0][44] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][44] ), .Q(\mem_r[0][44] ), .QN( ));
Q_FDP1 \mem_r_REG[0][45] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][45] ), .Q(\mem_r[0][45] ), .QN( ));
Q_FDP1 \mem_r_REG[0][46] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][46] ), .Q(\mem_r[0][46] ), .QN( ));
Q_FDP1 \mem_r_REG[0][47] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][47] ), .Q(\mem_r[0][47] ), .QN( ));
Q_FDP1 \mem_r_REG[0][48] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][48] ), .Q(\mem_r[0][48] ), .QN( ));
Q_FDP1 \mem_r_REG[0][49] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][49] ), .Q(\mem_r[0][49] ), .QN( ));
Q_FDP1 \mem_r_REG[0][50] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][50] ), .Q(\mem_r[0][50] ), .QN( ));
Q_FDP1 \mem_r_REG[0][51] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][51] ), .Q(\mem_r[0][51] ), .QN( ));
Q_FDP1 \mem_r_REG[0][52] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][52] ), .Q(\mem_r[0][52] ), .QN( ));
Q_FDP1 \mem_r_REG[0][53] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][53] ), .Q(\mem_r[0][53] ), .QN( ));
Q_FDP1 \mem_r_REG[0][54] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][54] ), .Q(\mem_r[0][54] ), .QN( ));
Q_FDP1 \mem_r_REG[0][55] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][55] ), .Q(\mem_r[0][55] ), .QN( ));
Q_FDP1 \mem_r_REG[0][56] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][56] ), .Q(\mem_r[0][56] ), .QN( ));
Q_FDP1 \mem_r_REG[0][57] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][57] ), .Q(\mem_r[0][57] ), .QN( ));
Q_FDP1 \mem_r_REG[0][58] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][58] ), .Q(\mem_r[0][58] ), .QN( ));
Q_FDP1 \mem_r_REG[0][59] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][59] ), .Q(\mem_r[0][59] ), .QN( ));
Q_FDP1 \mem_r_REG[0][60] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][60] ), .Q(\mem_r[0][60] ), .QN( ));
Q_FDP1 \mem_r_REG[0][61] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][61] ), .Q(\mem_r[0][61] ), .QN( ));
Q_FDP1 \mem_r_REG[0][62] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][62] ), .Q(\mem_r[0][62] ), .QN( ));
Q_FDP1 \mem_r_REG[0][63] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][63] ), .Q(\mem_r[0][63] ), .QN( ));
Q_FDP1 \mem_r_REG[0][64] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][64] ), .Q(\mem_r[0][64] ), .QN( ));
Q_FDP1 \mem_r_REG[0][65] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][65] ), .Q(\mem_r[0][65] ), .QN( ));
Q_FDP1 \mem_r_REG[0][66] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][66] ), .Q(\mem_r[0][66] ), .QN( ));
Q_FDP1 \mem_r_REG[0][67] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][67] ), .Q(\mem_r[0][67] ), .QN( ));
Q_FDP1 \mem_r_REG[0][68] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][68] ), .Q(\mem_r[0][68] ), .QN( ));
Q_FDP1 \mem_r_REG[0][69] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][69] ), .Q(\mem_r[0][69] ), .QN( ));
Q_FDP1 \mem_r_REG[0][70] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][70] ), .Q(\mem_r[0][70] ), .QN( ));
Q_FDP1 \mem_r_REG[0][71] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][71] ), .Q(\mem_r[0][71] ), .QN( ));
Q_FDP1 \mem_r_REG[0][72] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][72] ), .Q(\mem_r[0][72] ), .QN( ));
Q_FDP1 \mem_r_REG[0][73] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][73] ), .Q(\mem_r[0][73] ), .QN( ));
Q_FDP1 \mem_r_REG[0][74] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][74] ), .Q(\mem_r[0][74] ), .QN( ));
Q_FDP1 \mem_r_REG[0][75] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][75] ), .Q(\mem_r[0][75] ), .QN( ));
Q_FDP1 \mem_r_REG[0][76] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][76] ), .Q(\mem_r[0][76] ), .QN( ));
Q_FDP1 \mem_r_REG[0][77] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][77] ), .Q(\mem_r[0][77] ), .QN( ));
Q_FDP1 \mem_r_REG[0][78] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][78] ), .Q(\mem_r[0][78] ), .QN( ));
Q_FDP1 \mem_r_REG[0][79] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][79] ), .Q(\mem_r[0][79] ), .QN( ));
Q_FDP1 \mem_r_REG[0][80] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][80] ), .Q(\mem_r[0][80] ), .QN( ));
Q_FDP1 \mem_r_REG[0][81] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][81] ), .Q(\mem_r[0][81] ), .QN( ));
Q_FDP1 \mem_r_REG[0][82] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][82] ), .Q(\mem_r[0][82] ), .QN( ));
Q_FDP1 \mem_r_REG[0][83] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][83] ), .Q(\mem_r[0][83] ), .QN( ));
Q_FDP1 \mem_r_REG[0][84] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][84] ), .Q(\mem_r[0][84] ), .QN( ));
Q_FDP1 \mem_r_REG[0][85] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][85] ), .Q(\mem_r[0][85] ), .QN( ));
Q_FDP1 \mem_r_REG[0][86] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][86] ), .Q(\mem_r[0][86] ), .QN( ));
Q_FDP1 \mem_r_REG[0][87] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][87] ), .Q(\mem_r[0][87] ), .QN( ));
Q_FDP1 \mem_r_REG[0][88] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][88] ), .Q(\mem_r[0][88] ), .QN( ));
Q_FDP1 \mem_r_REG[0][89] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][89] ), .Q(\mem_r[0][89] ), .QN( ));
Q_FDP1 \mem_r_REG[0][90] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][90] ), .Q(\mem_r[0][90] ), .QN( ));
Q_FDP1 \mem_r_REG[0][91] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][91] ), .Q(\mem_r[0][91] ), .QN( ));
Q_FDP1 \mem_r_REG[0][92] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][92] ), .Q(\mem_r[0][92] ), .QN( ));
Q_FDP1 \mem_r_REG[0][93] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][93] ), .Q(\mem_r[0][93] ), .QN( ));
Q_FDP1 \mem_r_REG[0][94] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][94] ), .Q(\mem_r[0][94] ), .QN( ));
Q_FDP1 \mem_r_REG[0][95] ( .CK(clk), .R(rst_n), .D(\mem_nxt[0][95] ), .Q(\mem_r[0][95] ), .QN( ));
Q_AD01HF U1697 ( .A0(wr_ptr_r[1]), .B0(wr_ptr_r[0]), .S(n57), .CO(n58));
Q_AD01HF U1698 ( .A0(wr_ptr_r[2]), .B0(n58), .S(n59), .CO(n60));
Q_XOR2 U1699 ( .A0(wr_ptr_r[3]), .A1(n60), .Z(n61));
Q_AN02 U1700 ( .A0(n53), .A1(wr_ptr_r[0]), .Z(n62));
Q_MX02 U1701 ( .S(n66), .A0(n62), .A1(n40), .Z(wr_ptr_nxt[0]));
Q_AN02 U1702 ( .A0(n53), .A1(wr_ptr_r[1]), .Z(n63));
Q_MX02 U1703 ( .S(n66), .A0(n63), .A1(n57), .Z(wr_ptr_nxt[1]));
Q_AN02 U1704 ( .A0(n53), .A1(wr_ptr_r[2]), .Z(n64));
Q_MX02 U1705 ( .S(n66), .A0(n64), .A1(n59), .Z(wr_ptr_nxt[2]));
Q_XOR2 U1706 ( .A0(n44), .A1(wr_ptr_r[3]), .Z(n65));
Q_MX02 U1707 ( .S(n66), .A0(n65), .A1(n61), .Z(wr_ptr_nxt[3]));
Q_NR02 U1708 ( .A0(n67), .A1(n53), .Z(n66));
Q_AN03 U1709 ( .A0(n54), .A1(n69), .A2(n68), .Z(n67));
Q_NR02 U1710 ( .A0(n59), .A1(n57), .Z(n69));
Q_AN03 U1711 ( .A0(wr_en), .A1(n60), .A2(wr_ptr_r[0]), .Z(n68));
Q_AD01HF U1712 ( .A0(rd_ptr_r[1]), .B0(rd_ptr_r[0]), .S(n70), .CO(n71));
Q_AD01HF U1713 ( .A0(rd_ptr_r[2]), .B0(n71), .S(n72), .CO(n73));
Q_XOR2 U1714 ( .A0(rd_ptr_r[3]), .A1(n73), .Z(n74));
Q_AN02 U1715 ( .A0(n84), .A1(rd_ptr_r[0]), .Z(n75));
Q_MX02 U1716 ( .S(n85), .A0(n75), .A1(n86), .Z(rd_ptr_nxt[0]));
Q_AN02 U1717 ( .A0(n84), .A1(rd_ptr_r[1]), .Z(n76));
Q_MX02 U1718 ( .S(n85), .A0(n76), .A1(n70), .Z(rd_ptr_nxt[1]));
Q_AN02 U1719 ( .A0(n84), .A1(rd_ptr_r[2]), .Z(n77));
Q_MX02 U1720 ( .S(n85), .A0(n77), .A1(n72), .Z(rd_ptr_nxt[2]));
Q_XNR2 U1721 ( .A0(n84), .A1(rd_ptr_r[3]), .Z(n78));
Q_MX02 U1722 ( .S(n85), .A0(n78), .A1(n74), .Z(rd_ptr_nxt[3]));
Q_OR02 U1723 ( .A0(n79), .A1(empty_i), .Z(n84));
Q_INV U1724 ( .A(n84), .Z(n80));
Q_INV U1725 ( .A(rd_en), .Z(n79));
Q_OA21 U1726 ( .A0(n81), .A1(n82), .B0(n80), .Z(n85));
Q_INV U1727 ( .A(n73), .Z(n83));
Q_OR02 U1728 ( .A0(n83), .A1(n72), .Z(n81));
Q_OR02 U1729 ( .A0(n70), .A1(n86), .Z(n82));
Q_MX08 U1730 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][0] ), .A1(\mem_r[1][0] ), .A2(\mem_r[2][0] ), .A3(\mem_r[3][0] ), .A4(\mem_r[4][0] ), .A5(\mem_r[5][0] ), .A6(\mem_r[6][0] ), .A7(\mem_r[7][0] ), .Z(dout_i[0]));
Q_MX08 U1731 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][1] ), .A1(\mem_r[1][1] ), .A2(\mem_r[2][1] ), .A3(\mem_r[3][1] ), .A4(\mem_r[4][1] ), .A5(\mem_r[5][1] ), .A6(\mem_r[6][1] ), .A7(\mem_r[7][1] ), .Z(dout_i[1]));
Q_MX08 U1732 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][2] ), .A1(\mem_r[1][2] ), .A2(\mem_r[2][2] ), .A3(\mem_r[3][2] ), .A4(\mem_r[4][2] ), .A5(\mem_r[5][2] ), .A6(\mem_r[6][2] ), .A7(\mem_r[7][2] ), .Z(dout_i[2]));
Q_MX08 U1733 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][3] ), .A1(\mem_r[1][3] ), .A2(\mem_r[2][3] ), .A3(\mem_r[3][3] ), .A4(\mem_r[4][3] ), .A5(\mem_r[5][3] ), .A6(\mem_r[6][3] ), .A7(\mem_r[7][3] ), .Z(dout_i[3]));
Q_MX08 U1734 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][4] ), .A1(\mem_r[1][4] ), .A2(\mem_r[2][4] ), .A3(\mem_r[3][4] ), .A4(\mem_r[4][4] ), .A5(\mem_r[5][4] ), .A6(\mem_r[6][4] ), .A7(\mem_r[7][4] ), .Z(dout_i[4]));
Q_MX08 U1735 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][5] ), .A1(\mem_r[1][5] ), .A2(\mem_r[2][5] ), .A3(\mem_r[3][5] ), .A4(\mem_r[4][5] ), .A5(\mem_r[5][5] ), .A6(\mem_r[6][5] ), .A7(\mem_r[7][5] ), .Z(dout_i[5]));
Q_MX08 U1736 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][6] ), .A1(\mem_r[1][6] ), .A2(\mem_r[2][6] ), .A3(\mem_r[3][6] ), .A4(\mem_r[4][6] ), .A5(\mem_r[5][6] ), .A6(\mem_r[6][6] ), .A7(\mem_r[7][6] ), .Z(dout_i[6]));
Q_MX08 U1737 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][7] ), .A1(\mem_r[1][7] ), .A2(\mem_r[2][7] ), .A3(\mem_r[3][7] ), .A4(\mem_r[4][7] ), .A5(\mem_r[5][7] ), .A6(\mem_r[6][7] ), .A7(\mem_r[7][7] ), .Z(dout_i[7]));
Q_MX08 U1738 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][8] ), .A1(\mem_r[1][8] ), .A2(\mem_r[2][8] ), .A3(\mem_r[3][8] ), .A4(\mem_r[4][8] ), .A5(\mem_r[5][8] ), .A6(\mem_r[6][8] ), .A7(\mem_r[7][8] ), .Z(dout_i[8]));
Q_MX08 U1739 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][9] ), .A1(\mem_r[1][9] ), .A2(\mem_r[2][9] ), .A3(\mem_r[3][9] ), .A4(\mem_r[4][9] ), .A5(\mem_r[5][9] ), .A6(\mem_r[6][9] ), .A7(\mem_r[7][9] ), .Z(dout_i[9]));
Q_MX08 U1740 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][10] ), .A1(\mem_r[1][10] ), .A2(\mem_r[2][10] ), .A3(\mem_r[3][10] ), .A4(\mem_r[4][10] ), .A5(\mem_r[5][10] ), .A6(\mem_r[6][10] ), .A7(\mem_r[7][10] ), .Z(dout_i[10]));
Q_MX08 U1741 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][11] ), .A1(\mem_r[1][11] ), .A2(\mem_r[2][11] ), .A3(\mem_r[3][11] ), .A4(\mem_r[4][11] ), .A5(\mem_r[5][11] ), .A6(\mem_r[6][11] ), .A7(\mem_r[7][11] ), .Z(dout_i[11]));
Q_MX08 U1742 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][12] ), .A1(\mem_r[1][12] ), .A2(\mem_r[2][12] ), .A3(\mem_r[3][12] ), .A4(\mem_r[4][12] ), .A5(\mem_r[5][12] ), .A6(\mem_r[6][12] ), .A7(\mem_r[7][12] ), .Z(dout_i[12]));
Q_MX08 U1743 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][13] ), .A1(\mem_r[1][13] ), .A2(\mem_r[2][13] ), .A3(\mem_r[3][13] ), .A4(\mem_r[4][13] ), .A5(\mem_r[5][13] ), .A6(\mem_r[6][13] ), .A7(\mem_r[7][13] ), .Z(dout_i[13]));
Q_MX08 U1744 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][14] ), .A1(\mem_r[1][14] ), .A2(\mem_r[2][14] ), .A3(\mem_r[3][14] ), .A4(\mem_r[4][14] ), .A5(\mem_r[5][14] ), .A6(\mem_r[6][14] ), .A7(\mem_r[7][14] ), .Z(dout_i[14]));
Q_MX08 U1745 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][15] ), .A1(\mem_r[1][15] ), .A2(\mem_r[2][15] ), .A3(\mem_r[3][15] ), .A4(\mem_r[4][15] ), .A5(\mem_r[5][15] ), .A6(\mem_r[6][15] ), .A7(\mem_r[7][15] ), .Z(dout_i[15]));
Q_MX08 U1746 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][16] ), .A1(\mem_r[1][16] ), .A2(\mem_r[2][16] ), .A3(\mem_r[3][16] ), .A4(\mem_r[4][16] ), .A5(\mem_r[5][16] ), .A6(\mem_r[6][16] ), .A7(\mem_r[7][16] ), .Z(dout_i[16]));
Q_MX08 U1747 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][17] ), .A1(\mem_r[1][17] ), .A2(\mem_r[2][17] ), .A3(\mem_r[3][17] ), .A4(\mem_r[4][17] ), .A5(\mem_r[5][17] ), .A6(\mem_r[6][17] ), .A7(\mem_r[7][17] ), .Z(dout_i[17]));
Q_MX08 U1748 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][18] ), .A1(\mem_r[1][18] ), .A2(\mem_r[2][18] ), .A3(\mem_r[3][18] ), .A4(\mem_r[4][18] ), .A5(\mem_r[5][18] ), .A6(\mem_r[6][18] ), .A7(\mem_r[7][18] ), .Z(dout_i[18]));
Q_MX08 U1749 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][19] ), .A1(\mem_r[1][19] ), .A2(\mem_r[2][19] ), .A3(\mem_r[3][19] ), .A4(\mem_r[4][19] ), .A5(\mem_r[5][19] ), .A6(\mem_r[6][19] ), .A7(\mem_r[7][19] ), .Z(dout_i[19]));
Q_MX08 U1750 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][20] ), .A1(\mem_r[1][20] ), .A2(\mem_r[2][20] ), .A3(\mem_r[3][20] ), .A4(\mem_r[4][20] ), .A5(\mem_r[5][20] ), .A6(\mem_r[6][20] ), .A7(\mem_r[7][20] ), .Z(dout_i[20]));
Q_MX08 U1751 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][21] ), .A1(\mem_r[1][21] ), .A2(\mem_r[2][21] ), .A3(\mem_r[3][21] ), .A4(\mem_r[4][21] ), .A5(\mem_r[5][21] ), .A6(\mem_r[6][21] ), .A7(\mem_r[7][21] ), .Z(dout_i[21]));
Q_MX08 U1752 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][22] ), .A1(\mem_r[1][22] ), .A2(\mem_r[2][22] ), .A3(\mem_r[3][22] ), .A4(\mem_r[4][22] ), .A5(\mem_r[5][22] ), .A6(\mem_r[6][22] ), .A7(\mem_r[7][22] ), .Z(dout_i[22]));
Q_MX08 U1753 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][23] ), .A1(\mem_r[1][23] ), .A2(\mem_r[2][23] ), .A3(\mem_r[3][23] ), .A4(\mem_r[4][23] ), .A5(\mem_r[5][23] ), .A6(\mem_r[6][23] ), .A7(\mem_r[7][23] ), .Z(dout_i[23]));
Q_MX08 U1754 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][24] ), .A1(\mem_r[1][24] ), .A2(\mem_r[2][24] ), .A3(\mem_r[3][24] ), .A4(\mem_r[4][24] ), .A5(\mem_r[5][24] ), .A6(\mem_r[6][24] ), .A7(\mem_r[7][24] ), .Z(dout_i[24]));
Q_MX08 U1755 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][25] ), .A1(\mem_r[1][25] ), .A2(\mem_r[2][25] ), .A3(\mem_r[3][25] ), .A4(\mem_r[4][25] ), .A5(\mem_r[5][25] ), .A6(\mem_r[6][25] ), .A7(\mem_r[7][25] ), .Z(dout_i[25]));
Q_MX08 U1756 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][26] ), .A1(\mem_r[1][26] ), .A2(\mem_r[2][26] ), .A3(\mem_r[3][26] ), .A4(\mem_r[4][26] ), .A5(\mem_r[5][26] ), .A6(\mem_r[6][26] ), .A7(\mem_r[7][26] ), .Z(dout_i[26]));
Q_MX08 U1757 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][27] ), .A1(\mem_r[1][27] ), .A2(\mem_r[2][27] ), .A3(\mem_r[3][27] ), .A4(\mem_r[4][27] ), .A5(\mem_r[5][27] ), .A6(\mem_r[6][27] ), .A7(\mem_r[7][27] ), .Z(dout_i[27]));
Q_MX08 U1758 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][28] ), .A1(\mem_r[1][28] ), .A2(\mem_r[2][28] ), .A3(\mem_r[3][28] ), .A4(\mem_r[4][28] ), .A5(\mem_r[5][28] ), .A6(\mem_r[6][28] ), .A7(\mem_r[7][28] ), .Z(dout_i[28]));
Q_MX08 U1759 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][29] ), .A1(\mem_r[1][29] ), .A2(\mem_r[2][29] ), .A3(\mem_r[3][29] ), .A4(\mem_r[4][29] ), .A5(\mem_r[5][29] ), .A6(\mem_r[6][29] ), .A7(\mem_r[7][29] ), .Z(dout_i[29]));
Q_MX08 U1760 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][30] ), .A1(\mem_r[1][30] ), .A2(\mem_r[2][30] ), .A3(\mem_r[3][30] ), .A4(\mem_r[4][30] ), .A5(\mem_r[5][30] ), .A6(\mem_r[6][30] ), .A7(\mem_r[7][30] ), .Z(dout_i[30]));
Q_MX08 U1761 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][31] ), .A1(\mem_r[1][31] ), .A2(\mem_r[2][31] ), .A3(\mem_r[3][31] ), .A4(\mem_r[4][31] ), .A5(\mem_r[5][31] ), .A6(\mem_r[6][31] ), .A7(\mem_r[7][31] ), .Z(dout_i[31]));
Q_MX08 U1762 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][32] ), .A1(\mem_r[1][32] ), .A2(\mem_r[2][32] ), .A3(\mem_r[3][32] ), .A4(\mem_r[4][32] ), .A5(\mem_r[5][32] ), .A6(\mem_r[6][32] ), .A7(\mem_r[7][32] ), .Z(dout_i[32]));
Q_MX08 U1763 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][33] ), .A1(\mem_r[1][33] ), .A2(\mem_r[2][33] ), .A3(\mem_r[3][33] ), .A4(\mem_r[4][33] ), .A5(\mem_r[5][33] ), .A6(\mem_r[6][33] ), .A7(\mem_r[7][33] ), .Z(dout_i[33]));
Q_MX08 U1764 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][34] ), .A1(\mem_r[1][34] ), .A2(\mem_r[2][34] ), .A3(\mem_r[3][34] ), .A4(\mem_r[4][34] ), .A5(\mem_r[5][34] ), .A6(\mem_r[6][34] ), .A7(\mem_r[7][34] ), .Z(dout_i[34]));
Q_MX08 U1765 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][35] ), .A1(\mem_r[1][35] ), .A2(\mem_r[2][35] ), .A3(\mem_r[3][35] ), .A4(\mem_r[4][35] ), .A5(\mem_r[5][35] ), .A6(\mem_r[6][35] ), .A7(\mem_r[7][35] ), .Z(dout_i[35]));
Q_MX08 U1766 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][36] ), .A1(\mem_r[1][36] ), .A2(\mem_r[2][36] ), .A3(\mem_r[3][36] ), .A4(\mem_r[4][36] ), .A5(\mem_r[5][36] ), .A6(\mem_r[6][36] ), .A7(\mem_r[7][36] ), .Z(dout_i[36]));
Q_MX08 U1767 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][37] ), .A1(\mem_r[1][37] ), .A2(\mem_r[2][37] ), .A3(\mem_r[3][37] ), .A4(\mem_r[4][37] ), .A5(\mem_r[5][37] ), .A6(\mem_r[6][37] ), .A7(\mem_r[7][37] ), .Z(dout_i[37]));
Q_MX08 U1768 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][38] ), .A1(\mem_r[1][38] ), .A2(\mem_r[2][38] ), .A3(\mem_r[3][38] ), .A4(\mem_r[4][38] ), .A5(\mem_r[5][38] ), .A6(\mem_r[6][38] ), .A7(\mem_r[7][38] ), .Z(dout_i[38]));
Q_MX08 U1769 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][39] ), .A1(\mem_r[1][39] ), .A2(\mem_r[2][39] ), .A3(\mem_r[3][39] ), .A4(\mem_r[4][39] ), .A5(\mem_r[5][39] ), .A6(\mem_r[6][39] ), .A7(\mem_r[7][39] ), .Z(dout_i[39]));
Q_MX08 U1770 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][40] ), .A1(\mem_r[1][40] ), .A2(\mem_r[2][40] ), .A3(\mem_r[3][40] ), .A4(\mem_r[4][40] ), .A5(\mem_r[5][40] ), .A6(\mem_r[6][40] ), .A7(\mem_r[7][40] ), .Z(dout_i[40]));
Q_MX08 U1771 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][41] ), .A1(\mem_r[1][41] ), .A2(\mem_r[2][41] ), .A3(\mem_r[3][41] ), .A4(\mem_r[4][41] ), .A5(\mem_r[5][41] ), .A6(\mem_r[6][41] ), .A7(\mem_r[7][41] ), .Z(dout_i[41]));
Q_MX08 U1772 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][42] ), .A1(\mem_r[1][42] ), .A2(\mem_r[2][42] ), .A3(\mem_r[3][42] ), .A4(\mem_r[4][42] ), .A5(\mem_r[5][42] ), .A6(\mem_r[6][42] ), .A7(\mem_r[7][42] ), .Z(dout_i[42]));
Q_MX08 U1773 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][43] ), .A1(\mem_r[1][43] ), .A2(\mem_r[2][43] ), .A3(\mem_r[3][43] ), .A4(\mem_r[4][43] ), .A5(\mem_r[5][43] ), .A6(\mem_r[6][43] ), .A7(\mem_r[7][43] ), .Z(dout_i[43]));
Q_MX08 U1774 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][44] ), .A1(\mem_r[1][44] ), .A2(\mem_r[2][44] ), .A3(\mem_r[3][44] ), .A4(\mem_r[4][44] ), .A5(\mem_r[5][44] ), .A6(\mem_r[6][44] ), .A7(\mem_r[7][44] ), .Z(dout_i[44]));
Q_MX08 U1775 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][45] ), .A1(\mem_r[1][45] ), .A2(\mem_r[2][45] ), .A3(\mem_r[3][45] ), .A4(\mem_r[4][45] ), .A5(\mem_r[5][45] ), .A6(\mem_r[6][45] ), .A7(\mem_r[7][45] ), .Z(dout_i[45]));
Q_MX08 U1776 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][46] ), .A1(\mem_r[1][46] ), .A2(\mem_r[2][46] ), .A3(\mem_r[3][46] ), .A4(\mem_r[4][46] ), .A5(\mem_r[5][46] ), .A6(\mem_r[6][46] ), .A7(\mem_r[7][46] ), .Z(dout_i[46]));
Q_MX08 U1777 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][47] ), .A1(\mem_r[1][47] ), .A2(\mem_r[2][47] ), .A3(\mem_r[3][47] ), .A4(\mem_r[4][47] ), .A5(\mem_r[5][47] ), .A6(\mem_r[6][47] ), .A7(\mem_r[7][47] ), .Z(dout_i[47]));
Q_MX08 U1778 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][48] ), .A1(\mem_r[1][48] ), .A2(\mem_r[2][48] ), .A3(\mem_r[3][48] ), .A4(\mem_r[4][48] ), .A5(\mem_r[5][48] ), .A6(\mem_r[6][48] ), .A7(\mem_r[7][48] ), .Z(dout_i[48]));
Q_MX08 U1779 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][49] ), .A1(\mem_r[1][49] ), .A2(\mem_r[2][49] ), .A3(\mem_r[3][49] ), .A4(\mem_r[4][49] ), .A5(\mem_r[5][49] ), .A6(\mem_r[6][49] ), .A7(\mem_r[7][49] ), .Z(dout_i[49]));
Q_MX08 U1780 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][50] ), .A1(\mem_r[1][50] ), .A2(\mem_r[2][50] ), .A3(\mem_r[3][50] ), .A4(\mem_r[4][50] ), .A5(\mem_r[5][50] ), .A6(\mem_r[6][50] ), .A7(\mem_r[7][50] ), .Z(dout_i[50]));
Q_MX08 U1781 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][51] ), .A1(\mem_r[1][51] ), .A2(\mem_r[2][51] ), .A3(\mem_r[3][51] ), .A4(\mem_r[4][51] ), .A5(\mem_r[5][51] ), .A6(\mem_r[6][51] ), .A7(\mem_r[7][51] ), .Z(dout_i[51]));
Q_MX08 U1782 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][52] ), .A1(\mem_r[1][52] ), .A2(\mem_r[2][52] ), .A3(\mem_r[3][52] ), .A4(\mem_r[4][52] ), .A5(\mem_r[5][52] ), .A6(\mem_r[6][52] ), .A7(\mem_r[7][52] ), .Z(dout_i[52]));
Q_MX08 U1783 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][53] ), .A1(\mem_r[1][53] ), .A2(\mem_r[2][53] ), .A3(\mem_r[3][53] ), .A4(\mem_r[4][53] ), .A5(\mem_r[5][53] ), .A6(\mem_r[6][53] ), .A7(\mem_r[7][53] ), .Z(dout_i[53]));
Q_MX08 U1784 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][54] ), .A1(\mem_r[1][54] ), .A2(\mem_r[2][54] ), .A3(\mem_r[3][54] ), .A4(\mem_r[4][54] ), .A5(\mem_r[5][54] ), .A6(\mem_r[6][54] ), .A7(\mem_r[7][54] ), .Z(dout_i[54]));
Q_MX08 U1785 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][55] ), .A1(\mem_r[1][55] ), .A2(\mem_r[2][55] ), .A3(\mem_r[3][55] ), .A4(\mem_r[4][55] ), .A5(\mem_r[5][55] ), .A6(\mem_r[6][55] ), .A7(\mem_r[7][55] ), .Z(dout_i[55]));
Q_MX08 U1786 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][56] ), .A1(\mem_r[1][56] ), .A2(\mem_r[2][56] ), .A3(\mem_r[3][56] ), .A4(\mem_r[4][56] ), .A5(\mem_r[5][56] ), .A6(\mem_r[6][56] ), .A7(\mem_r[7][56] ), .Z(dout_i[56]));
Q_MX08 U1787 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][57] ), .A1(\mem_r[1][57] ), .A2(\mem_r[2][57] ), .A3(\mem_r[3][57] ), .A4(\mem_r[4][57] ), .A5(\mem_r[5][57] ), .A6(\mem_r[6][57] ), .A7(\mem_r[7][57] ), .Z(dout_i[57]));
Q_MX08 U1788 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][58] ), .A1(\mem_r[1][58] ), .A2(\mem_r[2][58] ), .A3(\mem_r[3][58] ), .A4(\mem_r[4][58] ), .A5(\mem_r[5][58] ), .A6(\mem_r[6][58] ), .A7(\mem_r[7][58] ), .Z(dout_i[58]));
Q_MX08 U1789 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][59] ), .A1(\mem_r[1][59] ), .A2(\mem_r[2][59] ), .A3(\mem_r[3][59] ), .A4(\mem_r[4][59] ), .A5(\mem_r[5][59] ), .A6(\mem_r[6][59] ), .A7(\mem_r[7][59] ), .Z(dout_i[59]));
Q_MX08 U1790 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][60] ), .A1(\mem_r[1][60] ), .A2(\mem_r[2][60] ), .A3(\mem_r[3][60] ), .A4(\mem_r[4][60] ), .A5(\mem_r[5][60] ), .A6(\mem_r[6][60] ), .A7(\mem_r[7][60] ), .Z(dout_i[60]));
Q_MX08 U1791 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][61] ), .A1(\mem_r[1][61] ), .A2(\mem_r[2][61] ), .A3(\mem_r[3][61] ), .A4(\mem_r[4][61] ), .A5(\mem_r[5][61] ), .A6(\mem_r[6][61] ), .A7(\mem_r[7][61] ), .Z(dout_i[61]));
Q_MX08 U1792 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][62] ), .A1(\mem_r[1][62] ), .A2(\mem_r[2][62] ), .A3(\mem_r[3][62] ), .A4(\mem_r[4][62] ), .A5(\mem_r[5][62] ), .A6(\mem_r[6][62] ), .A7(\mem_r[7][62] ), .Z(dout_i[62]));
Q_MX08 U1793 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][63] ), .A1(\mem_r[1][63] ), .A2(\mem_r[2][63] ), .A3(\mem_r[3][63] ), .A4(\mem_r[4][63] ), .A5(\mem_r[5][63] ), .A6(\mem_r[6][63] ), .A7(\mem_r[7][63] ), .Z(dout_i[63]));
Q_MX08 U1794 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][64] ), .A1(\mem_r[1][64] ), .A2(\mem_r[2][64] ), .A3(\mem_r[3][64] ), .A4(\mem_r[4][64] ), .A5(\mem_r[5][64] ), .A6(\mem_r[6][64] ), .A7(\mem_r[7][64] ), .Z(dout_i[64]));
Q_MX08 U1795 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][65] ), .A1(\mem_r[1][65] ), .A2(\mem_r[2][65] ), .A3(\mem_r[3][65] ), .A4(\mem_r[4][65] ), .A5(\mem_r[5][65] ), .A6(\mem_r[6][65] ), .A7(\mem_r[7][65] ), .Z(dout_i[65]));
Q_MX08 U1796 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][66] ), .A1(\mem_r[1][66] ), .A2(\mem_r[2][66] ), .A3(\mem_r[3][66] ), .A4(\mem_r[4][66] ), .A5(\mem_r[5][66] ), .A6(\mem_r[6][66] ), .A7(\mem_r[7][66] ), .Z(dout_i[66]));
Q_MX08 U1797 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][67] ), .A1(\mem_r[1][67] ), .A2(\mem_r[2][67] ), .A3(\mem_r[3][67] ), .A4(\mem_r[4][67] ), .A5(\mem_r[5][67] ), .A6(\mem_r[6][67] ), .A7(\mem_r[7][67] ), .Z(dout_i[67]));
Q_MX08 U1798 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][68] ), .A1(\mem_r[1][68] ), .A2(\mem_r[2][68] ), .A3(\mem_r[3][68] ), .A4(\mem_r[4][68] ), .A5(\mem_r[5][68] ), .A6(\mem_r[6][68] ), .A7(\mem_r[7][68] ), .Z(dout_i[68]));
Q_MX08 U1799 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][69] ), .A1(\mem_r[1][69] ), .A2(\mem_r[2][69] ), .A3(\mem_r[3][69] ), .A4(\mem_r[4][69] ), .A5(\mem_r[5][69] ), .A6(\mem_r[6][69] ), .A7(\mem_r[7][69] ), .Z(dout_i[69]));
Q_MX08 U1800 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][70] ), .A1(\mem_r[1][70] ), .A2(\mem_r[2][70] ), .A3(\mem_r[3][70] ), .A4(\mem_r[4][70] ), .A5(\mem_r[5][70] ), .A6(\mem_r[6][70] ), .A7(\mem_r[7][70] ), .Z(dout_i[70]));
Q_MX08 U1801 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][71] ), .A1(\mem_r[1][71] ), .A2(\mem_r[2][71] ), .A3(\mem_r[3][71] ), .A4(\mem_r[4][71] ), .A5(\mem_r[5][71] ), .A6(\mem_r[6][71] ), .A7(\mem_r[7][71] ), .Z(dout_i[71]));
Q_MX08 U1802 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][72] ), .A1(\mem_r[1][72] ), .A2(\mem_r[2][72] ), .A3(\mem_r[3][72] ), .A4(\mem_r[4][72] ), .A5(\mem_r[5][72] ), .A6(\mem_r[6][72] ), .A7(\mem_r[7][72] ), .Z(dout_i[72]));
Q_MX08 U1803 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][73] ), .A1(\mem_r[1][73] ), .A2(\mem_r[2][73] ), .A3(\mem_r[3][73] ), .A4(\mem_r[4][73] ), .A5(\mem_r[5][73] ), .A6(\mem_r[6][73] ), .A7(\mem_r[7][73] ), .Z(dout_i[73]));
Q_MX08 U1804 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][74] ), .A1(\mem_r[1][74] ), .A2(\mem_r[2][74] ), .A3(\mem_r[3][74] ), .A4(\mem_r[4][74] ), .A5(\mem_r[5][74] ), .A6(\mem_r[6][74] ), .A7(\mem_r[7][74] ), .Z(dout_i[74]));
Q_MX08 U1805 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][75] ), .A1(\mem_r[1][75] ), .A2(\mem_r[2][75] ), .A3(\mem_r[3][75] ), .A4(\mem_r[4][75] ), .A5(\mem_r[5][75] ), .A6(\mem_r[6][75] ), .A7(\mem_r[7][75] ), .Z(dout_i[75]));
Q_MX08 U1806 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][76] ), .A1(\mem_r[1][76] ), .A2(\mem_r[2][76] ), .A3(\mem_r[3][76] ), .A4(\mem_r[4][76] ), .A5(\mem_r[5][76] ), .A6(\mem_r[6][76] ), .A7(\mem_r[7][76] ), .Z(dout_i[76]));
Q_MX08 U1807 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][77] ), .A1(\mem_r[1][77] ), .A2(\mem_r[2][77] ), .A3(\mem_r[3][77] ), .A4(\mem_r[4][77] ), .A5(\mem_r[5][77] ), .A6(\mem_r[6][77] ), .A7(\mem_r[7][77] ), .Z(dout_i[77]));
Q_MX08 U1808 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][78] ), .A1(\mem_r[1][78] ), .A2(\mem_r[2][78] ), .A3(\mem_r[3][78] ), .A4(\mem_r[4][78] ), .A5(\mem_r[5][78] ), .A6(\mem_r[6][78] ), .A7(\mem_r[7][78] ), .Z(dout_i[78]));
Q_MX08 U1809 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][79] ), .A1(\mem_r[1][79] ), .A2(\mem_r[2][79] ), .A3(\mem_r[3][79] ), .A4(\mem_r[4][79] ), .A5(\mem_r[5][79] ), .A6(\mem_r[6][79] ), .A7(\mem_r[7][79] ), .Z(dout_i[79]));
Q_MX08 U1810 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][80] ), .A1(\mem_r[1][80] ), .A2(\mem_r[2][80] ), .A3(\mem_r[3][80] ), .A4(\mem_r[4][80] ), .A5(\mem_r[5][80] ), .A6(\mem_r[6][80] ), .A7(\mem_r[7][80] ), .Z(dout_i[80]));
Q_MX08 U1811 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][81] ), .A1(\mem_r[1][81] ), .A2(\mem_r[2][81] ), .A3(\mem_r[3][81] ), .A4(\mem_r[4][81] ), .A5(\mem_r[5][81] ), .A6(\mem_r[6][81] ), .A7(\mem_r[7][81] ), .Z(dout_i[81]));
Q_MX08 U1812 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][82] ), .A1(\mem_r[1][82] ), .A2(\mem_r[2][82] ), .A3(\mem_r[3][82] ), .A4(\mem_r[4][82] ), .A5(\mem_r[5][82] ), .A6(\mem_r[6][82] ), .A7(\mem_r[7][82] ), .Z(dout_i[82]));
Q_MX08 U1813 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][83] ), .A1(\mem_r[1][83] ), .A2(\mem_r[2][83] ), .A3(\mem_r[3][83] ), .A4(\mem_r[4][83] ), .A5(\mem_r[5][83] ), .A6(\mem_r[6][83] ), .A7(\mem_r[7][83] ), .Z(dout_i[83]));
Q_MX08 U1814 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][84] ), .A1(\mem_r[1][84] ), .A2(\mem_r[2][84] ), .A3(\mem_r[3][84] ), .A4(\mem_r[4][84] ), .A5(\mem_r[5][84] ), .A6(\mem_r[6][84] ), .A7(\mem_r[7][84] ), .Z(dout_i[84]));
Q_MX08 U1815 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][85] ), .A1(\mem_r[1][85] ), .A2(\mem_r[2][85] ), .A3(\mem_r[3][85] ), .A4(\mem_r[4][85] ), .A5(\mem_r[5][85] ), .A6(\mem_r[6][85] ), .A7(\mem_r[7][85] ), .Z(dout_i[85]));
Q_MX08 U1816 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][86] ), .A1(\mem_r[1][86] ), .A2(\mem_r[2][86] ), .A3(\mem_r[3][86] ), .A4(\mem_r[4][86] ), .A5(\mem_r[5][86] ), .A6(\mem_r[6][86] ), .A7(\mem_r[7][86] ), .Z(dout_i[86]));
Q_MX08 U1817 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][87] ), .A1(\mem_r[1][87] ), .A2(\mem_r[2][87] ), .A3(\mem_r[3][87] ), .A4(\mem_r[4][87] ), .A5(\mem_r[5][87] ), .A6(\mem_r[6][87] ), .A7(\mem_r[7][87] ), .Z(dout_i[87]));
Q_MX08 U1818 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][88] ), .A1(\mem_r[1][88] ), .A2(\mem_r[2][88] ), .A3(\mem_r[3][88] ), .A4(\mem_r[4][88] ), .A5(\mem_r[5][88] ), .A6(\mem_r[6][88] ), .A7(\mem_r[7][88] ), .Z(dout_i[88]));
Q_MX08 U1819 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][89] ), .A1(\mem_r[1][89] ), .A2(\mem_r[2][89] ), .A3(\mem_r[3][89] ), .A4(\mem_r[4][89] ), .A5(\mem_r[5][89] ), .A6(\mem_r[6][89] ), .A7(\mem_r[7][89] ), .Z(dout_i[89]));
Q_MX08 U1820 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][90] ), .A1(\mem_r[1][90] ), .A2(\mem_r[2][90] ), .A3(\mem_r[3][90] ), .A4(\mem_r[4][90] ), .A5(\mem_r[5][90] ), .A6(\mem_r[6][90] ), .A7(\mem_r[7][90] ), .Z(dout_i[90]));
Q_MX08 U1821 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][91] ), .A1(\mem_r[1][91] ), .A2(\mem_r[2][91] ), .A3(\mem_r[3][91] ), .A4(\mem_r[4][91] ), .A5(\mem_r[5][91] ), .A6(\mem_r[6][91] ), .A7(\mem_r[7][91] ), .Z(dout_i[91]));
Q_MX08 U1822 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][92] ), .A1(\mem_r[1][92] ), .A2(\mem_r[2][92] ), .A3(\mem_r[3][92] ), .A4(\mem_r[4][92] ), .A5(\mem_r[5][92] ), .A6(\mem_r[6][92] ), .A7(\mem_r[7][92] ), .Z(dout_i[92]));
Q_MX08 U1823 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][93] ), .A1(\mem_r[1][93] ), .A2(\mem_r[2][93] ), .A3(\mem_r[3][93] ), .A4(\mem_r[4][93] ), .A5(\mem_r[5][93] ), .A6(\mem_r[6][93] ), .A7(\mem_r[7][93] ), .Z(dout_i[93]));
Q_MX08 U1824 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][94] ), .A1(\mem_r[1][94] ), .A2(\mem_r[2][94] ), .A3(\mem_r[3][94] ), .A4(\mem_r[4][94] ), .A5(\mem_r[5][94] ), .A6(\mem_r[6][94] ), .A7(\mem_r[7][94] ), .Z(dout_i[94]));
Q_MX08 U1825 ( .S0(rd_ptr_r[0]), .S1(rd_ptr_r[1]), .S2(rd_ptr_r[2]), .A0(\mem_r[0][95] ), .A1(\mem_r[1][95] ), .A2(\mem_r[2][95] ), .A3(\mem_r[3][95] ), .A4(\mem_r[4][95] ), .A5(\mem_r[5][95] ), .A6(\mem_r[6][95] ), .A7(\mem_r[7][95] ), .Z(dout_i[95]));
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m1 "mem_nxt 1 95 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m2 "mem_r 1 95 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_NON_CMM "2"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_1 "-1 GEN_NO_RD_REG_MODE  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_0 "-1 genblk1  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "GEN_NO_RD_REG_MODE"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "genblk1"
endmodule
