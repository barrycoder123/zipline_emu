
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
`_2_ (* upf_always_on = 1 *) 
module ixc_context_write_1024 ( wdata);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
input [1023:0] wdata;
wire fclk;
wire writePending;
`_2_ wire [1024:0] wdataD;
`_2_ wire [0:0] header;
`_2_ wire [0:0] headerP;
supply0 n4;
supply1 n5;
Q_NOT_TOUCH _zzqnthw ( .sig());
ixc_rforce_1024 _zzfrcD ( wdata[1023:0], wdataD[1024:1], n6);
Q_AN02 U2 ( .A0(writePending), .A1(xc_top.callEmuPre), .Z(n6));
Q_XOR2 U3 ( .A0(header[0]), .A1(headerP[0]), .Z(writePending));
Q_LDN0 \header_REG[0] ( .G(xc_top.hotSwapOnPI), .D(wdataD[0]), .Q(header[0]), .QN( ));
Q_FDP0UA U5 ( .D(n2), .QTFCLK( ), .Q(headerP[0]));
Q_MX02 U6 ( .S(n6), .A0(headerP[0]), .A1(header[0]), .Z(n2));
`ifdef CBV

reg [511:0] _zymem [0:2];
initial begin: U7
  integer i;
  for (i=0; i<=2; i=i+1) _zymem[i] =
`ifdef CBV_MEM_INIT1
  {512{1'b1}};
`else
  512'b0;
`endif
end
reg [511:0] n10;
assign {wdataD[511], wdataD[510], wdataD[509], wdataD[508], wdataD[507], wdataD[506], wdataD[505],
wdataD[504], wdataD[503], wdataD[502], wdataD[501], wdataD[500], wdataD[499], wdataD[498], wdataD[497],
wdataD[496], wdataD[495], wdataD[494], wdataD[493], wdataD[492], wdataD[491], wdataD[490], wdataD[489],
wdataD[488], wdataD[487], wdataD[486], wdataD[485], wdataD[484], wdataD[483], wdataD[482], wdataD[481],
wdataD[480], wdataD[479], wdataD[478], wdataD[477], wdataD[476], wdataD[475], wdataD[474], wdataD[473],
wdataD[472], wdataD[471], wdataD[470], wdataD[469], wdataD[468], wdataD[467], wdataD[466], wdataD[465],
wdataD[464], wdataD[463], wdataD[462], wdataD[461], wdataD[460], wdataD[459], wdataD[458], wdataD[457],
wdataD[456], wdataD[455], wdataD[454], wdataD[453], wdataD[452], wdataD[451], wdataD[450], wdataD[449],
wdataD[448], wdataD[447], wdataD[446], wdataD[445], wdataD[444], wdataD[443], wdataD[442], wdataD[441],
wdataD[440], wdataD[439], wdataD[438], wdataD[437], wdataD[436], wdataD[435], wdataD[434], wdataD[433],
wdataD[432], wdataD[431], wdataD[430], wdataD[429], wdataD[428], wdataD[427], wdataD[426], wdataD[425],
wdataD[424], wdataD[423], wdataD[422], wdataD[421], wdataD[420], wdataD[419], wdataD[418], wdataD[417],
wdataD[416], wdataD[415], wdataD[414], wdataD[413], wdataD[412], wdataD[411], wdataD[410], wdataD[409],
wdataD[408], wdataD[407], wdataD[406], wdataD[405], wdataD[404], wdataD[403], wdataD[402], wdataD[401],
wdataD[400], wdataD[399], wdataD[398], wdataD[397], wdataD[396], wdataD[395], wdataD[394], wdataD[393],
wdataD[392], wdataD[391], wdataD[390], wdataD[389], wdataD[388], wdataD[387], wdataD[386], wdataD[385],
wdataD[384], wdataD[383], wdataD[382], wdataD[381], wdataD[380], wdataD[379], wdataD[378], wdataD[377],
wdataD[376], wdataD[375], wdataD[374], wdataD[373], wdataD[372], wdataD[371], wdataD[370], wdataD[369],
wdataD[368], wdataD[367], wdataD[366], wdataD[365], wdataD[364], wdataD[363], wdataD[362], wdataD[361],
wdataD[360], wdataD[359], wdataD[358], wdataD[357], wdataD[356], wdataD[355], wdataD[354], wdataD[353],
wdataD[352], wdataD[351], wdataD[350], wdataD[349], wdataD[348], wdataD[347], wdataD[346], wdataD[345],
wdataD[344], wdataD[343], wdataD[342], wdataD[341], wdataD[340], wdataD[339], wdataD[338], wdataD[337],
wdataD[336], wdataD[335], wdataD[334], wdataD[333], wdataD[332], wdataD[331], wdataD[330], wdataD[329],
wdataD[328], wdataD[327], wdataD[326], wdataD[325], wdataD[324], wdataD[323], wdataD[322], wdataD[321],
wdataD[320], wdataD[319], wdataD[318], wdataD[317], wdataD[316], wdataD[315], wdataD[314], wdataD[313],
wdataD[312], wdataD[311], wdataD[310], wdataD[309], wdataD[308], wdataD[307], wdataD[306], wdataD[305],
wdataD[304], wdataD[303], wdataD[302], wdataD[301], wdataD[300], wdataD[299], wdataD[298], wdataD[297],
wdataD[296], wdataD[295], wdataD[294], wdataD[293], wdataD[292], wdataD[291], wdataD[290], wdataD[289],
wdataD[288], wdataD[287], wdataD[286], wdataD[285], wdataD[284], wdataD[283], wdataD[282], wdataD[281],
wdataD[280], wdataD[279], wdataD[278], wdataD[277], wdataD[276], wdataD[275], wdataD[274], wdataD[273],
wdataD[272], wdataD[271], wdataD[270], wdataD[269], wdataD[268], wdataD[267], wdataD[266], wdataD[265],
wdataD[264], wdataD[263], wdataD[262], wdataD[261], wdataD[260], wdataD[259], wdataD[258], wdataD[257],
wdataD[256], wdataD[255], wdataD[254], wdataD[253], wdataD[252], wdataD[251], wdataD[250], wdataD[249],
wdataD[248], wdataD[247], wdataD[246], wdataD[245], wdataD[244], wdataD[243], wdataD[242], wdataD[241],
wdataD[240], wdataD[239], wdataD[238], wdataD[237], wdataD[236], wdataD[235], wdataD[234], wdataD[233],
wdataD[232], wdataD[231], wdataD[230], wdataD[229], wdataD[228], wdataD[227], wdataD[226], wdataD[225],
wdataD[224], wdataD[223], wdataD[222], wdataD[221], wdataD[220], wdataD[219], wdataD[218], wdataD[217],
wdataD[216], wdataD[215], wdataD[214], wdataD[213], wdataD[212], wdataD[211], wdataD[210], wdataD[209],
wdataD[208], wdataD[207], wdataD[206], wdataD[205], wdataD[204], wdataD[203], wdataD[202], wdataD[201],
wdataD[200], wdataD[199], wdataD[198], wdataD[197], wdataD[196], wdataD[195], wdataD[194], wdataD[193],
wdataD[192], wdataD[191], wdataD[190], wdataD[189], wdataD[188], wdataD[187], wdataD[186], wdataD[185],
wdataD[184], wdataD[183], wdataD[182], wdataD[181], wdataD[180], wdataD[179], wdataD[178], wdataD[177],
wdataD[176], wdataD[175], wdataD[174], wdataD[173], wdataD[172], wdataD[171], wdataD[170], wdataD[169],
wdataD[168], wdataD[167], wdataD[166], wdataD[165], wdataD[164], wdataD[163], wdataD[162], wdataD[161],
wdataD[160], wdataD[159], wdataD[158], wdataD[157], wdataD[156], wdataD[155], wdataD[154], wdataD[153],
wdataD[152], wdataD[151], wdataD[150], wdataD[149], wdataD[148], wdataD[147], wdataD[146], wdataD[145],
wdataD[144], wdataD[143], wdataD[142], wdataD[141], wdataD[140], wdataD[139], wdataD[138], wdataD[137],
wdataD[136], wdataD[135], wdataD[134], wdataD[133], wdataD[132], wdataD[131], wdataD[130], wdataD[129],
wdataD[128], wdataD[127], wdataD[126], wdataD[125], wdataD[124], wdataD[123], wdataD[122], wdataD[121],
wdataD[120], wdataD[119], wdataD[118], wdataD[117], wdataD[116], wdataD[115], wdataD[114], wdataD[113],
wdataD[112], wdataD[111], wdataD[110], wdataD[109], wdataD[108], wdataD[107], wdataD[106], wdataD[105],
wdataD[104], wdataD[103], wdataD[102], wdataD[101], wdataD[100], wdataD[99], wdataD[98], wdataD[97],
wdataD[96], wdataD[95], wdataD[94], wdataD[93], wdataD[92], wdataD[91], wdataD[90], wdataD[89],
wdataD[88], wdataD[87], wdataD[86], wdataD[85], wdataD[84], wdataD[83], wdataD[82], wdataD[81],
wdataD[80], wdataD[79], wdataD[78], wdataD[77], wdataD[76], wdataD[75], wdataD[74], wdataD[73],
wdataD[72], wdataD[71], wdataD[70], wdataD[69], wdataD[68], wdataD[67], wdataD[66], wdataD[65],
wdataD[64], wdataD[63], wdataD[62], wdataD[61], wdataD[60], wdataD[59], wdataD[58], wdataD[57],
wdataD[56], wdataD[55], wdataD[54], wdataD[53], wdataD[52], wdataD[51], wdataD[50], wdataD[49],
wdataD[48], wdataD[47], wdataD[46], wdataD[45], wdataD[44], wdataD[43], wdataD[42], wdataD[41],
wdataD[40], wdataD[39], wdataD[38], wdataD[37], wdataD[36], wdataD[35], wdataD[34], wdataD[33],
wdataD[32], wdataD[31], wdataD[30], wdataD[29], wdataD[28], wdataD[27], wdataD[26], wdataD[25],
wdataD[24], wdataD[23], wdataD[22], wdataD[21], wdataD[20], wdataD[19], wdataD[18], wdataD[17],
wdataD[16], wdataD[15], wdataD[14], wdataD[13], wdataD[12], wdataD[11], wdataD[10], wdataD[9],
wdataD[8], wdataD[7], wdataD[6], wdataD[5], wdataD[4], wdataD[3], wdataD[2], wdataD[1],
wdataD[0]} = n10; 
reg [511:0] n8;
assign {wdataD[1023], wdataD[1022], wdataD[1021], wdataD[1020], wdataD[1019], wdataD[1018], wdataD[1017],
wdataD[1016], wdataD[1015], wdataD[1014], wdataD[1013], wdataD[1012], wdataD[1011], wdataD[1010], wdataD[1009],
wdataD[1008], wdataD[1007], wdataD[1006], wdataD[1005], wdataD[1004], wdataD[1003], wdataD[1002], wdataD[1001],
wdataD[1000], wdataD[999], wdataD[998], wdataD[997], wdataD[996], wdataD[995], wdataD[994], wdataD[993],
wdataD[992], wdataD[991], wdataD[990], wdataD[989], wdataD[988], wdataD[987], wdataD[986], wdataD[985],
wdataD[984], wdataD[983], wdataD[982], wdataD[981], wdataD[980], wdataD[979], wdataD[978], wdataD[977],
wdataD[976], wdataD[975], wdataD[974], wdataD[973], wdataD[972], wdataD[971], wdataD[970], wdataD[969],
wdataD[968], wdataD[967], wdataD[966], wdataD[965], wdataD[964], wdataD[963], wdataD[962], wdataD[961],
wdataD[960], wdataD[959], wdataD[958], wdataD[957], wdataD[956], wdataD[955], wdataD[954], wdataD[953],
wdataD[952], wdataD[951], wdataD[950], wdataD[949], wdataD[948], wdataD[947], wdataD[946], wdataD[945],
wdataD[944], wdataD[943], wdataD[942], wdataD[941], wdataD[940], wdataD[939], wdataD[938], wdataD[937],
wdataD[936], wdataD[935], wdataD[934], wdataD[933], wdataD[932], wdataD[931], wdataD[930], wdataD[929],
wdataD[928], wdataD[927], wdataD[926], wdataD[925], wdataD[924], wdataD[923], wdataD[922], wdataD[921],
wdataD[920], wdataD[919], wdataD[918], wdataD[917], wdataD[916], wdataD[915], wdataD[914], wdataD[913],
wdataD[912], wdataD[911], wdataD[910], wdataD[909], wdataD[908], wdataD[907], wdataD[906], wdataD[905],
wdataD[904], wdataD[903], wdataD[902], wdataD[901], wdataD[900], wdataD[899], wdataD[898], wdataD[897],
wdataD[896], wdataD[895], wdataD[894], wdataD[893], wdataD[892], wdataD[891], wdataD[890], wdataD[889],
wdataD[888], wdataD[887], wdataD[886], wdataD[885], wdataD[884], wdataD[883], wdataD[882], wdataD[881],
wdataD[880], wdataD[879], wdataD[878], wdataD[877], wdataD[876], wdataD[875], wdataD[874], wdataD[873],
wdataD[872], wdataD[871], wdataD[870], wdataD[869], wdataD[868], wdataD[867], wdataD[866], wdataD[865],
wdataD[864], wdataD[863], wdataD[862], wdataD[861], wdataD[860], wdataD[859], wdataD[858], wdataD[857],
wdataD[856], wdataD[855], wdataD[854], wdataD[853], wdataD[852], wdataD[851], wdataD[850], wdataD[849],
wdataD[848], wdataD[847], wdataD[846], wdataD[845], wdataD[844], wdataD[843], wdataD[842], wdataD[841],
wdataD[840], wdataD[839], wdataD[838], wdataD[837], wdataD[836], wdataD[835], wdataD[834], wdataD[833],
wdataD[832], wdataD[831], wdataD[830], wdataD[829], wdataD[828], wdataD[827], wdataD[826], wdataD[825],
wdataD[824], wdataD[823], wdataD[822], wdataD[821], wdataD[820], wdataD[819], wdataD[818], wdataD[817],
wdataD[816], wdataD[815], wdataD[814], wdataD[813], wdataD[812], wdataD[811], wdataD[810], wdataD[809],
wdataD[808], wdataD[807], wdataD[806], wdataD[805], wdataD[804], wdataD[803], wdataD[802], wdataD[801],
wdataD[800], wdataD[799], wdataD[798], wdataD[797], wdataD[796], wdataD[795], wdataD[794], wdataD[793],
wdataD[792], wdataD[791], wdataD[790], wdataD[789], wdataD[788], wdataD[787], wdataD[786], wdataD[785],
wdataD[784], wdataD[783], wdataD[782], wdataD[781], wdataD[780], wdataD[779], wdataD[778], wdataD[777],
wdataD[776], wdataD[775], wdataD[774], wdataD[773], wdataD[772], wdataD[771], wdataD[770], wdataD[769],
wdataD[768], wdataD[767], wdataD[766], wdataD[765], wdataD[764], wdataD[763], wdataD[762], wdataD[761],
wdataD[760], wdataD[759], wdataD[758], wdataD[757], wdataD[756], wdataD[755], wdataD[754], wdataD[753],
wdataD[752], wdataD[751], wdataD[750], wdataD[749], wdataD[748], wdataD[747], wdataD[746], wdataD[745],
wdataD[744], wdataD[743], wdataD[742], wdataD[741], wdataD[740], wdataD[739], wdataD[738], wdataD[737],
wdataD[736], wdataD[735], wdataD[734], wdataD[733], wdataD[732], wdataD[731], wdataD[730], wdataD[729],
wdataD[728], wdataD[727], wdataD[726], wdataD[725], wdataD[724], wdataD[723], wdataD[722], wdataD[721],
wdataD[720], wdataD[719], wdataD[718], wdataD[717], wdataD[716], wdataD[715], wdataD[714], wdataD[713],
wdataD[712], wdataD[711], wdataD[710], wdataD[709], wdataD[708], wdataD[707], wdataD[706], wdataD[705],
wdataD[704], wdataD[703], wdataD[702], wdataD[701], wdataD[700], wdataD[699], wdataD[698], wdataD[697],
wdataD[696], wdataD[695], wdataD[694], wdataD[693], wdataD[692], wdataD[691], wdataD[690], wdataD[689],
wdataD[688], wdataD[687], wdataD[686], wdataD[685], wdataD[684], wdataD[683], wdataD[682], wdataD[681],
wdataD[680], wdataD[679], wdataD[678], wdataD[677], wdataD[676], wdataD[675], wdataD[674], wdataD[673],
wdataD[672], wdataD[671], wdataD[670], wdataD[669], wdataD[668], wdataD[667], wdataD[666], wdataD[665],
wdataD[664], wdataD[663], wdataD[662], wdataD[661], wdataD[660], wdataD[659], wdataD[658], wdataD[657],
wdataD[656], wdataD[655], wdataD[654], wdataD[653], wdataD[652], wdataD[651], wdataD[650], wdataD[649],
wdataD[648], wdataD[647], wdataD[646], wdataD[645], wdataD[644], wdataD[643], wdataD[642], wdataD[641],
wdataD[640], wdataD[639], wdataD[638], wdataD[637], wdataD[636], wdataD[635], wdataD[634], wdataD[633],
wdataD[632], wdataD[631], wdataD[630], wdataD[629], wdataD[628], wdataD[627], wdataD[626], wdataD[625],
wdataD[624], wdataD[623], wdataD[622], wdataD[621], wdataD[620], wdataD[619], wdataD[618], wdataD[617],
wdataD[616], wdataD[615], wdataD[614], wdataD[613], wdataD[612], wdataD[611], wdataD[610], wdataD[609],
wdataD[608], wdataD[607], wdataD[606], wdataD[605], wdataD[604], wdataD[603], wdataD[602], wdataD[601],
wdataD[600], wdataD[599], wdataD[598], wdataD[597], wdataD[596], wdataD[595], wdataD[594], wdataD[593],
wdataD[592], wdataD[591], wdataD[590], wdataD[589], wdataD[588], wdataD[587], wdataD[586], wdataD[585],
wdataD[584], wdataD[583], wdataD[582], wdataD[581], wdataD[580], wdataD[579], wdataD[578], wdataD[577],
wdataD[576], wdataD[575], wdataD[574], wdataD[573], wdataD[572], wdataD[571], wdataD[570], wdataD[569],
wdataD[568], wdataD[567], wdataD[566], wdataD[565], wdataD[564], wdataD[563], wdataD[562], wdataD[561],
wdataD[560], wdataD[559], wdataD[558], wdataD[557], wdataD[556], wdataD[555], wdataD[554], wdataD[553],
wdataD[552], wdataD[551], wdataD[550], wdataD[549], wdataD[548], wdataD[547], wdataD[546], wdataD[545],
wdataD[544], wdataD[543], wdataD[542], wdataD[541], wdataD[540], wdataD[539], wdataD[538], wdataD[537],
wdataD[536], wdataD[535], wdataD[534], wdataD[533], wdataD[532], wdataD[531], wdataD[530], wdataD[529],
wdataD[528], wdataD[527], wdataD[526], wdataD[525], wdataD[524], wdataD[523], wdataD[522], wdataD[521],
wdataD[520], wdataD[519], wdataD[518], wdataD[517], wdataD[516], wdataD[515], wdataD[514], wdataD[513],
wdataD[512]} = n8; 
reg [511:0] n9;
buf(wdataD[1024], n9[0]);
always @(n4 or n5)
#0 begin
n10 = _zymem[{n4, n4}];
n8 = _zymem[{n4, n5}];
n9 = _zymem[{n5, n4}];
end
`else

MPR4X512 _zymem ( .A1(n4), .A0(n4), .SYNC_IN(n4), .DO511(wdataD[511]), .DO510(wdataD[510]), .DO509(wdataD[509]),
 .DO508(wdataD[508]), .DO507(wdataD[507]), .DO506(wdataD[506]), .DO505(wdataD[505]), .DO504(wdataD[504]), .DO503(wdataD[503]), .DO502(wdataD[502]), .DO501(wdataD[501]),
 .DO500(wdataD[500]), .DO499(wdataD[499]), .DO498(wdataD[498]), .DO497(wdataD[497]), .DO496(wdataD[496]), .DO495(wdataD[495]), .DO494(wdataD[494]), .DO493(wdataD[493]),
 .DO492(wdataD[492]), .DO491(wdataD[491]), .DO490(wdataD[490]), .DO489(wdataD[489]), .DO488(wdataD[488]), .DO487(wdataD[487]), .DO486(wdataD[486]), .DO485(wdataD[485]),
 .DO484(wdataD[484]), .DO483(wdataD[483]), .DO482(wdataD[482]), .DO481(wdataD[481]), .DO480(wdataD[480]), .DO479(wdataD[479]), .DO478(wdataD[478]), .DO477(wdataD[477]),
 .DO476(wdataD[476]), .DO475(wdataD[475]), .DO474(wdataD[474]), .DO473(wdataD[473]), .DO472(wdataD[472]), .DO471(wdataD[471]), .DO470(wdataD[470]), .DO469(wdataD[469]),
 .DO468(wdataD[468]), .DO467(wdataD[467]), .DO466(wdataD[466]), .DO465(wdataD[465]), .DO464(wdataD[464]), .DO463(wdataD[463]), .DO462(wdataD[462]), .DO461(wdataD[461]),
 .DO460(wdataD[460]), .DO459(wdataD[459]), .DO458(wdataD[458]), .DO457(wdataD[457]), .DO456(wdataD[456]), .DO455(wdataD[455]), .DO454(wdataD[454]), .DO453(wdataD[453]),
 .DO452(wdataD[452]), .DO451(wdataD[451]), .DO450(wdataD[450]), .DO449(wdataD[449]), .DO448(wdataD[448]), .DO447(wdataD[447]), .DO446(wdataD[446]), .DO445(wdataD[445]),
 .DO444(wdataD[444]), .DO443(wdataD[443]), .DO442(wdataD[442]), .DO441(wdataD[441]), .DO440(wdataD[440]), .DO439(wdataD[439]), .DO438(wdataD[438]), .DO437(wdataD[437]),
 .DO436(wdataD[436]), .DO435(wdataD[435]), .DO434(wdataD[434]), .DO433(wdataD[433]), .DO432(wdataD[432]), .DO431(wdataD[431]), .DO430(wdataD[430]), .DO429(wdataD[429]),
 .DO428(wdataD[428]), .DO427(wdataD[427]), .DO426(wdataD[426]), .DO425(wdataD[425]), .DO424(wdataD[424]), .DO423(wdataD[423]), .DO422(wdataD[422]), .DO421(wdataD[421]),
 .DO420(wdataD[420]), .DO419(wdataD[419]), .DO418(wdataD[418]), .DO417(wdataD[417]), .DO416(wdataD[416]), .DO415(wdataD[415]), .DO414(wdataD[414]), .DO413(wdataD[413]),
 .DO412(wdataD[412]), .DO411(wdataD[411]), .DO410(wdataD[410]), .DO409(wdataD[409]), .DO408(wdataD[408]), .DO407(wdataD[407]), .DO406(wdataD[406]), .DO405(wdataD[405]),
 .DO404(wdataD[404]), .DO403(wdataD[403]), .DO402(wdataD[402]), .DO401(wdataD[401]), .DO400(wdataD[400]), .DO399(wdataD[399]), .DO398(wdataD[398]), .DO397(wdataD[397]),
 .DO396(wdataD[396]), .DO395(wdataD[395]), .DO394(wdataD[394]), .DO393(wdataD[393]), .DO392(wdataD[392]), .DO391(wdataD[391]), .DO390(wdataD[390]), .DO389(wdataD[389]),
 .DO388(wdataD[388]), .DO387(wdataD[387]), .DO386(wdataD[386]), .DO385(wdataD[385]), .DO384(wdataD[384]), .DO383(wdataD[383]), .DO382(wdataD[382]), .DO381(wdataD[381]),
 .DO380(wdataD[380]), .DO379(wdataD[379]), .DO378(wdataD[378]), .DO377(wdataD[377]), .DO376(wdataD[376]), .DO375(wdataD[375]), .DO374(wdataD[374]), .DO373(wdataD[373]),
 .DO372(wdataD[372]), .DO371(wdataD[371]), .DO370(wdataD[370]), .DO369(wdataD[369]), .DO368(wdataD[368]), .DO367(wdataD[367]), .DO366(wdataD[366]), .DO365(wdataD[365]),
 .DO364(wdataD[364]), .DO363(wdataD[363]), .DO362(wdataD[362]), .DO361(wdataD[361]), .DO360(wdataD[360]), .DO359(wdataD[359]), .DO358(wdataD[358]), .DO357(wdataD[357]),
 .DO356(wdataD[356]), .DO355(wdataD[355]), .DO354(wdataD[354]), .DO353(wdataD[353]), .DO352(wdataD[352]), .DO351(wdataD[351]), .DO350(wdataD[350]), .DO349(wdataD[349]),
 .DO348(wdataD[348]), .DO347(wdataD[347]), .DO346(wdataD[346]), .DO345(wdataD[345]), .DO344(wdataD[344]), .DO343(wdataD[343]), .DO342(wdataD[342]), .DO341(wdataD[341]),
 .DO340(wdataD[340]), .DO339(wdataD[339]), .DO338(wdataD[338]), .DO337(wdataD[337]), .DO336(wdataD[336]), .DO335(wdataD[335]), .DO334(wdataD[334]), .DO333(wdataD[333]),
 .DO332(wdataD[332]), .DO331(wdataD[331]), .DO330(wdataD[330]), .DO329(wdataD[329]), .DO328(wdataD[328]), .DO327(wdataD[327]), .DO326(wdataD[326]), .DO325(wdataD[325]),
 .DO324(wdataD[324]), .DO323(wdataD[323]), .DO322(wdataD[322]), .DO321(wdataD[321]), .DO320(wdataD[320]), .DO319(wdataD[319]), .DO318(wdataD[318]), .DO317(wdataD[317]),
 .DO316(wdataD[316]), .DO315(wdataD[315]), .DO314(wdataD[314]), .DO313(wdataD[313]), .DO312(wdataD[312]), .DO311(wdataD[311]), .DO310(wdataD[310]), .DO309(wdataD[309]),
 .DO308(wdataD[308]), .DO307(wdataD[307]), .DO306(wdataD[306]), .DO305(wdataD[305]), .DO304(wdataD[304]), .DO303(wdataD[303]), .DO302(wdataD[302]), .DO301(wdataD[301]),
 .DO300(wdataD[300]), .DO299(wdataD[299]), .DO298(wdataD[298]), .DO297(wdataD[297]), .DO296(wdataD[296]), .DO295(wdataD[295]), .DO294(wdataD[294]), .DO293(wdataD[293]),
 .DO292(wdataD[292]), .DO291(wdataD[291]), .DO290(wdataD[290]), .DO289(wdataD[289]), .DO288(wdataD[288]), .DO287(wdataD[287]), .DO286(wdataD[286]), .DO285(wdataD[285]),
 .DO284(wdataD[284]), .DO283(wdataD[283]), .DO282(wdataD[282]), .DO281(wdataD[281]), .DO280(wdataD[280]), .DO279(wdataD[279]), .DO278(wdataD[278]), .DO277(wdataD[277]),
 .DO276(wdataD[276]), .DO275(wdataD[275]), .DO274(wdataD[274]), .DO273(wdataD[273]), .DO272(wdataD[272]), .DO271(wdataD[271]), .DO270(wdataD[270]), .DO269(wdataD[269]),
 .DO268(wdataD[268]), .DO267(wdataD[267]), .DO266(wdataD[266]), .DO265(wdataD[265]), .DO264(wdataD[264]), .DO263(wdataD[263]), .DO262(wdataD[262]), .DO261(wdataD[261]),
 .DO260(wdataD[260]), .DO259(wdataD[259]), .DO258(wdataD[258]), .DO257(wdataD[257]), .DO256(wdataD[256]), .DO255(wdataD[255]), .DO254(wdataD[254]), .DO253(wdataD[253]),
 .DO252(wdataD[252]), .DO251(wdataD[251]), .DO250(wdataD[250]), .DO249(wdataD[249]), .DO248(wdataD[248]), .DO247(wdataD[247]), .DO246(wdataD[246]), .DO245(wdataD[245]),
 .DO244(wdataD[244]), .DO243(wdataD[243]), .DO242(wdataD[242]), .DO241(wdataD[241]), .DO240(wdataD[240]), .DO239(wdataD[239]), .DO238(wdataD[238]), .DO237(wdataD[237]),
 .DO236(wdataD[236]), .DO235(wdataD[235]), .DO234(wdataD[234]), .DO233(wdataD[233]), .DO232(wdataD[232]), .DO231(wdataD[231]), .DO230(wdataD[230]), .DO229(wdataD[229]),
 .DO228(wdataD[228]), .DO227(wdataD[227]), .DO226(wdataD[226]), .DO225(wdataD[225]), .DO224(wdataD[224]), .DO223(wdataD[223]), .DO222(wdataD[222]), .DO221(wdataD[221]),
 .DO220(wdataD[220]), .DO219(wdataD[219]), .DO218(wdataD[218]), .DO217(wdataD[217]), .DO216(wdataD[216]), .DO215(wdataD[215]), .DO214(wdataD[214]), .DO213(wdataD[213]),
 .DO212(wdataD[212]), .DO211(wdataD[211]), .DO210(wdataD[210]), .DO209(wdataD[209]), .DO208(wdataD[208]), .DO207(wdataD[207]), .DO206(wdataD[206]), .DO205(wdataD[205]),
 .DO204(wdataD[204]), .DO203(wdataD[203]), .DO202(wdataD[202]), .DO201(wdataD[201]), .DO200(wdataD[200]), .DO199(wdataD[199]), .DO198(wdataD[198]), .DO197(wdataD[197]),
 .DO196(wdataD[196]), .DO195(wdataD[195]), .DO194(wdataD[194]), .DO193(wdataD[193]), .DO192(wdataD[192]), .DO191(wdataD[191]), .DO190(wdataD[190]), .DO189(wdataD[189]),
 .DO188(wdataD[188]), .DO187(wdataD[187]), .DO186(wdataD[186]), .DO185(wdataD[185]), .DO184(wdataD[184]), .DO183(wdataD[183]), .DO182(wdataD[182]), .DO181(wdataD[181]),
 .DO180(wdataD[180]), .DO179(wdataD[179]), .DO178(wdataD[178]), .DO177(wdataD[177]), .DO176(wdataD[176]), .DO175(wdataD[175]), .DO174(wdataD[174]), .DO173(wdataD[173]),
 .DO172(wdataD[172]), .DO171(wdataD[171]), .DO170(wdataD[170]), .DO169(wdataD[169]), .DO168(wdataD[168]), .DO167(wdataD[167]), .DO166(wdataD[166]), .DO165(wdataD[165]),
 .DO164(wdataD[164]), .DO163(wdataD[163]), .DO162(wdataD[162]), .DO161(wdataD[161]), .DO160(wdataD[160]), .DO159(wdataD[159]), .DO158(wdataD[158]), .DO157(wdataD[157]),
 .DO156(wdataD[156]), .DO155(wdataD[155]), .DO154(wdataD[154]), .DO153(wdataD[153]), .DO152(wdataD[152]), .DO151(wdataD[151]), .DO150(wdataD[150]), .DO149(wdataD[149]),
 .DO148(wdataD[148]), .DO147(wdataD[147]), .DO146(wdataD[146]), .DO145(wdataD[145]), .DO144(wdataD[144]), .DO143(wdataD[143]), .DO142(wdataD[142]), .DO141(wdataD[141]),
 .DO140(wdataD[140]), .DO139(wdataD[139]), .DO138(wdataD[138]), .DO137(wdataD[137]), .DO136(wdataD[136]), .DO135(wdataD[135]), .DO134(wdataD[134]), .DO133(wdataD[133]),
 .DO132(wdataD[132]), .DO131(wdataD[131]), .DO130(wdataD[130]), .DO129(wdataD[129]), .DO128(wdataD[128]), .DO127(wdataD[127]), .DO126(wdataD[126]), .DO125(wdataD[125]),
 .DO124(wdataD[124]), .DO123(wdataD[123]), .DO122(wdataD[122]), .DO121(wdataD[121]), .DO120(wdataD[120]), .DO119(wdataD[119]), .DO118(wdataD[118]), .DO117(wdataD[117]),
 .DO116(wdataD[116]), .DO115(wdataD[115]), .DO114(wdataD[114]), .DO113(wdataD[113]), .DO112(wdataD[112]), .DO111(wdataD[111]), .DO110(wdataD[110]), .DO109(wdataD[109]),
 .DO108(wdataD[108]), .DO107(wdataD[107]), .DO106(wdataD[106]), .DO105(wdataD[105]), .DO104(wdataD[104]), .DO103(wdataD[103]), .DO102(wdataD[102]), .DO101(wdataD[101]),
 .DO100(wdataD[100]), .DO99(wdataD[99]), .DO98(wdataD[98]), .DO97(wdataD[97]), .DO96(wdataD[96]), .DO95(wdataD[95]), .DO94(wdataD[94]), .DO93(wdataD[93]),
 .DO92(wdataD[92]), .DO91(wdataD[91]), .DO90(wdataD[90]), .DO89(wdataD[89]), .DO88(wdataD[88]), .DO87(wdataD[87]), .DO86(wdataD[86]), .DO85(wdataD[85]),
 .DO84(wdataD[84]), .DO83(wdataD[83]), .DO82(wdataD[82]), .DO81(wdataD[81]), .DO80(wdataD[80]), .DO79(wdataD[79]), .DO78(wdataD[78]), .DO77(wdataD[77]),
 .DO76(wdataD[76]), .DO75(wdataD[75]), .DO74(wdataD[74]), .DO73(wdataD[73]), .DO72(wdataD[72]), .DO71(wdataD[71]), .DO70(wdataD[70]), .DO69(wdataD[69]),
 .DO68(wdataD[68]), .DO67(wdataD[67]), .DO66(wdataD[66]), .DO65(wdataD[65]), .DO64(wdataD[64]), .DO63(wdataD[63]), .DO62(wdataD[62]), .DO61(wdataD[61]),
 .DO60(wdataD[60]), .DO59(wdataD[59]), .DO58(wdataD[58]), .DO57(wdataD[57]), .DO56(wdataD[56]), .DO55(wdataD[55]), .DO54(wdataD[54]), .DO53(wdataD[53]),
 .DO52(wdataD[52]), .DO51(wdataD[51]), .DO50(wdataD[50]), .DO49(wdataD[49]), .DO48(wdataD[48]), .DO47(wdataD[47]), .DO46(wdataD[46]), .DO45(wdataD[45]),
 .DO44(wdataD[44]), .DO43(wdataD[43]), .DO42(wdataD[42]), .DO41(wdataD[41]), .DO40(wdataD[40]), .DO39(wdataD[39]), .DO38(wdataD[38]), .DO37(wdataD[37]),
 .DO36(wdataD[36]), .DO35(wdataD[35]), .DO34(wdataD[34]), .DO33(wdataD[33]), .DO32(wdataD[32]), .DO31(wdataD[31]), .DO30(wdataD[30]), .DO29(wdataD[29]),
 .DO28(wdataD[28]), .DO27(wdataD[27]), .DO26(wdataD[26]), .DO25(wdataD[25]), .DO24(wdataD[24]), .DO23(wdataD[23]), .DO22(wdataD[22]), .DO21(wdataD[21]),
 .DO20(wdataD[20]), .DO19(wdataD[19]), .DO18(wdataD[18]), .DO17(wdataD[17]), .DO16(wdataD[16]), .DO15(wdataD[15]), .DO14(wdataD[14]), .DO13(wdataD[13]),
 .DO12(wdataD[12]), .DO11(wdataD[11]), .DO10(wdataD[10]), .DO9(wdataD[9]), .DO8(wdataD[8]), .DO7(wdataD[7]), .DO6(wdataD[6]), .DO5(wdataD[5]),
 .DO4(wdataD[4]), .DO3(wdataD[3]), .DO2(wdataD[2]), .DO1(wdataD[1]), .DO0(wdataD[0]), .SYNC_OUT(n8));
// pragma CVASTRPROP INSTANCE "_zymem" HDL_MEMORY_DECL "1 511 0 0 2"
MPR4X512 U8 ( .A1(n4), .A0(n5), .SYNC_IN(n8), .DO511(wdataD[1023]), .DO510(wdataD[1022]), .DO509(wdataD[1021]),
 .DO508(wdataD[1020]), .DO507(wdataD[1019]), .DO506(wdataD[1018]), .DO505(wdataD[1017]), .DO504(wdataD[1016]), .DO503(wdataD[1015]), .DO502(wdataD[1014]), .DO501(wdataD[1013]),
 .DO500(wdataD[1012]), .DO499(wdataD[1011]), .DO498(wdataD[1010]), .DO497(wdataD[1009]), .DO496(wdataD[1008]), .DO495(wdataD[1007]), .DO494(wdataD[1006]), .DO493(wdataD[1005]),
 .DO492(wdataD[1004]), .DO491(wdataD[1003]), .DO490(wdataD[1002]), .DO489(wdataD[1001]), .DO488(wdataD[1000]), .DO487(wdataD[999]), .DO486(wdataD[998]), .DO485(wdataD[997]),
 .DO484(wdataD[996]), .DO483(wdataD[995]), .DO482(wdataD[994]), .DO481(wdataD[993]), .DO480(wdataD[992]), .DO479(wdataD[991]), .DO478(wdataD[990]), .DO477(wdataD[989]),
 .DO476(wdataD[988]), .DO475(wdataD[987]), .DO474(wdataD[986]), .DO473(wdataD[985]), .DO472(wdataD[984]), .DO471(wdataD[983]), .DO470(wdataD[982]), .DO469(wdataD[981]),
 .DO468(wdataD[980]), .DO467(wdataD[979]), .DO466(wdataD[978]), .DO465(wdataD[977]), .DO464(wdataD[976]), .DO463(wdataD[975]), .DO462(wdataD[974]), .DO461(wdataD[973]),
 .DO460(wdataD[972]), .DO459(wdataD[971]), .DO458(wdataD[970]), .DO457(wdataD[969]), .DO456(wdataD[968]), .DO455(wdataD[967]), .DO454(wdataD[966]), .DO453(wdataD[965]),
 .DO452(wdataD[964]), .DO451(wdataD[963]), .DO450(wdataD[962]), .DO449(wdataD[961]), .DO448(wdataD[960]), .DO447(wdataD[959]), .DO446(wdataD[958]), .DO445(wdataD[957]),
 .DO444(wdataD[956]), .DO443(wdataD[955]), .DO442(wdataD[954]), .DO441(wdataD[953]), .DO440(wdataD[952]), .DO439(wdataD[951]), .DO438(wdataD[950]), .DO437(wdataD[949]),
 .DO436(wdataD[948]), .DO435(wdataD[947]), .DO434(wdataD[946]), .DO433(wdataD[945]), .DO432(wdataD[944]), .DO431(wdataD[943]), .DO430(wdataD[942]), .DO429(wdataD[941]),
 .DO428(wdataD[940]), .DO427(wdataD[939]), .DO426(wdataD[938]), .DO425(wdataD[937]), .DO424(wdataD[936]), .DO423(wdataD[935]), .DO422(wdataD[934]), .DO421(wdataD[933]),
 .DO420(wdataD[932]), .DO419(wdataD[931]), .DO418(wdataD[930]), .DO417(wdataD[929]), .DO416(wdataD[928]), .DO415(wdataD[927]), .DO414(wdataD[926]), .DO413(wdataD[925]),
 .DO412(wdataD[924]), .DO411(wdataD[923]), .DO410(wdataD[922]), .DO409(wdataD[921]), .DO408(wdataD[920]), .DO407(wdataD[919]), .DO406(wdataD[918]), .DO405(wdataD[917]),
 .DO404(wdataD[916]), .DO403(wdataD[915]), .DO402(wdataD[914]), .DO401(wdataD[913]), .DO400(wdataD[912]), .DO399(wdataD[911]), .DO398(wdataD[910]), .DO397(wdataD[909]),
 .DO396(wdataD[908]), .DO395(wdataD[907]), .DO394(wdataD[906]), .DO393(wdataD[905]), .DO392(wdataD[904]), .DO391(wdataD[903]), .DO390(wdataD[902]), .DO389(wdataD[901]),
 .DO388(wdataD[900]), .DO387(wdataD[899]), .DO386(wdataD[898]), .DO385(wdataD[897]), .DO384(wdataD[896]), .DO383(wdataD[895]), .DO382(wdataD[894]), .DO381(wdataD[893]),
 .DO380(wdataD[892]), .DO379(wdataD[891]), .DO378(wdataD[890]), .DO377(wdataD[889]), .DO376(wdataD[888]), .DO375(wdataD[887]), .DO374(wdataD[886]), .DO373(wdataD[885]),
 .DO372(wdataD[884]), .DO371(wdataD[883]), .DO370(wdataD[882]), .DO369(wdataD[881]), .DO368(wdataD[880]), .DO367(wdataD[879]), .DO366(wdataD[878]), .DO365(wdataD[877]),
 .DO364(wdataD[876]), .DO363(wdataD[875]), .DO362(wdataD[874]), .DO361(wdataD[873]), .DO360(wdataD[872]), .DO359(wdataD[871]), .DO358(wdataD[870]), .DO357(wdataD[869]),
 .DO356(wdataD[868]), .DO355(wdataD[867]), .DO354(wdataD[866]), .DO353(wdataD[865]), .DO352(wdataD[864]), .DO351(wdataD[863]), .DO350(wdataD[862]), .DO349(wdataD[861]),
 .DO348(wdataD[860]), .DO347(wdataD[859]), .DO346(wdataD[858]), .DO345(wdataD[857]), .DO344(wdataD[856]), .DO343(wdataD[855]), .DO342(wdataD[854]), .DO341(wdataD[853]),
 .DO340(wdataD[852]), .DO339(wdataD[851]), .DO338(wdataD[850]), .DO337(wdataD[849]), .DO336(wdataD[848]), .DO335(wdataD[847]), .DO334(wdataD[846]), .DO333(wdataD[845]),
 .DO332(wdataD[844]), .DO331(wdataD[843]), .DO330(wdataD[842]), .DO329(wdataD[841]), .DO328(wdataD[840]), .DO327(wdataD[839]), .DO326(wdataD[838]), .DO325(wdataD[837]),
 .DO324(wdataD[836]), .DO323(wdataD[835]), .DO322(wdataD[834]), .DO321(wdataD[833]), .DO320(wdataD[832]), .DO319(wdataD[831]), .DO318(wdataD[830]), .DO317(wdataD[829]),
 .DO316(wdataD[828]), .DO315(wdataD[827]), .DO314(wdataD[826]), .DO313(wdataD[825]), .DO312(wdataD[824]), .DO311(wdataD[823]), .DO310(wdataD[822]), .DO309(wdataD[821]),
 .DO308(wdataD[820]), .DO307(wdataD[819]), .DO306(wdataD[818]), .DO305(wdataD[817]), .DO304(wdataD[816]), .DO303(wdataD[815]), .DO302(wdataD[814]), .DO301(wdataD[813]),
 .DO300(wdataD[812]), .DO299(wdataD[811]), .DO298(wdataD[810]), .DO297(wdataD[809]), .DO296(wdataD[808]), .DO295(wdataD[807]), .DO294(wdataD[806]), .DO293(wdataD[805]),
 .DO292(wdataD[804]), .DO291(wdataD[803]), .DO290(wdataD[802]), .DO289(wdataD[801]), .DO288(wdataD[800]), .DO287(wdataD[799]), .DO286(wdataD[798]), .DO285(wdataD[797]),
 .DO284(wdataD[796]), .DO283(wdataD[795]), .DO282(wdataD[794]), .DO281(wdataD[793]), .DO280(wdataD[792]), .DO279(wdataD[791]), .DO278(wdataD[790]), .DO277(wdataD[789]),
 .DO276(wdataD[788]), .DO275(wdataD[787]), .DO274(wdataD[786]), .DO273(wdataD[785]), .DO272(wdataD[784]), .DO271(wdataD[783]), .DO270(wdataD[782]), .DO269(wdataD[781]),
 .DO268(wdataD[780]), .DO267(wdataD[779]), .DO266(wdataD[778]), .DO265(wdataD[777]), .DO264(wdataD[776]), .DO263(wdataD[775]), .DO262(wdataD[774]), .DO261(wdataD[773]),
 .DO260(wdataD[772]), .DO259(wdataD[771]), .DO258(wdataD[770]), .DO257(wdataD[769]), .DO256(wdataD[768]), .DO255(wdataD[767]), .DO254(wdataD[766]), .DO253(wdataD[765]),
 .DO252(wdataD[764]), .DO251(wdataD[763]), .DO250(wdataD[762]), .DO249(wdataD[761]), .DO248(wdataD[760]), .DO247(wdataD[759]), .DO246(wdataD[758]), .DO245(wdataD[757]),
 .DO244(wdataD[756]), .DO243(wdataD[755]), .DO242(wdataD[754]), .DO241(wdataD[753]), .DO240(wdataD[752]), .DO239(wdataD[751]), .DO238(wdataD[750]), .DO237(wdataD[749]),
 .DO236(wdataD[748]), .DO235(wdataD[747]), .DO234(wdataD[746]), .DO233(wdataD[745]), .DO232(wdataD[744]), .DO231(wdataD[743]), .DO230(wdataD[742]), .DO229(wdataD[741]),
 .DO228(wdataD[740]), .DO227(wdataD[739]), .DO226(wdataD[738]), .DO225(wdataD[737]), .DO224(wdataD[736]), .DO223(wdataD[735]), .DO222(wdataD[734]), .DO221(wdataD[733]),
 .DO220(wdataD[732]), .DO219(wdataD[731]), .DO218(wdataD[730]), .DO217(wdataD[729]), .DO216(wdataD[728]), .DO215(wdataD[727]), .DO214(wdataD[726]), .DO213(wdataD[725]),
 .DO212(wdataD[724]), .DO211(wdataD[723]), .DO210(wdataD[722]), .DO209(wdataD[721]), .DO208(wdataD[720]), .DO207(wdataD[719]), .DO206(wdataD[718]), .DO205(wdataD[717]),
 .DO204(wdataD[716]), .DO203(wdataD[715]), .DO202(wdataD[714]), .DO201(wdataD[713]), .DO200(wdataD[712]), .DO199(wdataD[711]), .DO198(wdataD[710]), .DO197(wdataD[709]),
 .DO196(wdataD[708]), .DO195(wdataD[707]), .DO194(wdataD[706]), .DO193(wdataD[705]), .DO192(wdataD[704]), .DO191(wdataD[703]), .DO190(wdataD[702]), .DO189(wdataD[701]),
 .DO188(wdataD[700]), .DO187(wdataD[699]), .DO186(wdataD[698]), .DO185(wdataD[697]), .DO184(wdataD[696]), .DO183(wdataD[695]), .DO182(wdataD[694]), .DO181(wdataD[693]),
 .DO180(wdataD[692]), .DO179(wdataD[691]), .DO178(wdataD[690]), .DO177(wdataD[689]), .DO176(wdataD[688]), .DO175(wdataD[687]), .DO174(wdataD[686]), .DO173(wdataD[685]),
 .DO172(wdataD[684]), .DO171(wdataD[683]), .DO170(wdataD[682]), .DO169(wdataD[681]), .DO168(wdataD[680]), .DO167(wdataD[679]), .DO166(wdataD[678]), .DO165(wdataD[677]),
 .DO164(wdataD[676]), .DO163(wdataD[675]), .DO162(wdataD[674]), .DO161(wdataD[673]), .DO160(wdataD[672]), .DO159(wdataD[671]), .DO158(wdataD[670]), .DO157(wdataD[669]),
 .DO156(wdataD[668]), .DO155(wdataD[667]), .DO154(wdataD[666]), .DO153(wdataD[665]), .DO152(wdataD[664]), .DO151(wdataD[663]), .DO150(wdataD[662]), .DO149(wdataD[661]),
 .DO148(wdataD[660]), .DO147(wdataD[659]), .DO146(wdataD[658]), .DO145(wdataD[657]), .DO144(wdataD[656]), .DO143(wdataD[655]), .DO142(wdataD[654]), .DO141(wdataD[653]),
 .DO140(wdataD[652]), .DO139(wdataD[651]), .DO138(wdataD[650]), .DO137(wdataD[649]), .DO136(wdataD[648]), .DO135(wdataD[647]), .DO134(wdataD[646]), .DO133(wdataD[645]),
 .DO132(wdataD[644]), .DO131(wdataD[643]), .DO130(wdataD[642]), .DO129(wdataD[641]), .DO128(wdataD[640]), .DO127(wdataD[639]), .DO126(wdataD[638]), .DO125(wdataD[637]),
 .DO124(wdataD[636]), .DO123(wdataD[635]), .DO122(wdataD[634]), .DO121(wdataD[633]), .DO120(wdataD[632]), .DO119(wdataD[631]), .DO118(wdataD[630]), .DO117(wdataD[629]),
 .DO116(wdataD[628]), .DO115(wdataD[627]), .DO114(wdataD[626]), .DO113(wdataD[625]), .DO112(wdataD[624]), .DO111(wdataD[623]), .DO110(wdataD[622]), .DO109(wdataD[621]),
 .DO108(wdataD[620]), .DO107(wdataD[619]), .DO106(wdataD[618]), .DO105(wdataD[617]), .DO104(wdataD[616]), .DO103(wdataD[615]), .DO102(wdataD[614]), .DO101(wdataD[613]),
 .DO100(wdataD[612]), .DO99(wdataD[611]), .DO98(wdataD[610]), .DO97(wdataD[609]), .DO96(wdataD[608]), .DO95(wdataD[607]), .DO94(wdataD[606]), .DO93(wdataD[605]),
 .DO92(wdataD[604]), .DO91(wdataD[603]), .DO90(wdataD[602]), .DO89(wdataD[601]), .DO88(wdataD[600]), .DO87(wdataD[599]), .DO86(wdataD[598]), .DO85(wdataD[597]),
 .DO84(wdataD[596]), .DO83(wdataD[595]), .DO82(wdataD[594]), .DO81(wdataD[593]), .DO80(wdataD[592]), .DO79(wdataD[591]), .DO78(wdataD[590]), .DO77(wdataD[589]),
 .DO76(wdataD[588]), .DO75(wdataD[587]), .DO74(wdataD[586]), .DO73(wdataD[585]), .DO72(wdataD[584]), .DO71(wdataD[583]), .DO70(wdataD[582]), .DO69(wdataD[581]),
 .DO68(wdataD[580]), .DO67(wdataD[579]), .DO66(wdataD[578]), .DO65(wdataD[577]), .DO64(wdataD[576]), .DO63(wdataD[575]), .DO62(wdataD[574]), .DO61(wdataD[573]),
 .DO60(wdataD[572]), .DO59(wdataD[571]), .DO58(wdataD[570]), .DO57(wdataD[569]), .DO56(wdataD[568]), .DO55(wdataD[567]), .DO54(wdataD[566]), .DO53(wdataD[565]),
 .DO52(wdataD[564]), .DO51(wdataD[563]), .DO50(wdataD[562]), .DO49(wdataD[561]), .DO48(wdataD[560]), .DO47(wdataD[559]), .DO46(wdataD[558]), .DO45(wdataD[557]),
 .DO44(wdataD[556]), .DO43(wdataD[555]), .DO42(wdataD[554]), .DO41(wdataD[553]), .DO40(wdataD[552]), .DO39(wdataD[551]), .DO38(wdataD[550]), .DO37(wdataD[549]),
 .DO36(wdataD[548]), .DO35(wdataD[547]), .DO34(wdataD[546]), .DO33(wdataD[545]), .DO32(wdataD[544]), .DO31(wdataD[543]), .DO30(wdataD[542]), .DO29(wdataD[541]),
 .DO28(wdataD[540]), .DO27(wdataD[539]), .DO26(wdataD[538]), .DO25(wdataD[537]), .DO24(wdataD[536]), .DO23(wdataD[535]), .DO22(wdataD[534]), .DO21(wdataD[533]),
 .DO20(wdataD[532]), .DO19(wdataD[531]), .DO18(wdataD[530]), .DO17(wdataD[529]), .DO16(wdataD[528]), .DO15(wdataD[527]), .DO14(wdataD[526]), .DO13(wdataD[525]),
 .DO12(wdataD[524]), .DO11(wdataD[523]), .DO10(wdataD[522]), .DO9(wdataD[521]), .DO8(wdataD[520]), .DO7(wdataD[519]), .DO6(wdataD[518]), .DO5(wdataD[517]),
 .DO4(wdataD[516]), .DO3(wdataD[515]), .DO2(wdataD[514]), .DO1(wdataD[513]), .DO0(wdataD[512]), .SYNC_OUT(n9));
MPR4X512 U9 ( .A1(n5), .A0(n4), .SYNC_IN(n9), .DO511( ), .DO510( ), .DO509( ),
 .DO508( ), .DO507( ), .DO506( ), .DO505( ), .DO504( ), .DO503( ), .DO502( ), .DO501( ),
 .DO500( ), .DO499( ), .DO498( ), .DO497( ), .DO496( ), .DO495( ), .DO494( ), .DO493( ),
 .DO492( ), .DO491( ), .DO490( ), .DO489( ), .DO488( ), .DO487( ), .DO486( ), .DO485( ),
 .DO484( ), .DO483( ), .DO482( ), .DO481( ), .DO480( ), .DO479( ), .DO478( ), .DO477( ),
 .DO476( ), .DO475( ), .DO474( ), .DO473( ), .DO472( ), .DO471( ), .DO470( ), .DO469( ),
 .DO468( ), .DO467( ), .DO466( ), .DO465( ), .DO464( ), .DO463( ), .DO462( ), .DO461( ),
 .DO460( ), .DO459( ), .DO458( ), .DO457( ), .DO456( ), .DO455( ), .DO454( ), .DO453( ),
 .DO452( ), .DO451( ), .DO450( ), .DO449( ), .DO448( ), .DO447( ), .DO446( ), .DO445( ),
 .DO444( ), .DO443( ), .DO442( ), .DO441( ), .DO440( ), .DO439( ), .DO438( ), .DO437( ),
 .DO436( ), .DO435( ), .DO434( ), .DO433( ), .DO432( ), .DO431( ), .DO430( ), .DO429( ),
 .DO428( ), .DO427( ), .DO426( ), .DO425( ), .DO424( ), .DO423( ), .DO422( ), .DO421( ),
 .DO420( ), .DO419( ), .DO418( ), .DO417( ), .DO416( ), .DO415( ), .DO414( ), .DO413( ),
 .DO412( ), .DO411( ), .DO410( ), .DO409( ), .DO408( ), .DO407( ), .DO406( ), .DO405( ),
 .DO404( ), .DO403( ), .DO402( ), .DO401( ), .DO400( ), .DO399( ), .DO398( ), .DO397( ),
 .DO396( ), .DO395( ), .DO394( ), .DO393( ), .DO392( ), .DO391( ), .DO390( ), .DO389( ),
 .DO388( ), .DO387( ), .DO386( ), .DO385( ), .DO384( ), .DO383( ), .DO382( ), .DO381( ),
 .DO380( ), .DO379( ), .DO378( ), .DO377( ), .DO376( ), .DO375( ), .DO374( ), .DO373( ),
 .DO372( ), .DO371( ), .DO370( ), .DO369( ), .DO368( ), .DO367( ), .DO366( ), .DO365( ),
 .DO364( ), .DO363( ), .DO362( ), .DO361( ), .DO360( ), .DO359( ), .DO358( ), .DO357( ),
 .DO356( ), .DO355( ), .DO354( ), .DO353( ), .DO352( ), .DO351( ), .DO350( ), .DO349( ),
 .DO348( ), .DO347( ), .DO346( ), .DO345( ), .DO344( ), .DO343( ), .DO342( ), .DO341( ),
 .DO340( ), .DO339( ), .DO338( ), .DO337( ), .DO336( ), .DO335( ), .DO334( ), .DO333( ),
 .DO332( ), .DO331( ), .DO330( ), .DO329( ), .DO328( ), .DO327( ), .DO326( ), .DO325( ),
 .DO324( ), .DO323( ), .DO322( ), .DO321( ), .DO320( ), .DO319( ), .DO318( ), .DO317( ),
 .DO316( ), .DO315( ), .DO314( ), .DO313( ), .DO312( ), .DO311( ), .DO310( ), .DO309( ),
 .DO308( ), .DO307( ), .DO306( ), .DO305( ), .DO304( ), .DO303( ), .DO302( ), .DO301( ),
 .DO300( ), .DO299( ), .DO298( ), .DO297( ), .DO296( ), .DO295( ), .DO294( ), .DO293( ),
 .DO292( ), .DO291( ), .DO290( ), .DO289( ), .DO288( ), .DO287( ), .DO286( ), .DO285( ),
 .DO284( ), .DO283( ), .DO282( ), .DO281( ), .DO280( ), .DO279( ), .DO278( ), .DO277( ),
 .DO276( ), .DO275( ), .DO274( ), .DO273( ), .DO272( ), .DO271( ), .DO270( ), .DO269( ),
 .DO268( ), .DO267( ), .DO266( ), .DO265( ), .DO264( ), .DO263( ), .DO262( ), .DO261( ),
 .DO260( ), .DO259( ), .DO258( ), .DO257( ), .DO256( ), .DO255( ), .DO254( ), .DO253( ),
 .DO252( ), .DO251( ), .DO250( ), .DO249( ), .DO248( ), .DO247( ), .DO246( ), .DO245( ),
 .DO244( ), .DO243( ), .DO242( ), .DO241( ), .DO240( ), .DO239( ), .DO238( ), .DO237( ),
 .DO236( ), .DO235( ), .DO234( ), .DO233( ), .DO232( ), .DO231( ), .DO230( ), .DO229( ),
 .DO228( ), .DO227( ), .DO226( ), .DO225( ), .DO224( ), .DO223( ), .DO222( ), .DO221( ),
 .DO220( ), .DO219( ), .DO218( ), .DO217( ), .DO216( ), .DO215( ), .DO214( ), .DO213( ),
 .DO212( ), .DO211( ), .DO210( ), .DO209( ), .DO208( ), .DO207( ), .DO206( ), .DO205( ),
 .DO204( ), .DO203( ), .DO202( ), .DO201( ), .DO200( ), .DO199( ), .DO198( ), .DO197( ),
 .DO196( ), .DO195( ), .DO194( ), .DO193( ), .DO192( ), .DO191( ), .DO190( ), .DO189( ),
 .DO188( ), .DO187( ), .DO186( ), .DO185( ), .DO184( ), .DO183( ), .DO182( ), .DO181( ),
 .DO180( ), .DO179( ), .DO178( ), .DO177( ), .DO176( ), .DO175( ), .DO174( ), .DO173( ),
 .DO172( ), .DO171( ), .DO170( ), .DO169( ), .DO168( ), .DO167( ), .DO166( ), .DO165( ),
 .DO164( ), .DO163( ), .DO162( ), .DO161( ), .DO160( ), .DO159( ), .DO158( ), .DO157( ),
 .DO156( ), .DO155( ), .DO154( ), .DO153( ), .DO152( ), .DO151( ), .DO150( ), .DO149( ),
 .DO148( ), .DO147( ), .DO146( ), .DO145( ), .DO144( ), .DO143( ), .DO142( ), .DO141( ),
 .DO140( ), .DO139( ), .DO138( ), .DO137( ), .DO136( ), .DO135( ), .DO134( ), .DO133( ),
 .DO132( ), .DO131( ), .DO130( ), .DO129( ), .DO128( ), .DO127( ), .DO126( ), .DO125( ),
 .DO124( ), .DO123( ), .DO122( ), .DO121( ), .DO120( ), .DO119( ), .DO118( ), .DO117( ),
 .DO116( ), .DO115( ), .DO114( ), .DO113( ), .DO112( ), .DO111( ), .DO110( ), .DO109( ),
 .DO108( ), .DO107( ), .DO106( ), .DO105( ), .DO104( ), .DO103( ), .DO102( ), .DO101( ),
 .DO100( ), .DO99( ), .DO98( ), .DO97( ), .DO96( ), .DO95( ), .DO94( ), .DO93( ),
 .DO92( ), .DO91( ), .DO90( ), .DO89( ), .DO88( ), .DO87( ), .DO86( ), .DO85( ),
 .DO84( ), .DO83( ), .DO82( ), .DO81( ), .DO80( ), .DO79( ), .DO78( ), .DO77( ),
 .DO76( ), .DO75( ), .DO74( ), .DO73( ), .DO72( ), .DO71( ), .DO70( ), .DO69( ),
 .DO68( ), .DO67( ), .DO66( ), .DO65( ), .DO64( ), .DO63( ), .DO62( ), .DO61( ),
 .DO60( ), .DO59( ), .DO58( ), .DO57( ), .DO56( ), .DO55( ), .DO54( ), .DO53( ),
 .DO52( ), .DO51( ), .DO50( ), .DO49( ), .DO48( ), .DO47( ), .DO46( ), .DO45( ),
 .DO44( ), .DO43( ), .DO42( ), .DO41( ), .DO40( ), .DO39( ), .DO38( ), .DO37( ),
 .DO36( ), .DO35( ), .DO34( ), .DO33( ), .DO32( ), .DO31( ), .DO30( ), .DO29( ),
 .DO28( ), .DO27( ), .DO26( ), .DO25( ), .DO24( ), .DO23( ), .DO22( ), .DO21( ),
 .DO20( ), .DO19( ), .DO18( ), .DO17( ), .DO16( ), .DO15( ), .DO14( ), .DO13( ),
 .DO12( ), .DO11( ), .DO10( ), .DO9( ), .DO8( ), .DO7( ), .DO6( ), .DO5( ),
 .DO4( ), .DO3( ), .DO2( ), .DO1( ), .DO0(wdataD[1024]), .SYNC_OUT( ));
`endif
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "_zymem 1 511 0 0 2"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "1"
// pragma CVASTRPROP MODULE HDLICE CVAIUSNAMES_FORGEN_LABEL "genblk1"
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE "ixc_context_write"
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE_LIB "IXCOM_TEMP_LIBRARY"
// pragma CVASTRPROP MODULE HDLICE PROP_IXCOM_MOD TRUE
endmodule
`ifdef CBV
`else
`ifdef MPW4X512_MPR4X512
`else
module MPW4X512( A1, A0, DI511, DI510, DI509, DI508, DI507,
 DI506, DI505, DI504, DI503, DI502, DI501, DI500, DI499,
 DI498, DI497, DI496, DI495, DI494, DI493, DI492, DI491,
 DI490, DI489, DI488, DI487, DI486, DI485, DI484, DI483,
 DI482, DI481, DI480, DI479, DI478, DI477, DI476, DI475,
 DI474, DI473, DI472, DI471, DI470, DI469, DI468, DI467,
 DI466, DI465, DI464, DI463, DI462, DI461, DI460, DI459,
 DI458, DI457, DI456, DI455, DI454, DI453, DI452, DI451,
 DI450, DI449, DI448, DI447, DI446, DI445, DI444, DI443,
 DI442, DI441, DI440, DI439, DI438, DI437, DI436, DI435,
 DI434, DI433, DI432, DI431, DI430, DI429, DI428, DI427,
 DI426, DI425, DI424, DI423, DI422, DI421, DI420, DI419,
 DI418, DI417, DI416, DI415, DI414, DI413, DI412, DI411,
 DI410, DI409, DI408, DI407, DI406, DI405, DI404, DI403,
 DI402, DI401, DI400, DI399, DI398, DI397, DI396, DI395,
 DI394, DI393, DI392, DI391, DI390, DI389, DI388, DI387,
 DI386, DI385, DI384, DI383, DI382, DI381, DI380, DI379,
 DI378, DI377, DI376, DI375, DI374, DI373, DI372, DI371,
 DI370, DI369, DI368, DI367, DI366, DI365, DI364, DI363,
 DI362, DI361, DI360, DI359, DI358, DI357, DI356, DI355,
 DI354, DI353, DI352, DI351, DI350, DI349, DI348, DI347,
 DI346, DI345, DI344, DI343, DI342, DI341, DI340, DI339,
 DI338, DI337, DI336, DI335, DI334, DI333, DI332, DI331,
 DI330, DI329, DI328, DI327, DI326, DI325, DI324, DI323,
 DI322, DI321, DI320, DI319, DI318, DI317, DI316, DI315,
 DI314, DI313, DI312, DI311, DI310, DI309, DI308, DI307,
 DI306, DI305, DI304, DI303, DI302, DI301, DI300, DI299,
 DI298, DI297, DI296, DI295, DI294, DI293, DI292, DI291,
 DI290, DI289, DI288, DI287, DI286, DI285, DI284, DI283,
 DI282, DI281, DI280, DI279, DI278, DI277, DI276, DI275,
 DI274, DI273, DI272, DI271, DI270, DI269, DI268, DI267,
 DI266, DI265, DI264, DI263, DI262, DI261, DI260, DI259,
 DI258, DI257, DI256, DI255, DI254, DI253, DI252, DI251,
 DI250, DI249, DI248, DI247, DI246, DI245, DI244, DI243,
 DI242, DI241, DI240, DI239, DI238, DI237, DI236, DI235,
 DI234, DI233, DI232, DI231, DI230, DI229, DI228, DI227,
 DI226, DI225, DI224, DI223, DI222, DI221, DI220, DI219,
 DI218, DI217, DI216, DI215, DI214, DI213, DI212, DI211,
 DI210, DI209, DI208, DI207, DI206, DI205, DI204, DI203,
 DI202, DI201, DI200, DI199, DI198, DI197, DI196, DI195,
 DI194, DI193, DI192, DI191, DI190, DI189, DI188, DI187,
 DI186, DI185, DI184, DI183, DI182, DI181, DI180, DI179,
 DI178, DI177, DI176, DI175, DI174, DI173, DI172, DI171,
 DI170, DI169, DI168, DI167, DI166, DI165, DI164, DI163,
 DI162, DI161, DI160, DI159, DI158, DI157, DI156, DI155,
 DI154, DI153, DI152, DI151, DI150, DI149, DI148, DI147,
 DI146, DI145, DI144, DI143, DI142, DI141, DI140, DI139,
 DI138, DI137, DI136, DI135, DI134, DI133, DI132, DI131,
 DI130, DI129, DI128, DI127, DI126, DI125, DI124, DI123,
 DI122, DI121, DI120, DI119, DI118, DI117, DI116, DI115,
 DI114, DI113, DI112, DI111, DI110, DI109, DI108, DI107,
 DI106, DI105, DI104, DI103, DI102, DI101, DI100, DI99,
 DI98, DI97, DI96, DI95, DI94, DI93, DI92, DI91,
 DI90, DI89, DI88, DI87, DI86, DI85, DI84, DI83,
 DI82, DI81, DI80, DI79, DI78, DI77, DI76, DI75,
 DI74, DI73, DI72, DI71, DI70, DI69, DI68, DI67,
 DI66, DI65, DI64, DI63, DI62, DI61, DI60, DI59,
 DI58, DI57, DI56, DI55, DI54, DI53, DI52, DI51,
 DI50, DI49, DI48, DI47, DI46, DI45, DI44, DI43,
 DI42, DI41, DI40, DI39, DI38, DI37, DI36, DI35,
 DI34, DI33, DI32, DI31, DI30, DI29, DI28, DI27,
 DI26, DI25, DI24, DI23, DI22, DI21, DI20, DI19,
 DI18, DI17, DI16, DI15, DI14, DI13, DI12, DI11,
 DI10, DI9, DI8, DI7, DI6, DI5, DI4, DI3,
 DI2, DI1, DI0, WE, SYNC_IN, SYNC_OUT);
input  A1, A0, DI511, DI510, DI509, DI508, DI507, DI506,
 DI505, DI504, DI503, DI502, DI501, DI500, DI499, DI498, DI497, DI496,
 DI495, DI494, DI493, DI492, DI491, DI490, DI489, DI488, DI487, DI486,
 DI485, DI484, DI483, DI482, DI481, DI480, DI479, DI478, DI477, DI476,
 DI475, DI474, DI473, DI472, DI471, DI470, DI469, DI468, DI467, DI466,
 DI465, DI464, DI463, DI462, DI461, DI460, DI459, DI458, DI457, DI456,
 DI455, DI454, DI453, DI452, DI451, DI450, DI449, DI448, DI447, DI446,
 DI445, DI444, DI443, DI442, DI441, DI440, DI439, DI438, DI437, DI436,
 DI435, DI434, DI433, DI432, DI431, DI430, DI429, DI428, DI427, DI426,
 DI425, DI424, DI423, DI422, DI421, DI420, DI419, DI418, DI417, DI416,
 DI415, DI414, DI413, DI412, DI411, DI410, DI409, DI408, DI407, DI406,
 DI405, DI404, DI403, DI402, DI401, DI400, DI399, DI398, DI397, DI396,
 DI395, DI394, DI393, DI392, DI391, DI390, DI389, DI388, DI387, DI386,
 DI385, DI384, DI383, DI382, DI381, DI380, DI379, DI378, DI377, DI376,
 DI375, DI374, DI373, DI372, DI371, DI370, DI369, DI368, DI367, DI366,
 DI365, DI364, DI363, DI362, DI361, DI360, DI359, DI358, DI357, DI356,
 DI355, DI354, DI353, DI352, DI351, DI350, DI349, DI348, DI347, DI346,
 DI345, DI344, DI343, DI342, DI341, DI340, DI339, DI338, DI337, DI336,
 DI335, DI334, DI333, DI332, DI331, DI330, DI329, DI328, DI327, DI326,
 DI325, DI324, DI323, DI322, DI321, DI320, DI319, DI318, DI317, DI316,
 DI315, DI314, DI313, DI312, DI311, DI310, DI309, DI308, DI307, DI306,
 DI305, DI304, DI303, DI302, DI301, DI300, DI299, DI298, DI297, DI296,
 DI295, DI294, DI293, DI292, DI291, DI290, DI289, DI288, DI287, DI286,
 DI285, DI284, DI283, DI282, DI281, DI280, DI279, DI278, DI277, DI276,
 DI275, DI274, DI273, DI272, DI271, DI270, DI269, DI268, DI267, DI266,
 DI265, DI264, DI263, DI262, DI261, DI260, DI259, DI258, DI257, DI256,
 DI255, DI254, DI253, DI252, DI251, DI250, DI249, DI248, DI247, DI246,
 DI245, DI244, DI243, DI242, DI241, DI240, DI239, DI238, DI237, DI236,
 DI235, DI234, DI233, DI232, DI231, DI230, DI229, DI228, DI227, DI226,
 DI225, DI224, DI223, DI222, DI221, DI220, DI219, DI218, DI217, DI216,
 DI215, DI214, DI213, DI212, DI211, DI210, DI209, DI208, DI207, DI206,
 DI205, DI204, DI203, DI202, DI201, DI200, DI199, DI198, DI197, DI196,
 DI195, DI194, DI193, DI192, DI191, DI190, DI189, DI188, DI187, DI186,
 DI185, DI184, DI183, DI182, DI181, DI180, DI179, DI178, DI177, DI176,
 DI175, DI174, DI173, DI172, DI171, DI170, DI169, DI168, DI167, DI166,
 DI165, DI164, DI163, DI162, DI161, DI160, DI159, DI158, DI157, DI156,
 DI155, DI154, DI153, DI152, DI151, DI150, DI149, DI148, DI147, DI146,
 DI145, DI144, DI143, DI142, DI141, DI140, DI139, DI138, DI137, DI136,
 DI135, DI134, DI133, DI132, DI131, DI130, DI129, DI128, DI127, DI126,
 DI125, DI124, DI123, DI122, DI121, DI120, DI119, DI118, DI117, DI116,
 DI115, DI114, DI113, DI112, DI111, DI110, DI109, DI108, DI107, DI106,
 DI105, DI104, DI103, DI102, DI101, DI100, DI99, DI98, DI97, DI96,
 DI95, DI94, DI93, DI92, DI91, DI90, DI89, DI88, DI87, DI86,
 DI85, DI84, DI83, DI82, DI81, DI80, DI79, DI78, DI77, DI76,
 DI75, DI74, DI73, DI72, DI71, DI70, DI69, DI68, DI67, DI66,
 DI65, DI64, DI63, DI62, DI61, DI60, DI59, DI58, DI57, DI56,
 DI55, DI54, DI53, DI52, DI51, DI50, DI49, DI48, DI47, DI46,
 DI45, DI44, DI43, DI42, DI41, DI40, DI39, DI38, DI37, DI36,
 DI35, DI34, DI33, DI32, DI31, DI30, DI29, DI28, DI27, DI26,
 DI25, DI24, DI23, DI22, DI21, DI20, DI19, DI18, DI17, DI16,
 DI15, DI14, DI13, DI12, DI11, DI10, DI9, DI8, DI7, DI6,
 DI5, DI4, DI3, DI2, DI1, DI0, WE, SYNC_IN;
output  SYNC_OUT;
endmodule
`ifdef _MPR4X512_
`else
module MPR4X512( A1, A0, SYNC_IN, DO511, DO510, DO509, DO508,
 DO507, DO506, DO505, DO504, DO503, DO502, DO501, DO500,
 DO499, DO498, DO497, DO496, DO495, DO494, DO493, DO492,
 DO491, DO490, DO489, DO488, DO487, DO486, DO485, DO484,
 DO483, DO482, DO481, DO480, DO479, DO478, DO477, DO476,
 DO475, DO474, DO473, DO472, DO471, DO470, DO469, DO468,
 DO467, DO466, DO465, DO464, DO463, DO462, DO461, DO460,
 DO459, DO458, DO457, DO456, DO455, DO454, DO453, DO452,
 DO451, DO450, DO449, DO448, DO447, DO446, DO445, DO444,
 DO443, DO442, DO441, DO440, DO439, DO438, DO437, DO436,
 DO435, DO434, DO433, DO432, DO431, DO430, DO429, DO428,
 DO427, DO426, DO425, DO424, DO423, DO422, DO421, DO420,
 DO419, DO418, DO417, DO416, DO415, DO414, DO413, DO412,
 DO411, DO410, DO409, DO408, DO407, DO406, DO405, DO404,
 DO403, DO402, DO401, DO400, DO399, DO398, DO397, DO396,
 DO395, DO394, DO393, DO392, DO391, DO390, DO389, DO388,
 DO387, DO386, DO385, DO384, DO383, DO382, DO381, DO380,
 DO379, DO378, DO377, DO376, DO375, DO374, DO373, DO372,
 DO371, DO370, DO369, DO368, DO367, DO366, DO365, DO364,
 DO363, DO362, DO361, DO360, DO359, DO358, DO357, DO356,
 DO355, DO354, DO353, DO352, DO351, DO350, DO349, DO348,
 DO347, DO346, DO345, DO344, DO343, DO342, DO341, DO340,
 DO339, DO338, DO337, DO336, DO335, DO334, DO333, DO332,
 DO331, DO330, DO329, DO328, DO327, DO326, DO325, DO324,
 DO323, DO322, DO321, DO320, DO319, DO318, DO317, DO316,
 DO315, DO314, DO313, DO312, DO311, DO310, DO309, DO308,
 DO307, DO306, DO305, DO304, DO303, DO302, DO301, DO300,
 DO299, DO298, DO297, DO296, DO295, DO294, DO293, DO292,
 DO291, DO290, DO289, DO288, DO287, DO286, DO285, DO284,
 DO283, DO282, DO281, DO280, DO279, DO278, DO277, DO276,
 DO275, DO274, DO273, DO272, DO271, DO270, DO269, DO268,
 DO267, DO266, DO265, DO264, DO263, DO262, DO261, DO260,
 DO259, DO258, DO257, DO256, DO255, DO254, DO253, DO252,
 DO251, DO250, DO249, DO248, DO247, DO246, DO245, DO244,
 DO243, DO242, DO241, DO240, DO239, DO238, DO237, DO236,
 DO235, DO234, DO233, DO232, DO231, DO230, DO229, DO228,
 DO227, DO226, DO225, DO224, DO223, DO222, DO221, DO220,
 DO219, DO218, DO217, DO216, DO215, DO214, DO213, DO212,
 DO211, DO210, DO209, DO208, DO207, DO206, DO205, DO204,
 DO203, DO202, DO201, DO200, DO199, DO198, DO197, DO196,
 DO195, DO194, DO193, DO192, DO191, DO190, DO189, DO188,
 DO187, DO186, DO185, DO184, DO183, DO182, DO181, DO180,
 DO179, DO178, DO177, DO176, DO175, DO174, DO173, DO172,
 DO171, DO170, DO169, DO168, DO167, DO166, DO165, DO164,
 DO163, DO162, DO161, DO160, DO159, DO158, DO157, DO156,
 DO155, DO154, DO153, DO152, DO151, DO150, DO149, DO148,
 DO147, DO146, DO145, DO144, DO143, DO142, DO141, DO140,
 DO139, DO138, DO137, DO136, DO135, DO134, DO133, DO132,
 DO131, DO130, DO129, DO128, DO127, DO126, DO125, DO124,
 DO123, DO122, DO121, DO120, DO119, DO118, DO117, DO116,
 DO115, DO114, DO113, DO112, DO111, DO110, DO109, DO108,
 DO107, DO106, DO105, DO104, DO103, DO102, DO101, DO100,
 DO99, DO98, DO97, DO96, DO95, DO94, DO93, DO92,
 DO91, DO90, DO89, DO88, DO87, DO86, DO85, DO84,
 DO83, DO82, DO81, DO80, DO79, DO78, DO77, DO76,
 DO75, DO74, DO73, DO72, DO71, DO70, DO69, DO68,
 DO67, DO66, DO65, DO64, DO63, DO62, DO61, DO60,
 DO59, DO58, DO57, DO56, DO55, DO54, DO53, DO52,
 DO51, DO50, DO49, DO48, DO47, DO46, DO45, DO44,
 DO43, DO42, DO41, DO40, DO39, DO38, DO37, DO36,
 DO35, DO34, DO33, DO32, DO31, DO30, DO29, DO28,
 DO27, DO26, DO25, DO24, DO23, DO22, DO21, DO20,
 DO19, DO18, DO17, DO16, DO15, DO14, DO13, DO12,
 DO11, DO10, DO9, DO8, DO7, DO6, DO5, DO4,
 DO3, DO2, DO1, DO0, SYNC_OUT);
input  A1, A0, SYNC_IN;
output  DO511, DO510, DO509, DO508, DO507, DO506, DO505, DO504,
 DO503, DO502, DO501, DO500, DO499, DO498, DO497, DO496, DO495, DO494,
 DO493, DO492, DO491, DO490, DO489, DO488, DO487, DO486, DO485, DO484,
 DO483, DO482, DO481, DO480, DO479, DO478, DO477, DO476, DO475, DO474,
 DO473, DO472, DO471, DO470, DO469, DO468, DO467, DO466, DO465, DO464,
 DO463, DO462, DO461, DO460, DO459, DO458, DO457, DO456, DO455, DO454,
 DO453, DO452, DO451, DO450, DO449, DO448, DO447, DO446, DO445, DO444,
 DO443, DO442, DO441, DO440, DO439, DO438, DO437, DO436, DO435, DO434,
 DO433, DO432, DO431, DO430, DO429, DO428, DO427, DO426, DO425, DO424,
 DO423, DO422, DO421, DO420, DO419, DO418, DO417, DO416, DO415, DO414,
 DO413, DO412, DO411, DO410, DO409, DO408, DO407, DO406, DO405, DO404,
 DO403, DO402, DO401, DO400, DO399, DO398, DO397, DO396, DO395, DO394,
 DO393, DO392, DO391, DO390, DO389, DO388, DO387, DO386, DO385, DO384,
 DO383, DO382, DO381, DO380, DO379, DO378, DO377, DO376, DO375, DO374,
 DO373, DO372, DO371, DO370, DO369, DO368, DO367, DO366, DO365, DO364,
 DO363, DO362, DO361, DO360, DO359, DO358, DO357, DO356, DO355, DO354,
 DO353, DO352, DO351, DO350, DO349, DO348, DO347, DO346, DO345, DO344,
 DO343, DO342, DO341, DO340, DO339, DO338, DO337, DO336, DO335, DO334,
 DO333, DO332, DO331, DO330, DO329, DO328, DO327, DO326, DO325, DO324,
 DO323, DO322, DO321, DO320, DO319, DO318, DO317, DO316, DO315, DO314,
 DO313, DO312, DO311, DO310, DO309, DO308, DO307, DO306, DO305, DO304,
 DO303, DO302, DO301, DO300, DO299, DO298, DO297, DO296, DO295, DO294,
 DO293, DO292, DO291, DO290, DO289, DO288, DO287, DO286, DO285, DO284,
 DO283, DO282, DO281, DO280, DO279, DO278, DO277, DO276, DO275, DO274,
 DO273, DO272, DO271, DO270, DO269, DO268, DO267, DO266, DO265, DO264,
 DO263, DO262, DO261, DO260, DO259, DO258, DO257, DO256, DO255, DO254,
 DO253, DO252, DO251, DO250, DO249, DO248, DO247, DO246, DO245, DO244,
 DO243, DO242, DO241, DO240, DO239, DO238, DO237, DO236, DO235, DO234,
 DO233, DO232, DO231, DO230, DO229, DO228, DO227, DO226, DO225, DO224,
 DO223, DO222, DO221, DO220, DO219, DO218, DO217, DO216, DO215, DO214,
 DO213, DO212, DO211, DO210, DO209, DO208, DO207, DO206, DO205, DO204,
 DO203, DO202, DO201, DO200, DO199, DO198, DO197, DO196, DO195, DO194,
 DO193, DO192, DO191, DO190, DO189, DO188, DO187, DO186, DO185, DO184,
 DO183, DO182, DO181, DO180, DO179, DO178, DO177, DO176, DO175, DO174,
 DO173, DO172, DO171, DO170, DO169, DO168, DO167, DO166, DO165, DO164,
 DO163, DO162, DO161, DO160, DO159, DO158, DO157, DO156, DO155, DO154,
 DO153, DO152, DO151, DO150, DO149, DO148, DO147, DO146, DO145, DO144,
 DO143, DO142, DO141, DO140, DO139, DO138, DO137, DO136, DO135, DO134,
 DO133, DO132, DO131, DO130, DO129, DO128, DO127, DO126, DO125, DO124,
 DO123, DO122, DO121, DO120, DO119, DO118, DO117, DO116, DO115, DO114,
 DO113, DO112, DO111, DO110, DO109, DO108, DO107, DO106, DO105, DO104,
 DO103, DO102, DO101, DO100, DO99, DO98, DO97, DO96, DO95, DO94,
 DO93, DO92, DO91, DO90, DO89, DO88, DO87, DO86, DO85, DO84,
 DO83, DO82, DO81, DO80, DO79, DO78, DO77, DO76, DO75, DO74,
 DO73, DO72, DO71, DO70, DO69, DO68, DO67, DO66, DO65, DO64,
 DO63, DO62, DO61, DO60, DO59, DO58, DO57, DO56, DO55, DO54,
 DO53, DO52, DO51, DO50, DO49, DO48, DO47, DO46, DO45, DO44,
 DO43, DO42, DO41, DO40, DO39, DO38, DO37, DO36, DO35, DO34,
 DO33, DO32, DO31, DO30, DO29, DO28, DO27, DO26, DO25, DO24,
 DO23, DO22, DO21, DO20, DO19, DO18, DO17, DO16, DO15, DO14,
 DO13, DO12, DO11, DO10, DO9, DO8, DO7, DO6, DO5, DO4,
 DO3, DO2, DO1, DO0, SYNC_OUT;
endmodule
`define _MPR4X512_
`endif
`define MPW4X512_MPR4X512
`endif
`endif
