
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
(* upf_always_on = 1 *) 
module ixc_rforce_1024 ( L, V, en);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
input [1023:0] L;
input [1023:0] V;
input en;
wire fclk;
wire fen;
wire ren;
`_2_ wire _zzenr;
Q_NOT_TOUCH _zzqnthw ( .sig());
Q_RELEASE_WEAK \genblk1[1023].rrel ( .Q(L[1023]), .E(ren));
Q_REGFORCE \genblk1[1023].rfrc ( .Q(L[1023]), .A(V[1023]), .E(fen));
Q_RELEASE_WEAK \genblk1[1022].rrel ( .Q(L[1022]), .E(ren));
Q_REGFORCE \genblk1[1022].rfrc ( .Q(L[1022]), .A(V[1022]), .E(fen));
Q_RELEASE_WEAK \genblk1[1021].rrel ( .Q(L[1021]), .E(ren));
Q_REGFORCE \genblk1[1021].rfrc ( .Q(L[1021]), .A(V[1021]), .E(fen));
Q_RELEASE_WEAK \genblk1[1020].rrel ( .Q(L[1020]), .E(ren));
Q_REGFORCE \genblk1[1020].rfrc ( .Q(L[1020]), .A(V[1020]), .E(fen));
Q_RELEASE_WEAK \genblk1[1019].rrel ( .Q(L[1019]), .E(ren));
Q_REGFORCE \genblk1[1019].rfrc ( .Q(L[1019]), .A(V[1019]), .E(fen));
Q_RELEASE_WEAK \genblk1[1018].rrel ( .Q(L[1018]), .E(ren));
Q_REGFORCE \genblk1[1018].rfrc ( .Q(L[1018]), .A(V[1018]), .E(fen));
Q_RELEASE_WEAK \genblk1[1017].rrel ( .Q(L[1017]), .E(ren));
Q_REGFORCE \genblk1[1017].rfrc ( .Q(L[1017]), .A(V[1017]), .E(fen));
Q_RELEASE_WEAK \genblk1[1016].rrel ( .Q(L[1016]), .E(ren));
Q_REGFORCE \genblk1[1016].rfrc ( .Q(L[1016]), .A(V[1016]), .E(fen));
Q_RELEASE_WEAK \genblk1[1015].rrel ( .Q(L[1015]), .E(ren));
Q_REGFORCE \genblk1[1015].rfrc ( .Q(L[1015]), .A(V[1015]), .E(fen));
Q_RELEASE_WEAK \genblk1[1014].rrel ( .Q(L[1014]), .E(ren));
Q_REGFORCE \genblk1[1014].rfrc ( .Q(L[1014]), .A(V[1014]), .E(fen));
Q_RELEASE_WEAK \genblk1[1013].rrel ( .Q(L[1013]), .E(ren));
Q_REGFORCE \genblk1[1013].rfrc ( .Q(L[1013]), .A(V[1013]), .E(fen));
Q_RELEASE_WEAK \genblk1[1012].rrel ( .Q(L[1012]), .E(ren));
Q_REGFORCE \genblk1[1012].rfrc ( .Q(L[1012]), .A(V[1012]), .E(fen));
Q_RELEASE_WEAK \genblk1[1011].rrel ( .Q(L[1011]), .E(ren));
Q_REGFORCE \genblk1[1011].rfrc ( .Q(L[1011]), .A(V[1011]), .E(fen));
Q_RELEASE_WEAK \genblk1[1010].rrel ( .Q(L[1010]), .E(ren));
Q_REGFORCE \genblk1[1010].rfrc ( .Q(L[1010]), .A(V[1010]), .E(fen));
Q_RELEASE_WEAK \genblk1[1009].rrel ( .Q(L[1009]), .E(ren));
Q_REGFORCE \genblk1[1009].rfrc ( .Q(L[1009]), .A(V[1009]), .E(fen));
Q_RELEASE_WEAK \genblk1[1008].rrel ( .Q(L[1008]), .E(ren));
Q_REGFORCE \genblk1[1008].rfrc ( .Q(L[1008]), .A(V[1008]), .E(fen));
Q_RELEASE_WEAK \genblk1[1007].rrel ( .Q(L[1007]), .E(ren));
Q_REGFORCE \genblk1[1007].rfrc ( .Q(L[1007]), .A(V[1007]), .E(fen));
Q_RELEASE_WEAK \genblk1[1006].rrel ( .Q(L[1006]), .E(ren));
Q_REGFORCE \genblk1[1006].rfrc ( .Q(L[1006]), .A(V[1006]), .E(fen));
Q_RELEASE_WEAK \genblk1[1005].rrel ( .Q(L[1005]), .E(ren));
Q_REGFORCE \genblk1[1005].rfrc ( .Q(L[1005]), .A(V[1005]), .E(fen));
Q_RELEASE_WEAK \genblk1[1004].rrel ( .Q(L[1004]), .E(ren));
Q_REGFORCE \genblk1[1004].rfrc ( .Q(L[1004]), .A(V[1004]), .E(fen));
Q_RELEASE_WEAK \genblk1[1003].rrel ( .Q(L[1003]), .E(ren));
Q_REGFORCE \genblk1[1003].rfrc ( .Q(L[1003]), .A(V[1003]), .E(fen));
Q_RELEASE_WEAK \genblk1[1002].rrel ( .Q(L[1002]), .E(ren));
Q_REGFORCE \genblk1[1002].rfrc ( .Q(L[1002]), .A(V[1002]), .E(fen));
Q_RELEASE_WEAK \genblk1[1001].rrel ( .Q(L[1001]), .E(ren));
Q_REGFORCE \genblk1[1001].rfrc ( .Q(L[1001]), .A(V[1001]), .E(fen));
Q_RELEASE_WEAK \genblk1[1000].rrel ( .Q(L[1000]), .E(ren));
Q_REGFORCE \genblk1[1000].rfrc ( .Q(L[1000]), .A(V[1000]), .E(fen));
Q_RELEASE_WEAK \genblk1[999].rrel ( .Q(L[999]), .E(ren));
Q_REGFORCE \genblk1[999].rfrc ( .Q(L[999]), .A(V[999]), .E(fen));
Q_RELEASE_WEAK \genblk1[998].rrel ( .Q(L[998]), .E(ren));
Q_REGFORCE \genblk1[998].rfrc ( .Q(L[998]), .A(V[998]), .E(fen));
Q_RELEASE_WEAK \genblk1[997].rrel ( .Q(L[997]), .E(ren));
Q_REGFORCE \genblk1[997].rfrc ( .Q(L[997]), .A(V[997]), .E(fen));
Q_RELEASE_WEAK \genblk1[996].rrel ( .Q(L[996]), .E(ren));
Q_REGFORCE \genblk1[996].rfrc ( .Q(L[996]), .A(V[996]), .E(fen));
Q_RELEASE_WEAK \genblk1[995].rrel ( .Q(L[995]), .E(ren));
Q_REGFORCE \genblk1[995].rfrc ( .Q(L[995]), .A(V[995]), .E(fen));
Q_RELEASE_WEAK \genblk1[994].rrel ( .Q(L[994]), .E(ren));
Q_REGFORCE \genblk1[994].rfrc ( .Q(L[994]), .A(V[994]), .E(fen));
Q_RELEASE_WEAK \genblk1[993].rrel ( .Q(L[993]), .E(ren));
Q_REGFORCE \genblk1[993].rfrc ( .Q(L[993]), .A(V[993]), .E(fen));
Q_RELEASE_WEAK \genblk1[992].rrel ( .Q(L[992]), .E(ren));
Q_REGFORCE \genblk1[992].rfrc ( .Q(L[992]), .A(V[992]), .E(fen));
Q_RELEASE_WEAK \genblk1[991].rrel ( .Q(L[991]), .E(ren));
Q_REGFORCE \genblk1[991].rfrc ( .Q(L[991]), .A(V[991]), .E(fen));
Q_RELEASE_WEAK \genblk1[990].rrel ( .Q(L[990]), .E(ren));
Q_REGFORCE \genblk1[990].rfrc ( .Q(L[990]), .A(V[990]), .E(fen));
Q_RELEASE_WEAK \genblk1[989].rrel ( .Q(L[989]), .E(ren));
Q_REGFORCE \genblk1[989].rfrc ( .Q(L[989]), .A(V[989]), .E(fen));
Q_RELEASE_WEAK \genblk1[988].rrel ( .Q(L[988]), .E(ren));
Q_REGFORCE \genblk1[988].rfrc ( .Q(L[988]), .A(V[988]), .E(fen));
Q_RELEASE_WEAK \genblk1[987].rrel ( .Q(L[987]), .E(ren));
Q_REGFORCE \genblk1[987].rfrc ( .Q(L[987]), .A(V[987]), .E(fen));
Q_RELEASE_WEAK \genblk1[986].rrel ( .Q(L[986]), .E(ren));
Q_REGFORCE \genblk1[986].rfrc ( .Q(L[986]), .A(V[986]), .E(fen));
Q_RELEASE_WEAK \genblk1[985].rrel ( .Q(L[985]), .E(ren));
Q_REGFORCE \genblk1[985].rfrc ( .Q(L[985]), .A(V[985]), .E(fen));
Q_RELEASE_WEAK \genblk1[984].rrel ( .Q(L[984]), .E(ren));
Q_REGFORCE \genblk1[984].rfrc ( .Q(L[984]), .A(V[984]), .E(fen));
Q_RELEASE_WEAK \genblk1[983].rrel ( .Q(L[983]), .E(ren));
Q_REGFORCE \genblk1[983].rfrc ( .Q(L[983]), .A(V[983]), .E(fen));
Q_RELEASE_WEAK \genblk1[982].rrel ( .Q(L[982]), .E(ren));
Q_REGFORCE \genblk1[982].rfrc ( .Q(L[982]), .A(V[982]), .E(fen));
Q_RELEASE_WEAK \genblk1[981].rrel ( .Q(L[981]), .E(ren));
Q_REGFORCE \genblk1[981].rfrc ( .Q(L[981]), .A(V[981]), .E(fen));
Q_RELEASE_WEAK \genblk1[980].rrel ( .Q(L[980]), .E(ren));
Q_REGFORCE \genblk1[980].rfrc ( .Q(L[980]), .A(V[980]), .E(fen));
Q_RELEASE_WEAK \genblk1[979].rrel ( .Q(L[979]), .E(ren));
Q_REGFORCE \genblk1[979].rfrc ( .Q(L[979]), .A(V[979]), .E(fen));
Q_RELEASE_WEAK \genblk1[978].rrel ( .Q(L[978]), .E(ren));
Q_REGFORCE \genblk1[978].rfrc ( .Q(L[978]), .A(V[978]), .E(fen));
Q_RELEASE_WEAK \genblk1[977].rrel ( .Q(L[977]), .E(ren));
Q_REGFORCE \genblk1[977].rfrc ( .Q(L[977]), .A(V[977]), .E(fen));
Q_RELEASE_WEAK \genblk1[976].rrel ( .Q(L[976]), .E(ren));
Q_REGFORCE \genblk1[976].rfrc ( .Q(L[976]), .A(V[976]), .E(fen));
Q_RELEASE_WEAK \genblk1[975].rrel ( .Q(L[975]), .E(ren));
Q_REGFORCE \genblk1[975].rfrc ( .Q(L[975]), .A(V[975]), .E(fen));
Q_RELEASE_WEAK \genblk1[974].rrel ( .Q(L[974]), .E(ren));
Q_REGFORCE \genblk1[974].rfrc ( .Q(L[974]), .A(V[974]), .E(fen));
Q_RELEASE_WEAK \genblk1[973].rrel ( .Q(L[973]), .E(ren));
Q_REGFORCE \genblk1[973].rfrc ( .Q(L[973]), .A(V[973]), .E(fen));
Q_RELEASE_WEAK \genblk1[972].rrel ( .Q(L[972]), .E(ren));
Q_REGFORCE \genblk1[972].rfrc ( .Q(L[972]), .A(V[972]), .E(fen));
Q_RELEASE_WEAK \genblk1[971].rrel ( .Q(L[971]), .E(ren));
Q_REGFORCE \genblk1[971].rfrc ( .Q(L[971]), .A(V[971]), .E(fen));
Q_RELEASE_WEAK \genblk1[970].rrel ( .Q(L[970]), .E(ren));
Q_REGFORCE \genblk1[970].rfrc ( .Q(L[970]), .A(V[970]), .E(fen));
Q_RELEASE_WEAK \genblk1[969].rrel ( .Q(L[969]), .E(ren));
Q_REGFORCE \genblk1[969].rfrc ( .Q(L[969]), .A(V[969]), .E(fen));
Q_RELEASE_WEAK \genblk1[968].rrel ( .Q(L[968]), .E(ren));
Q_REGFORCE \genblk1[968].rfrc ( .Q(L[968]), .A(V[968]), .E(fen));
Q_RELEASE_WEAK \genblk1[967].rrel ( .Q(L[967]), .E(ren));
Q_REGFORCE \genblk1[967].rfrc ( .Q(L[967]), .A(V[967]), .E(fen));
Q_RELEASE_WEAK \genblk1[966].rrel ( .Q(L[966]), .E(ren));
Q_REGFORCE \genblk1[966].rfrc ( .Q(L[966]), .A(V[966]), .E(fen));
Q_RELEASE_WEAK \genblk1[965].rrel ( .Q(L[965]), .E(ren));
Q_REGFORCE \genblk1[965].rfrc ( .Q(L[965]), .A(V[965]), .E(fen));
Q_RELEASE_WEAK \genblk1[964].rrel ( .Q(L[964]), .E(ren));
Q_REGFORCE \genblk1[964].rfrc ( .Q(L[964]), .A(V[964]), .E(fen));
Q_RELEASE_WEAK \genblk1[963].rrel ( .Q(L[963]), .E(ren));
Q_REGFORCE \genblk1[963].rfrc ( .Q(L[963]), .A(V[963]), .E(fen));
Q_RELEASE_WEAK \genblk1[962].rrel ( .Q(L[962]), .E(ren));
Q_REGFORCE \genblk1[962].rfrc ( .Q(L[962]), .A(V[962]), .E(fen));
Q_RELEASE_WEAK \genblk1[961].rrel ( .Q(L[961]), .E(ren));
Q_REGFORCE \genblk1[961].rfrc ( .Q(L[961]), .A(V[961]), .E(fen));
Q_RELEASE_WEAK \genblk1[960].rrel ( .Q(L[960]), .E(ren));
Q_REGFORCE \genblk1[960].rfrc ( .Q(L[960]), .A(V[960]), .E(fen));
Q_RELEASE_WEAK \genblk1[959].rrel ( .Q(L[959]), .E(ren));
Q_REGFORCE \genblk1[959].rfrc ( .Q(L[959]), .A(V[959]), .E(fen));
Q_RELEASE_WEAK \genblk1[958].rrel ( .Q(L[958]), .E(ren));
Q_REGFORCE \genblk1[958].rfrc ( .Q(L[958]), .A(V[958]), .E(fen));
Q_RELEASE_WEAK \genblk1[957].rrel ( .Q(L[957]), .E(ren));
Q_REGFORCE \genblk1[957].rfrc ( .Q(L[957]), .A(V[957]), .E(fen));
Q_RELEASE_WEAK \genblk1[956].rrel ( .Q(L[956]), .E(ren));
Q_REGFORCE \genblk1[956].rfrc ( .Q(L[956]), .A(V[956]), .E(fen));
Q_RELEASE_WEAK \genblk1[955].rrel ( .Q(L[955]), .E(ren));
Q_REGFORCE \genblk1[955].rfrc ( .Q(L[955]), .A(V[955]), .E(fen));
Q_RELEASE_WEAK \genblk1[954].rrel ( .Q(L[954]), .E(ren));
Q_REGFORCE \genblk1[954].rfrc ( .Q(L[954]), .A(V[954]), .E(fen));
Q_RELEASE_WEAK \genblk1[953].rrel ( .Q(L[953]), .E(ren));
Q_REGFORCE \genblk1[953].rfrc ( .Q(L[953]), .A(V[953]), .E(fen));
Q_RELEASE_WEAK \genblk1[952].rrel ( .Q(L[952]), .E(ren));
Q_REGFORCE \genblk1[952].rfrc ( .Q(L[952]), .A(V[952]), .E(fen));
Q_RELEASE_WEAK \genblk1[951].rrel ( .Q(L[951]), .E(ren));
Q_REGFORCE \genblk1[951].rfrc ( .Q(L[951]), .A(V[951]), .E(fen));
Q_RELEASE_WEAK \genblk1[950].rrel ( .Q(L[950]), .E(ren));
Q_REGFORCE \genblk1[950].rfrc ( .Q(L[950]), .A(V[950]), .E(fen));
Q_RELEASE_WEAK \genblk1[949].rrel ( .Q(L[949]), .E(ren));
Q_REGFORCE \genblk1[949].rfrc ( .Q(L[949]), .A(V[949]), .E(fen));
Q_RELEASE_WEAK \genblk1[948].rrel ( .Q(L[948]), .E(ren));
Q_REGFORCE \genblk1[948].rfrc ( .Q(L[948]), .A(V[948]), .E(fen));
Q_RELEASE_WEAK \genblk1[947].rrel ( .Q(L[947]), .E(ren));
Q_REGFORCE \genblk1[947].rfrc ( .Q(L[947]), .A(V[947]), .E(fen));
Q_RELEASE_WEAK \genblk1[946].rrel ( .Q(L[946]), .E(ren));
Q_REGFORCE \genblk1[946].rfrc ( .Q(L[946]), .A(V[946]), .E(fen));
Q_RELEASE_WEAK \genblk1[945].rrel ( .Q(L[945]), .E(ren));
Q_REGFORCE \genblk1[945].rfrc ( .Q(L[945]), .A(V[945]), .E(fen));
Q_RELEASE_WEAK \genblk1[944].rrel ( .Q(L[944]), .E(ren));
Q_REGFORCE \genblk1[944].rfrc ( .Q(L[944]), .A(V[944]), .E(fen));
Q_RELEASE_WEAK \genblk1[943].rrel ( .Q(L[943]), .E(ren));
Q_REGFORCE \genblk1[943].rfrc ( .Q(L[943]), .A(V[943]), .E(fen));
Q_RELEASE_WEAK \genblk1[942].rrel ( .Q(L[942]), .E(ren));
Q_REGFORCE \genblk1[942].rfrc ( .Q(L[942]), .A(V[942]), .E(fen));
Q_RELEASE_WEAK \genblk1[941].rrel ( .Q(L[941]), .E(ren));
Q_REGFORCE \genblk1[941].rfrc ( .Q(L[941]), .A(V[941]), .E(fen));
Q_RELEASE_WEAK \genblk1[940].rrel ( .Q(L[940]), .E(ren));
Q_REGFORCE \genblk1[940].rfrc ( .Q(L[940]), .A(V[940]), .E(fen));
Q_RELEASE_WEAK \genblk1[939].rrel ( .Q(L[939]), .E(ren));
Q_REGFORCE \genblk1[939].rfrc ( .Q(L[939]), .A(V[939]), .E(fen));
Q_RELEASE_WEAK \genblk1[938].rrel ( .Q(L[938]), .E(ren));
Q_REGFORCE \genblk1[938].rfrc ( .Q(L[938]), .A(V[938]), .E(fen));
Q_RELEASE_WEAK \genblk1[937].rrel ( .Q(L[937]), .E(ren));
Q_REGFORCE \genblk1[937].rfrc ( .Q(L[937]), .A(V[937]), .E(fen));
Q_RELEASE_WEAK \genblk1[936].rrel ( .Q(L[936]), .E(ren));
Q_REGFORCE \genblk1[936].rfrc ( .Q(L[936]), .A(V[936]), .E(fen));
Q_RELEASE_WEAK \genblk1[935].rrel ( .Q(L[935]), .E(ren));
Q_REGFORCE \genblk1[935].rfrc ( .Q(L[935]), .A(V[935]), .E(fen));
Q_RELEASE_WEAK \genblk1[934].rrel ( .Q(L[934]), .E(ren));
Q_REGFORCE \genblk1[934].rfrc ( .Q(L[934]), .A(V[934]), .E(fen));
Q_RELEASE_WEAK \genblk1[933].rrel ( .Q(L[933]), .E(ren));
Q_REGFORCE \genblk1[933].rfrc ( .Q(L[933]), .A(V[933]), .E(fen));
Q_RELEASE_WEAK \genblk1[932].rrel ( .Q(L[932]), .E(ren));
Q_REGFORCE \genblk1[932].rfrc ( .Q(L[932]), .A(V[932]), .E(fen));
Q_RELEASE_WEAK \genblk1[931].rrel ( .Q(L[931]), .E(ren));
Q_REGFORCE \genblk1[931].rfrc ( .Q(L[931]), .A(V[931]), .E(fen));
Q_RELEASE_WEAK \genblk1[930].rrel ( .Q(L[930]), .E(ren));
Q_REGFORCE \genblk1[930].rfrc ( .Q(L[930]), .A(V[930]), .E(fen));
Q_RELEASE_WEAK \genblk1[929].rrel ( .Q(L[929]), .E(ren));
Q_REGFORCE \genblk1[929].rfrc ( .Q(L[929]), .A(V[929]), .E(fen));
Q_RELEASE_WEAK \genblk1[928].rrel ( .Q(L[928]), .E(ren));
Q_REGFORCE \genblk1[928].rfrc ( .Q(L[928]), .A(V[928]), .E(fen));
Q_RELEASE_WEAK \genblk1[927].rrel ( .Q(L[927]), .E(ren));
Q_REGFORCE \genblk1[927].rfrc ( .Q(L[927]), .A(V[927]), .E(fen));
Q_RELEASE_WEAK \genblk1[926].rrel ( .Q(L[926]), .E(ren));
Q_REGFORCE \genblk1[926].rfrc ( .Q(L[926]), .A(V[926]), .E(fen));
Q_RELEASE_WEAK \genblk1[925].rrel ( .Q(L[925]), .E(ren));
Q_REGFORCE \genblk1[925].rfrc ( .Q(L[925]), .A(V[925]), .E(fen));
Q_RELEASE_WEAK \genblk1[924].rrel ( .Q(L[924]), .E(ren));
Q_REGFORCE \genblk1[924].rfrc ( .Q(L[924]), .A(V[924]), .E(fen));
Q_RELEASE_WEAK \genblk1[923].rrel ( .Q(L[923]), .E(ren));
Q_REGFORCE \genblk1[923].rfrc ( .Q(L[923]), .A(V[923]), .E(fen));
Q_RELEASE_WEAK \genblk1[922].rrel ( .Q(L[922]), .E(ren));
Q_REGFORCE \genblk1[922].rfrc ( .Q(L[922]), .A(V[922]), .E(fen));
Q_RELEASE_WEAK \genblk1[921].rrel ( .Q(L[921]), .E(ren));
Q_REGFORCE \genblk1[921].rfrc ( .Q(L[921]), .A(V[921]), .E(fen));
Q_RELEASE_WEAK \genblk1[920].rrel ( .Q(L[920]), .E(ren));
Q_REGFORCE \genblk1[920].rfrc ( .Q(L[920]), .A(V[920]), .E(fen));
Q_RELEASE_WEAK \genblk1[919].rrel ( .Q(L[919]), .E(ren));
Q_REGFORCE \genblk1[919].rfrc ( .Q(L[919]), .A(V[919]), .E(fen));
Q_RELEASE_WEAK \genblk1[918].rrel ( .Q(L[918]), .E(ren));
Q_REGFORCE \genblk1[918].rfrc ( .Q(L[918]), .A(V[918]), .E(fen));
Q_RELEASE_WEAK \genblk1[917].rrel ( .Q(L[917]), .E(ren));
Q_REGFORCE \genblk1[917].rfrc ( .Q(L[917]), .A(V[917]), .E(fen));
Q_RELEASE_WEAK \genblk1[916].rrel ( .Q(L[916]), .E(ren));
Q_REGFORCE \genblk1[916].rfrc ( .Q(L[916]), .A(V[916]), .E(fen));
Q_RELEASE_WEAK \genblk1[915].rrel ( .Q(L[915]), .E(ren));
Q_REGFORCE \genblk1[915].rfrc ( .Q(L[915]), .A(V[915]), .E(fen));
Q_RELEASE_WEAK \genblk1[914].rrel ( .Q(L[914]), .E(ren));
Q_REGFORCE \genblk1[914].rfrc ( .Q(L[914]), .A(V[914]), .E(fen));
Q_RELEASE_WEAK \genblk1[913].rrel ( .Q(L[913]), .E(ren));
Q_REGFORCE \genblk1[913].rfrc ( .Q(L[913]), .A(V[913]), .E(fen));
Q_RELEASE_WEAK \genblk1[912].rrel ( .Q(L[912]), .E(ren));
Q_REGFORCE \genblk1[912].rfrc ( .Q(L[912]), .A(V[912]), .E(fen));
Q_RELEASE_WEAK \genblk1[911].rrel ( .Q(L[911]), .E(ren));
Q_REGFORCE \genblk1[911].rfrc ( .Q(L[911]), .A(V[911]), .E(fen));
Q_RELEASE_WEAK \genblk1[910].rrel ( .Q(L[910]), .E(ren));
Q_REGFORCE \genblk1[910].rfrc ( .Q(L[910]), .A(V[910]), .E(fen));
Q_RELEASE_WEAK \genblk1[909].rrel ( .Q(L[909]), .E(ren));
Q_REGFORCE \genblk1[909].rfrc ( .Q(L[909]), .A(V[909]), .E(fen));
Q_RELEASE_WEAK \genblk1[908].rrel ( .Q(L[908]), .E(ren));
Q_REGFORCE \genblk1[908].rfrc ( .Q(L[908]), .A(V[908]), .E(fen));
Q_RELEASE_WEAK \genblk1[907].rrel ( .Q(L[907]), .E(ren));
Q_REGFORCE \genblk1[907].rfrc ( .Q(L[907]), .A(V[907]), .E(fen));
Q_RELEASE_WEAK \genblk1[906].rrel ( .Q(L[906]), .E(ren));
Q_REGFORCE \genblk1[906].rfrc ( .Q(L[906]), .A(V[906]), .E(fen));
Q_RELEASE_WEAK \genblk1[905].rrel ( .Q(L[905]), .E(ren));
Q_REGFORCE \genblk1[905].rfrc ( .Q(L[905]), .A(V[905]), .E(fen));
Q_RELEASE_WEAK \genblk1[904].rrel ( .Q(L[904]), .E(ren));
Q_REGFORCE \genblk1[904].rfrc ( .Q(L[904]), .A(V[904]), .E(fen));
Q_RELEASE_WEAK \genblk1[903].rrel ( .Q(L[903]), .E(ren));
Q_REGFORCE \genblk1[903].rfrc ( .Q(L[903]), .A(V[903]), .E(fen));
Q_RELEASE_WEAK \genblk1[902].rrel ( .Q(L[902]), .E(ren));
Q_REGFORCE \genblk1[902].rfrc ( .Q(L[902]), .A(V[902]), .E(fen));
Q_RELEASE_WEAK \genblk1[901].rrel ( .Q(L[901]), .E(ren));
Q_REGFORCE \genblk1[901].rfrc ( .Q(L[901]), .A(V[901]), .E(fen));
Q_RELEASE_WEAK \genblk1[900].rrel ( .Q(L[900]), .E(ren));
Q_REGFORCE \genblk1[900].rfrc ( .Q(L[900]), .A(V[900]), .E(fen));
Q_RELEASE_WEAK \genblk1[899].rrel ( .Q(L[899]), .E(ren));
Q_REGFORCE \genblk1[899].rfrc ( .Q(L[899]), .A(V[899]), .E(fen));
Q_RELEASE_WEAK \genblk1[898].rrel ( .Q(L[898]), .E(ren));
Q_REGFORCE \genblk1[898].rfrc ( .Q(L[898]), .A(V[898]), .E(fen));
Q_RELEASE_WEAK \genblk1[897].rrel ( .Q(L[897]), .E(ren));
Q_REGFORCE \genblk1[897].rfrc ( .Q(L[897]), .A(V[897]), .E(fen));
Q_RELEASE_WEAK \genblk1[896].rrel ( .Q(L[896]), .E(ren));
Q_REGFORCE \genblk1[896].rfrc ( .Q(L[896]), .A(V[896]), .E(fen));
Q_RELEASE_WEAK \genblk1[895].rrel ( .Q(L[895]), .E(ren));
Q_REGFORCE \genblk1[895].rfrc ( .Q(L[895]), .A(V[895]), .E(fen));
Q_RELEASE_WEAK \genblk1[894].rrel ( .Q(L[894]), .E(ren));
Q_REGFORCE \genblk1[894].rfrc ( .Q(L[894]), .A(V[894]), .E(fen));
Q_RELEASE_WEAK \genblk1[893].rrel ( .Q(L[893]), .E(ren));
Q_REGFORCE \genblk1[893].rfrc ( .Q(L[893]), .A(V[893]), .E(fen));
Q_RELEASE_WEAK \genblk1[892].rrel ( .Q(L[892]), .E(ren));
Q_REGFORCE \genblk1[892].rfrc ( .Q(L[892]), .A(V[892]), .E(fen));
Q_RELEASE_WEAK \genblk1[891].rrel ( .Q(L[891]), .E(ren));
Q_REGFORCE \genblk1[891].rfrc ( .Q(L[891]), .A(V[891]), .E(fen));
Q_RELEASE_WEAK \genblk1[890].rrel ( .Q(L[890]), .E(ren));
Q_REGFORCE \genblk1[890].rfrc ( .Q(L[890]), .A(V[890]), .E(fen));
Q_RELEASE_WEAK \genblk1[889].rrel ( .Q(L[889]), .E(ren));
Q_REGFORCE \genblk1[889].rfrc ( .Q(L[889]), .A(V[889]), .E(fen));
Q_RELEASE_WEAK \genblk1[888].rrel ( .Q(L[888]), .E(ren));
Q_REGFORCE \genblk1[888].rfrc ( .Q(L[888]), .A(V[888]), .E(fen));
Q_RELEASE_WEAK \genblk1[887].rrel ( .Q(L[887]), .E(ren));
Q_REGFORCE \genblk1[887].rfrc ( .Q(L[887]), .A(V[887]), .E(fen));
Q_RELEASE_WEAK \genblk1[886].rrel ( .Q(L[886]), .E(ren));
Q_REGFORCE \genblk1[886].rfrc ( .Q(L[886]), .A(V[886]), .E(fen));
Q_RELEASE_WEAK \genblk1[885].rrel ( .Q(L[885]), .E(ren));
Q_REGFORCE \genblk1[885].rfrc ( .Q(L[885]), .A(V[885]), .E(fen));
Q_RELEASE_WEAK \genblk1[884].rrel ( .Q(L[884]), .E(ren));
Q_REGFORCE \genblk1[884].rfrc ( .Q(L[884]), .A(V[884]), .E(fen));
Q_RELEASE_WEAK \genblk1[883].rrel ( .Q(L[883]), .E(ren));
Q_REGFORCE \genblk1[883].rfrc ( .Q(L[883]), .A(V[883]), .E(fen));
Q_RELEASE_WEAK \genblk1[882].rrel ( .Q(L[882]), .E(ren));
Q_REGFORCE \genblk1[882].rfrc ( .Q(L[882]), .A(V[882]), .E(fen));
Q_RELEASE_WEAK \genblk1[881].rrel ( .Q(L[881]), .E(ren));
Q_REGFORCE \genblk1[881].rfrc ( .Q(L[881]), .A(V[881]), .E(fen));
Q_RELEASE_WEAK \genblk1[880].rrel ( .Q(L[880]), .E(ren));
Q_REGFORCE \genblk1[880].rfrc ( .Q(L[880]), .A(V[880]), .E(fen));
Q_RELEASE_WEAK \genblk1[879].rrel ( .Q(L[879]), .E(ren));
Q_REGFORCE \genblk1[879].rfrc ( .Q(L[879]), .A(V[879]), .E(fen));
Q_RELEASE_WEAK \genblk1[878].rrel ( .Q(L[878]), .E(ren));
Q_REGFORCE \genblk1[878].rfrc ( .Q(L[878]), .A(V[878]), .E(fen));
Q_RELEASE_WEAK \genblk1[877].rrel ( .Q(L[877]), .E(ren));
Q_REGFORCE \genblk1[877].rfrc ( .Q(L[877]), .A(V[877]), .E(fen));
Q_RELEASE_WEAK \genblk1[876].rrel ( .Q(L[876]), .E(ren));
Q_REGFORCE \genblk1[876].rfrc ( .Q(L[876]), .A(V[876]), .E(fen));
Q_RELEASE_WEAK \genblk1[875].rrel ( .Q(L[875]), .E(ren));
Q_REGFORCE \genblk1[875].rfrc ( .Q(L[875]), .A(V[875]), .E(fen));
Q_RELEASE_WEAK \genblk1[874].rrel ( .Q(L[874]), .E(ren));
Q_REGFORCE \genblk1[874].rfrc ( .Q(L[874]), .A(V[874]), .E(fen));
Q_RELEASE_WEAK \genblk1[873].rrel ( .Q(L[873]), .E(ren));
Q_REGFORCE \genblk1[873].rfrc ( .Q(L[873]), .A(V[873]), .E(fen));
Q_RELEASE_WEAK \genblk1[872].rrel ( .Q(L[872]), .E(ren));
Q_REGFORCE \genblk1[872].rfrc ( .Q(L[872]), .A(V[872]), .E(fen));
Q_RELEASE_WEAK \genblk1[871].rrel ( .Q(L[871]), .E(ren));
Q_REGFORCE \genblk1[871].rfrc ( .Q(L[871]), .A(V[871]), .E(fen));
Q_RELEASE_WEAK \genblk1[870].rrel ( .Q(L[870]), .E(ren));
Q_REGFORCE \genblk1[870].rfrc ( .Q(L[870]), .A(V[870]), .E(fen));
Q_RELEASE_WEAK \genblk1[869].rrel ( .Q(L[869]), .E(ren));
Q_REGFORCE \genblk1[869].rfrc ( .Q(L[869]), .A(V[869]), .E(fen));
Q_RELEASE_WEAK \genblk1[868].rrel ( .Q(L[868]), .E(ren));
Q_REGFORCE \genblk1[868].rfrc ( .Q(L[868]), .A(V[868]), .E(fen));
Q_RELEASE_WEAK \genblk1[867].rrel ( .Q(L[867]), .E(ren));
Q_REGFORCE \genblk1[867].rfrc ( .Q(L[867]), .A(V[867]), .E(fen));
Q_RELEASE_WEAK \genblk1[866].rrel ( .Q(L[866]), .E(ren));
Q_REGFORCE \genblk1[866].rfrc ( .Q(L[866]), .A(V[866]), .E(fen));
Q_RELEASE_WEAK \genblk1[865].rrel ( .Q(L[865]), .E(ren));
Q_REGFORCE \genblk1[865].rfrc ( .Q(L[865]), .A(V[865]), .E(fen));
Q_RELEASE_WEAK \genblk1[864].rrel ( .Q(L[864]), .E(ren));
Q_REGFORCE \genblk1[864].rfrc ( .Q(L[864]), .A(V[864]), .E(fen));
Q_RELEASE_WEAK \genblk1[863].rrel ( .Q(L[863]), .E(ren));
Q_REGFORCE \genblk1[863].rfrc ( .Q(L[863]), .A(V[863]), .E(fen));
Q_RELEASE_WEAK \genblk1[862].rrel ( .Q(L[862]), .E(ren));
Q_REGFORCE \genblk1[862].rfrc ( .Q(L[862]), .A(V[862]), .E(fen));
Q_RELEASE_WEAK \genblk1[861].rrel ( .Q(L[861]), .E(ren));
Q_REGFORCE \genblk1[861].rfrc ( .Q(L[861]), .A(V[861]), .E(fen));
Q_RELEASE_WEAK \genblk1[860].rrel ( .Q(L[860]), .E(ren));
Q_REGFORCE \genblk1[860].rfrc ( .Q(L[860]), .A(V[860]), .E(fen));
Q_RELEASE_WEAK \genblk1[859].rrel ( .Q(L[859]), .E(ren));
Q_REGFORCE \genblk1[859].rfrc ( .Q(L[859]), .A(V[859]), .E(fen));
Q_RELEASE_WEAK \genblk1[858].rrel ( .Q(L[858]), .E(ren));
Q_REGFORCE \genblk1[858].rfrc ( .Q(L[858]), .A(V[858]), .E(fen));
Q_RELEASE_WEAK \genblk1[857].rrel ( .Q(L[857]), .E(ren));
Q_REGFORCE \genblk1[857].rfrc ( .Q(L[857]), .A(V[857]), .E(fen));
Q_RELEASE_WEAK \genblk1[856].rrel ( .Q(L[856]), .E(ren));
Q_REGFORCE \genblk1[856].rfrc ( .Q(L[856]), .A(V[856]), .E(fen));
Q_RELEASE_WEAK \genblk1[855].rrel ( .Q(L[855]), .E(ren));
Q_REGFORCE \genblk1[855].rfrc ( .Q(L[855]), .A(V[855]), .E(fen));
Q_RELEASE_WEAK \genblk1[854].rrel ( .Q(L[854]), .E(ren));
Q_REGFORCE \genblk1[854].rfrc ( .Q(L[854]), .A(V[854]), .E(fen));
Q_RELEASE_WEAK \genblk1[853].rrel ( .Q(L[853]), .E(ren));
Q_REGFORCE \genblk1[853].rfrc ( .Q(L[853]), .A(V[853]), .E(fen));
Q_RELEASE_WEAK \genblk1[852].rrel ( .Q(L[852]), .E(ren));
Q_REGFORCE \genblk1[852].rfrc ( .Q(L[852]), .A(V[852]), .E(fen));
Q_RELEASE_WEAK \genblk1[851].rrel ( .Q(L[851]), .E(ren));
Q_REGFORCE \genblk1[851].rfrc ( .Q(L[851]), .A(V[851]), .E(fen));
Q_RELEASE_WEAK \genblk1[850].rrel ( .Q(L[850]), .E(ren));
Q_REGFORCE \genblk1[850].rfrc ( .Q(L[850]), .A(V[850]), .E(fen));
Q_RELEASE_WEAK \genblk1[849].rrel ( .Q(L[849]), .E(ren));
Q_REGFORCE \genblk1[849].rfrc ( .Q(L[849]), .A(V[849]), .E(fen));
Q_RELEASE_WEAK \genblk1[848].rrel ( .Q(L[848]), .E(ren));
Q_REGFORCE \genblk1[848].rfrc ( .Q(L[848]), .A(V[848]), .E(fen));
Q_RELEASE_WEAK \genblk1[847].rrel ( .Q(L[847]), .E(ren));
Q_REGFORCE \genblk1[847].rfrc ( .Q(L[847]), .A(V[847]), .E(fen));
Q_RELEASE_WEAK \genblk1[846].rrel ( .Q(L[846]), .E(ren));
Q_REGFORCE \genblk1[846].rfrc ( .Q(L[846]), .A(V[846]), .E(fen));
Q_RELEASE_WEAK \genblk1[845].rrel ( .Q(L[845]), .E(ren));
Q_REGFORCE \genblk1[845].rfrc ( .Q(L[845]), .A(V[845]), .E(fen));
Q_RELEASE_WEAK \genblk1[844].rrel ( .Q(L[844]), .E(ren));
Q_REGFORCE \genblk1[844].rfrc ( .Q(L[844]), .A(V[844]), .E(fen));
Q_RELEASE_WEAK \genblk1[843].rrel ( .Q(L[843]), .E(ren));
Q_REGFORCE \genblk1[843].rfrc ( .Q(L[843]), .A(V[843]), .E(fen));
Q_RELEASE_WEAK \genblk1[842].rrel ( .Q(L[842]), .E(ren));
Q_REGFORCE \genblk1[842].rfrc ( .Q(L[842]), .A(V[842]), .E(fen));
Q_RELEASE_WEAK \genblk1[841].rrel ( .Q(L[841]), .E(ren));
Q_REGFORCE \genblk1[841].rfrc ( .Q(L[841]), .A(V[841]), .E(fen));
Q_RELEASE_WEAK \genblk1[840].rrel ( .Q(L[840]), .E(ren));
Q_REGFORCE \genblk1[840].rfrc ( .Q(L[840]), .A(V[840]), .E(fen));
Q_RELEASE_WEAK \genblk1[839].rrel ( .Q(L[839]), .E(ren));
Q_REGFORCE \genblk1[839].rfrc ( .Q(L[839]), .A(V[839]), .E(fen));
Q_RELEASE_WEAK \genblk1[838].rrel ( .Q(L[838]), .E(ren));
Q_REGFORCE \genblk1[838].rfrc ( .Q(L[838]), .A(V[838]), .E(fen));
Q_RELEASE_WEAK \genblk1[837].rrel ( .Q(L[837]), .E(ren));
Q_REGFORCE \genblk1[837].rfrc ( .Q(L[837]), .A(V[837]), .E(fen));
Q_RELEASE_WEAK \genblk1[836].rrel ( .Q(L[836]), .E(ren));
Q_REGFORCE \genblk1[836].rfrc ( .Q(L[836]), .A(V[836]), .E(fen));
Q_RELEASE_WEAK \genblk1[835].rrel ( .Q(L[835]), .E(ren));
Q_REGFORCE \genblk1[835].rfrc ( .Q(L[835]), .A(V[835]), .E(fen));
Q_RELEASE_WEAK \genblk1[834].rrel ( .Q(L[834]), .E(ren));
Q_REGFORCE \genblk1[834].rfrc ( .Q(L[834]), .A(V[834]), .E(fen));
Q_RELEASE_WEAK \genblk1[833].rrel ( .Q(L[833]), .E(ren));
Q_REGFORCE \genblk1[833].rfrc ( .Q(L[833]), .A(V[833]), .E(fen));
Q_RELEASE_WEAK \genblk1[832].rrel ( .Q(L[832]), .E(ren));
Q_REGFORCE \genblk1[832].rfrc ( .Q(L[832]), .A(V[832]), .E(fen));
Q_RELEASE_WEAK \genblk1[831].rrel ( .Q(L[831]), .E(ren));
Q_REGFORCE \genblk1[831].rfrc ( .Q(L[831]), .A(V[831]), .E(fen));
Q_RELEASE_WEAK \genblk1[830].rrel ( .Q(L[830]), .E(ren));
Q_REGFORCE \genblk1[830].rfrc ( .Q(L[830]), .A(V[830]), .E(fen));
Q_RELEASE_WEAK \genblk1[829].rrel ( .Q(L[829]), .E(ren));
Q_REGFORCE \genblk1[829].rfrc ( .Q(L[829]), .A(V[829]), .E(fen));
Q_RELEASE_WEAK \genblk1[828].rrel ( .Q(L[828]), .E(ren));
Q_REGFORCE \genblk1[828].rfrc ( .Q(L[828]), .A(V[828]), .E(fen));
Q_RELEASE_WEAK \genblk1[827].rrel ( .Q(L[827]), .E(ren));
Q_REGFORCE \genblk1[827].rfrc ( .Q(L[827]), .A(V[827]), .E(fen));
Q_RELEASE_WEAK \genblk1[826].rrel ( .Q(L[826]), .E(ren));
Q_REGFORCE \genblk1[826].rfrc ( .Q(L[826]), .A(V[826]), .E(fen));
Q_RELEASE_WEAK \genblk1[825].rrel ( .Q(L[825]), .E(ren));
Q_REGFORCE \genblk1[825].rfrc ( .Q(L[825]), .A(V[825]), .E(fen));
Q_RELEASE_WEAK \genblk1[824].rrel ( .Q(L[824]), .E(ren));
Q_REGFORCE \genblk1[824].rfrc ( .Q(L[824]), .A(V[824]), .E(fen));
Q_RELEASE_WEAK \genblk1[823].rrel ( .Q(L[823]), .E(ren));
Q_REGFORCE \genblk1[823].rfrc ( .Q(L[823]), .A(V[823]), .E(fen));
Q_RELEASE_WEAK \genblk1[822].rrel ( .Q(L[822]), .E(ren));
Q_REGFORCE \genblk1[822].rfrc ( .Q(L[822]), .A(V[822]), .E(fen));
Q_RELEASE_WEAK \genblk1[821].rrel ( .Q(L[821]), .E(ren));
Q_REGFORCE \genblk1[821].rfrc ( .Q(L[821]), .A(V[821]), .E(fen));
Q_RELEASE_WEAK \genblk1[820].rrel ( .Q(L[820]), .E(ren));
Q_REGFORCE \genblk1[820].rfrc ( .Q(L[820]), .A(V[820]), .E(fen));
Q_RELEASE_WEAK \genblk1[819].rrel ( .Q(L[819]), .E(ren));
Q_REGFORCE \genblk1[819].rfrc ( .Q(L[819]), .A(V[819]), .E(fen));
Q_RELEASE_WEAK \genblk1[818].rrel ( .Q(L[818]), .E(ren));
Q_REGFORCE \genblk1[818].rfrc ( .Q(L[818]), .A(V[818]), .E(fen));
Q_RELEASE_WEAK \genblk1[817].rrel ( .Q(L[817]), .E(ren));
Q_REGFORCE \genblk1[817].rfrc ( .Q(L[817]), .A(V[817]), .E(fen));
Q_RELEASE_WEAK \genblk1[816].rrel ( .Q(L[816]), .E(ren));
Q_REGFORCE \genblk1[816].rfrc ( .Q(L[816]), .A(V[816]), .E(fen));
Q_RELEASE_WEAK \genblk1[815].rrel ( .Q(L[815]), .E(ren));
Q_REGFORCE \genblk1[815].rfrc ( .Q(L[815]), .A(V[815]), .E(fen));
Q_RELEASE_WEAK \genblk1[814].rrel ( .Q(L[814]), .E(ren));
Q_REGFORCE \genblk1[814].rfrc ( .Q(L[814]), .A(V[814]), .E(fen));
Q_RELEASE_WEAK \genblk1[813].rrel ( .Q(L[813]), .E(ren));
Q_REGFORCE \genblk1[813].rfrc ( .Q(L[813]), .A(V[813]), .E(fen));
Q_RELEASE_WEAK \genblk1[812].rrel ( .Q(L[812]), .E(ren));
Q_REGFORCE \genblk1[812].rfrc ( .Q(L[812]), .A(V[812]), .E(fen));
Q_RELEASE_WEAK \genblk1[811].rrel ( .Q(L[811]), .E(ren));
Q_REGFORCE \genblk1[811].rfrc ( .Q(L[811]), .A(V[811]), .E(fen));
Q_RELEASE_WEAK \genblk1[810].rrel ( .Q(L[810]), .E(ren));
Q_REGFORCE \genblk1[810].rfrc ( .Q(L[810]), .A(V[810]), .E(fen));
Q_RELEASE_WEAK \genblk1[809].rrel ( .Q(L[809]), .E(ren));
Q_REGFORCE \genblk1[809].rfrc ( .Q(L[809]), .A(V[809]), .E(fen));
Q_RELEASE_WEAK \genblk1[808].rrel ( .Q(L[808]), .E(ren));
Q_REGFORCE \genblk1[808].rfrc ( .Q(L[808]), .A(V[808]), .E(fen));
Q_RELEASE_WEAK \genblk1[807].rrel ( .Q(L[807]), .E(ren));
Q_REGFORCE \genblk1[807].rfrc ( .Q(L[807]), .A(V[807]), .E(fen));
Q_RELEASE_WEAK \genblk1[806].rrel ( .Q(L[806]), .E(ren));
Q_REGFORCE \genblk1[806].rfrc ( .Q(L[806]), .A(V[806]), .E(fen));
Q_RELEASE_WEAK \genblk1[805].rrel ( .Q(L[805]), .E(ren));
Q_REGFORCE \genblk1[805].rfrc ( .Q(L[805]), .A(V[805]), .E(fen));
Q_RELEASE_WEAK \genblk1[804].rrel ( .Q(L[804]), .E(ren));
Q_REGFORCE \genblk1[804].rfrc ( .Q(L[804]), .A(V[804]), .E(fen));
Q_RELEASE_WEAK \genblk1[803].rrel ( .Q(L[803]), .E(ren));
Q_REGFORCE \genblk1[803].rfrc ( .Q(L[803]), .A(V[803]), .E(fen));
Q_RELEASE_WEAK \genblk1[802].rrel ( .Q(L[802]), .E(ren));
Q_REGFORCE \genblk1[802].rfrc ( .Q(L[802]), .A(V[802]), .E(fen));
Q_RELEASE_WEAK \genblk1[801].rrel ( .Q(L[801]), .E(ren));
Q_REGFORCE \genblk1[801].rfrc ( .Q(L[801]), .A(V[801]), .E(fen));
Q_RELEASE_WEAK \genblk1[800].rrel ( .Q(L[800]), .E(ren));
Q_REGFORCE \genblk1[800].rfrc ( .Q(L[800]), .A(V[800]), .E(fen));
Q_RELEASE_WEAK \genblk1[799].rrel ( .Q(L[799]), .E(ren));
Q_REGFORCE \genblk1[799].rfrc ( .Q(L[799]), .A(V[799]), .E(fen));
Q_RELEASE_WEAK \genblk1[798].rrel ( .Q(L[798]), .E(ren));
Q_REGFORCE \genblk1[798].rfrc ( .Q(L[798]), .A(V[798]), .E(fen));
Q_RELEASE_WEAK \genblk1[797].rrel ( .Q(L[797]), .E(ren));
Q_REGFORCE \genblk1[797].rfrc ( .Q(L[797]), .A(V[797]), .E(fen));
Q_RELEASE_WEAK \genblk1[796].rrel ( .Q(L[796]), .E(ren));
Q_REGFORCE \genblk1[796].rfrc ( .Q(L[796]), .A(V[796]), .E(fen));
Q_RELEASE_WEAK \genblk1[795].rrel ( .Q(L[795]), .E(ren));
Q_REGFORCE \genblk1[795].rfrc ( .Q(L[795]), .A(V[795]), .E(fen));
Q_RELEASE_WEAK \genblk1[794].rrel ( .Q(L[794]), .E(ren));
Q_REGFORCE \genblk1[794].rfrc ( .Q(L[794]), .A(V[794]), .E(fen));
Q_RELEASE_WEAK \genblk1[793].rrel ( .Q(L[793]), .E(ren));
Q_REGFORCE \genblk1[793].rfrc ( .Q(L[793]), .A(V[793]), .E(fen));
Q_RELEASE_WEAK \genblk1[792].rrel ( .Q(L[792]), .E(ren));
Q_REGFORCE \genblk1[792].rfrc ( .Q(L[792]), .A(V[792]), .E(fen));
Q_RELEASE_WEAK \genblk1[791].rrel ( .Q(L[791]), .E(ren));
Q_REGFORCE \genblk1[791].rfrc ( .Q(L[791]), .A(V[791]), .E(fen));
Q_RELEASE_WEAK \genblk1[790].rrel ( .Q(L[790]), .E(ren));
Q_REGFORCE \genblk1[790].rfrc ( .Q(L[790]), .A(V[790]), .E(fen));
Q_RELEASE_WEAK \genblk1[789].rrel ( .Q(L[789]), .E(ren));
Q_REGFORCE \genblk1[789].rfrc ( .Q(L[789]), .A(V[789]), .E(fen));
Q_RELEASE_WEAK \genblk1[788].rrel ( .Q(L[788]), .E(ren));
Q_REGFORCE \genblk1[788].rfrc ( .Q(L[788]), .A(V[788]), .E(fen));
Q_RELEASE_WEAK \genblk1[787].rrel ( .Q(L[787]), .E(ren));
Q_REGFORCE \genblk1[787].rfrc ( .Q(L[787]), .A(V[787]), .E(fen));
Q_RELEASE_WEAK \genblk1[786].rrel ( .Q(L[786]), .E(ren));
Q_REGFORCE \genblk1[786].rfrc ( .Q(L[786]), .A(V[786]), .E(fen));
Q_RELEASE_WEAK \genblk1[785].rrel ( .Q(L[785]), .E(ren));
Q_REGFORCE \genblk1[785].rfrc ( .Q(L[785]), .A(V[785]), .E(fen));
Q_RELEASE_WEAK \genblk1[784].rrel ( .Q(L[784]), .E(ren));
Q_REGFORCE \genblk1[784].rfrc ( .Q(L[784]), .A(V[784]), .E(fen));
Q_RELEASE_WEAK \genblk1[783].rrel ( .Q(L[783]), .E(ren));
Q_REGFORCE \genblk1[783].rfrc ( .Q(L[783]), .A(V[783]), .E(fen));
Q_RELEASE_WEAK \genblk1[782].rrel ( .Q(L[782]), .E(ren));
Q_REGFORCE \genblk1[782].rfrc ( .Q(L[782]), .A(V[782]), .E(fen));
Q_RELEASE_WEAK \genblk1[781].rrel ( .Q(L[781]), .E(ren));
Q_REGFORCE \genblk1[781].rfrc ( .Q(L[781]), .A(V[781]), .E(fen));
Q_RELEASE_WEAK \genblk1[780].rrel ( .Q(L[780]), .E(ren));
Q_REGFORCE \genblk1[780].rfrc ( .Q(L[780]), .A(V[780]), .E(fen));
Q_RELEASE_WEAK \genblk1[779].rrel ( .Q(L[779]), .E(ren));
Q_REGFORCE \genblk1[779].rfrc ( .Q(L[779]), .A(V[779]), .E(fen));
Q_RELEASE_WEAK \genblk1[778].rrel ( .Q(L[778]), .E(ren));
Q_REGFORCE \genblk1[778].rfrc ( .Q(L[778]), .A(V[778]), .E(fen));
Q_RELEASE_WEAK \genblk1[777].rrel ( .Q(L[777]), .E(ren));
Q_REGFORCE \genblk1[777].rfrc ( .Q(L[777]), .A(V[777]), .E(fen));
Q_RELEASE_WEAK \genblk1[776].rrel ( .Q(L[776]), .E(ren));
Q_REGFORCE \genblk1[776].rfrc ( .Q(L[776]), .A(V[776]), .E(fen));
Q_RELEASE_WEAK \genblk1[775].rrel ( .Q(L[775]), .E(ren));
Q_REGFORCE \genblk1[775].rfrc ( .Q(L[775]), .A(V[775]), .E(fen));
Q_RELEASE_WEAK \genblk1[774].rrel ( .Q(L[774]), .E(ren));
Q_REGFORCE \genblk1[774].rfrc ( .Q(L[774]), .A(V[774]), .E(fen));
Q_RELEASE_WEAK \genblk1[773].rrel ( .Q(L[773]), .E(ren));
Q_REGFORCE \genblk1[773].rfrc ( .Q(L[773]), .A(V[773]), .E(fen));
Q_RELEASE_WEAK \genblk1[772].rrel ( .Q(L[772]), .E(ren));
Q_REGFORCE \genblk1[772].rfrc ( .Q(L[772]), .A(V[772]), .E(fen));
Q_RELEASE_WEAK \genblk1[771].rrel ( .Q(L[771]), .E(ren));
Q_REGFORCE \genblk1[771].rfrc ( .Q(L[771]), .A(V[771]), .E(fen));
Q_RELEASE_WEAK \genblk1[770].rrel ( .Q(L[770]), .E(ren));
Q_REGFORCE \genblk1[770].rfrc ( .Q(L[770]), .A(V[770]), .E(fen));
Q_RELEASE_WEAK \genblk1[769].rrel ( .Q(L[769]), .E(ren));
Q_REGFORCE \genblk1[769].rfrc ( .Q(L[769]), .A(V[769]), .E(fen));
Q_RELEASE_WEAK \genblk1[768].rrel ( .Q(L[768]), .E(ren));
Q_REGFORCE \genblk1[768].rfrc ( .Q(L[768]), .A(V[768]), .E(fen));
Q_RELEASE_WEAK \genblk1[767].rrel ( .Q(L[767]), .E(ren));
Q_REGFORCE \genblk1[767].rfrc ( .Q(L[767]), .A(V[767]), .E(fen));
Q_RELEASE_WEAK \genblk1[766].rrel ( .Q(L[766]), .E(ren));
Q_REGFORCE \genblk1[766].rfrc ( .Q(L[766]), .A(V[766]), .E(fen));
Q_RELEASE_WEAK \genblk1[765].rrel ( .Q(L[765]), .E(ren));
Q_REGFORCE \genblk1[765].rfrc ( .Q(L[765]), .A(V[765]), .E(fen));
Q_RELEASE_WEAK \genblk1[764].rrel ( .Q(L[764]), .E(ren));
Q_REGFORCE \genblk1[764].rfrc ( .Q(L[764]), .A(V[764]), .E(fen));
Q_RELEASE_WEAK \genblk1[763].rrel ( .Q(L[763]), .E(ren));
Q_REGFORCE \genblk1[763].rfrc ( .Q(L[763]), .A(V[763]), .E(fen));
Q_RELEASE_WEAK \genblk1[762].rrel ( .Q(L[762]), .E(ren));
Q_REGFORCE \genblk1[762].rfrc ( .Q(L[762]), .A(V[762]), .E(fen));
Q_RELEASE_WEAK \genblk1[761].rrel ( .Q(L[761]), .E(ren));
Q_REGFORCE \genblk1[761].rfrc ( .Q(L[761]), .A(V[761]), .E(fen));
Q_RELEASE_WEAK \genblk1[760].rrel ( .Q(L[760]), .E(ren));
Q_REGFORCE \genblk1[760].rfrc ( .Q(L[760]), .A(V[760]), .E(fen));
Q_RELEASE_WEAK \genblk1[759].rrel ( .Q(L[759]), .E(ren));
Q_REGFORCE \genblk1[759].rfrc ( .Q(L[759]), .A(V[759]), .E(fen));
Q_RELEASE_WEAK \genblk1[758].rrel ( .Q(L[758]), .E(ren));
Q_REGFORCE \genblk1[758].rfrc ( .Q(L[758]), .A(V[758]), .E(fen));
Q_RELEASE_WEAK \genblk1[757].rrel ( .Q(L[757]), .E(ren));
Q_REGFORCE \genblk1[757].rfrc ( .Q(L[757]), .A(V[757]), .E(fen));
Q_RELEASE_WEAK \genblk1[756].rrel ( .Q(L[756]), .E(ren));
Q_REGFORCE \genblk1[756].rfrc ( .Q(L[756]), .A(V[756]), .E(fen));
Q_RELEASE_WEAK \genblk1[755].rrel ( .Q(L[755]), .E(ren));
Q_REGFORCE \genblk1[755].rfrc ( .Q(L[755]), .A(V[755]), .E(fen));
Q_RELEASE_WEAK \genblk1[754].rrel ( .Q(L[754]), .E(ren));
Q_REGFORCE \genblk1[754].rfrc ( .Q(L[754]), .A(V[754]), .E(fen));
Q_RELEASE_WEAK \genblk1[753].rrel ( .Q(L[753]), .E(ren));
Q_REGFORCE \genblk1[753].rfrc ( .Q(L[753]), .A(V[753]), .E(fen));
Q_RELEASE_WEAK \genblk1[752].rrel ( .Q(L[752]), .E(ren));
Q_REGFORCE \genblk1[752].rfrc ( .Q(L[752]), .A(V[752]), .E(fen));
Q_RELEASE_WEAK \genblk1[751].rrel ( .Q(L[751]), .E(ren));
Q_REGFORCE \genblk1[751].rfrc ( .Q(L[751]), .A(V[751]), .E(fen));
Q_RELEASE_WEAK \genblk1[750].rrel ( .Q(L[750]), .E(ren));
Q_REGFORCE \genblk1[750].rfrc ( .Q(L[750]), .A(V[750]), .E(fen));
Q_RELEASE_WEAK \genblk1[749].rrel ( .Q(L[749]), .E(ren));
Q_REGFORCE \genblk1[749].rfrc ( .Q(L[749]), .A(V[749]), .E(fen));
Q_RELEASE_WEAK \genblk1[748].rrel ( .Q(L[748]), .E(ren));
Q_REGFORCE \genblk1[748].rfrc ( .Q(L[748]), .A(V[748]), .E(fen));
Q_RELEASE_WEAK \genblk1[747].rrel ( .Q(L[747]), .E(ren));
Q_REGFORCE \genblk1[747].rfrc ( .Q(L[747]), .A(V[747]), .E(fen));
Q_RELEASE_WEAK \genblk1[746].rrel ( .Q(L[746]), .E(ren));
Q_REGFORCE \genblk1[746].rfrc ( .Q(L[746]), .A(V[746]), .E(fen));
Q_RELEASE_WEAK \genblk1[745].rrel ( .Q(L[745]), .E(ren));
Q_REGFORCE \genblk1[745].rfrc ( .Q(L[745]), .A(V[745]), .E(fen));
Q_RELEASE_WEAK \genblk1[744].rrel ( .Q(L[744]), .E(ren));
Q_REGFORCE \genblk1[744].rfrc ( .Q(L[744]), .A(V[744]), .E(fen));
Q_RELEASE_WEAK \genblk1[743].rrel ( .Q(L[743]), .E(ren));
Q_REGFORCE \genblk1[743].rfrc ( .Q(L[743]), .A(V[743]), .E(fen));
Q_RELEASE_WEAK \genblk1[742].rrel ( .Q(L[742]), .E(ren));
Q_REGFORCE \genblk1[742].rfrc ( .Q(L[742]), .A(V[742]), .E(fen));
Q_RELEASE_WEAK \genblk1[741].rrel ( .Q(L[741]), .E(ren));
Q_REGFORCE \genblk1[741].rfrc ( .Q(L[741]), .A(V[741]), .E(fen));
Q_RELEASE_WEAK \genblk1[740].rrel ( .Q(L[740]), .E(ren));
Q_REGFORCE \genblk1[740].rfrc ( .Q(L[740]), .A(V[740]), .E(fen));
Q_RELEASE_WEAK \genblk1[739].rrel ( .Q(L[739]), .E(ren));
Q_REGFORCE \genblk1[739].rfrc ( .Q(L[739]), .A(V[739]), .E(fen));
Q_RELEASE_WEAK \genblk1[738].rrel ( .Q(L[738]), .E(ren));
Q_REGFORCE \genblk1[738].rfrc ( .Q(L[738]), .A(V[738]), .E(fen));
Q_RELEASE_WEAK \genblk1[737].rrel ( .Q(L[737]), .E(ren));
Q_REGFORCE \genblk1[737].rfrc ( .Q(L[737]), .A(V[737]), .E(fen));
Q_RELEASE_WEAK \genblk1[736].rrel ( .Q(L[736]), .E(ren));
Q_REGFORCE \genblk1[736].rfrc ( .Q(L[736]), .A(V[736]), .E(fen));
Q_RELEASE_WEAK \genblk1[735].rrel ( .Q(L[735]), .E(ren));
Q_REGFORCE \genblk1[735].rfrc ( .Q(L[735]), .A(V[735]), .E(fen));
Q_RELEASE_WEAK \genblk1[734].rrel ( .Q(L[734]), .E(ren));
Q_REGFORCE \genblk1[734].rfrc ( .Q(L[734]), .A(V[734]), .E(fen));
Q_RELEASE_WEAK \genblk1[733].rrel ( .Q(L[733]), .E(ren));
Q_REGFORCE \genblk1[733].rfrc ( .Q(L[733]), .A(V[733]), .E(fen));
Q_RELEASE_WEAK \genblk1[732].rrel ( .Q(L[732]), .E(ren));
Q_REGFORCE \genblk1[732].rfrc ( .Q(L[732]), .A(V[732]), .E(fen));
Q_RELEASE_WEAK \genblk1[731].rrel ( .Q(L[731]), .E(ren));
Q_REGFORCE \genblk1[731].rfrc ( .Q(L[731]), .A(V[731]), .E(fen));
Q_RELEASE_WEAK \genblk1[730].rrel ( .Q(L[730]), .E(ren));
Q_REGFORCE \genblk1[730].rfrc ( .Q(L[730]), .A(V[730]), .E(fen));
Q_RELEASE_WEAK \genblk1[729].rrel ( .Q(L[729]), .E(ren));
Q_REGFORCE \genblk1[729].rfrc ( .Q(L[729]), .A(V[729]), .E(fen));
Q_RELEASE_WEAK \genblk1[728].rrel ( .Q(L[728]), .E(ren));
Q_REGFORCE \genblk1[728].rfrc ( .Q(L[728]), .A(V[728]), .E(fen));
Q_RELEASE_WEAK \genblk1[727].rrel ( .Q(L[727]), .E(ren));
Q_REGFORCE \genblk1[727].rfrc ( .Q(L[727]), .A(V[727]), .E(fen));
Q_RELEASE_WEAK \genblk1[726].rrel ( .Q(L[726]), .E(ren));
Q_REGFORCE \genblk1[726].rfrc ( .Q(L[726]), .A(V[726]), .E(fen));
Q_RELEASE_WEAK \genblk1[725].rrel ( .Q(L[725]), .E(ren));
Q_REGFORCE \genblk1[725].rfrc ( .Q(L[725]), .A(V[725]), .E(fen));
Q_RELEASE_WEAK \genblk1[724].rrel ( .Q(L[724]), .E(ren));
Q_REGFORCE \genblk1[724].rfrc ( .Q(L[724]), .A(V[724]), .E(fen));
Q_RELEASE_WEAK \genblk1[723].rrel ( .Q(L[723]), .E(ren));
Q_REGFORCE \genblk1[723].rfrc ( .Q(L[723]), .A(V[723]), .E(fen));
Q_RELEASE_WEAK \genblk1[722].rrel ( .Q(L[722]), .E(ren));
Q_REGFORCE \genblk1[722].rfrc ( .Q(L[722]), .A(V[722]), .E(fen));
Q_RELEASE_WEAK \genblk1[721].rrel ( .Q(L[721]), .E(ren));
Q_REGFORCE \genblk1[721].rfrc ( .Q(L[721]), .A(V[721]), .E(fen));
Q_RELEASE_WEAK \genblk1[720].rrel ( .Q(L[720]), .E(ren));
Q_REGFORCE \genblk1[720].rfrc ( .Q(L[720]), .A(V[720]), .E(fen));
Q_RELEASE_WEAK \genblk1[719].rrel ( .Q(L[719]), .E(ren));
Q_REGFORCE \genblk1[719].rfrc ( .Q(L[719]), .A(V[719]), .E(fen));
Q_RELEASE_WEAK \genblk1[718].rrel ( .Q(L[718]), .E(ren));
Q_REGFORCE \genblk1[718].rfrc ( .Q(L[718]), .A(V[718]), .E(fen));
Q_RELEASE_WEAK \genblk1[717].rrel ( .Q(L[717]), .E(ren));
Q_REGFORCE \genblk1[717].rfrc ( .Q(L[717]), .A(V[717]), .E(fen));
Q_RELEASE_WEAK \genblk1[716].rrel ( .Q(L[716]), .E(ren));
Q_REGFORCE \genblk1[716].rfrc ( .Q(L[716]), .A(V[716]), .E(fen));
Q_RELEASE_WEAK \genblk1[715].rrel ( .Q(L[715]), .E(ren));
Q_REGFORCE \genblk1[715].rfrc ( .Q(L[715]), .A(V[715]), .E(fen));
Q_RELEASE_WEAK \genblk1[714].rrel ( .Q(L[714]), .E(ren));
Q_REGFORCE \genblk1[714].rfrc ( .Q(L[714]), .A(V[714]), .E(fen));
Q_RELEASE_WEAK \genblk1[713].rrel ( .Q(L[713]), .E(ren));
Q_REGFORCE \genblk1[713].rfrc ( .Q(L[713]), .A(V[713]), .E(fen));
Q_RELEASE_WEAK \genblk1[712].rrel ( .Q(L[712]), .E(ren));
Q_REGFORCE \genblk1[712].rfrc ( .Q(L[712]), .A(V[712]), .E(fen));
Q_RELEASE_WEAK \genblk1[711].rrel ( .Q(L[711]), .E(ren));
Q_REGFORCE \genblk1[711].rfrc ( .Q(L[711]), .A(V[711]), .E(fen));
Q_RELEASE_WEAK \genblk1[710].rrel ( .Q(L[710]), .E(ren));
Q_REGFORCE \genblk1[710].rfrc ( .Q(L[710]), .A(V[710]), .E(fen));
Q_RELEASE_WEAK \genblk1[709].rrel ( .Q(L[709]), .E(ren));
Q_REGFORCE \genblk1[709].rfrc ( .Q(L[709]), .A(V[709]), .E(fen));
Q_RELEASE_WEAK \genblk1[708].rrel ( .Q(L[708]), .E(ren));
Q_REGFORCE \genblk1[708].rfrc ( .Q(L[708]), .A(V[708]), .E(fen));
Q_RELEASE_WEAK \genblk1[707].rrel ( .Q(L[707]), .E(ren));
Q_REGFORCE \genblk1[707].rfrc ( .Q(L[707]), .A(V[707]), .E(fen));
Q_RELEASE_WEAK \genblk1[706].rrel ( .Q(L[706]), .E(ren));
Q_REGFORCE \genblk1[706].rfrc ( .Q(L[706]), .A(V[706]), .E(fen));
Q_RELEASE_WEAK \genblk1[705].rrel ( .Q(L[705]), .E(ren));
Q_REGFORCE \genblk1[705].rfrc ( .Q(L[705]), .A(V[705]), .E(fen));
Q_RELEASE_WEAK \genblk1[704].rrel ( .Q(L[704]), .E(ren));
Q_REGFORCE \genblk1[704].rfrc ( .Q(L[704]), .A(V[704]), .E(fen));
Q_RELEASE_WEAK \genblk1[703].rrel ( .Q(L[703]), .E(ren));
Q_REGFORCE \genblk1[703].rfrc ( .Q(L[703]), .A(V[703]), .E(fen));
Q_RELEASE_WEAK \genblk1[702].rrel ( .Q(L[702]), .E(ren));
Q_REGFORCE \genblk1[702].rfrc ( .Q(L[702]), .A(V[702]), .E(fen));
Q_RELEASE_WEAK \genblk1[701].rrel ( .Q(L[701]), .E(ren));
Q_REGFORCE \genblk1[701].rfrc ( .Q(L[701]), .A(V[701]), .E(fen));
Q_RELEASE_WEAK \genblk1[700].rrel ( .Q(L[700]), .E(ren));
Q_REGFORCE \genblk1[700].rfrc ( .Q(L[700]), .A(V[700]), .E(fen));
Q_RELEASE_WEAK \genblk1[699].rrel ( .Q(L[699]), .E(ren));
Q_REGFORCE \genblk1[699].rfrc ( .Q(L[699]), .A(V[699]), .E(fen));
Q_RELEASE_WEAK \genblk1[698].rrel ( .Q(L[698]), .E(ren));
Q_REGFORCE \genblk1[698].rfrc ( .Q(L[698]), .A(V[698]), .E(fen));
Q_RELEASE_WEAK \genblk1[697].rrel ( .Q(L[697]), .E(ren));
Q_REGFORCE \genblk1[697].rfrc ( .Q(L[697]), .A(V[697]), .E(fen));
Q_RELEASE_WEAK \genblk1[696].rrel ( .Q(L[696]), .E(ren));
Q_REGFORCE \genblk1[696].rfrc ( .Q(L[696]), .A(V[696]), .E(fen));
Q_RELEASE_WEAK \genblk1[695].rrel ( .Q(L[695]), .E(ren));
Q_REGFORCE \genblk1[695].rfrc ( .Q(L[695]), .A(V[695]), .E(fen));
Q_RELEASE_WEAK \genblk1[694].rrel ( .Q(L[694]), .E(ren));
Q_REGFORCE \genblk1[694].rfrc ( .Q(L[694]), .A(V[694]), .E(fen));
Q_RELEASE_WEAK \genblk1[693].rrel ( .Q(L[693]), .E(ren));
Q_REGFORCE \genblk1[693].rfrc ( .Q(L[693]), .A(V[693]), .E(fen));
Q_RELEASE_WEAK \genblk1[692].rrel ( .Q(L[692]), .E(ren));
Q_REGFORCE \genblk1[692].rfrc ( .Q(L[692]), .A(V[692]), .E(fen));
Q_RELEASE_WEAK \genblk1[691].rrel ( .Q(L[691]), .E(ren));
Q_REGFORCE \genblk1[691].rfrc ( .Q(L[691]), .A(V[691]), .E(fen));
Q_RELEASE_WEAK \genblk1[690].rrel ( .Q(L[690]), .E(ren));
Q_REGFORCE \genblk1[690].rfrc ( .Q(L[690]), .A(V[690]), .E(fen));
Q_RELEASE_WEAK \genblk1[689].rrel ( .Q(L[689]), .E(ren));
Q_REGFORCE \genblk1[689].rfrc ( .Q(L[689]), .A(V[689]), .E(fen));
Q_RELEASE_WEAK \genblk1[688].rrel ( .Q(L[688]), .E(ren));
Q_REGFORCE \genblk1[688].rfrc ( .Q(L[688]), .A(V[688]), .E(fen));
Q_RELEASE_WEAK \genblk1[687].rrel ( .Q(L[687]), .E(ren));
Q_REGFORCE \genblk1[687].rfrc ( .Q(L[687]), .A(V[687]), .E(fen));
Q_RELEASE_WEAK \genblk1[686].rrel ( .Q(L[686]), .E(ren));
Q_REGFORCE \genblk1[686].rfrc ( .Q(L[686]), .A(V[686]), .E(fen));
Q_RELEASE_WEAK \genblk1[685].rrel ( .Q(L[685]), .E(ren));
Q_REGFORCE \genblk1[685].rfrc ( .Q(L[685]), .A(V[685]), .E(fen));
Q_RELEASE_WEAK \genblk1[684].rrel ( .Q(L[684]), .E(ren));
Q_REGFORCE \genblk1[684].rfrc ( .Q(L[684]), .A(V[684]), .E(fen));
Q_RELEASE_WEAK \genblk1[683].rrel ( .Q(L[683]), .E(ren));
Q_REGFORCE \genblk1[683].rfrc ( .Q(L[683]), .A(V[683]), .E(fen));
Q_RELEASE_WEAK \genblk1[682].rrel ( .Q(L[682]), .E(ren));
Q_REGFORCE \genblk1[682].rfrc ( .Q(L[682]), .A(V[682]), .E(fen));
Q_RELEASE_WEAK \genblk1[681].rrel ( .Q(L[681]), .E(ren));
Q_REGFORCE \genblk1[681].rfrc ( .Q(L[681]), .A(V[681]), .E(fen));
Q_RELEASE_WEAK \genblk1[680].rrel ( .Q(L[680]), .E(ren));
Q_REGFORCE \genblk1[680].rfrc ( .Q(L[680]), .A(V[680]), .E(fen));
Q_RELEASE_WEAK \genblk1[679].rrel ( .Q(L[679]), .E(ren));
Q_REGFORCE \genblk1[679].rfrc ( .Q(L[679]), .A(V[679]), .E(fen));
Q_RELEASE_WEAK \genblk1[678].rrel ( .Q(L[678]), .E(ren));
Q_REGFORCE \genblk1[678].rfrc ( .Q(L[678]), .A(V[678]), .E(fen));
Q_RELEASE_WEAK \genblk1[677].rrel ( .Q(L[677]), .E(ren));
Q_REGFORCE \genblk1[677].rfrc ( .Q(L[677]), .A(V[677]), .E(fen));
Q_RELEASE_WEAK \genblk1[676].rrel ( .Q(L[676]), .E(ren));
Q_REGFORCE \genblk1[676].rfrc ( .Q(L[676]), .A(V[676]), .E(fen));
Q_RELEASE_WEAK \genblk1[675].rrel ( .Q(L[675]), .E(ren));
Q_REGFORCE \genblk1[675].rfrc ( .Q(L[675]), .A(V[675]), .E(fen));
Q_RELEASE_WEAK \genblk1[674].rrel ( .Q(L[674]), .E(ren));
Q_REGFORCE \genblk1[674].rfrc ( .Q(L[674]), .A(V[674]), .E(fen));
Q_RELEASE_WEAK \genblk1[673].rrel ( .Q(L[673]), .E(ren));
Q_REGFORCE \genblk1[673].rfrc ( .Q(L[673]), .A(V[673]), .E(fen));
Q_RELEASE_WEAK \genblk1[672].rrel ( .Q(L[672]), .E(ren));
Q_REGFORCE \genblk1[672].rfrc ( .Q(L[672]), .A(V[672]), .E(fen));
Q_RELEASE_WEAK \genblk1[671].rrel ( .Q(L[671]), .E(ren));
Q_REGFORCE \genblk1[671].rfrc ( .Q(L[671]), .A(V[671]), .E(fen));
Q_RELEASE_WEAK \genblk1[670].rrel ( .Q(L[670]), .E(ren));
Q_REGFORCE \genblk1[670].rfrc ( .Q(L[670]), .A(V[670]), .E(fen));
Q_RELEASE_WEAK \genblk1[669].rrel ( .Q(L[669]), .E(ren));
Q_REGFORCE \genblk1[669].rfrc ( .Q(L[669]), .A(V[669]), .E(fen));
Q_RELEASE_WEAK \genblk1[668].rrel ( .Q(L[668]), .E(ren));
Q_REGFORCE \genblk1[668].rfrc ( .Q(L[668]), .A(V[668]), .E(fen));
Q_RELEASE_WEAK \genblk1[667].rrel ( .Q(L[667]), .E(ren));
Q_REGFORCE \genblk1[667].rfrc ( .Q(L[667]), .A(V[667]), .E(fen));
Q_RELEASE_WEAK \genblk1[666].rrel ( .Q(L[666]), .E(ren));
Q_REGFORCE \genblk1[666].rfrc ( .Q(L[666]), .A(V[666]), .E(fen));
Q_RELEASE_WEAK \genblk1[665].rrel ( .Q(L[665]), .E(ren));
Q_REGFORCE \genblk1[665].rfrc ( .Q(L[665]), .A(V[665]), .E(fen));
Q_RELEASE_WEAK \genblk1[664].rrel ( .Q(L[664]), .E(ren));
Q_REGFORCE \genblk1[664].rfrc ( .Q(L[664]), .A(V[664]), .E(fen));
Q_RELEASE_WEAK \genblk1[663].rrel ( .Q(L[663]), .E(ren));
Q_REGFORCE \genblk1[663].rfrc ( .Q(L[663]), .A(V[663]), .E(fen));
Q_RELEASE_WEAK \genblk1[662].rrel ( .Q(L[662]), .E(ren));
Q_REGFORCE \genblk1[662].rfrc ( .Q(L[662]), .A(V[662]), .E(fen));
Q_RELEASE_WEAK \genblk1[661].rrel ( .Q(L[661]), .E(ren));
Q_REGFORCE \genblk1[661].rfrc ( .Q(L[661]), .A(V[661]), .E(fen));
Q_RELEASE_WEAK \genblk1[660].rrel ( .Q(L[660]), .E(ren));
Q_REGFORCE \genblk1[660].rfrc ( .Q(L[660]), .A(V[660]), .E(fen));
Q_RELEASE_WEAK \genblk1[659].rrel ( .Q(L[659]), .E(ren));
Q_REGFORCE \genblk1[659].rfrc ( .Q(L[659]), .A(V[659]), .E(fen));
Q_RELEASE_WEAK \genblk1[658].rrel ( .Q(L[658]), .E(ren));
Q_REGFORCE \genblk1[658].rfrc ( .Q(L[658]), .A(V[658]), .E(fen));
Q_RELEASE_WEAK \genblk1[657].rrel ( .Q(L[657]), .E(ren));
Q_REGFORCE \genblk1[657].rfrc ( .Q(L[657]), .A(V[657]), .E(fen));
Q_RELEASE_WEAK \genblk1[656].rrel ( .Q(L[656]), .E(ren));
Q_REGFORCE \genblk1[656].rfrc ( .Q(L[656]), .A(V[656]), .E(fen));
Q_RELEASE_WEAK \genblk1[655].rrel ( .Q(L[655]), .E(ren));
Q_REGFORCE \genblk1[655].rfrc ( .Q(L[655]), .A(V[655]), .E(fen));
Q_RELEASE_WEAK \genblk1[654].rrel ( .Q(L[654]), .E(ren));
Q_REGFORCE \genblk1[654].rfrc ( .Q(L[654]), .A(V[654]), .E(fen));
Q_RELEASE_WEAK \genblk1[653].rrel ( .Q(L[653]), .E(ren));
Q_REGFORCE \genblk1[653].rfrc ( .Q(L[653]), .A(V[653]), .E(fen));
Q_RELEASE_WEAK \genblk1[652].rrel ( .Q(L[652]), .E(ren));
Q_REGFORCE \genblk1[652].rfrc ( .Q(L[652]), .A(V[652]), .E(fen));
Q_RELEASE_WEAK \genblk1[651].rrel ( .Q(L[651]), .E(ren));
Q_REGFORCE \genblk1[651].rfrc ( .Q(L[651]), .A(V[651]), .E(fen));
Q_RELEASE_WEAK \genblk1[650].rrel ( .Q(L[650]), .E(ren));
Q_REGFORCE \genblk1[650].rfrc ( .Q(L[650]), .A(V[650]), .E(fen));
Q_RELEASE_WEAK \genblk1[649].rrel ( .Q(L[649]), .E(ren));
Q_REGFORCE \genblk1[649].rfrc ( .Q(L[649]), .A(V[649]), .E(fen));
Q_RELEASE_WEAK \genblk1[648].rrel ( .Q(L[648]), .E(ren));
Q_REGFORCE \genblk1[648].rfrc ( .Q(L[648]), .A(V[648]), .E(fen));
Q_RELEASE_WEAK \genblk1[647].rrel ( .Q(L[647]), .E(ren));
Q_REGFORCE \genblk1[647].rfrc ( .Q(L[647]), .A(V[647]), .E(fen));
Q_RELEASE_WEAK \genblk1[646].rrel ( .Q(L[646]), .E(ren));
Q_REGFORCE \genblk1[646].rfrc ( .Q(L[646]), .A(V[646]), .E(fen));
Q_RELEASE_WEAK \genblk1[645].rrel ( .Q(L[645]), .E(ren));
Q_REGFORCE \genblk1[645].rfrc ( .Q(L[645]), .A(V[645]), .E(fen));
Q_RELEASE_WEAK \genblk1[644].rrel ( .Q(L[644]), .E(ren));
Q_REGFORCE \genblk1[644].rfrc ( .Q(L[644]), .A(V[644]), .E(fen));
Q_RELEASE_WEAK \genblk1[643].rrel ( .Q(L[643]), .E(ren));
Q_REGFORCE \genblk1[643].rfrc ( .Q(L[643]), .A(V[643]), .E(fen));
Q_RELEASE_WEAK \genblk1[642].rrel ( .Q(L[642]), .E(ren));
Q_REGFORCE \genblk1[642].rfrc ( .Q(L[642]), .A(V[642]), .E(fen));
Q_RELEASE_WEAK \genblk1[641].rrel ( .Q(L[641]), .E(ren));
Q_REGFORCE \genblk1[641].rfrc ( .Q(L[641]), .A(V[641]), .E(fen));
Q_RELEASE_WEAK \genblk1[640].rrel ( .Q(L[640]), .E(ren));
Q_REGFORCE \genblk1[640].rfrc ( .Q(L[640]), .A(V[640]), .E(fen));
Q_RELEASE_WEAK \genblk1[639].rrel ( .Q(L[639]), .E(ren));
Q_REGFORCE \genblk1[639].rfrc ( .Q(L[639]), .A(V[639]), .E(fen));
Q_RELEASE_WEAK \genblk1[638].rrel ( .Q(L[638]), .E(ren));
Q_REGFORCE \genblk1[638].rfrc ( .Q(L[638]), .A(V[638]), .E(fen));
Q_RELEASE_WEAK \genblk1[637].rrel ( .Q(L[637]), .E(ren));
Q_REGFORCE \genblk1[637].rfrc ( .Q(L[637]), .A(V[637]), .E(fen));
Q_RELEASE_WEAK \genblk1[636].rrel ( .Q(L[636]), .E(ren));
Q_REGFORCE \genblk1[636].rfrc ( .Q(L[636]), .A(V[636]), .E(fen));
Q_RELEASE_WEAK \genblk1[635].rrel ( .Q(L[635]), .E(ren));
Q_REGFORCE \genblk1[635].rfrc ( .Q(L[635]), .A(V[635]), .E(fen));
Q_RELEASE_WEAK \genblk1[634].rrel ( .Q(L[634]), .E(ren));
Q_REGFORCE \genblk1[634].rfrc ( .Q(L[634]), .A(V[634]), .E(fen));
Q_RELEASE_WEAK \genblk1[633].rrel ( .Q(L[633]), .E(ren));
Q_REGFORCE \genblk1[633].rfrc ( .Q(L[633]), .A(V[633]), .E(fen));
Q_RELEASE_WEAK \genblk1[632].rrel ( .Q(L[632]), .E(ren));
Q_REGFORCE \genblk1[632].rfrc ( .Q(L[632]), .A(V[632]), .E(fen));
Q_RELEASE_WEAK \genblk1[631].rrel ( .Q(L[631]), .E(ren));
Q_REGFORCE \genblk1[631].rfrc ( .Q(L[631]), .A(V[631]), .E(fen));
Q_RELEASE_WEAK \genblk1[630].rrel ( .Q(L[630]), .E(ren));
Q_REGFORCE \genblk1[630].rfrc ( .Q(L[630]), .A(V[630]), .E(fen));
Q_RELEASE_WEAK \genblk1[629].rrel ( .Q(L[629]), .E(ren));
Q_REGFORCE \genblk1[629].rfrc ( .Q(L[629]), .A(V[629]), .E(fen));
Q_RELEASE_WEAK \genblk1[628].rrel ( .Q(L[628]), .E(ren));
Q_REGFORCE \genblk1[628].rfrc ( .Q(L[628]), .A(V[628]), .E(fen));
Q_RELEASE_WEAK \genblk1[627].rrel ( .Q(L[627]), .E(ren));
Q_REGFORCE \genblk1[627].rfrc ( .Q(L[627]), .A(V[627]), .E(fen));
Q_RELEASE_WEAK \genblk1[626].rrel ( .Q(L[626]), .E(ren));
Q_REGFORCE \genblk1[626].rfrc ( .Q(L[626]), .A(V[626]), .E(fen));
Q_RELEASE_WEAK \genblk1[625].rrel ( .Q(L[625]), .E(ren));
Q_REGFORCE \genblk1[625].rfrc ( .Q(L[625]), .A(V[625]), .E(fen));
Q_RELEASE_WEAK \genblk1[624].rrel ( .Q(L[624]), .E(ren));
Q_REGFORCE \genblk1[624].rfrc ( .Q(L[624]), .A(V[624]), .E(fen));
Q_RELEASE_WEAK \genblk1[623].rrel ( .Q(L[623]), .E(ren));
Q_REGFORCE \genblk1[623].rfrc ( .Q(L[623]), .A(V[623]), .E(fen));
Q_RELEASE_WEAK \genblk1[622].rrel ( .Q(L[622]), .E(ren));
Q_REGFORCE \genblk1[622].rfrc ( .Q(L[622]), .A(V[622]), .E(fen));
Q_RELEASE_WEAK \genblk1[621].rrel ( .Q(L[621]), .E(ren));
Q_REGFORCE \genblk1[621].rfrc ( .Q(L[621]), .A(V[621]), .E(fen));
Q_RELEASE_WEAK \genblk1[620].rrel ( .Q(L[620]), .E(ren));
Q_REGFORCE \genblk1[620].rfrc ( .Q(L[620]), .A(V[620]), .E(fen));
Q_RELEASE_WEAK \genblk1[619].rrel ( .Q(L[619]), .E(ren));
Q_REGFORCE \genblk1[619].rfrc ( .Q(L[619]), .A(V[619]), .E(fen));
Q_RELEASE_WEAK \genblk1[618].rrel ( .Q(L[618]), .E(ren));
Q_REGFORCE \genblk1[618].rfrc ( .Q(L[618]), .A(V[618]), .E(fen));
Q_RELEASE_WEAK \genblk1[617].rrel ( .Q(L[617]), .E(ren));
Q_REGFORCE \genblk1[617].rfrc ( .Q(L[617]), .A(V[617]), .E(fen));
Q_RELEASE_WEAK \genblk1[616].rrel ( .Q(L[616]), .E(ren));
Q_REGFORCE \genblk1[616].rfrc ( .Q(L[616]), .A(V[616]), .E(fen));
Q_RELEASE_WEAK \genblk1[615].rrel ( .Q(L[615]), .E(ren));
Q_REGFORCE \genblk1[615].rfrc ( .Q(L[615]), .A(V[615]), .E(fen));
Q_RELEASE_WEAK \genblk1[614].rrel ( .Q(L[614]), .E(ren));
Q_REGFORCE \genblk1[614].rfrc ( .Q(L[614]), .A(V[614]), .E(fen));
Q_RELEASE_WEAK \genblk1[613].rrel ( .Q(L[613]), .E(ren));
Q_REGFORCE \genblk1[613].rfrc ( .Q(L[613]), .A(V[613]), .E(fen));
Q_RELEASE_WEAK \genblk1[612].rrel ( .Q(L[612]), .E(ren));
Q_REGFORCE \genblk1[612].rfrc ( .Q(L[612]), .A(V[612]), .E(fen));
Q_RELEASE_WEAK \genblk1[611].rrel ( .Q(L[611]), .E(ren));
Q_REGFORCE \genblk1[611].rfrc ( .Q(L[611]), .A(V[611]), .E(fen));
Q_RELEASE_WEAK \genblk1[610].rrel ( .Q(L[610]), .E(ren));
Q_REGFORCE \genblk1[610].rfrc ( .Q(L[610]), .A(V[610]), .E(fen));
Q_RELEASE_WEAK \genblk1[609].rrel ( .Q(L[609]), .E(ren));
Q_REGFORCE \genblk1[609].rfrc ( .Q(L[609]), .A(V[609]), .E(fen));
Q_RELEASE_WEAK \genblk1[608].rrel ( .Q(L[608]), .E(ren));
Q_REGFORCE \genblk1[608].rfrc ( .Q(L[608]), .A(V[608]), .E(fen));
Q_RELEASE_WEAK \genblk1[607].rrel ( .Q(L[607]), .E(ren));
Q_REGFORCE \genblk1[607].rfrc ( .Q(L[607]), .A(V[607]), .E(fen));
Q_RELEASE_WEAK \genblk1[606].rrel ( .Q(L[606]), .E(ren));
Q_REGFORCE \genblk1[606].rfrc ( .Q(L[606]), .A(V[606]), .E(fen));
Q_RELEASE_WEAK \genblk1[605].rrel ( .Q(L[605]), .E(ren));
Q_REGFORCE \genblk1[605].rfrc ( .Q(L[605]), .A(V[605]), .E(fen));
Q_RELEASE_WEAK \genblk1[604].rrel ( .Q(L[604]), .E(ren));
Q_REGFORCE \genblk1[604].rfrc ( .Q(L[604]), .A(V[604]), .E(fen));
Q_RELEASE_WEAK \genblk1[603].rrel ( .Q(L[603]), .E(ren));
Q_REGFORCE \genblk1[603].rfrc ( .Q(L[603]), .A(V[603]), .E(fen));
Q_RELEASE_WEAK \genblk1[602].rrel ( .Q(L[602]), .E(ren));
Q_REGFORCE \genblk1[602].rfrc ( .Q(L[602]), .A(V[602]), .E(fen));
Q_RELEASE_WEAK \genblk1[601].rrel ( .Q(L[601]), .E(ren));
Q_REGFORCE \genblk1[601].rfrc ( .Q(L[601]), .A(V[601]), .E(fen));
Q_RELEASE_WEAK \genblk1[600].rrel ( .Q(L[600]), .E(ren));
Q_REGFORCE \genblk1[600].rfrc ( .Q(L[600]), .A(V[600]), .E(fen));
Q_RELEASE_WEAK \genblk1[599].rrel ( .Q(L[599]), .E(ren));
Q_REGFORCE \genblk1[599].rfrc ( .Q(L[599]), .A(V[599]), .E(fen));
Q_RELEASE_WEAK \genblk1[598].rrel ( .Q(L[598]), .E(ren));
Q_REGFORCE \genblk1[598].rfrc ( .Q(L[598]), .A(V[598]), .E(fen));
Q_RELEASE_WEAK \genblk1[597].rrel ( .Q(L[597]), .E(ren));
Q_REGFORCE \genblk1[597].rfrc ( .Q(L[597]), .A(V[597]), .E(fen));
Q_RELEASE_WEAK \genblk1[596].rrel ( .Q(L[596]), .E(ren));
Q_REGFORCE \genblk1[596].rfrc ( .Q(L[596]), .A(V[596]), .E(fen));
Q_RELEASE_WEAK \genblk1[595].rrel ( .Q(L[595]), .E(ren));
Q_REGFORCE \genblk1[595].rfrc ( .Q(L[595]), .A(V[595]), .E(fen));
Q_RELEASE_WEAK \genblk1[594].rrel ( .Q(L[594]), .E(ren));
Q_REGFORCE \genblk1[594].rfrc ( .Q(L[594]), .A(V[594]), .E(fen));
Q_RELEASE_WEAK \genblk1[593].rrel ( .Q(L[593]), .E(ren));
Q_REGFORCE \genblk1[593].rfrc ( .Q(L[593]), .A(V[593]), .E(fen));
Q_RELEASE_WEAK \genblk1[592].rrel ( .Q(L[592]), .E(ren));
Q_REGFORCE \genblk1[592].rfrc ( .Q(L[592]), .A(V[592]), .E(fen));
Q_RELEASE_WEAK \genblk1[591].rrel ( .Q(L[591]), .E(ren));
Q_REGFORCE \genblk1[591].rfrc ( .Q(L[591]), .A(V[591]), .E(fen));
Q_RELEASE_WEAK \genblk1[590].rrel ( .Q(L[590]), .E(ren));
Q_REGFORCE \genblk1[590].rfrc ( .Q(L[590]), .A(V[590]), .E(fen));
Q_RELEASE_WEAK \genblk1[589].rrel ( .Q(L[589]), .E(ren));
Q_REGFORCE \genblk1[589].rfrc ( .Q(L[589]), .A(V[589]), .E(fen));
Q_RELEASE_WEAK \genblk1[588].rrel ( .Q(L[588]), .E(ren));
Q_REGFORCE \genblk1[588].rfrc ( .Q(L[588]), .A(V[588]), .E(fen));
Q_RELEASE_WEAK \genblk1[587].rrel ( .Q(L[587]), .E(ren));
Q_REGFORCE \genblk1[587].rfrc ( .Q(L[587]), .A(V[587]), .E(fen));
Q_RELEASE_WEAK \genblk1[586].rrel ( .Q(L[586]), .E(ren));
Q_REGFORCE \genblk1[586].rfrc ( .Q(L[586]), .A(V[586]), .E(fen));
Q_RELEASE_WEAK \genblk1[585].rrel ( .Q(L[585]), .E(ren));
Q_REGFORCE \genblk1[585].rfrc ( .Q(L[585]), .A(V[585]), .E(fen));
Q_RELEASE_WEAK \genblk1[584].rrel ( .Q(L[584]), .E(ren));
Q_REGFORCE \genblk1[584].rfrc ( .Q(L[584]), .A(V[584]), .E(fen));
Q_RELEASE_WEAK \genblk1[583].rrel ( .Q(L[583]), .E(ren));
Q_REGFORCE \genblk1[583].rfrc ( .Q(L[583]), .A(V[583]), .E(fen));
Q_RELEASE_WEAK \genblk1[582].rrel ( .Q(L[582]), .E(ren));
Q_REGFORCE \genblk1[582].rfrc ( .Q(L[582]), .A(V[582]), .E(fen));
Q_RELEASE_WEAK \genblk1[581].rrel ( .Q(L[581]), .E(ren));
Q_REGFORCE \genblk1[581].rfrc ( .Q(L[581]), .A(V[581]), .E(fen));
Q_RELEASE_WEAK \genblk1[580].rrel ( .Q(L[580]), .E(ren));
Q_REGFORCE \genblk1[580].rfrc ( .Q(L[580]), .A(V[580]), .E(fen));
Q_RELEASE_WEAK \genblk1[579].rrel ( .Q(L[579]), .E(ren));
Q_REGFORCE \genblk1[579].rfrc ( .Q(L[579]), .A(V[579]), .E(fen));
Q_RELEASE_WEAK \genblk1[578].rrel ( .Q(L[578]), .E(ren));
Q_REGFORCE \genblk1[578].rfrc ( .Q(L[578]), .A(V[578]), .E(fen));
Q_RELEASE_WEAK \genblk1[577].rrel ( .Q(L[577]), .E(ren));
Q_REGFORCE \genblk1[577].rfrc ( .Q(L[577]), .A(V[577]), .E(fen));
Q_RELEASE_WEAK \genblk1[576].rrel ( .Q(L[576]), .E(ren));
Q_REGFORCE \genblk1[576].rfrc ( .Q(L[576]), .A(V[576]), .E(fen));
Q_RELEASE_WEAK \genblk1[575].rrel ( .Q(L[575]), .E(ren));
Q_REGFORCE \genblk1[575].rfrc ( .Q(L[575]), .A(V[575]), .E(fen));
Q_RELEASE_WEAK \genblk1[574].rrel ( .Q(L[574]), .E(ren));
Q_REGFORCE \genblk1[574].rfrc ( .Q(L[574]), .A(V[574]), .E(fen));
Q_RELEASE_WEAK \genblk1[573].rrel ( .Q(L[573]), .E(ren));
Q_REGFORCE \genblk1[573].rfrc ( .Q(L[573]), .A(V[573]), .E(fen));
Q_RELEASE_WEAK \genblk1[572].rrel ( .Q(L[572]), .E(ren));
Q_REGFORCE \genblk1[572].rfrc ( .Q(L[572]), .A(V[572]), .E(fen));
Q_RELEASE_WEAK \genblk1[571].rrel ( .Q(L[571]), .E(ren));
Q_REGFORCE \genblk1[571].rfrc ( .Q(L[571]), .A(V[571]), .E(fen));
Q_RELEASE_WEAK \genblk1[570].rrel ( .Q(L[570]), .E(ren));
Q_REGFORCE \genblk1[570].rfrc ( .Q(L[570]), .A(V[570]), .E(fen));
Q_RELEASE_WEAK \genblk1[569].rrel ( .Q(L[569]), .E(ren));
Q_REGFORCE \genblk1[569].rfrc ( .Q(L[569]), .A(V[569]), .E(fen));
Q_RELEASE_WEAK \genblk1[568].rrel ( .Q(L[568]), .E(ren));
Q_REGFORCE \genblk1[568].rfrc ( .Q(L[568]), .A(V[568]), .E(fen));
Q_RELEASE_WEAK \genblk1[567].rrel ( .Q(L[567]), .E(ren));
Q_REGFORCE \genblk1[567].rfrc ( .Q(L[567]), .A(V[567]), .E(fen));
Q_RELEASE_WEAK \genblk1[566].rrel ( .Q(L[566]), .E(ren));
Q_REGFORCE \genblk1[566].rfrc ( .Q(L[566]), .A(V[566]), .E(fen));
Q_RELEASE_WEAK \genblk1[565].rrel ( .Q(L[565]), .E(ren));
Q_REGFORCE \genblk1[565].rfrc ( .Q(L[565]), .A(V[565]), .E(fen));
Q_RELEASE_WEAK \genblk1[564].rrel ( .Q(L[564]), .E(ren));
Q_REGFORCE \genblk1[564].rfrc ( .Q(L[564]), .A(V[564]), .E(fen));
Q_RELEASE_WEAK \genblk1[563].rrel ( .Q(L[563]), .E(ren));
Q_REGFORCE \genblk1[563].rfrc ( .Q(L[563]), .A(V[563]), .E(fen));
Q_RELEASE_WEAK \genblk1[562].rrel ( .Q(L[562]), .E(ren));
Q_REGFORCE \genblk1[562].rfrc ( .Q(L[562]), .A(V[562]), .E(fen));
Q_RELEASE_WEAK \genblk1[561].rrel ( .Q(L[561]), .E(ren));
Q_REGFORCE \genblk1[561].rfrc ( .Q(L[561]), .A(V[561]), .E(fen));
Q_RELEASE_WEAK \genblk1[560].rrel ( .Q(L[560]), .E(ren));
Q_REGFORCE \genblk1[560].rfrc ( .Q(L[560]), .A(V[560]), .E(fen));
Q_RELEASE_WEAK \genblk1[559].rrel ( .Q(L[559]), .E(ren));
Q_REGFORCE \genblk1[559].rfrc ( .Q(L[559]), .A(V[559]), .E(fen));
Q_RELEASE_WEAK \genblk1[558].rrel ( .Q(L[558]), .E(ren));
Q_REGFORCE \genblk1[558].rfrc ( .Q(L[558]), .A(V[558]), .E(fen));
Q_RELEASE_WEAK \genblk1[557].rrel ( .Q(L[557]), .E(ren));
Q_REGFORCE \genblk1[557].rfrc ( .Q(L[557]), .A(V[557]), .E(fen));
Q_RELEASE_WEAK \genblk1[556].rrel ( .Q(L[556]), .E(ren));
Q_REGFORCE \genblk1[556].rfrc ( .Q(L[556]), .A(V[556]), .E(fen));
Q_RELEASE_WEAK \genblk1[555].rrel ( .Q(L[555]), .E(ren));
Q_REGFORCE \genblk1[555].rfrc ( .Q(L[555]), .A(V[555]), .E(fen));
Q_RELEASE_WEAK \genblk1[554].rrel ( .Q(L[554]), .E(ren));
Q_REGFORCE \genblk1[554].rfrc ( .Q(L[554]), .A(V[554]), .E(fen));
Q_RELEASE_WEAK \genblk1[553].rrel ( .Q(L[553]), .E(ren));
Q_REGFORCE \genblk1[553].rfrc ( .Q(L[553]), .A(V[553]), .E(fen));
Q_RELEASE_WEAK \genblk1[552].rrel ( .Q(L[552]), .E(ren));
Q_REGFORCE \genblk1[552].rfrc ( .Q(L[552]), .A(V[552]), .E(fen));
Q_RELEASE_WEAK \genblk1[551].rrel ( .Q(L[551]), .E(ren));
Q_REGFORCE \genblk1[551].rfrc ( .Q(L[551]), .A(V[551]), .E(fen));
Q_RELEASE_WEAK \genblk1[550].rrel ( .Q(L[550]), .E(ren));
Q_REGFORCE \genblk1[550].rfrc ( .Q(L[550]), .A(V[550]), .E(fen));
Q_RELEASE_WEAK \genblk1[549].rrel ( .Q(L[549]), .E(ren));
Q_REGFORCE \genblk1[549].rfrc ( .Q(L[549]), .A(V[549]), .E(fen));
Q_RELEASE_WEAK \genblk1[548].rrel ( .Q(L[548]), .E(ren));
Q_REGFORCE \genblk1[548].rfrc ( .Q(L[548]), .A(V[548]), .E(fen));
Q_RELEASE_WEAK \genblk1[547].rrel ( .Q(L[547]), .E(ren));
Q_REGFORCE \genblk1[547].rfrc ( .Q(L[547]), .A(V[547]), .E(fen));
Q_RELEASE_WEAK \genblk1[546].rrel ( .Q(L[546]), .E(ren));
Q_REGFORCE \genblk1[546].rfrc ( .Q(L[546]), .A(V[546]), .E(fen));
Q_RELEASE_WEAK \genblk1[545].rrel ( .Q(L[545]), .E(ren));
Q_REGFORCE \genblk1[545].rfrc ( .Q(L[545]), .A(V[545]), .E(fen));
Q_RELEASE_WEAK \genblk1[544].rrel ( .Q(L[544]), .E(ren));
Q_REGFORCE \genblk1[544].rfrc ( .Q(L[544]), .A(V[544]), .E(fen));
Q_RELEASE_WEAK \genblk1[543].rrel ( .Q(L[543]), .E(ren));
Q_REGFORCE \genblk1[543].rfrc ( .Q(L[543]), .A(V[543]), .E(fen));
Q_RELEASE_WEAK \genblk1[542].rrel ( .Q(L[542]), .E(ren));
Q_REGFORCE \genblk1[542].rfrc ( .Q(L[542]), .A(V[542]), .E(fen));
Q_RELEASE_WEAK \genblk1[541].rrel ( .Q(L[541]), .E(ren));
Q_REGFORCE \genblk1[541].rfrc ( .Q(L[541]), .A(V[541]), .E(fen));
Q_RELEASE_WEAK \genblk1[540].rrel ( .Q(L[540]), .E(ren));
Q_REGFORCE \genblk1[540].rfrc ( .Q(L[540]), .A(V[540]), .E(fen));
Q_RELEASE_WEAK \genblk1[539].rrel ( .Q(L[539]), .E(ren));
Q_REGFORCE \genblk1[539].rfrc ( .Q(L[539]), .A(V[539]), .E(fen));
Q_RELEASE_WEAK \genblk1[538].rrel ( .Q(L[538]), .E(ren));
Q_REGFORCE \genblk1[538].rfrc ( .Q(L[538]), .A(V[538]), .E(fen));
Q_RELEASE_WEAK \genblk1[537].rrel ( .Q(L[537]), .E(ren));
Q_REGFORCE \genblk1[537].rfrc ( .Q(L[537]), .A(V[537]), .E(fen));
Q_RELEASE_WEAK \genblk1[536].rrel ( .Q(L[536]), .E(ren));
Q_REGFORCE \genblk1[536].rfrc ( .Q(L[536]), .A(V[536]), .E(fen));
Q_RELEASE_WEAK \genblk1[535].rrel ( .Q(L[535]), .E(ren));
Q_REGFORCE \genblk1[535].rfrc ( .Q(L[535]), .A(V[535]), .E(fen));
Q_RELEASE_WEAK \genblk1[534].rrel ( .Q(L[534]), .E(ren));
Q_REGFORCE \genblk1[534].rfrc ( .Q(L[534]), .A(V[534]), .E(fen));
Q_RELEASE_WEAK \genblk1[533].rrel ( .Q(L[533]), .E(ren));
Q_REGFORCE \genblk1[533].rfrc ( .Q(L[533]), .A(V[533]), .E(fen));
Q_RELEASE_WEAK \genblk1[532].rrel ( .Q(L[532]), .E(ren));
Q_REGFORCE \genblk1[532].rfrc ( .Q(L[532]), .A(V[532]), .E(fen));
Q_RELEASE_WEAK \genblk1[531].rrel ( .Q(L[531]), .E(ren));
Q_REGFORCE \genblk1[531].rfrc ( .Q(L[531]), .A(V[531]), .E(fen));
Q_RELEASE_WEAK \genblk1[530].rrel ( .Q(L[530]), .E(ren));
Q_REGFORCE \genblk1[530].rfrc ( .Q(L[530]), .A(V[530]), .E(fen));
Q_RELEASE_WEAK \genblk1[529].rrel ( .Q(L[529]), .E(ren));
Q_REGFORCE \genblk1[529].rfrc ( .Q(L[529]), .A(V[529]), .E(fen));
Q_RELEASE_WEAK \genblk1[528].rrel ( .Q(L[528]), .E(ren));
Q_REGFORCE \genblk1[528].rfrc ( .Q(L[528]), .A(V[528]), .E(fen));
Q_RELEASE_WEAK \genblk1[527].rrel ( .Q(L[527]), .E(ren));
Q_REGFORCE \genblk1[527].rfrc ( .Q(L[527]), .A(V[527]), .E(fen));
Q_RELEASE_WEAK \genblk1[526].rrel ( .Q(L[526]), .E(ren));
Q_REGFORCE \genblk1[526].rfrc ( .Q(L[526]), .A(V[526]), .E(fen));
Q_RELEASE_WEAK \genblk1[525].rrel ( .Q(L[525]), .E(ren));
Q_REGFORCE \genblk1[525].rfrc ( .Q(L[525]), .A(V[525]), .E(fen));
Q_RELEASE_WEAK \genblk1[524].rrel ( .Q(L[524]), .E(ren));
Q_REGFORCE \genblk1[524].rfrc ( .Q(L[524]), .A(V[524]), .E(fen));
Q_RELEASE_WEAK \genblk1[523].rrel ( .Q(L[523]), .E(ren));
Q_REGFORCE \genblk1[523].rfrc ( .Q(L[523]), .A(V[523]), .E(fen));
Q_RELEASE_WEAK \genblk1[522].rrel ( .Q(L[522]), .E(ren));
Q_REGFORCE \genblk1[522].rfrc ( .Q(L[522]), .A(V[522]), .E(fen));
Q_RELEASE_WEAK \genblk1[521].rrel ( .Q(L[521]), .E(ren));
Q_REGFORCE \genblk1[521].rfrc ( .Q(L[521]), .A(V[521]), .E(fen));
Q_RELEASE_WEAK \genblk1[520].rrel ( .Q(L[520]), .E(ren));
Q_REGFORCE \genblk1[520].rfrc ( .Q(L[520]), .A(V[520]), .E(fen));
Q_RELEASE_WEAK \genblk1[519].rrel ( .Q(L[519]), .E(ren));
Q_REGFORCE \genblk1[519].rfrc ( .Q(L[519]), .A(V[519]), .E(fen));
Q_RELEASE_WEAK \genblk1[518].rrel ( .Q(L[518]), .E(ren));
Q_REGFORCE \genblk1[518].rfrc ( .Q(L[518]), .A(V[518]), .E(fen));
Q_RELEASE_WEAK \genblk1[517].rrel ( .Q(L[517]), .E(ren));
Q_REGFORCE \genblk1[517].rfrc ( .Q(L[517]), .A(V[517]), .E(fen));
Q_RELEASE_WEAK \genblk1[516].rrel ( .Q(L[516]), .E(ren));
Q_REGFORCE \genblk1[516].rfrc ( .Q(L[516]), .A(V[516]), .E(fen));
Q_RELEASE_WEAK \genblk1[515].rrel ( .Q(L[515]), .E(ren));
Q_REGFORCE \genblk1[515].rfrc ( .Q(L[515]), .A(V[515]), .E(fen));
Q_RELEASE_WEAK \genblk1[514].rrel ( .Q(L[514]), .E(ren));
Q_REGFORCE \genblk1[514].rfrc ( .Q(L[514]), .A(V[514]), .E(fen));
Q_RELEASE_WEAK \genblk1[513].rrel ( .Q(L[513]), .E(ren));
Q_REGFORCE \genblk1[513].rfrc ( .Q(L[513]), .A(V[513]), .E(fen));
Q_RELEASE_WEAK \genblk1[512].rrel ( .Q(L[512]), .E(ren));
Q_REGFORCE \genblk1[512].rfrc ( .Q(L[512]), .A(V[512]), .E(fen));
Q_RELEASE_WEAK \genblk1[511].rrel ( .Q(L[511]), .E(ren));
Q_REGFORCE \genblk1[511].rfrc ( .Q(L[511]), .A(V[511]), .E(fen));
Q_RELEASE_WEAK \genblk1[510].rrel ( .Q(L[510]), .E(ren));
Q_REGFORCE \genblk1[510].rfrc ( .Q(L[510]), .A(V[510]), .E(fen));
Q_RELEASE_WEAK \genblk1[509].rrel ( .Q(L[509]), .E(ren));
Q_REGFORCE \genblk1[509].rfrc ( .Q(L[509]), .A(V[509]), .E(fen));
Q_RELEASE_WEAK \genblk1[508].rrel ( .Q(L[508]), .E(ren));
Q_REGFORCE \genblk1[508].rfrc ( .Q(L[508]), .A(V[508]), .E(fen));
Q_RELEASE_WEAK \genblk1[507].rrel ( .Q(L[507]), .E(ren));
Q_REGFORCE \genblk1[507].rfrc ( .Q(L[507]), .A(V[507]), .E(fen));
Q_RELEASE_WEAK \genblk1[506].rrel ( .Q(L[506]), .E(ren));
Q_REGFORCE \genblk1[506].rfrc ( .Q(L[506]), .A(V[506]), .E(fen));
Q_RELEASE_WEAK \genblk1[505].rrel ( .Q(L[505]), .E(ren));
Q_REGFORCE \genblk1[505].rfrc ( .Q(L[505]), .A(V[505]), .E(fen));
Q_RELEASE_WEAK \genblk1[504].rrel ( .Q(L[504]), .E(ren));
Q_REGFORCE \genblk1[504].rfrc ( .Q(L[504]), .A(V[504]), .E(fen));
Q_RELEASE_WEAK \genblk1[503].rrel ( .Q(L[503]), .E(ren));
Q_REGFORCE \genblk1[503].rfrc ( .Q(L[503]), .A(V[503]), .E(fen));
Q_RELEASE_WEAK \genblk1[502].rrel ( .Q(L[502]), .E(ren));
Q_REGFORCE \genblk1[502].rfrc ( .Q(L[502]), .A(V[502]), .E(fen));
Q_RELEASE_WEAK \genblk1[501].rrel ( .Q(L[501]), .E(ren));
Q_REGFORCE \genblk1[501].rfrc ( .Q(L[501]), .A(V[501]), .E(fen));
Q_RELEASE_WEAK \genblk1[500].rrel ( .Q(L[500]), .E(ren));
Q_REGFORCE \genblk1[500].rfrc ( .Q(L[500]), .A(V[500]), .E(fen));
Q_RELEASE_WEAK \genblk1[499].rrel ( .Q(L[499]), .E(ren));
Q_REGFORCE \genblk1[499].rfrc ( .Q(L[499]), .A(V[499]), .E(fen));
Q_RELEASE_WEAK \genblk1[498].rrel ( .Q(L[498]), .E(ren));
Q_REGFORCE \genblk1[498].rfrc ( .Q(L[498]), .A(V[498]), .E(fen));
Q_RELEASE_WEAK \genblk1[497].rrel ( .Q(L[497]), .E(ren));
Q_REGFORCE \genblk1[497].rfrc ( .Q(L[497]), .A(V[497]), .E(fen));
Q_RELEASE_WEAK \genblk1[496].rrel ( .Q(L[496]), .E(ren));
Q_REGFORCE \genblk1[496].rfrc ( .Q(L[496]), .A(V[496]), .E(fen));
Q_RELEASE_WEAK \genblk1[495].rrel ( .Q(L[495]), .E(ren));
Q_REGFORCE \genblk1[495].rfrc ( .Q(L[495]), .A(V[495]), .E(fen));
Q_RELEASE_WEAK \genblk1[494].rrel ( .Q(L[494]), .E(ren));
Q_REGFORCE \genblk1[494].rfrc ( .Q(L[494]), .A(V[494]), .E(fen));
Q_RELEASE_WEAK \genblk1[493].rrel ( .Q(L[493]), .E(ren));
Q_REGFORCE \genblk1[493].rfrc ( .Q(L[493]), .A(V[493]), .E(fen));
Q_RELEASE_WEAK \genblk1[492].rrel ( .Q(L[492]), .E(ren));
Q_REGFORCE \genblk1[492].rfrc ( .Q(L[492]), .A(V[492]), .E(fen));
Q_RELEASE_WEAK \genblk1[491].rrel ( .Q(L[491]), .E(ren));
Q_REGFORCE \genblk1[491].rfrc ( .Q(L[491]), .A(V[491]), .E(fen));
Q_RELEASE_WEAK \genblk1[490].rrel ( .Q(L[490]), .E(ren));
Q_REGFORCE \genblk1[490].rfrc ( .Q(L[490]), .A(V[490]), .E(fen));
Q_RELEASE_WEAK \genblk1[489].rrel ( .Q(L[489]), .E(ren));
Q_REGFORCE \genblk1[489].rfrc ( .Q(L[489]), .A(V[489]), .E(fen));
Q_RELEASE_WEAK \genblk1[488].rrel ( .Q(L[488]), .E(ren));
Q_REGFORCE \genblk1[488].rfrc ( .Q(L[488]), .A(V[488]), .E(fen));
Q_RELEASE_WEAK \genblk1[487].rrel ( .Q(L[487]), .E(ren));
Q_REGFORCE \genblk1[487].rfrc ( .Q(L[487]), .A(V[487]), .E(fen));
Q_RELEASE_WEAK \genblk1[486].rrel ( .Q(L[486]), .E(ren));
Q_REGFORCE \genblk1[486].rfrc ( .Q(L[486]), .A(V[486]), .E(fen));
Q_RELEASE_WEAK \genblk1[485].rrel ( .Q(L[485]), .E(ren));
Q_REGFORCE \genblk1[485].rfrc ( .Q(L[485]), .A(V[485]), .E(fen));
Q_RELEASE_WEAK \genblk1[484].rrel ( .Q(L[484]), .E(ren));
Q_REGFORCE \genblk1[484].rfrc ( .Q(L[484]), .A(V[484]), .E(fen));
Q_RELEASE_WEAK \genblk1[483].rrel ( .Q(L[483]), .E(ren));
Q_REGFORCE \genblk1[483].rfrc ( .Q(L[483]), .A(V[483]), .E(fen));
Q_RELEASE_WEAK \genblk1[482].rrel ( .Q(L[482]), .E(ren));
Q_REGFORCE \genblk1[482].rfrc ( .Q(L[482]), .A(V[482]), .E(fen));
Q_RELEASE_WEAK \genblk1[481].rrel ( .Q(L[481]), .E(ren));
Q_REGFORCE \genblk1[481].rfrc ( .Q(L[481]), .A(V[481]), .E(fen));
Q_RELEASE_WEAK \genblk1[480].rrel ( .Q(L[480]), .E(ren));
Q_REGFORCE \genblk1[480].rfrc ( .Q(L[480]), .A(V[480]), .E(fen));
Q_RELEASE_WEAK \genblk1[479].rrel ( .Q(L[479]), .E(ren));
Q_REGFORCE \genblk1[479].rfrc ( .Q(L[479]), .A(V[479]), .E(fen));
Q_RELEASE_WEAK \genblk1[478].rrel ( .Q(L[478]), .E(ren));
Q_REGFORCE \genblk1[478].rfrc ( .Q(L[478]), .A(V[478]), .E(fen));
Q_RELEASE_WEAK \genblk1[477].rrel ( .Q(L[477]), .E(ren));
Q_REGFORCE \genblk1[477].rfrc ( .Q(L[477]), .A(V[477]), .E(fen));
Q_RELEASE_WEAK \genblk1[476].rrel ( .Q(L[476]), .E(ren));
Q_REGFORCE \genblk1[476].rfrc ( .Q(L[476]), .A(V[476]), .E(fen));
Q_RELEASE_WEAK \genblk1[475].rrel ( .Q(L[475]), .E(ren));
Q_REGFORCE \genblk1[475].rfrc ( .Q(L[475]), .A(V[475]), .E(fen));
Q_RELEASE_WEAK \genblk1[474].rrel ( .Q(L[474]), .E(ren));
Q_REGFORCE \genblk1[474].rfrc ( .Q(L[474]), .A(V[474]), .E(fen));
Q_RELEASE_WEAK \genblk1[473].rrel ( .Q(L[473]), .E(ren));
Q_REGFORCE \genblk1[473].rfrc ( .Q(L[473]), .A(V[473]), .E(fen));
Q_RELEASE_WEAK \genblk1[472].rrel ( .Q(L[472]), .E(ren));
Q_REGFORCE \genblk1[472].rfrc ( .Q(L[472]), .A(V[472]), .E(fen));
Q_RELEASE_WEAK \genblk1[471].rrel ( .Q(L[471]), .E(ren));
Q_REGFORCE \genblk1[471].rfrc ( .Q(L[471]), .A(V[471]), .E(fen));
Q_RELEASE_WEAK \genblk1[470].rrel ( .Q(L[470]), .E(ren));
Q_REGFORCE \genblk1[470].rfrc ( .Q(L[470]), .A(V[470]), .E(fen));
Q_RELEASE_WEAK \genblk1[469].rrel ( .Q(L[469]), .E(ren));
Q_REGFORCE \genblk1[469].rfrc ( .Q(L[469]), .A(V[469]), .E(fen));
Q_RELEASE_WEAK \genblk1[468].rrel ( .Q(L[468]), .E(ren));
Q_REGFORCE \genblk1[468].rfrc ( .Q(L[468]), .A(V[468]), .E(fen));
Q_RELEASE_WEAK \genblk1[467].rrel ( .Q(L[467]), .E(ren));
Q_REGFORCE \genblk1[467].rfrc ( .Q(L[467]), .A(V[467]), .E(fen));
Q_RELEASE_WEAK \genblk1[466].rrel ( .Q(L[466]), .E(ren));
Q_REGFORCE \genblk1[466].rfrc ( .Q(L[466]), .A(V[466]), .E(fen));
Q_RELEASE_WEAK \genblk1[465].rrel ( .Q(L[465]), .E(ren));
Q_REGFORCE \genblk1[465].rfrc ( .Q(L[465]), .A(V[465]), .E(fen));
Q_RELEASE_WEAK \genblk1[464].rrel ( .Q(L[464]), .E(ren));
Q_REGFORCE \genblk1[464].rfrc ( .Q(L[464]), .A(V[464]), .E(fen));
Q_RELEASE_WEAK \genblk1[463].rrel ( .Q(L[463]), .E(ren));
Q_REGFORCE \genblk1[463].rfrc ( .Q(L[463]), .A(V[463]), .E(fen));
Q_RELEASE_WEAK \genblk1[462].rrel ( .Q(L[462]), .E(ren));
Q_REGFORCE \genblk1[462].rfrc ( .Q(L[462]), .A(V[462]), .E(fen));
Q_RELEASE_WEAK \genblk1[461].rrel ( .Q(L[461]), .E(ren));
Q_REGFORCE \genblk1[461].rfrc ( .Q(L[461]), .A(V[461]), .E(fen));
Q_RELEASE_WEAK \genblk1[460].rrel ( .Q(L[460]), .E(ren));
Q_REGFORCE \genblk1[460].rfrc ( .Q(L[460]), .A(V[460]), .E(fen));
Q_RELEASE_WEAK \genblk1[459].rrel ( .Q(L[459]), .E(ren));
Q_REGFORCE \genblk1[459].rfrc ( .Q(L[459]), .A(V[459]), .E(fen));
Q_RELEASE_WEAK \genblk1[458].rrel ( .Q(L[458]), .E(ren));
Q_REGFORCE \genblk1[458].rfrc ( .Q(L[458]), .A(V[458]), .E(fen));
Q_RELEASE_WEAK \genblk1[457].rrel ( .Q(L[457]), .E(ren));
Q_REGFORCE \genblk1[457].rfrc ( .Q(L[457]), .A(V[457]), .E(fen));
Q_RELEASE_WEAK \genblk1[456].rrel ( .Q(L[456]), .E(ren));
Q_REGFORCE \genblk1[456].rfrc ( .Q(L[456]), .A(V[456]), .E(fen));
Q_RELEASE_WEAK \genblk1[455].rrel ( .Q(L[455]), .E(ren));
Q_REGFORCE \genblk1[455].rfrc ( .Q(L[455]), .A(V[455]), .E(fen));
Q_RELEASE_WEAK \genblk1[454].rrel ( .Q(L[454]), .E(ren));
Q_REGFORCE \genblk1[454].rfrc ( .Q(L[454]), .A(V[454]), .E(fen));
Q_RELEASE_WEAK \genblk1[453].rrel ( .Q(L[453]), .E(ren));
Q_REGFORCE \genblk1[453].rfrc ( .Q(L[453]), .A(V[453]), .E(fen));
Q_RELEASE_WEAK \genblk1[452].rrel ( .Q(L[452]), .E(ren));
Q_REGFORCE \genblk1[452].rfrc ( .Q(L[452]), .A(V[452]), .E(fen));
Q_RELEASE_WEAK \genblk1[451].rrel ( .Q(L[451]), .E(ren));
Q_REGFORCE \genblk1[451].rfrc ( .Q(L[451]), .A(V[451]), .E(fen));
Q_RELEASE_WEAK \genblk1[450].rrel ( .Q(L[450]), .E(ren));
Q_REGFORCE \genblk1[450].rfrc ( .Q(L[450]), .A(V[450]), .E(fen));
Q_RELEASE_WEAK \genblk1[449].rrel ( .Q(L[449]), .E(ren));
Q_REGFORCE \genblk1[449].rfrc ( .Q(L[449]), .A(V[449]), .E(fen));
Q_RELEASE_WEAK \genblk1[448].rrel ( .Q(L[448]), .E(ren));
Q_REGFORCE \genblk1[448].rfrc ( .Q(L[448]), .A(V[448]), .E(fen));
Q_RELEASE_WEAK \genblk1[447].rrel ( .Q(L[447]), .E(ren));
Q_REGFORCE \genblk1[447].rfrc ( .Q(L[447]), .A(V[447]), .E(fen));
Q_RELEASE_WEAK \genblk1[446].rrel ( .Q(L[446]), .E(ren));
Q_REGFORCE \genblk1[446].rfrc ( .Q(L[446]), .A(V[446]), .E(fen));
Q_RELEASE_WEAK \genblk1[445].rrel ( .Q(L[445]), .E(ren));
Q_REGFORCE \genblk1[445].rfrc ( .Q(L[445]), .A(V[445]), .E(fen));
Q_RELEASE_WEAK \genblk1[444].rrel ( .Q(L[444]), .E(ren));
Q_REGFORCE \genblk1[444].rfrc ( .Q(L[444]), .A(V[444]), .E(fen));
Q_RELEASE_WEAK \genblk1[443].rrel ( .Q(L[443]), .E(ren));
Q_REGFORCE \genblk1[443].rfrc ( .Q(L[443]), .A(V[443]), .E(fen));
Q_RELEASE_WEAK \genblk1[442].rrel ( .Q(L[442]), .E(ren));
Q_REGFORCE \genblk1[442].rfrc ( .Q(L[442]), .A(V[442]), .E(fen));
Q_RELEASE_WEAK \genblk1[441].rrel ( .Q(L[441]), .E(ren));
Q_REGFORCE \genblk1[441].rfrc ( .Q(L[441]), .A(V[441]), .E(fen));
Q_RELEASE_WEAK \genblk1[440].rrel ( .Q(L[440]), .E(ren));
Q_REGFORCE \genblk1[440].rfrc ( .Q(L[440]), .A(V[440]), .E(fen));
Q_RELEASE_WEAK \genblk1[439].rrel ( .Q(L[439]), .E(ren));
Q_REGFORCE \genblk1[439].rfrc ( .Q(L[439]), .A(V[439]), .E(fen));
Q_RELEASE_WEAK \genblk1[438].rrel ( .Q(L[438]), .E(ren));
Q_REGFORCE \genblk1[438].rfrc ( .Q(L[438]), .A(V[438]), .E(fen));
Q_RELEASE_WEAK \genblk1[437].rrel ( .Q(L[437]), .E(ren));
Q_REGFORCE \genblk1[437].rfrc ( .Q(L[437]), .A(V[437]), .E(fen));
Q_RELEASE_WEAK \genblk1[436].rrel ( .Q(L[436]), .E(ren));
Q_REGFORCE \genblk1[436].rfrc ( .Q(L[436]), .A(V[436]), .E(fen));
Q_RELEASE_WEAK \genblk1[435].rrel ( .Q(L[435]), .E(ren));
Q_REGFORCE \genblk1[435].rfrc ( .Q(L[435]), .A(V[435]), .E(fen));
Q_RELEASE_WEAK \genblk1[434].rrel ( .Q(L[434]), .E(ren));
Q_REGFORCE \genblk1[434].rfrc ( .Q(L[434]), .A(V[434]), .E(fen));
Q_RELEASE_WEAK \genblk1[433].rrel ( .Q(L[433]), .E(ren));
Q_REGFORCE \genblk1[433].rfrc ( .Q(L[433]), .A(V[433]), .E(fen));
Q_RELEASE_WEAK \genblk1[432].rrel ( .Q(L[432]), .E(ren));
Q_REGFORCE \genblk1[432].rfrc ( .Q(L[432]), .A(V[432]), .E(fen));
Q_RELEASE_WEAK \genblk1[431].rrel ( .Q(L[431]), .E(ren));
Q_REGFORCE \genblk1[431].rfrc ( .Q(L[431]), .A(V[431]), .E(fen));
Q_RELEASE_WEAK \genblk1[430].rrel ( .Q(L[430]), .E(ren));
Q_REGFORCE \genblk1[430].rfrc ( .Q(L[430]), .A(V[430]), .E(fen));
Q_RELEASE_WEAK \genblk1[429].rrel ( .Q(L[429]), .E(ren));
Q_REGFORCE \genblk1[429].rfrc ( .Q(L[429]), .A(V[429]), .E(fen));
Q_RELEASE_WEAK \genblk1[428].rrel ( .Q(L[428]), .E(ren));
Q_REGFORCE \genblk1[428].rfrc ( .Q(L[428]), .A(V[428]), .E(fen));
Q_RELEASE_WEAK \genblk1[427].rrel ( .Q(L[427]), .E(ren));
Q_REGFORCE \genblk1[427].rfrc ( .Q(L[427]), .A(V[427]), .E(fen));
Q_RELEASE_WEAK \genblk1[426].rrel ( .Q(L[426]), .E(ren));
Q_REGFORCE \genblk1[426].rfrc ( .Q(L[426]), .A(V[426]), .E(fen));
Q_RELEASE_WEAK \genblk1[425].rrel ( .Q(L[425]), .E(ren));
Q_REGFORCE \genblk1[425].rfrc ( .Q(L[425]), .A(V[425]), .E(fen));
Q_RELEASE_WEAK \genblk1[424].rrel ( .Q(L[424]), .E(ren));
Q_REGFORCE \genblk1[424].rfrc ( .Q(L[424]), .A(V[424]), .E(fen));
Q_RELEASE_WEAK \genblk1[423].rrel ( .Q(L[423]), .E(ren));
Q_REGFORCE \genblk1[423].rfrc ( .Q(L[423]), .A(V[423]), .E(fen));
Q_RELEASE_WEAK \genblk1[422].rrel ( .Q(L[422]), .E(ren));
Q_REGFORCE \genblk1[422].rfrc ( .Q(L[422]), .A(V[422]), .E(fen));
Q_RELEASE_WEAK \genblk1[421].rrel ( .Q(L[421]), .E(ren));
Q_REGFORCE \genblk1[421].rfrc ( .Q(L[421]), .A(V[421]), .E(fen));
Q_RELEASE_WEAK \genblk1[420].rrel ( .Q(L[420]), .E(ren));
Q_REGFORCE \genblk1[420].rfrc ( .Q(L[420]), .A(V[420]), .E(fen));
Q_RELEASE_WEAK \genblk1[419].rrel ( .Q(L[419]), .E(ren));
Q_REGFORCE \genblk1[419].rfrc ( .Q(L[419]), .A(V[419]), .E(fen));
Q_RELEASE_WEAK \genblk1[418].rrel ( .Q(L[418]), .E(ren));
Q_REGFORCE \genblk1[418].rfrc ( .Q(L[418]), .A(V[418]), .E(fen));
Q_RELEASE_WEAK \genblk1[417].rrel ( .Q(L[417]), .E(ren));
Q_REGFORCE \genblk1[417].rfrc ( .Q(L[417]), .A(V[417]), .E(fen));
Q_RELEASE_WEAK \genblk1[416].rrel ( .Q(L[416]), .E(ren));
Q_REGFORCE \genblk1[416].rfrc ( .Q(L[416]), .A(V[416]), .E(fen));
Q_RELEASE_WEAK \genblk1[415].rrel ( .Q(L[415]), .E(ren));
Q_REGFORCE \genblk1[415].rfrc ( .Q(L[415]), .A(V[415]), .E(fen));
Q_RELEASE_WEAK \genblk1[414].rrel ( .Q(L[414]), .E(ren));
Q_REGFORCE \genblk1[414].rfrc ( .Q(L[414]), .A(V[414]), .E(fen));
Q_RELEASE_WEAK \genblk1[413].rrel ( .Q(L[413]), .E(ren));
Q_REGFORCE \genblk1[413].rfrc ( .Q(L[413]), .A(V[413]), .E(fen));
Q_RELEASE_WEAK \genblk1[412].rrel ( .Q(L[412]), .E(ren));
Q_REGFORCE \genblk1[412].rfrc ( .Q(L[412]), .A(V[412]), .E(fen));
Q_RELEASE_WEAK \genblk1[411].rrel ( .Q(L[411]), .E(ren));
Q_REGFORCE \genblk1[411].rfrc ( .Q(L[411]), .A(V[411]), .E(fen));
Q_RELEASE_WEAK \genblk1[410].rrel ( .Q(L[410]), .E(ren));
Q_REGFORCE \genblk1[410].rfrc ( .Q(L[410]), .A(V[410]), .E(fen));
Q_RELEASE_WEAK \genblk1[409].rrel ( .Q(L[409]), .E(ren));
Q_REGFORCE \genblk1[409].rfrc ( .Q(L[409]), .A(V[409]), .E(fen));
Q_RELEASE_WEAK \genblk1[408].rrel ( .Q(L[408]), .E(ren));
Q_REGFORCE \genblk1[408].rfrc ( .Q(L[408]), .A(V[408]), .E(fen));
Q_RELEASE_WEAK \genblk1[407].rrel ( .Q(L[407]), .E(ren));
Q_REGFORCE \genblk1[407].rfrc ( .Q(L[407]), .A(V[407]), .E(fen));
Q_RELEASE_WEAK \genblk1[406].rrel ( .Q(L[406]), .E(ren));
Q_REGFORCE \genblk1[406].rfrc ( .Q(L[406]), .A(V[406]), .E(fen));
Q_RELEASE_WEAK \genblk1[405].rrel ( .Q(L[405]), .E(ren));
Q_REGFORCE \genblk1[405].rfrc ( .Q(L[405]), .A(V[405]), .E(fen));
Q_RELEASE_WEAK \genblk1[404].rrel ( .Q(L[404]), .E(ren));
Q_REGFORCE \genblk1[404].rfrc ( .Q(L[404]), .A(V[404]), .E(fen));
Q_RELEASE_WEAK \genblk1[403].rrel ( .Q(L[403]), .E(ren));
Q_REGFORCE \genblk1[403].rfrc ( .Q(L[403]), .A(V[403]), .E(fen));
Q_RELEASE_WEAK \genblk1[402].rrel ( .Q(L[402]), .E(ren));
Q_REGFORCE \genblk1[402].rfrc ( .Q(L[402]), .A(V[402]), .E(fen));
Q_RELEASE_WEAK \genblk1[401].rrel ( .Q(L[401]), .E(ren));
Q_REGFORCE \genblk1[401].rfrc ( .Q(L[401]), .A(V[401]), .E(fen));
Q_RELEASE_WEAK \genblk1[400].rrel ( .Q(L[400]), .E(ren));
Q_REGFORCE \genblk1[400].rfrc ( .Q(L[400]), .A(V[400]), .E(fen));
Q_RELEASE_WEAK \genblk1[399].rrel ( .Q(L[399]), .E(ren));
Q_REGFORCE \genblk1[399].rfrc ( .Q(L[399]), .A(V[399]), .E(fen));
Q_RELEASE_WEAK \genblk1[398].rrel ( .Q(L[398]), .E(ren));
Q_REGFORCE \genblk1[398].rfrc ( .Q(L[398]), .A(V[398]), .E(fen));
Q_RELEASE_WEAK \genblk1[397].rrel ( .Q(L[397]), .E(ren));
Q_REGFORCE \genblk1[397].rfrc ( .Q(L[397]), .A(V[397]), .E(fen));
Q_RELEASE_WEAK \genblk1[396].rrel ( .Q(L[396]), .E(ren));
Q_REGFORCE \genblk1[396].rfrc ( .Q(L[396]), .A(V[396]), .E(fen));
Q_RELEASE_WEAK \genblk1[395].rrel ( .Q(L[395]), .E(ren));
Q_REGFORCE \genblk1[395].rfrc ( .Q(L[395]), .A(V[395]), .E(fen));
Q_RELEASE_WEAK \genblk1[394].rrel ( .Q(L[394]), .E(ren));
Q_REGFORCE \genblk1[394].rfrc ( .Q(L[394]), .A(V[394]), .E(fen));
Q_RELEASE_WEAK \genblk1[393].rrel ( .Q(L[393]), .E(ren));
Q_REGFORCE \genblk1[393].rfrc ( .Q(L[393]), .A(V[393]), .E(fen));
Q_RELEASE_WEAK \genblk1[392].rrel ( .Q(L[392]), .E(ren));
Q_REGFORCE \genblk1[392].rfrc ( .Q(L[392]), .A(V[392]), .E(fen));
Q_RELEASE_WEAK \genblk1[391].rrel ( .Q(L[391]), .E(ren));
Q_REGFORCE \genblk1[391].rfrc ( .Q(L[391]), .A(V[391]), .E(fen));
Q_RELEASE_WEAK \genblk1[390].rrel ( .Q(L[390]), .E(ren));
Q_REGFORCE \genblk1[390].rfrc ( .Q(L[390]), .A(V[390]), .E(fen));
Q_RELEASE_WEAK \genblk1[389].rrel ( .Q(L[389]), .E(ren));
Q_REGFORCE \genblk1[389].rfrc ( .Q(L[389]), .A(V[389]), .E(fen));
Q_RELEASE_WEAK \genblk1[388].rrel ( .Q(L[388]), .E(ren));
Q_REGFORCE \genblk1[388].rfrc ( .Q(L[388]), .A(V[388]), .E(fen));
Q_RELEASE_WEAK \genblk1[387].rrel ( .Q(L[387]), .E(ren));
Q_REGFORCE \genblk1[387].rfrc ( .Q(L[387]), .A(V[387]), .E(fen));
Q_RELEASE_WEAK \genblk1[386].rrel ( .Q(L[386]), .E(ren));
Q_REGFORCE \genblk1[386].rfrc ( .Q(L[386]), .A(V[386]), .E(fen));
Q_RELEASE_WEAK \genblk1[385].rrel ( .Q(L[385]), .E(ren));
Q_REGFORCE \genblk1[385].rfrc ( .Q(L[385]), .A(V[385]), .E(fen));
Q_RELEASE_WEAK \genblk1[384].rrel ( .Q(L[384]), .E(ren));
Q_REGFORCE \genblk1[384].rfrc ( .Q(L[384]), .A(V[384]), .E(fen));
Q_RELEASE_WEAK \genblk1[383].rrel ( .Q(L[383]), .E(ren));
Q_REGFORCE \genblk1[383].rfrc ( .Q(L[383]), .A(V[383]), .E(fen));
Q_RELEASE_WEAK \genblk1[382].rrel ( .Q(L[382]), .E(ren));
Q_REGFORCE \genblk1[382].rfrc ( .Q(L[382]), .A(V[382]), .E(fen));
Q_RELEASE_WEAK \genblk1[381].rrel ( .Q(L[381]), .E(ren));
Q_REGFORCE \genblk1[381].rfrc ( .Q(L[381]), .A(V[381]), .E(fen));
Q_RELEASE_WEAK \genblk1[380].rrel ( .Q(L[380]), .E(ren));
Q_REGFORCE \genblk1[380].rfrc ( .Q(L[380]), .A(V[380]), .E(fen));
Q_RELEASE_WEAK \genblk1[379].rrel ( .Q(L[379]), .E(ren));
Q_REGFORCE \genblk1[379].rfrc ( .Q(L[379]), .A(V[379]), .E(fen));
Q_RELEASE_WEAK \genblk1[378].rrel ( .Q(L[378]), .E(ren));
Q_REGFORCE \genblk1[378].rfrc ( .Q(L[378]), .A(V[378]), .E(fen));
Q_RELEASE_WEAK \genblk1[377].rrel ( .Q(L[377]), .E(ren));
Q_REGFORCE \genblk1[377].rfrc ( .Q(L[377]), .A(V[377]), .E(fen));
Q_RELEASE_WEAK \genblk1[376].rrel ( .Q(L[376]), .E(ren));
Q_REGFORCE \genblk1[376].rfrc ( .Q(L[376]), .A(V[376]), .E(fen));
Q_RELEASE_WEAK \genblk1[375].rrel ( .Q(L[375]), .E(ren));
Q_REGFORCE \genblk1[375].rfrc ( .Q(L[375]), .A(V[375]), .E(fen));
Q_RELEASE_WEAK \genblk1[374].rrel ( .Q(L[374]), .E(ren));
Q_REGFORCE \genblk1[374].rfrc ( .Q(L[374]), .A(V[374]), .E(fen));
Q_RELEASE_WEAK \genblk1[373].rrel ( .Q(L[373]), .E(ren));
Q_REGFORCE \genblk1[373].rfrc ( .Q(L[373]), .A(V[373]), .E(fen));
Q_RELEASE_WEAK \genblk1[372].rrel ( .Q(L[372]), .E(ren));
Q_REGFORCE \genblk1[372].rfrc ( .Q(L[372]), .A(V[372]), .E(fen));
Q_RELEASE_WEAK \genblk1[371].rrel ( .Q(L[371]), .E(ren));
Q_REGFORCE \genblk1[371].rfrc ( .Q(L[371]), .A(V[371]), .E(fen));
Q_RELEASE_WEAK \genblk1[370].rrel ( .Q(L[370]), .E(ren));
Q_REGFORCE \genblk1[370].rfrc ( .Q(L[370]), .A(V[370]), .E(fen));
Q_RELEASE_WEAK \genblk1[369].rrel ( .Q(L[369]), .E(ren));
Q_REGFORCE \genblk1[369].rfrc ( .Q(L[369]), .A(V[369]), .E(fen));
Q_RELEASE_WEAK \genblk1[368].rrel ( .Q(L[368]), .E(ren));
Q_REGFORCE \genblk1[368].rfrc ( .Q(L[368]), .A(V[368]), .E(fen));
Q_RELEASE_WEAK \genblk1[367].rrel ( .Q(L[367]), .E(ren));
Q_REGFORCE \genblk1[367].rfrc ( .Q(L[367]), .A(V[367]), .E(fen));
Q_RELEASE_WEAK \genblk1[366].rrel ( .Q(L[366]), .E(ren));
Q_REGFORCE \genblk1[366].rfrc ( .Q(L[366]), .A(V[366]), .E(fen));
Q_RELEASE_WEAK \genblk1[365].rrel ( .Q(L[365]), .E(ren));
Q_REGFORCE \genblk1[365].rfrc ( .Q(L[365]), .A(V[365]), .E(fen));
Q_RELEASE_WEAK \genblk1[364].rrel ( .Q(L[364]), .E(ren));
Q_REGFORCE \genblk1[364].rfrc ( .Q(L[364]), .A(V[364]), .E(fen));
Q_RELEASE_WEAK \genblk1[363].rrel ( .Q(L[363]), .E(ren));
Q_REGFORCE \genblk1[363].rfrc ( .Q(L[363]), .A(V[363]), .E(fen));
Q_RELEASE_WEAK \genblk1[362].rrel ( .Q(L[362]), .E(ren));
Q_REGFORCE \genblk1[362].rfrc ( .Q(L[362]), .A(V[362]), .E(fen));
Q_RELEASE_WEAK \genblk1[361].rrel ( .Q(L[361]), .E(ren));
Q_REGFORCE \genblk1[361].rfrc ( .Q(L[361]), .A(V[361]), .E(fen));
Q_RELEASE_WEAK \genblk1[360].rrel ( .Q(L[360]), .E(ren));
Q_REGFORCE \genblk1[360].rfrc ( .Q(L[360]), .A(V[360]), .E(fen));
Q_RELEASE_WEAK \genblk1[359].rrel ( .Q(L[359]), .E(ren));
Q_REGFORCE \genblk1[359].rfrc ( .Q(L[359]), .A(V[359]), .E(fen));
Q_RELEASE_WEAK \genblk1[358].rrel ( .Q(L[358]), .E(ren));
Q_REGFORCE \genblk1[358].rfrc ( .Q(L[358]), .A(V[358]), .E(fen));
Q_RELEASE_WEAK \genblk1[357].rrel ( .Q(L[357]), .E(ren));
Q_REGFORCE \genblk1[357].rfrc ( .Q(L[357]), .A(V[357]), .E(fen));
Q_RELEASE_WEAK \genblk1[356].rrel ( .Q(L[356]), .E(ren));
Q_REGFORCE \genblk1[356].rfrc ( .Q(L[356]), .A(V[356]), .E(fen));
Q_RELEASE_WEAK \genblk1[355].rrel ( .Q(L[355]), .E(ren));
Q_REGFORCE \genblk1[355].rfrc ( .Q(L[355]), .A(V[355]), .E(fen));
Q_RELEASE_WEAK \genblk1[354].rrel ( .Q(L[354]), .E(ren));
Q_REGFORCE \genblk1[354].rfrc ( .Q(L[354]), .A(V[354]), .E(fen));
Q_RELEASE_WEAK \genblk1[353].rrel ( .Q(L[353]), .E(ren));
Q_REGFORCE \genblk1[353].rfrc ( .Q(L[353]), .A(V[353]), .E(fen));
Q_RELEASE_WEAK \genblk1[352].rrel ( .Q(L[352]), .E(ren));
Q_REGFORCE \genblk1[352].rfrc ( .Q(L[352]), .A(V[352]), .E(fen));
Q_RELEASE_WEAK \genblk1[351].rrel ( .Q(L[351]), .E(ren));
Q_REGFORCE \genblk1[351].rfrc ( .Q(L[351]), .A(V[351]), .E(fen));
Q_RELEASE_WEAK \genblk1[350].rrel ( .Q(L[350]), .E(ren));
Q_REGFORCE \genblk1[350].rfrc ( .Q(L[350]), .A(V[350]), .E(fen));
Q_RELEASE_WEAK \genblk1[349].rrel ( .Q(L[349]), .E(ren));
Q_REGFORCE \genblk1[349].rfrc ( .Q(L[349]), .A(V[349]), .E(fen));
Q_RELEASE_WEAK \genblk1[348].rrel ( .Q(L[348]), .E(ren));
Q_REGFORCE \genblk1[348].rfrc ( .Q(L[348]), .A(V[348]), .E(fen));
Q_RELEASE_WEAK \genblk1[347].rrel ( .Q(L[347]), .E(ren));
Q_REGFORCE \genblk1[347].rfrc ( .Q(L[347]), .A(V[347]), .E(fen));
Q_RELEASE_WEAK \genblk1[346].rrel ( .Q(L[346]), .E(ren));
Q_REGFORCE \genblk1[346].rfrc ( .Q(L[346]), .A(V[346]), .E(fen));
Q_RELEASE_WEAK \genblk1[345].rrel ( .Q(L[345]), .E(ren));
Q_REGFORCE \genblk1[345].rfrc ( .Q(L[345]), .A(V[345]), .E(fen));
Q_RELEASE_WEAK \genblk1[344].rrel ( .Q(L[344]), .E(ren));
Q_REGFORCE \genblk1[344].rfrc ( .Q(L[344]), .A(V[344]), .E(fen));
Q_RELEASE_WEAK \genblk1[343].rrel ( .Q(L[343]), .E(ren));
Q_REGFORCE \genblk1[343].rfrc ( .Q(L[343]), .A(V[343]), .E(fen));
Q_RELEASE_WEAK \genblk1[342].rrel ( .Q(L[342]), .E(ren));
Q_REGFORCE \genblk1[342].rfrc ( .Q(L[342]), .A(V[342]), .E(fen));
Q_RELEASE_WEAK \genblk1[341].rrel ( .Q(L[341]), .E(ren));
Q_REGFORCE \genblk1[341].rfrc ( .Q(L[341]), .A(V[341]), .E(fen));
Q_RELEASE_WEAK \genblk1[340].rrel ( .Q(L[340]), .E(ren));
Q_REGFORCE \genblk1[340].rfrc ( .Q(L[340]), .A(V[340]), .E(fen));
Q_RELEASE_WEAK \genblk1[339].rrel ( .Q(L[339]), .E(ren));
Q_REGFORCE \genblk1[339].rfrc ( .Q(L[339]), .A(V[339]), .E(fen));
Q_RELEASE_WEAK \genblk1[338].rrel ( .Q(L[338]), .E(ren));
Q_REGFORCE \genblk1[338].rfrc ( .Q(L[338]), .A(V[338]), .E(fen));
Q_RELEASE_WEAK \genblk1[337].rrel ( .Q(L[337]), .E(ren));
Q_REGFORCE \genblk1[337].rfrc ( .Q(L[337]), .A(V[337]), .E(fen));
Q_RELEASE_WEAK \genblk1[336].rrel ( .Q(L[336]), .E(ren));
Q_REGFORCE \genblk1[336].rfrc ( .Q(L[336]), .A(V[336]), .E(fen));
Q_RELEASE_WEAK \genblk1[335].rrel ( .Q(L[335]), .E(ren));
Q_REGFORCE \genblk1[335].rfrc ( .Q(L[335]), .A(V[335]), .E(fen));
Q_RELEASE_WEAK \genblk1[334].rrel ( .Q(L[334]), .E(ren));
Q_REGFORCE \genblk1[334].rfrc ( .Q(L[334]), .A(V[334]), .E(fen));
Q_RELEASE_WEAK \genblk1[333].rrel ( .Q(L[333]), .E(ren));
Q_REGFORCE \genblk1[333].rfrc ( .Q(L[333]), .A(V[333]), .E(fen));
Q_RELEASE_WEAK \genblk1[332].rrel ( .Q(L[332]), .E(ren));
Q_REGFORCE \genblk1[332].rfrc ( .Q(L[332]), .A(V[332]), .E(fen));
Q_RELEASE_WEAK \genblk1[331].rrel ( .Q(L[331]), .E(ren));
Q_REGFORCE \genblk1[331].rfrc ( .Q(L[331]), .A(V[331]), .E(fen));
Q_RELEASE_WEAK \genblk1[330].rrel ( .Q(L[330]), .E(ren));
Q_REGFORCE \genblk1[330].rfrc ( .Q(L[330]), .A(V[330]), .E(fen));
Q_RELEASE_WEAK \genblk1[329].rrel ( .Q(L[329]), .E(ren));
Q_REGFORCE \genblk1[329].rfrc ( .Q(L[329]), .A(V[329]), .E(fen));
Q_RELEASE_WEAK \genblk1[328].rrel ( .Q(L[328]), .E(ren));
Q_REGFORCE \genblk1[328].rfrc ( .Q(L[328]), .A(V[328]), .E(fen));
Q_RELEASE_WEAK \genblk1[327].rrel ( .Q(L[327]), .E(ren));
Q_REGFORCE \genblk1[327].rfrc ( .Q(L[327]), .A(V[327]), .E(fen));
Q_RELEASE_WEAK \genblk1[326].rrel ( .Q(L[326]), .E(ren));
Q_REGFORCE \genblk1[326].rfrc ( .Q(L[326]), .A(V[326]), .E(fen));
Q_RELEASE_WEAK \genblk1[325].rrel ( .Q(L[325]), .E(ren));
Q_REGFORCE \genblk1[325].rfrc ( .Q(L[325]), .A(V[325]), .E(fen));
Q_RELEASE_WEAK \genblk1[324].rrel ( .Q(L[324]), .E(ren));
Q_REGFORCE \genblk1[324].rfrc ( .Q(L[324]), .A(V[324]), .E(fen));
Q_RELEASE_WEAK \genblk1[323].rrel ( .Q(L[323]), .E(ren));
Q_REGFORCE \genblk1[323].rfrc ( .Q(L[323]), .A(V[323]), .E(fen));
Q_RELEASE_WEAK \genblk1[322].rrel ( .Q(L[322]), .E(ren));
Q_REGFORCE \genblk1[322].rfrc ( .Q(L[322]), .A(V[322]), .E(fen));
Q_RELEASE_WEAK \genblk1[321].rrel ( .Q(L[321]), .E(ren));
Q_REGFORCE \genblk1[321].rfrc ( .Q(L[321]), .A(V[321]), .E(fen));
Q_RELEASE_WEAK \genblk1[320].rrel ( .Q(L[320]), .E(ren));
Q_REGFORCE \genblk1[320].rfrc ( .Q(L[320]), .A(V[320]), .E(fen));
Q_RELEASE_WEAK \genblk1[319].rrel ( .Q(L[319]), .E(ren));
Q_REGFORCE \genblk1[319].rfrc ( .Q(L[319]), .A(V[319]), .E(fen));
Q_RELEASE_WEAK \genblk1[318].rrel ( .Q(L[318]), .E(ren));
Q_REGFORCE \genblk1[318].rfrc ( .Q(L[318]), .A(V[318]), .E(fen));
Q_RELEASE_WEAK \genblk1[317].rrel ( .Q(L[317]), .E(ren));
Q_REGFORCE \genblk1[317].rfrc ( .Q(L[317]), .A(V[317]), .E(fen));
Q_RELEASE_WEAK \genblk1[316].rrel ( .Q(L[316]), .E(ren));
Q_REGFORCE \genblk1[316].rfrc ( .Q(L[316]), .A(V[316]), .E(fen));
Q_RELEASE_WEAK \genblk1[315].rrel ( .Q(L[315]), .E(ren));
Q_REGFORCE \genblk1[315].rfrc ( .Q(L[315]), .A(V[315]), .E(fen));
Q_RELEASE_WEAK \genblk1[314].rrel ( .Q(L[314]), .E(ren));
Q_REGFORCE \genblk1[314].rfrc ( .Q(L[314]), .A(V[314]), .E(fen));
Q_RELEASE_WEAK \genblk1[313].rrel ( .Q(L[313]), .E(ren));
Q_REGFORCE \genblk1[313].rfrc ( .Q(L[313]), .A(V[313]), .E(fen));
Q_RELEASE_WEAK \genblk1[312].rrel ( .Q(L[312]), .E(ren));
Q_REGFORCE \genblk1[312].rfrc ( .Q(L[312]), .A(V[312]), .E(fen));
Q_RELEASE_WEAK \genblk1[311].rrel ( .Q(L[311]), .E(ren));
Q_REGFORCE \genblk1[311].rfrc ( .Q(L[311]), .A(V[311]), .E(fen));
Q_RELEASE_WEAK \genblk1[310].rrel ( .Q(L[310]), .E(ren));
Q_REGFORCE \genblk1[310].rfrc ( .Q(L[310]), .A(V[310]), .E(fen));
Q_RELEASE_WEAK \genblk1[309].rrel ( .Q(L[309]), .E(ren));
Q_REGFORCE \genblk1[309].rfrc ( .Q(L[309]), .A(V[309]), .E(fen));
Q_RELEASE_WEAK \genblk1[308].rrel ( .Q(L[308]), .E(ren));
Q_REGFORCE \genblk1[308].rfrc ( .Q(L[308]), .A(V[308]), .E(fen));
Q_RELEASE_WEAK \genblk1[307].rrel ( .Q(L[307]), .E(ren));
Q_REGFORCE \genblk1[307].rfrc ( .Q(L[307]), .A(V[307]), .E(fen));
Q_RELEASE_WEAK \genblk1[306].rrel ( .Q(L[306]), .E(ren));
Q_REGFORCE \genblk1[306].rfrc ( .Q(L[306]), .A(V[306]), .E(fen));
Q_RELEASE_WEAK \genblk1[305].rrel ( .Q(L[305]), .E(ren));
Q_REGFORCE \genblk1[305].rfrc ( .Q(L[305]), .A(V[305]), .E(fen));
Q_RELEASE_WEAK \genblk1[304].rrel ( .Q(L[304]), .E(ren));
Q_REGFORCE \genblk1[304].rfrc ( .Q(L[304]), .A(V[304]), .E(fen));
Q_RELEASE_WEAK \genblk1[303].rrel ( .Q(L[303]), .E(ren));
Q_REGFORCE \genblk1[303].rfrc ( .Q(L[303]), .A(V[303]), .E(fen));
Q_RELEASE_WEAK \genblk1[302].rrel ( .Q(L[302]), .E(ren));
Q_REGFORCE \genblk1[302].rfrc ( .Q(L[302]), .A(V[302]), .E(fen));
Q_RELEASE_WEAK \genblk1[301].rrel ( .Q(L[301]), .E(ren));
Q_REGFORCE \genblk1[301].rfrc ( .Q(L[301]), .A(V[301]), .E(fen));
Q_RELEASE_WEAK \genblk1[300].rrel ( .Q(L[300]), .E(ren));
Q_REGFORCE \genblk1[300].rfrc ( .Q(L[300]), .A(V[300]), .E(fen));
Q_RELEASE_WEAK \genblk1[299].rrel ( .Q(L[299]), .E(ren));
Q_REGFORCE \genblk1[299].rfrc ( .Q(L[299]), .A(V[299]), .E(fen));
Q_RELEASE_WEAK \genblk1[298].rrel ( .Q(L[298]), .E(ren));
Q_REGFORCE \genblk1[298].rfrc ( .Q(L[298]), .A(V[298]), .E(fen));
Q_RELEASE_WEAK \genblk1[297].rrel ( .Q(L[297]), .E(ren));
Q_REGFORCE \genblk1[297].rfrc ( .Q(L[297]), .A(V[297]), .E(fen));
Q_RELEASE_WEAK \genblk1[296].rrel ( .Q(L[296]), .E(ren));
Q_REGFORCE \genblk1[296].rfrc ( .Q(L[296]), .A(V[296]), .E(fen));
Q_RELEASE_WEAK \genblk1[295].rrel ( .Q(L[295]), .E(ren));
Q_REGFORCE \genblk1[295].rfrc ( .Q(L[295]), .A(V[295]), .E(fen));
Q_RELEASE_WEAK \genblk1[294].rrel ( .Q(L[294]), .E(ren));
Q_REGFORCE \genblk1[294].rfrc ( .Q(L[294]), .A(V[294]), .E(fen));
Q_RELEASE_WEAK \genblk1[293].rrel ( .Q(L[293]), .E(ren));
Q_REGFORCE \genblk1[293].rfrc ( .Q(L[293]), .A(V[293]), .E(fen));
Q_RELEASE_WEAK \genblk1[292].rrel ( .Q(L[292]), .E(ren));
Q_REGFORCE \genblk1[292].rfrc ( .Q(L[292]), .A(V[292]), .E(fen));
Q_RELEASE_WEAK \genblk1[291].rrel ( .Q(L[291]), .E(ren));
Q_REGFORCE \genblk1[291].rfrc ( .Q(L[291]), .A(V[291]), .E(fen));
Q_RELEASE_WEAK \genblk1[290].rrel ( .Q(L[290]), .E(ren));
Q_REGFORCE \genblk1[290].rfrc ( .Q(L[290]), .A(V[290]), .E(fen));
Q_RELEASE_WEAK \genblk1[289].rrel ( .Q(L[289]), .E(ren));
Q_REGFORCE \genblk1[289].rfrc ( .Q(L[289]), .A(V[289]), .E(fen));
Q_RELEASE_WEAK \genblk1[288].rrel ( .Q(L[288]), .E(ren));
Q_REGFORCE \genblk1[288].rfrc ( .Q(L[288]), .A(V[288]), .E(fen));
Q_RELEASE_WEAK \genblk1[287].rrel ( .Q(L[287]), .E(ren));
Q_REGFORCE \genblk1[287].rfrc ( .Q(L[287]), .A(V[287]), .E(fen));
Q_RELEASE_WEAK \genblk1[286].rrel ( .Q(L[286]), .E(ren));
Q_REGFORCE \genblk1[286].rfrc ( .Q(L[286]), .A(V[286]), .E(fen));
Q_RELEASE_WEAK \genblk1[285].rrel ( .Q(L[285]), .E(ren));
Q_REGFORCE \genblk1[285].rfrc ( .Q(L[285]), .A(V[285]), .E(fen));
Q_RELEASE_WEAK \genblk1[284].rrel ( .Q(L[284]), .E(ren));
Q_REGFORCE \genblk1[284].rfrc ( .Q(L[284]), .A(V[284]), .E(fen));
Q_RELEASE_WEAK \genblk1[283].rrel ( .Q(L[283]), .E(ren));
Q_REGFORCE \genblk1[283].rfrc ( .Q(L[283]), .A(V[283]), .E(fen));
Q_RELEASE_WEAK \genblk1[282].rrel ( .Q(L[282]), .E(ren));
Q_REGFORCE \genblk1[282].rfrc ( .Q(L[282]), .A(V[282]), .E(fen));
Q_RELEASE_WEAK \genblk1[281].rrel ( .Q(L[281]), .E(ren));
Q_REGFORCE \genblk1[281].rfrc ( .Q(L[281]), .A(V[281]), .E(fen));
Q_RELEASE_WEAK \genblk1[280].rrel ( .Q(L[280]), .E(ren));
Q_REGFORCE \genblk1[280].rfrc ( .Q(L[280]), .A(V[280]), .E(fen));
Q_RELEASE_WEAK \genblk1[279].rrel ( .Q(L[279]), .E(ren));
Q_REGFORCE \genblk1[279].rfrc ( .Q(L[279]), .A(V[279]), .E(fen));
Q_RELEASE_WEAK \genblk1[278].rrel ( .Q(L[278]), .E(ren));
Q_REGFORCE \genblk1[278].rfrc ( .Q(L[278]), .A(V[278]), .E(fen));
Q_RELEASE_WEAK \genblk1[277].rrel ( .Q(L[277]), .E(ren));
Q_REGFORCE \genblk1[277].rfrc ( .Q(L[277]), .A(V[277]), .E(fen));
Q_RELEASE_WEAK \genblk1[276].rrel ( .Q(L[276]), .E(ren));
Q_REGFORCE \genblk1[276].rfrc ( .Q(L[276]), .A(V[276]), .E(fen));
Q_RELEASE_WEAK \genblk1[275].rrel ( .Q(L[275]), .E(ren));
Q_REGFORCE \genblk1[275].rfrc ( .Q(L[275]), .A(V[275]), .E(fen));
Q_RELEASE_WEAK \genblk1[274].rrel ( .Q(L[274]), .E(ren));
Q_REGFORCE \genblk1[274].rfrc ( .Q(L[274]), .A(V[274]), .E(fen));
Q_RELEASE_WEAK \genblk1[273].rrel ( .Q(L[273]), .E(ren));
Q_REGFORCE \genblk1[273].rfrc ( .Q(L[273]), .A(V[273]), .E(fen));
Q_RELEASE_WEAK \genblk1[272].rrel ( .Q(L[272]), .E(ren));
Q_REGFORCE \genblk1[272].rfrc ( .Q(L[272]), .A(V[272]), .E(fen));
Q_RELEASE_WEAK \genblk1[271].rrel ( .Q(L[271]), .E(ren));
Q_REGFORCE \genblk1[271].rfrc ( .Q(L[271]), .A(V[271]), .E(fen));
Q_RELEASE_WEAK \genblk1[270].rrel ( .Q(L[270]), .E(ren));
Q_REGFORCE \genblk1[270].rfrc ( .Q(L[270]), .A(V[270]), .E(fen));
Q_RELEASE_WEAK \genblk1[269].rrel ( .Q(L[269]), .E(ren));
Q_REGFORCE \genblk1[269].rfrc ( .Q(L[269]), .A(V[269]), .E(fen));
Q_RELEASE_WEAK \genblk1[268].rrel ( .Q(L[268]), .E(ren));
Q_REGFORCE \genblk1[268].rfrc ( .Q(L[268]), .A(V[268]), .E(fen));
Q_RELEASE_WEAK \genblk1[267].rrel ( .Q(L[267]), .E(ren));
Q_REGFORCE \genblk1[267].rfrc ( .Q(L[267]), .A(V[267]), .E(fen));
Q_RELEASE_WEAK \genblk1[266].rrel ( .Q(L[266]), .E(ren));
Q_REGFORCE \genblk1[266].rfrc ( .Q(L[266]), .A(V[266]), .E(fen));
Q_RELEASE_WEAK \genblk1[265].rrel ( .Q(L[265]), .E(ren));
Q_REGFORCE \genblk1[265].rfrc ( .Q(L[265]), .A(V[265]), .E(fen));
Q_RELEASE_WEAK \genblk1[264].rrel ( .Q(L[264]), .E(ren));
Q_REGFORCE \genblk1[264].rfrc ( .Q(L[264]), .A(V[264]), .E(fen));
Q_RELEASE_WEAK \genblk1[263].rrel ( .Q(L[263]), .E(ren));
Q_REGFORCE \genblk1[263].rfrc ( .Q(L[263]), .A(V[263]), .E(fen));
Q_RELEASE_WEAK \genblk1[262].rrel ( .Q(L[262]), .E(ren));
Q_REGFORCE \genblk1[262].rfrc ( .Q(L[262]), .A(V[262]), .E(fen));
Q_RELEASE_WEAK \genblk1[261].rrel ( .Q(L[261]), .E(ren));
Q_REGFORCE \genblk1[261].rfrc ( .Q(L[261]), .A(V[261]), .E(fen));
Q_RELEASE_WEAK \genblk1[260].rrel ( .Q(L[260]), .E(ren));
Q_REGFORCE \genblk1[260].rfrc ( .Q(L[260]), .A(V[260]), .E(fen));
Q_RELEASE_WEAK \genblk1[259].rrel ( .Q(L[259]), .E(ren));
Q_REGFORCE \genblk1[259].rfrc ( .Q(L[259]), .A(V[259]), .E(fen));
Q_RELEASE_WEAK \genblk1[258].rrel ( .Q(L[258]), .E(ren));
Q_REGFORCE \genblk1[258].rfrc ( .Q(L[258]), .A(V[258]), .E(fen));
Q_RELEASE_WEAK \genblk1[257].rrel ( .Q(L[257]), .E(ren));
Q_REGFORCE \genblk1[257].rfrc ( .Q(L[257]), .A(V[257]), .E(fen));
Q_RELEASE_WEAK \genblk1[256].rrel ( .Q(L[256]), .E(ren));
Q_REGFORCE \genblk1[256].rfrc ( .Q(L[256]), .A(V[256]), .E(fen));
Q_RELEASE_WEAK \genblk1[255].rrel ( .Q(L[255]), .E(ren));
Q_REGFORCE \genblk1[255].rfrc ( .Q(L[255]), .A(V[255]), .E(fen));
Q_RELEASE_WEAK \genblk1[254].rrel ( .Q(L[254]), .E(ren));
Q_REGFORCE \genblk1[254].rfrc ( .Q(L[254]), .A(V[254]), .E(fen));
Q_RELEASE_WEAK \genblk1[253].rrel ( .Q(L[253]), .E(ren));
Q_REGFORCE \genblk1[253].rfrc ( .Q(L[253]), .A(V[253]), .E(fen));
Q_RELEASE_WEAK \genblk1[252].rrel ( .Q(L[252]), .E(ren));
Q_REGFORCE \genblk1[252].rfrc ( .Q(L[252]), .A(V[252]), .E(fen));
Q_RELEASE_WEAK \genblk1[251].rrel ( .Q(L[251]), .E(ren));
Q_REGFORCE \genblk1[251].rfrc ( .Q(L[251]), .A(V[251]), .E(fen));
Q_RELEASE_WEAK \genblk1[250].rrel ( .Q(L[250]), .E(ren));
Q_REGFORCE \genblk1[250].rfrc ( .Q(L[250]), .A(V[250]), .E(fen));
Q_RELEASE_WEAK \genblk1[249].rrel ( .Q(L[249]), .E(ren));
Q_REGFORCE \genblk1[249].rfrc ( .Q(L[249]), .A(V[249]), .E(fen));
Q_RELEASE_WEAK \genblk1[248].rrel ( .Q(L[248]), .E(ren));
Q_REGFORCE \genblk1[248].rfrc ( .Q(L[248]), .A(V[248]), .E(fen));
Q_RELEASE_WEAK \genblk1[247].rrel ( .Q(L[247]), .E(ren));
Q_REGFORCE \genblk1[247].rfrc ( .Q(L[247]), .A(V[247]), .E(fen));
Q_RELEASE_WEAK \genblk1[246].rrel ( .Q(L[246]), .E(ren));
Q_REGFORCE \genblk1[246].rfrc ( .Q(L[246]), .A(V[246]), .E(fen));
Q_RELEASE_WEAK \genblk1[245].rrel ( .Q(L[245]), .E(ren));
Q_REGFORCE \genblk1[245].rfrc ( .Q(L[245]), .A(V[245]), .E(fen));
Q_RELEASE_WEAK \genblk1[244].rrel ( .Q(L[244]), .E(ren));
Q_REGFORCE \genblk1[244].rfrc ( .Q(L[244]), .A(V[244]), .E(fen));
Q_RELEASE_WEAK \genblk1[243].rrel ( .Q(L[243]), .E(ren));
Q_REGFORCE \genblk1[243].rfrc ( .Q(L[243]), .A(V[243]), .E(fen));
Q_RELEASE_WEAK \genblk1[242].rrel ( .Q(L[242]), .E(ren));
Q_REGFORCE \genblk1[242].rfrc ( .Q(L[242]), .A(V[242]), .E(fen));
Q_RELEASE_WEAK \genblk1[241].rrel ( .Q(L[241]), .E(ren));
Q_REGFORCE \genblk1[241].rfrc ( .Q(L[241]), .A(V[241]), .E(fen));
Q_RELEASE_WEAK \genblk1[240].rrel ( .Q(L[240]), .E(ren));
Q_REGFORCE \genblk1[240].rfrc ( .Q(L[240]), .A(V[240]), .E(fen));
Q_RELEASE_WEAK \genblk1[239].rrel ( .Q(L[239]), .E(ren));
Q_REGFORCE \genblk1[239].rfrc ( .Q(L[239]), .A(V[239]), .E(fen));
Q_RELEASE_WEAK \genblk1[238].rrel ( .Q(L[238]), .E(ren));
Q_REGFORCE \genblk1[238].rfrc ( .Q(L[238]), .A(V[238]), .E(fen));
Q_RELEASE_WEAK \genblk1[237].rrel ( .Q(L[237]), .E(ren));
Q_REGFORCE \genblk1[237].rfrc ( .Q(L[237]), .A(V[237]), .E(fen));
Q_RELEASE_WEAK \genblk1[236].rrel ( .Q(L[236]), .E(ren));
Q_REGFORCE \genblk1[236].rfrc ( .Q(L[236]), .A(V[236]), .E(fen));
Q_RELEASE_WEAK \genblk1[235].rrel ( .Q(L[235]), .E(ren));
Q_REGFORCE \genblk1[235].rfrc ( .Q(L[235]), .A(V[235]), .E(fen));
Q_RELEASE_WEAK \genblk1[234].rrel ( .Q(L[234]), .E(ren));
Q_REGFORCE \genblk1[234].rfrc ( .Q(L[234]), .A(V[234]), .E(fen));
Q_RELEASE_WEAK \genblk1[233].rrel ( .Q(L[233]), .E(ren));
Q_REGFORCE \genblk1[233].rfrc ( .Q(L[233]), .A(V[233]), .E(fen));
Q_RELEASE_WEAK \genblk1[232].rrel ( .Q(L[232]), .E(ren));
Q_REGFORCE \genblk1[232].rfrc ( .Q(L[232]), .A(V[232]), .E(fen));
Q_RELEASE_WEAK \genblk1[231].rrel ( .Q(L[231]), .E(ren));
Q_REGFORCE \genblk1[231].rfrc ( .Q(L[231]), .A(V[231]), .E(fen));
Q_RELEASE_WEAK \genblk1[230].rrel ( .Q(L[230]), .E(ren));
Q_REGFORCE \genblk1[230].rfrc ( .Q(L[230]), .A(V[230]), .E(fen));
Q_RELEASE_WEAK \genblk1[229].rrel ( .Q(L[229]), .E(ren));
Q_REGFORCE \genblk1[229].rfrc ( .Q(L[229]), .A(V[229]), .E(fen));
Q_RELEASE_WEAK \genblk1[228].rrel ( .Q(L[228]), .E(ren));
Q_REGFORCE \genblk1[228].rfrc ( .Q(L[228]), .A(V[228]), .E(fen));
Q_RELEASE_WEAK \genblk1[227].rrel ( .Q(L[227]), .E(ren));
Q_REGFORCE \genblk1[227].rfrc ( .Q(L[227]), .A(V[227]), .E(fen));
Q_RELEASE_WEAK \genblk1[226].rrel ( .Q(L[226]), .E(ren));
Q_REGFORCE \genblk1[226].rfrc ( .Q(L[226]), .A(V[226]), .E(fen));
Q_RELEASE_WEAK \genblk1[225].rrel ( .Q(L[225]), .E(ren));
Q_REGFORCE \genblk1[225].rfrc ( .Q(L[225]), .A(V[225]), .E(fen));
Q_RELEASE_WEAK \genblk1[224].rrel ( .Q(L[224]), .E(ren));
Q_REGFORCE \genblk1[224].rfrc ( .Q(L[224]), .A(V[224]), .E(fen));
Q_RELEASE_WEAK \genblk1[223].rrel ( .Q(L[223]), .E(ren));
Q_REGFORCE \genblk1[223].rfrc ( .Q(L[223]), .A(V[223]), .E(fen));
Q_RELEASE_WEAK \genblk1[222].rrel ( .Q(L[222]), .E(ren));
Q_REGFORCE \genblk1[222].rfrc ( .Q(L[222]), .A(V[222]), .E(fen));
Q_RELEASE_WEAK \genblk1[221].rrel ( .Q(L[221]), .E(ren));
Q_REGFORCE \genblk1[221].rfrc ( .Q(L[221]), .A(V[221]), .E(fen));
Q_RELEASE_WEAK \genblk1[220].rrel ( .Q(L[220]), .E(ren));
Q_REGFORCE \genblk1[220].rfrc ( .Q(L[220]), .A(V[220]), .E(fen));
Q_RELEASE_WEAK \genblk1[219].rrel ( .Q(L[219]), .E(ren));
Q_REGFORCE \genblk1[219].rfrc ( .Q(L[219]), .A(V[219]), .E(fen));
Q_RELEASE_WEAK \genblk1[218].rrel ( .Q(L[218]), .E(ren));
Q_REGFORCE \genblk1[218].rfrc ( .Q(L[218]), .A(V[218]), .E(fen));
Q_RELEASE_WEAK \genblk1[217].rrel ( .Q(L[217]), .E(ren));
Q_REGFORCE \genblk1[217].rfrc ( .Q(L[217]), .A(V[217]), .E(fen));
Q_RELEASE_WEAK \genblk1[216].rrel ( .Q(L[216]), .E(ren));
Q_REGFORCE \genblk1[216].rfrc ( .Q(L[216]), .A(V[216]), .E(fen));
Q_RELEASE_WEAK \genblk1[215].rrel ( .Q(L[215]), .E(ren));
Q_REGFORCE \genblk1[215].rfrc ( .Q(L[215]), .A(V[215]), .E(fen));
Q_RELEASE_WEAK \genblk1[214].rrel ( .Q(L[214]), .E(ren));
Q_REGFORCE \genblk1[214].rfrc ( .Q(L[214]), .A(V[214]), .E(fen));
Q_RELEASE_WEAK \genblk1[213].rrel ( .Q(L[213]), .E(ren));
Q_REGFORCE \genblk1[213].rfrc ( .Q(L[213]), .A(V[213]), .E(fen));
Q_RELEASE_WEAK \genblk1[212].rrel ( .Q(L[212]), .E(ren));
Q_REGFORCE \genblk1[212].rfrc ( .Q(L[212]), .A(V[212]), .E(fen));
Q_RELEASE_WEAK \genblk1[211].rrel ( .Q(L[211]), .E(ren));
Q_REGFORCE \genblk1[211].rfrc ( .Q(L[211]), .A(V[211]), .E(fen));
Q_RELEASE_WEAK \genblk1[210].rrel ( .Q(L[210]), .E(ren));
Q_REGFORCE \genblk1[210].rfrc ( .Q(L[210]), .A(V[210]), .E(fen));
Q_RELEASE_WEAK \genblk1[209].rrel ( .Q(L[209]), .E(ren));
Q_REGFORCE \genblk1[209].rfrc ( .Q(L[209]), .A(V[209]), .E(fen));
Q_RELEASE_WEAK \genblk1[208].rrel ( .Q(L[208]), .E(ren));
Q_REGFORCE \genblk1[208].rfrc ( .Q(L[208]), .A(V[208]), .E(fen));
Q_RELEASE_WEAK \genblk1[207].rrel ( .Q(L[207]), .E(ren));
Q_REGFORCE \genblk1[207].rfrc ( .Q(L[207]), .A(V[207]), .E(fen));
Q_RELEASE_WEAK \genblk1[206].rrel ( .Q(L[206]), .E(ren));
Q_REGFORCE \genblk1[206].rfrc ( .Q(L[206]), .A(V[206]), .E(fen));
Q_RELEASE_WEAK \genblk1[205].rrel ( .Q(L[205]), .E(ren));
Q_REGFORCE \genblk1[205].rfrc ( .Q(L[205]), .A(V[205]), .E(fen));
Q_RELEASE_WEAK \genblk1[204].rrel ( .Q(L[204]), .E(ren));
Q_REGFORCE \genblk1[204].rfrc ( .Q(L[204]), .A(V[204]), .E(fen));
Q_RELEASE_WEAK \genblk1[203].rrel ( .Q(L[203]), .E(ren));
Q_REGFORCE \genblk1[203].rfrc ( .Q(L[203]), .A(V[203]), .E(fen));
Q_RELEASE_WEAK \genblk1[202].rrel ( .Q(L[202]), .E(ren));
Q_REGFORCE \genblk1[202].rfrc ( .Q(L[202]), .A(V[202]), .E(fen));
Q_RELEASE_WEAK \genblk1[201].rrel ( .Q(L[201]), .E(ren));
Q_REGFORCE \genblk1[201].rfrc ( .Q(L[201]), .A(V[201]), .E(fen));
Q_RELEASE_WEAK \genblk1[200].rrel ( .Q(L[200]), .E(ren));
Q_REGFORCE \genblk1[200].rfrc ( .Q(L[200]), .A(V[200]), .E(fen));
Q_RELEASE_WEAK \genblk1[199].rrel ( .Q(L[199]), .E(ren));
Q_REGFORCE \genblk1[199].rfrc ( .Q(L[199]), .A(V[199]), .E(fen));
Q_RELEASE_WEAK \genblk1[198].rrel ( .Q(L[198]), .E(ren));
Q_REGFORCE \genblk1[198].rfrc ( .Q(L[198]), .A(V[198]), .E(fen));
Q_RELEASE_WEAK \genblk1[197].rrel ( .Q(L[197]), .E(ren));
Q_REGFORCE \genblk1[197].rfrc ( .Q(L[197]), .A(V[197]), .E(fen));
Q_RELEASE_WEAK \genblk1[196].rrel ( .Q(L[196]), .E(ren));
Q_REGFORCE \genblk1[196].rfrc ( .Q(L[196]), .A(V[196]), .E(fen));
Q_RELEASE_WEAK \genblk1[195].rrel ( .Q(L[195]), .E(ren));
Q_REGFORCE \genblk1[195].rfrc ( .Q(L[195]), .A(V[195]), .E(fen));
Q_RELEASE_WEAK \genblk1[194].rrel ( .Q(L[194]), .E(ren));
Q_REGFORCE \genblk1[194].rfrc ( .Q(L[194]), .A(V[194]), .E(fen));
Q_RELEASE_WEAK \genblk1[193].rrel ( .Q(L[193]), .E(ren));
Q_REGFORCE \genblk1[193].rfrc ( .Q(L[193]), .A(V[193]), .E(fen));
Q_RELEASE_WEAK \genblk1[192].rrel ( .Q(L[192]), .E(ren));
Q_REGFORCE \genblk1[192].rfrc ( .Q(L[192]), .A(V[192]), .E(fen));
Q_RELEASE_WEAK \genblk1[191].rrel ( .Q(L[191]), .E(ren));
Q_REGFORCE \genblk1[191].rfrc ( .Q(L[191]), .A(V[191]), .E(fen));
Q_RELEASE_WEAK \genblk1[190].rrel ( .Q(L[190]), .E(ren));
Q_REGFORCE \genblk1[190].rfrc ( .Q(L[190]), .A(V[190]), .E(fen));
Q_RELEASE_WEAK \genblk1[189].rrel ( .Q(L[189]), .E(ren));
Q_REGFORCE \genblk1[189].rfrc ( .Q(L[189]), .A(V[189]), .E(fen));
Q_RELEASE_WEAK \genblk1[188].rrel ( .Q(L[188]), .E(ren));
Q_REGFORCE \genblk1[188].rfrc ( .Q(L[188]), .A(V[188]), .E(fen));
Q_RELEASE_WEAK \genblk1[187].rrel ( .Q(L[187]), .E(ren));
Q_REGFORCE \genblk1[187].rfrc ( .Q(L[187]), .A(V[187]), .E(fen));
Q_RELEASE_WEAK \genblk1[186].rrel ( .Q(L[186]), .E(ren));
Q_REGFORCE \genblk1[186].rfrc ( .Q(L[186]), .A(V[186]), .E(fen));
Q_RELEASE_WEAK \genblk1[185].rrel ( .Q(L[185]), .E(ren));
Q_REGFORCE \genblk1[185].rfrc ( .Q(L[185]), .A(V[185]), .E(fen));
Q_RELEASE_WEAK \genblk1[184].rrel ( .Q(L[184]), .E(ren));
Q_REGFORCE \genblk1[184].rfrc ( .Q(L[184]), .A(V[184]), .E(fen));
Q_RELEASE_WEAK \genblk1[183].rrel ( .Q(L[183]), .E(ren));
Q_REGFORCE \genblk1[183].rfrc ( .Q(L[183]), .A(V[183]), .E(fen));
Q_RELEASE_WEAK \genblk1[182].rrel ( .Q(L[182]), .E(ren));
Q_REGFORCE \genblk1[182].rfrc ( .Q(L[182]), .A(V[182]), .E(fen));
Q_RELEASE_WEAK \genblk1[181].rrel ( .Q(L[181]), .E(ren));
Q_REGFORCE \genblk1[181].rfrc ( .Q(L[181]), .A(V[181]), .E(fen));
Q_RELEASE_WEAK \genblk1[180].rrel ( .Q(L[180]), .E(ren));
Q_REGFORCE \genblk1[180].rfrc ( .Q(L[180]), .A(V[180]), .E(fen));
Q_RELEASE_WEAK \genblk1[179].rrel ( .Q(L[179]), .E(ren));
Q_REGFORCE \genblk1[179].rfrc ( .Q(L[179]), .A(V[179]), .E(fen));
Q_RELEASE_WEAK \genblk1[178].rrel ( .Q(L[178]), .E(ren));
Q_REGFORCE \genblk1[178].rfrc ( .Q(L[178]), .A(V[178]), .E(fen));
Q_RELEASE_WEAK \genblk1[177].rrel ( .Q(L[177]), .E(ren));
Q_REGFORCE \genblk1[177].rfrc ( .Q(L[177]), .A(V[177]), .E(fen));
Q_RELEASE_WEAK \genblk1[176].rrel ( .Q(L[176]), .E(ren));
Q_REGFORCE \genblk1[176].rfrc ( .Q(L[176]), .A(V[176]), .E(fen));
Q_RELEASE_WEAK \genblk1[175].rrel ( .Q(L[175]), .E(ren));
Q_REGFORCE \genblk1[175].rfrc ( .Q(L[175]), .A(V[175]), .E(fen));
Q_RELEASE_WEAK \genblk1[174].rrel ( .Q(L[174]), .E(ren));
Q_REGFORCE \genblk1[174].rfrc ( .Q(L[174]), .A(V[174]), .E(fen));
Q_RELEASE_WEAK \genblk1[173].rrel ( .Q(L[173]), .E(ren));
Q_REGFORCE \genblk1[173].rfrc ( .Q(L[173]), .A(V[173]), .E(fen));
Q_RELEASE_WEAK \genblk1[172].rrel ( .Q(L[172]), .E(ren));
Q_REGFORCE \genblk1[172].rfrc ( .Q(L[172]), .A(V[172]), .E(fen));
Q_RELEASE_WEAK \genblk1[171].rrel ( .Q(L[171]), .E(ren));
Q_REGFORCE \genblk1[171].rfrc ( .Q(L[171]), .A(V[171]), .E(fen));
Q_RELEASE_WEAK \genblk1[170].rrel ( .Q(L[170]), .E(ren));
Q_REGFORCE \genblk1[170].rfrc ( .Q(L[170]), .A(V[170]), .E(fen));
Q_RELEASE_WEAK \genblk1[169].rrel ( .Q(L[169]), .E(ren));
Q_REGFORCE \genblk1[169].rfrc ( .Q(L[169]), .A(V[169]), .E(fen));
Q_RELEASE_WEAK \genblk1[168].rrel ( .Q(L[168]), .E(ren));
Q_REGFORCE \genblk1[168].rfrc ( .Q(L[168]), .A(V[168]), .E(fen));
Q_RELEASE_WEAK \genblk1[167].rrel ( .Q(L[167]), .E(ren));
Q_REGFORCE \genblk1[167].rfrc ( .Q(L[167]), .A(V[167]), .E(fen));
Q_RELEASE_WEAK \genblk1[166].rrel ( .Q(L[166]), .E(ren));
Q_REGFORCE \genblk1[166].rfrc ( .Q(L[166]), .A(V[166]), .E(fen));
Q_RELEASE_WEAK \genblk1[165].rrel ( .Q(L[165]), .E(ren));
Q_REGFORCE \genblk1[165].rfrc ( .Q(L[165]), .A(V[165]), .E(fen));
Q_RELEASE_WEAK \genblk1[164].rrel ( .Q(L[164]), .E(ren));
Q_REGFORCE \genblk1[164].rfrc ( .Q(L[164]), .A(V[164]), .E(fen));
Q_RELEASE_WEAK \genblk1[163].rrel ( .Q(L[163]), .E(ren));
Q_REGFORCE \genblk1[163].rfrc ( .Q(L[163]), .A(V[163]), .E(fen));
Q_RELEASE_WEAK \genblk1[162].rrel ( .Q(L[162]), .E(ren));
Q_REGFORCE \genblk1[162].rfrc ( .Q(L[162]), .A(V[162]), .E(fen));
Q_RELEASE_WEAK \genblk1[161].rrel ( .Q(L[161]), .E(ren));
Q_REGFORCE \genblk1[161].rfrc ( .Q(L[161]), .A(V[161]), .E(fen));
Q_RELEASE_WEAK \genblk1[160].rrel ( .Q(L[160]), .E(ren));
Q_REGFORCE \genblk1[160].rfrc ( .Q(L[160]), .A(V[160]), .E(fen));
Q_RELEASE_WEAK \genblk1[159].rrel ( .Q(L[159]), .E(ren));
Q_REGFORCE \genblk1[159].rfrc ( .Q(L[159]), .A(V[159]), .E(fen));
Q_RELEASE_WEAK \genblk1[158].rrel ( .Q(L[158]), .E(ren));
Q_REGFORCE \genblk1[158].rfrc ( .Q(L[158]), .A(V[158]), .E(fen));
Q_RELEASE_WEAK \genblk1[157].rrel ( .Q(L[157]), .E(ren));
Q_REGFORCE \genblk1[157].rfrc ( .Q(L[157]), .A(V[157]), .E(fen));
Q_RELEASE_WEAK \genblk1[156].rrel ( .Q(L[156]), .E(ren));
Q_REGFORCE \genblk1[156].rfrc ( .Q(L[156]), .A(V[156]), .E(fen));
Q_RELEASE_WEAK \genblk1[155].rrel ( .Q(L[155]), .E(ren));
Q_REGFORCE \genblk1[155].rfrc ( .Q(L[155]), .A(V[155]), .E(fen));
Q_RELEASE_WEAK \genblk1[154].rrel ( .Q(L[154]), .E(ren));
Q_REGFORCE \genblk1[154].rfrc ( .Q(L[154]), .A(V[154]), .E(fen));
Q_RELEASE_WEAK \genblk1[153].rrel ( .Q(L[153]), .E(ren));
Q_REGFORCE \genblk1[153].rfrc ( .Q(L[153]), .A(V[153]), .E(fen));
Q_RELEASE_WEAK \genblk1[152].rrel ( .Q(L[152]), .E(ren));
Q_REGFORCE \genblk1[152].rfrc ( .Q(L[152]), .A(V[152]), .E(fen));
Q_RELEASE_WEAK \genblk1[151].rrel ( .Q(L[151]), .E(ren));
Q_REGFORCE \genblk1[151].rfrc ( .Q(L[151]), .A(V[151]), .E(fen));
Q_RELEASE_WEAK \genblk1[150].rrel ( .Q(L[150]), .E(ren));
Q_REGFORCE \genblk1[150].rfrc ( .Q(L[150]), .A(V[150]), .E(fen));
Q_RELEASE_WEAK \genblk1[149].rrel ( .Q(L[149]), .E(ren));
Q_REGFORCE \genblk1[149].rfrc ( .Q(L[149]), .A(V[149]), .E(fen));
Q_RELEASE_WEAK \genblk1[148].rrel ( .Q(L[148]), .E(ren));
Q_REGFORCE \genblk1[148].rfrc ( .Q(L[148]), .A(V[148]), .E(fen));
Q_RELEASE_WEAK \genblk1[147].rrel ( .Q(L[147]), .E(ren));
Q_REGFORCE \genblk1[147].rfrc ( .Q(L[147]), .A(V[147]), .E(fen));
Q_RELEASE_WEAK \genblk1[146].rrel ( .Q(L[146]), .E(ren));
Q_REGFORCE \genblk1[146].rfrc ( .Q(L[146]), .A(V[146]), .E(fen));
Q_RELEASE_WEAK \genblk1[145].rrel ( .Q(L[145]), .E(ren));
Q_REGFORCE \genblk1[145].rfrc ( .Q(L[145]), .A(V[145]), .E(fen));
Q_RELEASE_WEAK \genblk1[144].rrel ( .Q(L[144]), .E(ren));
Q_REGFORCE \genblk1[144].rfrc ( .Q(L[144]), .A(V[144]), .E(fen));
Q_RELEASE_WEAK \genblk1[143].rrel ( .Q(L[143]), .E(ren));
Q_REGFORCE \genblk1[143].rfrc ( .Q(L[143]), .A(V[143]), .E(fen));
Q_RELEASE_WEAK \genblk1[142].rrel ( .Q(L[142]), .E(ren));
Q_REGFORCE \genblk1[142].rfrc ( .Q(L[142]), .A(V[142]), .E(fen));
Q_RELEASE_WEAK \genblk1[141].rrel ( .Q(L[141]), .E(ren));
Q_REGFORCE \genblk1[141].rfrc ( .Q(L[141]), .A(V[141]), .E(fen));
Q_RELEASE_WEAK \genblk1[140].rrel ( .Q(L[140]), .E(ren));
Q_REGFORCE \genblk1[140].rfrc ( .Q(L[140]), .A(V[140]), .E(fen));
Q_RELEASE_WEAK \genblk1[139].rrel ( .Q(L[139]), .E(ren));
Q_REGFORCE \genblk1[139].rfrc ( .Q(L[139]), .A(V[139]), .E(fen));
Q_RELEASE_WEAK \genblk1[138].rrel ( .Q(L[138]), .E(ren));
Q_REGFORCE \genblk1[138].rfrc ( .Q(L[138]), .A(V[138]), .E(fen));
Q_RELEASE_WEAK \genblk1[137].rrel ( .Q(L[137]), .E(ren));
Q_REGFORCE \genblk1[137].rfrc ( .Q(L[137]), .A(V[137]), .E(fen));
Q_RELEASE_WEAK \genblk1[136].rrel ( .Q(L[136]), .E(ren));
Q_REGFORCE \genblk1[136].rfrc ( .Q(L[136]), .A(V[136]), .E(fen));
Q_RELEASE_WEAK \genblk1[135].rrel ( .Q(L[135]), .E(ren));
Q_REGFORCE \genblk1[135].rfrc ( .Q(L[135]), .A(V[135]), .E(fen));
Q_RELEASE_WEAK \genblk1[134].rrel ( .Q(L[134]), .E(ren));
Q_REGFORCE \genblk1[134].rfrc ( .Q(L[134]), .A(V[134]), .E(fen));
Q_RELEASE_WEAK \genblk1[133].rrel ( .Q(L[133]), .E(ren));
Q_REGFORCE \genblk1[133].rfrc ( .Q(L[133]), .A(V[133]), .E(fen));
Q_RELEASE_WEAK \genblk1[132].rrel ( .Q(L[132]), .E(ren));
Q_REGFORCE \genblk1[132].rfrc ( .Q(L[132]), .A(V[132]), .E(fen));
Q_RELEASE_WEAK \genblk1[131].rrel ( .Q(L[131]), .E(ren));
Q_REGFORCE \genblk1[131].rfrc ( .Q(L[131]), .A(V[131]), .E(fen));
Q_RELEASE_WEAK \genblk1[130].rrel ( .Q(L[130]), .E(ren));
Q_REGFORCE \genblk1[130].rfrc ( .Q(L[130]), .A(V[130]), .E(fen));
Q_RELEASE_WEAK \genblk1[129].rrel ( .Q(L[129]), .E(ren));
Q_REGFORCE \genblk1[129].rfrc ( .Q(L[129]), .A(V[129]), .E(fen));
Q_RELEASE_WEAK \genblk1[128].rrel ( .Q(L[128]), .E(ren));
Q_REGFORCE \genblk1[128].rfrc ( .Q(L[128]), .A(V[128]), .E(fen));
Q_RELEASE_WEAK \genblk1[127].rrel ( .Q(L[127]), .E(ren));
Q_REGFORCE \genblk1[127].rfrc ( .Q(L[127]), .A(V[127]), .E(fen));
Q_RELEASE_WEAK \genblk1[126].rrel ( .Q(L[126]), .E(ren));
Q_REGFORCE \genblk1[126].rfrc ( .Q(L[126]), .A(V[126]), .E(fen));
Q_RELEASE_WEAK \genblk1[125].rrel ( .Q(L[125]), .E(ren));
Q_REGFORCE \genblk1[125].rfrc ( .Q(L[125]), .A(V[125]), .E(fen));
Q_RELEASE_WEAK \genblk1[124].rrel ( .Q(L[124]), .E(ren));
Q_REGFORCE \genblk1[124].rfrc ( .Q(L[124]), .A(V[124]), .E(fen));
Q_RELEASE_WEAK \genblk1[123].rrel ( .Q(L[123]), .E(ren));
Q_REGFORCE \genblk1[123].rfrc ( .Q(L[123]), .A(V[123]), .E(fen));
Q_RELEASE_WEAK \genblk1[122].rrel ( .Q(L[122]), .E(ren));
Q_REGFORCE \genblk1[122].rfrc ( .Q(L[122]), .A(V[122]), .E(fen));
Q_RELEASE_WEAK \genblk1[121].rrel ( .Q(L[121]), .E(ren));
Q_REGFORCE \genblk1[121].rfrc ( .Q(L[121]), .A(V[121]), .E(fen));
Q_RELEASE_WEAK \genblk1[120].rrel ( .Q(L[120]), .E(ren));
Q_REGFORCE \genblk1[120].rfrc ( .Q(L[120]), .A(V[120]), .E(fen));
Q_RELEASE_WEAK \genblk1[119].rrel ( .Q(L[119]), .E(ren));
Q_REGFORCE \genblk1[119].rfrc ( .Q(L[119]), .A(V[119]), .E(fen));
Q_RELEASE_WEAK \genblk1[118].rrel ( .Q(L[118]), .E(ren));
Q_REGFORCE \genblk1[118].rfrc ( .Q(L[118]), .A(V[118]), .E(fen));
Q_RELEASE_WEAK \genblk1[117].rrel ( .Q(L[117]), .E(ren));
Q_REGFORCE \genblk1[117].rfrc ( .Q(L[117]), .A(V[117]), .E(fen));
Q_RELEASE_WEAK \genblk1[116].rrel ( .Q(L[116]), .E(ren));
Q_REGFORCE \genblk1[116].rfrc ( .Q(L[116]), .A(V[116]), .E(fen));
Q_RELEASE_WEAK \genblk1[115].rrel ( .Q(L[115]), .E(ren));
Q_REGFORCE \genblk1[115].rfrc ( .Q(L[115]), .A(V[115]), .E(fen));
Q_RELEASE_WEAK \genblk1[114].rrel ( .Q(L[114]), .E(ren));
Q_REGFORCE \genblk1[114].rfrc ( .Q(L[114]), .A(V[114]), .E(fen));
Q_RELEASE_WEAK \genblk1[113].rrel ( .Q(L[113]), .E(ren));
Q_REGFORCE \genblk1[113].rfrc ( .Q(L[113]), .A(V[113]), .E(fen));
Q_RELEASE_WEAK \genblk1[112].rrel ( .Q(L[112]), .E(ren));
Q_REGFORCE \genblk1[112].rfrc ( .Q(L[112]), .A(V[112]), .E(fen));
Q_RELEASE_WEAK \genblk1[111].rrel ( .Q(L[111]), .E(ren));
Q_REGFORCE \genblk1[111].rfrc ( .Q(L[111]), .A(V[111]), .E(fen));
Q_RELEASE_WEAK \genblk1[110].rrel ( .Q(L[110]), .E(ren));
Q_REGFORCE \genblk1[110].rfrc ( .Q(L[110]), .A(V[110]), .E(fen));
Q_RELEASE_WEAK \genblk1[109].rrel ( .Q(L[109]), .E(ren));
Q_REGFORCE \genblk1[109].rfrc ( .Q(L[109]), .A(V[109]), .E(fen));
Q_RELEASE_WEAK \genblk1[108].rrel ( .Q(L[108]), .E(ren));
Q_REGFORCE \genblk1[108].rfrc ( .Q(L[108]), .A(V[108]), .E(fen));
Q_RELEASE_WEAK \genblk1[107].rrel ( .Q(L[107]), .E(ren));
Q_REGFORCE \genblk1[107].rfrc ( .Q(L[107]), .A(V[107]), .E(fen));
Q_RELEASE_WEAK \genblk1[106].rrel ( .Q(L[106]), .E(ren));
Q_REGFORCE \genblk1[106].rfrc ( .Q(L[106]), .A(V[106]), .E(fen));
Q_RELEASE_WEAK \genblk1[105].rrel ( .Q(L[105]), .E(ren));
Q_REGFORCE \genblk1[105].rfrc ( .Q(L[105]), .A(V[105]), .E(fen));
Q_RELEASE_WEAK \genblk1[104].rrel ( .Q(L[104]), .E(ren));
Q_REGFORCE \genblk1[104].rfrc ( .Q(L[104]), .A(V[104]), .E(fen));
Q_RELEASE_WEAK \genblk1[103].rrel ( .Q(L[103]), .E(ren));
Q_REGFORCE \genblk1[103].rfrc ( .Q(L[103]), .A(V[103]), .E(fen));
Q_RELEASE_WEAK \genblk1[102].rrel ( .Q(L[102]), .E(ren));
Q_REGFORCE \genblk1[102].rfrc ( .Q(L[102]), .A(V[102]), .E(fen));
Q_RELEASE_WEAK \genblk1[101].rrel ( .Q(L[101]), .E(ren));
Q_REGFORCE \genblk1[101].rfrc ( .Q(L[101]), .A(V[101]), .E(fen));
Q_RELEASE_WEAK \genblk1[100].rrel ( .Q(L[100]), .E(ren));
Q_REGFORCE \genblk1[100].rfrc ( .Q(L[100]), .A(V[100]), .E(fen));
Q_RELEASE_WEAK \genblk1[99].rrel ( .Q(L[99]), .E(ren));
Q_REGFORCE \genblk1[99].rfrc ( .Q(L[99]), .A(V[99]), .E(fen));
Q_RELEASE_WEAK \genblk1[98].rrel ( .Q(L[98]), .E(ren));
Q_REGFORCE \genblk1[98].rfrc ( .Q(L[98]), .A(V[98]), .E(fen));
Q_RELEASE_WEAK \genblk1[97].rrel ( .Q(L[97]), .E(ren));
Q_REGFORCE \genblk1[97].rfrc ( .Q(L[97]), .A(V[97]), .E(fen));
Q_RELEASE_WEAK \genblk1[96].rrel ( .Q(L[96]), .E(ren));
Q_REGFORCE \genblk1[96].rfrc ( .Q(L[96]), .A(V[96]), .E(fen));
Q_RELEASE_WEAK \genblk1[95].rrel ( .Q(L[95]), .E(ren));
Q_REGFORCE \genblk1[95].rfrc ( .Q(L[95]), .A(V[95]), .E(fen));
Q_RELEASE_WEAK \genblk1[94].rrel ( .Q(L[94]), .E(ren));
Q_REGFORCE \genblk1[94].rfrc ( .Q(L[94]), .A(V[94]), .E(fen));
Q_RELEASE_WEAK \genblk1[93].rrel ( .Q(L[93]), .E(ren));
Q_REGFORCE \genblk1[93].rfrc ( .Q(L[93]), .A(V[93]), .E(fen));
Q_RELEASE_WEAK \genblk1[92].rrel ( .Q(L[92]), .E(ren));
Q_REGFORCE \genblk1[92].rfrc ( .Q(L[92]), .A(V[92]), .E(fen));
Q_RELEASE_WEAK \genblk1[91].rrel ( .Q(L[91]), .E(ren));
Q_REGFORCE \genblk1[91].rfrc ( .Q(L[91]), .A(V[91]), .E(fen));
Q_RELEASE_WEAK \genblk1[90].rrel ( .Q(L[90]), .E(ren));
Q_REGFORCE \genblk1[90].rfrc ( .Q(L[90]), .A(V[90]), .E(fen));
Q_RELEASE_WEAK \genblk1[89].rrel ( .Q(L[89]), .E(ren));
Q_REGFORCE \genblk1[89].rfrc ( .Q(L[89]), .A(V[89]), .E(fen));
Q_RELEASE_WEAK \genblk1[88].rrel ( .Q(L[88]), .E(ren));
Q_REGFORCE \genblk1[88].rfrc ( .Q(L[88]), .A(V[88]), .E(fen));
Q_RELEASE_WEAK \genblk1[87].rrel ( .Q(L[87]), .E(ren));
Q_REGFORCE \genblk1[87].rfrc ( .Q(L[87]), .A(V[87]), .E(fen));
Q_RELEASE_WEAK \genblk1[86].rrel ( .Q(L[86]), .E(ren));
Q_REGFORCE \genblk1[86].rfrc ( .Q(L[86]), .A(V[86]), .E(fen));
Q_RELEASE_WEAK \genblk1[85].rrel ( .Q(L[85]), .E(ren));
Q_REGFORCE \genblk1[85].rfrc ( .Q(L[85]), .A(V[85]), .E(fen));
Q_RELEASE_WEAK \genblk1[84].rrel ( .Q(L[84]), .E(ren));
Q_REGFORCE \genblk1[84].rfrc ( .Q(L[84]), .A(V[84]), .E(fen));
Q_RELEASE_WEAK \genblk1[83].rrel ( .Q(L[83]), .E(ren));
Q_REGFORCE \genblk1[83].rfrc ( .Q(L[83]), .A(V[83]), .E(fen));
Q_RELEASE_WEAK \genblk1[82].rrel ( .Q(L[82]), .E(ren));
Q_REGFORCE \genblk1[82].rfrc ( .Q(L[82]), .A(V[82]), .E(fen));
Q_RELEASE_WEAK \genblk1[81].rrel ( .Q(L[81]), .E(ren));
Q_REGFORCE \genblk1[81].rfrc ( .Q(L[81]), .A(V[81]), .E(fen));
Q_RELEASE_WEAK \genblk1[80].rrel ( .Q(L[80]), .E(ren));
Q_REGFORCE \genblk1[80].rfrc ( .Q(L[80]), .A(V[80]), .E(fen));
Q_RELEASE_WEAK \genblk1[79].rrel ( .Q(L[79]), .E(ren));
Q_REGFORCE \genblk1[79].rfrc ( .Q(L[79]), .A(V[79]), .E(fen));
Q_RELEASE_WEAK \genblk1[78].rrel ( .Q(L[78]), .E(ren));
Q_REGFORCE \genblk1[78].rfrc ( .Q(L[78]), .A(V[78]), .E(fen));
Q_RELEASE_WEAK \genblk1[77].rrel ( .Q(L[77]), .E(ren));
Q_REGFORCE \genblk1[77].rfrc ( .Q(L[77]), .A(V[77]), .E(fen));
Q_RELEASE_WEAK \genblk1[76].rrel ( .Q(L[76]), .E(ren));
Q_REGFORCE \genblk1[76].rfrc ( .Q(L[76]), .A(V[76]), .E(fen));
Q_RELEASE_WEAK \genblk1[75].rrel ( .Q(L[75]), .E(ren));
Q_REGFORCE \genblk1[75].rfrc ( .Q(L[75]), .A(V[75]), .E(fen));
Q_RELEASE_WEAK \genblk1[74].rrel ( .Q(L[74]), .E(ren));
Q_REGFORCE \genblk1[74].rfrc ( .Q(L[74]), .A(V[74]), .E(fen));
Q_RELEASE_WEAK \genblk1[73].rrel ( .Q(L[73]), .E(ren));
Q_REGFORCE \genblk1[73].rfrc ( .Q(L[73]), .A(V[73]), .E(fen));
Q_RELEASE_WEAK \genblk1[72].rrel ( .Q(L[72]), .E(ren));
Q_REGFORCE \genblk1[72].rfrc ( .Q(L[72]), .A(V[72]), .E(fen));
Q_RELEASE_WEAK \genblk1[71].rrel ( .Q(L[71]), .E(ren));
Q_REGFORCE \genblk1[71].rfrc ( .Q(L[71]), .A(V[71]), .E(fen));
Q_RELEASE_WEAK \genblk1[70].rrel ( .Q(L[70]), .E(ren));
Q_REGFORCE \genblk1[70].rfrc ( .Q(L[70]), .A(V[70]), .E(fen));
Q_RELEASE_WEAK \genblk1[69].rrel ( .Q(L[69]), .E(ren));
Q_REGFORCE \genblk1[69].rfrc ( .Q(L[69]), .A(V[69]), .E(fen));
Q_RELEASE_WEAK \genblk1[68].rrel ( .Q(L[68]), .E(ren));
Q_REGFORCE \genblk1[68].rfrc ( .Q(L[68]), .A(V[68]), .E(fen));
Q_RELEASE_WEAK \genblk1[67].rrel ( .Q(L[67]), .E(ren));
Q_REGFORCE \genblk1[67].rfrc ( .Q(L[67]), .A(V[67]), .E(fen));
Q_RELEASE_WEAK \genblk1[66].rrel ( .Q(L[66]), .E(ren));
Q_REGFORCE \genblk1[66].rfrc ( .Q(L[66]), .A(V[66]), .E(fen));
Q_RELEASE_WEAK \genblk1[65].rrel ( .Q(L[65]), .E(ren));
Q_REGFORCE \genblk1[65].rfrc ( .Q(L[65]), .A(V[65]), .E(fen));
Q_RELEASE_WEAK \genblk1[64].rrel ( .Q(L[64]), .E(ren));
Q_REGFORCE \genblk1[64].rfrc ( .Q(L[64]), .A(V[64]), .E(fen));
Q_RELEASE_WEAK \genblk1[63].rrel ( .Q(L[63]), .E(ren));
Q_REGFORCE \genblk1[63].rfrc ( .Q(L[63]), .A(V[63]), .E(fen));
Q_RELEASE_WEAK \genblk1[62].rrel ( .Q(L[62]), .E(ren));
Q_REGFORCE \genblk1[62].rfrc ( .Q(L[62]), .A(V[62]), .E(fen));
Q_RELEASE_WEAK \genblk1[61].rrel ( .Q(L[61]), .E(ren));
Q_REGFORCE \genblk1[61].rfrc ( .Q(L[61]), .A(V[61]), .E(fen));
Q_RELEASE_WEAK \genblk1[60].rrel ( .Q(L[60]), .E(ren));
Q_REGFORCE \genblk1[60].rfrc ( .Q(L[60]), .A(V[60]), .E(fen));
Q_RELEASE_WEAK \genblk1[59].rrel ( .Q(L[59]), .E(ren));
Q_REGFORCE \genblk1[59].rfrc ( .Q(L[59]), .A(V[59]), .E(fen));
Q_RELEASE_WEAK \genblk1[58].rrel ( .Q(L[58]), .E(ren));
Q_REGFORCE \genblk1[58].rfrc ( .Q(L[58]), .A(V[58]), .E(fen));
Q_RELEASE_WEAK \genblk1[57].rrel ( .Q(L[57]), .E(ren));
Q_REGFORCE \genblk1[57].rfrc ( .Q(L[57]), .A(V[57]), .E(fen));
Q_RELEASE_WEAK \genblk1[56].rrel ( .Q(L[56]), .E(ren));
Q_REGFORCE \genblk1[56].rfrc ( .Q(L[56]), .A(V[56]), .E(fen));
Q_RELEASE_WEAK \genblk1[55].rrel ( .Q(L[55]), .E(ren));
Q_REGFORCE \genblk1[55].rfrc ( .Q(L[55]), .A(V[55]), .E(fen));
Q_RELEASE_WEAK \genblk1[54].rrel ( .Q(L[54]), .E(ren));
Q_REGFORCE \genblk1[54].rfrc ( .Q(L[54]), .A(V[54]), .E(fen));
Q_RELEASE_WEAK \genblk1[53].rrel ( .Q(L[53]), .E(ren));
Q_REGFORCE \genblk1[53].rfrc ( .Q(L[53]), .A(V[53]), .E(fen));
Q_RELEASE_WEAK \genblk1[52].rrel ( .Q(L[52]), .E(ren));
Q_REGFORCE \genblk1[52].rfrc ( .Q(L[52]), .A(V[52]), .E(fen));
Q_RELEASE_WEAK \genblk1[51].rrel ( .Q(L[51]), .E(ren));
Q_REGFORCE \genblk1[51].rfrc ( .Q(L[51]), .A(V[51]), .E(fen));
Q_RELEASE_WEAK \genblk1[50].rrel ( .Q(L[50]), .E(ren));
Q_REGFORCE \genblk1[50].rfrc ( .Q(L[50]), .A(V[50]), .E(fen));
Q_RELEASE_WEAK \genblk1[49].rrel ( .Q(L[49]), .E(ren));
Q_REGFORCE \genblk1[49].rfrc ( .Q(L[49]), .A(V[49]), .E(fen));
Q_RELEASE_WEAK \genblk1[48].rrel ( .Q(L[48]), .E(ren));
Q_REGFORCE \genblk1[48].rfrc ( .Q(L[48]), .A(V[48]), .E(fen));
Q_RELEASE_WEAK \genblk1[47].rrel ( .Q(L[47]), .E(ren));
Q_REGFORCE \genblk1[47].rfrc ( .Q(L[47]), .A(V[47]), .E(fen));
Q_RELEASE_WEAK \genblk1[46].rrel ( .Q(L[46]), .E(ren));
Q_REGFORCE \genblk1[46].rfrc ( .Q(L[46]), .A(V[46]), .E(fen));
Q_RELEASE_WEAK \genblk1[45].rrel ( .Q(L[45]), .E(ren));
Q_REGFORCE \genblk1[45].rfrc ( .Q(L[45]), .A(V[45]), .E(fen));
Q_RELEASE_WEAK \genblk1[44].rrel ( .Q(L[44]), .E(ren));
Q_REGFORCE \genblk1[44].rfrc ( .Q(L[44]), .A(V[44]), .E(fen));
Q_RELEASE_WEAK \genblk1[43].rrel ( .Q(L[43]), .E(ren));
Q_REGFORCE \genblk1[43].rfrc ( .Q(L[43]), .A(V[43]), .E(fen));
Q_RELEASE_WEAK \genblk1[42].rrel ( .Q(L[42]), .E(ren));
Q_REGFORCE \genblk1[42].rfrc ( .Q(L[42]), .A(V[42]), .E(fen));
Q_RELEASE_WEAK \genblk1[41].rrel ( .Q(L[41]), .E(ren));
Q_REGFORCE \genblk1[41].rfrc ( .Q(L[41]), .A(V[41]), .E(fen));
Q_RELEASE_WEAK \genblk1[40].rrel ( .Q(L[40]), .E(ren));
Q_REGFORCE \genblk1[40].rfrc ( .Q(L[40]), .A(V[40]), .E(fen));
Q_RELEASE_WEAK \genblk1[39].rrel ( .Q(L[39]), .E(ren));
Q_REGFORCE \genblk1[39].rfrc ( .Q(L[39]), .A(V[39]), .E(fen));
Q_RELEASE_WEAK \genblk1[38].rrel ( .Q(L[38]), .E(ren));
Q_REGFORCE \genblk1[38].rfrc ( .Q(L[38]), .A(V[38]), .E(fen));
Q_RELEASE_WEAK \genblk1[37].rrel ( .Q(L[37]), .E(ren));
Q_REGFORCE \genblk1[37].rfrc ( .Q(L[37]), .A(V[37]), .E(fen));
Q_RELEASE_WEAK \genblk1[36].rrel ( .Q(L[36]), .E(ren));
Q_REGFORCE \genblk1[36].rfrc ( .Q(L[36]), .A(V[36]), .E(fen));
Q_RELEASE_WEAK \genblk1[35].rrel ( .Q(L[35]), .E(ren));
Q_REGFORCE \genblk1[35].rfrc ( .Q(L[35]), .A(V[35]), .E(fen));
Q_RELEASE_WEAK \genblk1[34].rrel ( .Q(L[34]), .E(ren));
Q_REGFORCE \genblk1[34].rfrc ( .Q(L[34]), .A(V[34]), .E(fen));
Q_RELEASE_WEAK \genblk1[33].rrel ( .Q(L[33]), .E(ren));
Q_REGFORCE \genblk1[33].rfrc ( .Q(L[33]), .A(V[33]), .E(fen));
Q_RELEASE_WEAK \genblk1[32].rrel ( .Q(L[32]), .E(ren));
Q_REGFORCE \genblk1[32].rfrc ( .Q(L[32]), .A(V[32]), .E(fen));
Q_RELEASE_WEAK \genblk1[31].rrel ( .Q(L[31]), .E(ren));
Q_REGFORCE \genblk1[31].rfrc ( .Q(L[31]), .A(V[31]), .E(fen));
Q_RELEASE_WEAK \genblk1[30].rrel ( .Q(L[30]), .E(ren));
Q_REGFORCE \genblk1[30].rfrc ( .Q(L[30]), .A(V[30]), .E(fen));
Q_RELEASE_WEAK \genblk1[29].rrel ( .Q(L[29]), .E(ren));
Q_REGFORCE \genblk1[29].rfrc ( .Q(L[29]), .A(V[29]), .E(fen));
Q_RELEASE_WEAK \genblk1[28].rrel ( .Q(L[28]), .E(ren));
Q_REGFORCE \genblk1[28].rfrc ( .Q(L[28]), .A(V[28]), .E(fen));
Q_RELEASE_WEAK \genblk1[27].rrel ( .Q(L[27]), .E(ren));
Q_REGFORCE \genblk1[27].rfrc ( .Q(L[27]), .A(V[27]), .E(fen));
Q_RELEASE_WEAK \genblk1[26].rrel ( .Q(L[26]), .E(ren));
Q_REGFORCE \genblk1[26].rfrc ( .Q(L[26]), .A(V[26]), .E(fen));
Q_RELEASE_WEAK \genblk1[25].rrel ( .Q(L[25]), .E(ren));
Q_REGFORCE \genblk1[25].rfrc ( .Q(L[25]), .A(V[25]), .E(fen));
Q_RELEASE_WEAK \genblk1[24].rrel ( .Q(L[24]), .E(ren));
Q_REGFORCE \genblk1[24].rfrc ( .Q(L[24]), .A(V[24]), .E(fen));
Q_RELEASE_WEAK \genblk1[23].rrel ( .Q(L[23]), .E(ren));
Q_REGFORCE \genblk1[23].rfrc ( .Q(L[23]), .A(V[23]), .E(fen));
Q_RELEASE_WEAK \genblk1[22].rrel ( .Q(L[22]), .E(ren));
Q_REGFORCE \genblk1[22].rfrc ( .Q(L[22]), .A(V[22]), .E(fen));
Q_RELEASE_WEAK \genblk1[21].rrel ( .Q(L[21]), .E(ren));
Q_REGFORCE \genblk1[21].rfrc ( .Q(L[21]), .A(V[21]), .E(fen));
Q_RELEASE_WEAK \genblk1[20].rrel ( .Q(L[20]), .E(ren));
Q_REGFORCE \genblk1[20].rfrc ( .Q(L[20]), .A(V[20]), .E(fen));
Q_RELEASE_WEAK \genblk1[19].rrel ( .Q(L[19]), .E(ren));
Q_REGFORCE \genblk1[19].rfrc ( .Q(L[19]), .A(V[19]), .E(fen));
Q_RELEASE_WEAK \genblk1[18].rrel ( .Q(L[18]), .E(ren));
Q_REGFORCE \genblk1[18].rfrc ( .Q(L[18]), .A(V[18]), .E(fen));
Q_RELEASE_WEAK \genblk1[17].rrel ( .Q(L[17]), .E(ren));
Q_REGFORCE \genblk1[17].rfrc ( .Q(L[17]), .A(V[17]), .E(fen));
Q_RELEASE_WEAK \genblk1[16].rrel ( .Q(L[16]), .E(ren));
Q_REGFORCE \genblk1[16].rfrc ( .Q(L[16]), .A(V[16]), .E(fen));
Q_RELEASE_WEAK \genblk1[15].rrel ( .Q(L[15]), .E(ren));
Q_REGFORCE \genblk1[15].rfrc ( .Q(L[15]), .A(V[15]), .E(fen));
Q_RELEASE_WEAK \genblk1[14].rrel ( .Q(L[14]), .E(ren));
Q_REGFORCE \genblk1[14].rfrc ( .Q(L[14]), .A(V[14]), .E(fen));
Q_RELEASE_WEAK \genblk1[13].rrel ( .Q(L[13]), .E(ren));
Q_REGFORCE \genblk1[13].rfrc ( .Q(L[13]), .A(V[13]), .E(fen));
Q_RELEASE_WEAK \genblk1[12].rrel ( .Q(L[12]), .E(ren));
Q_REGFORCE \genblk1[12].rfrc ( .Q(L[12]), .A(V[12]), .E(fen));
Q_RELEASE_WEAK \genblk1[11].rrel ( .Q(L[11]), .E(ren));
Q_REGFORCE \genblk1[11].rfrc ( .Q(L[11]), .A(V[11]), .E(fen));
Q_RELEASE_WEAK \genblk1[10].rrel ( .Q(L[10]), .E(ren));
Q_REGFORCE \genblk1[10].rfrc ( .Q(L[10]), .A(V[10]), .E(fen));
Q_RELEASE_WEAK \genblk1[9].rrel ( .Q(L[9]), .E(ren));
Q_REGFORCE \genblk1[9].rfrc ( .Q(L[9]), .A(V[9]), .E(fen));
Q_RELEASE_WEAK \genblk1[8].rrel ( .Q(L[8]), .E(ren));
Q_REGFORCE \genblk1[8].rfrc ( .Q(L[8]), .A(V[8]), .E(fen));
Q_RELEASE_WEAK \genblk1[7].rrel ( .Q(L[7]), .E(ren));
Q_REGFORCE \genblk1[7].rfrc ( .Q(L[7]), .A(V[7]), .E(fen));
Q_RELEASE_WEAK \genblk1[6].rrel ( .Q(L[6]), .E(ren));
Q_REGFORCE \genblk1[6].rfrc ( .Q(L[6]), .A(V[6]), .E(fen));
Q_RELEASE_WEAK \genblk1[5].rrel ( .Q(L[5]), .E(ren));
Q_REGFORCE \genblk1[5].rfrc ( .Q(L[5]), .A(V[5]), .E(fen));
Q_RELEASE_WEAK \genblk1[4].rrel ( .Q(L[4]), .E(ren));
Q_REGFORCE \genblk1[4].rfrc ( .Q(L[4]), .A(V[4]), .E(fen));
Q_RELEASE_WEAK \genblk1[3].rrel ( .Q(L[3]), .E(ren));
Q_REGFORCE \genblk1[3].rfrc ( .Q(L[3]), .A(V[3]), .E(fen));
Q_RELEASE_WEAK \genblk1[2].rrel ( .Q(L[2]), .E(ren));
Q_REGFORCE \genblk1[2].rfrc ( .Q(L[2]), .A(V[2]), .E(fen));
Q_RELEASE_WEAK \genblk1[1].rrel ( .Q(L[1]), .E(ren));
Q_REGFORCE \genblk1[1].rfrc ( .Q(L[1]), .A(V[1]), .E(fen));
Q_RELEASE_WEAK \genblk1[0].rrel ( .Q(L[0]), .E(ren));
Q_REGFORCE \genblk1[0].rfrc ( .Q(L[0]), .A(V[0]), .E(fen));
Q_AN02 U2049 ( .A0(_zzenr), .A1(n4), .Z(ren));
Q_INV U2050 ( .A(en), .Z(n4));
Q_AN02 U2051 ( .A0(n3), .A1(en), .Z(fen));
Q_INV U2052 ( .A(_zzenr), .Z(n3));
Q_FDP0UA U2053 ( .D(n5), .QTFCLK( ), .Q(_zzenr));
Q_XOR2 U2054 ( .A0(xc_top.hotSwapOnPI), .A1(en), .Z(n5));
// pragma CVASTRPROP MODULE HDLICE CVAIUSNAMES_FORGEN_LABEL "genblk1"
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE "ixc_rforce"
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE_LIB "ixcom_temp_library"
// pragma CVASTRPROP MODULE HDLICE PROP_IXCOM_MOD TRUE
endmodule
