library ieee, quickturn ;
use ieee.std_logic_1164.all ;
use quickturn.verilog.all ;
entity IXC_GFIFO is
  attribute _2_state_: integer;
  attribute upf_always_on : integer;
  attribute upf_always_on of IXC_GFIFO: entity is 1 ;
  attribute _2_state_ of IXC_GFIFO: entity is 1 ;
end IXC_GFIFO ;
