
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module cr_kme_kop_kdf_stream_pipe_xcm79 ( pipe_valid, pipe_data, 
	pipe_byte_count, clk, rst_n, cmd_valid, cmd_data_size, cmd_data, 
	pipe_ack, pipe_ack_num_bytes);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output [0:0] pipe_valid;
output [127:0] pipe_data;
output [5:0] pipe_byte_count;
input clk;
input rst_n;
input cmd_valid;
input [5:0] cmd_data_size;
input [295:0] cmd_data;
input [0:0] pipe_ack;
input [4:0] pipe_ack_num_bytes;
wire [0:5] _zy_simnet_pipe_byte_count_0_w$;
wire [295:0] cmd_data_q;
Q_ND02 U0 ( .A0(pipe_valid[0]), .A1(pipe_ack[0]), .Z(n2));
Q_INV U1 ( .A(cmd_valid), .Z(n1));
Q_AN02 U2 ( .A0(n1), .A1(n2), .Z(n3));
Q_MX02 U3 ( .S(cmd_valid), .A0(n306), .A1(cmd_data_size[5]), .Z(n4));
Q_MX02 U4 ( .S(cmd_valid), .A0(n308), .A1(cmd_data_size[4]), .Z(n5));
Q_MX02 U5 ( .S(cmd_valid), .A0(n309), .A1(cmd_data_size[3]), .Z(n6));
Q_MX02 U6 ( .S(cmd_valid), .A0(n311), .A1(cmd_data_size[2]), .Z(n7));
Q_MX02 U7 ( .S(cmd_valid), .A0(n312), .A1(cmd_data_size[1]), .Z(n8));
Q_MX02 U8 ( .S(cmd_valid), .A0(n314), .A1(cmd_data_size[0]), .Z(n9));
Q_MX02 U9 ( .S(cmd_valid), .A0(n611), .A1(cmd_data[295]), .Z(n10));
Q_MX02 U10 ( .S(cmd_valid), .A0(n610), .A1(cmd_data[294]), .Z(n11));
Q_MX02 U11 ( .S(cmd_valid), .A0(n609), .A1(cmd_data[293]), .Z(n12));
Q_MX02 U12 ( .S(cmd_valid), .A0(n608), .A1(cmd_data[292]), .Z(n13));
Q_MX02 U13 ( .S(cmd_valid), .A0(n607), .A1(cmd_data[291]), .Z(n14));
Q_MX02 U14 ( .S(cmd_valid), .A0(n606), .A1(cmd_data[290]), .Z(n15));
Q_MX02 U15 ( .S(cmd_valid), .A0(n605), .A1(cmd_data[289]), .Z(n16));
Q_MX02 U16 ( .S(cmd_valid), .A0(n604), .A1(cmd_data[288]), .Z(n17));
Q_MX02 U17 ( .S(cmd_valid), .A0(n603), .A1(cmd_data[287]), .Z(n18));
Q_MX02 U18 ( .S(cmd_valid), .A0(n602), .A1(cmd_data[286]), .Z(n19));
Q_MX02 U19 ( .S(cmd_valid), .A0(n601), .A1(cmd_data[285]), .Z(n20));
Q_MX02 U20 ( .S(cmd_valid), .A0(n600), .A1(cmd_data[284]), .Z(n21));
Q_MX02 U21 ( .S(cmd_valid), .A0(n599), .A1(cmd_data[283]), .Z(n22));
Q_MX02 U22 ( .S(cmd_valid), .A0(n598), .A1(cmd_data[282]), .Z(n23));
Q_MX02 U23 ( .S(cmd_valid), .A0(n597), .A1(cmd_data[281]), .Z(n24));
Q_MX02 U24 ( .S(cmd_valid), .A0(n596), .A1(cmd_data[280]), .Z(n25));
Q_MX02 U25 ( .S(cmd_valid), .A0(n595), .A1(cmd_data[279]), .Z(n26));
Q_MX02 U26 ( .S(cmd_valid), .A0(n594), .A1(cmd_data[278]), .Z(n27));
Q_MX02 U27 ( .S(cmd_valid), .A0(n593), .A1(cmd_data[277]), .Z(n28));
Q_MX02 U28 ( .S(cmd_valid), .A0(n592), .A1(cmd_data[276]), .Z(n29));
Q_MX02 U29 ( .S(cmd_valid), .A0(n591), .A1(cmd_data[275]), .Z(n30));
Q_MX02 U30 ( .S(cmd_valid), .A0(n590), .A1(cmd_data[274]), .Z(n31));
Q_MX02 U31 ( .S(cmd_valid), .A0(n589), .A1(cmd_data[273]), .Z(n32));
Q_MX02 U32 ( .S(cmd_valid), .A0(n588), .A1(cmd_data[272]), .Z(n33));
Q_MX02 U33 ( .S(cmd_valid), .A0(n587), .A1(cmd_data[271]), .Z(n34));
Q_MX02 U34 ( .S(cmd_valid), .A0(n586), .A1(cmd_data[270]), .Z(n35));
Q_MX02 U35 ( .S(cmd_valid), .A0(n585), .A1(cmd_data[269]), .Z(n36));
Q_MX02 U36 ( .S(cmd_valid), .A0(n584), .A1(cmd_data[268]), .Z(n37));
Q_MX02 U37 ( .S(cmd_valid), .A0(n583), .A1(cmd_data[267]), .Z(n38));
Q_MX02 U38 ( .S(cmd_valid), .A0(n582), .A1(cmd_data[266]), .Z(n39));
Q_MX02 U39 ( .S(cmd_valid), .A0(n581), .A1(cmd_data[265]), .Z(n40));
Q_MX02 U40 ( .S(cmd_valid), .A0(n580), .A1(cmd_data[264]), .Z(n41));
Q_MX02 U41 ( .S(cmd_valid), .A0(n579), .A1(cmd_data[263]), .Z(n42));
Q_MX02 U42 ( .S(cmd_valid), .A0(n578), .A1(cmd_data[262]), .Z(n43));
Q_MX02 U43 ( .S(cmd_valid), .A0(n577), .A1(cmd_data[261]), .Z(n44));
Q_MX02 U44 ( .S(cmd_valid), .A0(n576), .A1(cmd_data[260]), .Z(n45));
Q_MX02 U45 ( .S(cmd_valid), .A0(n575), .A1(cmd_data[259]), .Z(n46));
Q_MX02 U46 ( .S(cmd_valid), .A0(n574), .A1(cmd_data[258]), .Z(n47));
Q_MX02 U47 ( .S(cmd_valid), .A0(n573), .A1(cmd_data[257]), .Z(n48));
Q_MX02 U48 ( .S(cmd_valid), .A0(n572), .A1(cmd_data[256]), .Z(n49));
Q_MX02 U49 ( .S(cmd_valid), .A0(n571), .A1(cmd_data[255]), .Z(n50));
Q_MX02 U50 ( .S(cmd_valid), .A0(n570), .A1(cmd_data[254]), .Z(n51));
Q_MX02 U51 ( .S(cmd_valid), .A0(n569), .A1(cmd_data[253]), .Z(n52));
Q_MX02 U52 ( .S(cmd_valid), .A0(n568), .A1(cmd_data[252]), .Z(n53));
Q_MX02 U53 ( .S(cmd_valid), .A0(n567), .A1(cmd_data[251]), .Z(n54));
Q_MX02 U54 ( .S(cmd_valid), .A0(n566), .A1(cmd_data[250]), .Z(n55));
Q_MX02 U55 ( .S(cmd_valid), .A0(n565), .A1(cmd_data[249]), .Z(n56));
Q_MX02 U56 ( .S(cmd_valid), .A0(n564), .A1(cmd_data[248]), .Z(n57));
Q_MX02 U57 ( .S(cmd_valid), .A0(n563), .A1(cmd_data[247]), .Z(n58));
Q_MX02 U58 ( .S(cmd_valid), .A0(n562), .A1(cmd_data[246]), .Z(n59));
Q_MX02 U59 ( .S(cmd_valid), .A0(n561), .A1(cmd_data[245]), .Z(n60));
Q_MX02 U60 ( .S(cmd_valid), .A0(n560), .A1(cmd_data[244]), .Z(n61));
Q_MX02 U61 ( .S(cmd_valid), .A0(n559), .A1(cmd_data[243]), .Z(n62));
Q_MX02 U62 ( .S(cmd_valid), .A0(n558), .A1(cmd_data[242]), .Z(n63));
Q_MX02 U63 ( .S(cmd_valid), .A0(n557), .A1(cmd_data[241]), .Z(n64));
Q_MX02 U64 ( .S(cmd_valid), .A0(n556), .A1(cmd_data[240]), .Z(n65));
Q_MX02 U65 ( .S(cmd_valid), .A0(n555), .A1(cmd_data[239]), .Z(n66));
Q_MX02 U66 ( .S(cmd_valid), .A0(n554), .A1(cmd_data[238]), .Z(n67));
Q_MX02 U67 ( .S(cmd_valid), .A0(n553), .A1(cmd_data[237]), .Z(n68));
Q_MX02 U68 ( .S(cmd_valid), .A0(n552), .A1(cmd_data[236]), .Z(n69));
Q_MX02 U69 ( .S(cmd_valid), .A0(n551), .A1(cmd_data[235]), .Z(n70));
Q_MX02 U70 ( .S(cmd_valid), .A0(n550), .A1(cmd_data[234]), .Z(n71));
Q_MX02 U71 ( .S(cmd_valid), .A0(n549), .A1(cmd_data[233]), .Z(n72));
Q_MX02 U72 ( .S(cmd_valid), .A0(n548), .A1(cmd_data[232]), .Z(n73));
Q_MX02 U73 ( .S(cmd_valid), .A0(n547), .A1(cmd_data[231]), .Z(n74));
Q_MX02 U74 ( .S(cmd_valid), .A0(n546), .A1(cmd_data[230]), .Z(n75));
Q_MX02 U75 ( .S(cmd_valid), .A0(n545), .A1(cmd_data[229]), .Z(n76));
Q_MX02 U76 ( .S(cmd_valid), .A0(n544), .A1(cmd_data[228]), .Z(n77));
Q_MX02 U77 ( .S(cmd_valid), .A0(n543), .A1(cmd_data[227]), .Z(n78));
Q_MX02 U78 ( .S(cmd_valid), .A0(n542), .A1(cmd_data[226]), .Z(n79));
Q_MX02 U79 ( .S(cmd_valid), .A0(n541), .A1(cmd_data[225]), .Z(n80));
Q_MX02 U80 ( .S(cmd_valid), .A0(n540), .A1(cmd_data[224]), .Z(n81));
Q_MX02 U81 ( .S(cmd_valid), .A0(n539), .A1(cmd_data[223]), .Z(n82));
Q_MX02 U82 ( .S(cmd_valid), .A0(n538), .A1(cmd_data[222]), .Z(n83));
Q_MX02 U83 ( .S(cmd_valid), .A0(n537), .A1(cmd_data[221]), .Z(n84));
Q_MX02 U84 ( .S(cmd_valid), .A0(n536), .A1(cmd_data[220]), .Z(n85));
Q_MX02 U85 ( .S(cmd_valid), .A0(n535), .A1(cmd_data[219]), .Z(n86));
Q_MX02 U86 ( .S(cmd_valid), .A0(n534), .A1(cmd_data[218]), .Z(n87));
Q_MX02 U87 ( .S(cmd_valid), .A0(n533), .A1(cmd_data[217]), .Z(n88));
Q_MX02 U88 ( .S(cmd_valid), .A0(n532), .A1(cmd_data[216]), .Z(n89));
Q_MX02 U89 ( .S(cmd_valid), .A0(n531), .A1(cmd_data[215]), .Z(n90));
Q_MX02 U90 ( .S(cmd_valid), .A0(n530), .A1(cmd_data[214]), .Z(n91));
Q_MX02 U91 ( .S(cmd_valid), .A0(n529), .A1(cmd_data[213]), .Z(n92));
Q_MX02 U92 ( .S(cmd_valid), .A0(n528), .A1(cmd_data[212]), .Z(n93));
Q_MX02 U93 ( .S(cmd_valid), .A0(n527), .A1(cmd_data[211]), .Z(n94));
Q_MX02 U94 ( .S(cmd_valid), .A0(n526), .A1(cmd_data[210]), .Z(n95));
Q_MX02 U95 ( .S(cmd_valid), .A0(n525), .A1(cmd_data[209]), .Z(n96));
Q_MX02 U96 ( .S(cmd_valid), .A0(n524), .A1(cmd_data[208]), .Z(n97));
Q_MX02 U97 ( .S(cmd_valid), .A0(n523), .A1(cmd_data[207]), .Z(n98));
Q_MX02 U98 ( .S(cmd_valid), .A0(n522), .A1(cmd_data[206]), .Z(n99));
Q_MX02 U99 ( .S(cmd_valid), .A0(n521), .A1(cmd_data[205]), .Z(n100));
Q_MX02 U100 ( .S(cmd_valid), .A0(n520), .A1(cmd_data[204]), .Z(n101));
Q_MX02 U101 ( .S(cmd_valid), .A0(n519), .A1(cmd_data[203]), .Z(n102));
Q_MX02 U102 ( .S(cmd_valid), .A0(n518), .A1(cmd_data[202]), .Z(n103));
Q_MX02 U103 ( .S(cmd_valid), .A0(n517), .A1(cmd_data[201]), .Z(n104));
Q_MX02 U104 ( .S(cmd_valid), .A0(n516), .A1(cmd_data[200]), .Z(n105));
Q_MX02 U105 ( .S(cmd_valid), .A0(n515), .A1(cmd_data[199]), .Z(n106));
Q_MX02 U106 ( .S(cmd_valid), .A0(n514), .A1(cmd_data[198]), .Z(n107));
Q_MX02 U107 ( .S(cmd_valid), .A0(n513), .A1(cmd_data[197]), .Z(n108));
Q_MX02 U108 ( .S(cmd_valid), .A0(n512), .A1(cmd_data[196]), .Z(n109));
Q_MX02 U109 ( .S(cmd_valid), .A0(n511), .A1(cmd_data[195]), .Z(n110));
Q_MX02 U110 ( .S(cmd_valid), .A0(n510), .A1(cmd_data[194]), .Z(n111));
Q_MX02 U111 ( .S(cmd_valid), .A0(n509), .A1(cmd_data[193]), .Z(n112));
Q_MX02 U112 ( .S(cmd_valid), .A0(n508), .A1(cmd_data[192]), .Z(n113));
Q_MX02 U113 ( .S(cmd_valid), .A0(n507), .A1(cmd_data[191]), .Z(n114));
Q_MX02 U114 ( .S(cmd_valid), .A0(n506), .A1(cmd_data[190]), .Z(n115));
Q_MX02 U115 ( .S(cmd_valid), .A0(n505), .A1(cmd_data[189]), .Z(n116));
Q_MX02 U116 ( .S(cmd_valid), .A0(n504), .A1(cmd_data[188]), .Z(n117));
Q_MX02 U117 ( .S(cmd_valid), .A0(n503), .A1(cmd_data[187]), .Z(n118));
Q_MX02 U118 ( .S(cmd_valid), .A0(n502), .A1(cmd_data[186]), .Z(n119));
Q_MX02 U119 ( .S(cmd_valid), .A0(n501), .A1(cmd_data[185]), .Z(n120));
Q_MX02 U120 ( .S(cmd_valid), .A0(n500), .A1(cmd_data[184]), .Z(n121));
Q_MX02 U121 ( .S(cmd_valid), .A0(n499), .A1(cmd_data[183]), .Z(n122));
Q_MX02 U122 ( .S(cmd_valid), .A0(n498), .A1(cmd_data[182]), .Z(n123));
Q_MX02 U123 ( .S(cmd_valid), .A0(n497), .A1(cmd_data[181]), .Z(n124));
Q_MX02 U124 ( .S(cmd_valid), .A0(n496), .A1(cmd_data[180]), .Z(n125));
Q_MX02 U125 ( .S(cmd_valid), .A0(n495), .A1(cmd_data[179]), .Z(n126));
Q_MX02 U126 ( .S(cmd_valid), .A0(n494), .A1(cmd_data[178]), .Z(n127));
Q_MX02 U127 ( .S(cmd_valid), .A0(n493), .A1(cmd_data[177]), .Z(n128));
Q_MX02 U128 ( .S(cmd_valid), .A0(n492), .A1(cmd_data[176]), .Z(n129));
Q_MX02 U129 ( .S(cmd_valid), .A0(n491), .A1(cmd_data[175]), .Z(n130));
Q_MX02 U130 ( .S(cmd_valid), .A0(n490), .A1(cmd_data[174]), .Z(n131));
Q_MX02 U131 ( .S(cmd_valid), .A0(n489), .A1(cmd_data[173]), .Z(n132));
Q_MX02 U132 ( .S(cmd_valid), .A0(n488), .A1(cmd_data[172]), .Z(n133));
Q_MX02 U133 ( .S(cmd_valid), .A0(n487), .A1(cmd_data[171]), .Z(n134));
Q_MX02 U134 ( .S(cmd_valid), .A0(n486), .A1(cmd_data[170]), .Z(n135));
Q_MX02 U135 ( .S(cmd_valid), .A0(n485), .A1(cmd_data[169]), .Z(n136));
Q_MX02 U136 ( .S(cmd_valid), .A0(n484), .A1(cmd_data[168]), .Z(n137));
Q_MX02 U137 ( .S(cmd_valid), .A0(n483), .A1(cmd_data[167]), .Z(n138));
Q_MX02 U138 ( .S(cmd_valid), .A0(n482), .A1(cmd_data[166]), .Z(n139));
Q_MX02 U139 ( .S(cmd_valid), .A0(n481), .A1(cmd_data[165]), .Z(n140));
Q_MX02 U140 ( .S(cmd_valid), .A0(n480), .A1(cmd_data[164]), .Z(n141));
Q_MX02 U141 ( .S(cmd_valid), .A0(n479), .A1(cmd_data[163]), .Z(n142));
Q_MX02 U142 ( .S(cmd_valid), .A0(n478), .A1(cmd_data[162]), .Z(n143));
Q_MX02 U143 ( .S(cmd_valid), .A0(n477), .A1(cmd_data[161]), .Z(n144));
Q_MX02 U144 ( .S(cmd_valid), .A0(n476), .A1(cmd_data[160]), .Z(n145));
Q_MX02 U145 ( .S(cmd_valid), .A0(n475), .A1(cmd_data[159]), .Z(n146));
Q_MX02 U146 ( .S(cmd_valid), .A0(n474), .A1(cmd_data[158]), .Z(n147));
Q_MX02 U147 ( .S(cmd_valid), .A0(n473), .A1(cmd_data[157]), .Z(n148));
Q_MX02 U148 ( .S(cmd_valid), .A0(n472), .A1(cmd_data[156]), .Z(n149));
Q_MX02 U149 ( .S(cmd_valid), .A0(n471), .A1(cmd_data[155]), .Z(n150));
Q_MX02 U150 ( .S(cmd_valid), .A0(n470), .A1(cmd_data[154]), .Z(n151));
Q_MX02 U151 ( .S(cmd_valid), .A0(n469), .A1(cmd_data[153]), .Z(n152));
Q_MX02 U152 ( .S(cmd_valid), .A0(n468), .A1(cmd_data[152]), .Z(n153));
Q_MX02 U153 ( .S(cmd_valid), .A0(n467), .A1(cmd_data[151]), .Z(n154));
Q_MX02 U154 ( .S(cmd_valid), .A0(n466), .A1(cmd_data[150]), .Z(n155));
Q_MX02 U155 ( .S(cmd_valid), .A0(n465), .A1(cmd_data[149]), .Z(n156));
Q_MX02 U156 ( .S(cmd_valid), .A0(n464), .A1(cmd_data[148]), .Z(n157));
Q_MX02 U157 ( .S(cmd_valid), .A0(n463), .A1(cmd_data[147]), .Z(n158));
Q_MX02 U158 ( .S(cmd_valid), .A0(n462), .A1(cmd_data[146]), .Z(n159));
Q_MX02 U159 ( .S(cmd_valid), .A0(n461), .A1(cmd_data[145]), .Z(n160));
Q_MX02 U160 ( .S(cmd_valid), .A0(n460), .A1(cmd_data[144]), .Z(n161));
Q_MX02 U161 ( .S(cmd_valid), .A0(n459), .A1(cmd_data[143]), .Z(n162));
Q_MX02 U162 ( .S(cmd_valid), .A0(n458), .A1(cmd_data[142]), .Z(n163));
Q_MX02 U163 ( .S(cmd_valid), .A0(n457), .A1(cmd_data[141]), .Z(n164));
Q_MX02 U164 ( .S(cmd_valid), .A0(n456), .A1(cmd_data[140]), .Z(n165));
Q_MX02 U165 ( .S(cmd_valid), .A0(n455), .A1(cmd_data[139]), .Z(n166));
Q_MX02 U166 ( .S(cmd_valid), .A0(n454), .A1(cmd_data[138]), .Z(n167));
Q_MX02 U167 ( .S(cmd_valid), .A0(n453), .A1(cmd_data[137]), .Z(n168));
Q_MX02 U168 ( .S(cmd_valid), .A0(n452), .A1(cmd_data[136]), .Z(n169));
Q_MX02 U169 ( .S(cmd_valid), .A0(n451), .A1(cmd_data[135]), .Z(n170));
Q_MX02 U170 ( .S(cmd_valid), .A0(n450), .A1(cmd_data[134]), .Z(n171));
Q_MX02 U171 ( .S(cmd_valid), .A0(n449), .A1(cmd_data[133]), .Z(n172));
Q_MX02 U172 ( .S(cmd_valid), .A0(n448), .A1(cmd_data[132]), .Z(n173));
Q_MX02 U173 ( .S(cmd_valid), .A0(n447), .A1(cmd_data[131]), .Z(n174));
Q_MX02 U174 ( .S(cmd_valid), .A0(n446), .A1(cmd_data[130]), .Z(n175));
Q_MX02 U175 ( .S(cmd_valid), .A0(n445), .A1(cmd_data[129]), .Z(n176));
Q_MX02 U176 ( .S(cmd_valid), .A0(n444), .A1(cmd_data[128]), .Z(n177));
Q_MX02 U177 ( .S(cmd_valid), .A0(n442), .A1(cmd_data[127]), .Z(n178));
Q_MX02 U178 ( .S(cmd_valid), .A0(n441), .A1(cmd_data[126]), .Z(n179));
Q_MX02 U179 ( .S(cmd_valid), .A0(n440), .A1(cmd_data[125]), .Z(n180));
Q_MX02 U180 ( .S(cmd_valid), .A0(n439), .A1(cmd_data[124]), .Z(n181));
Q_MX02 U181 ( .S(cmd_valid), .A0(n438), .A1(cmd_data[123]), .Z(n182));
Q_MX02 U182 ( .S(cmd_valid), .A0(n437), .A1(cmd_data[122]), .Z(n183));
Q_MX02 U183 ( .S(cmd_valid), .A0(n436), .A1(cmd_data[121]), .Z(n184));
Q_MX02 U184 ( .S(cmd_valid), .A0(n435), .A1(cmd_data[120]), .Z(n185));
Q_MX02 U185 ( .S(cmd_valid), .A0(n434), .A1(cmd_data[119]), .Z(n186));
Q_MX02 U186 ( .S(cmd_valid), .A0(n433), .A1(cmd_data[118]), .Z(n187));
Q_MX02 U187 ( .S(cmd_valid), .A0(n432), .A1(cmd_data[117]), .Z(n188));
Q_MX02 U188 ( .S(cmd_valid), .A0(n431), .A1(cmd_data[116]), .Z(n189));
Q_MX02 U189 ( .S(cmd_valid), .A0(n430), .A1(cmd_data[115]), .Z(n190));
Q_MX02 U190 ( .S(cmd_valid), .A0(n429), .A1(cmd_data[114]), .Z(n191));
Q_MX02 U191 ( .S(cmd_valid), .A0(n428), .A1(cmd_data[113]), .Z(n192));
Q_MX02 U192 ( .S(cmd_valid), .A0(n427), .A1(cmd_data[112]), .Z(n193));
Q_MX02 U193 ( .S(cmd_valid), .A0(n426), .A1(cmd_data[111]), .Z(n194));
Q_MX02 U194 ( .S(cmd_valid), .A0(n425), .A1(cmd_data[110]), .Z(n195));
Q_MX02 U195 ( .S(cmd_valid), .A0(n424), .A1(cmd_data[109]), .Z(n196));
Q_MX02 U196 ( .S(cmd_valid), .A0(n423), .A1(cmd_data[108]), .Z(n197));
Q_MX02 U197 ( .S(cmd_valid), .A0(n422), .A1(cmd_data[107]), .Z(n198));
Q_MX02 U198 ( .S(cmd_valid), .A0(n421), .A1(cmd_data[106]), .Z(n199));
Q_MX02 U199 ( .S(cmd_valid), .A0(n420), .A1(cmd_data[105]), .Z(n200));
Q_MX02 U200 ( .S(cmd_valid), .A0(n419), .A1(cmd_data[104]), .Z(n201));
Q_MX02 U201 ( .S(cmd_valid), .A0(n418), .A1(cmd_data[103]), .Z(n202));
Q_MX02 U202 ( .S(cmd_valid), .A0(n417), .A1(cmd_data[102]), .Z(n203));
Q_MX02 U203 ( .S(cmd_valid), .A0(n416), .A1(cmd_data[101]), .Z(n204));
Q_MX02 U204 ( .S(cmd_valid), .A0(n415), .A1(cmd_data[100]), .Z(n205));
Q_MX02 U205 ( .S(cmd_valid), .A0(n414), .A1(cmd_data[99]), .Z(n206));
Q_MX02 U206 ( .S(cmd_valid), .A0(n413), .A1(cmd_data[98]), .Z(n207));
Q_MX02 U207 ( .S(cmd_valid), .A0(n412), .A1(cmd_data[97]), .Z(n208));
Q_MX02 U208 ( .S(cmd_valid), .A0(n411), .A1(cmd_data[96]), .Z(n209));
Q_MX02 U209 ( .S(cmd_valid), .A0(n410), .A1(cmd_data[95]), .Z(n210));
Q_MX02 U210 ( .S(cmd_valid), .A0(n409), .A1(cmd_data[94]), .Z(n211));
Q_MX02 U211 ( .S(cmd_valid), .A0(n408), .A1(cmd_data[93]), .Z(n212));
Q_MX02 U212 ( .S(cmd_valid), .A0(n407), .A1(cmd_data[92]), .Z(n213));
Q_MX02 U213 ( .S(cmd_valid), .A0(n406), .A1(cmd_data[91]), .Z(n214));
Q_MX02 U214 ( .S(cmd_valid), .A0(n405), .A1(cmd_data[90]), .Z(n215));
Q_MX02 U215 ( .S(cmd_valid), .A0(n404), .A1(cmd_data[89]), .Z(n216));
Q_MX02 U216 ( .S(cmd_valid), .A0(n403), .A1(cmd_data[88]), .Z(n217));
Q_MX02 U217 ( .S(cmd_valid), .A0(n402), .A1(cmd_data[87]), .Z(n218));
Q_MX02 U218 ( .S(cmd_valid), .A0(n401), .A1(cmd_data[86]), .Z(n219));
Q_MX02 U219 ( .S(cmd_valid), .A0(n400), .A1(cmd_data[85]), .Z(n220));
Q_MX02 U220 ( .S(cmd_valid), .A0(n399), .A1(cmd_data[84]), .Z(n221));
Q_MX02 U221 ( .S(cmd_valid), .A0(n398), .A1(cmd_data[83]), .Z(n222));
Q_MX02 U222 ( .S(cmd_valid), .A0(n397), .A1(cmd_data[82]), .Z(n223));
Q_MX02 U223 ( .S(cmd_valid), .A0(n396), .A1(cmd_data[81]), .Z(n224));
Q_MX02 U224 ( .S(cmd_valid), .A0(n395), .A1(cmd_data[80]), .Z(n225));
Q_MX02 U225 ( .S(cmd_valid), .A0(n394), .A1(cmd_data[79]), .Z(n226));
Q_MX02 U226 ( .S(cmd_valid), .A0(n393), .A1(cmd_data[78]), .Z(n227));
Q_MX02 U227 ( .S(cmd_valid), .A0(n392), .A1(cmd_data[77]), .Z(n228));
Q_MX02 U228 ( .S(cmd_valid), .A0(n391), .A1(cmd_data[76]), .Z(n229));
Q_MX02 U229 ( .S(cmd_valid), .A0(n390), .A1(cmd_data[75]), .Z(n230));
Q_MX02 U230 ( .S(cmd_valid), .A0(n389), .A1(cmd_data[74]), .Z(n231));
Q_MX02 U231 ( .S(cmd_valid), .A0(n388), .A1(cmd_data[73]), .Z(n232));
Q_MX02 U232 ( .S(cmd_valid), .A0(n387), .A1(cmd_data[72]), .Z(n233));
Q_MX02 U233 ( .S(cmd_valid), .A0(n386), .A1(cmd_data[71]), .Z(n234));
Q_MX02 U234 ( .S(cmd_valid), .A0(n385), .A1(cmd_data[70]), .Z(n235));
Q_MX02 U235 ( .S(cmd_valid), .A0(n384), .A1(cmd_data[69]), .Z(n236));
Q_MX02 U236 ( .S(cmd_valid), .A0(n383), .A1(cmd_data[68]), .Z(n237));
Q_MX02 U237 ( .S(cmd_valid), .A0(n382), .A1(cmd_data[67]), .Z(n238));
Q_MX02 U238 ( .S(cmd_valid), .A0(n381), .A1(cmd_data[66]), .Z(n239));
Q_MX02 U239 ( .S(cmd_valid), .A0(n380), .A1(cmd_data[65]), .Z(n240));
Q_MX02 U240 ( .S(cmd_valid), .A0(n379), .A1(cmd_data[64]), .Z(n241));
Q_MX02 U241 ( .S(cmd_valid), .A0(n378), .A1(cmd_data[63]), .Z(n242));
Q_MX02 U242 ( .S(cmd_valid), .A0(n377), .A1(cmd_data[62]), .Z(n243));
Q_MX02 U243 ( .S(cmd_valid), .A0(n376), .A1(cmd_data[61]), .Z(n244));
Q_MX02 U244 ( .S(cmd_valid), .A0(n375), .A1(cmd_data[60]), .Z(n245));
Q_MX02 U245 ( .S(cmd_valid), .A0(n374), .A1(cmd_data[59]), .Z(n246));
Q_MX02 U246 ( .S(cmd_valid), .A0(n373), .A1(cmd_data[58]), .Z(n247));
Q_MX02 U247 ( .S(cmd_valid), .A0(n372), .A1(cmd_data[57]), .Z(n248));
Q_MX02 U248 ( .S(cmd_valid), .A0(n371), .A1(cmd_data[56]), .Z(n249));
Q_MX02 U249 ( .S(cmd_valid), .A0(n370), .A1(cmd_data[55]), .Z(n250));
Q_MX02 U250 ( .S(cmd_valid), .A0(n369), .A1(cmd_data[54]), .Z(n251));
Q_MX02 U251 ( .S(cmd_valid), .A0(n368), .A1(cmd_data[53]), .Z(n252));
Q_MX02 U252 ( .S(cmd_valid), .A0(n367), .A1(cmd_data[52]), .Z(n253));
Q_MX02 U253 ( .S(cmd_valid), .A0(n366), .A1(cmd_data[51]), .Z(n254));
Q_MX02 U254 ( .S(cmd_valid), .A0(n365), .A1(cmd_data[50]), .Z(n255));
Q_MX02 U255 ( .S(cmd_valid), .A0(n364), .A1(cmd_data[49]), .Z(n256));
Q_MX02 U256 ( .S(cmd_valid), .A0(n363), .A1(cmd_data[48]), .Z(n257));
Q_MX02 U257 ( .S(cmd_valid), .A0(n362), .A1(cmd_data[47]), .Z(n258));
Q_MX02 U258 ( .S(cmd_valid), .A0(n361), .A1(cmd_data[46]), .Z(n259));
Q_MX02 U259 ( .S(cmd_valid), .A0(n360), .A1(cmd_data[45]), .Z(n260));
Q_MX02 U260 ( .S(cmd_valid), .A0(n359), .A1(cmd_data[44]), .Z(n261));
Q_MX02 U261 ( .S(cmd_valid), .A0(n358), .A1(cmd_data[43]), .Z(n262));
Q_MX02 U262 ( .S(cmd_valid), .A0(n357), .A1(cmd_data[42]), .Z(n263));
Q_MX02 U263 ( .S(cmd_valid), .A0(n356), .A1(cmd_data[41]), .Z(n264));
Q_MX02 U264 ( .S(cmd_valid), .A0(n355), .A1(cmd_data[40]), .Z(n265));
Q_MX02 U265 ( .S(cmd_valid), .A0(n354), .A1(cmd_data[39]), .Z(n266));
Q_MX02 U266 ( .S(cmd_valid), .A0(n353), .A1(cmd_data[38]), .Z(n267));
Q_MX02 U267 ( .S(cmd_valid), .A0(n352), .A1(cmd_data[37]), .Z(n268));
Q_MX02 U268 ( .S(cmd_valid), .A0(n351), .A1(cmd_data[36]), .Z(n269));
Q_MX02 U269 ( .S(cmd_valid), .A0(n350), .A1(cmd_data[35]), .Z(n270));
Q_MX02 U270 ( .S(cmd_valid), .A0(n349), .A1(cmd_data[34]), .Z(n271));
Q_MX02 U271 ( .S(cmd_valid), .A0(n348), .A1(cmd_data[33]), .Z(n272));
Q_MX02 U272 ( .S(cmd_valid), .A0(n347), .A1(cmd_data[32]), .Z(n273));
Q_MX02 U273 ( .S(cmd_valid), .A0(n346), .A1(cmd_data[31]), .Z(n274));
Q_MX02 U274 ( .S(cmd_valid), .A0(n345), .A1(cmd_data[30]), .Z(n275));
Q_MX02 U275 ( .S(cmd_valid), .A0(n344), .A1(cmd_data[29]), .Z(n276));
Q_MX02 U276 ( .S(cmd_valid), .A0(n343), .A1(cmd_data[28]), .Z(n277));
Q_MX02 U277 ( .S(cmd_valid), .A0(n342), .A1(cmd_data[27]), .Z(n278));
Q_MX02 U278 ( .S(cmd_valid), .A0(n341), .A1(cmd_data[26]), .Z(n279));
Q_MX02 U279 ( .S(cmd_valid), .A0(n340), .A1(cmd_data[25]), .Z(n280));
Q_MX02 U280 ( .S(cmd_valid), .A0(n339), .A1(cmd_data[24]), .Z(n281));
Q_MX02 U281 ( .S(cmd_valid), .A0(n338), .A1(cmd_data[23]), .Z(n282));
Q_MX02 U282 ( .S(cmd_valid), .A0(n337), .A1(cmd_data[22]), .Z(n283));
Q_MX02 U283 ( .S(cmd_valid), .A0(n336), .A1(cmd_data[21]), .Z(n284));
Q_MX02 U284 ( .S(cmd_valid), .A0(n335), .A1(cmd_data[20]), .Z(n285));
Q_MX02 U285 ( .S(cmd_valid), .A0(n334), .A1(cmd_data[19]), .Z(n286));
Q_MX02 U286 ( .S(cmd_valid), .A0(n333), .A1(cmd_data[18]), .Z(n287));
Q_MX02 U287 ( .S(cmd_valid), .A0(n332), .A1(cmd_data[17]), .Z(n288));
Q_MX02 U288 ( .S(cmd_valid), .A0(n331), .A1(cmd_data[16]), .Z(n289));
Q_MX02 U289 ( .S(cmd_valid), .A0(n330), .A1(cmd_data[15]), .Z(n290));
Q_MX02 U290 ( .S(cmd_valid), .A0(n329), .A1(cmd_data[14]), .Z(n291));
Q_MX02 U291 ( .S(cmd_valid), .A0(n328), .A1(cmd_data[13]), .Z(n292));
Q_MX02 U292 ( .S(cmd_valid), .A0(n327), .A1(cmd_data[12]), .Z(n293));
Q_MX02 U293 ( .S(cmd_valid), .A0(n326), .A1(cmd_data[11]), .Z(n294));
Q_MX02 U294 ( .S(cmd_valid), .A0(n325), .A1(cmd_data[10]), .Z(n295));
Q_MX02 U295 ( .S(cmd_valid), .A0(n324), .A1(cmd_data[9]), .Z(n296));
Q_MX02 U296 ( .S(cmd_valid), .A0(n323), .A1(cmd_data[8]), .Z(n297));
Q_MX02 U297 ( .S(cmd_valid), .A0(n322), .A1(cmd_data[7]), .Z(n298));
Q_MX02 U298 ( .S(cmd_valid), .A0(n321), .A1(cmd_data[6]), .Z(n299));
Q_MX02 U299 ( .S(cmd_valid), .A0(n320), .A1(cmd_data[5]), .Z(n300));
Q_MX02 U300 ( .S(cmd_valid), .A0(n319), .A1(cmd_data[4]), .Z(n301));
Q_MX02 U301 ( .S(cmd_valid), .A0(n318), .A1(cmd_data[3]), .Z(n302));
Q_MX02 U302 ( .S(cmd_valid), .A0(n317), .A1(cmd_data[2]), .Z(n303));
Q_MX02 U303 ( .S(cmd_valid), .A0(n316), .A1(cmd_data[1]), .Z(n304));
Q_MX02 U304 ( .S(cmd_valid), .A0(n315), .A1(cmd_data[0]), .Z(n305));
Q_XNR2 U305 ( .A0(pipe_byte_count[5]), .A1(n307), .Z(n306));
Q_AD02 U306 ( .CI(n310), .A0(pipe_byte_count[3]), .A1(pipe_byte_count[4]), .B0(n676), .B1(n443), .S0(n309), .S1(n308), .CO(n307));
Q_AD02 U307 ( .CI(n313), .A0(pipe_byte_count[1]), .A1(pipe_byte_count[2]), .B0(n1094), .B1(n813), .S0(n312), .S1(n311), .CO(n310));
Q_OR02 U308 ( .A0(pipe_byte_count[0]), .A1(n1351), .Z(n313));
Q_XNR2 U309 ( .A0(pipe_byte_count[0]), .A1(n1351), .Z(n314));
Q_AN02 U310 ( .A0(n443), .A1(n612), .Z(n315));
Q_AN02 U311 ( .A0(n443), .A1(n613), .Z(n316));
Q_AN02 U312 ( .A0(n443), .A1(n614), .Z(n317));
Q_AN02 U313 ( .A0(n443), .A1(n615), .Z(n318));
Q_AN02 U314 ( .A0(n443), .A1(n616), .Z(n319));
Q_AN02 U315 ( .A0(n443), .A1(n617), .Z(n320));
Q_AN02 U316 ( .A0(n443), .A1(n618), .Z(n321));
Q_AN02 U317 ( .A0(n443), .A1(n619), .Z(n322));
Q_AN02 U318 ( .A0(n443), .A1(n620), .Z(n323));
Q_AN02 U319 ( .A0(n443), .A1(n621), .Z(n324));
Q_AN02 U320 ( .A0(n443), .A1(n622), .Z(n325));
Q_AN02 U321 ( .A0(n443), .A1(n623), .Z(n326));
Q_AN02 U322 ( .A0(n443), .A1(n624), .Z(n327));
Q_AN02 U323 ( .A0(n443), .A1(n625), .Z(n328));
Q_AN02 U324 ( .A0(n443), .A1(n626), .Z(n329));
Q_AN02 U325 ( .A0(n443), .A1(n627), .Z(n330));
Q_AN02 U326 ( .A0(n443), .A1(n628), .Z(n331));
Q_AN02 U327 ( .A0(n443), .A1(n629), .Z(n332));
Q_AN02 U328 ( .A0(n443), .A1(n630), .Z(n333));
Q_AN02 U329 ( .A0(n443), .A1(n631), .Z(n334));
Q_AN02 U330 ( .A0(n443), .A1(n632), .Z(n335));
Q_AN02 U331 ( .A0(n443), .A1(n633), .Z(n336));
Q_AN02 U332 ( .A0(n443), .A1(n634), .Z(n337));
Q_AN02 U333 ( .A0(n443), .A1(n635), .Z(n338));
Q_AN02 U334 ( .A0(n443), .A1(n636), .Z(n339));
Q_AN02 U335 ( .A0(n443), .A1(n637), .Z(n340));
Q_AN02 U336 ( .A0(n443), .A1(n638), .Z(n341));
Q_AN02 U337 ( .A0(n443), .A1(n639), .Z(n342));
Q_AN02 U338 ( .A0(n443), .A1(n640), .Z(n343));
Q_AN02 U339 ( .A0(n443), .A1(n641), .Z(n344));
Q_AN02 U340 ( .A0(n443), .A1(n642), .Z(n345));
Q_AN02 U341 ( .A0(n443), .A1(n643), .Z(n346));
Q_AN02 U342 ( .A0(n443), .A1(n644), .Z(n347));
Q_AN02 U343 ( .A0(n443), .A1(n645), .Z(n348));
Q_AN02 U344 ( .A0(n443), .A1(n646), .Z(n349));
Q_AN02 U345 ( .A0(n443), .A1(n647), .Z(n350));
Q_AN02 U346 ( .A0(n443), .A1(n648), .Z(n351));
Q_AN02 U347 ( .A0(n443), .A1(n649), .Z(n352));
Q_AN02 U348 ( .A0(n443), .A1(n650), .Z(n353));
Q_AN02 U349 ( .A0(n443), .A1(n651), .Z(n354));
Q_AN02 U350 ( .A0(n443), .A1(n652), .Z(n355));
Q_AN02 U351 ( .A0(n443), .A1(n653), .Z(n356));
Q_AN02 U352 ( .A0(n443), .A1(n654), .Z(n357));
Q_AN02 U353 ( .A0(n443), .A1(n655), .Z(n358));
Q_AN02 U354 ( .A0(n443), .A1(n656), .Z(n359));
Q_AN02 U355 ( .A0(n443), .A1(n657), .Z(n360));
Q_AN02 U356 ( .A0(n443), .A1(n658), .Z(n361));
Q_AN02 U357 ( .A0(n443), .A1(n659), .Z(n362));
Q_AN02 U358 ( .A0(n443), .A1(n660), .Z(n363));
Q_AN02 U359 ( .A0(n443), .A1(n661), .Z(n364));
Q_AN02 U360 ( .A0(n443), .A1(n662), .Z(n365));
Q_AN02 U361 ( .A0(n443), .A1(n663), .Z(n366));
Q_AN02 U362 ( .A0(n443), .A1(n664), .Z(n367));
Q_AN02 U363 ( .A0(n443), .A1(n665), .Z(n368));
Q_AN02 U364 ( .A0(n443), .A1(n666), .Z(n369));
Q_AN02 U365 ( .A0(n443), .A1(n667), .Z(n370));
Q_AN02 U366 ( .A0(n443), .A1(n668), .Z(n371));
Q_AN02 U367 ( .A0(n443), .A1(n669), .Z(n372));
Q_AN02 U368 ( .A0(n443), .A1(n670), .Z(n373));
Q_AN02 U369 ( .A0(n443), .A1(n671), .Z(n374));
Q_AN02 U370 ( .A0(n443), .A1(n672), .Z(n375));
Q_AN02 U371 ( .A0(n443), .A1(n673), .Z(n376));
Q_AN02 U372 ( .A0(n443), .A1(n674), .Z(n377));
Q_AN02 U373 ( .A0(n443), .A1(n675), .Z(n378));
Q_AN02 U374 ( .A0(n443), .A1(n677), .Z(n379));
Q_AN02 U375 ( .A0(n443), .A1(n678), .Z(n380));
Q_AN02 U376 ( .A0(n443), .A1(n679), .Z(n381));
Q_AN02 U377 ( .A0(n443), .A1(n680), .Z(n382));
Q_AN02 U378 ( .A0(n443), .A1(n681), .Z(n383));
Q_AN02 U379 ( .A0(n443), .A1(n682), .Z(n384));
Q_AN02 U380 ( .A0(n443), .A1(n683), .Z(n385));
Q_AN02 U381 ( .A0(n443), .A1(n684), .Z(n386));
Q_AN02 U382 ( .A0(n443), .A1(n685), .Z(n387));
Q_AN02 U383 ( .A0(n443), .A1(n686), .Z(n388));
Q_AN02 U384 ( .A0(n443), .A1(n687), .Z(n389));
Q_AN02 U385 ( .A0(n443), .A1(n688), .Z(n390));
Q_AN02 U386 ( .A0(n443), .A1(n689), .Z(n391));
Q_AN02 U387 ( .A0(n443), .A1(n690), .Z(n392));
Q_AN02 U388 ( .A0(n443), .A1(n691), .Z(n393));
Q_AN02 U389 ( .A0(n443), .A1(n692), .Z(n394));
Q_AN02 U390 ( .A0(n443), .A1(n693), .Z(n395));
Q_AN02 U391 ( .A0(n443), .A1(n694), .Z(n396));
Q_AN02 U392 ( .A0(n443), .A1(n695), .Z(n397));
Q_AN02 U393 ( .A0(n443), .A1(n696), .Z(n398));
Q_AN02 U394 ( .A0(n443), .A1(n697), .Z(n399));
Q_AN02 U395 ( .A0(n443), .A1(n698), .Z(n400));
Q_AN02 U396 ( .A0(n443), .A1(n699), .Z(n401));
Q_AN02 U397 ( .A0(n443), .A1(n700), .Z(n402));
Q_AN02 U398 ( .A0(n443), .A1(n701), .Z(n403));
Q_AN02 U399 ( .A0(n443), .A1(n702), .Z(n404));
Q_AN02 U400 ( .A0(n443), .A1(n703), .Z(n405));
Q_AN02 U401 ( .A0(n443), .A1(n704), .Z(n406));
Q_AN02 U402 ( .A0(n443), .A1(n705), .Z(n407));
Q_AN02 U403 ( .A0(n443), .A1(n706), .Z(n408));
Q_AN02 U404 ( .A0(n443), .A1(n707), .Z(n409));
Q_AN02 U405 ( .A0(n443), .A1(n708), .Z(n410));
Q_AN02 U406 ( .A0(n443), .A1(n709), .Z(n411));
Q_AN02 U407 ( .A0(n443), .A1(n710), .Z(n412));
Q_AN02 U408 ( .A0(n443), .A1(n711), .Z(n413));
Q_AN02 U409 ( .A0(n443), .A1(n712), .Z(n414));
Q_AN02 U410 ( .A0(n443), .A1(n713), .Z(n415));
Q_AN02 U411 ( .A0(n443), .A1(n714), .Z(n416));
Q_AN02 U412 ( .A0(n443), .A1(n715), .Z(n417));
Q_AN02 U413 ( .A0(n443), .A1(n716), .Z(n418));
Q_AN02 U414 ( .A0(n443), .A1(n717), .Z(n419));
Q_AN02 U415 ( .A0(n443), .A1(n718), .Z(n420));
Q_AN02 U416 ( .A0(n443), .A1(n719), .Z(n421));
Q_AN02 U417 ( .A0(n443), .A1(n720), .Z(n422));
Q_AN02 U418 ( .A0(n443), .A1(n721), .Z(n423));
Q_AN02 U419 ( .A0(n443), .A1(n722), .Z(n424));
Q_AN02 U420 ( .A0(n443), .A1(n723), .Z(n425));
Q_AN02 U421 ( .A0(n443), .A1(n724), .Z(n426));
Q_AN02 U422 ( .A0(n443), .A1(n725), .Z(n427));
Q_AN02 U423 ( .A0(n443), .A1(n726), .Z(n428));
Q_AN02 U424 ( .A0(n443), .A1(n727), .Z(n429));
Q_AN02 U425 ( .A0(n443), .A1(n728), .Z(n430));
Q_AN02 U426 ( .A0(n443), .A1(n729), .Z(n431));
Q_AN02 U427 ( .A0(n443), .A1(n730), .Z(n432));
Q_AN02 U428 ( .A0(n443), .A1(n731), .Z(n433));
Q_AN02 U429 ( .A0(n443), .A1(n732), .Z(n434));
Q_AN02 U430 ( .A0(n443), .A1(n733), .Z(n435));
Q_AN02 U431 ( .A0(n443), .A1(n734), .Z(n436));
Q_AN02 U432 ( .A0(n443), .A1(n735), .Z(n437));
Q_AN02 U433 ( .A0(n443), .A1(n736), .Z(n438));
Q_AN02 U434 ( .A0(n443), .A1(n737), .Z(n439));
Q_AN02 U435 ( .A0(n443), .A1(n738), .Z(n440));
Q_AN02 U436 ( .A0(n443), .A1(n739), .Z(n441));
Q_AN02 U437 ( .A0(n443), .A1(n740), .Z(n442));
Q_INV U438 ( .A(pipe_ack_num_bytes[4]), .Z(n443));
Q_MX02 U439 ( .S(pipe_ack_num_bytes[4]), .A0(n741), .A1(n612), .Z(n444));
Q_MX02 U440 ( .S(pipe_ack_num_bytes[4]), .A0(n742), .A1(n613), .Z(n445));
Q_MX02 U441 ( .S(pipe_ack_num_bytes[4]), .A0(n743), .A1(n614), .Z(n446));
Q_MX02 U442 ( .S(pipe_ack_num_bytes[4]), .A0(n744), .A1(n615), .Z(n447));
Q_MX02 U443 ( .S(pipe_ack_num_bytes[4]), .A0(n745), .A1(n616), .Z(n448));
Q_MX02 U444 ( .S(pipe_ack_num_bytes[4]), .A0(n746), .A1(n617), .Z(n449));
Q_MX02 U445 ( .S(pipe_ack_num_bytes[4]), .A0(n747), .A1(n618), .Z(n450));
Q_MX02 U446 ( .S(pipe_ack_num_bytes[4]), .A0(n748), .A1(n619), .Z(n451));
Q_MX02 U447 ( .S(pipe_ack_num_bytes[4]), .A0(n749), .A1(n620), .Z(n452));
Q_MX02 U448 ( .S(pipe_ack_num_bytes[4]), .A0(n750), .A1(n621), .Z(n453));
Q_MX02 U449 ( .S(pipe_ack_num_bytes[4]), .A0(n751), .A1(n622), .Z(n454));
Q_MX02 U450 ( .S(pipe_ack_num_bytes[4]), .A0(n752), .A1(n623), .Z(n455));
Q_MX02 U451 ( .S(pipe_ack_num_bytes[4]), .A0(n753), .A1(n624), .Z(n456));
Q_MX02 U452 ( .S(pipe_ack_num_bytes[4]), .A0(n754), .A1(n625), .Z(n457));
Q_MX02 U453 ( .S(pipe_ack_num_bytes[4]), .A0(n755), .A1(n626), .Z(n458));
Q_MX02 U454 ( .S(pipe_ack_num_bytes[4]), .A0(n756), .A1(n627), .Z(n459));
Q_MX02 U455 ( .S(pipe_ack_num_bytes[4]), .A0(n757), .A1(n628), .Z(n460));
Q_MX02 U456 ( .S(pipe_ack_num_bytes[4]), .A0(n758), .A1(n629), .Z(n461));
Q_MX02 U457 ( .S(pipe_ack_num_bytes[4]), .A0(n759), .A1(n630), .Z(n462));
Q_MX02 U458 ( .S(pipe_ack_num_bytes[4]), .A0(n760), .A1(n631), .Z(n463));
Q_MX02 U459 ( .S(pipe_ack_num_bytes[4]), .A0(n761), .A1(n632), .Z(n464));
Q_MX02 U460 ( .S(pipe_ack_num_bytes[4]), .A0(n762), .A1(n633), .Z(n465));
Q_MX02 U461 ( .S(pipe_ack_num_bytes[4]), .A0(n763), .A1(n634), .Z(n466));
Q_MX02 U462 ( .S(pipe_ack_num_bytes[4]), .A0(n764), .A1(n635), .Z(n467));
Q_MX02 U463 ( .S(pipe_ack_num_bytes[4]), .A0(n765), .A1(n636), .Z(n468));
Q_MX02 U464 ( .S(pipe_ack_num_bytes[4]), .A0(n766), .A1(n637), .Z(n469));
Q_MX02 U465 ( .S(pipe_ack_num_bytes[4]), .A0(n767), .A1(n638), .Z(n470));
Q_MX02 U466 ( .S(pipe_ack_num_bytes[4]), .A0(n768), .A1(n639), .Z(n471));
Q_MX02 U467 ( .S(pipe_ack_num_bytes[4]), .A0(n769), .A1(n640), .Z(n472));
Q_MX02 U468 ( .S(pipe_ack_num_bytes[4]), .A0(n770), .A1(n641), .Z(n473));
Q_MX02 U469 ( .S(pipe_ack_num_bytes[4]), .A0(n771), .A1(n642), .Z(n474));
Q_MX02 U470 ( .S(pipe_ack_num_bytes[4]), .A0(n772), .A1(n643), .Z(n475));
Q_MX02 U471 ( .S(pipe_ack_num_bytes[4]), .A0(n773), .A1(n644), .Z(n476));
Q_MX02 U472 ( .S(pipe_ack_num_bytes[4]), .A0(n774), .A1(n645), .Z(n477));
Q_MX02 U473 ( .S(pipe_ack_num_bytes[4]), .A0(n775), .A1(n646), .Z(n478));
Q_MX02 U474 ( .S(pipe_ack_num_bytes[4]), .A0(n776), .A1(n647), .Z(n479));
Q_MX02 U475 ( .S(pipe_ack_num_bytes[4]), .A0(n777), .A1(n648), .Z(n480));
Q_MX02 U476 ( .S(pipe_ack_num_bytes[4]), .A0(n778), .A1(n649), .Z(n481));
Q_MX02 U477 ( .S(pipe_ack_num_bytes[4]), .A0(n779), .A1(n650), .Z(n482));
Q_MX02 U478 ( .S(pipe_ack_num_bytes[4]), .A0(n780), .A1(n651), .Z(n483));
Q_MX03 U479 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n950), .A1(n886), .A2(n652), .Z(n484));
Q_MX03 U480 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n951), .A1(n887), .A2(n653), .Z(n485));
Q_MX03 U481 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n952), .A1(n888), .A2(n654), .Z(n486));
Q_MX03 U482 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n953), .A1(n889), .A2(n655), .Z(n487));
Q_MX03 U483 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n954), .A1(n890), .A2(n656), .Z(n488));
Q_MX03 U484 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n955), .A1(n891), .A2(n657), .Z(n489));
Q_MX03 U485 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n956), .A1(n892), .A2(n658), .Z(n490));
Q_MX03 U486 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n957), .A1(n893), .A2(n659), .Z(n491));
Q_MX03 U487 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n958), .A1(n894), .A2(n660), .Z(n492));
Q_MX03 U488 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n959), .A1(n895), .A2(n661), .Z(n493));
Q_MX03 U489 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n960), .A1(n896), .A2(n662), .Z(n494));
Q_MX03 U490 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n961), .A1(n897), .A2(n663), .Z(n495));
Q_MX03 U491 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n962), .A1(n898), .A2(n664), .Z(n496));
Q_MX03 U492 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n963), .A1(n899), .A2(n665), .Z(n497));
Q_MX03 U493 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n964), .A1(n900), .A2(n666), .Z(n498));
Q_MX03 U494 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n965), .A1(n901), .A2(n667), .Z(n499));
Q_MX03 U495 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n966), .A1(n902), .A2(n668), .Z(n500));
Q_MX03 U496 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n967), .A1(n903), .A2(n669), .Z(n501));
Q_MX03 U497 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n968), .A1(n904), .A2(n670), .Z(n502));
Q_MX03 U498 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n969), .A1(n905), .A2(n671), .Z(n503));
Q_MX03 U499 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n970), .A1(n906), .A2(n672), .Z(n504));
Q_MX03 U500 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n971), .A1(n907), .A2(n673), .Z(n505));
Q_MX03 U501 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n972), .A1(n908), .A2(n674), .Z(n506));
Q_MX03 U502 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n973), .A1(n909), .A2(n675), .Z(n507));
Q_MX03 U503 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n974), .A1(n910), .A2(n677), .Z(n508));
Q_MX03 U504 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n975), .A1(n911), .A2(n678), .Z(n509));
Q_MX03 U505 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n976), .A1(n912), .A2(n679), .Z(n510));
Q_MX03 U506 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n977), .A1(n913), .A2(n680), .Z(n511));
Q_MX03 U507 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n978), .A1(n914), .A2(n681), .Z(n512));
Q_MX03 U508 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n979), .A1(n915), .A2(n682), .Z(n513));
Q_MX03 U509 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n980), .A1(n916), .A2(n683), .Z(n514));
Q_MX03 U510 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n981), .A1(n917), .A2(n684), .Z(n515));
Q_MX03 U511 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n982), .A1(n918), .A2(n685), .Z(n516));
Q_MX03 U512 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n983), .A1(n919), .A2(n686), .Z(n517));
Q_MX03 U513 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n984), .A1(n920), .A2(n687), .Z(n518));
Q_MX03 U514 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n985), .A1(n921), .A2(n688), .Z(n519));
Q_MX03 U515 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n986), .A1(n922), .A2(n689), .Z(n520));
Q_MX03 U516 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n987), .A1(n923), .A2(n690), .Z(n521));
Q_MX03 U517 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n988), .A1(n924), .A2(n691), .Z(n522));
Q_MX03 U518 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n989), .A1(n925), .A2(n692), .Z(n523));
Q_MX03 U519 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n990), .A1(n926), .A2(n693), .Z(n524));
Q_MX03 U520 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n991), .A1(n927), .A2(n694), .Z(n525));
Q_MX03 U521 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n992), .A1(n928), .A2(n695), .Z(n526));
Q_MX03 U522 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n993), .A1(n929), .A2(n696), .Z(n527));
Q_MX03 U523 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n994), .A1(n930), .A2(n697), .Z(n528));
Q_MX03 U524 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n995), .A1(n931), .A2(n698), .Z(n529));
Q_MX03 U525 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n996), .A1(n932), .A2(n699), .Z(n530));
Q_MX03 U526 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n997), .A1(n933), .A2(n700), .Z(n531));
Q_MX03 U527 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n998), .A1(n934), .A2(n701), .Z(n532));
Q_MX03 U528 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n999), .A1(n935), .A2(n702), .Z(n533));
Q_MX03 U529 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1000), .A1(n936), .A2(n703), .Z(n534));
Q_MX03 U530 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1001), .A1(n937), .A2(n704), .Z(n535));
Q_MX03 U531 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1002), .A1(n938), .A2(n705), .Z(n536));
Q_MX03 U532 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1003), .A1(n939), .A2(n706), .Z(n537));
Q_MX03 U533 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1004), .A1(n940), .A2(n707), .Z(n538));
Q_MX03 U534 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1005), .A1(n941), .A2(n708), .Z(n539));
Q_MX03 U535 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1006), .A1(n942), .A2(n709), .Z(n540));
Q_MX03 U536 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1007), .A1(n943), .A2(n710), .Z(n541));
Q_MX03 U537 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1008), .A1(n944), .A2(n711), .Z(n542));
Q_MX03 U538 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1009), .A1(n945), .A2(n712), .Z(n543));
Q_MX03 U539 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1010), .A1(n946), .A2(n713), .Z(n544));
Q_MX03 U540 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1011), .A1(n947), .A2(n714), .Z(n545));
Q_MX03 U541 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1012), .A1(n948), .A2(n715), .Z(n546));
Q_MX03 U542 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1013), .A1(n949), .A2(n716), .Z(n547));
Q_MX03 U543 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1014), .A1(n950), .A2(n717), .Z(n548));
Q_MX03 U544 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1015), .A1(n951), .A2(n718), .Z(n549));
Q_MX03 U545 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1016), .A1(n952), .A2(n719), .Z(n550));
Q_MX03 U546 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1017), .A1(n953), .A2(n720), .Z(n551));
Q_MX03 U547 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1018), .A1(n954), .A2(n721), .Z(n552));
Q_MX03 U548 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1019), .A1(n955), .A2(n722), .Z(n553));
Q_MX03 U549 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1020), .A1(n956), .A2(n723), .Z(n554));
Q_MX03 U550 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1021), .A1(n957), .A2(n724), .Z(n555));
Q_MX03 U551 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1022), .A1(n958), .A2(n725), .Z(n556));
Q_MX03 U552 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1023), .A1(n959), .A2(n726), .Z(n557));
Q_MX03 U553 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1024), .A1(n960), .A2(n727), .Z(n558));
Q_MX03 U554 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1025), .A1(n961), .A2(n728), .Z(n559));
Q_MX03 U555 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1026), .A1(n962), .A2(n729), .Z(n560));
Q_MX03 U556 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1027), .A1(n963), .A2(n730), .Z(n561));
Q_MX03 U557 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1028), .A1(n964), .A2(n731), .Z(n562));
Q_MX03 U558 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1029), .A1(n965), .A2(n732), .Z(n563));
Q_MX03 U559 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1030), .A1(n966), .A2(n733), .Z(n564));
Q_MX03 U560 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1031), .A1(n967), .A2(n734), .Z(n565));
Q_MX03 U561 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1032), .A1(n968), .A2(n735), .Z(n566));
Q_MX03 U562 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1033), .A1(n969), .A2(n736), .Z(n567));
Q_MX03 U563 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1034), .A1(n970), .A2(n737), .Z(n568));
Q_MX03 U564 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1035), .A1(n971), .A2(n738), .Z(n569));
Q_MX03 U565 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1036), .A1(n972), .A2(n739), .Z(n570));
Q_MX03 U566 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1037), .A1(n973), .A2(n740), .Z(n571));
Q_MX03 U567 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1038), .A1(n974), .A2(n741), .Z(n572));
Q_MX03 U568 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1039), .A1(n975), .A2(n742), .Z(n573));
Q_MX03 U569 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1040), .A1(n976), .A2(n743), .Z(n574));
Q_MX03 U570 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1041), .A1(n977), .A2(n744), .Z(n575));
Q_MX03 U571 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1042), .A1(n978), .A2(n745), .Z(n576));
Q_MX03 U572 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1043), .A1(n979), .A2(n746), .Z(n577));
Q_MX03 U573 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1044), .A1(n980), .A2(n747), .Z(n578));
Q_MX03 U574 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1045), .A1(n981), .A2(n748), .Z(n579));
Q_MX03 U575 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1046), .A1(n982), .A2(n749), .Z(n580));
Q_MX03 U576 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1047), .A1(n983), .A2(n750), .Z(n581));
Q_MX03 U577 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1048), .A1(n984), .A2(n751), .Z(n582));
Q_MX03 U578 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1049), .A1(n985), .A2(n752), .Z(n583));
Q_MX03 U579 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1050), .A1(n986), .A2(n753), .Z(n584));
Q_MX03 U580 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1051), .A1(n987), .A2(n754), .Z(n585));
Q_MX03 U581 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1052), .A1(n988), .A2(n755), .Z(n586));
Q_MX03 U582 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1053), .A1(n989), .A2(n756), .Z(n587));
Q_MX03 U583 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1054), .A1(n990), .A2(n757), .Z(n588));
Q_MX03 U584 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1055), .A1(n991), .A2(n758), .Z(n589));
Q_MX03 U585 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1056), .A1(n992), .A2(n759), .Z(n590));
Q_MX03 U586 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1057), .A1(n993), .A2(n760), .Z(n591));
Q_MX03 U587 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1058), .A1(n994), .A2(n761), .Z(n592));
Q_MX03 U588 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1059), .A1(n995), .A2(n762), .Z(n593));
Q_MX03 U589 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1060), .A1(n996), .A2(n763), .Z(n594));
Q_MX03 U590 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1061), .A1(n997), .A2(n764), .Z(n595));
Q_MX03 U591 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1062), .A1(n998), .A2(n765), .Z(n596));
Q_MX03 U592 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1063), .A1(n999), .A2(n766), .Z(n597));
Q_MX03 U593 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1064), .A1(n1000), .A2(n767), .Z(n598));
Q_MX03 U594 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1065), .A1(n1001), .A2(n768), .Z(n599));
Q_MX03 U595 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1066), .A1(n1002), .A2(n769), .Z(n600));
Q_MX03 U596 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1067), .A1(n1003), .A2(n770), .Z(n601));
Q_MX03 U597 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1068), .A1(n1004), .A2(n771), .Z(n602));
Q_MX03 U598 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1069), .A1(n1005), .A2(n772), .Z(n603));
Q_MX03 U599 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1070), .A1(n1006), .A2(n773), .Z(n604));
Q_MX03 U600 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1071), .A1(n1007), .A2(n774), .Z(n605));
Q_MX03 U601 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1072), .A1(n1008), .A2(n775), .Z(n606));
Q_MX03 U602 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1073), .A1(n1009), .A2(n776), .Z(n607));
Q_MX03 U603 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1074), .A1(n1010), .A2(n777), .Z(n608));
Q_MX03 U604 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1075), .A1(n1011), .A2(n778), .Z(n609));
Q_MX03 U605 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1076), .A1(n1012), .A2(n779), .Z(n610));
Q_MX03 U606 ( .S0(pipe_ack_num_bytes[3]), .S1(pipe_ack_num_bytes[4]), .A0(n1077), .A1(n1013), .A2(n780), .Z(n611));
Q_AN02 U607 ( .A0(n676), .A1(n781), .Z(n612));
Q_AN02 U608 ( .A0(n676), .A1(n782), .Z(n613));
Q_AN02 U609 ( .A0(n676), .A1(n783), .Z(n614));
Q_AN02 U610 ( .A0(n676), .A1(n784), .Z(n615));
Q_AN02 U611 ( .A0(n676), .A1(n785), .Z(n616));
Q_AN02 U612 ( .A0(n676), .A1(n786), .Z(n617));
Q_AN02 U613 ( .A0(n676), .A1(n787), .Z(n618));
Q_AN02 U614 ( .A0(n676), .A1(n788), .Z(n619));
Q_AN02 U615 ( .A0(n676), .A1(n789), .Z(n620));
Q_AN02 U616 ( .A0(n676), .A1(n790), .Z(n621));
Q_AN02 U617 ( .A0(n676), .A1(n791), .Z(n622));
Q_AN02 U618 ( .A0(n676), .A1(n792), .Z(n623));
Q_AN02 U619 ( .A0(n676), .A1(n793), .Z(n624));
Q_AN02 U620 ( .A0(n676), .A1(n794), .Z(n625));
Q_AN02 U621 ( .A0(n676), .A1(n795), .Z(n626));
Q_AN02 U622 ( .A0(n676), .A1(n796), .Z(n627));
Q_AN02 U623 ( .A0(n676), .A1(n797), .Z(n628));
Q_AN02 U624 ( .A0(n676), .A1(n798), .Z(n629));
Q_AN02 U625 ( .A0(n676), .A1(n799), .Z(n630));
Q_AN02 U626 ( .A0(n676), .A1(n800), .Z(n631));
Q_AN02 U627 ( .A0(n676), .A1(n801), .Z(n632));
Q_AN02 U628 ( .A0(n676), .A1(n802), .Z(n633));
Q_AN02 U629 ( .A0(n676), .A1(n803), .Z(n634));
Q_AN02 U630 ( .A0(n676), .A1(n804), .Z(n635));
Q_AN02 U631 ( .A0(n676), .A1(n805), .Z(n636));
Q_AN02 U632 ( .A0(n676), .A1(n806), .Z(n637));
Q_AN02 U633 ( .A0(n676), .A1(n807), .Z(n638));
Q_AN02 U634 ( .A0(n676), .A1(n808), .Z(n639));
Q_AN02 U635 ( .A0(n676), .A1(n809), .Z(n640));
Q_AN02 U636 ( .A0(n676), .A1(n810), .Z(n641));
Q_AN02 U637 ( .A0(n676), .A1(n811), .Z(n642));
Q_AN02 U638 ( .A0(n676), .A1(n812), .Z(n643));
Q_AN02 U639 ( .A0(n676), .A1(n814), .Z(n644));
Q_AN02 U640 ( .A0(n676), .A1(n815), .Z(n645));
Q_AN02 U641 ( .A0(n676), .A1(n816), .Z(n646));
Q_AN02 U642 ( .A0(n676), .A1(n817), .Z(n647));
Q_AN02 U643 ( .A0(n676), .A1(n818), .Z(n648));
Q_AN02 U644 ( .A0(n676), .A1(n819), .Z(n649));
Q_AN02 U645 ( .A0(n676), .A1(n820), .Z(n650));
Q_AN02 U646 ( .A0(n676), .A1(n821), .Z(n651));
Q_AN02 U647 ( .A0(n676), .A1(n822), .Z(n652));
Q_AN02 U648 ( .A0(n676), .A1(n823), .Z(n653));
Q_AN02 U649 ( .A0(n676), .A1(n824), .Z(n654));
Q_AN02 U650 ( .A0(n676), .A1(n825), .Z(n655));
Q_AN02 U651 ( .A0(n676), .A1(n826), .Z(n656));
Q_AN02 U652 ( .A0(n676), .A1(n827), .Z(n657));
Q_AN02 U653 ( .A0(n676), .A1(n828), .Z(n658));
Q_AN02 U654 ( .A0(n676), .A1(n829), .Z(n659));
Q_AN02 U655 ( .A0(n676), .A1(n830), .Z(n660));
Q_AN02 U656 ( .A0(n676), .A1(n831), .Z(n661));
Q_AN02 U657 ( .A0(n676), .A1(n832), .Z(n662));
Q_AN02 U658 ( .A0(n676), .A1(n833), .Z(n663));
Q_AN02 U659 ( .A0(n676), .A1(n834), .Z(n664));
Q_AN02 U660 ( .A0(n676), .A1(n835), .Z(n665));
Q_AN02 U661 ( .A0(n676), .A1(n836), .Z(n666));
Q_AN02 U662 ( .A0(n676), .A1(n837), .Z(n667));
Q_AN02 U663 ( .A0(n676), .A1(n838), .Z(n668));
Q_AN02 U664 ( .A0(n676), .A1(n839), .Z(n669));
Q_AN02 U665 ( .A0(n676), .A1(n840), .Z(n670));
Q_AN02 U666 ( .A0(n676), .A1(n841), .Z(n671));
Q_AN02 U667 ( .A0(n676), .A1(n842), .Z(n672));
Q_AN02 U668 ( .A0(n676), .A1(n843), .Z(n673));
Q_AN02 U669 ( .A0(n676), .A1(n844), .Z(n674));
Q_AN02 U670 ( .A0(n676), .A1(n845), .Z(n675));
Q_INV U671 ( .A(pipe_ack_num_bytes[3]), .Z(n676));
Q_MX02 U672 ( .S(pipe_ack_num_bytes[3]), .A0(n846), .A1(n781), .Z(n677));
Q_MX02 U673 ( .S(pipe_ack_num_bytes[3]), .A0(n847), .A1(n782), .Z(n678));
Q_MX02 U674 ( .S(pipe_ack_num_bytes[3]), .A0(n848), .A1(n783), .Z(n679));
Q_MX02 U675 ( .S(pipe_ack_num_bytes[3]), .A0(n849), .A1(n784), .Z(n680));
Q_MX02 U676 ( .S(pipe_ack_num_bytes[3]), .A0(n850), .A1(n785), .Z(n681));
Q_MX02 U677 ( .S(pipe_ack_num_bytes[3]), .A0(n851), .A1(n786), .Z(n682));
Q_MX02 U678 ( .S(pipe_ack_num_bytes[3]), .A0(n852), .A1(n787), .Z(n683));
Q_MX02 U679 ( .S(pipe_ack_num_bytes[3]), .A0(n853), .A1(n788), .Z(n684));
Q_MX02 U680 ( .S(pipe_ack_num_bytes[3]), .A0(n854), .A1(n789), .Z(n685));
Q_MX02 U681 ( .S(pipe_ack_num_bytes[3]), .A0(n855), .A1(n790), .Z(n686));
Q_MX02 U682 ( .S(pipe_ack_num_bytes[3]), .A0(n856), .A1(n791), .Z(n687));
Q_MX02 U683 ( .S(pipe_ack_num_bytes[3]), .A0(n857), .A1(n792), .Z(n688));
Q_MX02 U684 ( .S(pipe_ack_num_bytes[3]), .A0(n858), .A1(n793), .Z(n689));
Q_MX02 U685 ( .S(pipe_ack_num_bytes[3]), .A0(n859), .A1(n794), .Z(n690));
Q_MX02 U686 ( .S(pipe_ack_num_bytes[3]), .A0(n860), .A1(n795), .Z(n691));
Q_MX02 U687 ( .S(pipe_ack_num_bytes[3]), .A0(n861), .A1(n796), .Z(n692));
Q_MX02 U688 ( .S(pipe_ack_num_bytes[3]), .A0(n862), .A1(n797), .Z(n693));
Q_MX02 U689 ( .S(pipe_ack_num_bytes[3]), .A0(n863), .A1(n798), .Z(n694));
Q_MX02 U690 ( .S(pipe_ack_num_bytes[3]), .A0(n864), .A1(n799), .Z(n695));
Q_MX02 U691 ( .S(pipe_ack_num_bytes[3]), .A0(n865), .A1(n800), .Z(n696));
Q_MX02 U692 ( .S(pipe_ack_num_bytes[3]), .A0(n866), .A1(n801), .Z(n697));
Q_MX02 U693 ( .S(pipe_ack_num_bytes[3]), .A0(n867), .A1(n802), .Z(n698));
Q_MX02 U694 ( .S(pipe_ack_num_bytes[3]), .A0(n868), .A1(n803), .Z(n699));
Q_MX02 U695 ( .S(pipe_ack_num_bytes[3]), .A0(n869), .A1(n804), .Z(n700));
Q_MX02 U696 ( .S(pipe_ack_num_bytes[3]), .A0(n870), .A1(n805), .Z(n701));
Q_MX02 U697 ( .S(pipe_ack_num_bytes[3]), .A0(n871), .A1(n806), .Z(n702));
Q_MX02 U698 ( .S(pipe_ack_num_bytes[3]), .A0(n872), .A1(n807), .Z(n703));
Q_MX02 U699 ( .S(pipe_ack_num_bytes[3]), .A0(n873), .A1(n808), .Z(n704));
Q_MX02 U700 ( .S(pipe_ack_num_bytes[3]), .A0(n874), .A1(n809), .Z(n705));
Q_MX02 U701 ( .S(pipe_ack_num_bytes[3]), .A0(n875), .A1(n810), .Z(n706));
Q_MX02 U702 ( .S(pipe_ack_num_bytes[3]), .A0(n876), .A1(n811), .Z(n707));
Q_MX02 U703 ( .S(pipe_ack_num_bytes[3]), .A0(n877), .A1(n812), .Z(n708));
Q_MX02 U704 ( .S(pipe_ack_num_bytes[3]), .A0(n878), .A1(n814), .Z(n709));
Q_MX02 U705 ( .S(pipe_ack_num_bytes[3]), .A0(n879), .A1(n815), .Z(n710));
Q_MX02 U706 ( .S(pipe_ack_num_bytes[3]), .A0(n880), .A1(n816), .Z(n711));
Q_MX02 U707 ( .S(pipe_ack_num_bytes[3]), .A0(n881), .A1(n817), .Z(n712));
Q_MX02 U708 ( .S(pipe_ack_num_bytes[3]), .A0(n882), .A1(n818), .Z(n713));
Q_MX02 U709 ( .S(pipe_ack_num_bytes[3]), .A0(n883), .A1(n819), .Z(n714));
Q_MX02 U710 ( .S(pipe_ack_num_bytes[3]), .A0(n884), .A1(n820), .Z(n715));
Q_MX02 U711 ( .S(pipe_ack_num_bytes[3]), .A0(n885), .A1(n821), .Z(n716));
Q_MX02 U712 ( .S(pipe_ack_num_bytes[3]), .A0(n886), .A1(n822), .Z(n717));
Q_MX02 U713 ( .S(pipe_ack_num_bytes[3]), .A0(n887), .A1(n823), .Z(n718));
Q_MX02 U714 ( .S(pipe_ack_num_bytes[3]), .A0(n888), .A1(n824), .Z(n719));
Q_MX02 U715 ( .S(pipe_ack_num_bytes[3]), .A0(n889), .A1(n825), .Z(n720));
Q_MX02 U716 ( .S(pipe_ack_num_bytes[3]), .A0(n890), .A1(n826), .Z(n721));
Q_MX02 U717 ( .S(pipe_ack_num_bytes[3]), .A0(n891), .A1(n827), .Z(n722));
Q_MX02 U718 ( .S(pipe_ack_num_bytes[3]), .A0(n892), .A1(n828), .Z(n723));
Q_MX02 U719 ( .S(pipe_ack_num_bytes[3]), .A0(n893), .A1(n829), .Z(n724));
Q_MX02 U720 ( .S(pipe_ack_num_bytes[3]), .A0(n894), .A1(n830), .Z(n725));
Q_MX02 U721 ( .S(pipe_ack_num_bytes[3]), .A0(n895), .A1(n831), .Z(n726));
Q_MX02 U722 ( .S(pipe_ack_num_bytes[3]), .A0(n896), .A1(n832), .Z(n727));
Q_MX02 U723 ( .S(pipe_ack_num_bytes[3]), .A0(n897), .A1(n833), .Z(n728));
Q_MX02 U724 ( .S(pipe_ack_num_bytes[3]), .A0(n898), .A1(n834), .Z(n729));
Q_MX02 U725 ( .S(pipe_ack_num_bytes[3]), .A0(n899), .A1(n835), .Z(n730));
Q_MX02 U726 ( .S(pipe_ack_num_bytes[3]), .A0(n900), .A1(n836), .Z(n731));
Q_MX02 U727 ( .S(pipe_ack_num_bytes[3]), .A0(n901), .A1(n837), .Z(n732));
Q_MX02 U728 ( .S(pipe_ack_num_bytes[3]), .A0(n902), .A1(n838), .Z(n733));
Q_MX02 U729 ( .S(pipe_ack_num_bytes[3]), .A0(n903), .A1(n839), .Z(n734));
Q_MX02 U730 ( .S(pipe_ack_num_bytes[3]), .A0(n904), .A1(n840), .Z(n735));
Q_MX02 U731 ( .S(pipe_ack_num_bytes[3]), .A0(n905), .A1(n841), .Z(n736));
Q_MX02 U732 ( .S(pipe_ack_num_bytes[3]), .A0(n906), .A1(n842), .Z(n737));
Q_MX02 U733 ( .S(pipe_ack_num_bytes[3]), .A0(n907), .A1(n843), .Z(n738));
Q_MX02 U734 ( .S(pipe_ack_num_bytes[3]), .A0(n908), .A1(n844), .Z(n739));
Q_MX02 U735 ( .S(pipe_ack_num_bytes[3]), .A0(n909), .A1(n845), .Z(n740));
Q_MX02 U736 ( .S(pipe_ack_num_bytes[3]), .A0(n910), .A1(n846), .Z(n741));
Q_MX02 U737 ( .S(pipe_ack_num_bytes[3]), .A0(n911), .A1(n847), .Z(n742));
Q_MX02 U738 ( .S(pipe_ack_num_bytes[3]), .A0(n912), .A1(n848), .Z(n743));
Q_MX02 U739 ( .S(pipe_ack_num_bytes[3]), .A0(n913), .A1(n849), .Z(n744));
Q_MX02 U740 ( .S(pipe_ack_num_bytes[3]), .A0(n914), .A1(n850), .Z(n745));
Q_MX02 U741 ( .S(pipe_ack_num_bytes[3]), .A0(n915), .A1(n851), .Z(n746));
Q_MX02 U742 ( .S(pipe_ack_num_bytes[3]), .A0(n916), .A1(n852), .Z(n747));
Q_MX02 U743 ( .S(pipe_ack_num_bytes[3]), .A0(n917), .A1(n853), .Z(n748));
Q_MX02 U744 ( .S(pipe_ack_num_bytes[3]), .A0(n918), .A1(n854), .Z(n749));
Q_MX02 U745 ( .S(pipe_ack_num_bytes[3]), .A0(n919), .A1(n855), .Z(n750));
Q_MX02 U746 ( .S(pipe_ack_num_bytes[3]), .A0(n920), .A1(n856), .Z(n751));
Q_MX02 U747 ( .S(pipe_ack_num_bytes[3]), .A0(n921), .A1(n857), .Z(n752));
Q_MX02 U748 ( .S(pipe_ack_num_bytes[3]), .A0(n922), .A1(n858), .Z(n753));
Q_MX02 U749 ( .S(pipe_ack_num_bytes[3]), .A0(n923), .A1(n859), .Z(n754));
Q_MX02 U750 ( .S(pipe_ack_num_bytes[3]), .A0(n924), .A1(n860), .Z(n755));
Q_MX02 U751 ( .S(pipe_ack_num_bytes[3]), .A0(n925), .A1(n861), .Z(n756));
Q_MX02 U752 ( .S(pipe_ack_num_bytes[3]), .A0(n926), .A1(n862), .Z(n757));
Q_MX02 U753 ( .S(pipe_ack_num_bytes[3]), .A0(n927), .A1(n863), .Z(n758));
Q_MX02 U754 ( .S(pipe_ack_num_bytes[3]), .A0(n928), .A1(n864), .Z(n759));
Q_MX02 U755 ( .S(pipe_ack_num_bytes[3]), .A0(n929), .A1(n865), .Z(n760));
Q_MX02 U756 ( .S(pipe_ack_num_bytes[3]), .A0(n930), .A1(n866), .Z(n761));
Q_MX02 U757 ( .S(pipe_ack_num_bytes[3]), .A0(n931), .A1(n867), .Z(n762));
Q_MX02 U758 ( .S(pipe_ack_num_bytes[3]), .A0(n932), .A1(n868), .Z(n763));
Q_MX02 U759 ( .S(pipe_ack_num_bytes[3]), .A0(n933), .A1(n869), .Z(n764));
Q_MX02 U760 ( .S(pipe_ack_num_bytes[3]), .A0(n934), .A1(n870), .Z(n765));
Q_MX02 U761 ( .S(pipe_ack_num_bytes[3]), .A0(n935), .A1(n871), .Z(n766));
Q_MX02 U762 ( .S(pipe_ack_num_bytes[3]), .A0(n936), .A1(n872), .Z(n767));
Q_MX02 U763 ( .S(pipe_ack_num_bytes[3]), .A0(n937), .A1(n873), .Z(n768));
Q_MX02 U764 ( .S(pipe_ack_num_bytes[3]), .A0(n938), .A1(n874), .Z(n769));
Q_MX02 U765 ( .S(pipe_ack_num_bytes[3]), .A0(n939), .A1(n875), .Z(n770));
Q_MX02 U766 ( .S(pipe_ack_num_bytes[3]), .A0(n940), .A1(n876), .Z(n771));
Q_MX02 U767 ( .S(pipe_ack_num_bytes[3]), .A0(n941), .A1(n877), .Z(n772));
Q_MX02 U768 ( .S(pipe_ack_num_bytes[3]), .A0(n942), .A1(n878), .Z(n773));
Q_MX02 U769 ( .S(pipe_ack_num_bytes[3]), .A0(n943), .A1(n879), .Z(n774));
Q_MX02 U770 ( .S(pipe_ack_num_bytes[3]), .A0(n944), .A1(n880), .Z(n775));
Q_MX02 U771 ( .S(pipe_ack_num_bytes[3]), .A0(n945), .A1(n881), .Z(n776));
Q_MX02 U772 ( .S(pipe_ack_num_bytes[3]), .A0(n946), .A1(n882), .Z(n777));
Q_MX02 U773 ( .S(pipe_ack_num_bytes[3]), .A0(n947), .A1(n883), .Z(n778));
Q_MX02 U774 ( .S(pipe_ack_num_bytes[3]), .A0(n948), .A1(n884), .Z(n779));
Q_MX02 U775 ( .S(pipe_ack_num_bytes[3]), .A0(n949), .A1(n885), .Z(n780));
Q_AN02 U776 ( .A0(n813), .A1(n1078), .Z(n781));
Q_AN02 U777 ( .A0(n813), .A1(n1079), .Z(n782));
Q_AN02 U778 ( .A0(n813), .A1(n1080), .Z(n783));
Q_AN02 U779 ( .A0(n813), .A1(n1081), .Z(n784));
Q_AN02 U780 ( .A0(n813), .A1(n1082), .Z(n785));
Q_AN02 U781 ( .A0(n813), .A1(n1083), .Z(n786));
Q_AN02 U782 ( .A0(n813), .A1(n1084), .Z(n787));
Q_AN02 U783 ( .A0(n813), .A1(n1085), .Z(n788));
Q_AN02 U784 ( .A0(n813), .A1(n1086), .Z(n789));
Q_AN02 U785 ( .A0(n813), .A1(n1087), .Z(n790));
Q_AN02 U786 ( .A0(n813), .A1(n1088), .Z(n791));
Q_AN02 U787 ( .A0(n813), .A1(n1089), .Z(n792));
Q_AN02 U788 ( .A0(n813), .A1(n1090), .Z(n793));
Q_AN02 U789 ( .A0(n813), .A1(n1091), .Z(n794));
Q_AN02 U790 ( .A0(n813), .A1(n1092), .Z(n795));
Q_AN02 U791 ( .A0(n813), .A1(n1093), .Z(n796));
Q_AN02 U792 ( .A0(n813), .A1(n1095), .Z(n797));
Q_AN02 U793 ( .A0(n813), .A1(n1096), .Z(n798));
Q_AN02 U794 ( .A0(n813), .A1(n1097), .Z(n799));
Q_AN02 U795 ( .A0(n813), .A1(n1098), .Z(n800));
Q_AN02 U796 ( .A0(n813), .A1(n1099), .Z(n801));
Q_AN02 U797 ( .A0(n813), .A1(n1100), .Z(n802));
Q_AN02 U798 ( .A0(n813), .A1(n1101), .Z(n803));
Q_AN02 U799 ( .A0(n813), .A1(n1102), .Z(n804));
Q_AN02 U800 ( .A0(n813), .A1(n1103), .Z(n805));
Q_AN02 U801 ( .A0(n813), .A1(n1104), .Z(n806));
Q_AN02 U802 ( .A0(n813), .A1(n1105), .Z(n807));
Q_AN02 U803 ( .A0(n813), .A1(n1106), .Z(n808));
Q_AN02 U804 ( .A0(n813), .A1(n1107), .Z(n809));
Q_AN02 U805 ( .A0(n813), .A1(n1108), .Z(n810));
Q_AN02 U806 ( .A0(n813), .A1(n1109), .Z(n811));
Q_AN02 U807 ( .A0(n813), .A1(n1110), .Z(n812));
Q_INV U808 ( .A(pipe_ack_num_bytes[2]), .Z(n813));
Q_MX02 U809 ( .S(pipe_ack_num_bytes[2]), .A0(n1111), .A1(n1078), .Z(n814));
Q_MX02 U810 ( .S(pipe_ack_num_bytes[2]), .A0(n1112), .A1(n1079), .Z(n815));
Q_MX02 U811 ( .S(pipe_ack_num_bytes[2]), .A0(n1113), .A1(n1080), .Z(n816));
Q_MX02 U812 ( .S(pipe_ack_num_bytes[2]), .A0(n1114), .A1(n1081), .Z(n817));
Q_MX02 U813 ( .S(pipe_ack_num_bytes[2]), .A0(n1115), .A1(n1082), .Z(n818));
Q_MX02 U814 ( .S(pipe_ack_num_bytes[2]), .A0(n1116), .A1(n1083), .Z(n819));
Q_MX02 U815 ( .S(pipe_ack_num_bytes[2]), .A0(n1117), .A1(n1084), .Z(n820));
Q_MX02 U816 ( .S(pipe_ack_num_bytes[2]), .A0(n1118), .A1(n1085), .Z(n821));
Q_MX02 U817 ( .S(pipe_ack_num_bytes[2]), .A0(n1119), .A1(n1086), .Z(n822));
Q_MX02 U818 ( .S(pipe_ack_num_bytes[2]), .A0(n1120), .A1(n1087), .Z(n823));
Q_MX02 U819 ( .S(pipe_ack_num_bytes[2]), .A0(n1121), .A1(n1088), .Z(n824));
Q_MX02 U820 ( .S(pipe_ack_num_bytes[2]), .A0(n1122), .A1(n1089), .Z(n825));
Q_MX02 U821 ( .S(pipe_ack_num_bytes[2]), .A0(n1123), .A1(n1090), .Z(n826));
Q_MX02 U822 ( .S(pipe_ack_num_bytes[2]), .A0(n1124), .A1(n1091), .Z(n827));
Q_MX02 U823 ( .S(pipe_ack_num_bytes[2]), .A0(n1125), .A1(n1092), .Z(n828));
Q_MX02 U824 ( .S(pipe_ack_num_bytes[2]), .A0(n1126), .A1(n1093), .Z(n829));
Q_MX02 U825 ( .S(pipe_ack_num_bytes[2]), .A0(n1127), .A1(n1095), .Z(n830));
Q_MX02 U826 ( .S(pipe_ack_num_bytes[2]), .A0(n1128), .A1(n1096), .Z(n831));
Q_MX02 U827 ( .S(pipe_ack_num_bytes[2]), .A0(n1129), .A1(n1097), .Z(n832));
Q_MX02 U828 ( .S(pipe_ack_num_bytes[2]), .A0(n1130), .A1(n1098), .Z(n833));
Q_MX02 U829 ( .S(pipe_ack_num_bytes[2]), .A0(n1131), .A1(n1099), .Z(n834));
Q_MX02 U830 ( .S(pipe_ack_num_bytes[2]), .A0(n1132), .A1(n1100), .Z(n835));
Q_MX02 U831 ( .S(pipe_ack_num_bytes[2]), .A0(n1133), .A1(n1101), .Z(n836));
Q_MX02 U832 ( .S(pipe_ack_num_bytes[2]), .A0(n1134), .A1(n1102), .Z(n837));
Q_MX02 U833 ( .S(pipe_ack_num_bytes[2]), .A0(n1135), .A1(n1103), .Z(n838));
Q_MX02 U834 ( .S(pipe_ack_num_bytes[2]), .A0(n1136), .A1(n1104), .Z(n839));
Q_MX02 U835 ( .S(pipe_ack_num_bytes[2]), .A0(n1137), .A1(n1105), .Z(n840));
Q_MX02 U836 ( .S(pipe_ack_num_bytes[2]), .A0(n1138), .A1(n1106), .Z(n841));
Q_MX02 U837 ( .S(pipe_ack_num_bytes[2]), .A0(n1139), .A1(n1107), .Z(n842));
Q_MX02 U838 ( .S(pipe_ack_num_bytes[2]), .A0(n1140), .A1(n1108), .Z(n843));
Q_MX02 U839 ( .S(pipe_ack_num_bytes[2]), .A0(n1141), .A1(n1109), .Z(n844));
Q_MX02 U840 ( .S(pipe_ack_num_bytes[2]), .A0(n1142), .A1(n1110), .Z(n845));
Q_MX02 U841 ( .S(pipe_ack_num_bytes[2]), .A0(n1143), .A1(n1111), .Z(n846));
Q_MX02 U842 ( .S(pipe_ack_num_bytes[2]), .A0(n1144), .A1(n1112), .Z(n847));
Q_MX02 U843 ( .S(pipe_ack_num_bytes[2]), .A0(n1145), .A1(n1113), .Z(n848));
Q_MX02 U844 ( .S(pipe_ack_num_bytes[2]), .A0(n1146), .A1(n1114), .Z(n849));
Q_MX02 U845 ( .S(pipe_ack_num_bytes[2]), .A0(n1147), .A1(n1115), .Z(n850));
Q_MX02 U846 ( .S(pipe_ack_num_bytes[2]), .A0(n1148), .A1(n1116), .Z(n851));
Q_MX02 U847 ( .S(pipe_ack_num_bytes[2]), .A0(n1149), .A1(n1117), .Z(n852));
Q_MX02 U848 ( .S(pipe_ack_num_bytes[2]), .A0(n1150), .A1(n1118), .Z(n853));
Q_MX02 U849 ( .S(pipe_ack_num_bytes[2]), .A0(n1151), .A1(n1119), .Z(n854));
Q_MX02 U850 ( .S(pipe_ack_num_bytes[2]), .A0(n1152), .A1(n1120), .Z(n855));
Q_MX02 U851 ( .S(pipe_ack_num_bytes[2]), .A0(n1153), .A1(n1121), .Z(n856));
Q_MX02 U852 ( .S(pipe_ack_num_bytes[2]), .A0(n1154), .A1(n1122), .Z(n857));
Q_MX02 U853 ( .S(pipe_ack_num_bytes[2]), .A0(n1155), .A1(n1123), .Z(n858));
Q_MX02 U854 ( .S(pipe_ack_num_bytes[2]), .A0(n1156), .A1(n1124), .Z(n859));
Q_MX02 U855 ( .S(pipe_ack_num_bytes[2]), .A0(n1157), .A1(n1125), .Z(n860));
Q_MX02 U856 ( .S(pipe_ack_num_bytes[2]), .A0(n1158), .A1(n1126), .Z(n861));
Q_MX02 U857 ( .S(pipe_ack_num_bytes[2]), .A0(n1159), .A1(n1127), .Z(n862));
Q_MX02 U858 ( .S(pipe_ack_num_bytes[2]), .A0(n1160), .A1(n1128), .Z(n863));
Q_MX02 U859 ( .S(pipe_ack_num_bytes[2]), .A0(n1161), .A1(n1129), .Z(n864));
Q_MX02 U860 ( .S(pipe_ack_num_bytes[2]), .A0(n1162), .A1(n1130), .Z(n865));
Q_MX02 U861 ( .S(pipe_ack_num_bytes[2]), .A0(n1163), .A1(n1131), .Z(n866));
Q_MX02 U862 ( .S(pipe_ack_num_bytes[2]), .A0(n1164), .A1(n1132), .Z(n867));
Q_MX02 U863 ( .S(pipe_ack_num_bytes[2]), .A0(n1165), .A1(n1133), .Z(n868));
Q_MX02 U864 ( .S(pipe_ack_num_bytes[2]), .A0(n1166), .A1(n1134), .Z(n869));
Q_MX02 U865 ( .S(pipe_ack_num_bytes[2]), .A0(n1167), .A1(n1135), .Z(n870));
Q_MX02 U866 ( .S(pipe_ack_num_bytes[2]), .A0(n1168), .A1(n1136), .Z(n871));
Q_MX02 U867 ( .S(pipe_ack_num_bytes[2]), .A0(n1169), .A1(n1137), .Z(n872));
Q_MX02 U868 ( .S(pipe_ack_num_bytes[2]), .A0(n1170), .A1(n1138), .Z(n873));
Q_MX02 U869 ( .S(pipe_ack_num_bytes[2]), .A0(n1171), .A1(n1139), .Z(n874));
Q_MX02 U870 ( .S(pipe_ack_num_bytes[2]), .A0(n1172), .A1(n1140), .Z(n875));
Q_MX02 U871 ( .S(pipe_ack_num_bytes[2]), .A0(n1173), .A1(n1141), .Z(n876));
Q_MX02 U872 ( .S(pipe_ack_num_bytes[2]), .A0(n1174), .A1(n1142), .Z(n877));
Q_MX02 U873 ( .S(pipe_ack_num_bytes[2]), .A0(n1175), .A1(n1143), .Z(n878));
Q_MX02 U874 ( .S(pipe_ack_num_bytes[2]), .A0(n1176), .A1(n1144), .Z(n879));
Q_MX02 U875 ( .S(pipe_ack_num_bytes[2]), .A0(n1177), .A1(n1145), .Z(n880));
Q_MX02 U876 ( .S(pipe_ack_num_bytes[2]), .A0(n1178), .A1(n1146), .Z(n881));
Q_MX02 U877 ( .S(pipe_ack_num_bytes[2]), .A0(n1179), .A1(n1147), .Z(n882));
Q_MX02 U878 ( .S(pipe_ack_num_bytes[2]), .A0(n1180), .A1(n1148), .Z(n883));
Q_MX02 U879 ( .S(pipe_ack_num_bytes[2]), .A0(n1181), .A1(n1149), .Z(n884));
Q_MX02 U880 ( .S(pipe_ack_num_bytes[2]), .A0(n1182), .A1(n1150), .Z(n885));
Q_MX02 U881 ( .S(pipe_ack_num_bytes[2]), .A0(n1183), .A1(n1151), .Z(n886));
Q_MX02 U882 ( .S(pipe_ack_num_bytes[2]), .A0(n1184), .A1(n1152), .Z(n887));
Q_MX02 U883 ( .S(pipe_ack_num_bytes[2]), .A0(n1185), .A1(n1153), .Z(n888));
Q_MX02 U884 ( .S(pipe_ack_num_bytes[2]), .A0(n1186), .A1(n1154), .Z(n889));
Q_MX02 U885 ( .S(pipe_ack_num_bytes[2]), .A0(n1187), .A1(n1155), .Z(n890));
Q_MX02 U886 ( .S(pipe_ack_num_bytes[2]), .A0(n1188), .A1(n1156), .Z(n891));
Q_MX02 U887 ( .S(pipe_ack_num_bytes[2]), .A0(n1189), .A1(n1157), .Z(n892));
Q_MX02 U888 ( .S(pipe_ack_num_bytes[2]), .A0(n1190), .A1(n1158), .Z(n893));
Q_MX02 U889 ( .S(pipe_ack_num_bytes[2]), .A0(n1191), .A1(n1159), .Z(n894));
Q_MX02 U890 ( .S(pipe_ack_num_bytes[2]), .A0(n1192), .A1(n1160), .Z(n895));
Q_MX02 U891 ( .S(pipe_ack_num_bytes[2]), .A0(n1193), .A1(n1161), .Z(n896));
Q_MX02 U892 ( .S(pipe_ack_num_bytes[2]), .A0(n1194), .A1(n1162), .Z(n897));
Q_MX02 U893 ( .S(pipe_ack_num_bytes[2]), .A0(n1195), .A1(n1163), .Z(n898));
Q_MX02 U894 ( .S(pipe_ack_num_bytes[2]), .A0(n1196), .A1(n1164), .Z(n899));
Q_MX02 U895 ( .S(pipe_ack_num_bytes[2]), .A0(n1197), .A1(n1165), .Z(n900));
Q_MX02 U896 ( .S(pipe_ack_num_bytes[2]), .A0(n1198), .A1(n1166), .Z(n901));
Q_MX02 U897 ( .S(pipe_ack_num_bytes[2]), .A0(n1199), .A1(n1167), .Z(n902));
Q_MX02 U898 ( .S(pipe_ack_num_bytes[2]), .A0(n1200), .A1(n1168), .Z(n903));
Q_MX02 U899 ( .S(pipe_ack_num_bytes[2]), .A0(n1201), .A1(n1169), .Z(n904));
Q_MX02 U900 ( .S(pipe_ack_num_bytes[2]), .A0(n1202), .A1(n1170), .Z(n905));
Q_MX02 U901 ( .S(pipe_ack_num_bytes[2]), .A0(n1203), .A1(n1171), .Z(n906));
Q_MX02 U902 ( .S(pipe_ack_num_bytes[2]), .A0(n1204), .A1(n1172), .Z(n907));
Q_MX02 U903 ( .S(pipe_ack_num_bytes[2]), .A0(n1205), .A1(n1173), .Z(n908));
Q_MX02 U904 ( .S(pipe_ack_num_bytes[2]), .A0(n1206), .A1(n1174), .Z(n909));
Q_MX02 U905 ( .S(pipe_ack_num_bytes[2]), .A0(n1207), .A1(n1175), .Z(n910));
Q_MX02 U906 ( .S(pipe_ack_num_bytes[2]), .A0(n1208), .A1(n1176), .Z(n911));
Q_MX02 U907 ( .S(pipe_ack_num_bytes[2]), .A0(n1209), .A1(n1177), .Z(n912));
Q_MX02 U908 ( .S(pipe_ack_num_bytes[2]), .A0(n1210), .A1(n1178), .Z(n913));
Q_MX02 U909 ( .S(pipe_ack_num_bytes[2]), .A0(n1211), .A1(n1179), .Z(n914));
Q_MX02 U910 ( .S(pipe_ack_num_bytes[2]), .A0(n1212), .A1(n1180), .Z(n915));
Q_MX02 U911 ( .S(pipe_ack_num_bytes[2]), .A0(n1213), .A1(n1181), .Z(n916));
Q_MX02 U912 ( .S(pipe_ack_num_bytes[2]), .A0(n1214), .A1(n1182), .Z(n917));
Q_MX02 U913 ( .S(pipe_ack_num_bytes[2]), .A0(n1215), .A1(n1183), .Z(n918));
Q_MX02 U914 ( .S(pipe_ack_num_bytes[2]), .A0(n1216), .A1(n1184), .Z(n919));
Q_MX02 U915 ( .S(pipe_ack_num_bytes[2]), .A0(n1217), .A1(n1185), .Z(n920));
Q_MX02 U916 ( .S(pipe_ack_num_bytes[2]), .A0(n1218), .A1(n1186), .Z(n921));
Q_MX02 U917 ( .S(pipe_ack_num_bytes[2]), .A0(n1219), .A1(n1187), .Z(n922));
Q_MX02 U918 ( .S(pipe_ack_num_bytes[2]), .A0(n1220), .A1(n1188), .Z(n923));
Q_MX02 U919 ( .S(pipe_ack_num_bytes[2]), .A0(n1221), .A1(n1189), .Z(n924));
Q_MX02 U920 ( .S(pipe_ack_num_bytes[2]), .A0(n1222), .A1(n1190), .Z(n925));
Q_MX02 U921 ( .S(pipe_ack_num_bytes[2]), .A0(n1223), .A1(n1191), .Z(n926));
Q_MX02 U922 ( .S(pipe_ack_num_bytes[2]), .A0(n1224), .A1(n1192), .Z(n927));
Q_MX02 U923 ( .S(pipe_ack_num_bytes[2]), .A0(n1225), .A1(n1193), .Z(n928));
Q_MX02 U924 ( .S(pipe_ack_num_bytes[2]), .A0(n1226), .A1(n1194), .Z(n929));
Q_MX02 U925 ( .S(pipe_ack_num_bytes[2]), .A0(n1227), .A1(n1195), .Z(n930));
Q_MX02 U926 ( .S(pipe_ack_num_bytes[2]), .A0(n1228), .A1(n1196), .Z(n931));
Q_MX02 U927 ( .S(pipe_ack_num_bytes[2]), .A0(n1229), .A1(n1197), .Z(n932));
Q_MX02 U928 ( .S(pipe_ack_num_bytes[2]), .A0(n1230), .A1(n1198), .Z(n933));
Q_MX02 U929 ( .S(pipe_ack_num_bytes[2]), .A0(n1231), .A1(n1199), .Z(n934));
Q_MX02 U930 ( .S(pipe_ack_num_bytes[2]), .A0(n1232), .A1(n1200), .Z(n935));
Q_MX02 U931 ( .S(pipe_ack_num_bytes[2]), .A0(n1233), .A1(n1201), .Z(n936));
Q_MX02 U932 ( .S(pipe_ack_num_bytes[2]), .A0(n1234), .A1(n1202), .Z(n937));
Q_MX02 U933 ( .S(pipe_ack_num_bytes[2]), .A0(n1235), .A1(n1203), .Z(n938));
Q_MX02 U934 ( .S(pipe_ack_num_bytes[2]), .A0(n1236), .A1(n1204), .Z(n939));
Q_MX02 U935 ( .S(pipe_ack_num_bytes[2]), .A0(n1237), .A1(n1205), .Z(n940));
Q_MX02 U936 ( .S(pipe_ack_num_bytes[2]), .A0(n1238), .A1(n1206), .Z(n941));
Q_MX02 U937 ( .S(pipe_ack_num_bytes[2]), .A0(n1239), .A1(n1207), .Z(n942));
Q_MX02 U938 ( .S(pipe_ack_num_bytes[2]), .A0(n1240), .A1(n1208), .Z(n943));
Q_MX02 U939 ( .S(pipe_ack_num_bytes[2]), .A0(n1241), .A1(n1209), .Z(n944));
Q_MX02 U940 ( .S(pipe_ack_num_bytes[2]), .A0(n1242), .A1(n1210), .Z(n945));
Q_MX02 U941 ( .S(pipe_ack_num_bytes[2]), .A0(n1243), .A1(n1211), .Z(n946));
Q_MX02 U942 ( .S(pipe_ack_num_bytes[2]), .A0(n1244), .A1(n1212), .Z(n947));
Q_MX02 U943 ( .S(pipe_ack_num_bytes[2]), .A0(n1245), .A1(n1213), .Z(n948));
Q_MX02 U944 ( .S(pipe_ack_num_bytes[2]), .A0(n1246), .A1(n1214), .Z(n949));
Q_MX02 U945 ( .S(pipe_ack_num_bytes[2]), .A0(n1247), .A1(n1215), .Z(n950));
Q_MX02 U946 ( .S(pipe_ack_num_bytes[2]), .A0(n1248), .A1(n1216), .Z(n951));
Q_MX02 U947 ( .S(pipe_ack_num_bytes[2]), .A0(n1249), .A1(n1217), .Z(n952));
Q_MX02 U948 ( .S(pipe_ack_num_bytes[2]), .A0(n1250), .A1(n1218), .Z(n953));
Q_MX02 U949 ( .S(pipe_ack_num_bytes[2]), .A0(n1251), .A1(n1219), .Z(n954));
Q_MX02 U950 ( .S(pipe_ack_num_bytes[2]), .A0(n1252), .A1(n1220), .Z(n955));
Q_MX02 U951 ( .S(pipe_ack_num_bytes[2]), .A0(n1253), .A1(n1221), .Z(n956));
Q_MX02 U952 ( .S(pipe_ack_num_bytes[2]), .A0(n1254), .A1(n1222), .Z(n957));
Q_MX02 U953 ( .S(pipe_ack_num_bytes[2]), .A0(n1255), .A1(n1223), .Z(n958));
Q_MX02 U954 ( .S(pipe_ack_num_bytes[2]), .A0(n1256), .A1(n1224), .Z(n959));
Q_MX02 U955 ( .S(pipe_ack_num_bytes[2]), .A0(n1257), .A1(n1225), .Z(n960));
Q_MX02 U956 ( .S(pipe_ack_num_bytes[2]), .A0(n1258), .A1(n1226), .Z(n961));
Q_MX02 U957 ( .S(pipe_ack_num_bytes[2]), .A0(n1259), .A1(n1227), .Z(n962));
Q_MX02 U958 ( .S(pipe_ack_num_bytes[2]), .A0(n1260), .A1(n1228), .Z(n963));
Q_MX02 U959 ( .S(pipe_ack_num_bytes[2]), .A0(n1261), .A1(n1229), .Z(n964));
Q_MX02 U960 ( .S(pipe_ack_num_bytes[2]), .A0(n1262), .A1(n1230), .Z(n965));
Q_MX02 U961 ( .S(pipe_ack_num_bytes[2]), .A0(n1263), .A1(n1231), .Z(n966));
Q_MX02 U962 ( .S(pipe_ack_num_bytes[2]), .A0(n1264), .A1(n1232), .Z(n967));
Q_MX02 U963 ( .S(pipe_ack_num_bytes[2]), .A0(n1265), .A1(n1233), .Z(n968));
Q_MX02 U964 ( .S(pipe_ack_num_bytes[2]), .A0(n1266), .A1(n1234), .Z(n969));
Q_MX02 U965 ( .S(pipe_ack_num_bytes[2]), .A0(n1267), .A1(n1235), .Z(n970));
Q_MX02 U966 ( .S(pipe_ack_num_bytes[2]), .A0(n1268), .A1(n1236), .Z(n971));
Q_MX02 U967 ( .S(pipe_ack_num_bytes[2]), .A0(n1269), .A1(n1237), .Z(n972));
Q_MX02 U968 ( .S(pipe_ack_num_bytes[2]), .A0(n1270), .A1(n1238), .Z(n973));
Q_MX02 U969 ( .S(pipe_ack_num_bytes[2]), .A0(n1271), .A1(n1239), .Z(n974));
Q_MX02 U970 ( .S(pipe_ack_num_bytes[2]), .A0(n1272), .A1(n1240), .Z(n975));
Q_MX02 U971 ( .S(pipe_ack_num_bytes[2]), .A0(n1273), .A1(n1241), .Z(n976));
Q_MX02 U972 ( .S(pipe_ack_num_bytes[2]), .A0(n1274), .A1(n1242), .Z(n977));
Q_MX02 U973 ( .S(pipe_ack_num_bytes[2]), .A0(n1275), .A1(n1243), .Z(n978));
Q_MX02 U974 ( .S(pipe_ack_num_bytes[2]), .A0(n1276), .A1(n1244), .Z(n979));
Q_MX02 U975 ( .S(pipe_ack_num_bytes[2]), .A0(n1277), .A1(n1245), .Z(n980));
Q_MX02 U976 ( .S(pipe_ack_num_bytes[2]), .A0(n1278), .A1(n1246), .Z(n981));
Q_MX02 U977 ( .S(pipe_ack_num_bytes[2]), .A0(n1279), .A1(n1247), .Z(n982));
Q_MX02 U978 ( .S(pipe_ack_num_bytes[2]), .A0(n1280), .A1(n1248), .Z(n983));
Q_MX02 U979 ( .S(pipe_ack_num_bytes[2]), .A0(n1281), .A1(n1249), .Z(n984));
Q_MX02 U980 ( .S(pipe_ack_num_bytes[2]), .A0(n1282), .A1(n1250), .Z(n985));
Q_MX02 U981 ( .S(pipe_ack_num_bytes[2]), .A0(n1283), .A1(n1251), .Z(n986));
Q_MX02 U982 ( .S(pipe_ack_num_bytes[2]), .A0(n1284), .A1(n1252), .Z(n987));
Q_MX02 U983 ( .S(pipe_ack_num_bytes[2]), .A0(n1285), .A1(n1253), .Z(n988));
Q_MX02 U984 ( .S(pipe_ack_num_bytes[2]), .A0(n1286), .A1(n1254), .Z(n989));
Q_MX02 U985 ( .S(pipe_ack_num_bytes[2]), .A0(n1287), .A1(n1255), .Z(n990));
Q_MX02 U986 ( .S(pipe_ack_num_bytes[2]), .A0(n1288), .A1(n1256), .Z(n991));
Q_MX02 U987 ( .S(pipe_ack_num_bytes[2]), .A0(n1289), .A1(n1257), .Z(n992));
Q_MX02 U988 ( .S(pipe_ack_num_bytes[2]), .A0(n1290), .A1(n1258), .Z(n993));
Q_MX02 U989 ( .S(pipe_ack_num_bytes[2]), .A0(n1291), .A1(n1259), .Z(n994));
Q_MX02 U990 ( .S(pipe_ack_num_bytes[2]), .A0(n1292), .A1(n1260), .Z(n995));
Q_MX02 U991 ( .S(pipe_ack_num_bytes[2]), .A0(n1293), .A1(n1261), .Z(n996));
Q_MX02 U992 ( .S(pipe_ack_num_bytes[2]), .A0(n1294), .A1(n1262), .Z(n997));
Q_MX02 U993 ( .S(pipe_ack_num_bytes[2]), .A0(n1295), .A1(n1263), .Z(n998));
Q_MX02 U994 ( .S(pipe_ack_num_bytes[2]), .A0(n1296), .A1(n1264), .Z(n999));
Q_MX02 U995 ( .S(pipe_ack_num_bytes[2]), .A0(n1297), .A1(n1265), .Z(n1000));
Q_MX02 U996 ( .S(pipe_ack_num_bytes[2]), .A0(n1298), .A1(n1266), .Z(n1001));
Q_MX02 U997 ( .S(pipe_ack_num_bytes[2]), .A0(n1299), .A1(n1267), .Z(n1002));
Q_MX02 U998 ( .S(pipe_ack_num_bytes[2]), .A0(n1300), .A1(n1268), .Z(n1003));
Q_MX02 U999 ( .S(pipe_ack_num_bytes[2]), .A0(n1301), .A1(n1269), .Z(n1004));
Q_MX02 U1000 ( .S(pipe_ack_num_bytes[2]), .A0(n1302), .A1(n1270), .Z(n1005));
Q_MX02 U1001 ( .S(pipe_ack_num_bytes[2]), .A0(n1303), .A1(n1271), .Z(n1006));
Q_MX02 U1002 ( .S(pipe_ack_num_bytes[2]), .A0(n1304), .A1(n1272), .Z(n1007));
Q_MX02 U1003 ( .S(pipe_ack_num_bytes[2]), .A0(n1305), .A1(n1273), .Z(n1008));
Q_MX02 U1004 ( .S(pipe_ack_num_bytes[2]), .A0(n1306), .A1(n1274), .Z(n1009));
Q_MX02 U1005 ( .S(pipe_ack_num_bytes[2]), .A0(n1307), .A1(n1275), .Z(n1010));
Q_MX02 U1006 ( .S(pipe_ack_num_bytes[2]), .A0(n1308), .A1(n1276), .Z(n1011));
Q_MX02 U1007 ( .S(pipe_ack_num_bytes[2]), .A0(n1309), .A1(n1277), .Z(n1012));
Q_MX02 U1008 ( .S(pipe_ack_num_bytes[2]), .A0(n1310), .A1(n1278), .Z(n1013));
Q_MX02 U1009 ( .S(pipe_ack_num_bytes[2]), .A0(n1311), .A1(n1279), .Z(n1014));
Q_MX02 U1010 ( .S(pipe_ack_num_bytes[2]), .A0(n1312), .A1(n1280), .Z(n1015));
Q_MX02 U1011 ( .S(pipe_ack_num_bytes[2]), .A0(n1313), .A1(n1281), .Z(n1016));
Q_MX02 U1012 ( .S(pipe_ack_num_bytes[2]), .A0(n1314), .A1(n1282), .Z(n1017));
Q_MX02 U1013 ( .S(pipe_ack_num_bytes[2]), .A0(n1315), .A1(n1283), .Z(n1018));
Q_MX02 U1014 ( .S(pipe_ack_num_bytes[2]), .A0(n1316), .A1(n1284), .Z(n1019));
Q_MX02 U1015 ( .S(pipe_ack_num_bytes[2]), .A0(n1317), .A1(n1285), .Z(n1020));
Q_MX02 U1016 ( .S(pipe_ack_num_bytes[2]), .A0(n1318), .A1(n1286), .Z(n1021));
Q_MX02 U1017 ( .S(pipe_ack_num_bytes[2]), .A0(n1319), .A1(n1287), .Z(n1022));
Q_MX02 U1018 ( .S(pipe_ack_num_bytes[2]), .A0(n1320), .A1(n1288), .Z(n1023));
Q_MX02 U1019 ( .S(pipe_ack_num_bytes[2]), .A0(n1321), .A1(n1289), .Z(n1024));
Q_MX02 U1020 ( .S(pipe_ack_num_bytes[2]), .A0(n1322), .A1(n1290), .Z(n1025));
Q_MX02 U1021 ( .S(pipe_ack_num_bytes[2]), .A0(n1323), .A1(n1291), .Z(n1026));
Q_MX02 U1022 ( .S(pipe_ack_num_bytes[2]), .A0(n1324), .A1(n1292), .Z(n1027));
Q_MX02 U1023 ( .S(pipe_ack_num_bytes[2]), .A0(n1325), .A1(n1293), .Z(n1028));
Q_MX02 U1024 ( .S(pipe_ack_num_bytes[2]), .A0(n1326), .A1(n1294), .Z(n1029));
Q_MX02 U1025 ( .S(pipe_ack_num_bytes[2]), .A0(n1327), .A1(n1295), .Z(n1030));
Q_MX02 U1026 ( .S(pipe_ack_num_bytes[2]), .A0(n1328), .A1(n1296), .Z(n1031));
Q_MX02 U1027 ( .S(pipe_ack_num_bytes[2]), .A0(n1329), .A1(n1297), .Z(n1032));
Q_MX02 U1028 ( .S(pipe_ack_num_bytes[2]), .A0(n1330), .A1(n1298), .Z(n1033));
Q_MX02 U1029 ( .S(pipe_ack_num_bytes[2]), .A0(n1331), .A1(n1299), .Z(n1034));
Q_MX02 U1030 ( .S(pipe_ack_num_bytes[2]), .A0(n1332), .A1(n1300), .Z(n1035));
Q_MX02 U1031 ( .S(pipe_ack_num_bytes[2]), .A0(n1333), .A1(n1301), .Z(n1036));
Q_MX02 U1032 ( .S(pipe_ack_num_bytes[2]), .A0(n1334), .A1(n1302), .Z(n1037));
Q_MX02 U1033 ( .S(pipe_ack_num_bytes[2]), .A0(n1335), .A1(n1303), .Z(n1038));
Q_MX02 U1034 ( .S(pipe_ack_num_bytes[2]), .A0(n1336), .A1(n1304), .Z(n1039));
Q_MX02 U1035 ( .S(pipe_ack_num_bytes[2]), .A0(n1337), .A1(n1305), .Z(n1040));
Q_MX02 U1036 ( .S(pipe_ack_num_bytes[2]), .A0(n1338), .A1(n1306), .Z(n1041));
Q_MX02 U1037 ( .S(pipe_ack_num_bytes[2]), .A0(n1339), .A1(n1307), .Z(n1042));
Q_MX02 U1038 ( .S(pipe_ack_num_bytes[2]), .A0(n1340), .A1(n1308), .Z(n1043));
Q_MX02 U1039 ( .S(pipe_ack_num_bytes[2]), .A0(n1341), .A1(n1309), .Z(n1044));
Q_MX02 U1040 ( .S(pipe_ack_num_bytes[2]), .A0(n1342), .A1(n1310), .Z(n1045));
Q_MX03 U1041 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1608), .A1(n1592), .A2(n1311), .Z(n1046));
Q_MX03 U1042 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1609), .A1(n1593), .A2(n1312), .Z(n1047));
Q_MX03 U1043 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1610), .A1(n1594), .A2(n1313), .Z(n1048));
Q_MX03 U1044 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1611), .A1(n1595), .A2(n1314), .Z(n1049));
Q_MX03 U1045 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1612), .A1(n1596), .A2(n1315), .Z(n1050));
Q_MX03 U1046 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1613), .A1(n1597), .A2(n1316), .Z(n1051));
Q_MX03 U1047 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1614), .A1(n1598), .A2(n1317), .Z(n1052));
Q_MX03 U1048 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1615), .A1(n1599), .A2(n1318), .Z(n1053));
Q_MX03 U1049 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1616), .A1(n1600), .A2(n1319), .Z(n1054));
Q_MX03 U1050 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1617), .A1(n1601), .A2(n1320), .Z(n1055));
Q_MX03 U1051 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1618), .A1(n1602), .A2(n1321), .Z(n1056));
Q_MX03 U1052 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1619), .A1(n1603), .A2(n1322), .Z(n1057));
Q_MX03 U1053 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1620), .A1(n1604), .A2(n1323), .Z(n1058));
Q_MX03 U1054 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1621), .A1(n1605), .A2(n1324), .Z(n1059));
Q_MX03 U1055 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1622), .A1(n1606), .A2(n1325), .Z(n1060));
Q_MX03 U1056 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1623), .A1(n1607), .A2(n1326), .Z(n1061));
Q_MX03 U1057 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1624), .A1(n1608), .A2(n1327), .Z(n1062));
Q_MX03 U1058 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1625), .A1(n1609), .A2(n1328), .Z(n1063));
Q_MX03 U1059 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1626), .A1(n1610), .A2(n1329), .Z(n1064));
Q_MX03 U1060 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1627), .A1(n1611), .A2(n1330), .Z(n1065));
Q_MX03 U1061 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1628), .A1(n1612), .A2(n1331), .Z(n1066));
Q_MX03 U1062 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1629), .A1(n1613), .A2(n1332), .Z(n1067));
Q_MX03 U1063 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1630), .A1(n1614), .A2(n1333), .Z(n1068));
Q_MX03 U1064 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1631), .A1(n1615), .A2(n1334), .Z(n1069));
Q_MX03 U1065 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1632), .A1(n1616), .A2(n1335), .Z(n1070));
Q_MX03 U1066 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1633), .A1(n1617), .A2(n1336), .Z(n1071));
Q_MX03 U1067 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1634), .A1(n1618), .A2(n1337), .Z(n1072));
Q_MX03 U1068 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1635), .A1(n1619), .A2(n1338), .Z(n1073));
Q_MX03 U1069 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1636), .A1(n1620), .A2(n1339), .Z(n1074));
Q_MX03 U1070 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1637), .A1(n1621), .A2(n1340), .Z(n1075));
Q_MX03 U1071 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1638), .A1(n1622), .A2(n1341), .Z(n1076));
Q_MX03 U1072 ( .S0(pipe_ack_num_bytes[1]), .S1(pipe_ack_num_bytes[2]), .A0(n1639), .A1(n1623), .A2(n1342), .Z(n1077));
Q_AN02 U1073 ( .A0(n1094), .A1(n1343), .Z(n1078));
Q_AN02 U1074 ( .A0(n1094), .A1(n1344), .Z(n1079));
Q_AN02 U1075 ( .A0(n1094), .A1(n1345), .Z(n1080));
Q_AN02 U1076 ( .A0(n1094), .A1(n1346), .Z(n1081));
Q_AN02 U1077 ( .A0(n1094), .A1(n1347), .Z(n1082));
Q_AN02 U1078 ( .A0(n1094), .A1(n1348), .Z(n1083));
Q_AN02 U1079 ( .A0(n1094), .A1(n1349), .Z(n1084));
Q_AN02 U1080 ( .A0(n1094), .A1(n1350), .Z(n1085));
Q_AN02 U1081 ( .A0(n1094), .A1(n1352), .Z(n1086));
Q_AN02 U1082 ( .A0(n1094), .A1(n1353), .Z(n1087));
Q_AN02 U1083 ( .A0(n1094), .A1(n1354), .Z(n1088));
Q_AN02 U1084 ( .A0(n1094), .A1(n1355), .Z(n1089));
Q_AN02 U1085 ( .A0(n1094), .A1(n1356), .Z(n1090));
Q_AN02 U1086 ( .A0(n1094), .A1(n1357), .Z(n1091));
Q_AN02 U1087 ( .A0(n1094), .A1(n1358), .Z(n1092));
Q_AN02 U1088 ( .A0(n1094), .A1(n1359), .Z(n1093));
Q_INV U1089 ( .A(pipe_ack_num_bytes[1]), .Z(n1094));
Q_MX02 U1090 ( .S(pipe_ack_num_bytes[1]), .A0(n1360), .A1(n1343), .Z(n1095));
Q_MX02 U1091 ( .S(pipe_ack_num_bytes[1]), .A0(n1361), .A1(n1344), .Z(n1096));
Q_MX02 U1092 ( .S(pipe_ack_num_bytes[1]), .A0(n1362), .A1(n1345), .Z(n1097));
Q_MX02 U1093 ( .S(pipe_ack_num_bytes[1]), .A0(n1363), .A1(n1346), .Z(n1098));
Q_MX02 U1094 ( .S(pipe_ack_num_bytes[1]), .A0(n1364), .A1(n1347), .Z(n1099));
Q_MX02 U1095 ( .S(pipe_ack_num_bytes[1]), .A0(n1365), .A1(n1348), .Z(n1100));
Q_MX02 U1096 ( .S(pipe_ack_num_bytes[1]), .A0(n1366), .A1(n1349), .Z(n1101));
Q_MX02 U1097 ( .S(pipe_ack_num_bytes[1]), .A0(n1367), .A1(n1350), .Z(n1102));
Q_MX02 U1098 ( .S(pipe_ack_num_bytes[1]), .A0(n1368), .A1(n1352), .Z(n1103));
Q_MX02 U1099 ( .S(pipe_ack_num_bytes[1]), .A0(n1369), .A1(n1353), .Z(n1104));
Q_MX02 U1100 ( .S(pipe_ack_num_bytes[1]), .A0(n1370), .A1(n1354), .Z(n1105));
Q_MX02 U1101 ( .S(pipe_ack_num_bytes[1]), .A0(n1371), .A1(n1355), .Z(n1106));
Q_MX02 U1102 ( .S(pipe_ack_num_bytes[1]), .A0(n1372), .A1(n1356), .Z(n1107));
Q_MX02 U1103 ( .S(pipe_ack_num_bytes[1]), .A0(n1373), .A1(n1357), .Z(n1108));
Q_MX02 U1104 ( .S(pipe_ack_num_bytes[1]), .A0(n1374), .A1(n1358), .Z(n1109));
Q_MX02 U1105 ( .S(pipe_ack_num_bytes[1]), .A0(n1375), .A1(n1359), .Z(n1110));
Q_MX02 U1106 ( .S(pipe_ack_num_bytes[1]), .A0(n1376), .A1(n1360), .Z(n1111));
Q_MX02 U1107 ( .S(pipe_ack_num_bytes[1]), .A0(n1377), .A1(n1361), .Z(n1112));
Q_MX02 U1108 ( .S(pipe_ack_num_bytes[1]), .A0(n1378), .A1(n1362), .Z(n1113));
Q_MX02 U1109 ( .S(pipe_ack_num_bytes[1]), .A0(n1379), .A1(n1363), .Z(n1114));
Q_MX02 U1110 ( .S(pipe_ack_num_bytes[1]), .A0(n1380), .A1(n1364), .Z(n1115));
Q_MX02 U1111 ( .S(pipe_ack_num_bytes[1]), .A0(n1381), .A1(n1365), .Z(n1116));
Q_MX02 U1112 ( .S(pipe_ack_num_bytes[1]), .A0(n1382), .A1(n1366), .Z(n1117));
Q_MX02 U1113 ( .S(pipe_ack_num_bytes[1]), .A0(n1383), .A1(n1367), .Z(n1118));
Q_MX02 U1114 ( .S(pipe_ack_num_bytes[1]), .A0(n1384), .A1(n1368), .Z(n1119));
Q_MX02 U1115 ( .S(pipe_ack_num_bytes[1]), .A0(n1385), .A1(n1369), .Z(n1120));
Q_MX02 U1116 ( .S(pipe_ack_num_bytes[1]), .A0(n1386), .A1(n1370), .Z(n1121));
Q_MX02 U1117 ( .S(pipe_ack_num_bytes[1]), .A0(n1387), .A1(n1371), .Z(n1122));
Q_MX02 U1118 ( .S(pipe_ack_num_bytes[1]), .A0(n1388), .A1(n1372), .Z(n1123));
Q_MX02 U1119 ( .S(pipe_ack_num_bytes[1]), .A0(n1389), .A1(n1373), .Z(n1124));
Q_MX02 U1120 ( .S(pipe_ack_num_bytes[1]), .A0(n1390), .A1(n1374), .Z(n1125));
Q_MX02 U1121 ( .S(pipe_ack_num_bytes[1]), .A0(n1391), .A1(n1375), .Z(n1126));
Q_MX02 U1122 ( .S(pipe_ack_num_bytes[1]), .A0(n1392), .A1(n1376), .Z(n1127));
Q_MX02 U1123 ( .S(pipe_ack_num_bytes[1]), .A0(n1393), .A1(n1377), .Z(n1128));
Q_MX02 U1124 ( .S(pipe_ack_num_bytes[1]), .A0(n1394), .A1(n1378), .Z(n1129));
Q_MX02 U1125 ( .S(pipe_ack_num_bytes[1]), .A0(n1395), .A1(n1379), .Z(n1130));
Q_MX02 U1126 ( .S(pipe_ack_num_bytes[1]), .A0(n1396), .A1(n1380), .Z(n1131));
Q_MX02 U1127 ( .S(pipe_ack_num_bytes[1]), .A0(n1397), .A1(n1381), .Z(n1132));
Q_MX02 U1128 ( .S(pipe_ack_num_bytes[1]), .A0(n1398), .A1(n1382), .Z(n1133));
Q_MX02 U1129 ( .S(pipe_ack_num_bytes[1]), .A0(n1399), .A1(n1383), .Z(n1134));
Q_MX02 U1130 ( .S(pipe_ack_num_bytes[1]), .A0(n1400), .A1(n1384), .Z(n1135));
Q_MX02 U1131 ( .S(pipe_ack_num_bytes[1]), .A0(n1401), .A1(n1385), .Z(n1136));
Q_MX02 U1132 ( .S(pipe_ack_num_bytes[1]), .A0(n1402), .A1(n1386), .Z(n1137));
Q_MX02 U1133 ( .S(pipe_ack_num_bytes[1]), .A0(n1403), .A1(n1387), .Z(n1138));
Q_MX02 U1134 ( .S(pipe_ack_num_bytes[1]), .A0(n1404), .A1(n1388), .Z(n1139));
Q_MX02 U1135 ( .S(pipe_ack_num_bytes[1]), .A0(n1405), .A1(n1389), .Z(n1140));
Q_MX02 U1136 ( .S(pipe_ack_num_bytes[1]), .A0(n1406), .A1(n1390), .Z(n1141));
Q_MX02 U1137 ( .S(pipe_ack_num_bytes[1]), .A0(n1407), .A1(n1391), .Z(n1142));
Q_MX02 U1138 ( .S(pipe_ack_num_bytes[1]), .A0(n1408), .A1(n1392), .Z(n1143));
Q_MX02 U1139 ( .S(pipe_ack_num_bytes[1]), .A0(n1409), .A1(n1393), .Z(n1144));
Q_MX02 U1140 ( .S(pipe_ack_num_bytes[1]), .A0(n1410), .A1(n1394), .Z(n1145));
Q_MX02 U1141 ( .S(pipe_ack_num_bytes[1]), .A0(n1411), .A1(n1395), .Z(n1146));
Q_MX02 U1142 ( .S(pipe_ack_num_bytes[1]), .A0(n1412), .A1(n1396), .Z(n1147));
Q_MX02 U1143 ( .S(pipe_ack_num_bytes[1]), .A0(n1413), .A1(n1397), .Z(n1148));
Q_MX02 U1144 ( .S(pipe_ack_num_bytes[1]), .A0(n1414), .A1(n1398), .Z(n1149));
Q_MX02 U1145 ( .S(pipe_ack_num_bytes[1]), .A0(n1415), .A1(n1399), .Z(n1150));
Q_MX02 U1146 ( .S(pipe_ack_num_bytes[1]), .A0(n1416), .A1(n1400), .Z(n1151));
Q_MX02 U1147 ( .S(pipe_ack_num_bytes[1]), .A0(n1417), .A1(n1401), .Z(n1152));
Q_MX02 U1148 ( .S(pipe_ack_num_bytes[1]), .A0(n1418), .A1(n1402), .Z(n1153));
Q_MX02 U1149 ( .S(pipe_ack_num_bytes[1]), .A0(n1419), .A1(n1403), .Z(n1154));
Q_MX02 U1150 ( .S(pipe_ack_num_bytes[1]), .A0(n1420), .A1(n1404), .Z(n1155));
Q_MX02 U1151 ( .S(pipe_ack_num_bytes[1]), .A0(n1421), .A1(n1405), .Z(n1156));
Q_MX02 U1152 ( .S(pipe_ack_num_bytes[1]), .A0(n1422), .A1(n1406), .Z(n1157));
Q_MX02 U1153 ( .S(pipe_ack_num_bytes[1]), .A0(n1423), .A1(n1407), .Z(n1158));
Q_MX02 U1154 ( .S(pipe_ack_num_bytes[1]), .A0(n1424), .A1(n1408), .Z(n1159));
Q_MX02 U1155 ( .S(pipe_ack_num_bytes[1]), .A0(n1425), .A1(n1409), .Z(n1160));
Q_MX02 U1156 ( .S(pipe_ack_num_bytes[1]), .A0(n1426), .A1(n1410), .Z(n1161));
Q_MX02 U1157 ( .S(pipe_ack_num_bytes[1]), .A0(n1427), .A1(n1411), .Z(n1162));
Q_MX02 U1158 ( .S(pipe_ack_num_bytes[1]), .A0(n1428), .A1(n1412), .Z(n1163));
Q_MX02 U1159 ( .S(pipe_ack_num_bytes[1]), .A0(n1429), .A1(n1413), .Z(n1164));
Q_MX02 U1160 ( .S(pipe_ack_num_bytes[1]), .A0(n1430), .A1(n1414), .Z(n1165));
Q_MX02 U1161 ( .S(pipe_ack_num_bytes[1]), .A0(n1431), .A1(n1415), .Z(n1166));
Q_MX02 U1162 ( .S(pipe_ack_num_bytes[1]), .A0(n1432), .A1(n1416), .Z(n1167));
Q_MX02 U1163 ( .S(pipe_ack_num_bytes[1]), .A0(n1433), .A1(n1417), .Z(n1168));
Q_MX02 U1164 ( .S(pipe_ack_num_bytes[1]), .A0(n1434), .A1(n1418), .Z(n1169));
Q_MX02 U1165 ( .S(pipe_ack_num_bytes[1]), .A0(n1435), .A1(n1419), .Z(n1170));
Q_MX02 U1166 ( .S(pipe_ack_num_bytes[1]), .A0(n1436), .A1(n1420), .Z(n1171));
Q_MX02 U1167 ( .S(pipe_ack_num_bytes[1]), .A0(n1437), .A1(n1421), .Z(n1172));
Q_MX02 U1168 ( .S(pipe_ack_num_bytes[1]), .A0(n1438), .A1(n1422), .Z(n1173));
Q_MX02 U1169 ( .S(pipe_ack_num_bytes[1]), .A0(n1439), .A1(n1423), .Z(n1174));
Q_MX02 U1170 ( .S(pipe_ack_num_bytes[1]), .A0(n1440), .A1(n1424), .Z(n1175));
Q_MX02 U1171 ( .S(pipe_ack_num_bytes[1]), .A0(n1441), .A1(n1425), .Z(n1176));
Q_MX02 U1172 ( .S(pipe_ack_num_bytes[1]), .A0(n1442), .A1(n1426), .Z(n1177));
Q_MX02 U1173 ( .S(pipe_ack_num_bytes[1]), .A0(n1443), .A1(n1427), .Z(n1178));
Q_MX02 U1174 ( .S(pipe_ack_num_bytes[1]), .A0(n1444), .A1(n1428), .Z(n1179));
Q_MX02 U1175 ( .S(pipe_ack_num_bytes[1]), .A0(n1445), .A1(n1429), .Z(n1180));
Q_MX02 U1176 ( .S(pipe_ack_num_bytes[1]), .A0(n1446), .A1(n1430), .Z(n1181));
Q_MX02 U1177 ( .S(pipe_ack_num_bytes[1]), .A0(n1447), .A1(n1431), .Z(n1182));
Q_MX02 U1178 ( .S(pipe_ack_num_bytes[1]), .A0(n1448), .A1(n1432), .Z(n1183));
Q_MX02 U1179 ( .S(pipe_ack_num_bytes[1]), .A0(n1449), .A1(n1433), .Z(n1184));
Q_MX02 U1180 ( .S(pipe_ack_num_bytes[1]), .A0(n1450), .A1(n1434), .Z(n1185));
Q_MX02 U1181 ( .S(pipe_ack_num_bytes[1]), .A0(n1451), .A1(n1435), .Z(n1186));
Q_MX02 U1182 ( .S(pipe_ack_num_bytes[1]), .A0(n1452), .A1(n1436), .Z(n1187));
Q_MX02 U1183 ( .S(pipe_ack_num_bytes[1]), .A0(n1453), .A1(n1437), .Z(n1188));
Q_MX02 U1184 ( .S(pipe_ack_num_bytes[1]), .A0(n1454), .A1(n1438), .Z(n1189));
Q_MX02 U1185 ( .S(pipe_ack_num_bytes[1]), .A0(n1455), .A1(n1439), .Z(n1190));
Q_MX02 U1186 ( .S(pipe_ack_num_bytes[1]), .A0(n1456), .A1(n1440), .Z(n1191));
Q_MX02 U1187 ( .S(pipe_ack_num_bytes[1]), .A0(n1457), .A1(n1441), .Z(n1192));
Q_MX02 U1188 ( .S(pipe_ack_num_bytes[1]), .A0(n1458), .A1(n1442), .Z(n1193));
Q_MX02 U1189 ( .S(pipe_ack_num_bytes[1]), .A0(n1459), .A1(n1443), .Z(n1194));
Q_MX02 U1190 ( .S(pipe_ack_num_bytes[1]), .A0(n1460), .A1(n1444), .Z(n1195));
Q_MX02 U1191 ( .S(pipe_ack_num_bytes[1]), .A0(n1461), .A1(n1445), .Z(n1196));
Q_MX02 U1192 ( .S(pipe_ack_num_bytes[1]), .A0(n1462), .A1(n1446), .Z(n1197));
Q_MX02 U1193 ( .S(pipe_ack_num_bytes[1]), .A0(n1463), .A1(n1447), .Z(n1198));
Q_MX02 U1194 ( .S(pipe_ack_num_bytes[1]), .A0(n1464), .A1(n1448), .Z(n1199));
Q_MX02 U1195 ( .S(pipe_ack_num_bytes[1]), .A0(n1465), .A1(n1449), .Z(n1200));
Q_MX02 U1196 ( .S(pipe_ack_num_bytes[1]), .A0(n1466), .A1(n1450), .Z(n1201));
Q_MX02 U1197 ( .S(pipe_ack_num_bytes[1]), .A0(n1467), .A1(n1451), .Z(n1202));
Q_MX02 U1198 ( .S(pipe_ack_num_bytes[1]), .A0(n1468), .A1(n1452), .Z(n1203));
Q_MX02 U1199 ( .S(pipe_ack_num_bytes[1]), .A0(n1469), .A1(n1453), .Z(n1204));
Q_MX02 U1200 ( .S(pipe_ack_num_bytes[1]), .A0(n1470), .A1(n1454), .Z(n1205));
Q_MX02 U1201 ( .S(pipe_ack_num_bytes[1]), .A0(n1471), .A1(n1455), .Z(n1206));
Q_MX02 U1202 ( .S(pipe_ack_num_bytes[1]), .A0(n1472), .A1(n1456), .Z(n1207));
Q_MX02 U1203 ( .S(pipe_ack_num_bytes[1]), .A0(n1473), .A1(n1457), .Z(n1208));
Q_MX02 U1204 ( .S(pipe_ack_num_bytes[1]), .A0(n1474), .A1(n1458), .Z(n1209));
Q_MX02 U1205 ( .S(pipe_ack_num_bytes[1]), .A0(n1475), .A1(n1459), .Z(n1210));
Q_MX02 U1206 ( .S(pipe_ack_num_bytes[1]), .A0(n1476), .A1(n1460), .Z(n1211));
Q_MX02 U1207 ( .S(pipe_ack_num_bytes[1]), .A0(n1477), .A1(n1461), .Z(n1212));
Q_MX02 U1208 ( .S(pipe_ack_num_bytes[1]), .A0(n1478), .A1(n1462), .Z(n1213));
Q_MX02 U1209 ( .S(pipe_ack_num_bytes[1]), .A0(n1479), .A1(n1463), .Z(n1214));
Q_MX02 U1210 ( .S(pipe_ack_num_bytes[1]), .A0(n1480), .A1(n1464), .Z(n1215));
Q_MX02 U1211 ( .S(pipe_ack_num_bytes[1]), .A0(n1481), .A1(n1465), .Z(n1216));
Q_MX02 U1212 ( .S(pipe_ack_num_bytes[1]), .A0(n1482), .A1(n1466), .Z(n1217));
Q_MX02 U1213 ( .S(pipe_ack_num_bytes[1]), .A0(n1483), .A1(n1467), .Z(n1218));
Q_MX02 U1214 ( .S(pipe_ack_num_bytes[1]), .A0(n1484), .A1(n1468), .Z(n1219));
Q_MX02 U1215 ( .S(pipe_ack_num_bytes[1]), .A0(n1485), .A1(n1469), .Z(n1220));
Q_MX02 U1216 ( .S(pipe_ack_num_bytes[1]), .A0(n1486), .A1(n1470), .Z(n1221));
Q_MX02 U1217 ( .S(pipe_ack_num_bytes[1]), .A0(n1487), .A1(n1471), .Z(n1222));
Q_MX02 U1218 ( .S(pipe_ack_num_bytes[1]), .A0(n1488), .A1(n1472), .Z(n1223));
Q_MX02 U1219 ( .S(pipe_ack_num_bytes[1]), .A0(n1489), .A1(n1473), .Z(n1224));
Q_MX02 U1220 ( .S(pipe_ack_num_bytes[1]), .A0(n1490), .A1(n1474), .Z(n1225));
Q_MX02 U1221 ( .S(pipe_ack_num_bytes[1]), .A0(n1491), .A1(n1475), .Z(n1226));
Q_MX02 U1222 ( .S(pipe_ack_num_bytes[1]), .A0(n1492), .A1(n1476), .Z(n1227));
Q_MX02 U1223 ( .S(pipe_ack_num_bytes[1]), .A0(n1493), .A1(n1477), .Z(n1228));
Q_MX02 U1224 ( .S(pipe_ack_num_bytes[1]), .A0(n1494), .A1(n1478), .Z(n1229));
Q_MX02 U1225 ( .S(pipe_ack_num_bytes[1]), .A0(n1495), .A1(n1479), .Z(n1230));
Q_MX02 U1226 ( .S(pipe_ack_num_bytes[1]), .A0(n1496), .A1(n1480), .Z(n1231));
Q_MX02 U1227 ( .S(pipe_ack_num_bytes[1]), .A0(n1497), .A1(n1481), .Z(n1232));
Q_MX02 U1228 ( .S(pipe_ack_num_bytes[1]), .A0(n1498), .A1(n1482), .Z(n1233));
Q_MX02 U1229 ( .S(pipe_ack_num_bytes[1]), .A0(n1499), .A1(n1483), .Z(n1234));
Q_MX02 U1230 ( .S(pipe_ack_num_bytes[1]), .A0(n1500), .A1(n1484), .Z(n1235));
Q_MX02 U1231 ( .S(pipe_ack_num_bytes[1]), .A0(n1501), .A1(n1485), .Z(n1236));
Q_MX02 U1232 ( .S(pipe_ack_num_bytes[1]), .A0(n1502), .A1(n1486), .Z(n1237));
Q_MX02 U1233 ( .S(pipe_ack_num_bytes[1]), .A0(n1503), .A1(n1487), .Z(n1238));
Q_MX02 U1234 ( .S(pipe_ack_num_bytes[1]), .A0(n1504), .A1(n1488), .Z(n1239));
Q_MX02 U1235 ( .S(pipe_ack_num_bytes[1]), .A0(n1505), .A1(n1489), .Z(n1240));
Q_MX02 U1236 ( .S(pipe_ack_num_bytes[1]), .A0(n1506), .A1(n1490), .Z(n1241));
Q_MX02 U1237 ( .S(pipe_ack_num_bytes[1]), .A0(n1507), .A1(n1491), .Z(n1242));
Q_MX02 U1238 ( .S(pipe_ack_num_bytes[1]), .A0(n1508), .A1(n1492), .Z(n1243));
Q_MX02 U1239 ( .S(pipe_ack_num_bytes[1]), .A0(n1509), .A1(n1493), .Z(n1244));
Q_MX02 U1240 ( .S(pipe_ack_num_bytes[1]), .A0(n1510), .A1(n1494), .Z(n1245));
Q_MX02 U1241 ( .S(pipe_ack_num_bytes[1]), .A0(n1511), .A1(n1495), .Z(n1246));
Q_MX02 U1242 ( .S(pipe_ack_num_bytes[1]), .A0(n1512), .A1(n1496), .Z(n1247));
Q_MX02 U1243 ( .S(pipe_ack_num_bytes[1]), .A0(n1513), .A1(n1497), .Z(n1248));
Q_MX02 U1244 ( .S(pipe_ack_num_bytes[1]), .A0(n1514), .A1(n1498), .Z(n1249));
Q_MX02 U1245 ( .S(pipe_ack_num_bytes[1]), .A0(n1515), .A1(n1499), .Z(n1250));
Q_MX02 U1246 ( .S(pipe_ack_num_bytes[1]), .A0(n1516), .A1(n1500), .Z(n1251));
Q_MX02 U1247 ( .S(pipe_ack_num_bytes[1]), .A0(n1517), .A1(n1501), .Z(n1252));
Q_MX02 U1248 ( .S(pipe_ack_num_bytes[1]), .A0(n1518), .A1(n1502), .Z(n1253));
Q_MX02 U1249 ( .S(pipe_ack_num_bytes[1]), .A0(n1519), .A1(n1503), .Z(n1254));
Q_MX02 U1250 ( .S(pipe_ack_num_bytes[1]), .A0(n1520), .A1(n1504), .Z(n1255));
Q_MX02 U1251 ( .S(pipe_ack_num_bytes[1]), .A0(n1521), .A1(n1505), .Z(n1256));
Q_MX02 U1252 ( .S(pipe_ack_num_bytes[1]), .A0(n1522), .A1(n1506), .Z(n1257));
Q_MX02 U1253 ( .S(pipe_ack_num_bytes[1]), .A0(n1523), .A1(n1507), .Z(n1258));
Q_MX02 U1254 ( .S(pipe_ack_num_bytes[1]), .A0(n1524), .A1(n1508), .Z(n1259));
Q_MX02 U1255 ( .S(pipe_ack_num_bytes[1]), .A0(n1525), .A1(n1509), .Z(n1260));
Q_MX02 U1256 ( .S(pipe_ack_num_bytes[1]), .A0(n1526), .A1(n1510), .Z(n1261));
Q_MX02 U1257 ( .S(pipe_ack_num_bytes[1]), .A0(n1527), .A1(n1511), .Z(n1262));
Q_MX02 U1258 ( .S(pipe_ack_num_bytes[1]), .A0(n1528), .A1(n1512), .Z(n1263));
Q_MX02 U1259 ( .S(pipe_ack_num_bytes[1]), .A0(n1529), .A1(n1513), .Z(n1264));
Q_MX02 U1260 ( .S(pipe_ack_num_bytes[1]), .A0(n1530), .A1(n1514), .Z(n1265));
Q_MX02 U1261 ( .S(pipe_ack_num_bytes[1]), .A0(n1531), .A1(n1515), .Z(n1266));
Q_MX02 U1262 ( .S(pipe_ack_num_bytes[1]), .A0(n1532), .A1(n1516), .Z(n1267));
Q_MX02 U1263 ( .S(pipe_ack_num_bytes[1]), .A0(n1533), .A1(n1517), .Z(n1268));
Q_MX02 U1264 ( .S(pipe_ack_num_bytes[1]), .A0(n1534), .A1(n1518), .Z(n1269));
Q_MX02 U1265 ( .S(pipe_ack_num_bytes[1]), .A0(n1535), .A1(n1519), .Z(n1270));
Q_MX02 U1266 ( .S(pipe_ack_num_bytes[1]), .A0(n1536), .A1(n1520), .Z(n1271));
Q_MX02 U1267 ( .S(pipe_ack_num_bytes[1]), .A0(n1537), .A1(n1521), .Z(n1272));
Q_MX02 U1268 ( .S(pipe_ack_num_bytes[1]), .A0(n1538), .A1(n1522), .Z(n1273));
Q_MX02 U1269 ( .S(pipe_ack_num_bytes[1]), .A0(n1539), .A1(n1523), .Z(n1274));
Q_MX02 U1270 ( .S(pipe_ack_num_bytes[1]), .A0(n1540), .A1(n1524), .Z(n1275));
Q_MX02 U1271 ( .S(pipe_ack_num_bytes[1]), .A0(n1541), .A1(n1525), .Z(n1276));
Q_MX02 U1272 ( .S(pipe_ack_num_bytes[1]), .A0(n1542), .A1(n1526), .Z(n1277));
Q_MX02 U1273 ( .S(pipe_ack_num_bytes[1]), .A0(n1543), .A1(n1527), .Z(n1278));
Q_MX02 U1274 ( .S(pipe_ack_num_bytes[1]), .A0(n1544), .A1(n1528), .Z(n1279));
Q_MX02 U1275 ( .S(pipe_ack_num_bytes[1]), .A0(n1545), .A1(n1529), .Z(n1280));
Q_MX02 U1276 ( .S(pipe_ack_num_bytes[1]), .A0(n1546), .A1(n1530), .Z(n1281));
Q_MX02 U1277 ( .S(pipe_ack_num_bytes[1]), .A0(n1547), .A1(n1531), .Z(n1282));
Q_MX02 U1278 ( .S(pipe_ack_num_bytes[1]), .A0(n1548), .A1(n1532), .Z(n1283));
Q_MX02 U1279 ( .S(pipe_ack_num_bytes[1]), .A0(n1549), .A1(n1533), .Z(n1284));
Q_MX02 U1280 ( .S(pipe_ack_num_bytes[1]), .A0(n1550), .A1(n1534), .Z(n1285));
Q_MX02 U1281 ( .S(pipe_ack_num_bytes[1]), .A0(n1551), .A1(n1535), .Z(n1286));
Q_MX02 U1282 ( .S(pipe_ack_num_bytes[1]), .A0(n1552), .A1(n1536), .Z(n1287));
Q_MX02 U1283 ( .S(pipe_ack_num_bytes[1]), .A0(n1553), .A1(n1537), .Z(n1288));
Q_MX02 U1284 ( .S(pipe_ack_num_bytes[1]), .A0(n1554), .A1(n1538), .Z(n1289));
Q_MX02 U1285 ( .S(pipe_ack_num_bytes[1]), .A0(n1555), .A1(n1539), .Z(n1290));
Q_MX02 U1286 ( .S(pipe_ack_num_bytes[1]), .A0(n1556), .A1(n1540), .Z(n1291));
Q_MX02 U1287 ( .S(pipe_ack_num_bytes[1]), .A0(n1557), .A1(n1541), .Z(n1292));
Q_MX02 U1288 ( .S(pipe_ack_num_bytes[1]), .A0(n1558), .A1(n1542), .Z(n1293));
Q_MX02 U1289 ( .S(pipe_ack_num_bytes[1]), .A0(n1559), .A1(n1543), .Z(n1294));
Q_MX02 U1290 ( .S(pipe_ack_num_bytes[1]), .A0(n1560), .A1(n1544), .Z(n1295));
Q_MX02 U1291 ( .S(pipe_ack_num_bytes[1]), .A0(n1561), .A1(n1545), .Z(n1296));
Q_MX02 U1292 ( .S(pipe_ack_num_bytes[1]), .A0(n1562), .A1(n1546), .Z(n1297));
Q_MX02 U1293 ( .S(pipe_ack_num_bytes[1]), .A0(n1563), .A1(n1547), .Z(n1298));
Q_MX02 U1294 ( .S(pipe_ack_num_bytes[1]), .A0(n1564), .A1(n1548), .Z(n1299));
Q_MX02 U1295 ( .S(pipe_ack_num_bytes[1]), .A0(n1565), .A1(n1549), .Z(n1300));
Q_MX02 U1296 ( .S(pipe_ack_num_bytes[1]), .A0(n1566), .A1(n1550), .Z(n1301));
Q_MX02 U1297 ( .S(pipe_ack_num_bytes[1]), .A0(n1567), .A1(n1551), .Z(n1302));
Q_MX02 U1298 ( .S(pipe_ack_num_bytes[1]), .A0(n1568), .A1(n1552), .Z(n1303));
Q_MX02 U1299 ( .S(pipe_ack_num_bytes[1]), .A0(n1569), .A1(n1553), .Z(n1304));
Q_MX02 U1300 ( .S(pipe_ack_num_bytes[1]), .A0(n1570), .A1(n1554), .Z(n1305));
Q_MX02 U1301 ( .S(pipe_ack_num_bytes[1]), .A0(n1571), .A1(n1555), .Z(n1306));
Q_MX02 U1302 ( .S(pipe_ack_num_bytes[1]), .A0(n1572), .A1(n1556), .Z(n1307));
Q_MX02 U1303 ( .S(pipe_ack_num_bytes[1]), .A0(n1573), .A1(n1557), .Z(n1308));
Q_MX02 U1304 ( .S(pipe_ack_num_bytes[1]), .A0(n1574), .A1(n1558), .Z(n1309));
Q_MX02 U1305 ( .S(pipe_ack_num_bytes[1]), .A0(n1575), .A1(n1559), .Z(n1310));
Q_MX02 U1306 ( .S(pipe_ack_num_bytes[1]), .A0(n1576), .A1(n1560), .Z(n1311));
Q_MX02 U1307 ( .S(pipe_ack_num_bytes[1]), .A0(n1577), .A1(n1561), .Z(n1312));
Q_MX02 U1308 ( .S(pipe_ack_num_bytes[1]), .A0(n1578), .A1(n1562), .Z(n1313));
Q_MX02 U1309 ( .S(pipe_ack_num_bytes[1]), .A0(n1579), .A1(n1563), .Z(n1314));
Q_MX02 U1310 ( .S(pipe_ack_num_bytes[1]), .A0(n1580), .A1(n1564), .Z(n1315));
Q_MX02 U1311 ( .S(pipe_ack_num_bytes[1]), .A0(n1581), .A1(n1565), .Z(n1316));
Q_MX02 U1312 ( .S(pipe_ack_num_bytes[1]), .A0(n1582), .A1(n1566), .Z(n1317));
Q_MX02 U1313 ( .S(pipe_ack_num_bytes[1]), .A0(n1583), .A1(n1567), .Z(n1318));
Q_MX02 U1314 ( .S(pipe_ack_num_bytes[1]), .A0(n1584), .A1(n1568), .Z(n1319));
Q_MX02 U1315 ( .S(pipe_ack_num_bytes[1]), .A0(n1585), .A1(n1569), .Z(n1320));
Q_MX02 U1316 ( .S(pipe_ack_num_bytes[1]), .A0(n1586), .A1(n1570), .Z(n1321));
Q_MX02 U1317 ( .S(pipe_ack_num_bytes[1]), .A0(n1587), .A1(n1571), .Z(n1322));
Q_MX02 U1318 ( .S(pipe_ack_num_bytes[1]), .A0(n1588), .A1(n1572), .Z(n1323));
Q_MX02 U1319 ( .S(pipe_ack_num_bytes[1]), .A0(n1589), .A1(n1573), .Z(n1324));
Q_MX02 U1320 ( .S(pipe_ack_num_bytes[1]), .A0(n1590), .A1(n1574), .Z(n1325));
Q_MX02 U1321 ( .S(pipe_ack_num_bytes[1]), .A0(n1591), .A1(n1575), .Z(n1326));
Q_MX02 U1322 ( .S(pipe_ack_num_bytes[1]), .A0(n1592), .A1(n1576), .Z(n1327));
Q_MX02 U1323 ( .S(pipe_ack_num_bytes[1]), .A0(n1593), .A1(n1577), .Z(n1328));
Q_MX02 U1324 ( .S(pipe_ack_num_bytes[1]), .A0(n1594), .A1(n1578), .Z(n1329));
Q_MX02 U1325 ( .S(pipe_ack_num_bytes[1]), .A0(n1595), .A1(n1579), .Z(n1330));
Q_MX02 U1326 ( .S(pipe_ack_num_bytes[1]), .A0(n1596), .A1(n1580), .Z(n1331));
Q_MX02 U1327 ( .S(pipe_ack_num_bytes[1]), .A0(n1597), .A1(n1581), .Z(n1332));
Q_MX02 U1328 ( .S(pipe_ack_num_bytes[1]), .A0(n1598), .A1(n1582), .Z(n1333));
Q_MX02 U1329 ( .S(pipe_ack_num_bytes[1]), .A0(n1599), .A1(n1583), .Z(n1334));
Q_MX02 U1330 ( .S(pipe_ack_num_bytes[1]), .A0(n1600), .A1(n1584), .Z(n1335));
Q_MX02 U1331 ( .S(pipe_ack_num_bytes[1]), .A0(n1601), .A1(n1585), .Z(n1336));
Q_MX02 U1332 ( .S(pipe_ack_num_bytes[1]), .A0(n1602), .A1(n1586), .Z(n1337));
Q_MX02 U1333 ( .S(pipe_ack_num_bytes[1]), .A0(n1603), .A1(n1587), .Z(n1338));
Q_MX02 U1334 ( .S(pipe_ack_num_bytes[1]), .A0(n1604), .A1(n1588), .Z(n1339));
Q_MX02 U1335 ( .S(pipe_ack_num_bytes[1]), .A0(n1605), .A1(n1589), .Z(n1340));
Q_MX02 U1336 ( .S(pipe_ack_num_bytes[1]), .A0(n1606), .A1(n1590), .Z(n1341));
Q_MX02 U1337 ( .S(pipe_ack_num_bytes[1]), .A0(n1607), .A1(n1591), .Z(n1342));
Q_AN02 U1338 ( .A0(n1351), .A1(cmd_data_q[0]), .Z(n1343));
Q_AN02 U1339 ( .A0(n1351), .A1(cmd_data_q[1]), .Z(n1344));
Q_AN02 U1340 ( .A0(n1351), .A1(cmd_data_q[2]), .Z(n1345));
Q_AN02 U1341 ( .A0(n1351), .A1(cmd_data_q[3]), .Z(n1346));
Q_AN02 U1342 ( .A0(n1351), .A1(cmd_data_q[4]), .Z(n1347));
Q_AN02 U1343 ( .A0(n1351), .A1(cmd_data_q[5]), .Z(n1348));
Q_AN02 U1344 ( .A0(n1351), .A1(cmd_data_q[6]), .Z(n1349));
Q_AN02 U1345 ( .A0(n1351), .A1(cmd_data_q[7]), .Z(n1350));
Q_INV U1346 ( .A(pipe_ack_num_bytes[0]), .Z(n1351));
Q_MX02 U1347 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[8]), .A1(cmd_data_q[0]), .Z(n1352));
Q_MX02 U1348 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[9]), .A1(cmd_data_q[1]), .Z(n1353));
Q_MX02 U1349 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[10]), .A1(cmd_data_q[2]), .Z(n1354));
Q_MX02 U1350 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[11]), .A1(cmd_data_q[3]), .Z(n1355));
Q_MX02 U1351 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[12]), .A1(cmd_data_q[4]), .Z(n1356));
Q_MX02 U1352 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[13]), .A1(cmd_data_q[5]), .Z(n1357));
Q_MX02 U1353 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[14]), .A1(cmd_data_q[6]), .Z(n1358));
Q_MX02 U1354 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[15]), .A1(cmd_data_q[7]), .Z(n1359));
Q_MX02 U1355 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[16]), .A1(cmd_data_q[8]), .Z(n1360));
Q_MX02 U1356 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[17]), .A1(cmd_data_q[9]), .Z(n1361));
Q_MX02 U1357 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[18]), .A1(cmd_data_q[10]), .Z(n1362));
Q_MX02 U1358 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[19]), .A1(cmd_data_q[11]), .Z(n1363));
Q_MX02 U1359 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[20]), .A1(cmd_data_q[12]), .Z(n1364));
Q_MX02 U1360 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[21]), .A1(cmd_data_q[13]), .Z(n1365));
Q_MX02 U1361 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[22]), .A1(cmd_data_q[14]), .Z(n1366));
Q_MX02 U1362 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[23]), .A1(cmd_data_q[15]), .Z(n1367));
Q_MX02 U1363 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[24]), .A1(cmd_data_q[16]), .Z(n1368));
Q_MX02 U1364 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[25]), .A1(cmd_data_q[17]), .Z(n1369));
Q_MX02 U1365 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[26]), .A1(cmd_data_q[18]), .Z(n1370));
Q_MX02 U1366 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[27]), .A1(cmd_data_q[19]), .Z(n1371));
Q_MX02 U1367 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[28]), .A1(cmd_data_q[20]), .Z(n1372));
Q_MX02 U1368 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[29]), .A1(cmd_data_q[21]), .Z(n1373));
Q_MX02 U1369 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[30]), .A1(cmd_data_q[22]), .Z(n1374));
Q_MX02 U1370 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[31]), .A1(cmd_data_q[23]), .Z(n1375));
Q_MX02 U1371 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[32]), .A1(cmd_data_q[24]), .Z(n1376));
Q_MX02 U1372 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[33]), .A1(cmd_data_q[25]), .Z(n1377));
Q_MX02 U1373 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[34]), .A1(cmd_data_q[26]), .Z(n1378));
Q_MX02 U1374 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[35]), .A1(cmd_data_q[27]), .Z(n1379));
Q_MX02 U1375 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[36]), .A1(cmd_data_q[28]), .Z(n1380));
Q_MX02 U1376 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[37]), .A1(cmd_data_q[29]), .Z(n1381));
Q_MX02 U1377 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[38]), .A1(cmd_data_q[30]), .Z(n1382));
Q_MX02 U1378 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[39]), .A1(cmd_data_q[31]), .Z(n1383));
Q_MX02 U1379 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[40]), .A1(cmd_data_q[32]), .Z(n1384));
Q_MX02 U1380 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[41]), .A1(cmd_data_q[33]), .Z(n1385));
Q_MX02 U1381 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[42]), .A1(cmd_data_q[34]), .Z(n1386));
Q_MX02 U1382 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[43]), .A1(cmd_data_q[35]), .Z(n1387));
Q_MX02 U1383 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[44]), .A1(cmd_data_q[36]), .Z(n1388));
Q_MX02 U1384 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[45]), .A1(cmd_data_q[37]), .Z(n1389));
Q_MX02 U1385 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[46]), .A1(cmd_data_q[38]), .Z(n1390));
Q_MX02 U1386 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[47]), .A1(cmd_data_q[39]), .Z(n1391));
Q_MX02 U1387 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[48]), .A1(cmd_data_q[40]), .Z(n1392));
Q_MX02 U1388 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[49]), .A1(cmd_data_q[41]), .Z(n1393));
Q_MX02 U1389 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[50]), .A1(cmd_data_q[42]), .Z(n1394));
Q_MX02 U1390 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[51]), .A1(cmd_data_q[43]), .Z(n1395));
Q_MX02 U1391 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[52]), .A1(cmd_data_q[44]), .Z(n1396));
Q_MX02 U1392 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[53]), .A1(cmd_data_q[45]), .Z(n1397));
Q_MX02 U1393 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[54]), .A1(cmd_data_q[46]), .Z(n1398));
Q_MX02 U1394 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[55]), .A1(cmd_data_q[47]), .Z(n1399));
Q_MX02 U1395 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[56]), .A1(cmd_data_q[48]), .Z(n1400));
Q_MX02 U1396 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[57]), .A1(cmd_data_q[49]), .Z(n1401));
Q_MX02 U1397 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[58]), .A1(cmd_data_q[50]), .Z(n1402));
Q_MX02 U1398 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[59]), .A1(cmd_data_q[51]), .Z(n1403));
Q_MX02 U1399 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[60]), .A1(cmd_data_q[52]), .Z(n1404));
Q_MX02 U1400 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[61]), .A1(cmd_data_q[53]), .Z(n1405));
Q_MX02 U1401 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[62]), .A1(cmd_data_q[54]), .Z(n1406));
Q_MX02 U1402 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[63]), .A1(cmd_data_q[55]), .Z(n1407));
Q_MX02 U1403 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[64]), .A1(cmd_data_q[56]), .Z(n1408));
Q_MX02 U1404 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[65]), .A1(cmd_data_q[57]), .Z(n1409));
Q_MX02 U1405 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[66]), .A1(cmd_data_q[58]), .Z(n1410));
Q_MX02 U1406 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[67]), .A1(cmd_data_q[59]), .Z(n1411));
Q_MX02 U1407 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[68]), .A1(cmd_data_q[60]), .Z(n1412));
Q_MX02 U1408 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[69]), .A1(cmd_data_q[61]), .Z(n1413));
Q_MX02 U1409 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[70]), .A1(cmd_data_q[62]), .Z(n1414));
Q_MX02 U1410 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[71]), .A1(cmd_data_q[63]), .Z(n1415));
Q_MX02 U1411 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[72]), .A1(cmd_data_q[64]), .Z(n1416));
Q_MX02 U1412 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[73]), .A1(cmd_data_q[65]), .Z(n1417));
Q_MX02 U1413 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[74]), .A1(cmd_data_q[66]), .Z(n1418));
Q_MX02 U1414 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[75]), .A1(cmd_data_q[67]), .Z(n1419));
Q_MX02 U1415 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[76]), .A1(cmd_data_q[68]), .Z(n1420));
Q_MX02 U1416 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[77]), .A1(cmd_data_q[69]), .Z(n1421));
Q_MX02 U1417 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[78]), .A1(cmd_data_q[70]), .Z(n1422));
Q_MX02 U1418 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[79]), .A1(cmd_data_q[71]), .Z(n1423));
Q_MX02 U1419 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[80]), .A1(cmd_data_q[72]), .Z(n1424));
Q_MX02 U1420 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[81]), .A1(cmd_data_q[73]), .Z(n1425));
Q_MX02 U1421 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[82]), .A1(cmd_data_q[74]), .Z(n1426));
Q_MX02 U1422 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[83]), .A1(cmd_data_q[75]), .Z(n1427));
Q_MX02 U1423 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[84]), .A1(cmd_data_q[76]), .Z(n1428));
Q_MX02 U1424 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[85]), .A1(cmd_data_q[77]), .Z(n1429));
Q_MX02 U1425 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[86]), .A1(cmd_data_q[78]), .Z(n1430));
Q_MX02 U1426 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[87]), .A1(cmd_data_q[79]), .Z(n1431));
Q_MX02 U1427 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[88]), .A1(cmd_data_q[80]), .Z(n1432));
Q_MX02 U1428 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[89]), .A1(cmd_data_q[81]), .Z(n1433));
Q_MX02 U1429 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[90]), .A1(cmd_data_q[82]), .Z(n1434));
Q_MX02 U1430 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[91]), .A1(cmd_data_q[83]), .Z(n1435));
Q_MX02 U1431 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[92]), .A1(cmd_data_q[84]), .Z(n1436));
Q_MX02 U1432 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[93]), .A1(cmd_data_q[85]), .Z(n1437));
Q_MX02 U1433 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[94]), .A1(cmd_data_q[86]), .Z(n1438));
Q_MX02 U1434 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[95]), .A1(cmd_data_q[87]), .Z(n1439));
Q_MX02 U1435 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[96]), .A1(cmd_data_q[88]), .Z(n1440));
Q_MX02 U1436 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[97]), .A1(cmd_data_q[89]), .Z(n1441));
Q_MX02 U1437 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[98]), .A1(cmd_data_q[90]), .Z(n1442));
Q_MX02 U1438 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[99]), .A1(cmd_data_q[91]), .Z(n1443));
Q_MX02 U1439 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[100]), .A1(cmd_data_q[92]), .Z(n1444));
Q_MX02 U1440 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[101]), .A1(cmd_data_q[93]), .Z(n1445));
Q_MX02 U1441 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[102]), .A1(cmd_data_q[94]), .Z(n1446));
Q_MX02 U1442 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[103]), .A1(cmd_data_q[95]), .Z(n1447));
Q_MX02 U1443 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[104]), .A1(cmd_data_q[96]), .Z(n1448));
Q_MX02 U1444 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[105]), .A1(cmd_data_q[97]), .Z(n1449));
Q_MX02 U1445 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[106]), .A1(cmd_data_q[98]), .Z(n1450));
Q_MX02 U1446 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[107]), .A1(cmd_data_q[99]), .Z(n1451));
Q_MX02 U1447 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[108]), .A1(cmd_data_q[100]), .Z(n1452));
Q_MX02 U1448 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[109]), .A1(cmd_data_q[101]), .Z(n1453));
Q_MX02 U1449 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[110]), .A1(cmd_data_q[102]), .Z(n1454));
Q_MX02 U1450 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[111]), .A1(cmd_data_q[103]), .Z(n1455));
Q_MX02 U1451 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[112]), .A1(cmd_data_q[104]), .Z(n1456));
Q_MX02 U1452 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[113]), .A1(cmd_data_q[105]), .Z(n1457));
Q_MX02 U1453 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[114]), .A1(cmd_data_q[106]), .Z(n1458));
Q_MX02 U1454 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[115]), .A1(cmd_data_q[107]), .Z(n1459));
Q_MX02 U1455 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[116]), .A1(cmd_data_q[108]), .Z(n1460));
Q_MX02 U1456 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[117]), .A1(cmd_data_q[109]), .Z(n1461));
Q_MX02 U1457 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[118]), .A1(cmd_data_q[110]), .Z(n1462));
Q_MX02 U1458 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[119]), .A1(cmd_data_q[111]), .Z(n1463));
Q_MX02 U1459 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[120]), .A1(cmd_data_q[112]), .Z(n1464));
Q_MX02 U1460 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[121]), .A1(cmd_data_q[113]), .Z(n1465));
Q_MX02 U1461 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[122]), .A1(cmd_data_q[114]), .Z(n1466));
Q_MX02 U1462 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[123]), .A1(cmd_data_q[115]), .Z(n1467));
Q_MX02 U1463 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[124]), .A1(cmd_data_q[116]), .Z(n1468));
Q_MX02 U1464 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[125]), .A1(cmd_data_q[117]), .Z(n1469));
Q_MX02 U1465 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[126]), .A1(cmd_data_q[118]), .Z(n1470));
Q_MX02 U1466 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[127]), .A1(cmd_data_q[119]), .Z(n1471));
Q_MX02 U1467 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[128]), .A1(cmd_data_q[120]), .Z(n1472));
Q_MX02 U1468 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[129]), .A1(cmd_data_q[121]), .Z(n1473));
Q_MX02 U1469 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[130]), .A1(cmd_data_q[122]), .Z(n1474));
Q_MX02 U1470 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[131]), .A1(cmd_data_q[123]), .Z(n1475));
Q_MX02 U1471 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[132]), .A1(cmd_data_q[124]), .Z(n1476));
Q_MX02 U1472 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[133]), .A1(cmd_data_q[125]), .Z(n1477));
Q_MX02 U1473 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[134]), .A1(cmd_data_q[126]), .Z(n1478));
Q_MX02 U1474 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[135]), .A1(cmd_data_q[127]), .Z(n1479));
Q_MX02 U1475 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[136]), .A1(cmd_data_q[128]), .Z(n1480));
Q_MX02 U1476 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[137]), .A1(cmd_data_q[129]), .Z(n1481));
Q_MX02 U1477 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[138]), .A1(cmd_data_q[130]), .Z(n1482));
Q_MX02 U1478 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[139]), .A1(cmd_data_q[131]), .Z(n1483));
Q_MX02 U1479 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[140]), .A1(cmd_data_q[132]), .Z(n1484));
Q_MX02 U1480 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[141]), .A1(cmd_data_q[133]), .Z(n1485));
Q_MX02 U1481 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[142]), .A1(cmd_data_q[134]), .Z(n1486));
Q_MX02 U1482 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[143]), .A1(cmd_data_q[135]), .Z(n1487));
Q_MX02 U1483 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[144]), .A1(cmd_data_q[136]), .Z(n1488));
Q_MX02 U1484 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[145]), .A1(cmd_data_q[137]), .Z(n1489));
Q_MX02 U1485 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[146]), .A1(cmd_data_q[138]), .Z(n1490));
Q_MX02 U1486 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[147]), .A1(cmd_data_q[139]), .Z(n1491));
Q_MX02 U1487 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[148]), .A1(cmd_data_q[140]), .Z(n1492));
Q_MX02 U1488 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[149]), .A1(cmd_data_q[141]), .Z(n1493));
Q_MX02 U1489 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[150]), .A1(cmd_data_q[142]), .Z(n1494));
Q_MX02 U1490 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[151]), .A1(cmd_data_q[143]), .Z(n1495));
Q_MX02 U1491 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[152]), .A1(cmd_data_q[144]), .Z(n1496));
Q_MX02 U1492 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[153]), .A1(cmd_data_q[145]), .Z(n1497));
Q_MX02 U1493 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[154]), .A1(cmd_data_q[146]), .Z(n1498));
Q_MX02 U1494 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[155]), .A1(cmd_data_q[147]), .Z(n1499));
Q_MX02 U1495 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[156]), .A1(cmd_data_q[148]), .Z(n1500));
Q_MX02 U1496 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[157]), .A1(cmd_data_q[149]), .Z(n1501));
Q_MX02 U1497 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[158]), .A1(cmd_data_q[150]), .Z(n1502));
Q_MX02 U1498 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[159]), .A1(cmd_data_q[151]), .Z(n1503));
Q_MX02 U1499 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[160]), .A1(cmd_data_q[152]), .Z(n1504));
Q_MX02 U1500 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[161]), .A1(cmd_data_q[153]), .Z(n1505));
Q_MX02 U1501 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[162]), .A1(cmd_data_q[154]), .Z(n1506));
Q_MX02 U1502 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[163]), .A1(cmd_data_q[155]), .Z(n1507));
Q_MX02 U1503 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[164]), .A1(cmd_data_q[156]), .Z(n1508));
Q_MX02 U1504 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[165]), .A1(cmd_data_q[157]), .Z(n1509));
Q_MX02 U1505 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[166]), .A1(cmd_data_q[158]), .Z(n1510));
Q_MX02 U1506 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[167]), .A1(cmd_data_q[159]), .Z(n1511));
Q_MX02 U1507 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[168]), .A1(cmd_data_q[160]), .Z(n1512));
Q_MX02 U1508 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[169]), .A1(cmd_data_q[161]), .Z(n1513));
Q_MX02 U1509 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[170]), .A1(cmd_data_q[162]), .Z(n1514));
Q_MX02 U1510 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[171]), .A1(cmd_data_q[163]), .Z(n1515));
Q_MX02 U1511 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[172]), .A1(cmd_data_q[164]), .Z(n1516));
Q_MX02 U1512 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[173]), .A1(cmd_data_q[165]), .Z(n1517));
Q_MX02 U1513 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[174]), .A1(cmd_data_q[166]), .Z(n1518));
Q_MX02 U1514 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[175]), .A1(cmd_data_q[167]), .Z(n1519));
Q_MX02 U1515 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[176]), .A1(cmd_data_q[168]), .Z(n1520));
Q_MX02 U1516 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[177]), .A1(cmd_data_q[169]), .Z(n1521));
Q_MX02 U1517 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[178]), .A1(cmd_data_q[170]), .Z(n1522));
Q_MX02 U1518 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[179]), .A1(cmd_data_q[171]), .Z(n1523));
Q_MX02 U1519 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[180]), .A1(cmd_data_q[172]), .Z(n1524));
Q_MX02 U1520 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[181]), .A1(cmd_data_q[173]), .Z(n1525));
Q_MX02 U1521 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[182]), .A1(cmd_data_q[174]), .Z(n1526));
Q_MX02 U1522 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[183]), .A1(cmd_data_q[175]), .Z(n1527));
Q_MX02 U1523 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[184]), .A1(cmd_data_q[176]), .Z(n1528));
Q_MX02 U1524 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[185]), .A1(cmd_data_q[177]), .Z(n1529));
Q_MX02 U1525 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[186]), .A1(cmd_data_q[178]), .Z(n1530));
Q_MX02 U1526 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[187]), .A1(cmd_data_q[179]), .Z(n1531));
Q_MX02 U1527 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[188]), .A1(cmd_data_q[180]), .Z(n1532));
Q_MX02 U1528 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[189]), .A1(cmd_data_q[181]), .Z(n1533));
Q_MX02 U1529 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[190]), .A1(cmd_data_q[182]), .Z(n1534));
Q_MX02 U1530 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[191]), .A1(cmd_data_q[183]), .Z(n1535));
Q_MX02 U1531 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[192]), .A1(cmd_data_q[184]), .Z(n1536));
Q_MX02 U1532 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[193]), .A1(cmd_data_q[185]), .Z(n1537));
Q_MX02 U1533 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[194]), .A1(cmd_data_q[186]), .Z(n1538));
Q_MX02 U1534 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[195]), .A1(cmd_data_q[187]), .Z(n1539));
Q_MX02 U1535 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[196]), .A1(cmd_data_q[188]), .Z(n1540));
Q_MX02 U1536 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[197]), .A1(cmd_data_q[189]), .Z(n1541));
Q_MX02 U1537 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[198]), .A1(cmd_data_q[190]), .Z(n1542));
Q_MX02 U1538 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[199]), .A1(cmd_data_q[191]), .Z(n1543));
Q_MX02 U1539 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[200]), .A1(cmd_data_q[192]), .Z(n1544));
Q_MX02 U1540 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[201]), .A1(cmd_data_q[193]), .Z(n1545));
Q_MX02 U1541 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[202]), .A1(cmd_data_q[194]), .Z(n1546));
Q_MX02 U1542 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[203]), .A1(cmd_data_q[195]), .Z(n1547));
Q_MX02 U1543 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[204]), .A1(cmd_data_q[196]), .Z(n1548));
Q_MX02 U1544 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[205]), .A1(cmd_data_q[197]), .Z(n1549));
Q_MX02 U1545 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[206]), .A1(cmd_data_q[198]), .Z(n1550));
Q_MX02 U1546 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[207]), .A1(cmd_data_q[199]), .Z(n1551));
Q_MX02 U1547 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[208]), .A1(cmd_data_q[200]), .Z(n1552));
Q_MX02 U1548 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[209]), .A1(cmd_data_q[201]), .Z(n1553));
Q_MX02 U1549 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[210]), .A1(cmd_data_q[202]), .Z(n1554));
Q_MX02 U1550 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[211]), .A1(cmd_data_q[203]), .Z(n1555));
Q_MX02 U1551 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[212]), .A1(cmd_data_q[204]), .Z(n1556));
Q_MX02 U1552 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[213]), .A1(cmd_data_q[205]), .Z(n1557));
Q_MX02 U1553 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[214]), .A1(cmd_data_q[206]), .Z(n1558));
Q_MX02 U1554 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[215]), .A1(cmd_data_q[207]), .Z(n1559));
Q_MX02 U1555 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[216]), .A1(cmd_data_q[208]), .Z(n1560));
Q_MX02 U1556 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[217]), .A1(cmd_data_q[209]), .Z(n1561));
Q_MX02 U1557 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[218]), .A1(cmd_data_q[210]), .Z(n1562));
Q_MX02 U1558 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[219]), .A1(cmd_data_q[211]), .Z(n1563));
Q_MX02 U1559 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[220]), .A1(cmd_data_q[212]), .Z(n1564));
Q_MX02 U1560 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[221]), .A1(cmd_data_q[213]), .Z(n1565));
Q_MX02 U1561 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[222]), .A1(cmd_data_q[214]), .Z(n1566));
Q_MX02 U1562 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[223]), .A1(cmd_data_q[215]), .Z(n1567));
Q_MX02 U1563 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[224]), .A1(cmd_data_q[216]), .Z(n1568));
Q_MX02 U1564 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[225]), .A1(cmd_data_q[217]), .Z(n1569));
Q_MX02 U1565 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[226]), .A1(cmd_data_q[218]), .Z(n1570));
Q_MX02 U1566 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[227]), .A1(cmd_data_q[219]), .Z(n1571));
Q_MX02 U1567 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[228]), .A1(cmd_data_q[220]), .Z(n1572));
Q_MX02 U1568 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[229]), .A1(cmd_data_q[221]), .Z(n1573));
Q_MX02 U1569 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[230]), .A1(cmd_data_q[222]), .Z(n1574));
Q_MX02 U1570 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[231]), .A1(cmd_data_q[223]), .Z(n1575));
Q_MX02 U1571 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[232]), .A1(cmd_data_q[224]), .Z(n1576));
Q_MX02 U1572 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[233]), .A1(cmd_data_q[225]), .Z(n1577));
Q_MX02 U1573 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[234]), .A1(cmd_data_q[226]), .Z(n1578));
Q_MX02 U1574 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[235]), .A1(cmd_data_q[227]), .Z(n1579));
Q_MX02 U1575 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[236]), .A1(cmd_data_q[228]), .Z(n1580));
Q_MX02 U1576 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[237]), .A1(cmd_data_q[229]), .Z(n1581));
Q_MX02 U1577 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[238]), .A1(cmd_data_q[230]), .Z(n1582));
Q_MX02 U1578 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[239]), .A1(cmd_data_q[231]), .Z(n1583));
Q_MX02 U1579 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[240]), .A1(cmd_data_q[232]), .Z(n1584));
Q_MX02 U1580 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[241]), .A1(cmd_data_q[233]), .Z(n1585));
Q_MX02 U1581 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[242]), .A1(cmd_data_q[234]), .Z(n1586));
Q_MX02 U1582 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[243]), .A1(cmd_data_q[235]), .Z(n1587));
Q_MX02 U1583 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[244]), .A1(cmd_data_q[236]), .Z(n1588));
Q_MX02 U1584 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[245]), .A1(cmd_data_q[237]), .Z(n1589));
Q_MX02 U1585 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[246]), .A1(cmd_data_q[238]), .Z(n1590));
Q_MX02 U1586 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[247]), .A1(cmd_data_q[239]), .Z(n1591));
Q_MX02 U1587 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[248]), .A1(cmd_data_q[240]), .Z(n1592));
Q_MX02 U1588 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[249]), .A1(cmd_data_q[241]), .Z(n1593));
Q_MX02 U1589 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[250]), .A1(cmd_data_q[242]), .Z(n1594));
Q_MX02 U1590 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[251]), .A1(cmd_data_q[243]), .Z(n1595));
Q_MX02 U1591 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[252]), .A1(cmd_data_q[244]), .Z(n1596));
Q_MX02 U1592 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[253]), .A1(cmd_data_q[245]), .Z(n1597));
Q_MX02 U1593 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[254]), .A1(cmd_data_q[246]), .Z(n1598));
Q_MX02 U1594 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[255]), .A1(cmd_data_q[247]), .Z(n1599));
Q_MX02 U1595 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[256]), .A1(cmd_data_q[248]), .Z(n1600));
Q_MX02 U1596 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[257]), .A1(cmd_data_q[249]), .Z(n1601));
Q_MX02 U1597 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[258]), .A1(cmd_data_q[250]), .Z(n1602));
Q_MX02 U1598 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[259]), .A1(cmd_data_q[251]), .Z(n1603));
Q_MX02 U1599 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[260]), .A1(cmd_data_q[252]), .Z(n1604));
Q_MX02 U1600 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[261]), .A1(cmd_data_q[253]), .Z(n1605));
Q_MX02 U1601 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[262]), .A1(cmd_data_q[254]), .Z(n1606));
Q_MX02 U1602 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[263]), .A1(cmd_data_q[255]), .Z(n1607));
Q_MX02 U1603 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[264]), .A1(cmd_data_q[256]), .Z(n1608));
Q_MX02 U1604 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[265]), .A1(cmd_data_q[257]), .Z(n1609));
Q_MX02 U1605 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[266]), .A1(cmd_data_q[258]), .Z(n1610));
Q_MX02 U1606 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[267]), .A1(cmd_data_q[259]), .Z(n1611));
Q_MX02 U1607 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[268]), .A1(cmd_data_q[260]), .Z(n1612));
Q_MX02 U1608 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[269]), .A1(cmd_data_q[261]), .Z(n1613));
Q_MX02 U1609 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[270]), .A1(cmd_data_q[262]), .Z(n1614));
Q_MX02 U1610 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[271]), .A1(cmd_data_q[263]), .Z(n1615));
Q_MX02 U1611 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[272]), .A1(cmd_data_q[264]), .Z(n1616));
Q_MX02 U1612 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[273]), .A1(cmd_data_q[265]), .Z(n1617));
Q_MX02 U1613 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[274]), .A1(cmd_data_q[266]), .Z(n1618));
Q_MX02 U1614 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[275]), .A1(cmd_data_q[267]), .Z(n1619));
Q_MX02 U1615 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[276]), .A1(cmd_data_q[268]), .Z(n1620));
Q_MX02 U1616 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[277]), .A1(cmd_data_q[269]), .Z(n1621));
Q_MX02 U1617 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[278]), .A1(cmd_data_q[270]), .Z(n1622));
Q_MX02 U1618 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[279]), .A1(cmd_data_q[271]), .Z(n1623));
Q_MX02 U1619 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[280]), .A1(cmd_data_q[272]), .Z(n1624));
Q_MX02 U1620 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[281]), .A1(cmd_data_q[273]), .Z(n1625));
Q_MX02 U1621 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[282]), .A1(cmd_data_q[274]), .Z(n1626));
Q_MX02 U1622 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[283]), .A1(cmd_data_q[275]), .Z(n1627));
Q_MX02 U1623 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[284]), .A1(cmd_data_q[276]), .Z(n1628));
Q_MX02 U1624 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[285]), .A1(cmd_data_q[277]), .Z(n1629));
Q_MX02 U1625 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[286]), .A1(cmd_data_q[278]), .Z(n1630));
Q_MX02 U1626 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[287]), .A1(cmd_data_q[279]), .Z(n1631));
Q_MX02 U1627 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[288]), .A1(cmd_data_q[280]), .Z(n1632));
Q_MX02 U1628 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[289]), .A1(cmd_data_q[281]), .Z(n1633));
Q_MX02 U1629 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[290]), .A1(cmd_data_q[282]), .Z(n1634));
Q_MX02 U1630 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[291]), .A1(cmd_data_q[283]), .Z(n1635));
Q_MX02 U1631 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[292]), .A1(cmd_data_q[284]), .Z(n1636));
Q_MX02 U1632 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[293]), .A1(cmd_data_q[285]), .Z(n1637));
Q_MX02 U1633 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[294]), .A1(cmd_data_q[286]), .Z(n1638));
Q_MX02 U1634 ( .S(pipe_ack_num_bytes[0]), .A0(cmd_data_q[295]), .A1(cmd_data_q[287]), .Z(n1639));
ixc_assign_128 _zz_strnp_0 ( pipe_data[127:0], cmd_data_q[295:168]);
Q_OR03 U1636 ( .A0(pipe_byte_count[5]), .A1(pipe_byte_count[4]), .A2(pipe_byte_count[3]), .Z(n1641));
Q_OR03 U1637 ( .A0(pipe_byte_count[2]), .A1(pipe_byte_count[1]), .A2(pipe_byte_count[0]), .Z(n1640));
Q_OR02 U1638 ( .A0(n1641), .A1(n1640), .Z(pipe_valid[0]));
ixc_assign_6 _zz_strnp_1 ( _zy_simnet_pipe_byte_count_0_w$[0:5], 
	pipe_byte_count[5:0]);
Q_INV U1640 ( .A(n3), .Z(n1642));
Q_FDP4EP \pipe_byte_count_REG[5] ( .CK(clk), .CE(n1642), .R(n1643), .D(n4), .Q(pipe_byte_count[5]));
Q_INV U1642 ( .A(rst_n), .Z(n1643));
Q_FDP4EP \pipe_byte_count_REG[4] ( .CK(clk), .CE(n1642), .R(n1643), .D(n5), .Q(pipe_byte_count[4]));
Q_FDP4EP \pipe_byte_count_REG[3] ( .CK(clk), .CE(n1642), .R(n1643), .D(n6), .Q(pipe_byte_count[3]));
Q_FDP4EP \pipe_byte_count_REG[2] ( .CK(clk), .CE(n1642), .R(n1643), .D(n7), .Q(pipe_byte_count[2]));
Q_FDP4EP \pipe_byte_count_REG[1] ( .CK(clk), .CE(n1642), .R(n1643), .D(n8), .Q(pipe_byte_count[1]));
Q_FDP4EP \pipe_byte_count_REG[0] ( .CK(clk), .CE(n1642), .R(n1643), .D(n9), .Q(pipe_byte_count[0]));
Q_FDP4EP \cmd_data_q_REG[295] ( .CK(clk), .CE(n1642), .R(n1643), .D(n10), .Q(cmd_data_q[295]));
Q_FDP4EP \cmd_data_q_REG[294] ( .CK(clk), .CE(n1642), .R(n1643), .D(n11), .Q(cmd_data_q[294]));
Q_FDP4EP \cmd_data_q_REG[293] ( .CK(clk), .CE(n1642), .R(n1643), .D(n12), .Q(cmd_data_q[293]));
Q_FDP4EP \cmd_data_q_REG[292] ( .CK(clk), .CE(n1642), .R(n1643), .D(n13), .Q(cmd_data_q[292]));
Q_FDP4EP \cmd_data_q_REG[291] ( .CK(clk), .CE(n1642), .R(n1643), .D(n14), .Q(cmd_data_q[291]));
Q_FDP4EP \cmd_data_q_REG[290] ( .CK(clk), .CE(n1642), .R(n1643), .D(n15), .Q(cmd_data_q[290]));
Q_FDP4EP \cmd_data_q_REG[289] ( .CK(clk), .CE(n1642), .R(n1643), .D(n16), .Q(cmd_data_q[289]));
Q_FDP4EP \cmd_data_q_REG[288] ( .CK(clk), .CE(n1642), .R(n1643), .D(n17), .Q(cmd_data_q[288]));
Q_FDP4EP \cmd_data_q_REG[287] ( .CK(clk), .CE(n1642), .R(n1643), .D(n18), .Q(cmd_data_q[287]));
Q_FDP4EP \cmd_data_q_REG[286] ( .CK(clk), .CE(n1642), .R(n1643), .D(n19), .Q(cmd_data_q[286]));
Q_FDP4EP \cmd_data_q_REG[285] ( .CK(clk), .CE(n1642), .R(n1643), .D(n20), .Q(cmd_data_q[285]));
Q_FDP4EP \cmd_data_q_REG[284] ( .CK(clk), .CE(n1642), .R(n1643), .D(n21), .Q(cmd_data_q[284]));
Q_FDP4EP \cmd_data_q_REG[283] ( .CK(clk), .CE(n1642), .R(n1643), .D(n22), .Q(cmd_data_q[283]));
Q_FDP4EP \cmd_data_q_REG[282] ( .CK(clk), .CE(n1642), .R(n1643), .D(n23), .Q(cmd_data_q[282]));
Q_FDP4EP \cmd_data_q_REG[281] ( .CK(clk), .CE(n1642), .R(n1643), .D(n24), .Q(cmd_data_q[281]));
Q_FDP4EP \cmd_data_q_REG[280] ( .CK(clk), .CE(n1642), .R(n1643), .D(n25), .Q(cmd_data_q[280]));
Q_FDP4EP \cmd_data_q_REG[279] ( .CK(clk), .CE(n1642), .R(n1643), .D(n26), .Q(cmd_data_q[279]));
Q_FDP4EP \cmd_data_q_REG[278] ( .CK(clk), .CE(n1642), .R(n1643), .D(n27), .Q(cmd_data_q[278]));
Q_FDP4EP \cmd_data_q_REG[277] ( .CK(clk), .CE(n1642), .R(n1643), .D(n28), .Q(cmd_data_q[277]));
Q_FDP4EP \cmd_data_q_REG[276] ( .CK(clk), .CE(n1642), .R(n1643), .D(n29), .Q(cmd_data_q[276]));
Q_FDP4EP \cmd_data_q_REG[275] ( .CK(clk), .CE(n1642), .R(n1643), .D(n30), .Q(cmd_data_q[275]));
Q_FDP4EP \cmd_data_q_REG[274] ( .CK(clk), .CE(n1642), .R(n1643), .D(n31), .Q(cmd_data_q[274]));
Q_FDP4EP \cmd_data_q_REG[273] ( .CK(clk), .CE(n1642), .R(n1643), .D(n32), .Q(cmd_data_q[273]));
Q_FDP4EP \cmd_data_q_REG[272] ( .CK(clk), .CE(n1642), .R(n1643), .D(n33), .Q(cmd_data_q[272]));
Q_FDP4EP \cmd_data_q_REG[271] ( .CK(clk), .CE(n1642), .R(n1643), .D(n34), .Q(cmd_data_q[271]));
Q_FDP4EP \cmd_data_q_REG[270] ( .CK(clk), .CE(n1642), .R(n1643), .D(n35), .Q(cmd_data_q[270]));
Q_FDP4EP \cmd_data_q_REG[269] ( .CK(clk), .CE(n1642), .R(n1643), .D(n36), .Q(cmd_data_q[269]));
Q_FDP4EP \cmd_data_q_REG[268] ( .CK(clk), .CE(n1642), .R(n1643), .D(n37), .Q(cmd_data_q[268]));
Q_FDP4EP \cmd_data_q_REG[267] ( .CK(clk), .CE(n1642), .R(n1643), .D(n38), .Q(cmd_data_q[267]));
Q_FDP4EP \cmd_data_q_REG[266] ( .CK(clk), .CE(n1642), .R(n1643), .D(n39), .Q(cmd_data_q[266]));
Q_FDP4EP \cmd_data_q_REG[265] ( .CK(clk), .CE(n1642), .R(n1643), .D(n40), .Q(cmd_data_q[265]));
Q_FDP4EP \cmd_data_q_REG[264] ( .CK(clk), .CE(n1642), .R(n1643), .D(n41), .Q(cmd_data_q[264]));
Q_FDP4EP \cmd_data_q_REG[263] ( .CK(clk), .CE(n1642), .R(n1643), .D(n42), .Q(cmd_data_q[263]));
Q_FDP4EP \cmd_data_q_REG[262] ( .CK(clk), .CE(n1642), .R(n1643), .D(n43), .Q(cmd_data_q[262]));
Q_FDP4EP \cmd_data_q_REG[261] ( .CK(clk), .CE(n1642), .R(n1643), .D(n44), .Q(cmd_data_q[261]));
Q_FDP4EP \cmd_data_q_REG[260] ( .CK(clk), .CE(n1642), .R(n1643), .D(n45), .Q(cmd_data_q[260]));
Q_FDP4EP \cmd_data_q_REG[259] ( .CK(clk), .CE(n1642), .R(n1643), .D(n46), .Q(cmd_data_q[259]));
Q_FDP4EP \cmd_data_q_REG[258] ( .CK(clk), .CE(n1642), .R(n1643), .D(n47), .Q(cmd_data_q[258]));
Q_FDP4EP \cmd_data_q_REG[257] ( .CK(clk), .CE(n1642), .R(n1643), .D(n48), .Q(cmd_data_q[257]));
Q_FDP4EP \cmd_data_q_REG[256] ( .CK(clk), .CE(n1642), .R(n1643), .D(n49), .Q(cmd_data_q[256]));
Q_FDP4EP \cmd_data_q_REG[255] ( .CK(clk), .CE(n1642), .R(n1643), .D(n50), .Q(cmd_data_q[255]));
Q_FDP4EP \cmd_data_q_REG[254] ( .CK(clk), .CE(n1642), .R(n1643), .D(n51), .Q(cmd_data_q[254]));
Q_FDP4EP \cmd_data_q_REG[253] ( .CK(clk), .CE(n1642), .R(n1643), .D(n52), .Q(cmd_data_q[253]));
Q_FDP4EP \cmd_data_q_REG[252] ( .CK(clk), .CE(n1642), .R(n1643), .D(n53), .Q(cmd_data_q[252]));
Q_FDP4EP \cmd_data_q_REG[251] ( .CK(clk), .CE(n1642), .R(n1643), .D(n54), .Q(cmd_data_q[251]));
Q_FDP4EP \cmd_data_q_REG[250] ( .CK(clk), .CE(n1642), .R(n1643), .D(n55), .Q(cmd_data_q[250]));
Q_FDP4EP \cmd_data_q_REG[249] ( .CK(clk), .CE(n1642), .R(n1643), .D(n56), .Q(cmd_data_q[249]));
Q_FDP4EP \cmd_data_q_REG[248] ( .CK(clk), .CE(n1642), .R(n1643), .D(n57), .Q(cmd_data_q[248]));
Q_FDP4EP \cmd_data_q_REG[247] ( .CK(clk), .CE(n1642), .R(n1643), .D(n58), .Q(cmd_data_q[247]));
Q_FDP4EP \cmd_data_q_REG[246] ( .CK(clk), .CE(n1642), .R(n1643), .D(n59), .Q(cmd_data_q[246]));
Q_FDP4EP \cmd_data_q_REG[245] ( .CK(clk), .CE(n1642), .R(n1643), .D(n60), .Q(cmd_data_q[245]));
Q_FDP4EP \cmd_data_q_REG[244] ( .CK(clk), .CE(n1642), .R(n1643), .D(n61), .Q(cmd_data_q[244]));
Q_FDP4EP \cmd_data_q_REG[243] ( .CK(clk), .CE(n1642), .R(n1643), .D(n62), .Q(cmd_data_q[243]));
Q_FDP4EP \cmd_data_q_REG[242] ( .CK(clk), .CE(n1642), .R(n1643), .D(n63), .Q(cmd_data_q[242]));
Q_FDP4EP \cmd_data_q_REG[241] ( .CK(clk), .CE(n1642), .R(n1643), .D(n64), .Q(cmd_data_q[241]));
Q_FDP4EP \cmd_data_q_REG[240] ( .CK(clk), .CE(n1642), .R(n1643), .D(n65), .Q(cmd_data_q[240]));
Q_FDP4EP \cmd_data_q_REG[239] ( .CK(clk), .CE(n1642), .R(n1643), .D(n66), .Q(cmd_data_q[239]));
Q_FDP4EP \cmd_data_q_REG[238] ( .CK(clk), .CE(n1642), .R(n1643), .D(n67), .Q(cmd_data_q[238]));
Q_FDP4EP \cmd_data_q_REG[237] ( .CK(clk), .CE(n1642), .R(n1643), .D(n68), .Q(cmd_data_q[237]));
Q_FDP4EP \cmd_data_q_REG[236] ( .CK(clk), .CE(n1642), .R(n1643), .D(n69), .Q(cmd_data_q[236]));
Q_FDP4EP \cmd_data_q_REG[235] ( .CK(clk), .CE(n1642), .R(n1643), .D(n70), .Q(cmd_data_q[235]));
Q_FDP4EP \cmd_data_q_REG[234] ( .CK(clk), .CE(n1642), .R(n1643), .D(n71), .Q(cmd_data_q[234]));
Q_FDP4EP \cmd_data_q_REG[233] ( .CK(clk), .CE(n1642), .R(n1643), .D(n72), .Q(cmd_data_q[233]));
Q_FDP4EP \cmd_data_q_REG[232] ( .CK(clk), .CE(n1642), .R(n1643), .D(n73), .Q(cmd_data_q[232]));
Q_FDP4EP \cmd_data_q_REG[231] ( .CK(clk), .CE(n1642), .R(n1643), .D(n74), .Q(cmd_data_q[231]));
Q_FDP4EP \cmd_data_q_REG[230] ( .CK(clk), .CE(n1642), .R(n1643), .D(n75), .Q(cmd_data_q[230]));
Q_FDP4EP \cmd_data_q_REG[229] ( .CK(clk), .CE(n1642), .R(n1643), .D(n76), .Q(cmd_data_q[229]));
Q_FDP4EP \cmd_data_q_REG[228] ( .CK(clk), .CE(n1642), .R(n1643), .D(n77), .Q(cmd_data_q[228]));
Q_FDP4EP \cmd_data_q_REG[227] ( .CK(clk), .CE(n1642), .R(n1643), .D(n78), .Q(cmd_data_q[227]));
Q_FDP4EP \cmd_data_q_REG[226] ( .CK(clk), .CE(n1642), .R(n1643), .D(n79), .Q(cmd_data_q[226]));
Q_FDP4EP \cmd_data_q_REG[225] ( .CK(clk), .CE(n1642), .R(n1643), .D(n80), .Q(cmd_data_q[225]));
Q_FDP4EP \cmd_data_q_REG[224] ( .CK(clk), .CE(n1642), .R(n1643), .D(n81), .Q(cmd_data_q[224]));
Q_FDP4EP \cmd_data_q_REG[223] ( .CK(clk), .CE(n1642), .R(n1643), .D(n82), .Q(cmd_data_q[223]));
Q_FDP4EP \cmd_data_q_REG[222] ( .CK(clk), .CE(n1642), .R(n1643), .D(n83), .Q(cmd_data_q[222]));
Q_FDP4EP \cmd_data_q_REG[221] ( .CK(clk), .CE(n1642), .R(n1643), .D(n84), .Q(cmd_data_q[221]));
Q_FDP4EP \cmd_data_q_REG[220] ( .CK(clk), .CE(n1642), .R(n1643), .D(n85), .Q(cmd_data_q[220]));
Q_FDP4EP \cmd_data_q_REG[219] ( .CK(clk), .CE(n1642), .R(n1643), .D(n86), .Q(cmd_data_q[219]));
Q_FDP4EP \cmd_data_q_REG[218] ( .CK(clk), .CE(n1642), .R(n1643), .D(n87), .Q(cmd_data_q[218]));
Q_FDP4EP \cmd_data_q_REG[217] ( .CK(clk), .CE(n1642), .R(n1643), .D(n88), .Q(cmd_data_q[217]));
Q_FDP4EP \cmd_data_q_REG[216] ( .CK(clk), .CE(n1642), .R(n1643), .D(n89), .Q(cmd_data_q[216]));
Q_FDP4EP \cmd_data_q_REG[215] ( .CK(clk), .CE(n1642), .R(n1643), .D(n90), .Q(cmd_data_q[215]));
Q_FDP4EP \cmd_data_q_REG[214] ( .CK(clk), .CE(n1642), .R(n1643), .D(n91), .Q(cmd_data_q[214]));
Q_FDP4EP \cmd_data_q_REG[213] ( .CK(clk), .CE(n1642), .R(n1643), .D(n92), .Q(cmd_data_q[213]));
Q_FDP4EP \cmd_data_q_REG[212] ( .CK(clk), .CE(n1642), .R(n1643), .D(n93), .Q(cmd_data_q[212]));
Q_FDP4EP \cmd_data_q_REG[211] ( .CK(clk), .CE(n1642), .R(n1643), .D(n94), .Q(cmd_data_q[211]));
Q_FDP4EP \cmd_data_q_REG[210] ( .CK(clk), .CE(n1642), .R(n1643), .D(n95), .Q(cmd_data_q[210]));
Q_FDP4EP \cmd_data_q_REG[209] ( .CK(clk), .CE(n1642), .R(n1643), .D(n96), .Q(cmd_data_q[209]));
Q_FDP4EP \cmd_data_q_REG[208] ( .CK(clk), .CE(n1642), .R(n1643), .D(n97), .Q(cmd_data_q[208]));
Q_FDP4EP \cmd_data_q_REG[207] ( .CK(clk), .CE(n1642), .R(n1643), .D(n98), .Q(cmd_data_q[207]));
Q_FDP4EP \cmd_data_q_REG[206] ( .CK(clk), .CE(n1642), .R(n1643), .D(n99), .Q(cmd_data_q[206]));
Q_FDP4EP \cmd_data_q_REG[205] ( .CK(clk), .CE(n1642), .R(n1643), .D(n100), .Q(cmd_data_q[205]));
Q_FDP4EP \cmd_data_q_REG[204] ( .CK(clk), .CE(n1642), .R(n1643), .D(n101), .Q(cmd_data_q[204]));
Q_FDP4EP \cmd_data_q_REG[203] ( .CK(clk), .CE(n1642), .R(n1643), .D(n102), .Q(cmd_data_q[203]));
Q_FDP4EP \cmd_data_q_REG[202] ( .CK(clk), .CE(n1642), .R(n1643), .D(n103), .Q(cmd_data_q[202]));
Q_FDP4EP \cmd_data_q_REG[201] ( .CK(clk), .CE(n1642), .R(n1643), .D(n104), .Q(cmd_data_q[201]));
Q_FDP4EP \cmd_data_q_REG[200] ( .CK(clk), .CE(n1642), .R(n1643), .D(n105), .Q(cmd_data_q[200]));
Q_FDP4EP \cmd_data_q_REG[199] ( .CK(clk), .CE(n1642), .R(n1643), .D(n106), .Q(cmd_data_q[199]));
Q_FDP4EP \cmd_data_q_REG[198] ( .CK(clk), .CE(n1642), .R(n1643), .D(n107), .Q(cmd_data_q[198]));
Q_FDP4EP \cmd_data_q_REG[197] ( .CK(clk), .CE(n1642), .R(n1643), .D(n108), .Q(cmd_data_q[197]));
Q_FDP4EP \cmd_data_q_REG[196] ( .CK(clk), .CE(n1642), .R(n1643), .D(n109), .Q(cmd_data_q[196]));
Q_FDP4EP \cmd_data_q_REG[195] ( .CK(clk), .CE(n1642), .R(n1643), .D(n110), .Q(cmd_data_q[195]));
Q_FDP4EP \cmd_data_q_REG[194] ( .CK(clk), .CE(n1642), .R(n1643), .D(n111), .Q(cmd_data_q[194]));
Q_FDP4EP \cmd_data_q_REG[193] ( .CK(clk), .CE(n1642), .R(n1643), .D(n112), .Q(cmd_data_q[193]));
Q_FDP4EP \cmd_data_q_REG[192] ( .CK(clk), .CE(n1642), .R(n1643), .D(n113), .Q(cmd_data_q[192]));
Q_FDP4EP \cmd_data_q_REG[191] ( .CK(clk), .CE(n1642), .R(n1643), .D(n114), .Q(cmd_data_q[191]));
Q_FDP4EP \cmd_data_q_REG[190] ( .CK(clk), .CE(n1642), .R(n1643), .D(n115), .Q(cmd_data_q[190]));
Q_FDP4EP \cmd_data_q_REG[189] ( .CK(clk), .CE(n1642), .R(n1643), .D(n116), .Q(cmd_data_q[189]));
Q_FDP4EP \cmd_data_q_REG[188] ( .CK(clk), .CE(n1642), .R(n1643), .D(n117), .Q(cmd_data_q[188]));
Q_FDP4EP \cmd_data_q_REG[187] ( .CK(clk), .CE(n1642), .R(n1643), .D(n118), .Q(cmd_data_q[187]));
Q_FDP4EP \cmd_data_q_REG[186] ( .CK(clk), .CE(n1642), .R(n1643), .D(n119), .Q(cmd_data_q[186]));
Q_FDP4EP \cmd_data_q_REG[185] ( .CK(clk), .CE(n1642), .R(n1643), .D(n120), .Q(cmd_data_q[185]));
Q_FDP4EP \cmd_data_q_REG[184] ( .CK(clk), .CE(n1642), .R(n1643), .D(n121), .Q(cmd_data_q[184]));
Q_FDP4EP \cmd_data_q_REG[183] ( .CK(clk), .CE(n1642), .R(n1643), .D(n122), .Q(cmd_data_q[183]));
Q_FDP4EP \cmd_data_q_REG[182] ( .CK(clk), .CE(n1642), .R(n1643), .D(n123), .Q(cmd_data_q[182]));
Q_FDP4EP \cmd_data_q_REG[181] ( .CK(clk), .CE(n1642), .R(n1643), .D(n124), .Q(cmd_data_q[181]));
Q_FDP4EP \cmd_data_q_REG[180] ( .CK(clk), .CE(n1642), .R(n1643), .D(n125), .Q(cmd_data_q[180]));
Q_FDP4EP \cmd_data_q_REG[179] ( .CK(clk), .CE(n1642), .R(n1643), .D(n126), .Q(cmd_data_q[179]));
Q_FDP4EP \cmd_data_q_REG[178] ( .CK(clk), .CE(n1642), .R(n1643), .D(n127), .Q(cmd_data_q[178]));
Q_FDP4EP \cmd_data_q_REG[177] ( .CK(clk), .CE(n1642), .R(n1643), .D(n128), .Q(cmd_data_q[177]));
Q_FDP4EP \cmd_data_q_REG[176] ( .CK(clk), .CE(n1642), .R(n1643), .D(n129), .Q(cmd_data_q[176]));
Q_FDP4EP \cmd_data_q_REG[175] ( .CK(clk), .CE(n1642), .R(n1643), .D(n130), .Q(cmd_data_q[175]));
Q_FDP4EP \cmd_data_q_REG[174] ( .CK(clk), .CE(n1642), .R(n1643), .D(n131), .Q(cmd_data_q[174]));
Q_FDP4EP \cmd_data_q_REG[173] ( .CK(clk), .CE(n1642), .R(n1643), .D(n132), .Q(cmd_data_q[173]));
Q_FDP4EP \cmd_data_q_REG[172] ( .CK(clk), .CE(n1642), .R(n1643), .D(n133), .Q(cmd_data_q[172]));
Q_FDP4EP \cmd_data_q_REG[171] ( .CK(clk), .CE(n1642), .R(n1643), .D(n134), .Q(cmd_data_q[171]));
Q_FDP4EP \cmd_data_q_REG[170] ( .CK(clk), .CE(n1642), .R(n1643), .D(n135), .Q(cmd_data_q[170]));
Q_FDP4EP \cmd_data_q_REG[169] ( .CK(clk), .CE(n1642), .R(n1643), .D(n136), .Q(cmd_data_q[169]));
Q_FDP4EP \cmd_data_q_REG[168] ( .CK(clk), .CE(n1642), .R(n1643), .D(n137), .Q(cmd_data_q[168]));
Q_FDP4EP \cmd_data_q_REG[167] ( .CK(clk), .CE(n1642), .R(n1643), .D(n138), .Q(cmd_data_q[167]));
Q_FDP4EP \cmd_data_q_REG[166] ( .CK(clk), .CE(n1642), .R(n1643), .D(n139), .Q(cmd_data_q[166]));
Q_FDP4EP \cmd_data_q_REG[165] ( .CK(clk), .CE(n1642), .R(n1643), .D(n140), .Q(cmd_data_q[165]));
Q_FDP4EP \cmd_data_q_REG[164] ( .CK(clk), .CE(n1642), .R(n1643), .D(n141), .Q(cmd_data_q[164]));
Q_FDP4EP \cmd_data_q_REG[163] ( .CK(clk), .CE(n1642), .R(n1643), .D(n142), .Q(cmd_data_q[163]));
Q_FDP4EP \cmd_data_q_REG[162] ( .CK(clk), .CE(n1642), .R(n1643), .D(n143), .Q(cmd_data_q[162]));
Q_FDP4EP \cmd_data_q_REG[161] ( .CK(clk), .CE(n1642), .R(n1643), .D(n144), .Q(cmd_data_q[161]));
Q_FDP4EP \cmd_data_q_REG[160] ( .CK(clk), .CE(n1642), .R(n1643), .D(n145), .Q(cmd_data_q[160]));
Q_FDP4EP \cmd_data_q_REG[159] ( .CK(clk), .CE(n1642), .R(n1643), .D(n146), .Q(cmd_data_q[159]));
Q_FDP4EP \cmd_data_q_REG[158] ( .CK(clk), .CE(n1642), .R(n1643), .D(n147), .Q(cmd_data_q[158]));
Q_FDP4EP \cmd_data_q_REG[157] ( .CK(clk), .CE(n1642), .R(n1643), .D(n148), .Q(cmd_data_q[157]));
Q_FDP4EP \cmd_data_q_REG[156] ( .CK(clk), .CE(n1642), .R(n1643), .D(n149), .Q(cmd_data_q[156]));
Q_FDP4EP \cmd_data_q_REG[155] ( .CK(clk), .CE(n1642), .R(n1643), .D(n150), .Q(cmd_data_q[155]));
Q_FDP4EP \cmd_data_q_REG[154] ( .CK(clk), .CE(n1642), .R(n1643), .D(n151), .Q(cmd_data_q[154]));
Q_FDP4EP \cmd_data_q_REG[153] ( .CK(clk), .CE(n1642), .R(n1643), .D(n152), .Q(cmd_data_q[153]));
Q_FDP4EP \cmd_data_q_REG[152] ( .CK(clk), .CE(n1642), .R(n1643), .D(n153), .Q(cmd_data_q[152]));
Q_FDP4EP \cmd_data_q_REG[151] ( .CK(clk), .CE(n1642), .R(n1643), .D(n154), .Q(cmd_data_q[151]));
Q_FDP4EP \cmd_data_q_REG[150] ( .CK(clk), .CE(n1642), .R(n1643), .D(n155), .Q(cmd_data_q[150]));
Q_FDP4EP \cmd_data_q_REG[149] ( .CK(clk), .CE(n1642), .R(n1643), .D(n156), .Q(cmd_data_q[149]));
Q_FDP4EP \cmd_data_q_REG[148] ( .CK(clk), .CE(n1642), .R(n1643), .D(n157), .Q(cmd_data_q[148]));
Q_FDP4EP \cmd_data_q_REG[147] ( .CK(clk), .CE(n1642), .R(n1643), .D(n158), .Q(cmd_data_q[147]));
Q_FDP4EP \cmd_data_q_REG[146] ( .CK(clk), .CE(n1642), .R(n1643), .D(n159), .Q(cmd_data_q[146]));
Q_FDP4EP \cmd_data_q_REG[145] ( .CK(clk), .CE(n1642), .R(n1643), .D(n160), .Q(cmd_data_q[145]));
Q_FDP4EP \cmd_data_q_REG[144] ( .CK(clk), .CE(n1642), .R(n1643), .D(n161), .Q(cmd_data_q[144]));
Q_FDP4EP \cmd_data_q_REG[143] ( .CK(clk), .CE(n1642), .R(n1643), .D(n162), .Q(cmd_data_q[143]));
Q_FDP4EP \cmd_data_q_REG[142] ( .CK(clk), .CE(n1642), .R(n1643), .D(n163), .Q(cmd_data_q[142]));
Q_FDP4EP \cmd_data_q_REG[141] ( .CK(clk), .CE(n1642), .R(n1643), .D(n164), .Q(cmd_data_q[141]));
Q_FDP4EP \cmd_data_q_REG[140] ( .CK(clk), .CE(n1642), .R(n1643), .D(n165), .Q(cmd_data_q[140]));
Q_FDP4EP \cmd_data_q_REG[139] ( .CK(clk), .CE(n1642), .R(n1643), .D(n166), .Q(cmd_data_q[139]));
Q_FDP4EP \cmd_data_q_REG[138] ( .CK(clk), .CE(n1642), .R(n1643), .D(n167), .Q(cmd_data_q[138]));
Q_FDP4EP \cmd_data_q_REG[137] ( .CK(clk), .CE(n1642), .R(n1643), .D(n168), .Q(cmd_data_q[137]));
Q_FDP4EP \cmd_data_q_REG[136] ( .CK(clk), .CE(n1642), .R(n1643), .D(n169), .Q(cmd_data_q[136]));
Q_FDP4EP \cmd_data_q_REG[135] ( .CK(clk), .CE(n1642), .R(n1643), .D(n170), .Q(cmd_data_q[135]));
Q_FDP4EP \cmd_data_q_REG[134] ( .CK(clk), .CE(n1642), .R(n1643), .D(n171), .Q(cmd_data_q[134]));
Q_FDP4EP \cmd_data_q_REG[133] ( .CK(clk), .CE(n1642), .R(n1643), .D(n172), .Q(cmd_data_q[133]));
Q_FDP4EP \cmd_data_q_REG[132] ( .CK(clk), .CE(n1642), .R(n1643), .D(n173), .Q(cmd_data_q[132]));
Q_FDP4EP \cmd_data_q_REG[131] ( .CK(clk), .CE(n1642), .R(n1643), .D(n174), .Q(cmd_data_q[131]));
Q_FDP4EP \cmd_data_q_REG[130] ( .CK(clk), .CE(n1642), .R(n1643), .D(n175), .Q(cmd_data_q[130]));
Q_FDP4EP \cmd_data_q_REG[129] ( .CK(clk), .CE(n1642), .R(n1643), .D(n176), .Q(cmd_data_q[129]));
Q_FDP4EP \cmd_data_q_REG[128] ( .CK(clk), .CE(n1642), .R(n1643), .D(n177), .Q(cmd_data_q[128]));
Q_FDP4EP \cmd_data_q_REG[127] ( .CK(clk), .CE(n1642), .R(n1643), .D(n178), .Q(cmd_data_q[127]));
Q_FDP4EP \cmd_data_q_REG[126] ( .CK(clk), .CE(n1642), .R(n1643), .D(n179), .Q(cmd_data_q[126]));
Q_FDP4EP \cmd_data_q_REG[125] ( .CK(clk), .CE(n1642), .R(n1643), .D(n180), .Q(cmd_data_q[125]));
Q_FDP4EP \cmd_data_q_REG[124] ( .CK(clk), .CE(n1642), .R(n1643), .D(n181), .Q(cmd_data_q[124]));
Q_FDP4EP \cmd_data_q_REG[123] ( .CK(clk), .CE(n1642), .R(n1643), .D(n182), .Q(cmd_data_q[123]));
Q_FDP4EP \cmd_data_q_REG[122] ( .CK(clk), .CE(n1642), .R(n1643), .D(n183), .Q(cmd_data_q[122]));
Q_FDP4EP \cmd_data_q_REG[121] ( .CK(clk), .CE(n1642), .R(n1643), .D(n184), .Q(cmd_data_q[121]));
Q_FDP4EP \cmd_data_q_REG[120] ( .CK(clk), .CE(n1642), .R(n1643), .D(n185), .Q(cmd_data_q[120]));
Q_FDP4EP \cmd_data_q_REG[119] ( .CK(clk), .CE(n1642), .R(n1643), .D(n186), .Q(cmd_data_q[119]));
Q_FDP4EP \cmd_data_q_REG[118] ( .CK(clk), .CE(n1642), .R(n1643), .D(n187), .Q(cmd_data_q[118]));
Q_FDP4EP \cmd_data_q_REG[117] ( .CK(clk), .CE(n1642), .R(n1643), .D(n188), .Q(cmd_data_q[117]));
Q_FDP4EP \cmd_data_q_REG[116] ( .CK(clk), .CE(n1642), .R(n1643), .D(n189), .Q(cmd_data_q[116]));
Q_FDP4EP \cmd_data_q_REG[115] ( .CK(clk), .CE(n1642), .R(n1643), .D(n190), .Q(cmd_data_q[115]));
Q_FDP4EP \cmd_data_q_REG[114] ( .CK(clk), .CE(n1642), .R(n1643), .D(n191), .Q(cmd_data_q[114]));
Q_FDP4EP \cmd_data_q_REG[113] ( .CK(clk), .CE(n1642), .R(n1643), .D(n192), .Q(cmd_data_q[113]));
Q_FDP4EP \cmd_data_q_REG[112] ( .CK(clk), .CE(n1642), .R(n1643), .D(n193), .Q(cmd_data_q[112]));
Q_FDP4EP \cmd_data_q_REG[111] ( .CK(clk), .CE(n1642), .R(n1643), .D(n194), .Q(cmd_data_q[111]));
Q_FDP4EP \cmd_data_q_REG[110] ( .CK(clk), .CE(n1642), .R(n1643), .D(n195), .Q(cmd_data_q[110]));
Q_FDP4EP \cmd_data_q_REG[109] ( .CK(clk), .CE(n1642), .R(n1643), .D(n196), .Q(cmd_data_q[109]));
Q_FDP4EP \cmd_data_q_REG[108] ( .CK(clk), .CE(n1642), .R(n1643), .D(n197), .Q(cmd_data_q[108]));
Q_FDP4EP \cmd_data_q_REG[107] ( .CK(clk), .CE(n1642), .R(n1643), .D(n198), .Q(cmd_data_q[107]));
Q_FDP4EP \cmd_data_q_REG[106] ( .CK(clk), .CE(n1642), .R(n1643), .D(n199), .Q(cmd_data_q[106]));
Q_FDP4EP \cmd_data_q_REG[105] ( .CK(clk), .CE(n1642), .R(n1643), .D(n200), .Q(cmd_data_q[105]));
Q_FDP4EP \cmd_data_q_REG[104] ( .CK(clk), .CE(n1642), .R(n1643), .D(n201), .Q(cmd_data_q[104]));
Q_FDP4EP \cmd_data_q_REG[103] ( .CK(clk), .CE(n1642), .R(n1643), .D(n202), .Q(cmd_data_q[103]));
Q_FDP4EP \cmd_data_q_REG[102] ( .CK(clk), .CE(n1642), .R(n1643), .D(n203), .Q(cmd_data_q[102]));
Q_FDP4EP \cmd_data_q_REG[101] ( .CK(clk), .CE(n1642), .R(n1643), .D(n204), .Q(cmd_data_q[101]));
Q_FDP4EP \cmd_data_q_REG[100] ( .CK(clk), .CE(n1642), .R(n1643), .D(n205), .Q(cmd_data_q[100]));
Q_FDP4EP \cmd_data_q_REG[99] ( .CK(clk), .CE(n1642), .R(n1643), .D(n206), .Q(cmd_data_q[99]));
Q_FDP4EP \cmd_data_q_REG[98] ( .CK(clk), .CE(n1642), .R(n1643), .D(n207), .Q(cmd_data_q[98]));
Q_FDP4EP \cmd_data_q_REG[97] ( .CK(clk), .CE(n1642), .R(n1643), .D(n208), .Q(cmd_data_q[97]));
Q_FDP4EP \cmd_data_q_REG[96] ( .CK(clk), .CE(n1642), .R(n1643), .D(n209), .Q(cmd_data_q[96]));
Q_FDP4EP \cmd_data_q_REG[95] ( .CK(clk), .CE(n1642), .R(n1643), .D(n210), .Q(cmd_data_q[95]));
Q_FDP4EP \cmd_data_q_REG[94] ( .CK(clk), .CE(n1642), .R(n1643), .D(n211), .Q(cmd_data_q[94]));
Q_FDP4EP \cmd_data_q_REG[93] ( .CK(clk), .CE(n1642), .R(n1643), .D(n212), .Q(cmd_data_q[93]));
Q_FDP4EP \cmd_data_q_REG[92] ( .CK(clk), .CE(n1642), .R(n1643), .D(n213), .Q(cmd_data_q[92]));
Q_FDP4EP \cmd_data_q_REG[91] ( .CK(clk), .CE(n1642), .R(n1643), .D(n214), .Q(cmd_data_q[91]));
Q_FDP4EP \cmd_data_q_REG[90] ( .CK(clk), .CE(n1642), .R(n1643), .D(n215), .Q(cmd_data_q[90]));
Q_FDP4EP \cmd_data_q_REG[89] ( .CK(clk), .CE(n1642), .R(n1643), .D(n216), .Q(cmd_data_q[89]));
Q_FDP4EP \cmd_data_q_REG[88] ( .CK(clk), .CE(n1642), .R(n1643), .D(n217), .Q(cmd_data_q[88]));
Q_FDP4EP \cmd_data_q_REG[87] ( .CK(clk), .CE(n1642), .R(n1643), .D(n218), .Q(cmd_data_q[87]));
Q_FDP4EP \cmd_data_q_REG[86] ( .CK(clk), .CE(n1642), .R(n1643), .D(n219), .Q(cmd_data_q[86]));
Q_FDP4EP \cmd_data_q_REG[85] ( .CK(clk), .CE(n1642), .R(n1643), .D(n220), .Q(cmd_data_q[85]));
Q_FDP4EP \cmd_data_q_REG[84] ( .CK(clk), .CE(n1642), .R(n1643), .D(n221), .Q(cmd_data_q[84]));
Q_FDP4EP \cmd_data_q_REG[83] ( .CK(clk), .CE(n1642), .R(n1643), .D(n222), .Q(cmd_data_q[83]));
Q_FDP4EP \cmd_data_q_REG[82] ( .CK(clk), .CE(n1642), .R(n1643), .D(n223), .Q(cmd_data_q[82]));
Q_FDP4EP \cmd_data_q_REG[81] ( .CK(clk), .CE(n1642), .R(n1643), .D(n224), .Q(cmd_data_q[81]));
Q_FDP4EP \cmd_data_q_REG[80] ( .CK(clk), .CE(n1642), .R(n1643), .D(n225), .Q(cmd_data_q[80]));
Q_FDP4EP \cmd_data_q_REG[79] ( .CK(clk), .CE(n1642), .R(n1643), .D(n226), .Q(cmd_data_q[79]));
Q_FDP4EP \cmd_data_q_REG[78] ( .CK(clk), .CE(n1642), .R(n1643), .D(n227), .Q(cmd_data_q[78]));
Q_FDP4EP \cmd_data_q_REG[77] ( .CK(clk), .CE(n1642), .R(n1643), .D(n228), .Q(cmd_data_q[77]));
Q_FDP4EP \cmd_data_q_REG[76] ( .CK(clk), .CE(n1642), .R(n1643), .D(n229), .Q(cmd_data_q[76]));
Q_FDP4EP \cmd_data_q_REG[75] ( .CK(clk), .CE(n1642), .R(n1643), .D(n230), .Q(cmd_data_q[75]));
Q_FDP4EP \cmd_data_q_REG[74] ( .CK(clk), .CE(n1642), .R(n1643), .D(n231), .Q(cmd_data_q[74]));
Q_FDP4EP \cmd_data_q_REG[73] ( .CK(clk), .CE(n1642), .R(n1643), .D(n232), .Q(cmd_data_q[73]));
Q_FDP4EP \cmd_data_q_REG[72] ( .CK(clk), .CE(n1642), .R(n1643), .D(n233), .Q(cmd_data_q[72]));
Q_FDP4EP \cmd_data_q_REG[71] ( .CK(clk), .CE(n1642), .R(n1643), .D(n234), .Q(cmd_data_q[71]));
Q_FDP4EP \cmd_data_q_REG[70] ( .CK(clk), .CE(n1642), .R(n1643), .D(n235), .Q(cmd_data_q[70]));
Q_FDP4EP \cmd_data_q_REG[69] ( .CK(clk), .CE(n1642), .R(n1643), .D(n236), .Q(cmd_data_q[69]));
Q_FDP4EP \cmd_data_q_REG[68] ( .CK(clk), .CE(n1642), .R(n1643), .D(n237), .Q(cmd_data_q[68]));
Q_FDP4EP \cmd_data_q_REG[67] ( .CK(clk), .CE(n1642), .R(n1643), .D(n238), .Q(cmd_data_q[67]));
Q_FDP4EP \cmd_data_q_REG[66] ( .CK(clk), .CE(n1642), .R(n1643), .D(n239), .Q(cmd_data_q[66]));
Q_FDP4EP \cmd_data_q_REG[65] ( .CK(clk), .CE(n1642), .R(n1643), .D(n240), .Q(cmd_data_q[65]));
Q_FDP4EP \cmd_data_q_REG[64] ( .CK(clk), .CE(n1642), .R(n1643), .D(n241), .Q(cmd_data_q[64]));
Q_FDP4EP \cmd_data_q_REG[63] ( .CK(clk), .CE(n1642), .R(n1643), .D(n242), .Q(cmd_data_q[63]));
Q_FDP4EP \cmd_data_q_REG[62] ( .CK(clk), .CE(n1642), .R(n1643), .D(n243), .Q(cmd_data_q[62]));
Q_FDP4EP \cmd_data_q_REG[61] ( .CK(clk), .CE(n1642), .R(n1643), .D(n244), .Q(cmd_data_q[61]));
Q_FDP4EP \cmd_data_q_REG[60] ( .CK(clk), .CE(n1642), .R(n1643), .D(n245), .Q(cmd_data_q[60]));
Q_FDP4EP \cmd_data_q_REG[59] ( .CK(clk), .CE(n1642), .R(n1643), .D(n246), .Q(cmd_data_q[59]));
Q_FDP4EP \cmd_data_q_REG[58] ( .CK(clk), .CE(n1642), .R(n1643), .D(n247), .Q(cmd_data_q[58]));
Q_FDP4EP \cmd_data_q_REG[57] ( .CK(clk), .CE(n1642), .R(n1643), .D(n248), .Q(cmd_data_q[57]));
Q_FDP4EP \cmd_data_q_REG[56] ( .CK(clk), .CE(n1642), .R(n1643), .D(n249), .Q(cmd_data_q[56]));
Q_FDP4EP \cmd_data_q_REG[55] ( .CK(clk), .CE(n1642), .R(n1643), .D(n250), .Q(cmd_data_q[55]));
Q_FDP4EP \cmd_data_q_REG[54] ( .CK(clk), .CE(n1642), .R(n1643), .D(n251), .Q(cmd_data_q[54]));
Q_FDP4EP \cmd_data_q_REG[53] ( .CK(clk), .CE(n1642), .R(n1643), .D(n252), .Q(cmd_data_q[53]));
Q_FDP4EP \cmd_data_q_REG[52] ( .CK(clk), .CE(n1642), .R(n1643), .D(n253), .Q(cmd_data_q[52]));
Q_FDP4EP \cmd_data_q_REG[51] ( .CK(clk), .CE(n1642), .R(n1643), .D(n254), .Q(cmd_data_q[51]));
Q_FDP4EP \cmd_data_q_REG[50] ( .CK(clk), .CE(n1642), .R(n1643), .D(n255), .Q(cmd_data_q[50]));
Q_FDP4EP \cmd_data_q_REG[49] ( .CK(clk), .CE(n1642), .R(n1643), .D(n256), .Q(cmd_data_q[49]));
Q_FDP4EP \cmd_data_q_REG[48] ( .CK(clk), .CE(n1642), .R(n1643), .D(n257), .Q(cmd_data_q[48]));
Q_FDP4EP \cmd_data_q_REG[47] ( .CK(clk), .CE(n1642), .R(n1643), .D(n258), .Q(cmd_data_q[47]));
Q_FDP4EP \cmd_data_q_REG[46] ( .CK(clk), .CE(n1642), .R(n1643), .D(n259), .Q(cmd_data_q[46]));
Q_FDP4EP \cmd_data_q_REG[45] ( .CK(clk), .CE(n1642), .R(n1643), .D(n260), .Q(cmd_data_q[45]));
Q_FDP4EP \cmd_data_q_REG[44] ( .CK(clk), .CE(n1642), .R(n1643), .D(n261), .Q(cmd_data_q[44]));
Q_FDP4EP \cmd_data_q_REG[43] ( .CK(clk), .CE(n1642), .R(n1643), .D(n262), .Q(cmd_data_q[43]));
Q_FDP4EP \cmd_data_q_REG[42] ( .CK(clk), .CE(n1642), .R(n1643), .D(n263), .Q(cmd_data_q[42]));
Q_FDP4EP \cmd_data_q_REG[41] ( .CK(clk), .CE(n1642), .R(n1643), .D(n264), .Q(cmd_data_q[41]));
Q_FDP4EP \cmd_data_q_REG[40] ( .CK(clk), .CE(n1642), .R(n1643), .D(n265), .Q(cmd_data_q[40]));
Q_FDP4EP \cmd_data_q_REG[39] ( .CK(clk), .CE(n1642), .R(n1643), .D(n266), .Q(cmd_data_q[39]));
Q_FDP4EP \cmd_data_q_REG[38] ( .CK(clk), .CE(n1642), .R(n1643), .D(n267), .Q(cmd_data_q[38]));
Q_FDP4EP \cmd_data_q_REG[37] ( .CK(clk), .CE(n1642), .R(n1643), .D(n268), .Q(cmd_data_q[37]));
Q_FDP4EP \cmd_data_q_REG[36] ( .CK(clk), .CE(n1642), .R(n1643), .D(n269), .Q(cmd_data_q[36]));
Q_FDP4EP \cmd_data_q_REG[35] ( .CK(clk), .CE(n1642), .R(n1643), .D(n270), .Q(cmd_data_q[35]));
Q_FDP4EP \cmd_data_q_REG[34] ( .CK(clk), .CE(n1642), .R(n1643), .D(n271), .Q(cmd_data_q[34]));
Q_FDP4EP \cmd_data_q_REG[33] ( .CK(clk), .CE(n1642), .R(n1643), .D(n272), .Q(cmd_data_q[33]));
Q_FDP4EP \cmd_data_q_REG[32] ( .CK(clk), .CE(n1642), .R(n1643), .D(n273), .Q(cmd_data_q[32]));
Q_FDP4EP \cmd_data_q_REG[31] ( .CK(clk), .CE(n1642), .R(n1643), .D(n274), .Q(cmd_data_q[31]));
Q_FDP4EP \cmd_data_q_REG[30] ( .CK(clk), .CE(n1642), .R(n1643), .D(n275), .Q(cmd_data_q[30]));
Q_FDP4EP \cmd_data_q_REG[29] ( .CK(clk), .CE(n1642), .R(n1643), .D(n276), .Q(cmd_data_q[29]));
Q_FDP4EP \cmd_data_q_REG[28] ( .CK(clk), .CE(n1642), .R(n1643), .D(n277), .Q(cmd_data_q[28]));
Q_FDP4EP \cmd_data_q_REG[27] ( .CK(clk), .CE(n1642), .R(n1643), .D(n278), .Q(cmd_data_q[27]));
Q_FDP4EP \cmd_data_q_REG[26] ( .CK(clk), .CE(n1642), .R(n1643), .D(n279), .Q(cmd_data_q[26]));
Q_FDP4EP \cmd_data_q_REG[25] ( .CK(clk), .CE(n1642), .R(n1643), .D(n280), .Q(cmd_data_q[25]));
Q_FDP4EP \cmd_data_q_REG[24] ( .CK(clk), .CE(n1642), .R(n1643), .D(n281), .Q(cmd_data_q[24]));
Q_FDP4EP \cmd_data_q_REG[23] ( .CK(clk), .CE(n1642), .R(n1643), .D(n282), .Q(cmd_data_q[23]));
Q_FDP4EP \cmd_data_q_REG[22] ( .CK(clk), .CE(n1642), .R(n1643), .D(n283), .Q(cmd_data_q[22]));
Q_FDP4EP \cmd_data_q_REG[21] ( .CK(clk), .CE(n1642), .R(n1643), .D(n284), .Q(cmd_data_q[21]));
Q_FDP4EP \cmd_data_q_REG[20] ( .CK(clk), .CE(n1642), .R(n1643), .D(n285), .Q(cmd_data_q[20]));
Q_FDP4EP \cmd_data_q_REG[19] ( .CK(clk), .CE(n1642), .R(n1643), .D(n286), .Q(cmd_data_q[19]));
Q_FDP4EP \cmd_data_q_REG[18] ( .CK(clk), .CE(n1642), .R(n1643), .D(n287), .Q(cmd_data_q[18]));
Q_FDP4EP \cmd_data_q_REG[17] ( .CK(clk), .CE(n1642), .R(n1643), .D(n288), .Q(cmd_data_q[17]));
Q_FDP4EP \cmd_data_q_REG[16] ( .CK(clk), .CE(n1642), .R(n1643), .D(n289), .Q(cmd_data_q[16]));
Q_FDP4EP \cmd_data_q_REG[15] ( .CK(clk), .CE(n1642), .R(n1643), .D(n290), .Q(cmd_data_q[15]));
Q_FDP4EP \cmd_data_q_REG[14] ( .CK(clk), .CE(n1642), .R(n1643), .D(n291), .Q(cmd_data_q[14]));
Q_FDP4EP \cmd_data_q_REG[13] ( .CK(clk), .CE(n1642), .R(n1643), .D(n292), .Q(cmd_data_q[13]));
Q_FDP4EP \cmd_data_q_REG[12] ( .CK(clk), .CE(n1642), .R(n1643), .D(n293), .Q(cmd_data_q[12]));
Q_FDP4EP \cmd_data_q_REG[11] ( .CK(clk), .CE(n1642), .R(n1643), .D(n294), .Q(cmd_data_q[11]));
Q_FDP4EP \cmd_data_q_REG[10] ( .CK(clk), .CE(n1642), .R(n1643), .D(n295), .Q(cmd_data_q[10]));
Q_FDP4EP \cmd_data_q_REG[9] ( .CK(clk), .CE(n1642), .R(n1643), .D(n296), .Q(cmd_data_q[9]));
Q_FDP4EP \cmd_data_q_REG[8] ( .CK(clk), .CE(n1642), .R(n1643), .D(n297), .Q(cmd_data_q[8]));
Q_FDP4EP \cmd_data_q_REG[7] ( .CK(clk), .CE(n1642), .R(n1643), .D(n298), .Q(cmd_data_q[7]));
Q_FDP4EP \cmd_data_q_REG[6] ( .CK(clk), .CE(n1642), .R(n1643), .D(n299), .Q(cmd_data_q[6]));
Q_FDP4EP \cmd_data_q_REG[5] ( .CK(clk), .CE(n1642), .R(n1643), .D(n300), .Q(cmd_data_q[5]));
Q_FDP4EP \cmd_data_q_REG[4] ( .CK(clk), .CE(n1642), .R(n1643), .D(n301), .Q(cmd_data_q[4]));
Q_FDP4EP \cmd_data_q_REG[3] ( .CK(clk), .CE(n1642), .R(n1643), .D(n302), .Q(cmd_data_q[3]));
Q_FDP4EP \cmd_data_q_REG[2] ( .CK(clk), .CE(n1642), .R(n1643), .D(n303), .Q(cmd_data_q[2]));
Q_FDP4EP \cmd_data_q_REG[1] ( .CK(clk), .CE(n1642), .R(n1643), .D(n304), .Q(cmd_data_q[1]));
Q_FDP4EP \cmd_data_q_REG[0] ( .CK(clk), .CE(n1642), .R(n1643), .D(n305), .Q(cmd_data_q[0]));
endmodule
