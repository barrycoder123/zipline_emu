
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
(* celldefine = 1 *) 
module nx_fifo_xcm19 ( empty, full, underflow, overflow, used_slots, free_slots, 
	rdata, clk, rst_n, wen, ren, clear, wdata);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output empty;
output full;
output underflow;
output overflow;
output [1:0] used_slots;
output [1:0] free_slots;
output [105:0] rdata;
input clk;
input rst_n;
input wen;
input ren;
input clear;
input [105:0] wdata;
wire _zy_simnet_underflow_0_w$;
wire _zy_simnet_overflow_1_w$;
wire \depth_n._zy_simnet_overflow_3_w$ ;
wire \depth_n._zy_simnet_underflow_2_w$ ;
wire [0:0] \depth_n.wptr ;
wire [0:0] \depth_n.rptr ;
supply0 n113;
ixc_assign _zz_strnp_3 ( _zy_simnet_overflow_1_w$, overflow);
ixc_assign _zz_strnp_2 ( _zy_simnet_underflow_0_w$, underflow);
Q_MX02 U2 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][105] ), .A1(\depth_n.r_data[1][105] ), .Z(n1));
Q_MX02 U3 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][104] ), .A1(\depth_n.r_data[1][104] ), .Z(n2));
Q_MX02 U4 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][103] ), .A1(\depth_n.r_data[1][103] ), .Z(n3));
Q_MX02 U5 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][102] ), .A1(\depth_n.r_data[1][102] ), .Z(n4));
Q_MX02 U6 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][101] ), .A1(\depth_n.r_data[1][101] ), .Z(n5));
Q_MX02 U7 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][100] ), .A1(\depth_n.r_data[1][100] ), .Z(n6));
Q_MX02 U8 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][99] ), .A1(\depth_n.r_data[1][99] ), .Z(n7));
Q_MX02 U9 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][98] ), .A1(\depth_n.r_data[1][98] ), .Z(n8));
Q_MX02 U10 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][97] ), .A1(\depth_n.r_data[1][97] ), .Z(n9));
Q_MX02 U11 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][96] ), .A1(\depth_n.r_data[1][96] ), .Z(n10));
Q_MX02 U12 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][95] ), .A1(\depth_n.r_data[1][95] ), .Z(n11));
Q_MX02 U13 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][94] ), .A1(\depth_n.r_data[1][94] ), .Z(n12));
Q_MX02 U14 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][93] ), .A1(\depth_n.r_data[1][93] ), .Z(n13));
Q_MX02 U15 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][92] ), .A1(\depth_n.r_data[1][92] ), .Z(n14));
Q_MX02 U16 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][91] ), .A1(\depth_n.r_data[1][91] ), .Z(n15));
Q_MX02 U17 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][90] ), .A1(\depth_n.r_data[1][90] ), .Z(n16));
Q_MX02 U18 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][89] ), .A1(\depth_n.r_data[1][89] ), .Z(n17));
Q_MX02 U19 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][88] ), .A1(\depth_n.r_data[1][88] ), .Z(n18));
Q_MX02 U20 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][87] ), .A1(\depth_n.r_data[1][87] ), .Z(n19));
Q_MX02 U21 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][86] ), .A1(\depth_n.r_data[1][86] ), .Z(n20));
Q_MX02 U22 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][85] ), .A1(\depth_n.r_data[1][85] ), .Z(n21));
Q_MX02 U23 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][84] ), .A1(\depth_n.r_data[1][84] ), .Z(n22));
Q_MX02 U24 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][83] ), .A1(\depth_n.r_data[1][83] ), .Z(n23));
Q_MX02 U25 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][82] ), .A1(\depth_n.r_data[1][82] ), .Z(n24));
Q_MX02 U26 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][81] ), .A1(\depth_n.r_data[1][81] ), .Z(n25));
Q_MX02 U27 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][80] ), .A1(\depth_n.r_data[1][80] ), .Z(n26));
Q_MX02 U28 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][79] ), .A1(\depth_n.r_data[1][79] ), .Z(n27));
Q_MX02 U29 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][78] ), .A1(\depth_n.r_data[1][78] ), .Z(n28));
Q_MX02 U30 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][77] ), .A1(\depth_n.r_data[1][77] ), .Z(n29));
Q_MX02 U31 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][76] ), .A1(\depth_n.r_data[1][76] ), .Z(n30));
Q_MX02 U32 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][75] ), .A1(\depth_n.r_data[1][75] ), .Z(n31));
Q_MX02 U33 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][74] ), .A1(\depth_n.r_data[1][74] ), .Z(n32));
Q_MX02 U34 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][73] ), .A1(\depth_n.r_data[1][73] ), .Z(n33));
Q_MX02 U35 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][72] ), .A1(\depth_n.r_data[1][72] ), .Z(n34));
Q_MX02 U36 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][71] ), .A1(\depth_n.r_data[1][71] ), .Z(n35));
Q_MX02 U37 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][70] ), .A1(\depth_n.r_data[1][70] ), .Z(n36));
Q_MX02 U38 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][69] ), .A1(\depth_n.r_data[1][69] ), .Z(n37));
Q_MX02 U39 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][68] ), .A1(\depth_n.r_data[1][68] ), .Z(n38));
Q_MX02 U40 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][67] ), .A1(\depth_n.r_data[1][67] ), .Z(n39));
Q_MX02 U41 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][66] ), .A1(\depth_n.r_data[1][66] ), .Z(n40));
Q_MX02 U42 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][65] ), .A1(\depth_n.r_data[1][65] ), .Z(n41));
Q_MX02 U43 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][64] ), .A1(\depth_n.r_data[1][64] ), .Z(n42));
Q_MX02 U44 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][63] ), .A1(\depth_n.r_data[1][63] ), .Z(n43));
Q_MX02 U45 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][62] ), .A1(\depth_n.r_data[1][62] ), .Z(n44));
Q_MX02 U46 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][61] ), .A1(\depth_n.r_data[1][61] ), .Z(n45));
Q_MX02 U47 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][60] ), .A1(\depth_n.r_data[1][60] ), .Z(n46));
Q_MX02 U48 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][59] ), .A1(\depth_n.r_data[1][59] ), .Z(n47));
Q_MX02 U49 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][58] ), .A1(\depth_n.r_data[1][58] ), .Z(n48));
Q_MX02 U50 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][57] ), .A1(\depth_n.r_data[1][57] ), .Z(n49));
Q_MX02 U51 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][56] ), .A1(\depth_n.r_data[1][56] ), .Z(n50));
Q_MX02 U52 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][55] ), .A1(\depth_n.r_data[1][55] ), .Z(n51));
Q_MX02 U53 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][54] ), .A1(\depth_n.r_data[1][54] ), .Z(n52));
Q_MX02 U54 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][53] ), .A1(\depth_n.r_data[1][53] ), .Z(n53));
Q_MX02 U55 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][52] ), .A1(\depth_n.r_data[1][52] ), .Z(n54));
Q_MX02 U56 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][51] ), .A1(\depth_n.r_data[1][51] ), .Z(n55));
Q_MX02 U57 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][50] ), .A1(\depth_n.r_data[1][50] ), .Z(n56));
Q_MX02 U58 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][49] ), .A1(\depth_n.r_data[1][49] ), .Z(n57));
Q_MX02 U59 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][48] ), .A1(\depth_n.r_data[1][48] ), .Z(n58));
Q_MX02 U60 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][47] ), .A1(\depth_n.r_data[1][47] ), .Z(n59));
Q_MX02 U61 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][46] ), .A1(\depth_n.r_data[1][46] ), .Z(n60));
Q_MX02 U62 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][45] ), .A1(\depth_n.r_data[1][45] ), .Z(n61));
Q_MX02 U63 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][44] ), .A1(\depth_n.r_data[1][44] ), .Z(n62));
Q_MX02 U64 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][43] ), .A1(\depth_n.r_data[1][43] ), .Z(n63));
Q_MX02 U65 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][42] ), .A1(\depth_n.r_data[1][42] ), .Z(n64));
Q_MX02 U66 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][41] ), .A1(\depth_n.r_data[1][41] ), .Z(n65));
Q_MX02 U67 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][40] ), .A1(\depth_n.r_data[1][40] ), .Z(n66));
Q_MX02 U68 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][39] ), .A1(\depth_n.r_data[1][39] ), .Z(n67));
Q_MX02 U69 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][38] ), .A1(\depth_n.r_data[1][38] ), .Z(n68));
Q_MX02 U70 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][37] ), .A1(\depth_n.r_data[1][37] ), .Z(n69));
Q_MX02 U71 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][36] ), .A1(\depth_n.r_data[1][36] ), .Z(n70));
Q_MX02 U72 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][35] ), .A1(\depth_n.r_data[1][35] ), .Z(n71));
Q_MX02 U73 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][34] ), .A1(\depth_n.r_data[1][34] ), .Z(n72));
Q_MX02 U74 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][33] ), .A1(\depth_n.r_data[1][33] ), .Z(n73));
Q_MX02 U75 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][32] ), .A1(\depth_n.r_data[1][32] ), .Z(n74));
Q_MX02 U76 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][31] ), .A1(\depth_n.r_data[1][31] ), .Z(n75));
Q_MX02 U77 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][30] ), .A1(\depth_n.r_data[1][30] ), .Z(n76));
Q_MX02 U78 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][29] ), .A1(\depth_n.r_data[1][29] ), .Z(n77));
Q_MX02 U79 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][28] ), .A1(\depth_n.r_data[1][28] ), .Z(n78));
Q_MX02 U80 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][27] ), .A1(\depth_n.r_data[1][27] ), .Z(n79));
Q_MX02 U81 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][26] ), .A1(\depth_n.r_data[1][26] ), .Z(n80));
Q_MX02 U82 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][25] ), .A1(\depth_n.r_data[1][25] ), .Z(n81));
Q_MX02 U83 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][24] ), .A1(\depth_n.r_data[1][24] ), .Z(n82));
Q_MX02 U84 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][23] ), .A1(\depth_n.r_data[1][23] ), .Z(n83));
Q_MX02 U85 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][22] ), .A1(\depth_n.r_data[1][22] ), .Z(n84));
Q_MX02 U86 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][21] ), .A1(\depth_n.r_data[1][21] ), .Z(n85));
Q_MX02 U87 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][20] ), .A1(\depth_n.r_data[1][20] ), .Z(n86));
Q_MX02 U88 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][19] ), .A1(\depth_n.r_data[1][19] ), .Z(n87));
Q_MX02 U89 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][18] ), .A1(\depth_n.r_data[1][18] ), .Z(n88));
Q_MX02 U90 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][17] ), .A1(\depth_n.r_data[1][17] ), .Z(n89));
Q_MX02 U91 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][16] ), .A1(\depth_n.r_data[1][16] ), .Z(n90));
Q_MX02 U92 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][15] ), .A1(\depth_n.r_data[1][15] ), .Z(n91));
Q_MX02 U93 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][14] ), .A1(\depth_n.r_data[1][14] ), .Z(n92));
Q_MX02 U94 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][13] ), .A1(\depth_n.r_data[1][13] ), .Z(n93));
Q_MX02 U95 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][12] ), .A1(\depth_n.r_data[1][12] ), .Z(n94));
Q_MX02 U96 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][11] ), .A1(\depth_n.r_data[1][11] ), .Z(n95));
Q_MX02 U97 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][10] ), .A1(\depth_n.r_data[1][10] ), .Z(n96));
Q_MX02 U98 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][9] ), .A1(\depth_n.r_data[1][9] ), .Z(n97));
Q_MX02 U99 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][8] ), .A1(\depth_n.r_data[1][8] ), .Z(n98));
Q_MX02 U100 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][7] ), .A1(\depth_n.r_data[1][7] ), .Z(n99));
Q_MX02 U101 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][6] ), .A1(\depth_n.r_data[1][6] ), .Z(n100));
Q_MX02 U102 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][5] ), .A1(\depth_n.r_data[1][5] ), .Z(n101));
Q_MX02 U103 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][4] ), .A1(\depth_n.r_data[1][4] ), .Z(n102));
Q_MX02 U104 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][3] ), .A1(\depth_n.r_data[1][3] ), .Z(n103));
Q_MX02 U105 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][2] ), .A1(\depth_n.r_data[1][2] ), .Z(n104));
Q_MX02 U106 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][1] ), .A1(\depth_n.r_data[1][1] ), .Z(n105));
Q_MX02 U107 ( .S(\depth_n.rptr [0]), .A0(\depth_n.r_data[0][0] ), .A1(\depth_n.r_data[1][0] ), .Z(n106));
Q_AN02 U108 ( .A0(n108), .A1(n111), .Z(n107));
Q_INV U109 ( .A(n109), .Z(n108));
Q_AN02 U110 ( .A0(\depth_n.wptr [0]), .A1(n111), .Z(n109));
Q_INV U111 ( .A(empty), .Z(n110));
Q_AN02 U112 ( .A0(n110), .A1(n1), .Z(rdata[105]));
Q_AN02 U113 ( .A0(n110), .A1(n2), .Z(rdata[104]));
Q_AN02 U114 ( .A0(n110), .A1(n3), .Z(rdata[103]));
Q_AN02 U115 ( .A0(n110), .A1(n4), .Z(rdata[102]));
Q_AN02 U116 ( .A0(n110), .A1(n5), .Z(rdata[101]));
Q_AN02 U117 ( .A0(n110), .A1(n6), .Z(rdata[100]));
Q_AN02 U118 ( .A0(n110), .A1(n7), .Z(rdata[99]));
Q_AN02 U119 ( .A0(n110), .A1(n8), .Z(rdata[98]));
Q_AN02 U120 ( .A0(n110), .A1(n9), .Z(rdata[97]));
Q_AN02 U121 ( .A0(n110), .A1(n10), .Z(rdata[96]));
Q_AN02 U122 ( .A0(n110), .A1(n11), .Z(rdata[95]));
Q_AN02 U123 ( .A0(n110), .A1(n12), .Z(rdata[94]));
Q_AN02 U124 ( .A0(n110), .A1(n13), .Z(rdata[93]));
Q_AN02 U125 ( .A0(n110), .A1(n14), .Z(rdata[92]));
Q_AN02 U126 ( .A0(n110), .A1(n15), .Z(rdata[91]));
Q_AN02 U127 ( .A0(n110), .A1(n16), .Z(rdata[90]));
Q_AN02 U128 ( .A0(n110), .A1(n17), .Z(rdata[89]));
Q_AN02 U129 ( .A0(n110), .A1(n18), .Z(rdata[88]));
Q_AN02 U130 ( .A0(n110), .A1(n19), .Z(rdata[87]));
Q_AN02 U131 ( .A0(n110), .A1(n20), .Z(rdata[86]));
Q_AN02 U132 ( .A0(n110), .A1(n21), .Z(rdata[85]));
Q_AN02 U133 ( .A0(n110), .A1(n22), .Z(rdata[84]));
Q_AN02 U134 ( .A0(n110), .A1(n23), .Z(rdata[83]));
Q_AN02 U135 ( .A0(n110), .A1(n24), .Z(rdata[82]));
Q_AN02 U136 ( .A0(n110), .A1(n25), .Z(rdata[81]));
Q_AN02 U137 ( .A0(n110), .A1(n26), .Z(rdata[80]));
Q_AN02 U138 ( .A0(n110), .A1(n27), .Z(rdata[79]));
Q_AN02 U139 ( .A0(n110), .A1(n28), .Z(rdata[78]));
Q_AN02 U140 ( .A0(n110), .A1(n29), .Z(rdata[77]));
Q_AN02 U141 ( .A0(n110), .A1(n30), .Z(rdata[76]));
Q_AN02 U142 ( .A0(n110), .A1(n31), .Z(rdata[75]));
Q_AN02 U143 ( .A0(n110), .A1(n32), .Z(rdata[74]));
Q_AN02 U144 ( .A0(n110), .A1(n33), .Z(rdata[73]));
Q_AN02 U145 ( .A0(n110), .A1(n34), .Z(rdata[72]));
Q_AN02 U146 ( .A0(n110), .A1(n35), .Z(rdata[71]));
Q_AN02 U147 ( .A0(n110), .A1(n36), .Z(rdata[70]));
Q_AN02 U148 ( .A0(n110), .A1(n37), .Z(rdata[69]));
Q_AN02 U149 ( .A0(n110), .A1(n38), .Z(rdata[68]));
Q_AN02 U150 ( .A0(n110), .A1(n39), .Z(rdata[67]));
Q_AN02 U151 ( .A0(n110), .A1(n40), .Z(rdata[66]));
Q_AN02 U152 ( .A0(n110), .A1(n41), .Z(rdata[65]));
Q_AN02 U153 ( .A0(n110), .A1(n42), .Z(rdata[64]));
Q_AN02 U154 ( .A0(n110), .A1(n43), .Z(rdata[63]));
Q_AN02 U155 ( .A0(n110), .A1(n44), .Z(rdata[62]));
Q_AN02 U156 ( .A0(n110), .A1(n45), .Z(rdata[61]));
Q_AN02 U157 ( .A0(n110), .A1(n46), .Z(rdata[60]));
Q_AN02 U158 ( .A0(n110), .A1(n47), .Z(rdata[59]));
Q_AN02 U159 ( .A0(n110), .A1(n48), .Z(rdata[58]));
Q_AN02 U160 ( .A0(n110), .A1(n49), .Z(rdata[57]));
Q_AN02 U161 ( .A0(n110), .A1(n50), .Z(rdata[56]));
Q_AN02 U162 ( .A0(n110), .A1(n51), .Z(rdata[55]));
Q_AN02 U163 ( .A0(n110), .A1(n52), .Z(rdata[54]));
Q_AN02 U164 ( .A0(n110), .A1(n53), .Z(rdata[53]));
Q_AN02 U165 ( .A0(n110), .A1(n54), .Z(rdata[52]));
Q_AN02 U166 ( .A0(n110), .A1(n55), .Z(rdata[51]));
Q_AN02 U167 ( .A0(n110), .A1(n56), .Z(rdata[50]));
Q_AN02 U168 ( .A0(n110), .A1(n57), .Z(rdata[49]));
Q_AN02 U169 ( .A0(n110), .A1(n58), .Z(rdata[48]));
Q_AN02 U170 ( .A0(n110), .A1(n59), .Z(rdata[47]));
Q_AN02 U171 ( .A0(n110), .A1(n60), .Z(rdata[46]));
Q_AN02 U172 ( .A0(n110), .A1(n61), .Z(rdata[45]));
Q_AN02 U173 ( .A0(n110), .A1(n62), .Z(rdata[44]));
Q_AN02 U174 ( .A0(n110), .A1(n63), .Z(rdata[43]));
Q_AN02 U175 ( .A0(n110), .A1(n64), .Z(rdata[42]));
Q_AN02 U176 ( .A0(n110), .A1(n65), .Z(rdata[41]));
Q_AN02 U177 ( .A0(n110), .A1(n66), .Z(rdata[40]));
Q_AN02 U178 ( .A0(n110), .A1(n67), .Z(rdata[39]));
Q_AN02 U179 ( .A0(n110), .A1(n68), .Z(rdata[38]));
Q_AN02 U180 ( .A0(n110), .A1(n69), .Z(rdata[37]));
Q_AN02 U181 ( .A0(n110), .A1(n70), .Z(rdata[36]));
Q_AN02 U182 ( .A0(n110), .A1(n71), .Z(rdata[35]));
Q_AN02 U183 ( .A0(n110), .A1(n72), .Z(rdata[34]));
Q_AN02 U184 ( .A0(n110), .A1(n73), .Z(rdata[33]));
Q_AN02 U185 ( .A0(n110), .A1(n74), .Z(rdata[32]));
Q_AN02 U186 ( .A0(n110), .A1(n75), .Z(rdata[31]));
Q_AN02 U187 ( .A0(n110), .A1(n76), .Z(rdata[30]));
Q_AN02 U188 ( .A0(n110), .A1(n77), .Z(rdata[29]));
Q_AN02 U189 ( .A0(n110), .A1(n78), .Z(rdata[28]));
Q_AN02 U190 ( .A0(n110), .A1(n79), .Z(rdata[27]));
Q_AN02 U191 ( .A0(n110), .A1(n80), .Z(rdata[26]));
Q_AN02 U192 ( .A0(n110), .A1(n81), .Z(rdata[25]));
Q_AN02 U193 ( .A0(n110), .A1(n82), .Z(rdata[24]));
Q_AN02 U194 ( .A0(n110), .A1(n83), .Z(rdata[23]));
Q_AN02 U195 ( .A0(n110), .A1(n84), .Z(rdata[22]));
Q_AN02 U196 ( .A0(n110), .A1(n85), .Z(rdata[21]));
Q_AN02 U197 ( .A0(n110), .A1(n86), .Z(rdata[20]));
Q_AN02 U198 ( .A0(n110), .A1(n87), .Z(rdata[19]));
Q_AN02 U199 ( .A0(n110), .A1(n88), .Z(rdata[18]));
Q_AN02 U200 ( .A0(n110), .A1(n89), .Z(rdata[17]));
Q_AN02 U201 ( .A0(n110), .A1(n90), .Z(rdata[16]));
Q_AN02 U202 ( .A0(n110), .A1(n91), .Z(rdata[15]));
Q_AN02 U203 ( .A0(n110), .A1(n92), .Z(rdata[14]));
Q_AN02 U204 ( .A0(n110), .A1(n93), .Z(rdata[13]));
Q_AN02 U205 ( .A0(n110), .A1(n94), .Z(rdata[12]));
Q_AN02 U206 ( .A0(n110), .A1(n95), .Z(rdata[11]));
Q_AN02 U207 ( .A0(n110), .A1(n96), .Z(rdata[10]));
Q_AN02 U208 ( .A0(n110), .A1(n97), .Z(rdata[9]));
Q_AN02 U209 ( .A0(n110), .A1(n98), .Z(rdata[8]));
Q_AN02 U210 ( .A0(n110), .A1(n99), .Z(rdata[7]));
Q_AN02 U211 ( .A0(n110), .A1(n100), .Z(rdata[6]));
Q_AN02 U212 ( .A0(n110), .A1(n101), .Z(rdata[5]));
Q_AN02 U213 ( .A0(n110), .A1(n102), .Z(rdata[4]));
Q_AN02 U214 ( .A0(n110), .A1(n103), .Z(rdata[3]));
Q_AN02 U215 ( .A0(n110), .A1(n104), .Z(rdata[2]));
Q_AN02 U216 ( .A0(n110), .A1(n105), .Z(rdata[1]));
Q_AN02 U217 ( .A0(n110), .A1(n106), .Z(rdata[0]));
Q_INV U218 ( .A(full), .Z(n112));
Q_AN02 U219 ( .A0(wen), .A1(n112), .Z(n111));
nx_fifo_ctrl_xcm39 \depth_n.fifo_ctrl ( .empty( empty), .full( full), 
	.used_slots( used_slots[1:0]), .free_slots( free_slots[1:0]), 
	.rptr( \depth_n.rptr [0]), .wptr( \depth_n.wptr [0]), .underflow( 
	\depth_n._zy_simnet_underflow_2_w$ ), .overflow( 
	\depth_n._zy_simnet_overflow_3_w$ ), .clk( clk), .rst_n( rst_n), 
	.wen( wen), .ren( ren), .clear( clear));
ixc_assign \depth_n._zz_strnp_1 ( overflow, 
	\depth_n._zy_simnet_overflow_3_w$ );
ixc_assign \depth_n._zz_strnp_0 ( underflow, 
	\depth_n._zy_simnet_underflow_2_w$ );
Q_FDP4EP \depth_n.r_data_REG[0][0] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[0]), .Q(\depth_n.r_data[0][0] ));
Q_FDP4EP \depth_n.r_data_REG[0][1] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[1]), .Q(\depth_n.r_data[0][1] ));
Q_FDP4EP \depth_n.r_data_REG[0][2] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[2]), .Q(\depth_n.r_data[0][2] ));
Q_FDP4EP \depth_n.r_data_REG[0][3] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[3]), .Q(\depth_n.r_data[0][3] ));
Q_FDP4EP \depth_n.r_data_REG[0][4] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[4]), .Q(\depth_n.r_data[0][4] ));
Q_FDP4EP \depth_n.r_data_REG[0][5] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[5]), .Q(\depth_n.r_data[0][5] ));
Q_FDP4EP \depth_n.r_data_REG[0][6] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[6]), .Q(\depth_n.r_data[0][6] ));
Q_FDP4EP \depth_n.r_data_REG[0][7] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[7]), .Q(\depth_n.r_data[0][7] ));
Q_FDP4EP \depth_n.r_data_REG[0][8] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[8]), .Q(\depth_n.r_data[0][8] ));
Q_FDP4EP \depth_n.r_data_REG[0][9] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[9]), .Q(\depth_n.r_data[0][9] ));
Q_FDP4EP \depth_n.r_data_REG[0][10] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[10]), .Q(\depth_n.r_data[0][10] ));
Q_FDP4EP \depth_n.r_data_REG[0][11] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[11]), .Q(\depth_n.r_data[0][11] ));
Q_FDP4EP \depth_n.r_data_REG[0][12] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[12]), .Q(\depth_n.r_data[0][12] ));
Q_FDP4EP \depth_n.r_data_REG[0][13] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[13]), .Q(\depth_n.r_data[0][13] ));
Q_FDP4EP \depth_n.r_data_REG[0][14] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[14]), .Q(\depth_n.r_data[0][14] ));
Q_FDP4EP \depth_n.r_data_REG[0][15] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[15]), .Q(\depth_n.r_data[0][15] ));
Q_FDP4EP \depth_n.r_data_REG[0][16] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[16]), .Q(\depth_n.r_data[0][16] ));
Q_FDP4EP \depth_n.r_data_REG[0][17] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[17]), .Q(\depth_n.r_data[0][17] ));
Q_FDP4EP \depth_n.r_data_REG[0][18] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[18]), .Q(\depth_n.r_data[0][18] ));
Q_FDP4EP \depth_n.r_data_REG[0][19] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[19]), .Q(\depth_n.r_data[0][19] ));
Q_FDP4EP \depth_n.r_data_REG[0][20] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[20]), .Q(\depth_n.r_data[0][20] ));
Q_FDP4EP \depth_n.r_data_REG[0][21] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[21]), .Q(\depth_n.r_data[0][21] ));
Q_FDP4EP \depth_n.r_data_REG[0][22] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[22]), .Q(\depth_n.r_data[0][22] ));
Q_FDP4EP \depth_n.r_data_REG[0][23] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[23]), .Q(\depth_n.r_data[0][23] ));
Q_FDP4EP \depth_n.r_data_REG[0][24] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[24]), .Q(\depth_n.r_data[0][24] ));
Q_FDP4EP \depth_n.r_data_REG[0][25] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[25]), .Q(\depth_n.r_data[0][25] ));
Q_FDP4EP \depth_n.r_data_REG[0][26] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[26]), .Q(\depth_n.r_data[0][26] ));
Q_FDP4EP \depth_n.r_data_REG[0][27] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[27]), .Q(\depth_n.r_data[0][27] ));
Q_FDP4EP \depth_n.r_data_REG[0][28] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[28]), .Q(\depth_n.r_data[0][28] ));
Q_FDP4EP \depth_n.r_data_REG[0][29] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[29]), .Q(\depth_n.r_data[0][29] ));
Q_FDP4EP \depth_n.r_data_REG[0][30] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[30]), .Q(\depth_n.r_data[0][30] ));
Q_FDP4EP \depth_n.r_data_REG[0][31] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[31]), .Q(\depth_n.r_data[0][31] ));
Q_FDP4EP \depth_n.r_data_REG[0][32] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[32]), .Q(\depth_n.r_data[0][32] ));
Q_FDP4EP \depth_n.r_data_REG[0][33] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[33]), .Q(\depth_n.r_data[0][33] ));
Q_FDP4EP \depth_n.r_data_REG[0][34] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[34]), .Q(\depth_n.r_data[0][34] ));
Q_FDP4EP \depth_n.r_data_REG[0][35] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[35]), .Q(\depth_n.r_data[0][35] ));
Q_FDP4EP \depth_n.r_data_REG[0][36] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[36]), .Q(\depth_n.r_data[0][36] ));
Q_FDP4EP \depth_n.r_data_REG[0][37] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[37]), .Q(\depth_n.r_data[0][37] ));
Q_FDP4EP \depth_n.r_data_REG[0][38] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[38]), .Q(\depth_n.r_data[0][38] ));
Q_FDP4EP \depth_n.r_data_REG[0][39] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[39]), .Q(\depth_n.r_data[0][39] ));
Q_FDP4EP \depth_n.r_data_REG[0][40] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[40]), .Q(\depth_n.r_data[0][40] ));
Q_FDP4EP \depth_n.r_data_REG[0][41] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[41]), .Q(\depth_n.r_data[0][41] ));
Q_FDP4EP \depth_n.r_data_REG[0][42] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[42]), .Q(\depth_n.r_data[0][42] ));
Q_FDP4EP \depth_n.r_data_REG[0][43] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[43]), .Q(\depth_n.r_data[0][43] ));
Q_FDP4EP \depth_n.r_data_REG[0][44] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[44]), .Q(\depth_n.r_data[0][44] ));
Q_FDP4EP \depth_n.r_data_REG[0][45] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[45]), .Q(\depth_n.r_data[0][45] ));
Q_FDP4EP \depth_n.r_data_REG[0][46] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[46]), .Q(\depth_n.r_data[0][46] ));
Q_FDP4EP \depth_n.r_data_REG[0][47] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[47]), .Q(\depth_n.r_data[0][47] ));
Q_FDP4EP \depth_n.r_data_REG[0][48] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[48]), .Q(\depth_n.r_data[0][48] ));
Q_FDP4EP \depth_n.r_data_REG[0][49] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[49]), .Q(\depth_n.r_data[0][49] ));
Q_FDP4EP \depth_n.r_data_REG[0][50] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[50]), .Q(\depth_n.r_data[0][50] ));
Q_FDP4EP \depth_n.r_data_REG[0][51] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[51]), .Q(\depth_n.r_data[0][51] ));
Q_FDP4EP \depth_n.r_data_REG[0][52] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[52]), .Q(\depth_n.r_data[0][52] ));
Q_FDP4EP \depth_n.r_data_REG[0][53] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[53]), .Q(\depth_n.r_data[0][53] ));
Q_FDP4EP \depth_n.r_data_REG[0][54] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[54]), .Q(\depth_n.r_data[0][54] ));
Q_FDP4EP \depth_n.r_data_REG[0][55] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[55]), .Q(\depth_n.r_data[0][55] ));
Q_FDP4EP \depth_n.r_data_REG[0][56] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[56]), .Q(\depth_n.r_data[0][56] ));
Q_FDP4EP \depth_n.r_data_REG[0][57] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[57]), .Q(\depth_n.r_data[0][57] ));
Q_FDP4EP \depth_n.r_data_REG[0][58] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[58]), .Q(\depth_n.r_data[0][58] ));
Q_FDP4EP \depth_n.r_data_REG[0][59] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[59]), .Q(\depth_n.r_data[0][59] ));
Q_FDP4EP \depth_n.r_data_REG[0][60] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[60]), .Q(\depth_n.r_data[0][60] ));
Q_FDP4EP \depth_n.r_data_REG[0][61] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[61]), .Q(\depth_n.r_data[0][61] ));
Q_FDP4EP \depth_n.r_data_REG[0][62] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[62]), .Q(\depth_n.r_data[0][62] ));
Q_FDP4EP \depth_n.r_data_REG[0][63] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[63]), .Q(\depth_n.r_data[0][63] ));
Q_FDP4EP \depth_n.r_data_REG[0][64] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[64]), .Q(\depth_n.r_data[0][64] ));
Q_FDP4EP \depth_n.r_data_REG[0][65] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[65]), .Q(\depth_n.r_data[0][65] ));
Q_FDP4EP \depth_n.r_data_REG[0][66] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[66]), .Q(\depth_n.r_data[0][66] ));
Q_FDP4EP \depth_n.r_data_REG[0][67] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[67]), .Q(\depth_n.r_data[0][67] ));
Q_FDP4EP \depth_n.r_data_REG[0][68] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[68]), .Q(\depth_n.r_data[0][68] ));
Q_FDP4EP \depth_n.r_data_REG[0][69] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[69]), .Q(\depth_n.r_data[0][69] ));
Q_FDP4EP \depth_n.r_data_REG[0][70] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[70]), .Q(\depth_n.r_data[0][70] ));
Q_FDP4EP \depth_n.r_data_REG[0][71] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[71]), .Q(\depth_n.r_data[0][71] ));
Q_FDP4EP \depth_n.r_data_REG[0][72] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[72]), .Q(\depth_n.r_data[0][72] ));
Q_FDP4EP \depth_n.r_data_REG[0][73] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[73]), .Q(\depth_n.r_data[0][73] ));
Q_FDP4EP \depth_n.r_data_REG[0][74] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[74]), .Q(\depth_n.r_data[0][74] ));
Q_FDP4EP \depth_n.r_data_REG[0][75] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[75]), .Q(\depth_n.r_data[0][75] ));
Q_FDP4EP \depth_n.r_data_REG[0][76] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[76]), .Q(\depth_n.r_data[0][76] ));
Q_FDP4EP \depth_n.r_data_REG[0][77] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[77]), .Q(\depth_n.r_data[0][77] ));
Q_FDP4EP \depth_n.r_data_REG[0][78] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[78]), .Q(\depth_n.r_data[0][78] ));
Q_FDP4EP \depth_n.r_data_REG[0][79] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[79]), .Q(\depth_n.r_data[0][79] ));
Q_FDP4EP \depth_n.r_data_REG[0][80] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[80]), .Q(\depth_n.r_data[0][80] ));
Q_FDP4EP \depth_n.r_data_REG[0][81] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[81]), .Q(\depth_n.r_data[0][81] ));
Q_FDP4EP \depth_n.r_data_REG[0][82] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[82]), .Q(\depth_n.r_data[0][82] ));
Q_FDP4EP \depth_n.r_data_REG[0][83] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[83]), .Q(\depth_n.r_data[0][83] ));
Q_FDP4EP \depth_n.r_data_REG[0][84] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[84]), .Q(\depth_n.r_data[0][84] ));
Q_FDP4EP \depth_n.r_data_REG[0][85] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[85]), .Q(\depth_n.r_data[0][85] ));
Q_FDP4EP \depth_n.r_data_REG[0][86] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[86]), .Q(\depth_n.r_data[0][86] ));
Q_FDP4EP \depth_n.r_data_REG[0][87] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[87]), .Q(\depth_n.r_data[0][87] ));
Q_FDP4EP \depth_n.r_data_REG[0][88] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[88]), .Q(\depth_n.r_data[0][88] ));
Q_FDP4EP \depth_n.r_data_REG[0][89] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[89]), .Q(\depth_n.r_data[0][89] ));
Q_FDP4EP \depth_n.r_data_REG[0][90] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[90]), .Q(\depth_n.r_data[0][90] ));
Q_FDP4EP \depth_n.r_data_REG[0][91] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[91]), .Q(\depth_n.r_data[0][91] ));
Q_FDP4EP \depth_n.r_data_REG[0][92] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[92]), .Q(\depth_n.r_data[0][92] ));
Q_FDP4EP \depth_n.r_data_REG[0][93] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[93]), .Q(\depth_n.r_data[0][93] ));
Q_FDP4EP \depth_n.r_data_REG[0][94] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[94]), .Q(\depth_n.r_data[0][94] ));
Q_FDP4EP \depth_n.r_data_REG[0][95] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[95]), .Q(\depth_n.r_data[0][95] ));
Q_FDP4EP \depth_n.r_data_REG[0][96] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[96]), .Q(\depth_n.r_data[0][96] ));
Q_FDP4EP \depth_n.r_data_REG[0][97] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[97]), .Q(\depth_n.r_data[0][97] ));
Q_FDP4EP \depth_n.r_data_REG[0][98] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[98]), .Q(\depth_n.r_data[0][98] ));
Q_FDP4EP \depth_n.r_data_REG[0][99] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[99]), .Q(\depth_n.r_data[0][99] ));
Q_FDP4EP \depth_n.r_data_REG[0][100] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[100]), .Q(\depth_n.r_data[0][100] ));
Q_FDP4EP \depth_n.r_data_REG[0][101] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[101]), .Q(\depth_n.r_data[0][101] ));
Q_FDP4EP \depth_n.r_data_REG[0][102] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[102]), .Q(\depth_n.r_data[0][102] ));
Q_FDP4EP \depth_n.r_data_REG[0][103] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[103]), .Q(\depth_n.r_data[0][103] ));
Q_FDP4EP \depth_n.r_data_REG[0][104] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[104]), .Q(\depth_n.r_data[0][104] ));
Q_FDP4EP \depth_n.r_data_REG[0][105] ( .CK(clk), .CE(n107), .R(n113), .D(wdata[105]), .Q(\depth_n.r_data[0][105] ));
Q_FDP4EP \depth_n.r_data_REG[1][0] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[0]), .Q(\depth_n.r_data[1][0] ));
Q_FDP4EP \depth_n.r_data_REG[1][1] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[1]), .Q(\depth_n.r_data[1][1] ));
Q_FDP4EP \depth_n.r_data_REG[1][2] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[2]), .Q(\depth_n.r_data[1][2] ));
Q_FDP4EP \depth_n.r_data_REG[1][3] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[3]), .Q(\depth_n.r_data[1][3] ));
Q_FDP4EP \depth_n.r_data_REG[1][4] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[4]), .Q(\depth_n.r_data[1][4] ));
Q_FDP4EP \depth_n.r_data_REG[1][5] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[5]), .Q(\depth_n.r_data[1][5] ));
Q_FDP4EP \depth_n.r_data_REG[1][6] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[6]), .Q(\depth_n.r_data[1][6] ));
Q_FDP4EP \depth_n.r_data_REG[1][7] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[7]), .Q(\depth_n.r_data[1][7] ));
Q_FDP4EP \depth_n.r_data_REG[1][8] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[8]), .Q(\depth_n.r_data[1][8] ));
Q_FDP4EP \depth_n.r_data_REG[1][9] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[9]), .Q(\depth_n.r_data[1][9] ));
Q_FDP4EP \depth_n.r_data_REG[1][10] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[10]), .Q(\depth_n.r_data[1][10] ));
Q_FDP4EP \depth_n.r_data_REG[1][11] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[11]), .Q(\depth_n.r_data[1][11] ));
Q_FDP4EP \depth_n.r_data_REG[1][12] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[12]), .Q(\depth_n.r_data[1][12] ));
Q_FDP4EP \depth_n.r_data_REG[1][13] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[13]), .Q(\depth_n.r_data[1][13] ));
Q_FDP4EP \depth_n.r_data_REG[1][14] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[14]), .Q(\depth_n.r_data[1][14] ));
Q_FDP4EP \depth_n.r_data_REG[1][15] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[15]), .Q(\depth_n.r_data[1][15] ));
Q_FDP4EP \depth_n.r_data_REG[1][16] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[16]), .Q(\depth_n.r_data[1][16] ));
Q_FDP4EP \depth_n.r_data_REG[1][17] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[17]), .Q(\depth_n.r_data[1][17] ));
Q_FDP4EP \depth_n.r_data_REG[1][18] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[18]), .Q(\depth_n.r_data[1][18] ));
Q_FDP4EP \depth_n.r_data_REG[1][19] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[19]), .Q(\depth_n.r_data[1][19] ));
Q_FDP4EP \depth_n.r_data_REG[1][20] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[20]), .Q(\depth_n.r_data[1][20] ));
Q_FDP4EP \depth_n.r_data_REG[1][21] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[21]), .Q(\depth_n.r_data[1][21] ));
Q_FDP4EP \depth_n.r_data_REG[1][22] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[22]), .Q(\depth_n.r_data[1][22] ));
Q_FDP4EP \depth_n.r_data_REG[1][23] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[23]), .Q(\depth_n.r_data[1][23] ));
Q_FDP4EP \depth_n.r_data_REG[1][24] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[24]), .Q(\depth_n.r_data[1][24] ));
Q_FDP4EP \depth_n.r_data_REG[1][25] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[25]), .Q(\depth_n.r_data[1][25] ));
Q_FDP4EP \depth_n.r_data_REG[1][26] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[26]), .Q(\depth_n.r_data[1][26] ));
Q_FDP4EP \depth_n.r_data_REG[1][27] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[27]), .Q(\depth_n.r_data[1][27] ));
Q_FDP4EP \depth_n.r_data_REG[1][28] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[28]), .Q(\depth_n.r_data[1][28] ));
Q_FDP4EP \depth_n.r_data_REG[1][29] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[29]), .Q(\depth_n.r_data[1][29] ));
Q_FDP4EP \depth_n.r_data_REG[1][30] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[30]), .Q(\depth_n.r_data[1][30] ));
Q_FDP4EP \depth_n.r_data_REG[1][31] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[31]), .Q(\depth_n.r_data[1][31] ));
Q_FDP4EP \depth_n.r_data_REG[1][32] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[32]), .Q(\depth_n.r_data[1][32] ));
Q_FDP4EP \depth_n.r_data_REG[1][33] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[33]), .Q(\depth_n.r_data[1][33] ));
Q_FDP4EP \depth_n.r_data_REG[1][34] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[34]), .Q(\depth_n.r_data[1][34] ));
Q_FDP4EP \depth_n.r_data_REG[1][35] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[35]), .Q(\depth_n.r_data[1][35] ));
Q_FDP4EP \depth_n.r_data_REG[1][36] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[36]), .Q(\depth_n.r_data[1][36] ));
Q_FDP4EP \depth_n.r_data_REG[1][37] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[37]), .Q(\depth_n.r_data[1][37] ));
Q_FDP4EP \depth_n.r_data_REG[1][38] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[38]), .Q(\depth_n.r_data[1][38] ));
Q_FDP4EP \depth_n.r_data_REG[1][39] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[39]), .Q(\depth_n.r_data[1][39] ));
Q_FDP4EP \depth_n.r_data_REG[1][40] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[40]), .Q(\depth_n.r_data[1][40] ));
Q_FDP4EP \depth_n.r_data_REG[1][41] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[41]), .Q(\depth_n.r_data[1][41] ));
Q_FDP4EP \depth_n.r_data_REG[1][42] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[42]), .Q(\depth_n.r_data[1][42] ));
Q_FDP4EP \depth_n.r_data_REG[1][43] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[43]), .Q(\depth_n.r_data[1][43] ));
Q_FDP4EP \depth_n.r_data_REG[1][44] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[44]), .Q(\depth_n.r_data[1][44] ));
Q_FDP4EP \depth_n.r_data_REG[1][45] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[45]), .Q(\depth_n.r_data[1][45] ));
Q_FDP4EP \depth_n.r_data_REG[1][46] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[46]), .Q(\depth_n.r_data[1][46] ));
Q_FDP4EP \depth_n.r_data_REG[1][47] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[47]), .Q(\depth_n.r_data[1][47] ));
Q_FDP4EP \depth_n.r_data_REG[1][48] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[48]), .Q(\depth_n.r_data[1][48] ));
Q_FDP4EP \depth_n.r_data_REG[1][49] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[49]), .Q(\depth_n.r_data[1][49] ));
Q_FDP4EP \depth_n.r_data_REG[1][50] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[50]), .Q(\depth_n.r_data[1][50] ));
Q_FDP4EP \depth_n.r_data_REG[1][51] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[51]), .Q(\depth_n.r_data[1][51] ));
Q_FDP4EP \depth_n.r_data_REG[1][52] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[52]), .Q(\depth_n.r_data[1][52] ));
Q_FDP4EP \depth_n.r_data_REG[1][53] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[53]), .Q(\depth_n.r_data[1][53] ));
Q_FDP4EP \depth_n.r_data_REG[1][54] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[54]), .Q(\depth_n.r_data[1][54] ));
Q_FDP4EP \depth_n.r_data_REG[1][55] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[55]), .Q(\depth_n.r_data[1][55] ));
Q_FDP4EP \depth_n.r_data_REG[1][56] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[56]), .Q(\depth_n.r_data[1][56] ));
Q_FDP4EP \depth_n.r_data_REG[1][57] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[57]), .Q(\depth_n.r_data[1][57] ));
Q_FDP4EP \depth_n.r_data_REG[1][58] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[58]), .Q(\depth_n.r_data[1][58] ));
Q_FDP4EP \depth_n.r_data_REG[1][59] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[59]), .Q(\depth_n.r_data[1][59] ));
Q_FDP4EP \depth_n.r_data_REG[1][60] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[60]), .Q(\depth_n.r_data[1][60] ));
Q_FDP4EP \depth_n.r_data_REG[1][61] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[61]), .Q(\depth_n.r_data[1][61] ));
Q_FDP4EP \depth_n.r_data_REG[1][62] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[62]), .Q(\depth_n.r_data[1][62] ));
Q_FDP4EP \depth_n.r_data_REG[1][63] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[63]), .Q(\depth_n.r_data[1][63] ));
Q_FDP4EP \depth_n.r_data_REG[1][64] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[64]), .Q(\depth_n.r_data[1][64] ));
Q_FDP4EP \depth_n.r_data_REG[1][65] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[65]), .Q(\depth_n.r_data[1][65] ));
Q_FDP4EP \depth_n.r_data_REG[1][66] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[66]), .Q(\depth_n.r_data[1][66] ));
Q_FDP4EP \depth_n.r_data_REG[1][67] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[67]), .Q(\depth_n.r_data[1][67] ));
Q_FDP4EP \depth_n.r_data_REG[1][68] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[68]), .Q(\depth_n.r_data[1][68] ));
Q_FDP4EP \depth_n.r_data_REG[1][69] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[69]), .Q(\depth_n.r_data[1][69] ));
Q_FDP4EP \depth_n.r_data_REG[1][70] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[70]), .Q(\depth_n.r_data[1][70] ));
Q_FDP4EP \depth_n.r_data_REG[1][71] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[71]), .Q(\depth_n.r_data[1][71] ));
Q_FDP4EP \depth_n.r_data_REG[1][72] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[72]), .Q(\depth_n.r_data[1][72] ));
Q_FDP4EP \depth_n.r_data_REG[1][73] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[73]), .Q(\depth_n.r_data[1][73] ));
Q_FDP4EP \depth_n.r_data_REG[1][74] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[74]), .Q(\depth_n.r_data[1][74] ));
Q_FDP4EP \depth_n.r_data_REG[1][75] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[75]), .Q(\depth_n.r_data[1][75] ));
Q_FDP4EP \depth_n.r_data_REG[1][76] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[76]), .Q(\depth_n.r_data[1][76] ));
Q_FDP4EP \depth_n.r_data_REG[1][77] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[77]), .Q(\depth_n.r_data[1][77] ));
Q_FDP4EP \depth_n.r_data_REG[1][78] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[78]), .Q(\depth_n.r_data[1][78] ));
Q_FDP4EP \depth_n.r_data_REG[1][79] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[79]), .Q(\depth_n.r_data[1][79] ));
Q_FDP4EP \depth_n.r_data_REG[1][80] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[80]), .Q(\depth_n.r_data[1][80] ));
Q_FDP4EP \depth_n.r_data_REG[1][81] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[81]), .Q(\depth_n.r_data[1][81] ));
Q_FDP4EP \depth_n.r_data_REG[1][82] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[82]), .Q(\depth_n.r_data[1][82] ));
Q_FDP4EP \depth_n.r_data_REG[1][83] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[83]), .Q(\depth_n.r_data[1][83] ));
Q_FDP4EP \depth_n.r_data_REG[1][84] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[84]), .Q(\depth_n.r_data[1][84] ));
Q_FDP4EP \depth_n.r_data_REG[1][85] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[85]), .Q(\depth_n.r_data[1][85] ));
Q_FDP4EP \depth_n.r_data_REG[1][86] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[86]), .Q(\depth_n.r_data[1][86] ));
Q_FDP4EP \depth_n.r_data_REG[1][87] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[87]), .Q(\depth_n.r_data[1][87] ));
Q_FDP4EP \depth_n.r_data_REG[1][88] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[88]), .Q(\depth_n.r_data[1][88] ));
Q_FDP4EP \depth_n.r_data_REG[1][89] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[89]), .Q(\depth_n.r_data[1][89] ));
Q_FDP4EP \depth_n.r_data_REG[1][90] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[90]), .Q(\depth_n.r_data[1][90] ));
Q_FDP4EP \depth_n.r_data_REG[1][91] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[91]), .Q(\depth_n.r_data[1][91] ));
Q_FDP4EP \depth_n.r_data_REG[1][92] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[92]), .Q(\depth_n.r_data[1][92] ));
Q_FDP4EP \depth_n.r_data_REG[1][93] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[93]), .Q(\depth_n.r_data[1][93] ));
Q_FDP4EP \depth_n.r_data_REG[1][94] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[94]), .Q(\depth_n.r_data[1][94] ));
Q_FDP4EP \depth_n.r_data_REG[1][95] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[95]), .Q(\depth_n.r_data[1][95] ));
Q_FDP4EP \depth_n.r_data_REG[1][96] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[96]), .Q(\depth_n.r_data[1][96] ));
Q_FDP4EP \depth_n.r_data_REG[1][97] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[97]), .Q(\depth_n.r_data[1][97] ));
Q_FDP4EP \depth_n.r_data_REG[1][98] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[98]), .Q(\depth_n.r_data[1][98] ));
Q_FDP4EP \depth_n.r_data_REG[1][99] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[99]), .Q(\depth_n.r_data[1][99] ));
Q_FDP4EP \depth_n.r_data_REG[1][100] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[100]), .Q(\depth_n.r_data[1][100] ));
Q_FDP4EP \depth_n.r_data_REG[1][101] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[101]), .Q(\depth_n.r_data[1][101] ));
Q_FDP4EP \depth_n.r_data_REG[1][102] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[102]), .Q(\depth_n.r_data[1][102] ));
Q_FDP4EP \depth_n.r_data_REG[1][103] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[103]), .Q(\depth_n.r_data[1][103] ));
Q_FDP4EP \depth_n.r_data_REG[1][104] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[104]), .Q(\depth_n.r_data[1][104] ));
Q_FDP4EP \depth_n.r_data_REG[1][105] ( .CK(clk), .CE(n109), .R(n113), .D(wdata[105]), .Q(\depth_n.r_data[1][105] ));
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m1 "\depth_n.r_data  1 105 0 1 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_NON_CMM "1"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_1 "0 genblk1  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_0 "-1 depth_n  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "depth_n.genblk1"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "depth_n"
endmodule
