// xc_work/v/WORK/svPkg1n.sv
// /home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kmePKG.svp:14
package cr_kmePKG;
import cr_kme_regsPKG::* ;
endpackage

