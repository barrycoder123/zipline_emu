// xc_work/v/150.sv
// /home/ibarry/Project-Zipline-master/dv/KME/run/tb_top.sv:0
// NOTE: This file corresponds to a module in the Hardware/DUT partition.
`timescale 1ps/1ps
module _ixc_isc;
// external : tb_top.kme_tb_dut._zyixc_port_0_0_isf (resolved )  (var)  
// external : xcva_top.IXC_GFIFO.ISF.pvec (resolved )  (var)  
wire  [0:0] _zz_dummy_0 ;
// quickturn name_map   _zz_dummy_0   xcva_top.IXC_GFIFO.ISF.pvec
// external : tb_top.kme_tb_dut._zyixc_port_0_0_osf (resolved )  (var)  
// external : xcva_top.IXC_GFIFO.OSF.pvecEv (resolved )  (var)  
bit [0:0] _zz_dummy_1 ;
// quickturn name_map   _zz_dummy_1   xcva_top.IXC_GFIFO.OSF.pvecEv
// external : xcva_top.tb_top.kme_tb_dut.kme_dut.u_cr_kme_core.kme_is_core.txc_axi_intf.u_cr_fifo_wrap2.ram_fifo.u_nx_fifo_ram_1r1w.fifo_ctrl._zyixc_port_1_0_osf (resolved )  (var)  
// external : xcva_top.IXC_GFIFO.OSF1.pvecEv (resolved )  (var)  
bit [19:0] _zz_dummy_2 ;
// quickturn name_map   _zz_dummy_2   xcva_top.IXC_GFIFO.OSF1.pvecEv
// external : xcva_top.tb_top.kme_tb_dut.kme_dut.u_cr_kme_core.kme_is_core.cceip_encrypt_kop_fifo.ram_fifo.ram_fifo.u_nx_fifo_ram_1r1w.fifo_ctrl._zyixc_port_1_0_osf (resolved )  (var)  
// external : xcva_top.tb_top.kme_tb_dut.kme_dut.u_cr_kme_core.kme_is_core.cceip_validate_kop_fifo.ram_fifo.ram_fifo.u_nx_fifo_ram_1r1w.fifo_ctrl._zyixc_port_1_0_osf (resolved )  (var)  
// external : xcva_top.tb_top.kme_tb_dut.kme_dut.u_cr_kme_core.kme_is_core.cceip0_key_tlv_rsm.u_cr_tlvp2_rsm.u_cr_fifo_wrap2_tob.ram_fifo.u_nx_fifo_ram_1r1w.fifo_ctrl._zyixc_port_1_0_osf (resolved )  (var)  
// external : tb_top.kme_tb_dut.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cceip0.u_nx_credit_manager._zyixc_port_1_0_osf (resolved )  (var)  
// external : tb_top.kme_tb_dut.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cceip0.u_nx_credit_manager._zyixc_port_1_1_osf (resolved )  (var)  
// external : tb_top.kme_tb_dut.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cceip1.u_nx_credit_manager._zyixc_port_1_0_osf (resolved )  (var)  
// external : tb_top.kme_tb_dut.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cceip1.u_nx_credit_manager._zyixc_port_1_1_osf (resolved )  (var)  
// external : tb_top.kme_tb_dut.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cceip2.u_nx_credit_manager._zyixc_port_1_0_osf (resolved )  (var)  
// external : tb_top.kme_tb_dut.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cceip2.u_nx_credit_manager._zyixc_port_1_1_osf (resolved )  (var)  
// external : tb_top.kme_tb_dut.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cceip3.u_nx_credit_manager._zyixc_port_1_0_osf (resolved )  (var)  
// external : tb_top.kme_tb_dut.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cceip3.u_nx_credit_manager._zyixc_port_1_1_osf (resolved )  (var)  
// external : tb_top.kme_tb_dut.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cddip0.u_nx_credit_manager._zyixc_port_1_0_osf (resolved )  (var)  
// external : tb_top.kme_tb_dut.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cddip0.u_nx_credit_manager._zyixc_port_1_1_osf (resolved )  (var)  
// external : tb_top.kme_tb_dut.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cddip1.u_nx_credit_manager._zyixc_port_1_0_osf (resolved )  (var)  
// external : tb_top.kme_tb_dut.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cddip1.u_nx_credit_manager._zyixc_port_1_1_osf (resolved )  (var)  
// external : tb_top.kme_tb_dut.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cddip2.u_nx_credit_manager._zyixc_port_1_0_osf (resolved )  (var)  
// external : tb_top.kme_tb_dut.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cddip2.u_nx_credit_manager._zyixc_port_1_1_osf (resolved )  (var)  
// external : tb_top.kme_tb_dut.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cddip3.u_nx_credit_manager._zyixc_port_1_0_osf (resolved )  (var)  
// external : tb_top.kme_tb_dut.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cddip3.u_nx_credit_manager._zyixc_port_1_1_osf (resolved )  (var)  
wire  assertion_coverage_on;
reg assertion_global_off_s = 0;
// quickturn keep_net assertion_global_off_s
// quickturn external_ref assertion_global_off_s
reg assertion_global_on_s = 1;
// quickturn keep_net assertion_global_on_s
// quickturn external_ref assertion_global_on_s
reg assertion_global_off_sD = 0;
// quickturn keep_net assertion_global_off_sD
reg assertion_global_on_sD = 1;
// quickturn keep_net assertion_global_on_sD
reg assertion_global_off_ev;
reg assertion_global_on_ev;
// synopsys translate_off
wire  assertion_global_off_p;
// quickturn keep_net assertion_global_off_p
wire  assertion_global_on_p;
// quickturn keep_net assertion_global_on_p
reg assertion_global_deposit_on;
reg assertion_global_copy_t = 1;
reg _zy_svaTrigger;
reg _zy_svaKill;
reg _zy_svaOn;
// synopsys translate_on
wire  assertUCF;
int _zy_ixcg_mdh_L0_0;
int _zy_ixcg_mdh_L0_1;

reg xc_top_eventOn;
// quickturn name_map xc_top_eventOn xc_top.eventOn
wire fclk;
// quickturn fast_clock fclk

always@(posedge fclk)
  if (xc_top_eventOn) begin
    assertion_global_off_sD <= assertion_global_off_s;
    assertion_global_on_sD <= assertion_global_on_s;
  end

always @(*)
  assertion_global_on_ev = xc_top_eventOn & (assertion_global_on_s != assertion_global_on_sD);

always @(*)
  assertion_global_off_ev = xc_top_eventOn & (assertion_global_off_s != assertion_global_off_sD);

pulldown(assertion_global_on_p);
pulldown(assertion_global_off_p);

assign assertion_global_on_p = (assertion_global_on_ev & assertion_global_on_s & ~assertion_global_off_s) ? 1'b1: 1'bz;
assign assertion_global_off_p = (assertion_global_off_ev & assertion_global_off_s & ~assertion_global_on_s) ? 1'b1: 1'bz;

// pragma CVASTRPROP MODULE _ixc_isc PROP_IXCOM_MOD TRUE
endmodule

