library ieee, quickturn ;
use ieee.std_logic_1164.all ;
use quickturn.verilog.all ;
use work.cr_kme_regfilePKG.all ;
entity cr_kme_kop_tlv_inspector_xcm69 is
  generic (
    CCEIP_ENCRYPT_KOP : integer := 0;
    subtype gcm_op_e is std_logic_vector(2 downto 0) ;
    constant PT_CKV : gcm_op_e := std_logic_vector'("000") ;
    constant PT_KEY_BLOB : gcm_op_e := std_logic_vector'("001") ;
    constant DECRYPT_DEK256 : gcm_op_e := std_logic_vector'("010") ;
    constant DECRYPT_DEK512 : gcm_op_e := std_logic_vector'("011") ;
    constant DECRYPT_DAK : gcm_op_e := std_logic_vector'("100") ;
    constant DECRYPT_DEK256_COMB : gcm_op_e := std_logic_vector'("101") ;
    constant DECRYPT_DEK512_COMB : gcm_op_e := std_logic_vector'("110") ;
    constant DECRYPT_DAK_COMB : gcm_op_e := std_logic_vector'("111");
    type $_gcm_cmd_t is
    record
      key0 : std_logic_vector(255 downto 0) ;
      key1 : std_logic_vector(255 downto 0) ;
      iv : std_logic_vector(95 downto 0) ;
      op : gcm_op_e ;
    end record ;
    subtype gcm_cmd_t is $_gcm_cmd_t std_logic_vector(610 downto 0);
    type $_keyfilter_cmd_t is
    record
      combo_mode : std_logic_vector(0 downto 0) ;
    end record ;
    subtype keyfilter_cmd_t is $_keyfilter_cmd_t std_logic_vector(0 downto 0);
    type $_kdfstream_cmd_t is
    record
      combo_mode : std_logic_vector(0 downto 0) ;
      skip : std_logic_vector(0 downto 0) ;
      guid : std_logic_vector(255 downto 0) ;
      label_index : std_logic_vector(2 downto 0) ;
      num_iter : std_logic_vector(1 downto 0) ;
    end record ;
    subtype kdfstream_cmd_t is $_kdfstream_cmd_t std_logic_vector(262 downto 0);
    subtype aux_key_op_e is std_logic_vector(0 downto 0) ;
    constant NOOP : aux_key_op_e := "0" ;
    constant KDF : aux_key_op_e := "1";
    type $_kdf_cmd_t is
    record
      kdf_dek_iter : std_logic_vector(0 downto 0) ;
      combo_mode : std_logic_vector(0 downto 0) ;
      dek_key_op : aux_key_op_e ;
      dak_key_op : aux_key_op_e ;
    end record ;
    subtype kdf_cmd_t is $_kdf_cmd_t std_logic_vector(3 downto 0);
    type $_label_t is
    record
      guid_size : std_logic_vector(0 downto 0) ;
      label_size : std_logic_vector(5 downto 0) ;
      DUMMY1 : std_logic_vector(255 downto 0) ;
      delimiter_valid : std_logic_vector(0 downto 0) ;
      delimiter : std_logic_vector(7 downto 0) ;
    end record ;
    subtype label_t is $_label_t std_logic_vector(271 downto 0);
    type DUMMY2 is array(integer range <>) of label_t;
    subtype kme_internal_id is std_logic_vector(3 downto 0) ;
    constant KME_WORD0 : kme_internal_id := std_logic_vector'("0000") ;
    constant KME_DEBUG_KEYHDR : kme_internal_id := std_logic_vector'("0001") ;
    constant KME_IVTWEAK : kme_internal_id := std_logic_vector'("0010") ;
    constant KME_GUID : kme_internal_id := std_logic_vector'("0011") ;
    constant KME_KIM : kme_internal_id := std_logic_vector'("0100") ;
    constant KME_DEK_CKV0 : kme_internal_id := std_logic_vector'("0101") ;
    constant KME_DEK_CKV1 : kme_internal_id := std_logic_vector'("0110") ;
    constant KME_DAK_CKV : kme_internal_id := std_logic_vector'("0111") ;
    constant KME_EIV : kme_internal_id := std_logic_vector'("1000") ;
    constant KME_DEK0 : kme_internal_id := std_logic_vector'("1001") ;
    constant KME_DEK1 : kme_internal_id := std_logic_vector'("1010") ;
    constant KME_ETAG : kme_internal_id := std_logic_vector'("1011") ;
    constant KME_AIV : kme_internal_id := std_logic_vector'("1100") ;
    constant KME_DAK : kme_internal_id := std_logic_vector'("1101") ;
    constant KME_ATAG : kme_internal_id := std_logic_vector'("1110") ;
    constant KME_ERROR : kme_internal_id := std_logic_vector'("1111");
    type $_kme_internal_t is
    record
      sot : std_logic_vector(0 downto 0) ;
      eoi : std_logic_vector(0 downto 0) ;
      eot : std_logic_vector(0 downto 0) ;
      id : kme_internal_id ;
      tdata : std_logic_vector(63 downto 0) ;
    end record ;
    subtype kme_internal_t is $_kme_internal_t std_logic_vector(70 downto 0)
  ) ;
  port (
    kme_internal_out_ack : out std_logic ;
    gcm_cmd_in : out gcm_cmd_t ;
    gcm_cmd_in_valid : out std_logic ;
    gcm_tag_data_in : out std_logic_vector(95 downto 0) ;
    gcm_tag_data_in_valid : out std_logic ;
    inspector_upsizer_valid : out std_logic ;
    inspector_upsizer_eof : out std_logic ;
    inspector_upsizer_data : out std_logic_vector(63 downto 0) ;
    keyfilter_cmd_in : out keyfilter_cmd_t ;
    keyfilter_cmd_in_valid : out std_logic ;
    kdfstream_cmd_in : out kdfstream_cmd_t ;
    kdfstream_cmd_in_valid : out std_logic ;
    kdf_cmd_in : out kdf_cmd_t ;
    kdf_cmd_in_valid : out std_logic ;
    tlv_sb_data_in : out std_logic_vector(63 downto 0) ;
    tlv_sb_data_in_valid : out std_logic ;
    clk : in std_logic ;
    rst_n : in std_logic ;
    labels : in DUMMY2(7 downto 0) ;
    -- quickturn array_with_packed_dim labels 2 0
    kme_internal_out : in kme_internal_t ;
    kme_internal_out_valid : in std_logic ;
    gcm_cmd_in_stall : in std_logic ;
    gcm_tag_data_in_stall : in std_logic ;
    upsizer_inspector_stall : in std_logic ;
    keyfilter_cmd_in_stall : in std_logic ;
    kdfstream_cmd_in_stall : in std_logic ;
    kdf_cmd_in_stall : in std_logic ;
  tlv_sb_data_in_stall : in std_logic ) ;
  attribute _2_state_: integer;
  constant CKV_NUM_ENTRIES : integer := 32768 ;
  constant CKV_DATA_WIDTH : integer := 64 ;
  constant KIM_NUM_ENTRIES : integer := 16384 ;
  constant KIM_DATA_WIDTH : integer := 38 ;
  subtype pkt_hdr_e is std_logic_vector(1 downto 0) ;
  constant ENET : pkt_hdr_e := "00" ;
  constant IPV4 : pkt_hdr_e := "01" ;
  constant IPV6 : pkt_hdr_e := "10" ;
  constant MPLS : pkt_hdr_e := "11" ;
  subtype cmd_compound_cmd_frm_size_e is std_logic_vector(3 downto 0) ;
  constant CMD_SIMPLE : cmd_compound_cmd_frm_size_e := "0000" ;
  constant COMPND_4K : cmd_compound_cmd_frm_size_e := "0101" ;
  constant COMPND_8K : cmd_compound_cmd_frm_size_e := "0110" ;
  constant COMPND_RSV : cmd_compound_cmd_frm_size_e := "1111" ;
  subtype cmd_guid_present_e is std_logic_vector(0 downto 0) ;
  constant GUID_NOT_PRESENT : cmd_guid_present_e := "0" ;
  constant GUID_PRESENT : cmd_guid_present_e := "1" ;
  subtype cmd_frmd_crc_in_e is std_logic_vector(0 downto 0) ;
  constant CRC_NOT_PRESENT : cmd_frmd_crc_in_e := "0" ;
  constant CRC_PRESENT : cmd_frmd_crc_in_e := "1" ;
  subtype cceip_cmd_frmd_in_type_e is std_logic_vector(6 downto 0) ;
  constant CCEIP_FRMD_USER_NULL : cceip_cmd_frmd_in_type_e := "0001011" ;
  constant CCEIP_FRMD_USER_PI16 : cceip_cmd_frmd_in_type_e := "0001100" ;
  constant CCEIP_FRMD_USER_PI64 : cceip_cmd_frmd_in_type_e := "0001101" ;
  constant CCEIP_FRMD_USER_VM : cceip_cmd_frmd_in_type_e := "0001110" ;
  constant CCEIP_TYPE_IN_RSV : cceip_cmd_frmd_in_type_e := "1111111" ;
  subtype cddip_cmd_frmd_in_type_e is std_logic_vector(6 downto 0) ;
  constant CDDIP_FRMD_INT_APP : cddip_cmd_frmd_in_type_e := "0001111" ;
  constant CDDIP_FRMD_INT_SIP : cddip_cmd_frmd_in_type_e := "0010000" ;
  constant CDDIP_FRMD_INT_LIP : cddip_cmd_frmd_in_type_e := "0010001" ;
  constant CDDIP_FRMD_INT_VM : cddip_cmd_frmd_in_type_e := "0010010" ;
  constant CDDIP_FRMD_INT_VM_SHORT : cddip_cmd_frmd_in_type_e := "0010110" ;
  constant CDDIP_TYPE_IN_RSV : cddip_cmd_frmd_in_type_e := "1111111" ;
  subtype cceip_cmd_frmd_out_type_e is std_logic_vector(6 downto 0) ;
  constant CCEIP_FRMD_INT_APP : cceip_cmd_frmd_out_type_e := "0001111" ;
  constant CCEIP_FRMD_INT_SIP : cceip_cmd_frmd_out_type_e := "0010000" ;
  constant CCEIP_FRMD_INT_LIP : cceip_cmd_frmd_out_type_e := "0010001" ;
  constant CCEIP_FRMD_INT_VM : cceip_cmd_frmd_out_type_e := "0010010" ;
  constant CCEIP_FRMD_INT_VM_SHORT : cceip_cmd_frmd_out_type_e := "0010110" ;
  constant CCEIP_TYPE_OUT_RSV : cceip_cmd_frmd_out_type_e := "1111111" ;
  subtype cddip_cmd_frmd_out_type_e is std_logic_vector(6 downto 0) ;
  constant CDDIP_FRMD_USER_NULL : cddip_cmd_frmd_out_type_e := "0001011" ;
  constant CDDIP_FRMD_USER_PI16 : cddip_cmd_frmd_out_type_e := "0001100" ;
  constant CDDIP_FRMD_USER_PI64 : cddip_cmd_frmd_out_type_e := "0001101" ;
  constant CDDIP_FRMD_USER_VM : cddip_cmd_frmd_out_type_e := "0001110" ;
  constant CDDIP_TYPE_OUT_RSV : cddip_cmd_frmd_out_type_e := "1111111" ;
  subtype cmd_frmd_out_crc_e is std_logic_vector(0 downto 0) ;
  constant NOT_GEN : cmd_frmd_out_crc_e := "0" ;
  constant GEN : cmd_frmd_out_crc_e := "1" ;
  subtype cmd_frmd_out_crc_type_e is std_logic_vector(1 downto 0) ;
  constant FRMD_T10_DIX : cmd_frmd_out_crc_type_e := "00" ;
  constant FRMD_CRC64 : cmd_frmd_out_crc_type_e := "01" ;
  constant FRMD_CRC64E : cmd_frmd_out_crc_type_e := "10" ;
  constant FRMD_CRC_RSV : cmd_frmd_out_crc_type_e := "11" ;
  subtype cmd_md_type_e is std_logic_vector(1 downto 0) ;
  constant NO_CRC : cmd_md_type_e := "00" ;
  constant CRC_8B_CRC64 : cmd_md_type_e := "01" ;
  constant CRC_8B_CRC64E : cmd_md_type_e := "10" ;
  constant MD_TYPE_RSV : cmd_md_type_e := "11" ;
  subtype cmd_md_op_e is std_logic_vector(1 downto 0) ;
  constant CRC_GEN_VERIFY : cmd_md_op_e := "00" ;
  constant CRC_RSV1 : cmd_md_op_e := "01" ;
  constant CRC_RSV2 : cmd_md_op_e := "10" ;
  constant CRC_RSV3 : cmd_md_op_e := "11" ;
  subtype cmd_frmd_raw_mac_sel_e is std_logic_vector(0 downto 0) ;
  constant FRMD_MAC_NOP : cmd_frmd_raw_mac_sel_e := "0" ;
  constant FRMD_MAC_CAL : cmd_frmd_raw_mac_sel_e := "1" ;
  subtype cmd_chu_append_e is std_logic_vector(0 downto 0) ;
  constant CHU_NORMAL : cmd_chu_append_e := "0" ;
  constant CHU_APPEND : cmd_chu_append_e := "1" ;
  subtype cmd_comp_mode_e is std_logic_vector(3 downto 0) ;
  constant NONE : cmd_comp_mode_e := "0000" ;
  constant ZLIB : cmd_comp_mode_e := "0001" ;
  constant GZIP : cmd_comp_mode_e := "0010" ;
  constant XP9 : cmd_comp_mode_e := "0011" ;
  constant XP10 : cmd_comp_mode_e := "0100" ;
  constant CHU4K : cmd_comp_mode_e := "0101" ;
  constant CHU8K : cmd_comp_mode_e := "0110" ;
  constant RSV_MODE : cmd_comp_mode_e := "1111" ;
  subtype cmd_lz77_win_size_e is std_logic_vector(3 downto 0) ;
  constant WIN_32B : cmd_lz77_win_size_e := "0000" ;
  constant WIN_4K : cmd_lz77_win_size_e := "0001" ;
  constant WIN_8K : cmd_lz77_win_size_e := "0010" ;
  constant WIN_16K : cmd_lz77_win_size_e := "0011" ;
  constant WIN_32K : cmd_lz77_win_size_e := "0100" ;
  constant WIN_64K : cmd_lz77_win_size_e := "0101" ;
  constant RSV_WIN : cmd_lz77_win_size_e := "1111" ;
  subtype cmd_lz77_dly_match_win_e is std_logic_vector(1 downto 0) ;
  constant NO_MATCH : cmd_lz77_dly_match_win_e := "00" ;
  constant CHAR_1 : cmd_lz77_dly_match_win_e := "01" ;
  constant CHAR_2 : cmd_lz77_dly_match_win_e := "10" ;
  constant RSV_DLY : cmd_lz77_dly_match_win_e := "11" ;
  subtype cmd_lz77_min_match_len_e is std_logic_vector(0 downto 0) ;
  constant CHAR_3 : cmd_lz77_min_match_len_e := "0" ;
  constant CHAR_4 : cmd_lz77_min_match_len_e := "1" ;
  subtype cmd_lz77_max_symb_len_e is std_logic_vector(1 downto 0) ;
  constant LEN_LZ77_WIN : cmd_lz77_max_symb_len_e := "00" ;
  constant LEN_256B : cmd_lz77_max_symb_len_e := "01" ;
  constant MIN_MTCH_14 : cmd_lz77_max_symb_len_e := "10" ;
  constant LEN_64B : cmd_lz77_max_symb_len_e := "11" ;
  subtype cmd_xp10_prefix_mode_e is std_logic_vector(1 downto 0) ;
  constant NO_PREFIX : cmd_xp10_prefix_mode_e := "00" ;
  constant USER_PREFIX : cmd_xp10_prefix_mode_e := "01" ;
  constant PREDEF_PREFIX : cmd_xp10_prefix_mode_e := "10" ;
  constant PREDET_HUFF : cmd_xp10_prefix_mode_e := "11" ;
  subtype cmd_xp10_crc_mode_e is std_logic_vector(0 downto 0) ;
  constant CRC32 : cmd_xp10_crc_mode_e := "0" ;
  constant CRC64 : cmd_xp10_crc_mode_e := "1" ;
  subtype cmd_chu_comp_thrsh_e is std_logic_vector(1 downto 0) ;
  constant FRM : cmd_chu_comp_thrsh_e := "00" ;
  constant FRM_LESS_16 : cmd_chu_comp_thrsh_e := "01" ;
  constant INF : cmd_chu_comp_thrsh_e := "10" ;
  constant RSV_THRSH : cmd_chu_comp_thrsh_e := "11" ;
  subtype cmd_cipher_mode_e is std_logic_vector(0 downto 0) ;
  constant NO_CIPHER : cmd_cipher_mode_e := "0" ;
  constant CIPHER : cmd_cipher_mode_e := "1" ;
  subtype cmd_auth_op_e is std_logic_vector(3 downto 0) ;
  constant AUTH_NULL : cmd_auth_op_e := "0000" ;
  constant SHA2 : cmd_auth_op_e := "0001" ;
  constant HMAC_SHA2 : cmd_auth_op_e := "0010" ;
  constant AUTH_RSVD : cmd_auth_op_e := "1111" ;
  subtype cmd_cipher_op_e is std_logic_vector(3 downto 0) ;
  constant CPH_NULL : cmd_cipher_op_e := "0000" ;
  constant AES_GCM : cmd_cipher_op_e := "0001" ;
  constant AES_XTS_XEX : cmd_cipher_op_e := "0010" ;
  constant AES_GMAC : cmd_cipher_op_e := "0011" ;
  constant CPH_RSVD : cmd_cipher_op_e := "1111" ;
  subtype cmd_iv_src_e is std_logic_vector(1 downto 0) ;
  constant IV_NONE : cmd_iv_src_e := "00" ;
  constant IV_AUX_CMD : cmd_iv_src_e := "01" ;
  constant IV_KEYS : cmd_iv_src_e := "10" ;
  constant IV_AUX_FRMD : cmd_iv_src_e := "11" ;
  subtype cmd_iv_op_e is std_logic_vector(1 downto 0) ;
  constant IV_SRC : cmd_iv_op_e := "00" ;
  constant IV_RND : cmd_iv_op_e := "01" ;
  constant IV_INC : cmd_iv_op_e := "10" ;
  constant IV_RSV : cmd_iv_op_e := "11" ;
  subtype cmd_cipher_pad_e is std_logic_vector(0 downto 0) ;
  constant NO_PAD : cmd_cipher_pad_e := "0" ;
  constant PAD_16B : cmd_cipher_pad_e := "1" ;
  subtype cmd_digest_size_e is std_logic_vector(0 downto 0) ;
  constant DGST_256 : cmd_digest_size_e := "0" ;
  constant DGST_64 : cmd_digest_size_e := "1" ;
  subtype rqe_frame_type_e is std_logic_vector(0 downto 0) ;
  constant SIMPLE : rqe_frame_type_e := "0" ;
  constant COMPOUND : rqe_frame_type_e := "1" ;
  subtype rqe_trace_e is std_logic_vector(0 downto 0) ;
  constant TRACE_OFF : rqe_trace_e := "0" ;
  constant TRACE_ON : rqe_trace_e := "1" ;
  subtype rqe_frame_size_e is std_logic_vector(3 downto 0) ;
  constant RQE_SIMPLE : rqe_frame_size_e := "0000" ;
  constant RQE_COMPOUND_4K : rqe_frame_size_e := "0101" ;
  constant RQE_COMPOUND_8K : rqe_frame_size_e := "0110" ;
  constant RQE_RSV_FRAME_SIZE : rqe_frame_size_e := "1111" ;
  subtype frmd_coding_e is std_logic_vector(1 downto 0) ;
  constant PARSEABLE : frmd_coding_e := "00" ;
  constant RAW : frmd_coding_e := "01" ;
  constant XP10CFH4K : frmd_coding_e := "10" ;
  constant XP10CFH8K : frmd_coding_e := "11" ;
  subtype frmd_mac_size_e is std_logic_vector(1 downto 0) ;
  constant DIGEST_64b : frmd_mac_size_e := "00" ;
  constant DIGEST_128b : frmd_mac_size_e := "01" ;
  constant DIGEST_256b : frmd_mac_size_e := "10" ;
  constant DIGEST_0b : frmd_mac_size_e := "11" ;
  subtype tlv_types_e is std_logic_vector(7 downto 0) ;
  constant RQE : tlv_types_e := "00000000" ;
  constant CMD : tlv_types_e := "00000001" ;
  constant KEY : tlv_types_e := "00000010" ;
  constant PHD : tlv_types_e := "00000011" ;
  constant PFD : tlv_types_e := "00000100" ;
  constant DATA_UNK : tlv_types_e := "00000101" ;
  constant FTR : tlv_types_e := "00000110" ;
  constant LZ77 : tlv_types_e := "00000111" ;
  constant STAT : tlv_types_e := "00001000" ;
  constant CQE : tlv_types_e := "00001001" ;
  constant GUID : tlv_types_e := "00001010" ;
  constant FRMD_USER_NULL : tlv_types_e := "00001011" ;
  constant FRMD_USER_PI16 : tlv_types_e := "00001100" ;
  constant FRMD_USER_PI64 : tlv_types_e := "00001101" ;
  constant FRMD_USER_VM : tlv_types_e := "00001110" ;
  constant FRMD_INT_APP : tlv_types_e := "00001111" ;
  constant FRMD_INT_SIP : tlv_types_e := "00010000" ;
  constant FRMD_INT_LIP : tlv_types_e := "00010001" ;
  constant FRMD_INT_VM : tlv_types_e := "00010010" ;
  constant DATA : tlv_types_e := "00010011" ;
  constant CR_IV : tlv_types_e := "00010100" ;
  constant AUX_CMD : tlv_types_e := "00010101" ;
  constant FRMD_INT_VM_SHORT : tlv_types_e := "00010110" ;
  constant AUX_CMD_IV : tlv_types_e := "00010111" ;
  constant AUX_CMD_GUID : tlv_types_e := "00011000" ;
  constant AUX_CMD_GUID_IV : tlv_types_e := "00011001" ;
  constant SCH : tlv_types_e := "00011010" ;
  constant RSV_TLV : tlv_types_e := "11111111" ;
  subtype tlv_parse_action_e is std_logic_vector(1 downto 0) ;
  constant REP : tlv_parse_action_e := "00" ;
  constant PASS : tlv_parse_action_e := "01" ;
  constant MODIFY : tlv_parse_action_e := "10" ;
  constant DELETE : tlv_parse_action_e := "11" ;
  subtype tlvp_corrupt_e is std_logic_vector(0 downto 0) ;
  constant USER : tlvp_corrupt_e := "0" ;
  constant TLVP : tlvp_corrupt_e := "1" ;
  subtype cmd_type_e is std_logic_vector(0 downto 0) ;
  constant DATAPATH_CORRUPT : cmd_type_e := "0" ;
  constant FUNCTIONAL_ERROR : cmd_type_e := "1" ;
  subtype cmd_mode_e is std_logic_vector(1 downto 0) ;
  constant SINGLE_ERR : cmd_mode_e := "00" ;
  constant CONTINUOUS_ERROR : cmd_mode_e := "01" ;
  constant STOP : cmd_mode_e := "10" ;
  constant EOT : cmd_mode_e := "11" ;
  subtype aux_key_type_e is std_logic_vector(5 downto 0) ;
  constant NO_AUX_KEY : aux_key_type_e := "000000" ;
  constant AUX_KEY_ONLY : aux_key_type_e := "000001" ;
  constant DEK256 : aux_key_type_e := "000010" ;
  constant DEK512 : aux_key_type_e := "000011" ;
  constant DAK : aux_key_type_e := "000100" ;
  constant DEK256_DAK : aux_key_type_e := "000101" ;
  constant DEK512_DAK : aux_key_type_e := "000110" ;
  constant ENC_DEK256 : aux_key_type_e := "000111" ;
  constant ENC_DEK512 : aux_key_type_e := "001000" ;
  constant ENC_DAK : aux_key_type_e := "001001" ;
  constant ENC_DEK256_DAK : aux_key_type_e := "001010" ;
  constant ENC_DEK512_DAK : aux_key_type_e := "001011" ;
  constant ENC_DEK256_DAK_COMB : aux_key_type_e := "001100" ;
  constant ENC_DEK512_DAK_COMB : aux_key_type_e := "001101" ;
  constant KEY_TYPE_RSV : aux_key_type_e := "111111" ;
  subtype aux_kdf_mode_e is std_logic_vector(1 downto 0) ;
  constant KDF_MODE_GUID : aux_kdf_mode_e := "00" ;
  constant KDF_MODE_RGUID : aux_kdf_mode_e := "01" ;
  constant KDF_MODE_COMB_GUID : aux_kdf_mode_e := "10" ;
  constant KDF_MODE_COMB_RGUID : aux_kdf_mode_e := "11" ;
  subtype cceip_stats_e is std_logic_vector(9 downto 0) ;
  constant CKMIC_IV_MISMATCH_FRAME : cceip_stats_e := "0000000000" ;
  constant CKMIC_ENGINE_ID_MISMATCH_FRAME : cceip_stats_e := "0000000001" ;
  constant CKMIC_SEQ_ID_MISMATCH_FRAME : cceip_stats_e := "0000000010" ;
  constant CKMIC_HMAC_SHA256_TAG_FAIL_FRAME : cceip_stats_e := "0000000011" ;
  constant CKMIC_SHA256_TAG_FAIL_FRAME : cceip_stats_e := "0000000100" ;
  constant CKMIC_GMAC_TAG_FAIL_FRAME : cceip_stats_e := "0000000101" ;
  constant CKMIC_GCM_TAG_FAIL_FRAME : cceip_stats_e := "0000000110" ;
  constant CKMIC_AUTH_NOP_FRAME : cceip_stats_e := "0000000111" ;
  constant CKMIC_AUTH_HMAC_SHA256_FRAME : cceip_stats_e := "0000001000" ;
  constant CKMIC_AUTH_SHA256_FRAME : cceip_stats_e := "0000001001" ;
  constant CKMIC_AUTH_AES_GMAC_FRAME : cceip_stats_e := "0000001010" ;
  constant CKMIC_CIPH_NOP_FRAME : cceip_stats_e := "0000001011" ;
  constant CKMIC_CIPH_AES_XEX_FRAME : cceip_stats_e := "0000001100" ;
  constant CKMIC_CIPH_AES_XTS_FRAME : cceip_stats_e := "0000001101" ;
  constant CKMIC_CIPH_AES_GCM_FRAME : cceip_stats_e := "0000001110" ;
  constant CRCG0_RAW_CHSUM_GOOD_TOTAL : cceip_stats_e := "0001000000" ;
  constant CRCG0_RAW_CHSUM_ERROR_TOTAL : cceip_stats_e := "0001000001" ;
  constant CRCG0_CRC64E_CHSUM_GOOD_TOTAL : cceip_stats_e := "0001000010" ;
  constant CRCG0_CRC64E_CHSUM_ERROR_TOTAL : cceip_stats_e := "0001000011" ;
  constant CRCG0_ENC_CHSUM_GOOD_TOTAL : cceip_stats_e := "0001000100" ;
  constant CRCG0_ENC_CHSUM_ERROR_TOTAL : cceip_stats_e := "0001000101" ;
  constant CRCG0_NVME_CHSUM_GOOD_TOTAL : cceip_stats_e := "0001000110" ;
  constant CRCG0_NVME_CHSUM_ERROR_TOTAL : cceip_stats_e := "0001000111" ;
  constant CRCGC0_RAW_CHSUM_GOOD_TOTAL : cceip_stats_e := "0001001000" ;
  constant CRCGC0_RAW_CHSUM_ERROR_TOTAL : cceip_stats_e := "0001001001" ;
  constant CRCGC0_CRC64E_CHSUM_GOOD_TOTAL : cceip_stats_e := "0001001010" ;
  constant CRCGC0_CRC64E_CHSUM_ERROR_TOTAL : cceip_stats_e := "0001001011" ;
  constant CRCGC0_ENC_CHSUM_GOOD_TOTAL : cceip_stats_e := "0001001100" ;
  constant CRCGC0_ENC_CHSUM_ERROR_TOTAL : cceip_stats_e := "0001001101" ;
  constant CRCGC0_NVME_CHSUM_GOOD_TOTAL : cceip_stats_e := "0001001110" ;
  constant CRCGC0_NVME_CHSUM_ERROR_TOTAL : cceip_stats_e := "0001001111" ;
  constant CRCC1_RAW_CHSUM_GOOD_TOTAL : cceip_stats_e := "0001010000" ;
  constant CRCC1_RAW_CHSUM_ERROR_TOTAL : cceip_stats_e := "0001010001" ;
  constant CRCC1_CRC64E_CHSUM_GOOD_TOTAL : cceip_stats_e := "0001010010" ;
  constant CRCC1_CRC64E_CHSUM_ERROR_TOTAL : cceip_stats_e := "0001010011" ;
  constant CRCC1_ENC_CHSUM_GOOD_TOTAL : cceip_stats_e := "0001010100" ;
  constant CRCC1_ENC_CHSUM_ERROR_TOTAL : cceip_stats_e := "0001010101" ;
  constant CRCC1_NVME_CHSUM_GOOD_TOTAL : cceip_stats_e := "0001010110" ;
  constant CRCC1_NVME_CHSUM_ERROR_TOTAL : cceip_stats_e := "0001010111" ;
  constant CRCC0_RAW_CHSUM_GOOD_TOTAL : cceip_stats_e := "0001011000" ;
  constant CRCC0_RAW_CHSUM_ERROR_TOTAL : cceip_stats_e := "0001011001" ;
  constant CRCC0_CRC64E_CHSUM_GOOD_TOTAL : cceip_stats_e := "0001011010" ;
  constant CRCC0_CRC64E_CHSUM_ERROR_TOTAL : cceip_stats_e := "0001011011" ;
  constant CRCC0_ENC_CHSUM_GOOD_TOTAL : cceip_stats_e := "0001011100" ;
  constant CRCC0_ENC_CHSUM_ERROR_TOTAL : cceip_stats_e := "0001011101" ;
  constant CRCC0_NVME_CHSUM_GOOD_TOTAL : cceip_stats_e := "0001011110" ;
  constant CRCC0_NVME_CHSUM_ERROR_TOTAL : cceip_stats_e := "0001011111" ;
  constant CG_ENGINE_ERROR_COMMAND : cceip_stats_e := "0001100000" ;
  constant CG_SELECT_ENGINE_ERROR_COMMAND : cceip_stats_e := "0001100001" ;
  constant CG_SYSTEM_ERROR_COMMAND : cceip_stats_e := "0001100010" ;
  constant CG_CQE_OUTPUT_COMMAND : cceip_stats_e := "0001100011" ;
  constant HUFD_FE_XP9_FRM_TOTAL : cceip_stats_e := "0101000000" ;
  constant HUFD_FE_XP9_BLK_TOTAL : cceip_stats_e := "0101000001" ;
  constant HUFD_FE_XP9_RAW_FRM_TOTAL : cceip_stats_e := "0101000010" ;
  constant HUFD_FE_XP10_FRM_TOTAL : cceip_stats_e := "0101000011" ;
  constant HUFD_FE_XP10_FRM_PFX_TOTAL : cceip_stats_e := "0101000100" ;
  constant HUFD_FE_XP10_FRM_PDH_TOTAL : cceip_stats_e := "0101000101" ;
  constant HUFD_FE_XP10_BLK_TOTAL : cceip_stats_e := "0101000110" ;
  constant HUFD_FE_XP10_RAW_BLK_TOTAL : cceip_stats_e := "0101000111" ;
  constant HUFD_FE_GZIP_FRM_TOTAL : cceip_stats_e := "0101001000" ;
  constant HUFD_FE_GZIP_BLK_TOTAL : cceip_stats_e := "0101001001" ;
  constant HUFD_FE_GZIP_RAW_BLK_TOTAL : cceip_stats_e := "0101001010" ;
  constant HUFD_FE_ZLIB_FRM_TOTAL : cceip_stats_e := "0101001011" ;
  constant HUFD_FE_ZLIB_BLK_TOTAL : cceip_stats_e := "0101001100" ;
  constant HUFD_FE_ZLIB_RAW_BLK_TOTAL : cceip_stats_e := "0101001101" ;
  constant HUFD_FE_CHU4K_TOTAL : cceip_stats_e := "0101001110" ;
  constant HUFD_FE_CHU8K_TOTAL : cceip_stats_e := "0101001111" ;
  constant HUFD_FE_CHU4K_RAW_TOTAL : cceip_stats_e := "0101010000" ;
  constant HUFD_FE_CHU8K_RAW_TOTAL : cceip_stats_e := "0101010001" ;
  constant HUFD_FE_PFX_CRC_ERR_TOTAL : cceip_stats_e := "0101010010" ;
  constant HUFD_FE_PHD_CRC_ERR_TOTAL : cceip_stats_e := "0101010011" ;
  constant HUFD_FE_XP9_CRC_ERR_TOTAL : cceip_stats_e := "0101010100" ;
  constant HUFD_HTF_XP9_SIMPLE_SHORT_BLK_TOTAL : cceip_stats_e := "0101010101" ;
  constant HUFD_HTF_XP9_RETRO_SHORT_BLK_TOTAL : cceip_stats_e := "0101010110" ;
  constant HUFD_HTF_XP9_SIMPLE_LONG_BLK_TOTAL : cceip_stats_e := "0101010111" ;
  constant HUFD_HTF_XP9_RETRO_LONG_BLK_TOTAL : cceip_stats_e := "0101011000" ;
  constant HUFD_HTF_XP10_SIMPLE_SHORT_BLK_TOTAL : cceip_stats_e := "0101011001"
   ;
  constant HUFD_HTF_XP10_RETRO_SHORT_BLK_TOTAL : cceip_stats_e := "0101011010" ;
  constant HUFD_HTF_XP10_PREDEF_SHORT_BLK_TOTAL : cceip_stats_e := "0101011011"
   ;
  constant HUFD_HTF_XP10_SIMPLE_LONG_BLK_TOTAL : cceip_stats_e := "0101011100" ;
  constant HUFD_HTF_XP10_RETRO_LONG_BLK_TOTAL : cceip_stats_e := "0101011101" ;
  constant HUFD_HTF_XP10_PREDEF_LONG_BLK_TOTAL : cceip_stats_e := "0101011110" ;
  constant HUFD_HTF_CHU4K_SIMPLE_SHORT_BLK_TOTAL : cceip_stats_e := "0101011111"
   ;
  constant HUFD_HTF_CHU4K_RETRO_SHORT_BLK_TOTAL : cceip_stats_e := "0101100000"
   ;
  constant HUFD_HTF_CHU4K_PREDEF_SHORT_BLK_TOTAL : cceip_stats_e := "0101100001"
   ;
  constant HUFD_HTF_CHU4K_SIMPLE_LONG_BLK_TOTAL : cceip_stats_e := "0101100010"
   ;
  constant HUFD_HTF_CHU4K_RETRO_LONG_BLK_TOTAL : cceip_stats_e := "0101100011" ;
  constant HUFD_HTF_CHU4K_PREDEF_LONG_BLK_TOTAL : cceip_stats_e := "0101100100"
   ;
  constant HUFD_HTF_CHU8K_SIMPLE_SHORT_BLK_TOTAL : cceip_stats_e := "0101100101"
   ;
  constant HUFD_HTF_CHU8K_RETRO_SHORT_BLK_TOTAL : cceip_stats_e := "0101100110"
   ;
  constant HUFD_HTF_CHU8K_PREDEF_SHORT_BLK_TOTAL : cceip_stats_e := "0101100111"
   ;
  constant HUFD_HTF_CHU8K_SIMPLE_LONG_BLK_TOTAL : cceip_stats_e := "0101101000"
   ;
  constant HUFD_HTF_CHU8K_RETRO_LONG_BLK_TOTAL : cceip_stats_e := "0101101001" ;
  constant HUFD_HTF_CHU8K_PREDEF_LONG_BLK_TOTAL : cceip_stats_e := "0101101010"
   ;
  constant HUFD_HTF_DEFLATE_DYNAMIC_BLK_TOTAL : cceip_stats_e := "0101101011" ;
  constant HUFD_HTF_DEFLATE_FIXED_BLK_TOTAL : cceip_stats_e := "0101101100" ;
  constant HUFD_MTF_0_TOTAL : cceip_stats_e := "0101101101" ;
  constant HUFD_MTF_1_TOTAL : cceip_stats_e := "0101101110" ;
  constant HUFD_MTF_2_TOTAL : cceip_stats_e := "0101101111" ;
  constant HUFD_MTF_3_TOTAL : cceip_stats_e := "0101110000" ;
  constant HUFD_FE_FHP_STALL_TOTAL : cceip_stats_e := "0101110001" ;
  constant HUFD_FE_LFA_STALL_TOTAL : cceip_stats_e := "0101110010" ;
  constant HUFD_HTF_PREDEF_STALL_TOTAL : cceip_stats_e := "0101110011" ;
  constant HUFD_HTF_HDR_DATA_STALL_TOTAL : cceip_stats_e := "0101110100" ;
  constant HUFD_HTF_HDR_INFO_STALL_TOTAL : cceip_stats_e := "0101110101" ;
  constant HUFD_SDD_INPUT_STALL_TOTAL : cceip_stats_e := "0101110110" ;
  constant HUFD_SDD_BUF_FULL_STALL_TOTAL : cceip_stats_e := "0101110111" ;
  constant LZ77D_PTR_LEN_256_TOTAL : cceip_stats_e := "0110000000" ;
  constant LZ77D_PTR_LEN_128_TOTAL : cceip_stats_e := "0110000001" ;
  constant LZ77D_PTR_LEN_64_TOTAL : cceip_stats_e := "0110000010" ;
  constant LZ77D_PTR_LEN_32_TOTAL : cceip_stats_e := "0110000011" ;
  constant LZ77D_PTR_LEN_11_TOTAL : cceip_stats_e := "0110000100" ;
  constant LZ77D_PTR_LEN_10_TOTAL : cceip_stats_e := "0110000101" ;
  constant LZ77D_PTR_LEN_9_TOTAL : cceip_stats_e := "0110000110" ;
  constant LZ77D_PTR_LEN_8_TOTAL : cceip_stats_e := "0110000111" ;
  constant LZ77D_PTR_LEN_7_TOTAL : cceip_stats_e := "0110001000" ;
  constant LZ77D_PTR_LEN_6_TOTAL : cceip_stats_e := "0110001001" ;
  constant LZ77D_PTR_LEN_5_TOTAL : cceip_stats_e := "0110001010" ;
  constant LZ77D_PTR_LEN_4_TOTAL : cceip_stats_e := "0110001011" ;
  constant LZ77D_PTR_LEN_3_TOTAL : cceip_stats_e := "0110001100" ;
  constant LZ77D_LANE_1_LITERALS_TOTAL : cceip_stats_e := "0110001101" ;
  constant LZ77D_LANE_2_LITERALS_TOTAL : cceip_stats_e := "0110001110" ;
  constant LZ77D_LANE_3_LITERALS_TOTAL : cceip_stats_e := "0110001111" ;
  constant LZ77D_LANE_4_LITERALS_TOTAL : cceip_stats_e := "0110010000" ;
  constant LZ77D_PTRS_TOTAL : cceip_stats_e := "0110010001" ;
  constant LZ77D_FRM_IN_TOTAL : cceip_stats_e := "0110010010" ;
  constant LZ77D_FRM_OUT_TOTAL : cceip_stats_e := "0110010011" ;
  constant LZ77D_STALL_TOTAL : cceip_stats_e := "0110010100" ;
  constant DECRYPT_IV_MISMATCH_FRAME : cceip_stats_e := "0111000000" ;
  constant DECRYPT_ENGINE_ID_MISMATCH_FRAME : cceip_stats_e := "0111000001" ;
  constant DECRYPT_SEQ_ID_MISMATCH_FRAME : cceip_stats_e := "0111000010" ;
  constant DECRYPT_HMAC_SHA256_TAG_FAIL_FRAME : cceip_stats_e := "0111000011" ;
  constant DECRYPT_SHA256_TAG_FAIL_FRAME : cceip_stats_e := "0111000100" ;
  constant DECRYPT_GMAC_TAG_FAIL_FRAME : cceip_stats_e := "0111000101" ;
  constant DECRYPT_GCM_TAG_FAIL_FRAME : cceip_stats_e := "0111000110" ;
  constant DECRYPT_AUTH_NOP_FRAME : cceip_stats_e := "0111000111" ;
  constant DECRYPT_AUTH_HMAC_SHA256_FRAME : cceip_stats_e := "0111001000" ;
  constant DECRYPT_AUTH_SHA256_FRAME : cceip_stats_e := "0111001001" ;
  constant DECRYPT_AUTH_AES_GMAC_FRAME : cceip_stats_e := "0111001010" ;
  constant DECRYPT_CIPH_NOP_FRAME : cceip_stats_e := "0111001011" ;
  constant DECRYPT_CIPH_AES_XEX_FRAME : cceip_stats_e := "0111001100" ;
  constant DECRYPT_CIPH_AES_XTS_FRAME : cceip_stats_e := "0111001101" ;
  constant DECRYPT_CIPH_AES_GCM_FRAME : cceip_stats_e := "0111001110" ;
  constant OSF_DATA_INPUT_STALL_TOTAL : cceip_stats_e := "1000000000" ;
  constant OSF_CG_INPUT_STALL_TOTAL : cceip_stats_e := "1000000001" ;
  constant OSF_OUTPUT_BACKPRESSURE_TOTAL : cceip_stats_e := "1000000010" ;
  constant OSF_OUTPUT_STALL_TOTAL : cceip_stats_e := "1000000011" ;
  constant ENCRYPT_IV_MISMATCH_FRAME : cceip_stats_e := "1001000000" ;
  constant ENCRYPT_ENGINE_ID_MISMATCH_FRAME : cceip_stats_e := "1001000001" ;
  constant ENCRYPT_SEQ_ID_MISMATCH_FRAME : cceip_stats_e := "1001000010" ;
  constant ENCRYPT_HMAC_SHA256_TAG_FAIL_FRAME : cceip_stats_e := "1001000011" ;
  constant ENCRYPT_SHA256_TAG_FAIL_FRAME : cceip_stats_e := "1001000100" ;
  constant ENCRYPT_GMAC_TAG_FAIL_FRAME : cceip_stats_e := "1001000101" ;
  constant ENCRYPT_GCM_TAG_FAIL_FRAME : cceip_stats_e := "1001000110" ;
  constant ENCRYPT_AUTH_NOP_FRAME : cceip_stats_e := "1001000111" ;
  constant ENCRYPT_AUTH_HMAC_SHA256_FRAME : cceip_stats_e := "1001001000" ;
  constant ENCRYPT_AUTH_SHA256_FRAME : cceip_stats_e := "1001001001" ;
  constant ENCRYPT_AUTH_AES_GMAC_FRAME : cceip_stats_e := "1001001010" ;
  constant ENCRYPT_CIPH_NOP_FRAME : cceip_stats_e := "1001001011" ;
  constant ENCRYPT_CIPH_AES_XEX_FRAME : cceip_stats_e := "1001001100" ;
  constant ENCRYPT_CIPH_AES_XTS_FRAME : cceip_stats_e := "1001001101" ;
  constant ENCRYPT_CIPH_AES_GCM_FRAME : cceip_stats_e := "1001001110" ;
  constant SHORT_MAP_ERR_TOTAL : cceip_stats_e := "1010000000" ;
  constant LONG_MAP_ERR_TOTAL : cceip_stats_e := "1010000001" ;
  constant XP9_BLK_COMP_TOTAL : cceip_stats_e := "1010000010" ;
  constant XP9_FRM_RAW_TOTAL : cceip_stats_e := "1010000011" ;
  constant XP9_FRM_TOTAL : cceip_stats_e := "1010000100" ;
  constant XP9_BLK_SHORT_SIM_TOTAL : cceip_stats_e := "1010000101" ;
  constant XP9_BLK_LONG_SIM_TOTAL : cceip_stats_e := "1010000110" ;
  constant XP9_BLK_SHORT_RET_TOTAL : cceip_stats_e := "1010000111" ;
  constant XP9_BLK_LONG_RET_TOTAL : cceip_stats_e := "1010001000" ;
  constant XP10_BLK_COMP_TOTAL : cceip_stats_e := "1010001001" ;
  constant XP10_BLK_RAW_TOTAL : cceip_stats_e := "1010001010" ;
  constant XP10_BLK_SHORT_SIM_TOTAL : cceip_stats_e := "1010001011" ;
  constant XP10_BLK_LONG_SIM_TOTAL : cceip_stats_e := "1010001100" ;
  constant XP10_BLK_SHORT_RET_TOTAL : cceip_stats_e := "1010001101" ;
  constant XP10_BLK_LONG_RET_TOTAL : cceip_stats_e := "1010001110" ;
  constant XP10_BLK_SHORT_PRE_TOTAL : cceip_stats_e := "1010001111" ;
  constant XP10_BLK_LONG_PRE_TOTAL : cceip_stats_e := "1010010000" ;
  constant XP10_FRM_TOTAL : cceip_stats_e := "1010010001" ;
  constant CHU8_FRM_RAW_TOTAL : cceip_stats_e := "1010010010" ;
  constant CHU8_FRM_COMP_TOTAL : cceip_stats_e := "1010010011" ;
  constant CHU8_FRM_SHORT_SIM_TOTAL : cceip_stats_e := "1010010100" ;
  constant CHU8_FRM_LONG_SIM_TOTAL : cceip_stats_e := "1010010101" ;
  constant CHU8_FRM_SHORT_RET_TOTAL : cceip_stats_e := "1010010110" ;
  constant CHU8_FRM_LONG_RET_TOTAL : cceip_stats_e := "1010010111" ;
  constant CHU8_FRM_SHORT_PRE_TOTAL : cceip_stats_e := "1010011000" ;
  constant CHU8_FRM_LONG_PRE_TOTAL : cceip_stats_e := "1010011001" ;
  constant CHU8_CMD_TOTAL : cceip_stats_e := "1010011010" ;
  constant CHU4_FRM_RAW_TOTAL : cceip_stats_e := "1010011011" ;
  constant CHU4_FRM_COMP_TOTAL : cceip_stats_e := "1010011100" ;
  constant CHU4_FRM_SHORT_SIM_TOTAL : cceip_stats_e := "1010011101" ;
  constant CHU4_FRM_LONG_SIM_TOTAL : cceip_stats_e := "1010011110" ;
  constant CHU4_FRM_SHORT_RET_TOTAL : cceip_stats_e := "1010011111" ;
  constant CHU4_FRM_LONG_RET_TOTAL : cceip_stats_e := "1010100000" ;
  constant CHU4_FRM_SHORT_PRE_TOTAL : cceip_stats_e := "1010100001" ;
  constant CHU4_FRM_LONG_PRE_TOTAL : cceip_stats_e := "1010100010" ;
  constant CHU4_CMD_TOTAL : cceip_stats_e := "1010100011" ;
  constant DF_BLK_COMP_TOTAL : cceip_stats_e := "1010100100" ;
  constant DF_BLK_RAW_TOTAL : cceip_stats_e := "1010100101" ;
  constant DF_BLK_SHORT_SIM_TOTAL : cceip_stats_e := "1010100110" ;
  constant DF_BLK_LONG_SIM_TOTAL : cceip_stats_e := "1010100111" ;
  constant DF_BLK_SHORT_RET_TOTAL : cceip_stats_e := "1010101000" ;
  constant DF_BLK_LONG_RET_TOTAL : cceip_stats_e := "1010101001" ;
  constant DF_FRM_TOTAL : cceip_stats_e := "1010101010" ;
  constant PASS_THRU_FRM_TOTAL : cceip_stats_e := "1010101011" ;
  constant BYTE_0_TOTAL : cceip_stats_e := "1010101100" ;
  constant BYTE_1_TOTAL : cceip_stats_e := "1010101101" ;
  constant BYTE_2_TOTAL : cceip_stats_e := "1010101110" ;
  constant BYTE_3_TOTAL : cceip_stats_e := "1010101111" ;
  constant BYTE_4_TOTAL : cceip_stats_e := "1010110000" ;
  constant BYTE_5_TOTAL : cceip_stats_e := "1010110001" ;
  constant BYTE_6_TOTAL : cceip_stats_e := "1010110010" ;
  constant BYTE_7_TOTAL : cceip_stats_e := "1010110011" ;
  constant ENCRYPT_STALL_TOTAL : cceip_stats_e := "1010110100" ;
  constant LZ77_STALL_TOTAL : cceip_stats_e := "1010110101" ;
  constant LZ77C_eof_FRAME : cceip_stats_e := "1011000000" ;
  constant LZ77C_bypass_FRAME : cceip_stats_e := "1011000001" ;
  constant LZ77C_mtf_3_TOTAL : cceip_stats_e := "1011000010" ;
  constant LZ77C_mtf_2_TOTAL : cceip_stats_e := "1011000011" ;
  constant LZ77C_mtf_1_TOTAL : cceip_stats_e := "1011000100" ;
  constant LZ77C_mtf_0_TOTAL : cceip_stats_e := "1011000101" ;
  constant LZ77C_run_256_nup_TOTAL : cceip_stats_e := "1011000110" ;
  constant LZ77C_run_128_255_TOTAL : cceip_stats_e := "1011000111" ;
  constant LZ77C_run_64_127_TOTAL : cceip_stats_e := "1011001000" ;
  constant LZ77C_run_32_63_TOTAL : cceip_stats_e := "1011001001" ;
  constant LZ77C_run_11_31_TOTAL : cceip_stats_e := "1011001010" ;
  constant LZ77C_run_10_TOTAL : cceip_stats_e := "1011001011" ;
  constant LZ77C_run_9_TOTAL : cceip_stats_e := "1011001100" ;
  constant LZ77C_run_8_TOTAL : cceip_stats_e := "1011001101" ;
  constant LZ77C_run_7_TOTAL : cceip_stats_e := "1011001110" ;
  constant LZ77C_run_6_TOTAL : cceip_stats_e := "1011001111" ;
  constant LZ77C_run_5_TOTAL : cceip_stats_e := "1011010000" ;
  constant LZ77C_run_4_TOTAL : cceip_stats_e := "1011010001" ;
  constant LZ77C_run_3_TOTAL : cceip_stats_e := "1011010010" ;
  constant LZ77C_mtf_TOTAL : cceip_stats_e := "1011010011" ;
  constant LZ77C_ptr_TOTAL : cceip_stats_e := "1011010100" ;
  constant LZ77C_four_lit_TOTAL : cceip_stats_e := "1011010101" ;
  constant LZ77C_three_lit_TOTAL : cceip_stats_e := "1011010110" ;
  constant LZ77C_two_lit_TOTAL : cceip_stats_e := "1011010111" ;
  constant LZ77C_one_lit_TOTAL : cceip_stats_e := "1011011000" ;
  constant LZ77C_throttled_FRAME : cceip_stats_e := "1011011001" ;
  constant PREFIX_NUM_0_TOTAL : cceip_stats_e := "1101000000" ;
  constant PREFIX_NUM_1_TOTAL : cceip_stats_e := "1101000001" ;
  constant PREFIX_NUM_2_TOTAL : cceip_stats_e := "1101000010" ;
  constant PREFIX_NUM_3_TOTAL : cceip_stats_e := "1101000011" ;
  constant PREFIX_NUM_4_TOTAL : cceip_stats_e := "1101000100" ;
  constant PREFIX_NUM_5_TOTAL : cceip_stats_e := "1101000101" ;
  constant PREFIX_NUM_6_TOTAL : cceip_stats_e := "1101000110" ;
  constant PREFIX_NUM_7_TOTAL : cceip_stats_e := "1101000111" ;
  constant PREFIX_NUM_8_TOTAL : cceip_stats_e := "1101001000" ;
  constant PREFIX_NUM_9_TOTAL : cceip_stats_e := "1101001001" ;
  constant PREFIX_NUM_10_TOTAL : cceip_stats_e := "1101001010" ;
  constant PREFIX_NUM_11_TOTAL : cceip_stats_e := "1101001011" ;
  constant PREFIX_NUM_12_TOTAL : cceip_stats_e := "1101001100" ;
  constant PREFIX_NUM_13_TOTAL : cceip_stats_e := "1101001101" ;
  constant PREFIX_NUM_14_TOTAL : cceip_stats_e := "1101001110" ;
  constant PREFIX_NUM_15_TOTAL : cceip_stats_e := "1101001111" ;
  constant PREFIX_NUM_16_TOTAL : cceip_stats_e := "1101010000" ;
  constant PREFIX_NUM_17_TOTAL : cceip_stats_e := "1101010001" ;
  constant PREFIX_NUM_18_TOTAL : cceip_stats_e := "1101010010" ;
  constant PREFIX_NUM_19_TOTAL : cceip_stats_e := "1101010011" ;
  constant PREFIX_NUM_20_TOTAL : cceip_stats_e := "1101010100" ;
  constant PREFIX_NUM_21_TOTAL : cceip_stats_e := "1101010101" ;
  constant PREFIX_NUM_22_TOTAL : cceip_stats_e := "1101010110" ;
  constant PREFIX_NUM_23_TOTAL : cceip_stats_e := "1101010111" ;
  constant PREFIX_NUM_24_TOTAL : cceip_stats_e := "1101011000" ;
  constant PREFIX_NUM_25_TOTAL : cceip_stats_e := "1101011001" ;
  constant PREFIX_NUM_26_TOTAL : cceip_stats_e := "1101011010" ;
  constant PREFIX_NUM_27_TOTAL : cceip_stats_e := "1101011011" ;
  constant PREFIX_NUM_28_TOTAL : cceip_stats_e := "1101011100" ;
  constant PREFIX_NUM_29_TOTAL : cceip_stats_e := "1101011101" ;
  constant PREFIX_NUM_30_TOTAL : cceip_stats_e := "1101011110" ;
  constant PREFIX_NUM_31_TOTAL : cceip_stats_e := "1101011111" ;
  constant PREFIX_NUM_32_TOTAL : cceip_stats_e := "1101100000" ;
  constant PREFIX_NUM_33_TOTAL : cceip_stats_e := "1101100001" ;
  constant PREFIX_NUM_34_TOTAL : cceip_stats_e := "1101100010" ;
  constant PREFIX_NUM_35_TOTAL : cceip_stats_e := "1101100011" ;
  constant PREFIX_NUM_36_TOTAL : cceip_stats_e := "1101100100" ;
  constant PREFIX_NUM_37_TOTAL : cceip_stats_e := "1101100101" ;
  constant PREFIX_NUM_38_TOTAL : cceip_stats_e := "1101100110" ;
  constant PREFIX_NUM_39_TOTAL : cceip_stats_e := "1101100111" ;
  constant PREFIX_NUM_40_TOTAL : cceip_stats_e := "1101101000" ;
  constant PREFIX_NUM_41_TOTAL : cceip_stats_e := "1101101001" ;
  constant PREFIX_NUM_42_TOTAL : cceip_stats_e := "1101101010" ;
  constant PREFIX_NUM_43_TOTAL : cceip_stats_e := "1101101011" ;
  constant PREFIX_NUM_44_TOTAL : cceip_stats_e := "1101101100" ;
  constant PREFIX_NUM_45_TOTAL : cceip_stats_e := "1101101101" ;
  constant PREFIX_NUM_46_TOTAL : cceip_stats_e := "1101101110" ;
  constant PREFIX_NUM_47_TOTAL : cceip_stats_e := "1101101111" ;
  constant PREFIX_NUM_48_TOTAL : cceip_stats_e := "1101110000" ;
  constant PREFIX_NUM_49_TOTAL : cceip_stats_e := "1101110001" ;
  constant PREFIX_NUM_50_TOTAL : cceip_stats_e := "1101110010" ;
  constant PREFIX_NUM_51_TOTAL : cceip_stats_e := "1101110011" ;
  constant PREFIX_NUM_52_TOTAL : cceip_stats_e := "1101110100" ;
  constant PREFIX_NUM_53_TOTAL : cceip_stats_e := "1101110101" ;
  constant PREFIX_NUM_54_TOTAL : cceip_stats_e := "1101110110" ;
  constant PREFIX_NUM_55_TOTAL : cceip_stats_e := "1101110111" ;
  constant PREFIX_NUM_56_TOTAL : cceip_stats_e := "1101111000" ;
  constant PREFIX_NUM_57_TOTAL : cceip_stats_e := "1101111001" ;
  constant PREFIX_NUM_58_TOTAL : cceip_stats_e := "1101111010" ;
  constant PREFIX_NUM_59_TOTAL : cceip_stats_e := "1101111011" ;
  constant PREFIX_NUM_60_TOTAL : cceip_stats_e := "1101111100" ;
  constant PREFIX_NUM_61_TOTAL : cceip_stats_e := "1101111101" ;
  constant PREFIX_NUM_62_TOTAL : cceip_stats_e := "1101111110" ;
  constant PREFIX_NUM_63_TOTAL : cceip_stats_e := "1101111111" ;
  constant ISF_INPUT_COMMANDS : cceip_stats_e := "1110000000" ;
  constant ISF_INPUT_FRAMES : cceip_stats_e := "1110000001" ;
  constant ISF_INPUT_STALL_TOTAL : cceip_stats_e := "1110000010" ;
  constant ISF_INPUT_SYSTEM_STALL_TOTAL : cceip_stats_e := "1110000011" ;
  constant ISF_OUTPUT_BACKPRESSURE_TOTAL : cceip_stats_e := "1110000100" ;
  constant ISF_AUX_CMD_COMPRESS_CTL_MATCH_COMMAND_0 : cceip_stats_e :=
   "1110000101" ;
  constant ISF_AUX_CMD_COMPRESS_CTL_MATCH_COMMAND_1 : cceip_stats_e :=
   "1110000110" ;
  constant ISF_AUX_CMD_COMPRESS_CTL_MATCH_COMMAND_2 : cceip_stats_e :=
   "1110000111" ;
  constant ISF_AUX_CMD_COMPRESS_CTL_MATCH_COMMAND_3 : cceip_stats_e :=
   "1110001000" ;
  constant HUF_COMP_LZ77D_PTR_LEN_256_TOTAL : cceip_stats_e := "1111000000" ;
  constant HUF_COMP_LZ77D_PTR_LEN_128_TOTAL : cceip_stats_e := "1111000001" ;
  constant HUF_COMP_LZ77D_PTR_LEN_64_TOTAL : cceip_stats_e := "1111000010" ;
  constant HUF_COMP_LZ77D_PTR_LEN_32_TOTAL : cceip_stats_e := "1111000011" ;
  constant HUF_COMP_LZ77D_PTR_LEN_11_TOTAL : cceip_stats_e := "1111000100" ;
  constant HUF_COMP_LZ77D_PTR_LEN_10_TOTAL : cceip_stats_e := "1111000101" ;
  constant HUF_COMP_LZ77D_PTR_LEN_9_TOTAL : cceip_stats_e := "1111000110" ;
  constant HUF_COMP_LZ77D_PTR_LEN_8_TOTAL : cceip_stats_e := "1111000111" ;
  constant HUF_COMP_LZ77D_PTR_LEN_7_TOTAL : cceip_stats_e := "1111001000" ;
  constant HUF_COMP_LZ77D_PTR_LEN_6_TOTAL : cceip_stats_e := "1111001001" ;
  constant HUF_COMP_LZ77D_PTR_LEN_5_TOTAL : cceip_stats_e := "1111001010" ;
  constant HUF_COMP_LZ77D_PTR_LEN_4_TOTAL : cceip_stats_e := "1111001011" ;
  constant HUF_COMP_LZ77D_PTR_LEN_3_TOTAL : cceip_stats_e := "1111001100" ;
  constant HUF_COMP_LZ77D_LANE_4_LITERALS_TOTAL : cceip_stats_e := "1111001101"
   ;
  constant HUF_COMP_LZ77D_LANE_3_LITERALS_TOTAL : cceip_stats_e := "1111001110"
   ;
  constant HUF_COMP_LZ77D_LANE_2_LITERALS_TOTAL : cceip_stats_e := "1111001111"
   ;
  constant HUF_COMP_LZ77D_LANE_1_LITERALS_TOTAL : cceip_stats_e := "1111010000"
   ;
  constant HUF_COMP_LZ77D_PTRS_TOTAL : cceip_stats_e := "1111010001" ;
  constant HUF_COMP_LZ77D_FRM_IN_TOTAL : cceip_stats_e := "1111010010" ;
  constant HUF_COMP_LZ77D_FRM_OUT_TOTAL : cceip_stats_e := "1111010011" ;
  constant HUF_COMP_LZ77D_STALL_STB_TOTAL : cceip_stats_e := "1111010100" ;
  constant CCEIP_STATS_RESERVED : cceip_stats_e := "1111111111" ;
  subtype zipline_error_e is std_logic_vector(7 downto 0) ;
  constant NO_ERRORS : zipline_error_e := "00000000" ;
  constant CRCCG_CRC_ERROR : zipline_error_e := "00110010" ;
  constant CRCC0_CRC_ERROR : zipline_error_e := "00110011" ;
  constant CRCC1_CRC_ERROR : zipline_error_e := "00110100" ;
  constant CRCG0_CRC_ERROR : zipline_error_e := "00110101" ;
  constant CRCGC0_CRC_ERROR : zipline_error_e := "00110110" ;
  constant CRCDG0_CRC_ERROR : zipline_error_e := "00110111" ;
  constant CRCDC0_CRC_ERROR : zipline_error_e := "00111000" ;
  constant PREFIX_PC_OVERRUN_ERROR : zipline_error_e := "10010110" ;
  constant PREFIX_NUM_WR_ERROR : zipline_error_e := "10010111" ;
  constant PREFIX_ILLEGAL_OPCODE : zipline_error_e := "10011000" ;
  constant PREFIX_REC_US_SW_EN_ERROR : zipline_error_e := "10011001" ;
  constant PREFIX_ATTACH_PHD_CRC_ERROR : zipline_error_e := "10011011" ;
  constant PREFIX_ATTACH_PFD_CRC_ERROR : zipline_error_e := "10011100" ;
  constant LZ77_COMP_PREFIX_CRC_ERROR : zipline_error_e := "01000000" ;
  constant LZ77_COMP_INVALID_COMP_ALG : zipline_error_e := "01000001" ;
  constant LZ77_COMP_INVALID_WIN_SIZE : zipline_error_e := "01000010" ;
  constant LZ77_COMP_INVALID_MIN_LEN : zipline_error_e := "01000011" ;
  constant LZ77_COMP_INVALID_NUM_MTF : zipline_error_e := "01000100" ;
  constant LZ77_COMP_INVALID_MAX_LEN : zipline_error_e := "01000101" ;
  constant LZ77_COMP_INVALID_DMW_SIZE : zipline_error_e := "01000110" ;
  constant LZ77_COMP_LZ_ERROR : zipline_error_e := "01000111" ;
  constant HE_MEM_ECC : zipline_error_e := "01010000" ;
  constant HE_PDH_CRC : zipline_error_e := "01010001" ;
  constant HE_PFX_CRC : zipline_error_e := "01010010" ;
  constant HE_SYM_MAP_ERR : zipline_error_e := "01010011" ;
  constant CRYPTO_ENC_DRNG_HEALTH_FAIL : zipline_error_e := "01101100" ;
  constant CRYPTO_ENC_AAD_LEN_ERROR : zipline_error_e := "01101011" ;
  constant CRYPTO_ENC_XTS_LEN_ERROR : zipline_error_e := "01101010" ;
  constant CRYPTO_ENC_MAL_CMD : zipline_error_e := "01101001" ;
  constant CRYPTO_ENC_KEY_TLV_CRC_ERROR : zipline_error_e := "01101000" ;
  constant CRYPTO_ENC_INVALID_ENGINE_ID : zipline_error_e := "01100111" ;
  constant CRYPTO_ENC_INVALID_SEQNUM : zipline_error_e := "01100110" ;
  constant CRYPTO_ENC_IV_MISSING : zipline_error_e := "01100101" ;
  constant CRYPTO_ENC_SEED_EXPIRED : zipline_error_e := "01100100" ;
  constant CRYPTO_DEC_AAD_LEN_ERROR : zipline_error_e := "01110110" ;
  constant CRYPTO_DEC_XTS_LEN_ERROR : zipline_error_e := "01110101" ;
  constant CRYPTO_DEC_MAL_CMD : zipline_error_e := "01110100" ;
  constant CRYPTO_DEC_KEY_TLV_CRC_ERROR : zipline_error_e := "01110011" ;
  constant CRYPTO_DEC_INVALID_ENGINE_ID : zipline_error_e := "01110010" ;
  constant CRYPTO_DEC_INVALID_SEQNUM : zipline_error_e := "01110001" ;
  constant CRYPTO_DEC_IV_MISSING : zipline_error_e := "01110000" ;
  constant CRYPTO_DEC_TAG_MISCOMPARE : zipline_error_e := "01101110" ;
  constant CRYPTO_INT_KEY_TLV_CRC_ERROR : zipline_error_e := "01111011" ;
  constant CRYPTO_INT_INVALID_ENGINE_ID : zipline_error_e := "01111010" ;
  constant CRYPTO_INT_INVALID_SEQNUM : zipline_error_e := "01111001" ;
  constant CRYPTO_INT_TAG_MISCOMPARE : zipline_error_e := "01111000" ;
  constant KME_DAK_INV_KIM : zipline_error_e := "10000010" ;
  constant KME_DAK_PF_VF_VAL_ERR : zipline_error_e := "10000011" ;
  constant KME_DEK_INV_KIM : zipline_error_e := "10000100" ;
  constant KME_DEK_PF_VF_VAL_ERR : zipline_error_e := "10000101" ;
  constant KME_SEED_EXPIRED : zipline_error_e := "10000110" ;
  constant KME_DEK_GCM_TAG_FAIL : zipline_error_e := "10000111" ;
  constant KME_DAK_GCM_TAG_FAIL : zipline_error_e := "10001000" ;
  constant KME_ECC_FAIL : zipline_error_e := "10001001" ;
  constant KME_UNSUPPORTED_KEY_TYPE : zipline_error_e := "10001010" ;
  constant KME_DEK_ILLEGAL_KEK_USAGE : zipline_error_e := "10001011" ;
  constant KME_DAK_ILLEGAL_KEK_USAGE : zipline_error_e := "10001100" ;
  constant KME_DRNG_HEALTH_FAIL : zipline_error_e := "10001101" ;
  constant HD_MEM_ECC : zipline_error_e := "00000001" ;
  constant HD_FHP_PFX_CRC : zipline_error_e := "00000010" ;
  constant HD_FHP_PFX_DATA_ABSENT : zipline_error_e := "00000011" ;
  constant HD_FHP_PHD_CRC : zipline_error_e := "00000100" ;
  constant HD_FHP_BAD_FORMAT : zipline_error_e := "00000101" ;
  constant HD_BHP_INVALID_WSIZE : zipline_error_e := "00000110" ;
  constant HD_BHP_BLK_CRC : zipline_error_e := "00000111" ;
  constant HD_BHP_HDR_INVALID : zipline_error_e := "00001000" ;
  constant HD_BHP_XP9_HDR_SEQ : zipline_error_e := "00001001" ;
  constant HD_BHP_XP10_XTRA_FLAG_PRSNT : zipline_error_e := "00001010" ;
  constant HD_BHP_ZLIB_FDICT_PRSNT : zipline_error_e := "00001011" ;
  constant HD_BHP_GZ_CM_NOT_DEFLATE : zipline_error_e := "00001100" ;
  constant HD_BHP_ZLIB_CINFO_RANGE : zipline_error_e := "00001101" ;
  constant HD_BHP_ZLIB_FCHECK : zipline_error_e := "00001110" ;
  constant HD_BHP_DFLATE_LEN_CHECK : zipline_error_e := "00001111" ;
  constant HD_LFA_REWIND_FAIL : zipline_error_e := "00010000" ;
  constant HD_LFA_PREMATURE_EOF : zipline_error_e := "00010001" ;
  constant HD_LFA_LATE_EOF : zipline_error_e := "00010010" ;
  constant HD_LFA_MISSING_EOF : zipline_error_e := "00010011" ;
  constant HD_HTF_XP9_RESERVED_SYMBOL_TABLE_ENCODING : zipline_error_e :=
   "00010100" ;
  constant HD_HTF_XP10_RESERVED_SYMBOL_TABLE_ENCODING : zipline_error_e :=
   "00010101" ;
  constant HD_HTF_XP10_PREDEF_SYMBOL_TABLE_ENCODING : zipline_error_e :=
   "00010110" ;
  constant HD_HTF_XP9_ILLEGAL_NONZERO_BL : zipline_error_e := "00010111" ;
  constant HD_HTF_RLE_OVERRUN : zipline_error_e := "00011000" ;
  constant HD_HTF_BAD_HUFFMAN_CODE : zipline_error_e := "00011001" ;
  constant HD_HTF_ILLEGAL_SMALL_HUFFTREE : zipline_error_e := "00011010" ;
  constant HD_HTF_ILLEGAL_HUFFTREE : zipline_error_e := "00011011" ;
  constant HD_HTF_HDR_UNDERRUN : zipline_error_e := "00011100" ;
  constant HD_BHP_STBL_SIZE_ERR : zipline_error_e := "00011101" ;
  constant HD_SDD_INVALID_SYMBOL : zipline_error_e := "00100000" ;
  constant HD_SDD_END_MISMATCH : zipline_error_e := "00100001" ;
  constant HD_SDD_MISSING_EOB_SYM : zipline_error_e := "00100010" ;
  constant HD_MTF_XP9_MTF3_AFTER_BACKREF : zipline_error_e := "00100011" ;
  constant HD_MTF_XP10_MISSING_MTF : zipline_error_e := "00100100" ;
  constant HD_BHP_ILLEGAL_MTF_SZ : zipline_error_e := "00100101" ;
  constant HD_LZ_HBIF_SOFT_OFLOW : zipline_error_e := "00100110" ;
  constant HD_BE_FRM_CRC : zipline_error_e := "00100111" ;
  constant HD_BE_OLIMIT : zipline_error_e := "00101000" ;
  constant HD_BE_SZ_MISMATCH : zipline_error_e := "00101001" ;
  constant CG_UNDEF_FRMD_OUT : zipline_error_e := "10101010" ;
  constant ISF_PREFIX_ERR : zipline_error_e := "10110100" ;
  constant TLVP_BIP2_ERROR : zipline_error_e := "11111111" ;
  subtype kme_internal_idx is std_logic_vector(5 downto 0) ;
  constant IDX_KME_WORD0 : kme_internal_idx := std_logic_vector'("000000") ;
  constant IDX_KME_DEBUG_KEYHDR : kme_internal_idx := std_logic_vector'("000001"
  ) ;
  constant IDX_KME_GUID : kme_internal_idx := std_logic_vector'("000010") ;
  constant IDX_KME_IVTWEAK : kme_internal_idx := std_logic_vector'("000110") ;
  constant IDX_KME_KIM : kme_internal_idx := std_logic_vector'("001000") ;
  constant IDX_KME_DEK_CKV0 : kme_internal_idx := std_logic_vector'("001010") ;
  constant IDX_KME_DEK_CKV1 : kme_internal_idx := std_logic_vector'("001110") ;
  constant IDX_KME_DAK_CKV : kme_internal_idx := std_logic_vector'("010010") ;
  constant IDX_KME_EIV : kme_internal_idx := std_logic_vector'("010110") ;
  constant IDX_KME_DEK0 : kme_internal_idx := std_logic_vector'("011000") ;
  constant IDX_KME_DEK1 : kme_internal_idx := std_logic_vector'("011100") ;
  constant IDX_KME_ETAG : kme_internal_idx := std_logic_vector'("100000") ;
  constant IDX_KME_AIV : kme_internal_idx := std_logic_vector'("100010") ;
  constant IDX_KME_DAK : kme_internal_idx := std_logic_vector'("100100") ;
  constant IDX_KME_ATAG : kme_internal_idx := std_logic_vector'("101000") ;
  constant IDX_KME_ERROR : kme_internal_idx := std_logic_vector'("101010") ;
end cr_kme_kop_tlv_inspector_xcm69 ;
