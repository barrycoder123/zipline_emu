architecture module of ixc_assign is

begin

  process --:o53
  (*)
  begin
    L <= R ;
  end process ;
end module;
