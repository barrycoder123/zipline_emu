// xc_work/v/1.sv
// /home/ibarry/Project-Zipline-master/dv/KME/run/kme_tb.sv:12
// NOTE: This file corresponds to a module in the Software/TB partition.
`timescale 1ns/1ns
module kme_tb;
// external : kme_tb.kme_dut.clock_1 (resolved )  (var)  :(R)  
// external : apb_xactor.read (resolved )  (task)  
// external : apb_xactor.write (resolved )  (task)  
apb_xactor apb_xactor(,,,,,,,,,); 
cr_kme kme_dut(,,,,,,,,,,
  ,,,,,,,,,,
  ,,,,,,,,,,
  ,,,); 
endmodule

