library ieee, quickturn ;
use ieee.std_logic_1164.all ;
use quickturn.verilog.all ;
entity gfifo_conns is
  attribute _2_state_: integer;
end gfifo_conns ;
