ARCHITECTURE module OF ixc_assign_34 IS

BEGIN

  PROCESS --:o53
  (*)
  BEGIN
    L <= R ;
  END PROCESS ;
END module;