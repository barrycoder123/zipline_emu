
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module ixc_assign_296 ( L, R);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output [295:0] L;
input [295:0] R;
Q_ASSIGN U0 ( .B(R[0]), .A(L[0]));
Q_ASSIGN U1 ( .B(R[1]), .A(L[1]));
Q_ASSIGN U2 ( .B(R[2]), .A(L[2]));
Q_ASSIGN U3 ( .B(R[3]), .A(L[3]));
Q_ASSIGN U4 ( .B(R[4]), .A(L[4]));
Q_ASSIGN U5 ( .B(R[5]), .A(L[5]));
Q_ASSIGN U6 ( .B(R[6]), .A(L[6]));
Q_ASSIGN U7 ( .B(R[7]), .A(L[7]));
Q_ASSIGN U8 ( .B(R[8]), .A(L[8]));
Q_ASSIGN U9 ( .B(R[9]), .A(L[9]));
Q_ASSIGN U10 ( .B(R[10]), .A(L[10]));
Q_ASSIGN U11 ( .B(R[11]), .A(L[11]));
Q_ASSIGN U12 ( .B(R[12]), .A(L[12]));
Q_ASSIGN U13 ( .B(R[13]), .A(L[13]));
Q_ASSIGN U14 ( .B(R[14]), .A(L[14]));
Q_ASSIGN U15 ( .B(R[15]), .A(L[15]));
Q_ASSIGN U16 ( .B(R[16]), .A(L[16]));
Q_ASSIGN U17 ( .B(R[17]), .A(L[17]));
Q_ASSIGN U18 ( .B(R[18]), .A(L[18]));
Q_ASSIGN U19 ( .B(R[19]), .A(L[19]));
Q_ASSIGN U20 ( .B(R[20]), .A(L[20]));
Q_ASSIGN U21 ( .B(R[21]), .A(L[21]));
Q_ASSIGN U22 ( .B(R[22]), .A(L[22]));
Q_ASSIGN U23 ( .B(R[23]), .A(L[23]));
Q_ASSIGN U24 ( .B(R[24]), .A(L[24]));
Q_ASSIGN U25 ( .B(R[25]), .A(L[25]));
Q_ASSIGN U26 ( .B(R[26]), .A(L[26]));
Q_ASSIGN U27 ( .B(R[27]), .A(L[27]));
Q_ASSIGN U28 ( .B(R[28]), .A(L[28]));
Q_ASSIGN U29 ( .B(R[29]), .A(L[29]));
Q_ASSIGN U30 ( .B(R[30]), .A(L[30]));
Q_ASSIGN U31 ( .B(R[31]), .A(L[31]));
Q_ASSIGN U32 ( .B(R[32]), .A(L[32]));
Q_ASSIGN U33 ( .B(R[33]), .A(L[33]));
Q_ASSIGN U34 ( .B(R[34]), .A(L[34]));
Q_ASSIGN U35 ( .B(R[35]), .A(L[35]));
Q_ASSIGN U36 ( .B(R[36]), .A(L[36]));
Q_ASSIGN U37 ( .B(R[37]), .A(L[37]));
Q_ASSIGN U38 ( .B(R[38]), .A(L[38]));
Q_ASSIGN U39 ( .B(R[39]), .A(L[39]));
Q_ASSIGN U40 ( .B(R[40]), .A(L[40]));
Q_ASSIGN U41 ( .B(R[41]), .A(L[41]));
Q_ASSIGN U42 ( .B(R[42]), .A(L[42]));
Q_ASSIGN U43 ( .B(R[43]), .A(L[43]));
Q_ASSIGN U44 ( .B(R[44]), .A(L[44]));
Q_ASSIGN U45 ( .B(R[45]), .A(L[45]));
Q_ASSIGN U46 ( .B(R[46]), .A(L[46]));
Q_ASSIGN U47 ( .B(R[47]), .A(L[47]));
Q_ASSIGN U48 ( .B(R[48]), .A(L[48]));
Q_ASSIGN U49 ( .B(R[49]), .A(L[49]));
Q_ASSIGN U50 ( .B(R[50]), .A(L[50]));
Q_ASSIGN U51 ( .B(R[51]), .A(L[51]));
Q_ASSIGN U52 ( .B(R[52]), .A(L[52]));
Q_ASSIGN U53 ( .B(R[53]), .A(L[53]));
Q_ASSIGN U54 ( .B(R[54]), .A(L[54]));
Q_ASSIGN U55 ( .B(R[55]), .A(L[55]));
Q_ASSIGN U56 ( .B(R[56]), .A(L[56]));
Q_ASSIGN U57 ( .B(R[57]), .A(L[57]));
Q_ASSIGN U58 ( .B(R[58]), .A(L[58]));
Q_ASSIGN U59 ( .B(R[59]), .A(L[59]));
Q_ASSIGN U60 ( .B(R[60]), .A(L[60]));
Q_ASSIGN U61 ( .B(R[61]), .A(L[61]));
Q_ASSIGN U62 ( .B(R[62]), .A(L[62]));
Q_ASSIGN U63 ( .B(R[63]), .A(L[63]));
Q_ASSIGN U64 ( .B(R[64]), .A(L[64]));
Q_ASSIGN U65 ( .B(R[65]), .A(L[65]));
Q_ASSIGN U66 ( .B(R[66]), .A(L[66]));
Q_ASSIGN U67 ( .B(R[67]), .A(L[67]));
Q_ASSIGN U68 ( .B(R[68]), .A(L[68]));
Q_ASSIGN U69 ( .B(R[69]), .A(L[69]));
Q_ASSIGN U70 ( .B(R[70]), .A(L[70]));
Q_ASSIGN U71 ( .B(R[71]), .A(L[71]));
Q_ASSIGN U72 ( .B(R[72]), .A(L[72]));
Q_ASSIGN U73 ( .B(R[73]), .A(L[73]));
Q_ASSIGN U74 ( .B(R[74]), .A(L[74]));
Q_ASSIGN U75 ( .B(R[75]), .A(L[75]));
Q_ASSIGN U76 ( .B(R[76]), .A(L[76]));
Q_ASSIGN U77 ( .B(R[77]), .A(L[77]));
Q_ASSIGN U78 ( .B(R[78]), .A(L[78]));
Q_ASSIGN U79 ( .B(R[79]), .A(L[79]));
Q_ASSIGN U80 ( .B(R[80]), .A(L[80]));
Q_ASSIGN U81 ( .B(R[81]), .A(L[81]));
Q_ASSIGN U82 ( .B(R[82]), .A(L[82]));
Q_ASSIGN U83 ( .B(R[83]), .A(L[83]));
Q_ASSIGN U84 ( .B(R[84]), .A(L[84]));
Q_ASSIGN U85 ( .B(R[85]), .A(L[85]));
Q_ASSIGN U86 ( .B(R[86]), .A(L[86]));
Q_ASSIGN U87 ( .B(R[87]), .A(L[87]));
Q_ASSIGN U88 ( .B(R[88]), .A(L[88]));
Q_ASSIGN U89 ( .B(R[89]), .A(L[89]));
Q_ASSIGN U90 ( .B(R[90]), .A(L[90]));
Q_ASSIGN U91 ( .B(R[91]), .A(L[91]));
Q_ASSIGN U92 ( .B(R[92]), .A(L[92]));
Q_ASSIGN U93 ( .B(R[93]), .A(L[93]));
Q_ASSIGN U94 ( .B(R[94]), .A(L[94]));
Q_ASSIGN U95 ( .B(R[95]), .A(L[95]));
Q_ASSIGN U96 ( .B(R[96]), .A(L[96]));
Q_ASSIGN U97 ( .B(R[97]), .A(L[97]));
Q_ASSIGN U98 ( .B(R[98]), .A(L[98]));
Q_ASSIGN U99 ( .B(R[99]), .A(L[99]));
Q_ASSIGN U100 ( .B(R[100]), .A(L[100]));
Q_ASSIGN U101 ( .B(R[101]), .A(L[101]));
Q_ASSIGN U102 ( .B(R[102]), .A(L[102]));
Q_ASSIGN U103 ( .B(R[103]), .A(L[103]));
Q_ASSIGN U104 ( .B(R[104]), .A(L[104]));
Q_ASSIGN U105 ( .B(R[105]), .A(L[105]));
Q_ASSIGN U106 ( .B(R[106]), .A(L[106]));
Q_ASSIGN U107 ( .B(R[107]), .A(L[107]));
Q_ASSIGN U108 ( .B(R[108]), .A(L[108]));
Q_ASSIGN U109 ( .B(R[109]), .A(L[109]));
Q_ASSIGN U110 ( .B(R[110]), .A(L[110]));
Q_ASSIGN U111 ( .B(R[111]), .A(L[111]));
Q_ASSIGN U112 ( .B(R[112]), .A(L[112]));
Q_ASSIGN U113 ( .B(R[113]), .A(L[113]));
Q_ASSIGN U114 ( .B(R[114]), .A(L[114]));
Q_ASSIGN U115 ( .B(R[115]), .A(L[115]));
Q_ASSIGN U116 ( .B(R[116]), .A(L[116]));
Q_ASSIGN U117 ( .B(R[117]), .A(L[117]));
Q_ASSIGN U118 ( .B(R[118]), .A(L[118]));
Q_ASSIGN U119 ( .B(R[119]), .A(L[119]));
Q_ASSIGN U120 ( .B(R[120]), .A(L[120]));
Q_ASSIGN U121 ( .B(R[121]), .A(L[121]));
Q_ASSIGN U122 ( .B(R[122]), .A(L[122]));
Q_ASSIGN U123 ( .B(R[123]), .A(L[123]));
Q_ASSIGN U124 ( .B(R[124]), .A(L[124]));
Q_ASSIGN U125 ( .B(R[125]), .A(L[125]));
Q_ASSIGN U126 ( .B(R[126]), .A(L[126]));
Q_ASSIGN U127 ( .B(R[127]), .A(L[127]));
Q_ASSIGN U128 ( .B(R[128]), .A(L[128]));
Q_ASSIGN U129 ( .B(R[129]), .A(L[129]));
Q_ASSIGN U130 ( .B(R[130]), .A(L[130]));
Q_ASSIGN U131 ( .B(R[131]), .A(L[131]));
Q_ASSIGN U132 ( .B(R[132]), .A(L[132]));
Q_ASSIGN U133 ( .B(R[133]), .A(L[133]));
Q_ASSIGN U134 ( .B(R[134]), .A(L[134]));
Q_ASSIGN U135 ( .B(R[135]), .A(L[135]));
Q_ASSIGN U136 ( .B(R[136]), .A(L[136]));
Q_ASSIGN U137 ( .B(R[137]), .A(L[137]));
Q_ASSIGN U138 ( .B(R[138]), .A(L[138]));
Q_ASSIGN U139 ( .B(R[139]), .A(L[139]));
Q_ASSIGN U140 ( .B(R[140]), .A(L[140]));
Q_ASSIGN U141 ( .B(R[141]), .A(L[141]));
Q_ASSIGN U142 ( .B(R[142]), .A(L[142]));
Q_ASSIGN U143 ( .B(R[143]), .A(L[143]));
Q_ASSIGN U144 ( .B(R[144]), .A(L[144]));
Q_ASSIGN U145 ( .B(R[145]), .A(L[145]));
Q_ASSIGN U146 ( .B(R[146]), .A(L[146]));
Q_ASSIGN U147 ( .B(R[147]), .A(L[147]));
Q_ASSIGN U148 ( .B(R[148]), .A(L[148]));
Q_ASSIGN U149 ( .B(R[149]), .A(L[149]));
Q_ASSIGN U150 ( .B(R[150]), .A(L[150]));
Q_ASSIGN U151 ( .B(R[151]), .A(L[151]));
Q_ASSIGN U152 ( .B(R[152]), .A(L[152]));
Q_ASSIGN U153 ( .B(R[153]), .A(L[153]));
Q_ASSIGN U154 ( .B(R[154]), .A(L[154]));
Q_ASSIGN U155 ( .B(R[155]), .A(L[155]));
Q_ASSIGN U156 ( .B(R[156]), .A(L[156]));
Q_ASSIGN U157 ( .B(R[157]), .A(L[157]));
Q_ASSIGN U158 ( .B(R[158]), .A(L[158]));
Q_ASSIGN U159 ( .B(R[159]), .A(L[159]));
Q_ASSIGN U160 ( .B(R[160]), .A(L[160]));
Q_ASSIGN U161 ( .B(R[161]), .A(L[161]));
Q_ASSIGN U162 ( .B(R[162]), .A(L[162]));
Q_ASSIGN U163 ( .B(R[163]), .A(L[163]));
Q_ASSIGN U164 ( .B(R[164]), .A(L[164]));
Q_ASSIGN U165 ( .B(R[165]), .A(L[165]));
Q_ASSIGN U166 ( .B(R[166]), .A(L[166]));
Q_ASSIGN U167 ( .B(R[167]), .A(L[167]));
Q_ASSIGN U168 ( .B(R[168]), .A(L[168]));
Q_ASSIGN U169 ( .B(R[169]), .A(L[169]));
Q_ASSIGN U170 ( .B(R[170]), .A(L[170]));
Q_ASSIGN U171 ( .B(R[171]), .A(L[171]));
Q_ASSIGN U172 ( .B(R[172]), .A(L[172]));
Q_ASSIGN U173 ( .B(R[173]), .A(L[173]));
Q_ASSIGN U174 ( .B(R[174]), .A(L[174]));
Q_ASSIGN U175 ( .B(R[175]), .A(L[175]));
Q_ASSIGN U176 ( .B(R[176]), .A(L[176]));
Q_ASSIGN U177 ( .B(R[177]), .A(L[177]));
Q_ASSIGN U178 ( .B(R[178]), .A(L[178]));
Q_ASSIGN U179 ( .B(R[179]), .A(L[179]));
Q_ASSIGN U180 ( .B(R[180]), .A(L[180]));
Q_ASSIGN U181 ( .B(R[181]), .A(L[181]));
Q_ASSIGN U182 ( .B(R[182]), .A(L[182]));
Q_ASSIGN U183 ( .B(R[183]), .A(L[183]));
Q_ASSIGN U184 ( .B(R[184]), .A(L[184]));
Q_ASSIGN U185 ( .B(R[185]), .A(L[185]));
Q_ASSIGN U186 ( .B(R[186]), .A(L[186]));
Q_ASSIGN U187 ( .B(R[187]), .A(L[187]));
Q_ASSIGN U188 ( .B(R[188]), .A(L[188]));
Q_ASSIGN U189 ( .B(R[189]), .A(L[189]));
Q_ASSIGN U190 ( .B(R[190]), .A(L[190]));
Q_ASSIGN U191 ( .B(R[191]), .A(L[191]));
Q_ASSIGN U192 ( .B(R[192]), .A(L[192]));
Q_ASSIGN U193 ( .B(R[193]), .A(L[193]));
Q_ASSIGN U194 ( .B(R[194]), .A(L[194]));
Q_ASSIGN U195 ( .B(R[195]), .A(L[195]));
Q_ASSIGN U196 ( .B(R[196]), .A(L[196]));
Q_ASSIGN U197 ( .B(R[197]), .A(L[197]));
Q_ASSIGN U198 ( .B(R[198]), .A(L[198]));
Q_ASSIGN U199 ( .B(R[199]), .A(L[199]));
Q_ASSIGN U200 ( .B(R[200]), .A(L[200]));
Q_ASSIGN U201 ( .B(R[201]), .A(L[201]));
Q_ASSIGN U202 ( .B(R[202]), .A(L[202]));
Q_ASSIGN U203 ( .B(R[203]), .A(L[203]));
Q_ASSIGN U204 ( .B(R[204]), .A(L[204]));
Q_ASSIGN U205 ( .B(R[205]), .A(L[205]));
Q_ASSIGN U206 ( .B(R[206]), .A(L[206]));
Q_ASSIGN U207 ( .B(R[207]), .A(L[207]));
Q_ASSIGN U208 ( .B(R[208]), .A(L[208]));
Q_ASSIGN U209 ( .B(R[209]), .A(L[209]));
Q_ASSIGN U210 ( .B(R[210]), .A(L[210]));
Q_ASSIGN U211 ( .B(R[211]), .A(L[211]));
Q_ASSIGN U212 ( .B(R[212]), .A(L[212]));
Q_ASSIGN U213 ( .B(R[213]), .A(L[213]));
Q_ASSIGN U214 ( .B(R[214]), .A(L[214]));
Q_ASSIGN U215 ( .B(R[215]), .A(L[215]));
Q_ASSIGN U216 ( .B(R[216]), .A(L[216]));
Q_ASSIGN U217 ( .B(R[217]), .A(L[217]));
Q_ASSIGN U218 ( .B(R[218]), .A(L[218]));
Q_ASSIGN U219 ( .B(R[219]), .A(L[219]));
Q_ASSIGN U220 ( .B(R[220]), .A(L[220]));
Q_ASSIGN U221 ( .B(R[221]), .A(L[221]));
Q_ASSIGN U222 ( .B(R[222]), .A(L[222]));
Q_ASSIGN U223 ( .B(R[223]), .A(L[223]));
Q_ASSIGN U224 ( .B(R[224]), .A(L[224]));
Q_ASSIGN U225 ( .B(R[225]), .A(L[225]));
Q_ASSIGN U226 ( .B(R[226]), .A(L[226]));
Q_ASSIGN U227 ( .B(R[227]), .A(L[227]));
Q_ASSIGN U228 ( .B(R[228]), .A(L[228]));
Q_ASSIGN U229 ( .B(R[229]), .A(L[229]));
Q_ASSIGN U230 ( .B(R[230]), .A(L[230]));
Q_ASSIGN U231 ( .B(R[231]), .A(L[231]));
Q_ASSIGN U232 ( .B(R[232]), .A(L[232]));
Q_ASSIGN U233 ( .B(R[233]), .A(L[233]));
Q_ASSIGN U234 ( .B(R[234]), .A(L[234]));
Q_ASSIGN U235 ( .B(R[235]), .A(L[235]));
Q_ASSIGN U236 ( .B(R[236]), .A(L[236]));
Q_ASSIGN U237 ( .B(R[237]), .A(L[237]));
Q_ASSIGN U238 ( .B(R[238]), .A(L[238]));
Q_ASSIGN U239 ( .B(R[239]), .A(L[239]));
Q_ASSIGN U240 ( .B(R[240]), .A(L[240]));
Q_ASSIGN U241 ( .B(R[241]), .A(L[241]));
Q_ASSIGN U242 ( .B(R[242]), .A(L[242]));
Q_ASSIGN U243 ( .B(R[243]), .A(L[243]));
Q_ASSIGN U244 ( .B(R[244]), .A(L[244]));
Q_ASSIGN U245 ( .B(R[245]), .A(L[245]));
Q_ASSIGN U246 ( .B(R[246]), .A(L[246]));
Q_ASSIGN U247 ( .B(R[247]), .A(L[247]));
Q_ASSIGN U248 ( .B(R[248]), .A(L[248]));
Q_ASSIGN U249 ( .B(R[249]), .A(L[249]));
Q_ASSIGN U250 ( .B(R[250]), .A(L[250]));
Q_ASSIGN U251 ( .B(R[251]), .A(L[251]));
Q_ASSIGN U252 ( .B(R[252]), .A(L[252]));
Q_ASSIGN U253 ( .B(R[253]), .A(L[253]));
Q_ASSIGN U254 ( .B(R[254]), .A(L[254]));
Q_ASSIGN U255 ( .B(R[255]), .A(L[255]));
Q_ASSIGN U256 ( .B(R[256]), .A(L[256]));
Q_ASSIGN U257 ( .B(R[257]), .A(L[257]));
Q_ASSIGN U258 ( .B(R[258]), .A(L[258]));
Q_ASSIGN U259 ( .B(R[259]), .A(L[259]));
Q_ASSIGN U260 ( .B(R[260]), .A(L[260]));
Q_ASSIGN U261 ( .B(R[261]), .A(L[261]));
Q_ASSIGN U262 ( .B(R[262]), .A(L[262]));
Q_ASSIGN U263 ( .B(R[263]), .A(L[263]));
Q_ASSIGN U264 ( .B(R[264]), .A(L[264]));
Q_ASSIGN U265 ( .B(R[265]), .A(L[265]));
Q_ASSIGN U266 ( .B(R[266]), .A(L[266]));
Q_ASSIGN U267 ( .B(R[267]), .A(L[267]));
Q_ASSIGN U268 ( .B(R[268]), .A(L[268]));
Q_ASSIGN U269 ( .B(R[269]), .A(L[269]));
Q_ASSIGN U270 ( .B(R[270]), .A(L[270]));
Q_ASSIGN U271 ( .B(R[271]), .A(L[271]));
Q_ASSIGN U272 ( .B(R[272]), .A(L[272]));
Q_ASSIGN U273 ( .B(R[273]), .A(L[273]));
Q_ASSIGN U274 ( .B(R[274]), .A(L[274]));
Q_ASSIGN U275 ( .B(R[275]), .A(L[275]));
Q_ASSIGN U276 ( .B(R[276]), .A(L[276]));
Q_ASSIGN U277 ( .B(R[277]), .A(L[277]));
Q_ASSIGN U278 ( .B(R[278]), .A(L[278]));
Q_ASSIGN U279 ( .B(R[279]), .A(L[279]));
Q_ASSIGN U280 ( .B(R[280]), .A(L[280]));
Q_ASSIGN U281 ( .B(R[281]), .A(L[281]));
Q_ASSIGN U282 ( .B(R[282]), .A(L[282]));
Q_ASSIGN U283 ( .B(R[283]), .A(L[283]));
Q_ASSIGN U284 ( .B(R[284]), .A(L[284]));
Q_ASSIGN U285 ( .B(R[285]), .A(L[285]));
Q_ASSIGN U286 ( .B(R[286]), .A(L[286]));
Q_ASSIGN U287 ( .B(R[287]), .A(L[287]));
Q_ASSIGN U288 ( .B(R[288]), .A(L[288]));
Q_ASSIGN U289 ( .B(R[289]), .A(L[289]));
Q_ASSIGN U290 ( .B(R[290]), .A(L[290]));
Q_ASSIGN U291 ( .B(R[291]), .A(L[291]));
Q_ASSIGN U292 ( .B(R[292]), .A(L[292]));
Q_ASSIGN U293 ( .B(R[293]), .A(L[293]));
Q_ASSIGN U294 ( .B(R[294]), .A(L[294]));
Q_ASSIGN U295 ( .B(R[295]), .A(L[295]));
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE "ixc_assign"
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE_LIB "IXCOM_TEMP_LIBRARY"
endmodule
