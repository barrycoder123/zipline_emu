
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
(* celldefine = 1 *) 
module nx_indirect_access_cntrl_xcm111 ( clk, rst_n, wr_stb, reg_addr, cmnd_op, 
	cmnd_addr, cmnd_table_id, stat_code, stat_datawords, stat_addr, 
	stat_table_id, capability_lst, capability_type, enable, .addr_limit( {
	\addr_limit[0][4] , \addr_limit[0][3] , \addr_limit[0][2] , 
	\addr_limit[0][1] , \addr_limit[0][0] } ), wr_dat, rd_dat, sw_cs, 
	sw_ce, sw_we, sw_add, sw_wdat, sw_rdat, sw_match, sw_aindex, grant, 
	yield, reset);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
input clk;
input rst_n;
input wr_stb;
input [10:0] reg_addr;
input [3:0] cmnd_op;
input [4:0] cmnd_addr;
input [0:0] cmnd_table_id;
output [2:0] stat_code;
output [4:0] stat_datawords;
output [4:0] stat_addr;
output [0:0] stat_table_id;
output [15:0] capability_lst;
output [3:0] capability_type;
output enable;
input \addr_limit[0][4] ;
input \addr_limit[0][3] ;
input \addr_limit[0][2] ;
input \addr_limit[0][1] ;
input \addr_limit[0][0] ;
input [31:0] wr_dat;
output [31:0] rd_dat;
output sw_cs;
output sw_ce;
output sw_we;
output [4:0] sw_add;
output [31:0] sw_wdat;
input [31:0] sw_rdat;
input sw_match;
input [3:0] sw_aindex;
input grant;
output yield;
output reset;
wire [0:2] _zy_simnet_stat_code_0_w$;
wire [0:4] _zy_simnet_stat_datawords_1_w$;
wire [0:4] _zy_simnet_stat_addr_2_w$;
wire _zy_simnet_stat_table_id_3_w$;
wire [0:15] _zy_simnet_capability_lst_4_w$;
wire [0:3] _zy_simnet_capability_type_5_w$;
wire _zy_simnet_enable_6_w$;
wire [0:31] _zy_simnet_rd_dat_7_w$;
wire _zy_simnet_sw_cs_8_w$;
wire _zy_simnet_sw_ce_9_w$;
wire _zy_simnet_sw_we_10_w$;
wire [0:4] _zy_simnet_sw_add_11_w$;
wire [0:31] _zy_simnet_sw_wdat_12_w$;
wire _zy_simnet_yield_13_w$;
wire _zy_simnet_reset_14_w$;
wire [3:0] cmnd;
wire init_r;
wire [0:0] inc_r;
wire init_inc_r;
wire sw_cs_r;
wire sw_ce_r;
wire rst_r;
wire rst_or_ini_r;
wire [4:0] rst_addr_r;
wire sw_we_r;
wire cmnd_rd_stb;
wire cmnd_wr_stb;
wire cmnd_ena_stb;
wire cmnd_dis_stb;
wire cmnd_rst_stb;
wire cmnd_ini_stb;
wire cmnd_inc_stb;
wire cmnd_sis_stb;
wire cmnd_tmo_stb;
wire cmnd_cmp_stb;
wire cmnd_issued;
wire ack_error;
wire unsupported_op;
wire [3:0] state_r;
wire [0:0] timer_r;
wire timeout;
wire sim_tmo_r;
wire [4:0] maxaddr;
wire badaddr;
wire igrant;
wire [2:0] stat;
supply0 n1;
supply1 n2;
Q_BUF U0 ( .A(timer_r[0]), .Z(timeout));
Q_BUF U1 ( .A(n1), .Z(stat_datawords[0]));
Q_BUF U2 ( .A(n1), .Z(stat_datawords[1]));
Q_BUF U3 ( .A(n1), .Z(stat_datawords[2]));
Q_BUF U4 ( .A(n1), .Z(stat_datawords[3]));
Q_BUF U5 ( .A(n1), .Z(stat_datawords[4]));
Q_BUF U6 ( .A(n1), .Z(capability_type[0]));
Q_BUF U7 ( .A(n2), .Z(capability_type[1]));
Q_BUF U8 ( .A(n1), .Z(capability_type[2]));
Q_BUF U9 ( .A(n1), .Z(capability_type[3]));
Q_BUF U10 ( .A(n2), .Z(capability_lst[0]));
Q_BUF U11 ( .A(n2), .Z(capability_lst[1]));
Q_BUF U12 ( .A(n2), .Z(capability_lst[2]));
Q_BUF U13 ( .A(n1), .Z(capability_lst[3]));
Q_BUF U14 ( .A(n1), .Z(capability_lst[4]));
Q_BUF U15 ( .A(n2), .Z(capability_lst[5]));
Q_BUF U16 ( .A(n1), .Z(capability_lst[6]));
Q_BUF U17 ( .A(n1), .Z(capability_lst[7]));
Q_BUF U18 ( .A(n1), .Z(capability_lst[8]));
Q_BUF U19 ( .A(n1), .Z(capability_lst[9]));
Q_BUF U20 ( .A(n1), .Z(capability_lst[10]));
Q_BUF U21 ( .A(n1), .Z(capability_lst[11]));
Q_BUF U22 ( .A(n1), .Z(capability_lst[12]));
Q_BUF U23 ( .A(n1), .Z(capability_lst[13]));
Q_BUF U24 ( .A(n1), .Z(capability_lst[14]));
Q_BUF U25 ( .A(n2), .Z(capability_lst[15]));
Q_BUF U26 ( .A(n1), .Z(stat_table_id[0]));
ixc_assign_3 _zz_strnp_7 ( stat[2:0], stat_code[2:0]);
ixc_assign_4 _zz_strnp_1 ( cmnd[3:0], cmnd_op[3:0]);
ixc_assign \genblk1._zz_strnp_0 ( reset, rst_r);
ixc_context_read_6 _zzixc_ctxrd_0 ( { stat_code[2], stat_code[1], 
	stat_code[0], stat[2], stat[1], stat[0]});
ixc_assign _zz_strnp_22 ( _zy_simnet_reset_14_w$, reset);
ixc_assign _zz_strnp_21 ( _zy_simnet_yield_13_w$, yield);
ixc_assign_32 _zz_strnp_20 ( _zy_simnet_sw_wdat_12_w$[0:31], sw_wdat[31:0]);
ixc_assign_5 _zz_strnp_19 ( _zy_simnet_sw_add_11_w$[0:4], sw_add[4:0]);
ixc_assign _zz_strnp_18 ( _zy_simnet_sw_we_10_w$, sw_we);
ixc_assign _zz_strnp_17 ( _zy_simnet_sw_ce_9_w$, sw_ce);
ixc_assign _zz_strnp_16 ( _zy_simnet_sw_cs_8_w$, sw_cs);
ixc_assign_32 _zz_strnp_15 ( _zy_simnet_rd_dat_7_w$[0:31], rd_dat[31:0]);
ixc_assign _zz_strnp_14 ( _zy_simnet_enable_6_w$, enable);
ixc_assign_4 _zz_strnp_13 ( _zy_simnet_capability_type_5_w$[0:3], { n1, n1, 
	n2, n1});
ixc_assign_16 _zz_strnp_12 ( _zy_simnet_capability_lst_4_w$[0:15], { n2, n1, 
	n1, n1, n1, n1, n1, n1, n1, n1, n2, n1, n1, n2, n2, n2});
ixc_assign _zz_strnp_11 ( _zy_simnet_stat_table_id_3_w$, n1);
ixc_assign_5 _zz_strnp_10 ( _zy_simnet_stat_addr_2_w$[0:4], stat_addr[4:0]);
ixc_assign_5 _zz_strnp_9 ( _zy_simnet_stat_datawords_1_w$[0:4], { n1, n1, n1, 
	n1, n1});
ixc_assign_3 _zz_strnp_8 ( _zy_simnet_stat_code_0_w$[0:2], stat_code[2:0]);
ixc_assign_5 _zz_strnp_6 ( stat_addr[4:0], maxaddr[4:0]);
Q_AN02 U47 ( .A0(n19), .A1(grant), .Z(igrant));
Q_AN02 U48 ( .A0(cmnd_issued), .A1(n18), .Z(badaddr));
Q_AO21 U49 ( .A0(n15), .A1(n17), .B0(n14), .Z(n18));
Q_AN02 U50 ( .A0(cmnd_addr[0]), .A1(n16), .Z(n17));
Q_INV U51 ( .A(maxaddr[0]), .Z(n16));
Q_OR03 U52 ( .A0(n11), .A1(n10), .A2(n13), .Z(n14));
Q_OA21 U53 ( .A0(cmnd_addr[1]), .A1(n7), .B0(n9), .Z(n15));
Q_AN03 U54 ( .A0(cmnd_addr[1]), .A1(n7), .A2(n9), .Z(n10));
Q_INV U55 ( .A(maxaddr[1]), .Z(n7));
Q_OA21 U56 ( .A0(cmnd_addr[2]), .A1(n6), .B0(n8), .Z(n9));
Q_AN03 U57 ( .A0(cmnd_addr[2]), .A1(n6), .A2(n8), .Z(n11));
Q_INV U58 ( .A(maxaddr[2]), .Z(n6));
Q_OA21 U59 ( .A0(cmnd_addr[3]), .A1(n5), .B0(n4), .Z(n8));
Q_AN03 U60 ( .A0(cmnd_addr[3]), .A1(n5), .A2(n4), .Z(n12));
Q_INV U61 ( .A(maxaddr[3]), .Z(n5));
Q_OR02 U62 ( .A0(cmnd_addr[4]), .A1(n3), .Z(n4));
Q_AO21 U63 ( .A0(cmnd_addr[4]), .A1(n3), .B0(n12), .Z(n13));
Q_INV U64 ( .A(maxaddr[4]), .Z(n3));
ixc_assign _zz_strnp_5 ( yield, timeout);
ixc_assign _zz_strnp_4 ( sw_we, sw_we_r);
ixc_assign _zz_strnp_3 ( sw_ce, sw_ce_r);
ixc_assign _zz_strnp_2 ( sw_cs, sw_cs_r);
Q_MX02 U69 ( .S(rst_or_ini_r), .A0(cmnd_addr[0]), .A1(rst_addr_r[0]), .Z(sw_add[0]));
Q_MX02 U70 ( .S(rst_or_ini_r), .A0(cmnd_addr[1]), .A1(rst_addr_r[1]), .Z(sw_add[1]));
Q_MX02 U71 ( .S(rst_or_ini_r), .A0(cmnd_addr[2]), .A1(rst_addr_r[2]), .Z(sw_add[2]));
Q_MX02 U72 ( .S(rst_or_ini_r), .A0(cmnd_addr[3]), .A1(rst_addr_r[3]), .Z(sw_add[3]));
Q_MX02 U73 ( .S(rst_or_ini_r), .A0(cmnd_addr[4]), .A1(rst_addr_r[4]), .Z(sw_add[4]));
Q_AN02 U74 ( .A0(enable), .A1(\addr_limit[0][0] ), .Z(maxaddr[0]));
Q_AN02 U75 ( .A0(enable), .A1(\addr_limit[0][1] ), .Z(maxaddr[1]));
Q_AN02 U76 ( .A0(enable), .A1(\addr_limit[0][2] ), .Z(maxaddr[2]));
Q_AN02 U77 ( .A0(enable), .A1(\addr_limit[0][3] ), .Z(maxaddr[3]));
Q_AN02 U78 ( .A0(enable), .A1(\addr_limit[0][4] ), .Z(maxaddr[4]));
Q_INV U79 ( .A(reg_addr[2]), .Z(n20));
Q_INV U80 ( .A(reg_addr[4]), .Z(n21));
Q_INV U81 ( .A(reg_addr[6]), .Z(n22));
Q_INV U82 ( .A(reg_addr[10]), .Z(n23));
Q_OR03 U83 ( .A0(n23), .A1(reg_addr[9]), .A2(reg_addr[8]), .Z(n24));
Q_OR03 U84 ( .A0(reg_addr[7]), .A1(n22), .A2(reg_addr[5]), .Z(n25));
Q_OR03 U85 ( .A0(n21), .A1(reg_addr[3]), .A2(n20), .Z(n26));
Q_OR03 U86 ( .A0(reg_addr[1]), .A1(reg_addr[0]), .A2(n24), .Z(n27));
Q_NR03 U87 ( .A0(n25), .A1(n26), .A2(n27), .Z(n28));
Q_AN02 U88 ( .A0(wr_stb), .A1(n28), .Z(n52));
Q_INV U89 ( .A(n47), .Z(cmnd_issued));
Q_INV U90 ( .A(unsupported_op), .Z(n46));
Q_OA21 U91 ( .A0(n30), .A1(n31), .B0(n29), .Z(unsupported_op));
Q_AN02 U92 ( .A0(n29), .A1(n32), .Z(ack_error));
Q_AO21 U93 ( .A0(n34), .A1(n35), .B0(n33), .Z(n47));
Q_INV U94 ( .A(n52), .Z(n33));
Q_MX02 U95 ( .S(cmnd[3]), .A0(n38), .A1(n36), .Z(n34));
Q_INV U96 ( .A(cmnd_cmp_stb), .Z(n48));
Q_AN02 U97 ( .A0(n29), .A1(n39), .Z(cmnd_cmp_stb));
Q_AN02 U98 ( .A0(n29), .A1(n40), .Z(cmnd_tmo_stb));
Q_AN03 U99 ( .A0(n29), .A1(n35), .A2(n38), .Z(cmnd_sis_stb));
Q_AN02 U100 ( .A0(n52), .A1(cmnd[3]), .Z(n29));
Q_AN02 U101 ( .A0(n41), .A1(n32), .Z(cmnd_inc_stb));
Q_AN02 U102 ( .A0(n36), .A1(cmnd[0]), .Z(n32));
Q_AN02 U103 ( .A0(n41), .A1(n40), .Z(cmnd_ini_stb));
Q_AN02 U104 ( .A0(n36), .A1(n35), .Z(n40));
Q_AN02 U105 ( .A0(cmnd[2]), .A1(cmnd[1]), .Z(n36));
Q_INV U106 ( .A(cmnd_rst_stb), .Z(n49));
Q_AN02 U107 ( .A0(n31), .A1(n42), .Z(cmnd_rst_stb));
Q_AN02 U108 ( .A0(n41), .A1(cmnd[0]), .Z(n42));
Q_AN02 U109 ( .A0(n31), .A1(n43), .Z(cmnd_dis_stb));
Q_AN02 U110 ( .A0(n41), .A1(n35), .Z(n43));
Q_AN02 U111 ( .A0(cmnd[2]), .A1(n44), .Z(n31));
Q_AN02 U112 ( .A0(n30), .A1(n42), .Z(cmnd_ena_stb));
Q_INV U113 ( .A(cmnd_wr_stb), .Z(n50));
Q_AN02 U114 ( .A0(n30), .A1(n43), .Z(cmnd_wr_stb));
Q_INV U115 ( .A(cmnd[0]), .Z(n35));
Q_AN02 U116 ( .A0(n45), .A1(cmnd[1]), .Z(n30));
Q_INV U117 ( .A(cmnd_rd_stb), .Z(n51));
Q_AN02 U118 ( .A0(n41), .A1(n39), .Z(cmnd_rd_stb));
Q_AN02 U119 ( .A0(n38), .A1(cmnd[0]), .Z(n39));
Q_NR02 U120 ( .A0(cmnd[2]), .A1(cmnd[1]), .Z(n38));
Q_INV U121 ( .A(cmnd[1]), .Z(n44));
Q_INV U122 ( .A(cmnd[2]), .Z(n45));
Q_AN02 U123 ( .A0(n52), .A1(n37), .Z(n41));
Q_INV U124 ( .A(cmnd[3]), .Z(n37));
Q_OR02 U125 ( .A0(cmnd_ini_stb), .A1(cmnd_inc_stb), .Z(n320));
Q_XNR2 U126 ( .A0(rst_addr_r[0]), .A1(cmnd_addr[0]), .Z(n54));
Q_XNR2 U127 ( .A0(rst_addr_r[1]), .A1(cmnd_addr[1]), .Z(n55));
Q_XNR2 U128 ( .A0(rst_addr_r[2]), .A1(cmnd_addr[2]), .Z(n56));
Q_XNR2 U129 ( .A0(rst_addr_r[3]), .A1(cmnd_addr[3]), .Z(n57));
Q_XNR2 U130 ( .A0(rst_addr_r[4]), .A1(cmnd_addr[4]), .Z(n58));
Q_AN03 U131 ( .A0(n58), .A1(n57), .A2(n56), .Z(n59));
Q_AN03 U132 ( .A0(n55), .A1(n54), .A2(n59), .Z(n321));
Q_AN02 U133 ( .A0(init_inc_r), .A1(igrant), .Z(n60));
Q_XOR2 U134 ( .A0(inc_r[0]), .A1(n60), .Z(n61));
Q_AD01HF U135 ( .A0(rst_addr_r[0]), .B0(igrant), .S(n62), .CO(n63));
Q_AD01HF U136 ( .A0(rst_addr_r[1]), .B0(n63), .S(n64), .CO(n65));
Q_AD01HF U137 ( .A0(rst_addr_r[2]), .B0(n65), .S(n66), .CO(n67));
Q_AD01HF U138 ( .A0(rst_addr_r[3]), .B0(n67), .S(n68), .CO(n69));
Q_XOR2 U139 ( .A0(rst_addr_r[4]), .A1(n69), .Z(n70));
Q_MX02 U140 ( .S(n239), .A0(n76), .A1(n72), .Z(n71));
Q_ND02 U141 ( .A0(n73), .A1(n74), .Z(n72));
Q_ND02 U142 ( .A0(n298), .A1(n204), .Z(n74));
Q_OR02 U143 ( .A0(n75), .A1(n204), .Z(n73));
Q_OR02 U144 ( .A0(n204), .A1(n300), .Z(n76));
Q_INV U145 ( .A(n77), .Z(n78));
Q_MX02 U146 ( .S(n239), .A0(n73), .A1(n79), .Z(n77));
Q_INV U147 ( .A(n80), .Z(n79));
Q_INV U148 ( .A(n81), .Z(n82));
Q_MX02 U149 ( .S(n239), .A0(n88), .A1(n83), .Z(n81));
Q_INV U150 ( .A(n84), .Z(n83));
Q_MX02 U151 ( .S(n204), .A0(n80), .A1(n85), .Z(n84));
Q_INV U152 ( .A(n86), .Z(n85));
Q_XOR2 U153 ( .A0(n298), .A1(n87), .Z(n80));
Q_OR02 U154 ( .A0(n299), .A1(n75), .Z(n88));
Q_OR02 U155 ( .A0(n298), .A1(n300), .Z(n75));
Q_NR02 U156 ( .A0(n301), .A1(n90), .Z(n89));
Q_MX02 U157 ( .S(n204), .A0(n86), .A1(n300), .Z(n90));
Q_OR02 U158 ( .A0(n298), .A1(n87), .Z(n86));
Q_INV U159 ( .A(n300), .Z(n87));
Q_AN03 U160 ( .A0(n299), .A1(n298), .A2(n301), .Z(n91));
Q_AO21 U161 ( .A0(n91), .A1(state_r[3]), .B0(n89), .Z(n325));
Q_AO21 U162 ( .A0(n91), .A1(state_r[2]), .B0(n82), .Z(n324));
Q_AO21 U163 ( .A0(n91), .A1(state_r[1]), .B0(n78), .Z(n323));
Q_AO21 U164 ( .A0(n91), .A1(state_r[0]), .B0(n71), .Z(n322));
Q_AN02 U165 ( .A0(n303), .A1(cmnd_addr[0]), .Z(n93));
Q_MX02 U166 ( .S(n304), .A0(n93), .A1(n62), .Z(n94));
Q_AN02 U167 ( .A0(n303), .A1(cmnd_addr[1]), .Z(n95));
Q_MX02 U168 ( .S(n304), .A0(n95), .A1(n64), .Z(n96));
Q_AN02 U169 ( .A0(n303), .A1(cmnd_addr[2]), .Z(n97));
Q_MX02 U170 ( .S(n304), .A0(n97), .A1(n66), .Z(n98));
Q_AN02 U171 ( .A0(n303), .A1(cmnd_addr[3]), .Z(n99));
Q_MX02 U172 ( .S(n304), .A0(n99), .A1(n68), .Z(n100));
Q_AN02 U173 ( .A0(n303), .A1(cmnd_addr[4]), .Z(n101));
Q_MX02 U174 ( .S(n304), .A0(n101), .A1(n70), .Z(n102));
Q_AN02 U175 ( .A0(n309), .A1(n61), .Z(n103));
Q_MX03 U176 ( .S0(n311), .S1(n312), .A0(sw_aindex[0]), .A1(wr_dat[0]), .A2(sw_rdat[0]), .Z(n104));
Q_MX03 U177 ( .S0(n311), .S1(n312), .A0(sw_aindex[1]), .A1(wr_dat[1]), .A2(sw_rdat[1]), .Z(n105));
Q_MX03 U178 ( .S0(n311), .S1(n312), .A0(sw_aindex[2]), .A1(wr_dat[2]), .A2(sw_rdat[2]), .Z(n106));
Q_MX03 U179 ( .S0(n311), .S1(n312), .A0(sw_aindex[3]), .A1(wr_dat[3]), .A2(sw_rdat[3]), .Z(n107));
Q_MX03 U180 ( .S0(n311), .S1(n312), .A0(sw_match), .A1(wr_dat[4]), .A2(sw_rdat[4]), .Z(n108));
Q_AN02 U181 ( .A0(n311), .A1(wr_dat[5]), .Z(n109));
Q_MX02 U182 ( .S(n312), .A0(n109), .A1(sw_rdat[5]), .Z(n110));
Q_AN02 U183 ( .A0(n311), .A1(wr_dat[6]), .Z(n111));
Q_MX02 U184 ( .S(n312), .A0(n111), .A1(sw_rdat[6]), .Z(n112));
Q_AN02 U185 ( .A0(n311), .A1(wr_dat[7]), .Z(n113));
Q_MX02 U186 ( .S(n312), .A0(n113), .A1(sw_rdat[7]), .Z(n114));
Q_AN02 U187 ( .A0(n311), .A1(wr_dat[8]), .Z(n115));
Q_MX02 U188 ( .S(n312), .A0(n115), .A1(sw_rdat[8]), .Z(n116));
Q_AN02 U189 ( .A0(n311), .A1(wr_dat[9]), .Z(n117));
Q_MX02 U190 ( .S(n312), .A0(n117), .A1(sw_rdat[9]), .Z(n118));
Q_AN02 U191 ( .A0(n311), .A1(wr_dat[10]), .Z(n119));
Q_MX02 U192 ( .S(n312), .A0(n119), .A1(sw_rdat[10]), .Z(n120));
Q_AN02 U193 ( .A0(n311), .A1(wr_dat[11]), .Z(n121));
Q_MX02 U194 ( .S(n312), .A0(n121), .A1(sw_rdat[11]), .Z(n122));
Q_AN02 U195 ( .A0(n311), .A1(wr_dat[12]), .Z(n123));
Q_MX02 U196 ( .S(n312), .A0(n123), .A1(sw_rdat[12]), .Z(n124));
Q_AN02 U197 ( .A0(n311), .A1(wr_dat[13]), .Z(n125));
Q_MX02 U198 ( .S(n312), .A0(n125), .A1(sw_rdat[13]), .Z(n126));
Q_AN02 U199 ( .A0(n311), .A1(wr_dat[14]), .Z(n127));
Q_MX02 U200 ( .S(n312), .A0(n127), .A1(sw_rdat[14]), .Z(n128));
Q_AN02 U201 ( .A0(n311), .A1(wr_dat[15]), .Z(n129));
Q_MX02 U202 ( .S(n312), .A0(n129), .A1(sw_rdat[15]), .Z(n130));
Q_AN02 U203 ( .A0(n311), .A1(wr_dat[16]), .Z(n131));
Q_MX02 U204 ( .S(n312), .A0(n131), .A1(sw_rdat[16]), .Z(n132));
Q_AN02 U205 ( .A0(n311), .A1(wr_dat[17]), .Z(n133));
Q_MX02 U206 ( .S(n312), .A0(n133), .A1(sw_rdat[17]), .Z(n134));
Q_AN02 U207 ( .A0(n311), .A1(wr_dat[18]), .Z(n135));
Q_MX02 U208 ( .S(n312), .A0(n135), .A1(sw_rdat[18]), .Z(n136));
Q_AN02 U209 ( .A0(n311), .A1(wr_dat[19]), .Z(n137));
Q_MX02 U210 ( .S(n312), .A0(n137), .A1(sw_rdat[19]), .Z(n138));
Q_AN02 U211 ( .A0(n311), .A1(wr_dat[20]), .Z(n139));
Q_MX02 U212 ( .S(n312), .A0(n139), .A1(sw_rdat[20]), .Z(n140));
Q_AN02 U213 ( .A0(n311), .A1(wr_dat[21]), .Z(n141));
Q_MX02 U214 ( .S(n312), .A0(n141), .A1(sw_rdat[21]), .Z(n142));
Q_AN02 U215 ( .A0(n311), .A1(wr_dat[22]), .Z(n143));
Q_MX02 U216 ( .S(n312), .A0(n143), .A1(sw_rdat[22]), .Z(n144));
Q_AN02 U217 ( .A0(n311), .A1(wr_dat[23]), .Z(n145));
Q_MX02 U218 ( .S(n312), .A0(n145), .A1(sw_rdat[23]), .Z(n146));
Q_AN02 U219 ( .A0(n311), .A1(wr_dat[24]), .Z(n147));
Q_MX02 U220 ( .S(n312), .A0(n147), .A1(sw_rdat[24]), .Z(n148));
Q_AN02 U221 ( .A0(n311), .A1(wr_dat[25]), .Z(n149));
Q_MX02 U222 ( .S(n312), .A0(n149), .A1(sw_rdat[25]), .Z(n150));
Q_AN02 U223 ( .A0(n311), .A1(wr_dat[26]), .Z(n151));
Q_MX02 U224 ( .S(n312), .A0(n151), .A1(sw_rdat[26]), .Z(n152));
Q_AN02 U225 ( .A0(n311), .A1(wr_dat[27]), .Z(n153));
Q_MX02 U226 ( .S(n312), .A0(n153), .A1(sw_rdat[27]), .Z(n154));
Q_AN02 U227 ( .A0(n311), .A1(wr_dat[28]), .Z(n155));
Q_MX02 U228 ( .S(n312), .A0(n155), .A1(sw_rdat[28]), .Z(n156));
Q_AN02 U229 ( .A0(n311), .A1(wr_dat[29]), .Z(n157));
Q_MX02 U230 ( .S(n312), .A0(n157), .A1(sw_rdat[29]), .Z(n158));
Q_AN02 U231 ( .A0(n311), .A1(wr_dat[30]), .Z(n159));
Q_MX02 U232 ( .S(n312), .A0(n159), .A1(sw_rdat[30]), .Z(n160));
Q_AN02 U233 ( .A0(n311), .A1(wr_dat[31]), .Z(n161));
Q_MX02 U234 ( .S(n312), .A0(n161), .A1(sw_rdat[31]), .Z(n162));
Q_FDP1 \state_r_REG[3] ( .CK(clk), .R(rst_n), .D(n325), .Q(state_r[3]), .QN(n179));
Q_FDP1 \state_r_REG[2] ( .CK(clk), .R(rst_n), .D(n324), .Q(state_r[2]), .QN(n287));
Q_FDP1 \state_r_REG[1] ( .CK(clk), .R(rst_n), .D(n323), .Q(state_r[1]), .QN(n195));
Q_FDP2 \state_r_REG[0] ( .CK(clk), .S(rst_n), .D(n322), .Q(state_r[0]), .QN(n184));
Q_FDP1 \timer_r_REG[0] ( .CK(clk), .R(rst_n), .D(n92), .Q(timer_r[0]), .QN(n53));
Q_ND02 U240 ( .A0(n164), .A1(n165), .Z(n163));
Q_ND02 U241 ( .A0(n166), .A1(n270), .Z(n165));
Q_OR02 U242 ( .A0(n167), .A1(n314), .Z(n166));
Q_INV U243 ( .A(n313), .Z(n167));
Q_ND02 U244 ( .A0(n164), .A1(n169), .Z(n168));
Q_ND02 U245 ( .A0(n313), .A1(n270), .Z(n169));
Q_OR03 U246 ( .A0(n313), .A1(n314), .A2(n270), .Z(n164));
Q_MX02 U247 ( .S(n270), .A0(n313), .A1(n314), .Z(n170));
Q_FDP1 sw_cs_r_REG  ( .CK(clk), .R(rst_n), .D(n308), .Q(sw_cs_r), .QN( ));
Q_FDP1 sw_ce_r_REG  ( .CK(clk), .R(rst_n), .D(n307), .Q(sw_ce_r), .QN( ));
Q_FDP1 rst_r_REG  ( .CK(clk), .R(rst_n), .D(n306), .Q(rst_r), .QN(n326));
Q_FDP1 rst_or_ini_r_REG  ( .CK(clk), .R(rst_n), .D(n305), .Q(rst_or_ini_r), .QN( ));
Q_FDP1 sw_we_r_REG  ( .CK(clk), .R(rst_n), .D(n302), .Q(sw_we_r), .QN( ));
Q_OA21 U253 ( .A0(n172), .A1(n173), .B0(n171), .Z(n298));
Q_OR03 U254 ( .A0(n175), .A1(n176), .A2(n174), .Z(n173));
Q_AN03 U255 ( .A0(n179), .A1(n180), .A2(n177), .Z(n178));
Q_AN02 U256 ( .A0(n50), .A1(cmnd_rd_stb), .Z(n180));
Q_AO21 U257 ( .A0(n179), .A1(n181), .B0(n178), .Z(n176));
Q_AN02 U258 ( .A0(n182), .A1(n183), .Z(n181));
Q_NR02 U259 ( .A0(state_r[0]), .A1(cmnd_ena_stb), .Z(n183));
Q_OA21 U260 ( .A0(n186), .A1(n187), .B0(n185), .Z(n175));
Q_AN03 U261 ( .A0(state_r[3]), .A1(n189), .A2(n188), .Z(n187));
Q_OA21 U262 ( .A0(n191), .A1(n192), .B0(n190), .Z(n186));
Q_NR02 U263 ( .A0(n196), .A1(igrant), .Z(n192));
Q_AN02 U264 ( .A0(n193), .A1(n194), .Z(n191));
Q_INV U265 ( .A(n321), .Z(n194));
Q_NR02 U266 ( .A0(state_r[1]), .A1(state_r[0]), .Z(n193));
Q_AN03 U267 ( .A0(n200), .A1(n48), .A2(n198), .Z(n199));
Q_AN02 U268 ( .A0(cmnd_rst_stb), .A1(n179), .Z(n200));
Q_OR03 U269 ( .A0(n201), .A1(n199), .A2(n197), .Z(n172));
Q_AN03 U270 ( .A0(n202), .A1(n203), .A2(n188), .Z(n201));
Q_INV U271 ( .A(n204), .Z(n299));
Q_OA21 U272 ( .A0(n205), .A1(n174), .B0(n171), .Z(n204));
Q_AO21 U273 ( .A0(n177), .A1(n207), .B0(n206), .Z(n205));
Q_AN02 U274 ( .A0(n179), .A1(cmnd_wr_stb), .Z(n207));
Q_AN02 U275 ( .A0(n209), .A1(n210), .Z(n211));
Q_NR02 U276 ( .A0(state_r[3]), .A1(n290), .Z(n210));
Q_MX02 U277 ( .S(state_r[1]), .A0(cmnd_ena_stb), .A1(n213), .Z(n209));
Q_OR03 U278 ( .A0(n214), .A1(n211), .A2(n208), .Z(n174));
Q_AN02 U279 ( .A0(n53), .A1(n47), .Z(n185));
Q_AN03 U280 ( .A0(n216), .A1(n217), .A2(n215), .Z(n214));
Q_NR02 U281 ( .A0(cmnd_dis_stb), .A1(unsupported_op), .Z(n217));
Q_OA21 U282 ( .A0(n218), .A1(n219), .B0(n185), .Z(n208));
Q_OA21 U283 ( .A0(n220), .A1(n221), .B0(state_r[3]), .Z(n219));
Q_AN02 U284 ( .A0(state_r[2]), .A1(n213), .Z(n221));
Q_AN02 U285 ( .A0(n190), .A1(igrant), .Z(n223));
Q_AN02 U286 ( .A0(n179), .A1(state_r[2]), .Z(n190));
Q_AO21 U287 ( .A0(n224), .A1(n196), .B0(n222), .Z(n218));
Q_OA21 U288 ( .A0(state_r[0]), .A1(n225), .B0(n223), .Z(n222));
Q_AN02 U289 ( .A0(n195), .A1(n321), .Z(n225));
Q_OR02 U290 ( .A0(n179), .A1(n213), .Z(n224));
Q_AN02 U291 ( .A0(ack_error), .A1(enable), .Z(n213));
Q_OA21 U292 ( .A0(n226), .A1(n227), .B0(n182), .Z(n206));
Q_AN02 U293 ( .A0(n229), .A1(n48), .Z(n228));
Q_AN03 U294 ( .A0(n230), .A1(n231), .A2(n228), .Z(n227));
Q_AN02 U295 ( .A0(n179), .A1(state_r[0]), .Z(n230));
Q_AN02 U296 ( .A0(n232), .A1(n233), .Z(n226));
Q_AN03 U297 ( .A0(n235), .A1(n236), .A2(n234), .Z(n300));
Q_AO21 U298 ( .A0(n229), .A1(n238), .B0(n237), .Z(n234));
Q_INV U299 ( .A(n237), .Z(n238));
Q_INV U300 ( .A(n239), .Z(n301));
Q_OA21 U301 ( .A0(n240), .A1(n197), .B0(n171), .Z(n239));
Q_AN03 U302 ( .A0(n237), .A1(n179), .A2(n236), .Z(n241));
Q_AN02 U303 ( .A0(n177), .A1(n50), .Z(n236));
Q_AO21 U304 ( .A0(n51), .A1(cmnd_cmp_stb), .B0(cmnd_rd_stb), .Z(n237));
Q_AN03 U305 ( .A0(n229), .A1(n243), .A2(n198), .Z(n242));
Q_NR02 U306 ( .A0(state_r[3]), .A1(cmnd_cmp_stb), .Z(n243));
Q_AO21 U307 ( .A0(n49), .A1(n320), .B0(cmnd_rst_stb), .Z(n229));
Q_AN02 U308 ( .A0(n232), .A1(n47), .Z(n245));
Q_AN03 U309 ( .A0(n202), .A1(n182), .A2(n245), .Z(n246));
Q_OR03 U310 ( .A0(n246), .A1(n244), .A2(n241), .Z(n240));
Q_AO21 U311 ( .A0(n247), .A1(n248), .B0(n242), .Z(n244));
Q_AN02 U312 ( .A0(igrant), .A1(n47), .Z(n203));
Q_AN02 U313 ( .A0(n249), .A1(n203), .Z(n247));
Q_AN02 U314 ( .A0(n250), .A1(n184), .Z(n248));
Q_NR02 U315 ( .A0(timeout), .A1(state_r[3]), .Z(n250));
Q_AN02 U316 ( .A0(ack_error), .A1(init_r), .Z(n252));
Q_AO21 U317 ( .A0(n215), .A1(n253), .B0(n251), .Z(n197));
Q_AN02 U318 ( .A0(n216), .A1(cmnd_dis_stb), .Z(n253));
Q_NR02 U319 ( .A0(cmnd_cmp_stb), .A1(n320), .Z(n216));
Q_AN02 U320 ( .A0(n254), .A1(n198), .Z(n215));
Q_AN02 U321 ( .A0(n177), .A1(n231), .Z(n198));
Q_NR02 U322 ( .A0(cmnd_wr_stb), .A1(cmnd_rd_stb), .Z(n231));
Q_NR02 U323 ( .A0(cmnd_rst_stb), .A1(state_r[3]), .Z(n254));
Q_OA21 U324 ( .A0(n255), .A1(n256), .B0(n252), .Z(n251));
Q_AN02 U325 ( .A0(n202), .A1(n47), .Z(n233));
Q_AN02 U326 ( .A0(n53), .A1(state_r[3]), .Z(n202));
Q_OA21 U327 ( .A0(state_r[2]), .A1(n196), .B0(n233), .Z(n255));
Q_AN02 U328 ( .A0(state_r[1]), .A1(state_r[0]), .Z(n196));
Q_AO21 U329 ( .A0(n184), .A1(igrant), .B0(state_r[0]), .Z(n232));
Q_AN03 U330 ( .A0(n189), .A1(n308), .A2(n53), .Z(n92));
Q_INV U331 ( .A(igrant), .Z(n189));
Q_OA21 U332 ( .A0(n258), .A1(n259), .B0(n257), .Z(n302));
Q_AN02 U333 ( .A0(cmnd_sis_stb), .A1(n260), .Z(n303));
Q_INV U334 ( .A(n304), .Z(n260));
Q_OA21 U335 ( .A0(n258), .A1(n261), .B0(n257), .Z(n305));
Q_AN02 U336 ( .A0(n259), .A1(n262), .Z(n261));
Q_AN02 U337 ( .A0(n324), .A1(n263), .Z(n259));
Q_AN02 U338 ( .A0(n257), .A1(n258), .Z(n306));
Q_AN02 U339 ( .A0(n264), .A1(n322), .Z(n258));
Q_OR03 U340 ( .A0(n306), .A1(n265), .A2(n307), .Z(n308));
Q_AN02 U341 ( .A0(n325), .A1(n266), .Z(n307));
Q_AN03 U342 ( .A0(n257), .A1(n324), .A2(n267), .Z(n265));
Q_INV U343 ( .A(n268), .Z(n267));
Q_INV U344 ( .A(n269), .Z(n309));
Q_AN02 U345 ( .A0(n249), .A1(n230), .Z(n312));
Q_AN02 U346 ( .A0(state_r[2]), .A1(state_r[1]), .Z(n249));
Q_AN02 U347 ( .A0(n272), .A1(n273), .Z(n274));
Q_INV U348 ( .A(n275), .Z(n272));
Q_OR03 U349 ( .A0(n276), .A1(n274), .A2(n271), .Z(n270));
Q_AN03 U350 ( .A0(n278), .A1(n46), .A2(n277), .Z(n271));
Q_OR02 U351 ( .A0(n268), .A1(n279), .Z(n276));
Q_AN02 U352 ( .A0(n323), .A1(n322), .Z(n268));
Q_INV U353 ( .A(n280), .Z(n279));
Q_AN02 U354 ( .A0(n257), .A1(n281), .Z(n273));
Q_NR02 U355 ( .A0(n324), .A1(n322), .Z(n281));
Q_OA21 U356 ( .A0(n283), .A1(n263), .B0(n273), .Z(n313));
Q_AN02 U357 ( .A0(n46), .A1(n323), .Z(n275));
Q_OA21 U358 ( .A0(n278), .A1(badaddr), .B0(n275), .Z(n283));
Q_AN02 U359 ( .A0(timeout), .A1(n171), .Z(n278));
Q_NR02 U360 ( .A0(n325), .A1(n324), .Z(n280));
Q_OA21 U361 ( .A0(n284), .A1(n263), .B0(n280), .Z(n314));
Q_AN03 U362 ( .A0(n323), .A1(n262), .A2(unsupported_op), .Z(n284));
Q_ND02 U363 ( .A0(n256), .A1(n277), .Z(n285));
Q_AN02 U364 ( .A0(n264), .A1(n286), .Z(n277));
Q_NR02 U365 ( .A0(n325), .A1(n322), .Z(n286));
Q_AN02 U366 ( .A0(n282), .A1(n323), .Z(n264));
Q_AN02 U367 ( .A0(n179), .A1(n220), .Z(n256));
Q_AN03 U368 ( .A0(n287), .A1(state_r[1]), .A2(n184), .Z(n220));
Q_OA21 U369 ( .A0(n311), .A1(n288), .B0(n171), .Z(n315));
Q_AN02 U370 ( .A0(n289), .A1(state_r[1]), .Z(n288));
Q_INV U371 ( .A(n310), .Z(n311));
Q_AN02 U372 ( .A0(n182), .A1(n184), .Z(n188));
Q_MX02 U373 ( .S(state_r[3]), .A0(n291), .A1(n212), .Z(n289));
Q_INV U374 ( .A(n290), .Z(n212));
Q_AN02 U375 ( .A0(state_r[2]), .A1(state_r[0]), .Z(n291));
Q_AN03 U376 ( .A0(n310), .A1(n257), .A2(n266), .Z(n292));
Q_AN02 U377 ( .A0(n293), .A1(n262), .Z(n266));
Q_INV U378 ( .A(n322), .Z(n262));
Q_NR02 U379 ( .A0(n324), .A1(n323), .Z(n293));
Q_INV U380 ( .A(n323), .Z(n263));
Q_INV U381 ( .A(n324), .Z(n282));
Q_INV U382 ( .A(n325), .Z(n257));
Q_AO21 U383 ( .A0(n235), .A1(n294), .B0(n292), .Z(n316));
Q_AN03 U384 ( .A0(n184), .A1(cmnd_ena_stb), .A2(n182), .Z(n294));
Q_OR03 U385 ( .A0(state_r[3]), .A1(state_r[1]), .A2(n290), .Z(n310));
Q_OR02 U386 ( .A0(state_r[2]), .A1(state_r[0]), .Z(n290));
Q_AN03 U387 ( .A0(n235), .A1(n195), .A2(n295), .Z(n317));
Q_AO21 U388 ( .A0(state_r[2]), .A1(n184), .B0(n269), .Z(n295));
Q_AN02 U389 ( .A0(n287), .A1(state_r[0]), .Z(n269));
Q_ND02 U390 ( .A0(n235), .A1(n177), .Z(n318));
Q_AN02 U391 ( .A0(n182), .A1(state_r[0]), .Z(n177));
Q_NR02 U392 ( .A0(state_r[2]), .A1(state_r[1]), .Z(n182));
Q_AN02 U393 ( .A0(n235), .A1(n184), .Z(n296));
Q_AN03 U394 ( .A0(state_r[2]), .A1(n195), .A2(n296), .Z(n304));
Q_NR02 U395 ( .A0(badaddr), .A1(state_r[3]), .Z(n235));
Q_INV U396 ( .A(badaddr), .Z(n171));
Q_OR03 U397 ( .A0(cmnd_rst_stb), .A1(cmnd_sis_stb), .A2(n304), .Z(n319));
Q_OR02 U398 ( .A0(cmnd_tmo_stb), .A1(timeout), .Z(n297));
Q_AN02 U399 ( .A0(n326), .A1(wr_dat[0]), .Z(sw_wdat[0]));
Q_AN02 U400 ( .A0(n326), .A1(wr_dat[1]), .Z(sw_wdat[1]));
Q_AN02 U401 ( .A0(n326), .A1(wr_dat[2]), .Z(sw_wdat[2]));
Q_AN02 U402 ( .A0(n326), .A1(wr_dat[3]), .Z(sw_wdat[3]));
Q_AN02 U403 ( .A0(n326), .A1(wr_dat[4]), .Z(sw_wdat[4]));
Q_AN02 U404 ( .A0(n326), .A1(wr_dat[5]), .Z(sw_wdat[5]));
Q_AN02 U405 ( .A0(n326), .A1(wr_dat[6]), .Z(sw_wdat[6]));
Q_AN02 U406 ( .A0(n326), .A1(wr_dat[7]), .Z(sw_wdat[7]));
Q_AN02 U407 ( .A0(n326), .A1(wr_dat[8]), .Z(sw_wdat[8]));
Q_AN02 U408 ( .A0(n326), .A1(wr_dat[9]), .Z(sw_wdat[9]));
Q_AN02 U409 ( .A0(n326), .A1(wr_dat[10]), .Z(sw_wdat[10]));
Q_AN02 U410 ( .A0(n326), .A1(wr_dat[11]), .Z(sw_wdat[11]));
Q_AN02 U411 ( .A0(n326), .A1(wr_dat[12]), .Z(sw_wdat[12]));
Q_AN02 U412 ( .A0(n326), .A1(wr_dat[13]), .Z(sw_wdat[13]));
Q_AN02 U413 ( .A0(n326), .A1(wr_dat[14]), .Z(sw_wdat[14]));
Q_AN02 U414 ( .A0(n326), .A1(wr_dat[15]), .Z(sw_wdat[15]));
Q_AN02 U415 ( .A0(n326), .A1(wr_dat[16]), .Z(sw_wdat[16]));
Q_AN02 U416 ( .A0(n326), .A1(wr_dat[17]), .Z(sw_wdat[17]));
Q_AN02 U417 ( .A0(n326), .A1(wr_dat[18]), .Z(sw_wdat[18]));
Q_AN02 U418 ( .A0(n326), .A1(wr_dat[19]), .Z(sw_wdat[19]));
Q_AN02 U419 ( .A0(n326), .A1(wr_dat[20]), .Z(sw_wdat[20]));
Q_AN02 U420 ( .A0(n326), .A1(wr_dat[21]), .Z(sw_wdat[21]));
Q_AN02 U421 ( .A0(n326), .A1(wr_dat[22]), .Z(sw_wdat[22]));
Q_AN02 U422 ( .A0(n326), .A1(wr_dat[23]), .Z(sw_wdat[23]));
Q_AN02 U423 ( .A0(n326), .A1(wr_dat[24]), .Z(sw_wdat[24]));
Q_AN02 U424 ( .A0(n326), .A1(wr_dat[25]), .Z(sw_wdat[25]));
Q_AN02 U425 ( .A0(n326), .A1(wr_dat[26]), .Z(sw_wdat[26]));
Q_AN02 U426 ( .A0(n326), .A1(wr_dat[27]), .Z(sw_wdat[27]));
Q_AN02 U427 ( .A0(n326), .A1(wr_dat[28]), .Z(sw_wdat[28]));
Q_AN02 U428 ( .A0(n326), .A1(wr_dat[29]), .Z(sw_wdat[29]));
Q_AN02 U429 ( .A0(n326), .A1(wr_dat[30]), .Z(sw_wdat[30]));
Q_AN02 U430 ( .A0(n326), .A1(wr_dat[31]), .Z(sw_wdat[31]));
Q_FDP4EP sim_tmo_r_REG  ( .CK(clk), .CE(n297), .R(n327), .D(cmnd_tmo_stb), .Q(sim_tmo_r));
Q_INV U432 ( .A(rst_n), .Z(n327));
Q_INV U433 ( .A(sim_tmo_r), .Z(n19));
Q_FDP4EP init_r_REG  ( .CK(clk), .CE(n316), .R(n327), .D(n310), .Q(init_r));
Q_INV U435 ( .A(init_r), .Z(enable));
Q_FDP4EP \stat_code_REG[0] ( .CK(clk), .CE(n285), .R(n327), .D(n163), .Q(stat_code[0]));
Q_FDP4EP \stat_code_REG[1] ( .CK(clk), .CE(n285), .R(n327), .D(n168), .Q(stat_code[1]));
Q_FDP4EP \stat_code_REG[2] ( .CK(clk), .CE(n285), .R(n327), .D(n170), .Q(stat_code[2]));
Q_FDP4EP \rst_addr_r_REG[0] ( .CK(clk), .CE(n319), .R(n327), .D(n94), .Q(rst_addr_r[0]));
Q_FDP4EP \rst_addr_r_REG[1] ( .CK(clk), .CE(n319), .R(n327), .D(n96), .Q(rst_addr_r[1]));
Q_FDP4EP \rst_addr_r_REG[2] ( .CK(clk), .CE(n319), .R(n327), .D(n98), .Q(rst_addr_r[2]));
Q_FDP4EP \rst_addr_r_REG[3] ( .CK(clk), .CE(n319), .R(n327), .D(n100), .Q(rst_addr_r[3]));
Q_FDP4EP \rst_addr_r_REG[4] ( .CK(clk), .CE(n319), .R(n327), .D(n102), .Q(rst_addr_r[4]));
Q_FDP4EP \inc_r_REG[0] ( .CK(clk), .CE(n317), .R(n327), .D(n103), .Q(inc_r[0]));
Q_FDP4EP \rd_dat_REG[0] ( .CK(clk), .CE(n315), .R(n327), .D(n104), .Q(rd_dat[0]));
Q_FDP4EP \rd_dat_REG[1] ( .CK(clk), .CE(n315), .R(n327), .D(n105), .Q(rd_dat[1]));
Q_FDP4EP \rd_dat_REG[2] ( .CK(clk), .CE(n315), .R(n327), .D(n106), .Q(rd_dat[2]));
Q_FDP4EP \rd_dat_REG[3] ( .CK(clk), .CE(n315), .R(n327), .D(n107), .Q(rd_dat[3]));
Q_FDP4EP \rd_dat_REG[4] ( .CK(clk), .CE(n315), .R(n327), .D(n108), .Q(rd_dat[4]));
Q_FDP4EP \rd_dat_REG[5] ( .CK(clk), .CE(n315), .R(n327), .D(n110), .Q(rd_dat[5]));
Q_FDP4EP \rd_dat_REG[6] ( .CK(clk), .CE(n315), .R(n327), .D(n112), .Q(rd_dat[6]));
Q_FDP4EP \rd_dat_REG[7] ( .CK(clk), .CE(n315), .R(n327), .D(n114), .Q(rd_dat[7]));
Q_FDP4EP \rd_dat_REG[8] ( .CK(clk), .CE(n315), .R(n327), .D(n116), .Q(rd_dat[8]));
Q_FDP4EP \rd_dat_REG[9] ( .CK(clk), .CE(n315), .R(n327), .D(n118), .Q(rd_dat[9]));
Q_FDP4EP \rd_dat_REG[10] ( .CK(clk), .CE(n315), .R(n327), .D(n120), .Q(rd_dat[10]));
Q_FDP4EP \rd_dat_REG[11] ( .CK(clk), .CE(n315), .R(n327), .D(n122), .Q(rd_dat[11]));
Q_FDP4EP \rd_dat_REG[12] ( .CK(clk), .CE(n315), .R(n327), .D(n124), .Q(rd_dat[12]));
Q_FDP4EP \rd_dat_REG[13] ( .CK(clk), .CE(n315), .R(n327), .D(n126), .Q(rd_dat[13]));
Q_FDP4EP \rd_dat_REG[14] ( .CK(clk), .CE(n315), .R(n327), .D(n128), .Q(rd_dat[14]));
Q_FDP4EP \rd_dat_REG[15] ( .CK(clk), .CE(n315), .R(n327), .D(n130), .Q(rd_dat[15]));
Q_FDP4EP \rd_dat_REG[16] ( .CK(clk), .CE(n315), .R(n327), .D(n132), .Q(rd_dat[16]));
Q_FDP4EP \rd_dat_REG[17] ( .CK(clk), .CE(n315), .R(n327), .D(n134), .Q(rd_dat[17]));
Q_FDP4EP \rd_dat_REG[18] ( .CK(clk), .CE(n315), .R(n327), .D(n136), .Q(rd_dat[18]));
Q_FDP4EP \rd_dat_REG[19] ( .CK(clk), .CE(n315), .R(n327), .D(n138), .Q(rd_dat[19]));
Q_FDP4EP \rd_dat_REG[20] ( .CK(clk), .CE(n315), .R(n327), .D(n140), .Q(rd_dat[20]));
Q_FDP4EP \rd_dat_REG[21] ( .CK(clk), .CE(n315), .R(n327), .D(n142), .Q(rd_dat[21]));
Q_FDP4EP \rd_dat_REG[22] ( .CK(clk), .CE(n315), .R(n327), .D(n144), .Q(rd_dat[22]));
Q_FDP4EP \rd_dat_REG[23] ( .CK(clk), .CE(n315), .R(n327), .D(n146), .Q(rd_dat[23]));
Q_FDP4EP \rd_dat_REG[24] ( .CK(clk), .CE(n315), .R(n327), .D(n148), .Q(rd_dat[24]));
Q_FDP4EP \rd_dat_REG[25] ( .CK(clk), .CE(n315), .R(n327), .D(n150), .Q(rd_dat[25]));
Q_FDP4EP \rd_dat_REG[26] ( .CK(clk), .CE(n315), .R(n327), .D(n152), .Q(rd_dat[26]));
Q_FDP4EP \rd_dat_REG[27] ( .CK(clk), .CE(n315), .R(n327), .D(n154), .Q(rd_dat[27]));
Q_FDP4EP \rd_dat_REG[28] ( .CK(clk), .CE(n315), .R(n327), .D(n156), .Q(rd_dat[28]));
Q_FDP4EP \rd_dat_REG[29] ( .CK(clk), .CE(n315), .R(n327), .D(n158), .Q(rd_dat[29]));
Q_FDP4EP \rd_dat_REG[30] ( .CK(clk), .CE(n315), .R(n327), .D(n160), .Q(rd_dat[30]));
Q_FDP4EP \rd_dat_REG[31] ( .CK(clk), .CE(n315), .R(n327), .D(n162), .Q(rd_dat[31]));
Q_INV U477 ( .A(n318), .Z(n328));
Q_FDP4EP init_inc_r_REG  ( .CK(clk), .CE(n328), .R(n327), .D(n1), .Q(init_inc_r));
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "addr_limit (2,0) 1 4 0 0 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "1"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_1 "-1 genblk2  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_0 "-1 genblk1  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "genblk2"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "genblk1"
endmodule
