
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module cr_kme_kop_keybuilder ( tlv_sb_data_out_ack, keybuilder_kdf_stall, 
	gcm_status_data_out_ack, key_tlv_ob_wr, .key_tlv_ob_tlv( {
	\key_tlv_ob_tlv.insert , \key_tlv_ob_tlv.ordern [12], 
	\key_tlv_ob_tlv.ordern [11], \key_tlv_ob_tlv.ordern [10], 
	\key_tlv_ob_tlv.ordern [9], \key_tlv_ob_tlv.ordern [8], 
	\key_tlv_ob_tlv.ordern [7], \key_tlv_ob_tlv.ordern [6], 
	\key_tlv_ob_tlv.ordern [5], \key_tlv_ob_tlv.ordern [4], 
	\key_tlv_ob_tlv.ordern [3], \key_tlv_ob_tlv.ordern [2], 
	\key_tlv_ob_tlv.ordern [1], \key_tlv_ob_tlv.ordern [0], 
	\key_tlv_ob_tlv.typen [7], \key_tlv_ob_tlv.typen [6], 
	\key_tlv_ob_tlv.typen [5], \key_tlv_ob_tlv.typen [4], 
	\key_tlv_ob_tlv.typen [3], \key_tlv_ob_tlv.typen [2], 
	\key_tlv_ob_tlv.typen [1], \key_tlv_ob_tlv.typen [0], 
	\key_tlv_ob_tlv.sot , \key_tlv_ob_tlv.eot , \key_tlv_ob_tlv.tlast , 
	\key_tlv_ob_tlv.tid [0], \key_tlv_ob_tlv.tstrb [7], 
	\key_tlv_ob_tlv.tstrb [6], \key_tlv_ob_tlv.tstrb [5], 
	\key_tlv_ob_tlv.tstrb [4], \key_tlv_ob_tlv.tstrb [3], 
	\key_tlv_ob_tlv.tstrb [2], \key_tlv_ob_tlv.tstrb [1], 
	\key_tlv_ob_tlv.tstrb [0], \key_tlv_ob_tlv.tuser [7], 
	\key_tlv_ob_tlv.tuser [6], \key_tlv_ob_tlv.tuser [5], 
	\key_tlv_ob_tlv.tuser [4], \key_tlv_ob_tlv.tuser [3], 
	\key_tlv_ob_tlv.tuser [2], \key_tlv_ob_tlv.tuser [1], 
	\key_tlv_ob_tlv.tuser [0], \key_tlv_ob_tlv.tdata [63], 
	\key_tlv_ob_tlv.tdata [62], \key_tlv_ob_tlv.tdata [61], 
	\key_tlv_ob_tlv.tdata [60], \key_tlv_ob_tlv.tdata [59], 
	\key_tlv_ob_tlv.tdata [58], \key_tlv_ob_tlv.tdata [57], 
	\key_tlv_ob_tlv.tdata [56], \key_tlv_ob_tlv.tdata [55], 
	\key_tlv_ob_tlv.tdata [54], \key_tlv_ob_tlv.tdata [53], 
	\key_tlv_ob_tlv.tdata [52], \key_tlv_ob_tlv.tdata [51], 
	\key_tlv_ob_tlv.tdata [50], \key_tlv_ob_tlv.tdata [49], 
	\key_tlv_ob_tlv.tdata [48], \key_tlv_ob_tlv.tdata [47], 
	\key_tlv_ob_tlv.tdata [46], \key_tlv_ob_tlv.tdata [45], 
	\key_tlv_ob_tlv.tdata [44], \key_tlv_ob_tlv.tdata [43], 
	\key_tlv_ob_tlv.tdata [42], \key_tlv_ob_tlv.tdata [41], 
	\key_tlv_ob_tlv.tdata [40], \key_tlv_ob_tlv.tdata [39], 
	\key_tlv_ob_tlv.tdata [38], \key_tlv_ob_tlv.tdata [37], 
	\key_tlv_ob_tlv.tdata [36], \key_tlv_ob_tlv.tdata [35], 
	\key_tlv_ob_tlv.tdata [34], \key_tlv_ob_tlv.tdata [33], 
	\key_tlv_ob_tlv.tdata [32], \key_tlv_ob_tlv.tdata [31], 
	\key_tlv_ob_tlv.tdata [30], \key_tlv_ob_tlv.tdata [29], 
	\key_tlv_ob_tlv.tdata [28], \key_tlv_ob_tlv.tdata [27], 
	\key_tlv_ob_tlv.tdata [26], \key_tlv_ob_tlv.tdata [25], 
	\key_tlv_ob_tlv.tdata [24], \key_tlv_ob_tlv.tdata [23], 
	\key_tlv_ob_tlv.tdata [22], \key_tlv_ob_tlv.tdata [21], 
	\key_tlv_ob_tlv.tdata [20], \key_tlv_ob_tlv.tdata [19], 
	\key_tlv_ob_tlv.tdata [18], \key_tlv_ob_tlv.tdata [17], 
	\key_tlv_ob_tlv.tdata [16], \key_tlv_ob_tlv.tdata [15], 
	\key_tlv_ob_tlv.tdata [14], \key_tlv_ob_tlv.tdata [13], 
	\key_tlv_ob_tlv.tdata [12], \key_tlv_ob_tlv.tdata [11], 
	\key_tlv_ob_tlv.tdata [10], \key_tlv_ob_tlv.tdata [9], 
	\key_tlv_ob_tlv.tdata [8], \key_tlv_ob_tlv.tdata [7], 
	\key_tlv_ob_tlv.tdata [6], \key_tlv_ob_tlv.tdata [5], 
	\key_tlv_ob_tlv.tdata [4], \key_tlv_ob_tlv.tdata [3], 
	\key_tlv_ob_tlv.tdata [2], \key_tlv_ob_tlv.tdata [1], 
	\key_tlv_ob_tlv.tdata [0]} ), clk, rst_n, tlv_sb_data_out, 
	tlv_sb_data_out_valid, kdf_keybuilder_data, kdf_keybuilder_valid, 
	gcm_status_data_out_valid, .gcm_status_data_out( {
	\gcm_status_data_out.tag_mismatch [0]} ), key_tlv_ob_full, 
	key_tlv_ob_afull);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output tlv_sb_data_out_ack;
output keybuilder_kdf_stall;
output gcm_status_data_out_ack;
output key_tlv_ob_wr;
output \key_tlv_ob_tlv.insert ;
output [12:0] \key_tlv_ob_tlv.ordern ;
output [7:0] \key_tlv_ob_tlv.typen ;
output \key_tlv_ob_tlv.sot ;
output \key_tlv_ob_tlv.eot ;
output \key_tlv_ob_tlv.tlast ;
output [0:0] \key_tlv_ob_tlv.tid ;
output [7:0] \key_tlv_ob_tlv.tstrb ;
output [7:0] \key_tlv_ob_tlv.tuser ;
output [63:0] \key_tlv_ob_tlv.tdata ;
wire [105:0] key_tlv_ob_tlv;
input clk;
input rst_n;
input [63:0] tlv_sb_data_out;
input tlv_sb_data_out_valid;
input [63:0] kdf_keybuilder_data;
input kdf_keybuilder_valid;
input gcm_status_data_out_valid;
input [0:0] \gcm_status_data_out.tag_mismatch ;
wire [0:0] gcm_status_data_out;
input key_tlv_ob_full;
input key_tlv_ob_afull;
wire init;
wire data_valid;
wire [31:0] crc;
wire _zy_simnet_tlv_sb_data_out_ack_0_w$;
wire _zy_simnet_keybuilder_kdf_stall_1_w$;
wire _zy_simnet_gcm_status_data_out_ack_2_w$;
wire _zy_simnet_key_tlv_ob_wr_3_w$;
wire [0:105] _zy_simnet_key_tlv_ob_tlv_4_w$;
wire [0:63] _zy_simnet_key_tlv_ob_tlv_5_w$;
wire [0:7] _zy_simnet_cio_6;
wire _zy_simnet_cio_7;
wire [0:31] _zy_simnet_cio_8;
wire [63:0] key_tlv_word0;
wire [63:0] key_tlv_word19;
wire [63:0] key_tlv_word20;
wire [63:0] int_tlv_word0;
wire [55:0] int_tlv_word42;
wire [2:0] key_tlv_beat_num;
wire [2:0] cur_state;
wire [2:0] nxt_state;
wire dek_gcm_err;
wire nxt_dek_gcm_err;
wire dak_gcm_err;
wire nxt_dak_gcm_err;
wire corrupt_crc;
wire nxt_corrupt_crc;
wire needs_dek;
wire nxt_needs_dek;
wire needs_dak;
wire nxt_needs_dak;
supply0 n314;
supply1 n315;
wire [1:0] \key_tlv_word0.tlv_bip2 ;
wire [18:0] \key_tlv_word0.resv0 ;
wire [10:0] \key_tlv_word0.tlv_frame_num ;
wire [3:0] \key_tlv_word0.resv1 ;
wire [3:0] \key_tlv_word0.tlv_eng_id ;
wire [7:0] \key_tlv_word0.tlv_seq_num ;
wire [7:0] \key_tlv_word0.tlv_len ;
wire [7:0] \key_tlv_word0.tlv_type ;
wire [55:0] \key_tlv_word19.rsvd ;
wire [7:0] \key_tlv_word19.kme_errors ;
wire [31:0] \key_tlv_word20.rsvd ;
wire [31:0] \key_tlv_word20.crc32 ;
wire [1:0] \int_tlv_word0.tlv_bip2 ;
wire [12:0] \int_tlv_word0.resv0 ;
wire [0:0] \int_tlv_word0.kdf_dek_iter ;
wire [0:0] \int_tlv_word0.keyless_algos ;
wire [0:0] \int_tlv_word0.needs_dek ;
wire [0:0] \int_tlv_word0.needs_dak ;
wire [5:0] \int_tlv_word0.key_type ;
wire [10:0] \int_tlv_word0.tlv_frame_num ;
wire [3:0] \int_tlv_word0.tlv_eng_id ;
wire [7:0] \int_tlv_word0.tlv_seq_num ;
wire [7:0] \int_tlv_word0.tlv_len ;
wire [7:0] \int_tlv_word0.tlv_type ;
wire [0:0] \int_tlv_word42.corrupt_crc32 ;
wire [46:0] \int_tlv_word42.unused ;
wire [7:0] \int_tlv_word42.error_code ;
tran (key_tlv_ob_tlv[105], \key_tlv_ob_tlv.insert );
tran (key_tlv_ob_tlv[104], \key_tlv_ob_tlv.ordern [12]);
tran (key_tlv_ob_tlv[103], \key_tlv_ob_tlv.ordern [11]);
tran (key_tlv_ob_tlv[102], \key_tlv_ob_tlv.ordern [10]);
tran (key_tlv_ob_tlv[101], \key_tlv_ob_tlv.ordern [9]);
tran (key_tlv_ob_tlv[100], \key_tlv_ob_tlv.ordern [8]);
tran (key_tlv_ob_tlv[99], \key_tlv_ob_tlv.ordern [7]);
tran (key_tlv_ob_tlv[98], \key_tlv_ob_tlv.ordern [6]);
tran (key_tlv_ob_tlv[97], \key_tlv_ob_tlv.ordern [5]);
tran (key_tlv_ob_tlv[96], \key_tlv_ob_tlv.ordern [4]);
tran (key_tlv_ob_tlv[95], \key_tlv_ob_tlv.ordern [3]);
tran (key_tlv_ob_tlv[94], \key_tlv_ob_tlv.ordern [2]);
tran (key_tlv_ob_tlv[93], \key_tlv_ob_tlv.ordern [1]);
tran (key_tlv_ob_tlv[92], \key_tlv_ob_tlv.ordern [0]);
tran (key_tlv_ob_tlv[91], \key_tlv_ob_tlv.typen [7]);
tran (key_tlv_ob_tlv[90], \key_tlv_ob_tlv.typen [6]);
tran (key_tlv_ob_tlv[89], \key_tlv_ob_tlv.typen [5]);
tran (key_tlv_ob_tlv[88], \key_tlv_ob_tlv.typen [4]);
tran (key_tlv_ob_tlv[87], \key_tlv_ob_tlv.typen [3]);
tran (key_tlv_ob_tlv[86], \key_tlv_ob_tlv.typen [2]);
tran (key_tlv_ob_tlv[85], \key_tlv_ob_tlv.typen [1]);
tran (key_tlv_ob_tlv[84], \key_tlv_ob_tlv.typen [0]);
tran (key_tlv_ob_tlv[83], \key_tlv_ob_tlv.sot );
tran (key_tlv_ob_tlv[82], \key_tlv_ob_tlv.eot );
tran (key_tlv_ob_tlv[81], \key_tlv_ob_tlv.tlast );
tran (key_tlv_ob_tlv[80], \key_tlv_ob_tlv.tid [0]);
tran (key_tlv_ob_tlv[79], \key_tlv_ob_tlv.tstrb [7]);
tran (key_tlv_ob_tlv[78], \key_tlv_ob_tlv.tstrb [6]);
tran (key_tlv_ob_tlv[77], \key_tlv_ob_tlv.tstrb [5]);
tran (key_tlv_ob_tlv[76], \key_tlv_ob_tlv.tstrb [4]);
tran (key_tlv_ob_tlv[75], \key_tlv_ob_tlv.tstrb [3]);
tran (key_tlv_ob_tlv[74], \key_tlv_ob_tlv.tstrb [2]);
tran (key_tlv_ob_tlv[73], \key_tlv_ob_tlv.tstrb [1]);
tran (key_tlv_ob_tlv[72], \key_tlv_ob_tlv.tstrb [0]);
tran (key_tlv_ob_tlv[71], \key_tlv_ob_tlv.tuser [7]);
tran (key_tlv_ob_tlv[70], \key_tlv_ob_tlv.tuser [6]);
tran (key_tlv_ob_tlv[69], \key_tlv_ob_tlv.tuser [5]);
tran (key_tlv_ob_tlv[68], \key_tlv_ob_tlv.tuser [4]);
tran (key_tlv_ob_tlv[67], \key_tlv_ob_tlv.tuser [3]);
tran (key_tlv_ob_tlv[66], \key_tlv_ob_tlv.tuser [2]);
tran (key_tlv_ob_tlv[65], \key_tlv_ob_tlv.tuser [1]);
tran (key_tlv_ob_tlv[64], \key_tlv_ob_tlv.tuser [0]);
tran (key_tlv_ob_tlv[63], \key_tlv_ob_tlv.tdata [63]);
tran (key_tlv_ob_tlv[62], \key_tlv_ob_tlv.tdata [62]);
tran (key_tlv_ob_tlv[61], \key_tlv_ob_tlv.tdata [61]);
tran (key_tlv_ob_tlv[60], \key_tlv_ob_tlv.tdata [60]);
tran (key_tlv_ob_tlv[59], \key_tlv_ob_tlv.tdata [59]);
tran (key_tlv_ob_tlv[58], \key_tlv_ob_tlv.tdata [58]);
tran (key_tlv_ob_tlv[57], \key_tlv_ob_tlv.tdata [57]);
tran (key_tlv_ob_tlv[56], \key_tlv_ob_tlv.tdata [56]);
tran (key_tlv_ob_tlv[55], \key_tlv_ob_tlv.tdata [55]);
tran (key_tlv_ob_tlv[54], \key_tlv_ob_tlv.tdata [54]);
tran (key_tlv_ob_tlv[53], \key_tlv_ob_tlv.tdata [53]);
tran (key_tlv_ob_tlv[52], \key_tlv_ob_tlv.tdata [52]);
tran (key_tlv_ob_tlv[51], \key_tlv_ob_tlv.tdata [51]);
tran (key_tlv_ob_tlv[50], \key_tlv_ob_tlv.tdata [50]);
tran (key_tlv_ob_tlv[49], \key_tlv_ob_tlv.tdata [49]);
tran (key_tlv_ob_tlv[48], \key_tlv_ob_tlv.tdata [48]);
tran (key_tlv_ob_tlv[47], \key_tlv_ob_tlv.tdata [47]);
tran (key_tlv_ob_tlv[46], \key_tlv_ob_tlv.tdata [46]);
tran (key_tlv_ob_tlv[45], \key_tlv_ob_tlv.tdata [45]);
tran (key_tlv_ob_tlv[44], \key_tlv_ob_tlv.tdata [44]);
tran (key_tlv_ob_tlv[43], \key_tlv_ob_tlv.tdata [43]);
tran (key_tlv_ob_tlv[42], \key_tlv_ob_tlv.tdata [42]);
tran (key_tlv_ob_tlv[41], \key_tlv_ob_tlv.tdata [41]);
tran (key_tlv_ob_tlv[40], \key_tlv_ob_tlv.tdata [40]);
tran (key_tlv_ob_tlv[39], \key_tlv_ob_tlv.tdata [39]);
tran (key_tlv_ob_tlv[38], \key_tlv_ob_tlv.tdata [38]);
tran (key_tlv_ob_tlv[37], \key_tlv_ob_tlv.tdata [37]);
tran (key_tlv_ob_tlv[36], \key_tlv_ob_tlv.tdata [36]);
tran (key_tlv_ob_tlv[35], \key_tlv_ob_tlv.tdata [35]);
tran (key_tlv_ob_tlv[34], \key_tlv_ob_tlv.tdata [34]);
tran (key_tlv_ob_tlv[33], \key_tlv_ob_tlv.tdata [33]);
tran (key_tlv_ob_tlv[32], \key_tlv_ob_tlv.tdata [32]);
tran (key_tlv_ob_tlv[31], \key_tlv_ob_tlv.tdata [31]);
tran (key_tlv_ob_tlv[30], \key_tlv_ob_tlv.tdata [30]);
tran (key_tlv_ob_tlv[29], \key_tlv_ob_tlv.tdata [29]);
tran (key_tlv_ob_tlv[28], \key_tlv_ob_tlv.tdata [28]);
tran (key_tlv_ob_tlv[27], \key_tlv_ob_tlv.tdata [27]);
tran (key_tlv_ob_tlv[26], \key_tlv_ob_tlv.tdata [26]);
tran (key_tlv_ob_tlv[25], \key_tlv_ob_tlv.tdata [25]);
tran (key_tlv_ob_tlv[24], \key_tlv_ob_tlv.tdata [24]);
tran (key_tlv_ob_tlv[23], \key_tlv_ob_tlv.tdata [23]);
tran (key_tlv_ob_tlv[22], \key_tlv_ob_tlv.tdata [22]);
tran (key_tlv_ob_tlv[21], \key_tlv_ob_tlv.tdata [21]);
tran (key_tlv_ob_tlv[20], \key_tlv_ob_tlv.tdata [20]);
tran (key_tlv_ob_tlv[19], \key_tlv_ob_tlv.tdata [19]);
tran (key_tlv_ob_tlv[18], \key_tlv_ob_tlv.tdata [18]);
tran (key_tlv_ob_tlv[17], \key_tlv_ob_tlv.tdata [17]);
tran (key_tlv_ob_tlv[16], \key_tlv_ob_tlv.tdata [16]);
tran (key_tlv_ob_tlv[15], \key_tlv_ob_tlv.tdata [15]);
tran (key_tlv_ob_tlv[14], \key_tlv_ob_tlv.tdata [14]);
tran (key_tlv_ob_tlv[13], \key_tlv_ob_tlv.tdata [13]);
tran (key_tlv_ob_tlv[12], \key_tlv_ob_tlv.tdata [12]);
tran (key_tlv_ob_tlv[11], \key_tlv_ob_tlv.tdata [11]);
tran (key_tlv_ob_tlv[10], \key_tlv_ob_tlv.tdata [10]);
tran (key_tlv_ob_tlv[9], \key_tlv_ob_tlv.tdata [9]);
tran (key_tlv_ob_tlv[8], \key_tlv_ob_tlv.tdata [8]);
tran (key_tlv_ob_tlv[7], \key_tlv_ob_tlv.tdata [7]);
tran (key_tlv_ob_tlv[6], \key_tlv_ob_tlv.tdata [6]);
tran (key_tlv_ob_tlv[5], \key_tlv_ob_tlv.tdata [5]);
tran (key_tlv_ob_tlv[4], \key_tlv_ob_tlv.tdata [4]);
tran (key_tlv_ob_tlv[3], \key_tlv_ob_tlv.tdata [3]);
tran (key_tlv_ob_tlv[2], \key_tlv_ob_tlv.tdata [2]);
tran (key_tlv_ob_tlv[1], \key_tlv_ob_tlv.tdata [1]);
tran (key_tlv_ob_tlv[0], \key_tlv_ob_tlv.tdata [0]);
tran (gcm_status_data_out[0], \gcm_status_data_out.tag_mismatch [0]);
tran (int_tlv_word0[63], \int_tlv_word0.tlv_bip2 [1]);
tran (int_tlv_word0[62], \int_tlv_word0.tlv_bip2 [0]);
tran (int_tlv_word0[61], \int_tlv_word0.resv0 [12]);
tran (int_tlv_word0[60], \int_tlv_word0.resv0 [11]);
tran (int_tlv_word0[59], \int_tlv_word0.resv0 [10]);
tran (int_tlv_word0[58], \int_tlv_word0.resv0 [9]);
tran (int_tlv_word0[57], \int_tlv_word0.resv0 [8]);
tran (int_tlv_word0[56], \int_tlv_word0.resv0 [7]);
tran (int_tlv_word0[55], \int_tlv_word0.resv0 [6]);
tran (int_tlv_word42[55], \int_tlv_word42.corrupt_crc32 [0]);
tran (int_tlv_word0[54], \int_tlv_word0.resv0 [5]);
tran (int_tlv_word42[54], \int_tlv_word42.unused [46]);
tran (int_tlv_word0[53], \int_tlv_word0.resv0 [4]);
tran (int_tlv_word42[53], \int_tlv_word42.unused [45]);
tran (int_tlv_word0[52], \int_tlv_word0.resv0 [3]);
tran (int_tlv_word42[52], \int_tlv_word42.unused [44]);
tran (int_tlv_word0[51], \int_tlv_word0.resv0 [2]);
tran (int_tlv_word42[51], \int_tlv_word42.unused [43]);
tran (int_tlv_word0[50], \int_tlv_word0.resv0 [1]);
tran (int_tlv_word42[50], \int_tlv_word42.unused [42]);
tran (int_tlv_word0[49], \int_tlv_word0.resv0 [0]);
tran (int_tlv_word42[49], \int_tlv_word42.unused [41]);
tran (int_tlv_word0[48], \int_tlv_word0.kdf_dek_iter [0]);
tran (int_tlv_word42[48], \int_tlv_word42.unused [40]);
tran (int_tlv_word0[47], \int_tlv_word0.keyless_algos [0]);
tran (int_tlv_word42[47], \int_tlv_word42.unused [39]);
tran (int_tlv_word0[46], \int_tlv_word0.needs_dek [0]);
tran (int_tlv_word42[46], \int_tlv_word42.unused [38]);
tran (int_tlv_word0[45], \int_tlv_word0.needs_dak [0]);
tran (int_tlv_word42[45], \int_tlv_word42.unused [37]);
tran (int_tlv_word0[44], \int_tlv_word0.key_type [5]);
tran (int_tlv_word42[44], \int_tlv_word42.unused [36]);
tran (int_tlv_word0[43], \int_tlv_word0.key_type [4]);
tran (int_tlv_word42[43], \int_tlv_word42.unused [35]);
tran (int_tlv_word0[42], \int_tlv_word0.key_type [3]);
tran (int_tlv_word42[42], \int_tlv_word42.unused [34]);
tran (int_tlv_word0[41], \int_tlv_word0.key_type [2]);
tran (int_tlv_word42[41], \int_tlv_word42.unused [33]);
tran (int_tlv_word0[40], \int_tlv_word0.key_type [1]);
tran (int_tlv_word42[40], \int_tlv_word42.unused [32]);
tran (int_tlv_word0[39], \int_tlv_word0.key_type [0]);
tran (int_tlv_word42[39], \int_tlv_word42.unused [31]);
tran (key_tlv_word0[42], \key_tlv_word0.tlv_frame_num [10]);
tran (int_tlv_word0[38], \int_tlv_word0.tlv_frame_num [10]);
tran (int_tlv_word42[38], \int_tlv_word42.unused [30]);
tran (key_tlv_word0[41], \key_tlv_word0.tlv_frame_num [9]);
tran (int_tlv_word0[37], \int_tlv_word0.tlv_frame_num [9]);
tran (int_tlv_word42[37], \int_tlv_word42.unused [29]);
tran (key_tlv_word0[40], \key_tlv_word0.tlv_frame_num [8]);
tran (int_tlv_word0[36], \int_tlv_word0.tlv_frame_num [8]);
tran (int_tlv_word42[36], \int_tlv_word42.unused [28]);
tran (key_tlv_word0[39], \key_tlv_word0.tlv_frame_num [7]);
tran (int_tlv_word0[35], \int_tlv_word0.tlv_frame_num [7]);
tran (int_tlv_word42[35], \int_tlv_word42.unused [27]);
tran (key_tlv_word0[38], \key_tlv_word0.tlv_frame_num [6]);
tran (int_tlv_word0[34], \int_tlv_word0.tlv_frame_num [6]);
tran (int_tlv_word42[34], \int_tlv_word42.unused [26]);
tran (key_tlv_word0[37], \key_tlv_word0.tlv_frame_num [5]);
tran (int_tlv_word0[33], \int_tlv_word0.tlv_frame_num [5]);
tran (int_tlv_word42[33], \int_tlv_word42.unused [25]);
tran (key_tlv_word0[36], \key_tlv_word0.tlv_frame_num [4]);
tran (int_tlv_word0[32], \int_tlv_word0.tlv_frame_num [4]);
tran (int_tlv_word42[32], \int_tlv_word42.unused [24]);
tran (key_tlv_word0[35], \key_tlv_word0.tlv_frame_num [3]);
tran (int_tlv_word0[31], \int_tlv_word0.tlv_frame_num [3]);
tran (int_tlv_word42[31], \int_tlv_word42.unused [23]);
tran (key_tlv_word0[34], \key_tlv_word0.tlv_frame_num [2]);
tran (int_tlv_word0[30], \int_tlv_word0.tlv_frame_num [2]);
tran (int_tlv_word42[30], \int_tlv_word42.unused [22]);
tran (key_tlv_word0[33], \key_tlv_word0.tlv_frame_num [1]);
tran (int_tlv_word0[29], \int_tlv_word0.tlv_frame_num [1]);
tran (int_tlv_word42[29], \int_tlv_word42.unused [21]);
tran (key_tlv_word0[32], \key_tlv_word0.tlv_frame_num [0]);
tran (int_tlv_word0[28], \int_tlv_word0.tlv_frame_num [0]);
tran (int_tlv_word42[28], \int_tlv_word42.unused [20]);
tran (key_tlv_word0[27], \key_tlv_word0.tlv_eng_id [3]);
tran (int_tlv_word0[27], \int_tlv_word0.tlv_eng_id [3]);
tran (int_tlv_word42[27], \int_tlv_word42.unused [19]);
tran (key_tlv_word0[26], \key_tlv_word0.tlv_eng_id [2]);
tran (int_tlv_word0[26], \int_tlv_word0.tlv_eng_id [2]);
tran (int_tlv_word42[26], \int_tlv_word42.unused [18]);
tran (key_tlv_word0[25], \key_tlv_word0.tlv_eng_id [1]);
tran (int_tlv_word0[25], \int_tlv_word0.tlv_eng_id [1]);
tran (int_tlv_word42[25], \int_tlv_word42.unused [17]);
tran (key_tlv_word0[24], \key_tlv_word0.tlv_eng_id [0]);
tran (int_tlv_word0[24], \int_tlv_word0.tlv_eng_id [0]);
tran (int_tlv_word42[24], \int_tlv_word42.unused [16]);
tran (key_tlv_word0[23], \key_tlv_word0.tlv_seq_num [7]);
tran (int_tlv_word0[23], \int_tlv_word0.tlv_seq_num [7]);
tran (int_tlv_word42[23], \int_tlv_word42.unused [15]);
tran (key_tlv_word0[22], \key_tlv_word0.tlv_seq_num [6]);
tran (int_tlv_word0[22], \int_tlv_word0.tlv_seq_num [6]);
tran (int_tlv_word42[22], \int_tlv_word42.unused [14]);
tran (key_tlv_word0[21], \key_tlv_word0.tlv_seq_num [5]);
tran (int_tlv_word0[21], \int_tlv_word0.tlv_seq_num [5]);
tran (int_tlv_word42[21], \int_tlv_word42.unused [13]);
tran (key_tlv_word0[20], \key_tlv_word0.tlv_seq_num [4]);
tran (int_tlv_word0[20], \int_tlv_word0.tlv_seq_num [4]);
tran (int_tlv_word42[20], \int_tlv_word42.unused [12]);
tran (key_tlv_word0[19], \key_tlv_word0.tlv_seq_num [3]);
tran (int_tlv_word0[19], \int_tlv_word0.tlv_seq_num [3]);
tran (int_tlv_word42[19], \int_tlv_word42.unused [11]);
tran (key_tlv_word0[18], \key_tlv_word0.tlv_seq_num [2]);
tran (int_tlv_word0[18], \int_tlv_word0.tlv_seq_num [2]);
tran (int_tlv_word42[18], \int_tlv_word42.unused [10]);
tran (key_tlv_word0[17], \key_tlv_word0.tlv_seq_num [1]);
tran (int_tlv_word0[17], \int_tlv_word0.tlv_seq_num [1]);
tran (int_tlv_word42[17], \int_tlv_word42.unused [9]);
tran (key_tlv_word0[16], \key_tlv_word0.tlv_seq_num [0]);
tran (int_tlv_word0[16], \int_tlv_word0.tlv_seq_num [0]);
tran (int_tlv_word42[16], \int_tlv_word42.unused [8]);
tran (int_tlv_word0[15], \int_tlv_word0.tlv_len [7]);
tran (int_tlv_word42[15], \int_tlv_word42.unused [7]);
tran (int_tlv_word0[14], \int_tlv_word0.tlv_len [6]);
tran (int_tlv_word42[14], \int_tlv_word42.unused [6]);
tran (int_tlv_word0[13], \int_tlv_word0.tlv_len [5]);
tran (int_tlv_word42[13], \int_tlv_word42.unused [5]);
tran (int_tlv_word0[12], \int_tlv_word0.tlv_len [4]);
tran (int_tlv_word42[12], \int_tlv_word42.unused [4]);
tran (int_tlv_word0[11], \int_tlv_word0.tlv_len [3]);
tran (int_tlv_word42[11], \int_tlv_word42.unused [3]);
tran (int_tlv_word0[10], \int_tlv_word0.tlv_len [2]);
tran (int_tlv_word42[10], \int_tlv_word42.unused [2]);
tran (int_tlv_word0[9], \int_tlv_word0.tlv_len [1]);
tran (int_tlv_word42[9], \int_tlv_word42.unused [1]);
tran (int_tlv_word0[8], \int_tlv_word0.tlv_len [0]);
tran (int_tlv_word42[8], \int_tlv_word42.unused [0]);
tran (int_tlv_word0[7], \int_tlv_word0.tlv_type [7]);
tran (int_tlv_word42[7], \int_tlv_word42.error_code [7]);
tran (int_tlv_word0[6], \int_tlv_word0.tlv_type [6]);
tran (int_tlv_word42[6], \int_tlv_word42.error_code [6]);
tran (int_tlv_word0[5], \int_tlv_word0.tlv_type [5]);
tran (int_tlv_word42[5], \int_tlv_word42.error_code [5]);
tran (int_tlv_word0[4], \int_tlv_word0.tlv_type [4]);
tran (int_tlv_word42[4], \int_tlv_word42.error_code [4]);
tran (int_tlv_word0[3], \int_tlv_word0.tlv_type [3]);
tran (int_tlv_word42[3], \int_tlv_word42.error_code [3]);
tran (int_tlv_word0[2], \int_tlv_word0.tlv_type [2]);
tran (int_tlv_word42[2], \int_tlv_word42.error_code [2]);
tran (int_tlv_word0[1], \int_tlv_word0.tlv_type [1]);
tran (int_tlv_word42[1], \int_tlv_word42.error_code [1]);
tran (int_tlv_word0[0], \int_tlv_word0.tlv_type [0]);
tran (int_tlv_word42[0], \int_tlv_word42.error_code [0]);
tran (key_tlv_word20[0], \key_tlv_word20.crc32 [0]);
tran (key_tlv_word20[1], \key_tlv_word20.crc32 [1]);
tran (key_tlv_word20[2], \key_tlv_word20.crc32 [2]);
tran (key_tlv_word20[3], \key_tlv_word20.crc32 [3]);
tran (key_tlv_word20[4], \key_tlv_word20.crc32 [4]);
tran (key_tlv_word20[5], \key_tlv_word20.crc32 [5]);
tran (key_tlv_word20[6], \key_tlv_word20.crc32 [6]);
tran (key_tlv_word20[7], \key_tlv_word20.crc32 [7]);
tran (key_tlv_word20[8], \key_tlv_word20.crc32 [8]);
tran (key_tlv_word20[9], \key_tlv_word20.crc32 [9]);
tran (key_tlv_word20[10], \key_tlv_word20.crc32 [10]);
tran (key_tlv_word20[11], \key_tlv_word20.crc32 [11]);
tran (key_tlv_word20[12], \key_tlv_word20.crc32 [12]);
tran (key_tlv_word20[13], \key_tlv_word20.crc32 [13]);
tran (key_tlv_word20[14], \key_tlv_word20.crc32 [14]);
tran (key_tlv_word20[15], \key_tlv_word20.crc32 [15]);
tran (key_tlv_word20[16], \key_tlv_word20.crc32 [16]);
tran (key_tlv_word20[17], \key_tlv_word20.crc32 [17]);
tran (key_tlv_word20[18], \key_tlv_word20.crc32 [18]);
tran (key_tlv_word20[19], \key_tlv_word20.crc32 [19]);
tran (key_tlv_word20[20], \key_tlv_word20.crc32 [20]);
tran (key_tlv_word20[21], \key_tlv_word20.crc32 [21]);
tran (key_tlv_word20[22], \key_tlv_word20.crc32 [22]);
tran (key_tlv_word20[23], \key_tlv_word20.crc32 [23]);
tran (key_tlv_word20[24], \key_tlv_word20.crc32 [24]);
tran (key_tlv_word20[25], \key_tlv_word20.crc32 [25]);
tran (key_tlv_word20[26], \key_tlv_word20.crc32 [26]);
tran (key_tlv_word20[27], \key_tlv_word20.crc32 [27]);
tran (key_tlv_word20[28], \key_tlv_word20.crc32 [28]);
tran (key_tlv_word20[29], \key_tlv_word20.crc32 [29]);
tran (key_tlv_word20[30], \key_tlv_word20.crc32 [30]);
tran (key_tlv_word20[31], \key_tlv_word20.crc32 [31]);
tran (key_tlv_word20[32], \key_tlv_word20.rsvd [0]);
tran (key_tlv_word20[33], \key_tlv_word20.rsvd [1]);
tran (key_tlv_word20[34], \key_tlv_word20.rsvd [2]);
tran (key_tlv_word20[35], \key_tlv_word20.rsvd [3]);
tran (key_tlv_word20[36], \key_tlv_word20.rsvd [4]);
tran (key_tlv_word20[37], \key_tlv_word20.rsvd [5]);
tran (key_tlv_word20[38], \key_tlv_word20.rsvd [6]);
tran (key_tlv_word20[39], \key_tlv_word20.rsvd [7]);
tran (key_tlv_word20[40], \key_tlv_word20.rsvd [8]);
tran (key_tlv_word20[41], \key_tlv_word20.rsvd [9]);
tran (key_tlv_word20[42], \key_tlv_word20.rsvd [10]);
tran (key_tlv_word20[43], \key_tlv_word20.rsvd [11]);
tran (key_tlv_word20[44], \key_tlv_word20.rsvd [12]);
tran (key_tlv_word20[45], \key_tlv_word20.rsvd [13]);
tran (key_tlv_word20[46], \key_tlv_word20.rsvd [14]);
tran (key_tlv_word20[47], \key_tlv_word20.rsvd [15]);
tran (key_tlv_word20[48], \key_tlv_word20.rsvd [16]);
tran (key_tlv_word20[49], \key_tlv_word20.rsvd [17]);
tran (key_tlv_word20[50], \key_tlv_word20.rsvd [18]);
tran (key_tlv_word20[51], \key_tlv_word20.rsvd [19]);
tran (key_tlv_word20[52], \key_tlv_word20.rsvd [20]);
tran (key_tlv_word20[53], \key_tlv_word20.rsvd [21]);
tran (key_tlv_word20[54], \key_tlv_word20.rsvd [22]);
tran (key_tlv_word20[55], \key_tlv_word20.rsvd [23]);
tran (key_tlv_word20[56], \key_tlv_word20.rsvd [24]);
tran (key_tlv_word20[57], \key_tlv_word20.rsvd [25]);
tran (key_tlv_word20[58], \key_tlv_word20.rsvd [26]);
tran (key_tlv_word20[59], \key_tlv_word20.rsvd [27]);
tran (key_tlv_word20[60], \key_tlv_word20.rsvd [28]);
tran (key_tlv_word20[61], \key_tlv_word20.rsvd [29]);
tran (key_tlv_word20[62], \key_tlv_word20.rsvd [30]);
tran (key_tlv_word20[63], \key_tlv_word20.rsvd [31]);
tran (key_tlv_word19[0], \key_tlv_word19.kme_errors [0]);
tran (key_tlv_word19[1], \key_tlv_word19.kme_errors [1]);
tran (key_tlv_word19[2], \key_tlv_word19.kme_errors [2]);
tran (key_tlv_word19[3], \key_tlv_word19.kme_errors [3]);
tran (key_tlv_word19[4], \key_tlv_word19.kme_errors [4]);
tran (key_tlv_word19[5], \key_tlv_word19.kme_errors [5]);
tran (key_tlv_word19[6], \key_tlv_word19.kme_errors [6]);
tran (key_tlv_word19[7], \key_tlv_word19.kme_errors [7]);
tran (key_tlv_word19[8], \key_tlv_word19.rsvd [0]);
tran (key_tlv_word19[9], \key_tlv_word19.rsvd [1]);
tran (key_tlv_word19[10], \key_tlv_word19.rsvd [2]);
tran (key_tlv_word19[11], \key_tlv_word19.rsvd [3]);
tran (key_tlv_word19[12], \key_tlv_word19.rsvd [4]);
tran (key_tlv_word19[13], \key_tlv_word19.rsvd [5]);
tran (key_tlv_word19[14], \key_tlv_word19.rsvd [6]);
tran (key_tlv_word19[15], \key_tlv_word19.rsvd [7]);
tran (key_tlv_word19[16], \key_tlv_word19.rsvd [8]);
tran (key_tlv_word19[17], \key_tlv_word19.rsvd [9]);
tran (key_tlv_word19[18], \key_tlv_word19.rsvd [10]);
tran (key_tlv_word19[19], \key_tlv_word19.rsvd [11]);
tran (key_tlv_word19[20], \key_tlv_word19.rsvd [12]);
tran (key_tlv_word19[21], \key_tlv_word19.rsvd [13]);
tran (key_tlv_word19[22], \key_tlv_word19.rsvd [14]);
tran (key_tlv_word19[23], \key_tlv_word19.rsvd [15]);
tran (key_tlv_word19[24], \key_tlv_word19.rsvd [16]);
tran (key_tlv_word19[25], \key_tlv_word19.rsvd [17]);
tran (key_tlv_word19[26], \key_tlv_word19.rsvd [18]);
tran (key_tlv_word19[27], \key_tlv_word19.rsvd [19]);
tran (key_tlv_word19[28], \key_tlv_word19.rsvd [20]);
tran (key_tlv_word19[29], \key_tlv_word19.rsvd [21]);
tran (key_tlv_word19[30], \key_tlv_word19.rsvd [22]);
tran (key_tlv_word19[31], \key_tlv_word19.rsvd [23]);
tran (key_tlv_word19[32], \key_tlv_word19.rsvd [24]);
tran (key_tlv_word19[33], \key_tlv_word19.rsvd [25]);
tran (key_tlv_word19[34], \key_tlv_word19.rsvd [26]);
tran (key_tlv_word19[35], \key_tlv_word19.rsvd [27]);
tran (key_tlv_word19[36], \key_tlv_word19.rsvd [28]);
tran (key_tlv_word19[37], \key_tlv_word19.rsvd [29]);
tran (key_tlv_word19[38], \key_tlv_word19.rsvd [30]);
tran (key_tlv_word19[39], \key_tlv_word19.rsvd [31]);
tran (key_tlv_word19[40], \key_tlv_word19.rsvd [32]);
tran (key_tlv_word19[41], \key_tlv_word19.rsvd [33]);
tran (key_tlv_word19[42], \key_tlv_word19.rsvd [34]);
tran (key_tlv_word19[43], \key_tlv_word19.rsvd [35]);
tran (key_tlv_word19[44], \key_tlv_word19.rsvd [36]);
tran (key_tlv_word19[45], \key_tlv_word19.rsvd [37]);
tran (key_tlv_word19[46], \key_tlv_word19.rsvd [38]);
tran (key_tlv_word19[47], \key_tlv_word19.rsvd [39]);
tran (key_tlv_word19[48], \key_tlv_word19.rsvd [40]);
tran (key_tlv_word19[49], \key_tlv_word19.rsvd [41]);
tran (key_tlv_word19[50], \key_tlv_word19.rsvd [42]);
tran (key_tlv_word19[51], \key_tlv_word19.rsvd [43]);
tran (key_tlv_word19[52], \key_tlv_word19.rsvd [44]);
tran (key_tlv_word19[53], \key_tlv_word19.rsvd [45]);
tran (key_tlv_word19[54], \key_tlv_word19.rsvd [46]);
tran (key_tlv_word19[55], \key_tlv_word19.rsvd [47]);
tran (key_tlv_word19[56], \key_tlv_word19.rsvd [48]);
tran (key_tlv_word19[57], \key_tlv_word19.rsvd [49]);
tran (key_tlv_word19[58], \key_tlv_word19.rsvd [50]);
tran (key_tlv_word19[59], \key_tlv_word19.rsvd [51]);
tran (key_tlv_word19[60], \key_tlv_word19.rsvd [52]);
tran (key_tlv_word19[61], \key_tlv_word19.rsvd [53]);
tran (key_tlv_word19[62], \key_tlv_word19.rsvd [54]);
tran (key_tlv_word19[63], \key_tlv_word19.rsvd [55]);
tran (key_tlv_word0[0], \key_tlv_word0.tlv_type [0]);
tran (key_tlv_word0[1], \key_tlv_word0.tlv_type [1]);
tran (key_tlv_word0[2], \key_tlv_word0.tlv_type [2]);
tran (key_tlv_word0[3], \key_tlv_word0.tlv_type [3]);
tran (key_tlv_word0[4], \key_tlv_word0.tlv_type [4]);
tran (key_tlv_word0[5], \key_tlv_word0.tlv_type [5]);
tran (key_tlv_word0[6], \key_tlv_word0.tlv_type [6]);
tran (key_tlv_word0[7], \key_tlv_word0.tlv_type [7]);
tran (key_tlv_word0[8], \key_tlv_word0.tlv_len [0]);
tran (key_tlv_word0[9], \key_tlv_word0.tlv_len [1]);
tran (key_tlv_word0[10], \key_tlv_word0.tlv_len [2]);
tran (key_tlv_word0[11], \key_tlv_word0.tlv_len [3]);
tran (key_tlv_word0[12], \key_tlv_word0.tlv_len [4]);
tran (key_tlv_word0[13], \key_tlv_word0.tlv_len [5]);
tran (key_tlv_word0[14], \key_tlv_word0.tlv_len [6]);
tran (key_tlv_word0[15], \key_tlv_word0.tlv_len [7]);
tran (key_tlv_word0[28], \key_tlv_word0.resv1 [0]);
tran (key_tlv_word0[29], \key_tlv_word0.resv1 [1]);
tran (key_tlv_word0[30], \key_tlv_word0.resv1 [2]);
tran (key_tlv_word0[31], \key_tlv_word0.resv1 [3]);
tran (key_tlv_word0[43], \key_tlv_word0.resv0 [0]);
tran (key_tlv_word0[44], \key_tlv_word0.resv0 [1]);
tran (key_tlv_word0[45], \key_tlv_word0.resv0 [2]);
tran (key_tlv_word0[46], \key_tlv_word0.resv0 [3]);
tran (key_tlv_word0[47], \key_tlv_word0.resv0 [4]);
tran (key_tlv_word0[48], \key_tlv_word0.resv0 [5]);
tran (key_tlv_word0[49], \key_tlv_word0.resv0 [6]);
tran (key_tlv_word0[50], \key_tlv_word0.resv0 [7]);
tran (key_tlv_word0[51], \key_tlv_word0.resv0 [8]);
tran (key_tlv_word0[52], \key_tlv_word0.resv0 [9]);
tran (key_tlv_word0[53], \key_tlv_word0.resv0 [10]);
tran (key_tlv_word0[54], \key_tlv_word0.resv0 [11]);
tran (key_tlv_word0[55], \key_tlv_word0.resv0 [12]);
tran (key_tlv_word0[56], \key_tlv_word0.resv0 [13]);
tran (key_tlv_word0[57], \key_tlv_word0.resv0 [14]);
tran (key_tlv_word0[58], \key_tlv_word0.resv0 [15]);
tran (key_tlv_word0[59], \key_tlv_word0.resv0 [16]);
tran (key_tlv_word0[60], \key_tlv_word0.resv0 [17]);
tran (key_tlv_word0[61], \key_tlv_word0.resv0 [18]);
tran (key_tlv_word0[62], \key_tlv_word0.tlv_bip2 [0]);
tran (key_tlv_word0[63], \key_tlv_word0.tlv_bip2 [1]);
Q_BUF U0 ( .A(n314), .Z(key_tlv_word0[63]));
Q_BUF U1 ( .A(n314), .Z(key_tlv_word0[62]));
Q_BUF U2 ( .A(n314), .Z(key_tlv_word0[61]));
Q_BUF U3 ( .A(n314), .Z(key_tlv_word0[60]));
Q_BUF U4 ( .A(n314), .Z(key_tlv_word0[59]));
Q_BUF U5 ( .A(n314), .Z(key_tlv_word0[58]));
Q_BUF U6 ( .A(n314), .Z(key_tlv_word0[57]));
Q_BUF U7 ( .A(n314), .Z(key_tlv_word0[56]));
Q_BUF U8 ( .A(n314), .Z(key_tlv_word0[55]));
Q_BUF U9 ( .A(n314), .Z(key_tlv_word0[54]));
Q_BUF U10 ( .A(n314), .Z(key_tlv_word0[53]));
Q_BUF U11 ( .A(n314), .Z(key_tlv_word0[52]));
Q_BUF U12 ( .A(n314), .Z(key_tlv_word0[51]));
Q_BUF U13 ( .A(n314), .Z(key_tlv_word0[50]));
Q_BUF U14 ( .A(n314), .Z(key_tlv_word0[49]));
Q_BUF U15 ( .A(n314), .Z(key_tlv_word0[48]));
Q_BUF U16 ( .A(n314), .Z(key_tlv_word0[47]));
Q_BUF U17 ( .A(n314), .Z(key_tlv_word0[46]));
Q_BUF U18 ( .A(n314), .Z(key_tlv_word0[45]));
Q_BUF U19 ( .A(n314), .Z(key_tlv_word0[44]));
Q_BUF U20 ( .A(n314), .Z(key_tlv_word0[43]));
Q_BUF U21 ( .A(n314), .Z(key_tlv_word0[31]));
Q_BUF U22 ( .A(n314), .Z(key_tlv_word0[30]));
Q_BUF U23 ( .A(n314), .Z(key_tlv_word0[29]));
Q_BUF U24 ( .A(n314), .Z(key_tlv_word0[28]));
Q_BUF U25 ( .A(n315), .Z(key_tlv_word0[15]));
Q_BUF U26 ( .A(n314), .Z(key_tlv_word0[14]));
Q_BUF U27 ( .A(n315), .Z(key_tlv_word0[13]));
Q_BUF U28 ( .A(n314), .Z(key_tlv_word0[12]));
Q_BUF U29 ( .A(n315), .Z(key_tlv_word0[11]));
Q_BUF U30 ( .A(n314), .Z(key_tlv_word0[10]));
Q_BUF U31 ( .A(n314), .Z(key_tlv_word0[9]));
Q_BUF U32 ( .A(n314), .Z(key_tlv_word0[8]));
Q_BUF U33 ( .A(n314), .Z(key_tlv_word0[7]));
Q_BUF U34 ( .A(n314), .Z(key_tlv_word0[6]));
Q_BUF U35 ( .A(n314), .Z(key_tlv_word0[5]));
Q_BUF U36 ( .A(n314), .Z(key_tlv_word0[4]));
Q_BUF U37 ( .A(n314), .Z(key_tlv_word0[3]));
Q_BUF U38 ( .A(n314), .Z(key_tlv_word0[2]));
Q_BUF U39 ( .A(n315), .Z(key_tlv_word0[1]));
Q_BUF U40 ( .A(n314), .Z(key_tlv_word0[0]));
Q_BUF U41 ( .A(n314), .Z(key_tlv_word19[63]));
Q_BUF U42 ( .A(n314), .Z(key_tlv_word19[62]));
Q_BUF U43 ( .A(n314), .Z(key_tlv_word19[61]));
Q_BUF U44 ( .A(n314), .Z(key_tlv_word19[60]));
Q_BUF U45 ( .A(n314), .Z(key_tlv_word19[59]));
Q_BUF U46 ( .A(n314), .Z(key_tlv_word19[58]));
Q_BUF U47 ( .A(n314), .Z(key_tlv_word19[57]));
Q_BUF U48 ( .A(n314), .Z(key_tlv_word19[56]));
Q_BUF U49 ( .A(n314), .Z(key_tlv_word19[55]));
Q_BUF U50 ( .A(n314), .Z(key_tlv_word19[54]));
Q_BUF U51 ( .A(n314), .Z(key_tlv_word19[53]));
Q_BUF U52 ( .A(n314), .Z(key_tlv_word19[52]));
Q_BUF U53 ( .A(n314), .Z(key_tlv_word19[51]));
Q_BUF U54 ( .A(n314), .Z(key_tlv_word19[50]));
Q_BUF U55 ( .A(n314), .Z(key_tlv_word19[49]));
Q_BUF U56 ( .A(n314), .Z(key_tlv_word19[48]));
Q_BUF U57 ( .A(n314), .Z(key_tlv_word19[47]));
Q_BUF U58 ( .A(n314), .Z(key_tlv_word19[46]));
Q_BUF U59 ( .A(n314), .Z(key_tlv_word19[45]));
Q_BUF U60 ( .A(n314), .Z(key_tlv_word19[44]));
Q_BUF U61 ( .A(n314), .Z(key_tlv_word19[43]));
Q_BUF U62 ( .A(n314), .Z(key_tlv_word19[42]));
Q_BUF U63 ( .A(n314), .Z(key_tlv_word19[41]));
Q_BUF U64 ( .A(n314), .Z(key_tlv_word19[40]));
Q_BUF U65 ( .A(n314), .Z(key_tlv_word19[39]));
Q_BUF U66 ( .A(n314), .Z(key_tlv_word19[38]));
Q_BUF U67 ( .A(n314), .Z(key_tlv_word19[37]));
Q_BUF U68 ( .A(n314), .Z(key_tlv_word19[36]));
Q_BUF U69 ( .A(n314), .Z(key_tlv_word19[35]));
Q_BUF U70 ( .A(n314), .Z(key_tlv_word19[34]));
Q_BUF U71 ( .A(n314), .Z(key_tlv_word19[33]));
Q_BUF U72 ( .A(n314), .Z(key_tlv_word19[32]));
Q_BUF U73 ( .A(n314), .Z(key_tlv_word19[31]));
Q_BUF U74 ( .A(n314), .Z(key_tlv_word19[30]));
Q_BUF U75 ( .A(n314), .Z(key_tlv_word19[29]));
Q_BUF U76 ( .A(n314), .Z(key_tlv_word19[28]));
Q_BUF U77 ( .A(n314), .Z(key_tlv_word19[27]));
Q_BUF U78 ( .A(n314), .Z(key_tlv_word19[26]));
Q_BUF U79 ( .A(n314), .Z(key_tlv_word19[25]));
Q_BUF U80 ( .A(n314), .Z(key_tlv_word19[24]));
Q_BUF U81 ( .A(n314), .Z(key_tlv_word19[23]));
Q_BUF U82 ( .A(n314), .Z(key_tlv_word19[22]));
Q_BUF U83 ( .A(n314), .Z(key_tlv_word19[21]));
Q_BUF U84 ( .A(n314), .Z(key_tlv_word19[20]));
Q_BUF U85 ( .A(n314), .Z(key_tlv_word19[19]));
Q_BUF U86 ( .A(n314), .Z(key_tlv_word19[18]));
Q_BUF U87 ( .A(n314), .Z(key_tlv_word19[17]));
Q_BUF U88 ( .A(n314), .Z(key_tlv_word19[16]));
Q_BUF U89 ( .A(n314), .Z(key_tlv_word19[15]));
Q_BUF U90 ( .A(n314), .Z(key_tlv_word19[14]));
Q_BUF U91 ( .A(n314), .Z(key_tlv_word19[13]));
Q_BUF U92 ( .A(n314), .Z(key_tlv_word19[12]));
Q_BUF U93 ( .A(n314), .Z(key_tlv_word19[11]));
Q_BUF U94 ( .A(n314), .Z(key_tlv_word19[10]));
Q_BUF U95 ( .A(n314), .Z(key_tlv_word19[9]));
Q_BUF U96 ( .A(n314), .Z(key_tlv_word19[8]));
Q_BUF U97 ( .A(n314), .Z(key_tlv_word20[63]));
Q_BUF U98 ( .A(n314), .Z(key_tlv_word20[62]));
Q_BUF U99 ( .A(n314), .Z(key_tlv_word20[61]));
Q_BUF U100 ( .A(n314), .Z(key_tlv_word20[60]));
Q_BUF U101 ( .A(n314), .Z(key_tlv_word20[59]));
Q_BUF U102 ( .A(n314), .Z(key_tlv_word20[58]));
Q_BUF U103 ( .A(n314), .Z(key_tlv_word20[57]));
Q_BUF U104 ( .A(n314), .Z(key_tlv_word20[56]));
Q_BUF U105 ( .A(n314), .Z(key_tlv_word20[55]));
Q_BUF U106 ( .A(n314), .Z(key_tlv_word20[54]));
Q_BUF U107 ( .A(n314), .Z(key_tlv_word20[53]));
Q_BUF U108 ( .A(n314), .Z(key_tlv_word20[52]));
Q_BUF U109 ( .A(n314), .Z(key_tlv_word20[51]));
Q_BUF U110 ( .A(n314), .Z(key_tlv_word20[50]));
Q_BUF U111 ( .A(n314), .Z(key_tlv_word20[49]));
Q_BUF U112 ( .A(n314), .Z(key_tlv_word20[48]));
Q_BUF U113 ( .A(n314), .Z(key_tlv_word20[47]));
Q_BUF U114 ( .A(n314), .Z(key_tlv_word20[46]));
Q_BUF U115 ( .A(n314), .Z(key_tlv_word20[45]));
Q_BUF U116 ( .A(n314), .Z(key_tlv_word20[44]));
Q_BUF U117 ( .A(n314), .Z(key_tlv_word20[43]));
Q_BUF U118 ( .A(n314), .Z(key_tlv_word20[42]));
Q_BUF U119 ( .A(n314), .Z(key_tlv_word20[41]));
Q_BUF U120 ( .A(n314), .Z(key_tlv_word20[40]));
Q_BUF U121 ( .A(n314), .Z(key_tlv_word20[39]));
Q_BUF U122 ( .A(n314), .Z(key_tlv_word20[38]));
Q_BUF U123 ( .A(n314), .Z(key_tlv_word20[37]));
Q_BUF U124 ( .A(n314), .Z(key_tlv_word20[36]));
Q_BUF U125 ( .A(n314), .Z(key_tlv_word20[35]));
Q_BUF U126 ( .A(n314), .Z(key_tlv_word20[34]));
Q_BUF U127 ( .A(n314), .Z(key_tlv_word20[33]));
Q_BUF U128 ( .A(n314), .Z(key_tlv_word20[32]));
Q_BUF U129 ( .A(n315), .Z(_zy_simnet_cio_6[0]));
Q_BUF U130 ( .A(n315), .Z(_zy_simnet_cio_6[1]));
Q_BUF U131 ( .A(n315), .Z(_zy_simnet_cio_6[2]));
Q_BUF U132 ( .A(n315), .Z(_zy_simnet_cio_6[3]));
Q_BUF U133 ( .A(n315), .Z(_zy_simnet_cio_6[4]));
Q_BUF U134 ( .A(n315), .Z(_zy_simnet_cio_6[5]));
Q_BUF U135 ( .A(n315), .Z(_zy_simnet_cio_6[6]));
Q_BUF U136 ( .A(n315), .Z(_zy_simnet_cio_6[7]));
Q_BUF U137 ( .A(n315), .Z(_zy_simnet_cio_7));
Q_BUF U138 ( .A(n315), .Z(_zy_simnet_cio_8[0]));
Q_BUF U139 ( .A(n315), .Z(_zy_simnet_cio_8[1]));
Q_BUF U140 ( .A(n315), .Z(_zy_simnet_cio_8[2]));
Q_BUF U141 ( .A(n315), .Z(_zy_simnet_cio_8[3]));
Q_BUF U142 ( .A(n315), .Z(_zy_simnet_cio_8[4]));
Q_BUF U143 ( .A(n315), .Z(_zy_simnet_cio_8[5]));
Q_BUF U144 ( .A(n315), .Z(_zy_simnet_cio_8[6]));
Q_BUF U145 ( .A(n315), .Z(_zy_simnet_cio_8[7]));
Q_BUF U146 ( .A(n315), .Z(_zy_simnet_cio_8[8]));
Q_BUF U147 ( .A(n315), .Z(_zy_simnet_cio_8[9]));
Q_BUF U148 ( .A(n315), .Z(_zy_simnet_cio_8[10]));
Q_BUF U149 ( .A(n315), .Z(_zy_simnet_cio_8[11]));
Q_BUF U150 ( .A(n315), .Z(_zy_simnet_cio_8[12]));
Q_BUF U151 ( .A(n315), .Z(_zy_simnet_cio_8[13]));
Q_BUF U152 ( .A(n315), .Z(_zy_simnet_cio_8[14]));
Q_BUF U153 ( .A(n315), .Z(_zy_simnet_cio_8[15]));
Q_BUF U154 ( .A(n315), .Z(_zy_simnet_cio_8[16]));
Q_BUF U155 ( .A(n315), .Z(_zy_simnet_cio_8[17]));
Q_BUF U156 ( .A(n315), .Z(_zy_simnet_cio_8[18]));
Q_BUF U157 ( .A(n315), .Z(_zy_simnet_cio_8[19]));
Q_BUF U158 ( .A(n315), .Z(_zy_simnet_cio_8[20]));
Q_BUF U159 ( .A(n315), .Z(_zy_simnet_cio_8[21]));
Q_BUF U160 ( .A(n315), .Z(_zy_simnet_cio_8[22]));
Q_BUF U161 ( .A(n315), .Z(_zy_simnet_cio_8[23]));
Q_BUF U162 ( .A(n315), .Z(_zy_simnet_cio_8[24]));
Q_BUF U163 ( .A(n315), .Z(_zy_simnet_cio_8[25]));
Q_BUF U164 ( .A(n315), .Z(_zy_simnet_cio_8[26]));
Q_BUF U165 ( .A(n315), .Z(_zy_simnet_cio_8[27]));
Q_BUF U166 ( .A(n315), .Z(_zy_simnet_cio_8[28]));
Q_BUF U167 ( .A(n315), .Z(_zy_simnet_cio_8[29]));
Q_BUF U168 ( .A(n315), .Z(_zy_simnet_cio_8[30]));
Q_BUF U169 ( .A(n315), .Z(_zy_simnet_cio_8[31]));
Q_ASSIGN U170 ( .B(tlv_sb_data_out[63]), .A(int_tlv_word0[63]));
Q_ASSIGN U171 ( .B(tlv_sb_data_out[62]), .A(int_tlv_word0[62]));
Q_ASSIGN U172 ( .B(tlv_sb_data_out[61]), .A(int_tlv_word0[61]));
Q_ASSIGN U173 ( .B(tlv_sb_data_out[60]), .A(int_tlv_word0[60]));
Q_ASSIGN U174 ( .B(tlv_sb_data_out[59]), .A(int_tlv_word0[59]));
Q_ASSIGN U175 ( .B(tlv_sb_data_out[58]), .A(int_tlv_word0[58]));
Q_ASSIGN U176 ( .B(tlv_sb_data_out[57]), .A(int_tlv_word0[57]));
Q_ASSIGN U177 ( .B(tlv_sb_data_out[56]), .A(int_tlv_word0[56]));
Q_ASSIGN U178 ( .B(tlv_sb_data_out[55]), .A(int_tlv_word0[55]));
Q_ASSIGN U179 ( .B(tlv_sb_data_out[55]), .A(int_tlv_word42[55]));
Q_ASSIGN U180 ( .B(tlv_sb_data_out[54]), .A(int_tlv_word0[54]));
Q_ASSIGN U181 ( .B(tlv_sb_data_out[54]), .A(int_tlv_word42[54]));
Q_ASSIGN U182 ( .B(tlv_sb_data_out[53]), .A(int_tlv_word0[53]));
Q_ASSIGN U183 ( .B(tlv_sb_data_out[53]), .A(int_tlv_word42[53]));
Q_ASSIGN U184 ( .B(tlv_sb_data_out[52]), .A(int_tlv_word0[52]));
Q_ASSIGN U185 ( .B(tlv_sb_data_out[52]), .A(int_tlv_word42[52]));
Q_ASSIGN U186 ( .B(tlv_sb_data_out[51]), .A(int_tlv_word0[51]));
Q_ASSIGN U187 ( .B(tlv_sb_data_out[51]), .A(int_tlv_word42[51]));
Q_ASSIGN U188 ( .B(tlv_sb_data_out[50]), .A(int_tlv_word0[50]));
Q_ASSIGN U189 ( .B(tlv_sb_data_out[50]), .A(int_tlv_word42[50]));
Q_ASSIGN U190 ( .B(tlv_sb_data_out[49]), .A(int_tlv_word0[49]));
Q_ASSIGN U191 ( .B(tlv_sb_data_out[49]), .A(int_tlv_word42[49]));
Q_ASSIGN U192 ( .B(tlv_sb_data_out[48]), .A(int_tlv_word0[48]));
Q_ASSIGN U193 ( .B(tlv_sb_data_out[48]), .A(int_tlv_word42[48]));
Q_ASSIGN U194 ( .B(tlv_sb_data_out[47]), .A(int_tlv_word0[47]));
Q_ASSIGN U195 ( .B(tlv_sb_data_out[47]), .A(int_tlv_word42[47]));
Q_ASSIGN U196 ( .B(tlv_sb_data_out[46]), .A(int_tlv_word0[46]));
Q_ASSIGN U197 ( .B(tlv_sb_data_out[46]), .A(int_tlv_word42[46]));
Q_ASSIGN U198 ( .B(tlv_sb_data_out[45]), .A(int_tlv_word0[45]));
Q_ASSIGN U199 ( .B(tlv_sb_data_out[45]), .A(int_tlv_word42[45]));
Q_ASSIGN U200 ( .B(tlv_sb_data_out[44]), .A(int_tlv_word0[44]));
Q_ASSIGN U201 ( .B(tlv_sb_data_out[44]), .A(int_tlv_word42[44]));
Q_ASSIGN U202 ( .B(tlv_sb_data_out[43]), .A(int_tlv_word0[43]));
Q_ASSIGN U203 ( .B(tlv_sb_data_out[43]), .A(int_tlv_word42[43]));
Q_ASSIGN U204 ( .B(tlv_sb_data_out[42]), .A(int_tlv_word0[42]));
Q_ASSIGN U205 ( .B(tlv_sb_data_out[42]), .A(int_tlv_word42[42]));
Q_ASSIGN U206 ( .B(tlv_sb_data_out[41]), .A(int_tlv_word0[41]));
Q_ASSIGN U207 ( .B(tlv_sb_data_out[41]), .A(int_tlv_word42[41]));
Q_ASSIGN U208 ( .B(tlv_sb_data_out[40]), .A(int_tlv_word0[40]));
Q_ASSIGN U209 ( .B(tlv_sb_data_out[40]), .A(int_tlv_word42[40]));
Q_ASSIGN U210 ( .B(tlv_sb_data_out[39]), .A(int_tlv_word0[39]));
Q_ASSIGN U211 ( .B(tlv_sb_data_out[39]), .A(int_tlv_word42[39]));
Q_ASSIGN U212 ( .B(tlv_sb_data_out[38]), .A(key_tlv_word0[42]));
Q_ASSIGN U213 ( .B(tlv_sb_data_out[38]), .A(int_tlv_word0[38]));
Q_ASSIGN U214 ( .B(tlv_sb_data_out[38]), .A(int_tlv_word42[38]));
Q_ASSIGN U215 ( .B(tlv_sb_data_out[37]), .A(key_tlv_word0[41]));
Q_ASSIGN U216 ( .B(tlv_sb_data_out[37]), .A(int_tlv_word0[37]));
Q_ASSIGN U217 ( .B(tlv_sb_data_out[37]), .A(int_tlv_word42[37]));
Q_ASSIGN U218 ( .B(tlv_sb_data_out[36]), .A(key_tlv_word0[40]));
Q_ASSIGN U219 ( .B(tlv_sb_data_out[36]), .A(int_tlv_word0[36]));
Q_ASSIGN U220 ( .B(tlv_sb_data_out[36]), .A(int_tlv_word42[36]));
Q_ASSIGN U221 ( .B(tlv_sb_data_out[35]), .A(key_tlv_word0[39]));
Q_ASSIGN U222 ( .B(tlv_sb_data_out[35]), .A(int_tlv_word0[35]));
Q_ASSIGN U223 ( .B(tlv_sb_data_out[35]), .A(int_tlv_word42[35]));
Q_ASSIGN U224 ( .B(tlv_sb_data_out[34]), .A(key_tlv_word0[38]));
Q_ASSIGN U225 ( .B(tlv_sb_data_out[34]), .A(int_tlv_word0[34]));
Q_ASSIGN U226 ( .B(tlv_sb_data_out[34]), .A(int_tlv_word42[34]));
Q_ASSIGN U227 ( .B(tlv_sb_data_out[33]), .A(key_tlv_word0[37]));
Q_ASSIGN U228 ( .B(tlv_sb_data_out[33]), .A(int_tlv_word0[33]));
Q_ASSIGN U229 ( .B(tlv_sb_data_out[33]), .A(int_tlv_word42[33]));
Q_ASSIGN U230 ( .B(tlv_sb_data_out[32]), .A(key_tlv_word0[36]));
Q_ASSIGN U231 ( .B(tlv_sb_data_out[32]), .A(int_tlv_word0[32]));
Q_ASSIGN U232 ( .B(tlv_sb_data_out[32]), .A(int_tlv_word42[32]));
Q_ASSIGN U233 ( .B(tlv_sb_data_out[31]), .A(key_tlv_word0[35]));
Q_ASSIGN U234 ( .B(tlv_sb_data_out[31]), .A(int_tlv_word0[31]));
Q_ASSIGN U235 ( .B(tlv_sb_data_out[31]), .A(int_tlv_word42[31]));
Q_ASSIGN U236 ( .B(tlv_sb_data_out[30]), .A(key_tlv_word0[34]));
Q_ASSIGN U237 ( .B(tlv_sb_data_out[30]), .A(int_tlv_word0[30]));
Q_ASSIGN U238 ( .B(tlv_sb_data_out[30]), .A(int_tlv_word42[30]));
Q_ASSIGN U239 ( .B(tlv_sb_data_out[29]), .A(key_tlv_word0[33]));
Q_ASSIGN U240 ( .B(tlv_sb_data_out[29]), .A(int_tlv_word0[29]));
Q_ASSIGN U241 ( .B(tlv_sb_data_out[29]), .A(int_tlv_word42[29]));
Q_ASSIGN U242 ( .B(tlv_sb_data_out[28]), .A(key_tlv_word0[32]));
Q_ASSIGN U243 ( .B(tlv_sb_data_out[28]), .A(int_tlv_word0[28]));
Q_ASSIGN U244 ( .B(tlv_sb_data_out[28]), .A(int_tlv_word42[28]));
Q_ASSIGN U245 ( .B(tlv_sb_data_out[27]), .A(key_tlv_word0[27]));
Q_ASSIGN U246 ( .B(tlv_sb_data_out[27]), .A(int_tlv_word0[27]));
Q_ASSIGN U247 ( .B(tlv_sb_data_out[27]), .A(int_tlv_word42[27]));
Q_ASSIGN U248 ( .B(tlv_sb_data_out[26]), .A(key_tlv_word0[26]));
Q_ASSIGN U249 ( .B(tlv_sb_data_out[26]), .A(int_tlv_word0[26]));
Q_ASSIGN U250 ( .B(tlv_sb_data_out[26]), .A(int_tlv_word42[26]));
Q_ASSIGN U251 ( .B(tlv_sb_data_out[25]), .A(key_tlv_word0[25]));
Q_ASSIGN U252 ( .B(tlv_sb_data_out[25]), .A(int_tlv_word0[25]));
Q_ASSIGN U253 ( .B(tlv_sb_data_out[25]), .A(int_tlv_word42[25]));
Q_ASSIGN U254 ( .B(tlv_sb_data_out[24]), .A(key_tlv_word0[24]));
Q_ASSIGN U255 ( .B(tlv_sb_data_out[24]), .A(int_tlv_word0[24]));
Q_ASSIGN U256 ( .B(tlv_sb_data_out[24]), .A(int_tlv_word42[24]));
Q_ASSIGN U257 ( .B(tlv_sb_data_out[23]), .A(key_tlv_word0[23]));
Q_ASSIGN U258 ( .B(tlv_sb_data_out[23]), .A(int_tlv_word0[23]));
Q_ASSIGN U259 ( .B(tlv_sb_data_out[23]), .A(int_tlv_word42[23]));
Q_ASSIGN U260 ( .B(tlv_sb_data_out[22]), .A(key_tlv_word0[22]));
Q_ASSIGN U261 ( .B(tlv_sb_data_out[22]), .A(int_tlv_word0[22]));
Q_ASSIGN U262 ( .B(tlv_sb_data_out[22]), .A(int_tlv_word42[22]));
Q_ASSIGN U263 ( .B(tlv_sb_data_out[21]), .A(key_tlv_word0[21]));
Q_ASSIGN U264 ( .B(tlv_sb_data_out[21]), .A(int_tlv_word0[21]));
Q_ASSIGN U265 ( .B(tlv_sb_data_out[21]), .A(int_tlv_word42[21]));
Q_ASSIGN U266 ( .B(tlv_sb_data_out[20]), .A(key_tlv_word0[20]));
Q_ASSIGN U267 ( .B(tlv_sb_data_out[20]), .A(int_tlv_word0[20]));
Q_ASSIGN U268 ( .B(tlv_sb_data_out[20]), .A(int_tlv_word42[20]));
Q_ASSIGN U269 ( .B(tlv_sb_data_out[19]), .A(key_tlv_word0[19]));
Q_ASSIGN U270 ( .B(tlv_sb_data_out[19]), .A(int_tlv_word0[19]));
Q_ASSIGN U271 ( .B(tlv_sb_data_out[19]), .A(int_tlv_word42[19]));
Q_ASSIGN U272 ( .B(tlv_sb_data_out[18]), .A(key_tlv_word0[18]));
Q_ASSIGN U273 ( .B(tlv_sb_data_out[18]), .A(int_tlv_word0[18]));
Q_ASSIGN U274 ( .B(tlv_sb_data_out[18]), .A(int_tlv_word42[18]));
Q_ASSIGN U275 ( .B(tlv_sb_data_out[17]), .A(key_tlv_word0[17]));
Q_ASSIGN U276 ( .B(tlv_sb_data_out[17]), .A(int_tlv_word0[17]));
Q_ASSIGN U277 ( .B(tlv_sb_data_out[17]), .A(int_tlv_word42[17]));
Q_ASSIGN U278 ( .B(tlv_sb_data_out[16]), .A(key_tlv_word0[16]));
Q_ASSIGN U279 ( .B(tlv_sb_data_out[16]), .A(int_tlv_word0[16]));
Q_ASSIGN U280 ( .B(tlv_sb_data_out[16]), .A(int_tlv_word42[16]));
Q_ASSIGN U281 ( .B(tlv_sb_data_out[15]), .A(int_tlv_word0[15]));
Q_ASSIGN U282 ( .B(tlv_sb_data_out[15]), .A(int_tlv_word42[15]));
Q_ASSIGN U283 ( .B(tlv_sb_data_out[14]), .A(int_tlv_word0[14]));
Q_ASSIGN U284 ( .B(tlv_sb_data_out[14]), .A(int_tlv_word42[14]));
Q_ASSIGN U285 ( .B(tlv_sb_data_out[13]), .A(int_tlv_word0[13]));
Q_ASSIGN U286 ( .B(tlv_sb_data_out[13]), .A(int_tlv_word42[13]));
Q_ASSIGN U287 ( .B(tlv_sb_data_out[12]), .A(int_tlv_word0[12]));
Q_ASSIGN U288 ( .B(tlv_sb_data_out[12]), .A(int_tlv_word42[12]));
Q_ASSIGN U289 ( .B(tlv_sb_data_out[11]), .A(int_tlv_word0[11]));
Q_ASSIGN U290 ( .B(tlv_sb_data_out[11]), .A(int_tlv_word42[11]));
Q_ASSIGN U291 ( .B(tlv_sb_data_out[10]), .A(int_tlv_word0[10]));
Q_ASSIGN U292 ( .B(tlv_sb_data_out[10]), .A(int_tlv_word42[10]));
Q_ASSIGN U293 ( .B(tlv_sb_data_out[9]), .A(int_tlv_word0[9]));
Q_ASSIGN U294 ( .B(tlv_sb_data_out[9]), .A(int_tlv_word42[9]));
Q_ASSIGN U295 ( .B(tlv_sb_data_out[8]), .A(int_tlv_word0[8]));
Q_ASSIGN U296 ( .B(tlv_sb_data_out[8]), .A(int_tlv_word42[8]));
Q_ASSIGN U297 ( .B(tlv_sb_data_out[7]), .A(int_tlv_word0[7]));
Q_ASSIGN U298 ( .B(tlv_sb_data_out[7]), .A(int_tlv_word42[7]));
Q_ASSIGN U299 ( .B(tlv_sb_data_out[6]), .A(int_tlv_word0[6]));
Q_ASSIGN U300 ( .B(tlv_sb_data_out[6]), .A(int_tlv_word42[6]));
Q_ASSIGN U301 ( .B(tlv_sb_data_out[5]), .A(int_tlv_word0[5]));
Q_ASSIGN U302 ( .B(tlv_sb_data_out[5]), .A(int_tlv_word42[5]));
Q_ASSIGN U303 ( .B(tlv_sb_data_out[4]), .A(int_tlv_word0[4]));
Q_ASSIGN U304 ( .B(tlv_sb_data_out[4]), .A(int_tlv_word42[4]));
Q_ASSIGN U305 ( .B(tlv_sb_data_out[3]), .A(int_tlv_word0[3]));
Q_ASSIGN U306 ( .B(tlv_sb_data_out[3]), .A(int_tlv_word42[3]));
Q_ASSIGN U307 ( .B(tlv_sb_data_out[2]), .A(int_tlv_word0[2]));
Q_ASSIGN U308 ( .B(tlv_sb_data_out[2]), .A(int_tlv_word42[2]));
Q_ASSIGN U309 ( .B(tlv_sb_data_out[1]), .A(int_tlv_word0[1]));
Q_ASSIGN U310 ( .B(tlv_sb_data_out[1]), .A(int_tlv_word42[1]));
Q_ASSIGN U311 ( .B(tlv_sb_data_out[0]), .A(int_tlv_word0[0]));
Q_ASSIGN U312 ( .B(tlv_sb_data_out[0]), .A(int_tlv_word42[0]));
Q_BUF U313 ( .A(n314), .Z(key_tlv_ob_tlv[105]));
Q_BUF U314 ( .A(n314), .Z(key_tlv_ob_tlv[104]));
Q_BUF U315 ( .A(n314), .Z(key_tlv_ob_tlv[103]));
Q_BUF U316 ( .A(n314), .Z(key_tlv_ob_tlv[102]));
Q_BUF U317 ( .A(n314), .Z(key_tlv_ob_tlv[101]));
Q_BUF U318 ( .A(n314), .Z(key_tlv_ob_tlv[100]));
Q_BUF U319 ( .A(n314), .Z(key_tlv_ob_tlv[99]));
Q_BUF U320 ( .A(n314), .Z(key_tlv_ob_tlv[98]));
Q_BUF U321 ( .A(n314), .Z(key_tlv_ob_tlv[97]));
Q_BUF U322 ( .A(n314), .Z(key_tlv_ob_tlv[96]));
Q_BUF U323 ( .A(n314), .Z(key_tlv_ob_tlv[95]));
Q_BUF U324 ( .A(n314), .Z(key_tlv_ob_tlv[94]));
Q_BUF U325 ( .A(n314), .Z(key_tlv_ob_tlv[93]));
Q_BUF U326 ( .A(n314), .Z(key_tlv_ob_tlv[92]));
Q_BUF U327 ( .A(n314), .Z(key_tlv_ob_tlv[91]));
Q_BUF U328 ( .A(n314), .Z(key_tlv_ob_tlv[90]));
Q_BUF U329 ( .A(n314), .Z(key_tlv_ob_tlv[89]));
Q_BUF U330 ( .A(n314), .Z(key_tlv_ob_tlv[88]));
Q_BUF U331 ( .A(n314), .Z(key_tlv_ob_tlv[87]));
Q_BUF U332 ( .A(n314), .Z(key_tlv_ob_tlv[86]));
Q_BUF U333 ( .A(n315), .Z(key_tlv_ob_tlv[85]));
Q_BUF U334 ( .A(n314), .Z(key_tlv_ob_tlv[84]));
Q_BUF U335 ( .A(key_tlv_ob_tlv[83]), .Z(key_tlv_ob_tlv[64]));
Q_BUF U336 ( .A(n314), .Z(key_tlv_ob_tlv[81]));
Q_BUF U337 ( .A(n314), .Z(key_tlv_ob_tlv[80]));
Q_BUF U338 ( .A(n315), .Z(key_tlv_ob_tlv[79]));
Q_BUF U339 ( .A(n315), .Z(key_tlv_ob_tlv[78]));
Q_BUF U340 ( .A(n315), .Z(key_tlv_ob_tlv[77]));
Q_BUF U341 ( .A(n315), .Z(key_tlv_ob_tlv[76]));
Q_BUF U342 ( .A(n315), .Z(key_tlv_ob_tlv[75]));
Q_BUF U343 ( .A(n315), .Z(key_tlv_ob_tlv[74]));
Q_BUF U344 ( .A(n315), .Z(key_tlv_ob_tlv[73]));
Q_BUF U345 ( .A(n315), .Z(key_tlv_ob_tlv[72]));
Q_BUF U346 ( .A(n314), .Z(key_tlv_ob_tlv[71]));
Q_BUF U347 ( .A(n314), .Z(key_tlv_ob_tlv[70]));
Q_BUF U348 ( .A(n314), .Z(key_tlv_ob_tlv[69]));
Q_BUF U349 ( .A(n314), .Z(key_tlv_ob_tlv[68]));
Q_BUF U350 ( .A(n314), .Z(key_tlv_ob_tlv[67]));
Q_BUF U351 ( .A(n314), .Z(key_tlv_ob_tlv[66]));
Q_AN02 U352 ( .A0(n275), .A1(n294), .Z(n1));
Q_AN02 U353 ( .A0(n282), .A1(n294), .Z(n2));
Q_ND02 U354 ( .A0(cur_state[1]), .A1(cur_state[0]), .Z(n22));
Q_AN02 U355 ( .A0(n22), .A1(n33), .Z(n16));
Q_AN02 U356 ( .A0(cur_state[2]), .A1(n277), .Z(n30));
Q_OA21 U357 ( .A0(n16), .A1(n30), .B0(n44), .Z(tlv_sb_data_out_ack));
Q_INV U358 ( .A(key_tlv_ob_full), .Z(n44));
Q_NR02 U359 ( .A0(cur_state[2]), .A1(n22), .Z(n24));
Q_NR02 U360 ( .A0(cur_state[1]), .A1(cur_state[0]), .Z(n32));
Q_AN02 U361 ( .A0(cur_state[2]), .A1(n32), .Z(n25));
Q_OR02 U362 ( .A0(n24), .A1(n25), .Z(n41));
Q_AN02 U363 ( .A0(tlv_sb_data_out_valid), .A1(gcm_status_data_out_valid), .Z(n39));
Q_AN03 U364 ( .A0(n44), .A1(n39), .A2(n41), .Z(n6));
Q_INV U365 ( .A(n6), .Z(keybuilder_kdf_stall));
Q_OA21 U366 ( .A0(n16), .A1(n281), .B0(n44), .Z(n7));
Q_NR02 U367 ( .A0(key_tlv_ob_full), .A1(cur_state[2]), .Z(n23));
Q_AN03 U368 ( .A0(n23), .A1(n32), .A2(tlv_sb_data_out_valid), .Z(key_tlv_ob_tlv[83]));
Q_AN02 U369 ( .A0(n44), .A1(cur_state[2]), .Z(n46));
Q_AN02 U370 ( .A0(n46), .A1(n276), .Z(key_tlv_ob_tlv[82]));
Q_AN02 U371 ( .A0(cur_state[2]), .A1(cur_state[1]), .Z(n19));
Q_NR02 U372 ( .A0(cur_state[2]), .A1(cur_state[1]), .Z(n17));
Q_AN02 U373 ( .A0(n17), .A1(tlv_sb_data_out_valid), .Z(n18));
Q_OA21 U374 ( .A0(n19), .A1(n18), .B0(n20), .Z(n21));
Q_NR02 U375 ( .A0(key_tlv_ob_full), .A1(cur_state[0]), .Z(n20));
Q_AN03 U376 ( .A0(tlv_sb_data_out_valid), .A1(n22), .A2(n23), .Z(n8));
Q_AO21 U377 ( .A0(n24), .A1(needs_dek), .B0(n26), .Z(n31));
Q_AN02 U378 ( .A0(n25), .A1(needs_dak), .Z(n26));
Q_AN03 U379 ( .A0(gcm_status_data_out_valid), .A1(n4), .A2(n31), .Z(n28));
Q_AN02 U380 ( .A0(n290), .A1(n276), .Z(n27));
Q_OA21 U381 ( .A0(n28), .A1(n27), .B0(tlv_sb_data_out_valid), .Z(n29));
Q_OA21 U382 ( .A0(n30), .A1(n29), .B0(n44), .Z(n9));
Q_AN02 U383 ( .A0(cur_state[2]), .A1(n276), .Z(n42));
Q_AN03 U384 ( .A0(n39), .A1(n4), .A2(n31), .Z(n34));
Q_AN02 U385 ( .A0(n290), .A1(tlv_sb_data_out_valid), .Z(n33));
Q_AO21 U386 ( .A0(n33), .A1(n32), .B0(n42), .Z(n35));
Q_OA21 U387 ( .A0(n35), .A1(n34), .B0(n44), .Z(n10));
Q_AN03 U388 ( .A0(n44), .A1(n36), .A2(n41), .Z(n11));
Q_AO21 U389 ( .A0(n41), .A1(n36), .B0(n42), .Z(n37));
Q_ND02 U390 ( .A0(n44), .A1(n37), .Z(n38));
Q_AN02 U391 ( .A0(n39), .A1(n5), .Z(n40));
Q_AN03 U392 ( .A0(n44), .A1(n40), .A2(n41), .Z(n12));
Q_AO21 U393 ( .A0(n41), .A1(n40), .B0(n42), .Z(n43));
Q_ND02 U394 ( .A0(n44), .A1(n43), .Z(n45));
Q_AN02 U395 ( .A0(n46), .A1(n277), .Z(n13));
Q_ND02 U396 ( .A0(n46), .A1(n272), .Z(n47));
Q_AN02 U397 ( .A0(n48), .A1(dak_gcm_err), .Z(n49));
Q_OA21 U398 ( .A0(n49), .A1(dek_gcm_err), .B0(n3), .Z(n50));
Q_INV U399 ( .A(n50), .Z(n14));
Q_AN02 U400 ( .A0(n3), .A1(dek_gcm_err), .Z(n15));
Q_XOR2 U401 ( .A0(n21), .A1(key_tlv_ob_tlv[83]), .Z(key_tlv_ob_tlv[65]));
Q_AN02 U402 ( .A0(n6), .A1(n260), .Z(gcm_status_data_out_ack));
Q_MX02 U403 ( .S(n6), .A0(n7), .A1(kdf_keybuilder_valid), .Z(key_tlv_ob_wr));
Q_MX02 U404 ( .S(n8), .A0(n51), .A1(n52), .Z(key_tlv_ob_tlv[63]));
Q_AN03 U405 ( .A0(n10), .A1(kdf_keybuilder_data[7]), .A2(n9), .Z(n51));
Q_MX02 U406 ( .S(n9), .A0(n53), .A1(int_tlv_word0[63]), .Z(n52));
Q_AN02 U407 ( .A0(n244), .A1(tlv_sb_data_out[7]), .Z(n53));
Q_MX02 U408 ( .S(n8), .A0(n54), .A1(n55), .Z(key_tlv_ob_tlv[62]));
Q_AN03 U409 ( .A0(n10), .A1(kdf_keybuilder_data[6]), .A2(n9), .Z(n54));
Q_MX02 U410 ( .S(n9), .A0(n56), .A1(int_tlv_word0[62]), .Z(n55));
Q_AN02 U411 ( .A0(n244), .A1(tlv_sb_data_out[6]), .Z(n56));
Q_MX02 U412 ( .S(n8), .A0(n57), .A1(n58), .Z(key_tlv_ob_tlv[61]));
Q_AN03 U413 ( .A0(n10), .A1(kdf_keybuilder_data[5]), .A2(n9), .Z(n57));
Q_MX02 U414 ( .S(n9), .A0(n59), .A1(int_tlv_word0[61]), .Z(n58));
Q_AN02 U415 ( .A0(n244), .A1(tlv_sb_data_out[5]), .Z(n59));
Q_MX02 U416 ( .S(n8), .A0(n60), .A1(n61), .Z(key_tlv_ob_tlv[60]));
Q_AN03 U417 ( .A0(n10), .A1(kdf_keybuilder_data[4]), .A2(n9), .Z(n60));
Q_MX02 U418 ( .S(n9), .A0(n62), .A1(int_tlv_word0[60]), .Z(n61));
Q_AN02 U419 ( .A0(n244), .A1(tlv_sb_data_out[4]), .Z(n62));
Q_MX02 U420 ( .S(n8), .A0(n63), .A1(n64), .Z(key_tlv_ob_tlv[59]));
Q_AN03 U421 ( .A0(n10), .A1(kdf_keybuilder_data[3]), .A2(n9), .Z(n63));
Q_MX02 U422 ( .S(n9), .A0(n65), .A1(int_tlv_word0[59]), .Z(n64));
Q_AN02 U423 ( .A0(n244), .A1(tlv_sb_data_out[3]), .Z(n65));
Q_MX02 U424 ( .S(n8), .A0(n66), .A1(n67), .Z(key_tlv_ob_tlv[58]));
Q_AN03 U425 ( .A0(n10), .A1(kdf_keybuilder_data[2]), .A2(n9), .Z(n66));
Q_MX02 U426 ( .S(n9), .A0(n68), .A1(int_tlv_word0[58]), .Z(n67));
Q_AN02 U427 ( .A0(n244), .A1(tlv_sb_data_out[2]), .Z(n68));
Q_MX02 U428 ( .S(n8), .A0(n69), .A1(n70), .Z(key_tlv_ob_tlv[57]));
Q_AN03 U429 ( .A0(n10), .A1(kdf_keybuilder_data[1]), .A2(n9), .Z(n69));
Q_MX02 U430 ( .S(n9), .A0(n71), .A1(int_tlv_word0[57]), .Z(n70));
Q_AN02 U431 ( .A0(n244), .A1(tlv_sb_data_out[1]), .Z(n71));
Q_MX02 U432 ( .S(n8), .A0(n72), .A1(n73), .Z(key_tlv_ob_tlv[56]));
Q_AN03 U433 ( .A0(n10), .A1(kdf_keybuilder_data[0]), .A2(n9), .Z(n72));
Q_MX02 U434 ( .S(n9), .A0(n74), .A1(int_tlv_word0[56]), .Z(n73));
Q_AN02 U435 ( .A0(n244), .A1(tlv_sb_data_out[0]), .Z(n74));
Q_MX02 U436 ( .S(n8), .A0(n75), .A1(n76), .Z(key_tlv_ob_tlv[55]));
Q_AN03 U437 ( .A0(n10), .A1(kdf_keybuilder_data[15]), .A2(n9), .Z(n75));
Q_MX02 U438 ( .S(n9), .A0(n77), .A1(tlv_sb_data_out[55]), .Z(n76));
Q_AN02 U439 ( .A0(n244), .A1(tlv_sb_data_out[15]), .Z(n77));
Q_MX02 U440 ( .S(n8), .A0(n78), .A1(n79), .Z(key_tlv_ob_tlv[54]));
Q_AN03 U441 ( .A0(n10), .A1(kdf_keybuilder_data[14]), .A2(n9), .Z(n78));
Q_MX02 U442 ( .S(n9), .A0(n80), .A1(tlv_sb_data_out[54]), .Z(n79));
Q_AN02 U443 ( .A0(n244), .A1(tlv_sb_data_out[14]), .Z(n80));
Q_MX02 U444 ( .S(n8), .A0(n81), .A1(n82), .Z(key_tlv_ob_tlv[53]));
Q_AN03 U445 ( .A0(n10), .A1(kdf_keybuilder_data[13]), .A2(n9), .Z(n81));
Q_MX02 U446 ( .S(n9), .A0(n83), .A1(tlv_sb_data_out[53]), .Z(n82));
Q_AN02 U447 ( .A0(n244), .A1(tlv_sb_data_out[13]), .Z(n83));
Q_MX02 U448 ( .S(n8), .A0(n84), .A1(n85), .Z(key_tlv_ob_tlv[52]));
Q_AN03 U449 ( .A0(n10), .A1(kdf_keybuilder_data[12]), .A2(n9), .Z(n84));
Q_MX02 U450 ( .S(n9), .A0(n86), .A1(tlv_sb_data_out[52]), .Z(n85));
Q_AN02 U451 ( .A0(n244), .A1(tlv_sb_data_out[12]), .Z(n86));
Q_MX02 U452 ( .S(n8), .A0(n87), .A1(n88), .Z(key_tlv_ob_tlv[51]));
Q_AN03 U453 ( .A0(n10), .A1(kdf_keybuilder_data[11]), .A2(n9), .Z(n87));
Q_MX02 U454 ( .S(n9), .A0(n89), .A1(tlv_sb_data_out[51]), .Z(n88));
Q_AN02 U455 ( .A0(n244), .A1(tlv_sb_data_out[11]), .Z(n89));
Q_MX02 U456 ( .S(n8), .A0(n90), .A1(n91), .Z(key_tlv_ob_tlv[50]));
Q_AN03 U457 ( .A0(n10), .A1(kdf_keybuilder_data[10]), .A2(n9), .Z(n90));
Q_MX02 U458 ( .S(n9), .A0(n92), .A1(tlv_sb_data_out[50]), .Z(n91));
Q_AN02 U459 ( .A0(n244), .A1(tlv_sb_data_out[10]), .Z(n92));
Q_MX02 U460 ( .S(n8), .A0(n93), .A1(n94), .Z(key_tlv_ob_tlv[49]));
Q_AN03 U461 ( .A0(n10), .A1(kdf_keybuilder_data[9]), .A2(n9), .Z(n93));
Q_MX02 U462 ( .S(n9), .A0(n95), .A1(tlv_sb_data_out[49]), .Z(n94));
Q_AN02 U463 ( .A0(n244), .A1(tlv_sb_data_out[9]), .Z(n95));
Q_MX02 U464 ( .S(n8), .A0(n96), .A1(n97), .Z(key_tlv_ob_tlv[48]));
Q_AN03 U465 ( .A0(n10), .A1(kdf_keybuilder_data[8]), .A2(n9), .Z(n96));
Q_MX02 U466 ( .S(n9), .A0(n98), .A1(tlv_sb_data_out[48]), .Z(n97));
Q_AN02 U467 ( .A0(n244), .A1(tlv_sb_data_out[8]), .Z(n98));
Q_MX02 U468 ( .S(n8), .A0(n99), .A1(n100), .Z(key_tlv_ob_tlv[47]));
Q_AN03 U469 ( .A0(n10), .A1(kdf_keybuilder_data[23]), .A2(n9), .Z(n99));
Q_MX02 U470 ( .S(n9), .A0(n101), .A1(tlv_sb_data_out[47]), .Z(n100));
Q_AN02 U471 ( .A0(n244), .A1(tlv_sb_data_out[23]), .Z(n101));
Q_MX02 U472 ( .S(n8), .A0(n102), .A1(n103), .Z(key_tlv_ob_tlv[46]));
Q_AN03 U473 ( .A0(n10), .A1(kdf_keybuilder_data[22]), .A2(n9), .Z(n102));
Q_MX02 U474 ( .S(n9), .A0(n104), .A1(tlv_sb_data_out[46]), .Z(n103));
Q_AN02 U475 ( .A0(n244), .A1(tlv_sb_data_out[22]), .Z(n104));
Q_MX02 U476 ( .S(n8), .A0(n105), .A1(n106), .Z(key_tlv_ob_tlv[45]));
Q_AN03 U477 ( .A0(n10), .A1(kdf_keybuilder_data[21]), .A2(n9), .Z(n105));
Q_MX02 U478 ( .S(n9), .A0(n107), .A1(tlv_sb_data_out[45]), .Z(n106));
Q_AN02 U479 ( .A0(n244), .A1(tlv_sb_data_out[21]), .Z(n107));
Q_MX02 U480 ( .S(n8), .A0(n108), .A1(n109), .Z(key_tlv_ob_tlv[44]));
Q_AN03 U481 ( .A0(n10), .A1(kdf_keybuilder_data[20]), .A2(n9), .Z(n108));
Q_MX02 U482 ( .S(n9), .A0(n110), .A1(tlv_sb_data_out[44]), .Z(n109));
Q_AN02 U483 ( .A0(n244), .A1(tlv_sb_data_out[20]), .Z(n110));
Q_MX02 U484 ( .S(n8), .A0(n111), .A1(n112), .Z(key_tlv_ob_tlv[43]));
Q_AN03 U485 ( .A0(n10), .A1(kdf_keybuilder_data[19]), .A2(n9), .Z(n111));
Q_MX02 U486 ( .S(n9), .A0(n113), .A1(tlv_sb_data_out[43]), .Z(n112));
Q_AN02 U487 ( .A0(n244), .A1(tlv_sb_data_out[19]), .Z(n113));
Q_MX02 U488 ( .S(n8), .A0(n114), .A1(n115), .Z(key_tlv_ob_tlv[42]));
Q_AN03 U489 ( .A0(n10), .A1(kdf_keybuilder_data[18]), .A2(n9), .Z(n114));
Q_MX03 U490 ( .S0(n10), .S1(n9), .A0(tlv_sb_data_out[18]), .A1(tlv_sb_data_out[38]), .A2(tlv_sb_data_out[42]), .Z(n115));
Q_MX02 U491 ( .S(n8), .A0(n116), .A1(n117), .Z(key_tlv_ob_tlv[41]));
Q_AN03 U492 ( .A0(n10), .A1(kdf_keybuilder_data[17]), .A2(n9), .Z(n116));
Q_MX03 U493 ( .S0(n10), .S1(n9), .A0(tlv_sb_data_out[17]), .A1(tlv_sb_data_out[37]), .A2(tlv_sb_data_out[41]), .Z(n117));
Q_MX02 U494 ( .S(n8), .A0(n118), .A1(n119), .Z(key_tlv_ob_tlv[40]));
Q_AN03 U495 ( .A0(n10), .A1(kdf_keybuilder_data[16]), .A2(n9), .Z(n118));
Q_MX03 U496 ( .S0(n10), .S1(n9), .A0(tlv_sb_data_out[16]), .A1(tlv_sb_data_out[36]), .A2(tlv_sb_data_out[40]), .Z(n119));
Q_MX02 U497 ( .S(n8), .A0(n120), .A1(n121), .Z(key_tlv_ob_tlv[39]));
Q_AN03 U498 ( .A0(n10), .A1(kdf_keybuilder_data[31]), .A2(n9), .Z(n120));
Q_MX03 U499 ( .S0(n10), .S1(n9), .A0(tlv_sb_data_out[31]), .A1(tlv_sb_data_out[35]), .A2(tlv_sb_data_out[39]), .Z(n121));
Q_MX02 U500 ( .S(n8), .A0(n122), .A1(n123), .Z(key_tlv_ob_tlv[38]));
Q_AN03 U501 ( .A0(n10), .A1(kdf_keybuilder_data[30]), .A2(n9), .Z(n122));
Q_MX03 U502 ( .S0(n10), .S1(n9), .A0(tlv_sb_data_out[30]), .A1(tlv_sb_data_out[34]), .A2(tlv_sb_data_out[38]), .Z(n123));
Q_MX02 U503 ( .S(n8), .A0(n124), .A1(n125), .Z(key_tlv_ob_tlv[37]));
Q_AN03 U504 ( .A0(n10), .A1(kdf_keybuilder_data[29]), .A2(n9), .Z(n124));
Q_MX03 U505 ( .S0(n10), .S1(n9), .A0(tlv_sb_data_out[29]), .A1(tlv_sb_data_out[33]), .A2(tlv_sb_data_out[37]), .Z(n125));
Q_MX02 U506 ( .S(n8), .A0(n126), .A1(n127), .Z(key_tlv_ob_tlv[36]));
Q_AN03 U507 ( .A0(n10), .A1(kdf_keybuilder_data[28]), .A2(n9), .Z(n126));
Q_MX03 U508 ( .S0(n10), .S1(n9), .A0(tlv_sb_data_out[28]), .A1(tlv_sb_data_out[32]), .A2(tlv_sb_data_out[36]), .Z(n127));
Q_MX02 U509 ( .S(n8), .A0(n128), .A1(n129), .Z(key_tlv_ob_tlv[35]));
Q_AN03 U510 ( .A0(n10), .A1(kdf_keybuilder_data[27]), .A2(n9), .Z(n128));
Q_MX03 U511 ( .S0(n10), .S1(n9), .A0(tlv_sb_data_out[27]), .A1(tlv_sb_data_out[31]), .A2(tlv_sb_data_out[35]), .Z(n129));
Q_MX02 U512 ( .S(n8), .A0(n130), .A1(n131), .Z(key_tlv_ob_tlv[34]));
Q_AN03 U513 ( .A0(n10), .A1(kdf_keybuilder_data[26]), .A2(n9), .Z(n130));
Q_MX03 U514 ( .S0(n10), .S1(n9), .A0(tlv_sb_data_out[26]), .A1(tlv_sb_data_out[30]), .A2(tlv_sb_data_out[34]), .Z(n131));
Q_MX02 U515 ( .S(n8), .A0(n132), .A1(n133), .Z(key_tlv_ob_tlv[33]));
Q_AN03 U516 ( .A0(n10), .A1(kdf_keybuilder_data[25]), .A2(n9), .Z(n132));
Q_MX03 U517 ( .S0(n10), .S1(n9), .A0(tlv_sb_data_out[25]), .A1(tlv_sb_data_out[29]), .A2(tlv_sb_data_out[33]), .Z(n133));
Q_MX02 U518 ( .S(n8), .A0(n134), .A1(n135), .Z(key_tlv_ob_tlv[32]));
Q_AN03 U519 ( .A0(n10), .A1(kdf_keybuilder_data[24]), .A2(n9), .Z(n134));
Q_MX03 U520 ( .S0(n10), .S1(n9), .A0(tlv_sb_data_out[24]), .A1(tlv_sb_data_out[28]), .A2(tlv_sb_data_out[32]), .Z(n135));
Q_MX02 U521 ( .S(n8), .A0(n136), .A1(n138), .Z(key_tlv_ob_tlv[31]));
Q_AN02 U522 ( .A0(n10), .A1(n137), .Z(n136));
Q_MX02 U523 ( .S(n9), .A0(crc[31]), .A1(kdf_keybuilder_data[39]), .Z(n137));
Q_MX02 U524 ( .S(n9), .A0(n139), .A1(tlv_sb_data_out[31]), .Z(n138));
Q_AN02 U525 ( .A0(n244), .A1(tlv_sb_data_out[39]), .Z(n139));
Q_MX02 U526 ( .S(n8), .A0(n140), .A1(n142), .Z(key_tlv_ob_tlv[30]));
Q_AN02 U527 ( .A0(n10), .A1(n141), .Z(n140));
Q_MX02 U528 ( .S(n9), .A0(crc[30]), .A1(kdf_keybuilder_data[38]), .Z(n141));
Q_MX02 U529 ( .S(n9), .A0(n143), .A1(tlv_sb_data_out[30]), .Z(n142));
Q_AN02 U530 ( .A0(n244), .A1(tlv_sb_data_out[38]), .Z(n143));
Q_MX02 U531 ( .S(n8), .A0(n144), .A1(n146), .Z(key_tlv_ob_tlv[29]));
Q_AN02 U532 ( .A0(n10), .A1(n145), .Z(n144));
Q_MX02 U533 ( .S(n9), .A0(crc[29]), .A1(kdf_keybuilder_data[37]), .Z(n145));
Q_MX02 U534 ( .S(n9), .A0(n147), .A1(tlv_sb_data_out[29]), .Z(n146));
Q_AN02 U535 ( .A0(n244), .A1(tlv_sb_data_out[37]), .Z(n147));
Q_MX02 U536 ( .S(n8), .A0(n148), .A1(n150), .Z(key_tlv_ob_tlv[28]));
Q_AN02 U537 ( .A0(n10), .A1(n149), .Z(n148));
Q_MX02 U538 ( .S(n9), .A0(crc[28]), .A1(kdf_keybuilder_data[36]), .Z(n149));
Q_MX02 U539 ( .S(n9), .A0(n151), .A1(tlv_sb_data_out[28]), .Z(n150));
Q_AN02 U540 ( .A0(n244), .A1(tlv_sb_data_out[36]), .Z(n151));
Q_MX02 U541 ( .S(n8), .A0(n152), .A1(n154), .Z(key_tlv_ob_tlv[27]));
Q_AN02 U542 ( .A0(n10), .A1(n153), .Z(n152));
Q_MX02 U543 ( .S(n9), .A0(crc[27]), .A1(kdf_keybuilder_data[35]), .Z(n153));
Q_MX02 U544 ( .S(n316), .A0(tlv_sb_data_out[35]), .A1(tlv_sb_data_out[27]), .Z(n154));
Q_MX02 U545 ( .S(n8), .A0(n155), .A1(n157), .Z(key_tlv_ob_tlv[26]));
Q_AN02 U546 ( .A0(n10), .A1(n156), .Z(n155));
Q_MX02 U547 ( .S(n9), .A0(crc[26]), .A1(kdf_keybuilder_data[34]), .Z(n156));
Q_MX02 U548 ( .S(n316), .A0(tlv_sb_data_out[34]), .A1(tlv_sb_data_out[26]), .Z(n157));
Q_MX02 U549 ( .S(n8), .A0(n158), .A1(n160), .Z(key_tlv_ob_tlv[25]));
Q_AN02 U550 ( .A0(n10), .A1(n159), .Z(n158));
Q_MX02 U551 ( .S(n9), .A0(crc[25]), .A1(kdf_keybuilder_data[33]), .Z(n159));
Q_MX02 U552 ( .S(n316), .A0(tlv_sb_data_out[33]), .A1(tlv_sb_data_out[25]), .Z(n160));
Q_MX02 U553 ( .S(n8), .A0(n161), .A1(n163), .Z(key_tlv_ob_tlv[24]));
Q_AN02 U554 ( .A0(n10), .A1(n162), .Z(n161));
Q_MX02 U555 ( .S(n9), .A0(crc[24]), .A1(kdf_keybuilder_data[32]), .Z(n162));
Q_MX02 U556 ( .S(n316), .A0(tlv_sb_data_out[32]), .A1(tlv_sb_data_out[24]), .Z(n163));
Q_MX02 U557 ( .S(n8), .A0(n164), .A1(n166), .Z(key_tlv_ob_tlv[23]));
Q_AN02 U558 ( .A0(n10), .A1(n165), .Z(n164));
Q_MX02 U559 ( .S(n9), .A0(crc[23]), .A1(kdf_keybuilder_data[47]), .Z(n165));
Q_MX02 U560 ( .S(n316), .A0(tlv_sb_data_out[47]), .A1(tlv_sb_data_out[23]), .Z(n166));
Q_MX02 U561 ( .S(n8), .A0(n167), .A1(n169), .Z(key_tlv_ob_tlv[22]));
Q_AN02 U562 ( .A0(n10), .A1(n168), .Z(n167));
Q_MX02 U563 ( .S(n9), .A0(crc[22]), .A1(kdf_keybuilder_data[46]), .Z(n168));
Q_MX02 U564 ( .S(n316), .A0(tlv_sb_data_out[46]), .A1(tlv_sb_data_out[22]), .Z(n169));
Q_MX02 U565 ( .S(n8), .A0(n170), .A1(n172), .Z(key_tlv_ob_tlv[21]));
Q_AN02 U566 ( .A0(n10), .A1(n171), .Z(n170));
Q_MX02 U567 ( .S(n9), .A0(crc[21]), .A1(kdf_keybuilder_data[45]), .Z(n171));
Q_MX02 U568 ( .S(n316), .A0(tlv_sb_data_out[45]), .A1(tlv_sb_data_out[21]), .Z(n172));
Q_MX02 U569 ( .S(n8), .A0(n173), .A1(n175), .Z(key_tlv_ob_tlv[20]));
Q_AN02 U570 ( .A0(n10), .A1(n174), .Z(n173));
Q_MX02 U571 ( .S(n9), .A0(crc[20]), .A1(kdf_keybuilder_data[44]), .Z(n174));
Q_MX02 U572 ( .S(n316), .A0(tlv_sb_data_out[44]), .A1(tlv_sb_data_out[20]), .Z(n175));
Q_MX02 U573 ( .S(n8), .A0(n176), .A1(n178), .Z(key_tlv_ob_tlv[19]));
Q_AN02 U574 ( .A0(n10), .A1(n177), .Z(n176));
Q_MX02 U575 ( .S(n9), .A0(crc[19]), .A1(kdf_keybuilder_data[43]), .Z(n177));
Q_MX02 U576 ( .S(n316), .A0(tlv_sb_data_out[43]), .A1(tlv_sb_data_out[19]), .Z(n178));
Q_MX02 U577 ( .S(n8), .A0(n179), .A1(n181), .Z(key_tlv_ob_tlv[18]));
Q_AN02 U578 ( .A0(n10), .A1(n180), .Z(n179));
Q_MX02 U579 ( .S(n9), .A0(crc[18]), .A1(kdf_keybuilder_data[42]), .Z(n180));
Q_MX02 U580 ( .S(n316), .A0(tlv_sb_data_out[42]), .A1(tlv_sb_data_out[18]), .Z(n181));
Q_MX02 U581 ( .S(n8), .A0(n182), .A1(n184), .Z(key_tlv_ob_tlv[17]));
Q_AN02 U582 ( .A0(n10), .A1(n183), .Z(n182));
Q_MX02 U583 ( .S(n9), .A0(crc[17]), .A1(kdf_keybuilder_data[41]), .Z(n183));
Q_MX02 U584 ( .S(n316), .A0(tlv_sb_data_out[41]), .A1(tlv_sb_data_out[17]), .Z(n184));
Q_MX02 U585 ( .S(n8), .A0(n185), .A1(n187), .Z(key_tlv_ob_tlv[16]));
Q_AN02 U586 ( .A0(n10), .A1(n186), .Z(n185));
Q_MX02 U587 ( .S(n9), .A0(crc[16]), .A1(kdf_keybuilder_data[40]), .Z(n186));
Q_MX02 U588 ( .S(n316), .A0(tlv_sb_data_out[40]), .A1(tlv_sb_data_out[16]), .Z(n187));
Q_MX02 U589 ( .S(n8), .A0(n188), .A1(n190), .Z(key_tlv_ob_tlv[15]));
Q_AN02 U590 ( .A0(n10), .A1(n189), .Z(n188));
Q_MX02 U591 ( .S(n9), .A0(crc[15]), .A1(kdf_keybuilder_data[55]), .Z(n189));
Q_MX02 U592 ( .S(n9), .A0(n191), .A1(tlv_sb_data_out[15]), .Z(n190));
Q_OR02 U593 ( .A0(n10), .A1(tlv_sb_data_out[55]), .Z(n191));
Q_MX02 U594 ( .S(n8), .A0(n192), .A1(n194), .Z(key_tlv_ob_tlv[14]));
Q_AN02 U595 ( .A0(n10), .A1(n193), .Z(n192));
Q_MX02 U596 ( .S(n9), .A0(crc[14]), .A1(kdf_keybuilder_data[54]), .Z(n193));
Q_MX02 U597 ( .S(n9), .A0(n195), .A1(tlv_sb_data_out[14]), .Z(n194));
Q_AN02 U598 ( .A0(n244), .A1(tlv_sb_data_out[54]), .Z(n195));
Q_MX02 U599 ( .S(n8), .A0(n196), .A1(n198), .Z(key_tlv_ob_tlv[13]));
Q_AN02 U600 ( .A0(n10), .A1(n197), .Z(n196));
Q_MX02 U601 ( .S(n9), .A0(crc[13]), .A1(kdf_keybuilder_data[53]), .Z(n197));
Q_MX02 U602 ( .S(n9), .A0(n199), .A1(tlv_sb_data_out[13]), .Z(n198));
Q_OR02 U603 ( .A0(n10), .A1(tlv_sb_data_out[53]), .Z(n199));
Q_MX02 U604 ( .S(n8), .A0(n200), .A1(n202), .Z(key_tlv_ob_tlv[12]));
Q_AN02 U605 ( .A0(n10), .A1(n201), .Z(n200));
Q_MX02 U606 ( .S(n9), .A0(crc[12]), .A1(kdf_keybuilder_data[52]), .Z(n201));
Q_MX02 U607 ( .S(n9), .A0(n203), .A1(tlv_sb_data_out[12]), .Z(n202));
Q_AN02 U608 ( .A0(n244), .A1(tlv_sb_data_out[52]), .Z(n203));
Q_MX02 U609 ( .S(n8), .A0(n204), .A1(n206), .Z(key_tlv_ob_tlv[11]));
Q_AN02 U610 ( .A0(n10), .A1(n205), .Z(n204));
Q_MX02 U611 ( .S(n9), .A0(crc[11]), .A1(kdf_keybuilder_data[51]), .Z(n205));
Q_MX02 U612 ( .S(n9), .A0(n207), .A1(tlv_sb_data_out[11]), .Z(n206));
Q_OR02 U613 ( .A0(n10), .A1(tlv_sb_data_out[51]), .Z(n207));
Q_MX02 U614 ( .S(n8), .A0(n208), .A1(n210), .Z(key_tlv_ob_tlv[10]));
Q_AN02 U615 ( .A0(n10), .A1(n209), .Z(n208));
Q_MX02 U616 ( .S(n9), .A0(crc[10]), .A1(kdf_keybuilder_data[50]), .Z(n209));
Q_MX02 U617 ( .S(n9), .A0(n211), .A1(tlv_sb_data_out[10]), .Z(n210));
Q_AN02 U618 ( .A0(n244), .A1(tlv_sb_data_out[50]), .Z(n211));
Q_MX02 U619 ( .S(n8), .A0(n212), .A1(n214), .Z(key_tlv_ob_tlv[9]));
Q_AN02 U620 ( .A0(n10), .A1(n213), .Z(n212));
Q_MX02 U621 ( .S(n9), .A0(crc[9]), .A1(kdf_keybuilder_data[49]), .Z(n213));
Q_MX02 U622 ( .S(n9), .A0(n215), .A1(tlv_sb_data_out[9]), .Z(n214));
Q_AN02 U623 ( .A0(n244), .A1(tlv_sb_data_out[49]), .Z(n215));
Q_MX02 U624 ( .S(n8), .A0(n216), .A1(n218), .Z(key_tlv_ob_tlv[8]));
Q_AN02 U625 ( .A0(n10), .A1(n217), .Z(n216));
Q_MX02 U626 ( .S(n9), .A0(crc[8]), .A1(kdf_keybuilder_data[48]), .Z(n217));
Q_MX02 U627 ( .S(n9), .A0(n219), .A1(tlv_sb_data_out[8]), .Z(n218));
Q_AN02 U628 ( .A0(n244), .A1(tlv_sb_data_out[48]), .Z(n219));
Q_MX04 U629 ( .S0(n9), .S1(n8), .A0(n220), .A1(n221), .A2(n222), .A3(tlv_sb_data_out[7]), .Z(key_tlv_ob_tlv[7]));
Q_AN02 U630 ( .A0(n10), .A1(crc[7]), .Z(n220));
Q_MX02 U631 ( .S(n10), .A0(n248), .A1(kdf_keybuilder_data[63]), .Z(n221));
Q_AN02 U632 ( .A0(n244), .A1(int_tlv_word0[63]), .Z(n222));
Q_MX04 U633 ( .S0(n9), .S1(n8), .A0(n223), .A1(n224), .A2(n225), .A3(tlv_sb_data_out[6]), .Z(key_tlv_ob_tlv[6]));
Q_AN02 U634 ( .A0(n10), .A1(crc[6]), .Z(n223));
Q_MX02 U635 ( .S(n10), .A0(n249), .A1(kdf_keybuilder_data[62]), .Z(n224));
Q_AN02 U636 ( .A0(n244), .A1(int_tlv_word0[62]), .Z(n225));
Q_MX04 U637 ( .S0(n9), .S1(n8), .A0(n226), .A1(n227), .A2(n228), .A3(tlv_sb_data_out[5]), .Z(key_tlv_ob_tlv[5]));
Q_AN02 U638 ( .A0(n10), .A1(crc[5]), .Z(n226));
Q_MX02 U639 ( .S(n10), .A0(n250), .A1(kdf_keybuilder_data[61]), .Z(n227));
Q_AN02 U640 ( .A0(n244), .A1(int_tlv_word0[61]), .Z(n228));
Q_MX04 U641 ( .S0(n9), .S1(n8), .A0(n229), .A1(n230), .A2(n231), .A3(tlv_sb_data_out[4]), .Z(key_tlv_ob_tlv[4]));
Q_AN02 U642 ( .A0(n10), .A1(crc[4]), .Z(n229));
Q_MX02 U643 ( .S(n10), .A0(n251), .A1(kdf_keybuilder_data[60]), .Z(n230));
Q_AN02 U644 ( .A0(n244), .A1(int_tlv_word0[60]), .Z(n231));
Q_MX04 U645 ( .S0(n9), .S1(n8), .A0(n232), .A1(n233), .A2(n234), .A3(tlv_sb_data_out[3]), .Z(key_tlv_ob_tlv[3]));
Q_AN02 U646 ( .A0(n10), .A1(crc[3]), .Z(n232));
Q_MX02 U647 ( .S(n10), .A0(n252), .A1(kdf_keybuilder_data[59]), .Z(n233));
Q_AN02 U648 ( .A0(n244), .A1(int_tlv_word0[59]), .Z(n234));
Q_MX04 U649 ( .S0(n9), .S1(n8), .A0(n235), .A1(n236), .A2(n237), .A3(tlv_sb_data_out[2]), .Z(key_tlv_ob_tlv[2]));
Q_AN02 U650 ( .A0(n10), .A1(crc[2]), .Z(n235));
Q_MX02 U651 ( .S(n10), .A0(n254), .A1(kdf_keybuilder_data[58]), .Z(n236));
Q_AN02 U652 ( .A0(n244), .A1(int_tlv_word0[58]), .Z(n237));
Q_MX04 U653 ( .S0(n9), .S1(n8), .A0(n238), .A1(n239), .A2(n240), .A3(tlv_sb_data_out[1]), .Z(key_tlv_ob_tlv[1]));
Q_AN02 U654 ( .A0(n10), .A1(crc[1]), .Z(n238));
Q_MX02 U655 ( .S(n10), .A0(n255), .A1(kdf_keybuilder_data[57]), .Z(n239));
Q_OR02 U656 ( .A0(n10), .A1(int_tlv_word0[57]), .Z(n240));
Q_MX04 U657 ( .S0(n9), .S1(n8), .A0(n241), .A1(n242), .A2(n243), .A3(tlv_sb_data_out[0]), .Z(key_tlv_ob_tlv[0]));
Q_AN02 U658 ( .A0(n10), .A1(n257), .Z(n241));
Q_MX02 U659 ( .S(n10), .A0(n256), .A1(kdf_keybuilder_data[56]), .Z(n242));
Q_AN02 U660 ( .A0(n244), .A1(int_tlv_word0[56]), .Z(n243));
Q_INV U661 ( .A(n10), .Z(n244));
Q_MX02 U662 ( .S(n11), .A0(n245), .A1(gcm_status_data_out[0]), .Z(nxt_dek_gcm_err));
Q_AN02 U663 ( .A0(n38), .A1(dek_gcm_err), .Z(n245));
Q_MX02 U664 ( .S(n12), .A0(n246), .A1(gcm_status_data_out[0]), .Z(nxt_dak_gcm_err));
Q_AN02 U665 ( .A0(n45), .A1(dak_gcm_err), .Z(n246));
Q_MX02 U666 ( .S(n13), .A0(n247), .A1(tlv_sb_data_out[55]), .Z(nxt_corrupt_crc));
Q_AN02 U667 ( .A0(n47), .A1(corrupt_crc), .Z(n247));
Q_MX02 U668 ( .S(key_tlv_ob_tlv[83]), .A0(needs_dek), .A1(tlv_sb_data_out[46]), .Z(nxt_needs_dek));
Q_MX02 U669 ( .S(key_tlv_ob_tlv[83]), .A0(needs_dak), .A1(tlv_sb_data_out[45]), .Z(nxt_needs_dak));
Q_AN02 U670 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[31]), .Z(key_tlv_word20[31]));
Q_AN02 U671 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[30]), .Z(key_tlv_word20[30]));
Q_AN02 U672 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[29]), .Z(key_tlv_word20[29]));
Q_AN02 U673 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[28]), .Z(key_tlv_word20[28]));
Q_AN02 U674 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[27]), .Z(key_tlv_word20[27]));
Q_AN02 U675 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[26]), .Z(key_tlv_word20[26]));
Q_AN02 U676 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[25]), .Z(key_tlv_word20[25]));
Q_AN02 U677 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[24]), .Z(key_tlv_word20[24]));
Q_AN02 U678 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[23]), .Z(key_tlv_word20[23]));
Q_AN02 U679 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[22]), .Z(key_tlv_word20[22]));
Q_AN02 U680 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[21]), .Z(key_tlv_word20[21]));
Q_AN02 U681 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[20]), .Z(key_tlv_word20[20]));
Q_AN02 U682 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[19]), .Z(key_tlv_word20[19]));
Q_AN02 U683 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[18]), .Z(key_tlv_word20[18]));
Q_AN02 U684 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[17]), .Z(key_tlv_word20[17]));
Q_AN02 U685 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[16]), .Z(key_tlv_word20[16]));
Q_AN02 U686 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[15]), .Z(key_tlv_word20[15]));
Q_AN02 U687 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[14]), .Z(key_tlv_word20[14]));
Q_AN02 U688 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[13]), .Z(key_tlv_word20[13]));
Q_AN02 U689 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[12]), .Z(key_tlv_word20[12]));
Q_AN02 U690 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[11]), .Z(key_tlv_word20[11]));
Q_AN02 U691 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[10]), .Z(key_tlv_word20[10]));
Q_AN02 U692 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[9]), .Z(key_tlv_word20[9]));
Q_AN02 U693 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[8]), .Z(key_tlv_word20[8]));
Q_AN02 U694 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[7]), .Z(key_tlv_word20[7]));
Q_AN02 U695 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[6]), .Z(key_tlv_word20[6]));
Q_AN02 U696 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[5]), .Z(key_tlv_word20[5]));
Q_AN02 U697 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[4]), .Z(key_tlv_word20[4]));
Q_AN02 U698 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[3]), .Z(key_tlv_word20[3]));
Q_AN02 U699 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[2]), .Z(key_tlv_word20[2]));
Q_AN02 U700 ( .A0(key_tlv_ob_tlv[82]), .A1(crc[1]), .Z(key_tlv_word20[1]));
Q_AN02 U701 ( .A0(key_tlv_ob_tlv[82]), .A1(n257), .Z(key_tlv_word20[0]));
Q_AN02 U702 ( .A0(n13), .A1(n248), .Z(key_tlv_word19[7]));
Q_AN02 U703 ( .A0(n13), .A1(n249), .Z(key_tlv_word19[6]));
Q_AN02 U704 ( .A0(n13), .A1(n250), .Z(key_tlv_word19[5]));
Q_AN02 U705 ( .A0(n13), .A1(n251), .Z(key_tlv_word19[4]));
Q_AN02 U706 ( .A0(n13), .A1(n252), .Z(key_tlv_word19[3]));
Q_AN02 U707 ( .A0(n13), .A1(n254), .Z(key_tlv_word19[2]));
Q_AN02 U708 ( .A0(n13), .A1(n255), .Z(key_tlv_word19[1]));
Q_AN02 U709 ( .A0(n13), .A1(n256), .Z(key_tlv_word19[0]));
Q_OR02 U710 ( .A0(n50), .A1(tlv_sb_data_out[7]), .Z(n248));
Q_AN02 U711 ( .A0(n14), .A1(tlv_sb_data_out[6]), .Z(n249));
Q_AN02 U712 ( .A0(n14), .A1(tlv_sb_data_out[5]), .Z(n250));
Q_AN02 U713 ( .A0(n14), .A1(tlv_sb_data_out[4]), .Z(n251));
Q_MX02 U714 ( .S(n50), .A0(tlv_sb_data_out[3]), .A1(n253), .Z(n252));
Q_INV U715 ( .A(n15), .Z(n253));
Q_MX02 U716 ( .S(n50), .A0(tlv_sb_data_out[2]), .A1(n15), .Z(n254));
Q_MX02 U717 ( .S(n50), .A0(tlv_sb_data_out[1]), .A1(n15), .Z(n255));
Q_MX02 U718 ( .S(n50), .A0(tlv_sb_data_out[0]), .A1(n15), .Z(n256));
Q_XOR2 U719 ( .A0(crc[0]), .A1(corrupt_crc), .Z(n257));
Q_NR02 U720 ( .A0(n258), .A1(n301), .Z(n5));
Q_OR03 U721 ( .A0(cur_state[0]), .A1(cur_state[1]), .A2(n290), .Z(n258));
Q_AN03 U722 ( .A0(n259), .A1(n260), .A2(n39), .Z(n36));
Q_AN03 U723 ( .A0(cur_state[0]), .A1(cur_state[1]), .A2(n290), .Z(n259));
Q_INV U724 ( .A(n301), .Z(n260));
Q_NR02 U725 ( .A0(n261), .A1(gcm_status_data_out[0]), .Z(n4));
Q_INV U726 ( .A(n261), .Z(n3));
Q_OR02 U727 ( .A0(n263), .A1(n262), .Z(n261));
Q_OR03 U728 ( .A0(tlv_sb_data_out[1]), .A1(tlv_sb_data_out[0]), .A2(n264), .Z(n262));
Q_OR03 U729 ( .A0(tlv_sb_data_out[4]), .A1(tlv_sb_data_out[3]), .A2(tlv_sb_data_out[2]), .Z(n263));
Q_OR03 U730 ( .A0(tlv_sb_data_out[7]), .A1(tlv_sb_data_out[6]), .A2(tlv_sb_data_out[5]), .Z(n264));
Q_AN02 U731 ( .A0(cur_state[1]), .A1(n292), .Z(n276));
Q_AN02 U732 ( .A0(n288), .A1(cur_state[0]), .Z(n277));
Q_OR02 U733 ( .A0(n276), .A1(n277), .Z(n272));
Q_AN03 U734 ( .A0(cur_state[2]), .A1(n288), .A2(n268), .Z(n271));
Q_NR02 U735 ( .A0(cur_state[0]), .A1(key_tlv_beat_num[2]), .Z(n268));
Q_AN03 U736 ( .A0(n290), .A1(cur_state[1]), .A2(n269), .Z(n270));
Q_AN02 U737 ( .A0(cur_state[0]), .A1(key_tlv_beat_num[2]), .Z(n269));
Q_OA21 U738 ( .A0(n271), .A1(n270), .B0(n273), .Z(n274));
Q_AN02 U739 ( .A0(n272), .A1(cur_state[2]), .Z(n281));
Q_AN02 U740 ( .A0(key_tlv_beat_num[1]), .A1(key_tlv_beat_num[0]), .Z(n273));
Q_OA21 U741 ( .A0(n281), .A1(n274), .B0(key_tlv_ob_wr), .Z(n275));
Q_INV U742 ( .A(n275), .Z(n265));
Q_MX02 U743 ( .S(key_tlv_beat_num[1]), .A0(n276), .A1(n277), .Z(n279));
Q_AN02 U744 ( .A0(n285), .A1(key_tlv_beat_num[0]), .Z(n278));
Q_AN03 U745 ( .A0(n290), .A1(n278), .A2(n279), .Z(n280));
Q_OA21 U746 ( .A0(n281), .A1(n280), .B0(key_tlv_ob_wr), .Z(n282));
Q_INV U747 ( .A(n282), .Z(n266));
Q_AN02 U748 ( .A0(n285), .A1(key_tlv_beat_num[1]), .Z(n284));
Q_AN02 U749 ( .A0(n288), .A1(key_tlv_beat_num[0]), .Z(n283));
Q_AO21 U750 ( .A0(n284), .A1(n283), .B0(cur_state[1]), .Z(n289));
Q_NR02 U751 ( .A0(key_tlv_beat_num[2]), .A1(key_tlv_beat_num[1]), .Z(n287));
Q_AN02 U752 ( .A0(cur_state[1]), .A1(key_tlv_beat_num[0]), .Z(n286));
Q_AO21 U753 ( .A0(n287), .A1(n286), .B0(n288), .Z(n291));
Q_MX02 U754 ( .S(cur_state[2]), .A0(n291), .A1(n289), .Z(n293));
Q_AN03 U755 ( .A0(n292), .A1(key_tlv_ob_wr), .A2(n293), .Z(n294));
Q_INV U756 ( .A(n294), .Z(n267));
Q_AN02 U757 ( .A0(n296), .A1(cur_state[0]), .Z(n295));
Q_AO21 U758 ( .A0(n296), .A1(cur_state[1]), .B0(n299), .Z(nxt_state[1]));
Q_AO21 U759 ( .A0(n296), .A1(cur_state[2]), .B0(n298), .Z(nxt_state[2]));
Q_NR02 U760 ( .A0(n282), .A1(n275), .Z(n297));
Q_AN02 U761 ( .A0(n267), .A1(n297), .Z(n296));
Q_NR02 U762 ( .A0(n2), .A1(n265), .Z(n298));
Q_NR02 U763 ( .A0(n266), .A1(n1), .Z(n299));
Q_ND02 U764 ( .A0(n282), .A1(n275), .Z(n300));
Q_AO21 U765 ( .A0(n294), .A1(n300), .B0(n295), .Z(nxt_state[0]));
Q_INV U766 ( .A(key_tlv_ob_wr), .Z(n302));
Q_ND02 U767 ( .A0(n301), .A1(n302), .Z(n303));
Q_AN02 U768 ( .A0(n301), .A1(n307), .Z(n304));
Q_AN02 U769 ( .A0(n301), .A1(n308), .Z(n305));
Q_AN02 U770 ( .A0(n301), .A1(n309), .Z(n306));
Q_XOR2 U771 ( .A0(key_tlv_beat_num[2]), .A1(n273), .Z(n307));
Q_AN03 U772 ( .A0(n312), .A1(n311), .A2(n310), .Z(n301));
Q_XNR2 U773 ( .A0(cur_state[2]), .A1(nxt_state[2]), .Z(n310));
Q_XNR2 U774 ( .A0(cur_state[1]), .A1(nxt_state[1]), .Z(n311));
Q_XNR2 U775 ( .A0(cur_state[0]), .A1(nxt_state[0]), .Z(n312));
Q_FDP1 needs_dak_REG  ( .CK(clk), .R(rst_n), .D(nxt_needs_dak), .Q(needs_dak), .QN( ));
Q_FDP1 needs_dek_REG  ( .CK(clk), .R(rst_n), .D(nxt_needs_dek), .Q(needs_dek), .QN( ));
Q_FDP1 corrupt_crc_REG  ( .CK(clk), .R(rst_n), .D(nxt_corrupt_crc), .Q(corrupt_crc), .QN( ));
Q_FDP1 dak_gcm_err_REG  ( .CK(clk), .R(rst_n), .D(nxt_dak_gcm_err), .Q(dak_gcm_err), .QN( ));
Q_FDP1 dek_gcm_err_REG  ( .CK(clk), .R(rst_n), .D(nxt_dek_gcm_err), .Q(dek_gcm_err), .QN(n48));
Q_FDP1 \cur_state_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_state[0]), .Q(cur_state[0]), .QN(n292));
Q_FDP1 \cur_state_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_state[1]), .Q(cur_state[1]), .QN(n288));
Q_FDP1 \cur_state_REG[2] ( .CK(clk), .R(rst_n), .D(nxt_state[2]), .Q(cur_state[2]), .QN(n290));
Q_AN02 U784 ( .A0(key_tlv_ob_wr), .A1(key_tlv_ob_tlv[83]), .Z(init));
Q_NR02 U785 ( .A0(key_tlv_ob_tlv[83]), .A1(key_tlv_ob_tlv[82]), .Z(n313));
Q_AN02 U786 ( .A0(key_tlv_ob_wr), .A1(n313), .Z(data_valid));
ixc_assign _zz_strnp_0 ( _zy_simnet_tlv_sb_data_out_ack_0_w$, 
	tlv_sb_data_out_ack);
ixc_assign _zz_strnp_1 ( _zy_simnet_keybuilder_kdf_stall_1_w$, 
	keybuilder_kdf_stall);
ixc_assign _zz_strnp_2 ( _zy_simnet_gcm_status_data_out_ack_2_w$, 
	gcm_status_data_out_ack);
ixc_assign _zz_strnp_3 ( _zy_simnet_key_tlv_ob_wr_3_w$, key_tlv_ob_wr);
ixc_assign_106 _zz_strnp_4 ( _zy_simnet_key_tlv_ob_tlv_4_w$[0:105], { n314, 
	n314, n314, n314, n314, n314, n314, n314, n314, n314, n314, n314, 
	n314, n314, n314, n314, n314, n314, n314, n314, n315, n314, 
	key_tlv_ob_tlv[83], key_tlv_ob_tlv[82], n314, n314, n315, n315, n315, 
	n315, n315, n315, n315, n315, n314, n314, n314, n314, n314, n314, 
	key_tlv_ob_tlv[65], key_tlv_ob_tlv[83], key_tlv_ob_tlv[63], 
	key_tlv_ob_tlv[62], key_tlv_ob_tlv[61], key_tlv_ob_tlv[60], 
	key_tlv_ob_tlv[59], key_tlv_ob_tlv[58], key_tlv_ob_tlv[57], 
	key_tlv_ob_tlv[56], key_tlv_ob_tlv[55], key_tlv_ob_tlv[54], 
	key_tlv_ob_tlv[53], key_tlv_ob_tlv[52], key_tlv_ob_tlv[51], 
	key_tlv_ob_tlv[50], key_tlv_ob_tlv[49], key_tlv_ob_tlv[48], 
	key_tlv_ob_tlv[47], key_tlv_ob_tlv[46], key_tlv_ob_tlv[45], 
	key_tlv_ob_tlv[44], key_tlv_ob_tlv[43], key_tlv_ob_tlv[42], 
	key_tlv_ob_tlv[41], key_tlv_ob_tlv[40], key_tlv_ob_tlv[39], 
	key_tlv_ob_tlv[38], key_tlv_ob_tlv[37], key_tlv_ob_tlv[36], 
	key_tlv_ob_tlv[35], key_tlv_ob_tlv[34], key_tlv_ob_tlv[33], 
	key_tlv_ob_tlv[32], key_tlv_ob_tlv[31], key_tlv_ob_tlv[30], 
	key_tlv_ob_tlv[29], key_tlv_ob_tlv[28], key_tlv_ob_tlv[27], 
	key_tlv_ob_tlv[26], key_tlv_ob_tlv[25], key_tlv_ob_tlv[24], 
	key_tlv_ob_tlv[23], key_tlv_ob_tlv[22], key_tlv_ob_tlv[21], 
	key_tlv_ob_tlv[20], key_tlv_ob_tlv[19], key_tlv_ob_tlv[18], 
	key_tlv_ob_tlv[17], key_tlv_ob_tlv[16], key_tlv_ob_tlv[15], 
	key_tlv_ob_tlv[14], key_tlv_ob_tlv[13], key_tlv_ob_tlv[12], 
	key_tlv_ob_tlv[11], key_tlv_ob_tlv[10], key_tlv_ob_tlv[9], 
	key_tlv_ob_tlv[8], key_tlv_ob_tlv[7], key_tlv_ob_tlv[6], 
	key_tlv_ob_tlv[5], key_tlv_ob_tlv[4], key_tlv_ob_tlv[3], 
	key_tlv_ob_tlv[2], key_tlv_ob_tlv[1], key_tlv_ob_tlv[0]});
ixc_assign_64 _zz_strnp_5 ( _zy_simnet_key_tlv_ob_tlv_5_w$[0:63], 
	key_tlv_ob_tlv[63:0]);
cr_crc crc32 ( .crc( crc[31:0]), .clk( clk), .rst_n( rst_n), .data_in( 
	_zy_simnet_key_tlv_ob_tlv_5_w$[0:63]), .data_valid( data_valid), 
	.data_vbytes( _zy_simnet_cio_6[0:7]), .enable( _zy_simnet_cio_7), 
	.init_value( _zy_simnet_cio_8[0:31]), .init( init));
Q_OR02 U794 ( .A0(n10), .A1(n9), .Z(n316));
Q_XOR2 U795 ( .A0(key_tlv_beat_num[1]), .A1(key_tlv_beat_num[0]), .Z(n308));
Q_FDP4EP \key_tlv_beat_num_REG[2] ( .CK(clk), .CE(n303), .R(n317), .D(n304), .Q(key_tlv_beat_num[2]));
Q_INV U797 ( .A(rst_n), .Z(n317));
Q_INV U798 ( .A(key_tlv_beat_num[2]), .Z(n285));
Q_FDP4EP \key_tlv_beat_num_REG[1] ( .CK(clk), .CE(n303), .R(n317), .D(n305), .Q(key_tlv_beat_num[1]));
Q_FDP4EP \key_tlv_beat_num_REG[0] ( .CK(clk), .CE(n303), .R(n317), .D(n306), .Q(key_tlv_beat_num[0]));
Q_INV U801 ( .A(key_tlv_beat_num[0]), .Z(n309));
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "\key_tlv_ob_tlv.ordern  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m2 "\key_tlv_ob_tlv.typen  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m3 "\key_tlv_ob_tlv.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m4 "\key_tlv_ob_tlv.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m5 "\key_tlv_ob_tlv.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m6 "\key_tlv_ob_tlv.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m7 "\gcm_status_data_out.tag_mismatch  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m8 "\key_tlv_word0.tlv_bip2  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m9 "\key_tlv_word0.resv0  (1,0) 1 18 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m10 "\key_tlv_word0.tlv_frame_num  (1,0) 1 10 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m11 "\key_tlv_word0.resv1  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m12 "\key_tlv_word0.tlv_eng_id  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m13 "\key_tlv_word0.tlv_seq_num  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m14 "\key_tlv_word0.tlv_len  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m15 "\key_tlv_word0.tlv_type  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m16 "\key_tlv_word19.rsvd  (1,0) 1 55 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m17 "\key_tlv_word19.kme_errors  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m18 "\key_tlv_word20.rsvd  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m19 "\key_tlv_word20.crc32  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m20 "\int_tlv_word0.tlv_bip2  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m21 "\int_tlv_word0.resv0  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m22 "\int_tlv_word0.kdf_dek_iter  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m23 "\int_tlv_word0.keyless_algos  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m24 "\int_tlv_word0.needs_dek  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m25 "\int_tlv_word0.needs_dak  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m26 "\int_tlv_word0.key_type  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m27 "\int_tlv_word0.tlv_frame_num  (1,0) 1 10 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m28 "\int_tlv_word0.tlv_eng_id  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m29 "\int_tlv_word0.tlv_seq_num  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m30 "\int_tlv_word0.tlv_len  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m31 "\int_tlv_word0.tlv_type  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m32 "\int_tlv_word42.corrupt_crc32  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m33 "\int_tlv_word42.unused  (1,0) 1 46 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m34 "\int_tlv_word42.error_code  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "34"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r1 "key_tlv_ob_tlv 10 \key_tlv_ob_tlv.insert  \key_tlv_ob_tlv.ordern  \key_tlv_ob_tlv.typen  \key_tlv_ob_tlv.sot  \key_tlv_ob_tlv.eot  \key_tlv_ob_tlv.tlast  \key_tlv_ob_tlv.tid  \key_tlv_ob_tlv.tstrb  \key_tlv_ob_tlv.tuser  \key_tlv_ob_tlv.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r2 "gcm_status_data_out 1 \gcm_status_data_out.tag_mismatch "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r3 "key_tlv_word0 8 \key_tlv_word0.tlv_bip2  \key_tlv_word0.resv0  \key_tlv_word0.tlv_frame_num  \key_tlv_word0.resv1  \key_tlv_word0.tlv_eng_id  \key_tlv_word0.tlv_seq_num  \key_tlv_word0.tlv_len  \key_tlv_word0.tlv_type "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r4 "key_tlv_word19 2 \key_tlv_word19.rsvd  \key_tlv_word19.kme_errors "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r5 "key_tlv_word20 2 \key_tlv_word20.rsvd  \key_tlv_word20.crc32 "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r6 "int_tlv_word0 12 \int_tlv_word0.tlv_bip2  \int_tlv_word0.resv0  \int_tlv_word0.kdf_dek_iter  \int_tlv_word0.keyless_algos  \int_tlv_word0.needs_dek  \int_tlv_word0.needs_dak  \int_tlv_word0.key_type  \int_tlv_word0.tlv_frame_num  \int_tlv_word0.tlv_eng_id  \int_tlv_word0.tlv_seq_num  \int_tlv_word0.tlv_len  \int_tlv_word0.tlv_type "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r7 "int_tlv_word42 3 \int_tlv_word42.corrupt_crc32  \int_tlv_word42.unused  \int_tlv_word42.error_code "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_NUM "7"
endmodule
