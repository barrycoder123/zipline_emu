
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
(* celldefine = 1 *) 
module nx_fifo_xcm28 ( empty, full, underflow, overflow, used_slots, free_slots, 
	rdata, clk, rst_n, wen, ren, clear, wdata);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output empty;
output full;
output underflow;
output overflow;
output [2:0] used_slots;
output [2:0] free_slots;
output [255:0] rdata;
input clk;
input rst_n;
input wen;
input ren;
input clear;
input [255:0] wdata;
wire _zy_simnet_underflow_0_w$;
wire _zy_simnet_overflow_1_w$;
wire \depth_n._zy_simnet_overflow_3_w$ ;
wire \depth_n._zy_simnet_underflow_2_w$ ;
wire [1:0] \depth_n.wptr ;
wire [1:0] \depth_n.rptr ;
supply0 n525;
ixc_assign _zz_strnp_3 ( _zy_simnet_overflow_1_w$, overflow);
ixc_assign _zz_strnp_2 ( _zy_simnet_underflow_0_w$, underflow);
Q_FDP0 U2 ( .CK(clk), .D(wdata[255]), .Q(n524), .QN( ));
Q_FDP0 U3 ( .CK(clk), .D(wdata[254]), .Q(n523), .QN( ));
Q_FDP0 U4 ( .CK(clk), .D(wdata[253]), .Q(n522), .QN( ));
Q_FDP0 U5 ( .CK(clk), .D(wdata[252]), .Q(n521), .QN( ));
Q_FDP0 U6 ( .CK(clk), .D(wdata[251]), .Q(n520), .QN( ));
Q_FDP0 U7 ( .CK(clk), .D(wdata[250]), .Q(n519), .QN( ));
Q_FDP0 U8 ( .CK(clk), .D(wdata[249]), .Q(n518), .QN( ));
Q_FDP0 U9 ( .CK(clk), .D(wdata[248]), .Q(n517), .QN( ));
Q_FDP0 U10 ( .CK(clk), .D(wdata[247]), .Q(n516), .QN( ));
Q_FDP0 U11 ( .CK(clk), .D(wdata[246]), .Q(n515), .QN( ));
Q_FDP0 U12 ( .CK(clk), .D(wdata[245]), .Q(n514), .QN( ));
Q_FDP0 U13 ( .CK(clk), .D(wdata[244]), .Q(n513), .QN( ));
Q_FDP0 U14 ( .CK(clk), .D(wdata[243]), .Q(n512), .QN( ));
Q_FDP0 U15 ( .CK(clk), .D(wdata[242]), .Q(n511), .QN( ));
Q_FDP0 U16 ( .CK(clk), .D(wdata[241]), .Q(n510), .QN( ));
Q_FDP0 U17 ( .CK(clk), .D(wdata[240]), .Q(n509), .QN( ));
Q_FDP0 U18 ( .CK(clk), .D(wdata[239]), .Q(n508), .QN( ));
Q_FDP0 U19 ( .CK(clk), .D(wdata[238]), .Q(n507), .QN( ));
Q_FDP0 U20 ( .CK(clk), .D(wdata[237]), .Q(n506), .QN( ));
Q_FDP0 U21 ( .CK(clk), .D(wdata[236]), .Q(n505), .QN( ));
Q_FDP0 U22 ( .CK(clk), .D(wdata[235]), .Q(n504), .QN( ));
Q_FDP0 U23 ( .CK(clk), .D(wdata[234]), .Q(n503), .QN( ));
Q_FDP0 U24 ( .CK(clk), .D(wdata[233]), .Q(n502), .QN( ));
Q_FDP0 U25 ( .CK(clk), .D(wdata[232]), .Q(n501), .QN( ));
Q_FDP0 U26 ( .CK(clk), .D(wdata[231]), .Q(n500), .QN( ));
Q_FDP0 U27 ( .CK(clk), .D(wdata[230]), .Q(n499), .QN( ));
Q_FDP0 U28 ( .CK(clk), .D(wdata[229]), .Q(n498), .QN( ));
Q_FDP0 U29 ( .CK(clk), .D(wdata[228]), .Q(n497), .QN( ));
Q_FDP0 U30 ( .CK(clk), .D(wdata[227]), .Q(n496), .QN( ));
Q_FDP0 U31 ( .CK(clk), .D(wdata[226]), .Q(n495), .QN( ));
Q_FDP0 U32 ( .CK(clk), .D(wdata[225]), .Q(n494), .QN( ));
Q_FDP0 U33 ( .CK(clk), .D(wdata[224]), .Q(n493), .QN( ));
Q_FDP0 U34 ( .CK(clk), .D(wdata[223]), .Q(n492), .QN( ));
Q_FDP0 U35 ( .CK(clk), .D(wdata[222]), .Q(n491), .QN( ));
Q_FDP0 U36 ( .CK(clk), .D(wdata[221]), .Q(n490), .QN( ));
Q_FDP0 U37 ( .CK(clk), .D(wdata[220]), .Q(n489), .QN( ));
Q_FDP0 U38 ( .CK(clk), .D(wdata[219]), .Q(n488), .QN( ));
Q_FDP0 U39 ( .CK(clk), .D(wdata[218]), .Q(n487), .QN( ));
Q_FDP0 U40 ( .CK(clk), .D(wdata[217]), .Q(n486), .QN( ));
Q_FDP0 U41 ( .CK(clk), .D(wdata[216]), .Q(n485), .QN( ));
Q_FDP0 U42 ( .CK(clk), .D(wdata[215]), .Q(n484), .QN( ));
Q_FDP0 U43 ( .CK(clk), .D(wdata[214]), .Q(n483), .QN( ));
Q_FDP0 U44 ( .CK(clk), .D(wdata[213]), .Q(n482), .QN( ));
Q_FDP0 U45 ( .CK(clk), .D(wdata[212]), .Q(n481), .QN( ));
Q_FDP0 U46 ( .CK(clk), .D(wdata[211]), .Q(n480), .QN( ));
Q_FDP0 U47 ( .CK(clk), .D(wdata[210]), .Q(n479), .QN( ));
Q_FDP0 U48 ( .CK(clk), .D(wdata[209]), .Q(n478), .QN( ));
Q_FDP0 U49 ( .CK(clk), .D(wdata[208]), .Q(n477), .QN( ));
Q_FDP0 U50 ( .CK(clk), .D(wdata[207]), .Q(n476), .QN( ));
Q_FDP0 U51 ( .CK(clk), .D(wdata[206]), .Q(n475), .QN( ));
Q_FDP0 U52 ( .CK(clk), .D(wdata[205]), .Q(n474), .QN( ));
Q_FDP0 U53 ( .CK(clk), .D(wdata[204]), .Q(n473), .QN( ));
Q_FDP0 U54 ( .CK(clk), .D(wdata[203]), .Q(n472), .QN( ));
Q_FDP0 U55 ( .CK(clk), .D(wdata[202]), .Q(n471), .QN( ));
Q_FDP0 U56 ( .CK(clk), .D(wdata[201]), .Q(n470), .QN( ));
Q_FDP0 U57 ( .CK(clk), .D(wdata[200]), .Q(n469), .QN( ));
Q_FDP0 U58 ( .CK(clk), .D(wdata[199]), .Q(n468), .QN( ));
Q_FDP0 U59 ( .CK(clk), .D(wdata[198]), .Q(n467), .QN( ));
Q_FDP0 U60 ( .CK(clk), .D(wdata[197]), .Q(n466), .QN( ));
Q_FDP0 U61 ( .CK(clk), .D(wdata[196]), .Q(n465), .QN( ));
Q_FDP0 U62 ( .CK(clk), .D(wdata[195]), .Q(n464), .QN( ));
Q_FDP0 U63 ( .CK(clk), .D(wdata[194]), .Q(n463), .QN( ));
Q_FDP0 U64 ( .CK(clk), .D(wdata[193]), .Q(n462), .QN( ));
Q_FDP0 U65 ( .CK(clk), .D(wdata[192]), .Q(n461), .QN( ));
Q_FDP0 U66 ( .CK(clk), .D(wdata[191]), .Q(n460), .QN( ));
Q_FDP0 U67 ( .CK(clk), .D(wdata[190]), .Q(n459), .QN( ));
Q_FDP0 U68 ( .CK(clk), .D(wdata[189]), .Q(n458), .QN( ));
Q_FDP0 U69 ( .CK(clk), .D(wdata[188]), .Q(n457), .QN( ));
Q_FDP0 U70 ( .CK(clk), .D(wdata[187]), .Q(n456), .QN( ));
Q_FDP0 U71 ( .CK(clk), .D(wdata[186]), .Q(n455), .QN( ));
Q_FDP0 U72 ( .CK(clk), .D(wdata[185]), .Q(n454), .QN( ));
Q_FDP0 U73 ( .CK(clk), .D(wdata[184]), .Q(n453), .QN( ));
Q_FDP0 U74 ( .CK(clk), .D(wdata[183]), .Q(n452), .QN( ));
Q_FDP0 U75 ( .CK(clk), .D(wdata[182]), .Q(n451), .QN( ));
Q_FDP0 U76 ( .CK(clk), .D(wdata[181]), .Q(n450), .QN( ));
Q_FDP0 U77 ( .CK(clk), .D(wdata[180]), .Q(n449), .QN( ));
Q_FDP0 U78 ( .CK(clk), .D(wdata[179]), .Q(n448), .QN( ));
Q_FDP0 U79 ( .CK(clk), .D(wdata[178]), .Q(n447), .QN( ));
Q_FDP0 U80 ( .CK(clk), .D(wdata[177]), .Q(n446), .QN( ));
Q_FDP0 U81 ( .CK(clk), .D(wdata[176]), .Q(n445), .QN( ));
Q_FDP0 U82 ( .CK(clk), .D(wdata[175]), .Q(n444), .QN( ));
Q_FDP0 U83 ( .CK(clk), .D(wdata[174]), .Q(n443), .QN( ));
Q_FDP0 U84 ( .CK(clk), .D(wdata[173]), .Q(n442), .QN( ));
Q_FDP0 U85 ( .CK(clk), .D(wdata[172]), .Q(n441), .QN( ));
Q_FDP0 U86 ( .CK(clk), .D(wdata[171]), .Q(n440), .QN( ));
Q_FDP0 U87 ( .CK(clk), .D(wdata[170]), .Q(n439), .QN( ));
Q_FDP0 U88 ( .CK(clk), .D(wdata[169]), .Q(n438), .QN( ));
Q_FDP0 U89 ( .CK(clk), .D(wdata[168]), .Q(n437), .QN( ));
Q_FDP0 U90 ( .CK(clk), .D(wdata[167]), .Q(n436), .QN( ));
Q_FDP0 U91 ( .CK(clk), .D(wdata[166]), .Q(n435), .QN( ));
Q_FDP0 U92 ( .CK(clk), .D(wdata[165]), .Q(n434), .QN( ));
Q_FDP0 U93 ( .CK(clk), .D(wdata[164]), .Q(n433), .QN( ));
Q_FDP0 U94 ( .CK(clk), .D(wdata[163]), .Q(n432), .QN( ));
Q_FDP0 U95 ( .CK(clk), .D(wdata[162]), .Q(n431), .QN( ));
Q_FDP0 U96 ( .CK(clk), .D(wdata[161]), .Q(n430), .QN( ));
Q_FDP0 U97 ( .CK(clk), .D(wdata[160]), .Q(n429), .QN( ));
Q_FDP0 U98 ( .CK(clk), .D(wdata[159]), .Q(n428), .QN( ));
Q_FDP0 U99 ( .CK(clk), .D(wdata[158]), .Q(n427), .QN( ));
Q_FDP0 U100 ( .CK(clk), .D(wdata[157]), .Q(n426), .QN( ));
Q_FDP0 U101 ( .CK(clk), .D(wdata[156]), .Q(n425), .QN( ));
Q_FDP0 U102 ( .CK(clk), .D(wdata[155]), .Q(n424), .QN( ));
Q_FDP0 U103 ( .CK(clk), .D(wdata[154]), .Q(n423), .QN( ));
Q_FDP0 U104 ( .CK(clk), .D(wdata[153]), .Q(n422), .QN( ));
Q_FDP0 U105 ( .CK(clk), .D(wdata[152]), .Q(n421), .QN( ));
Q_FDP0 U106 ( .CK(clk), .D(wdata[151]), .Q(n420), .QN( ));
Q_FDP0 U107 ( .CK(clk), .D(wdata[150]), .Q(n419), .QN( ));
Q_FDP0 U108 ( .CK(clk), .D(wdata[149]), .Q(n418), .QN( ));
Q_FDP0 U109 ( .CK(clk), .D(wdata[148]), .Q(n417), .QN( ));
Q_FDP0 U110 ( .CK(clk), .D(wdata[147]), .Q(n416), .QN( ));
Q_FDP0 U111 ( .CK(clk), .D(wdata[146]), .Q(n415), .QN( ));
Q_FDP0 U112 ( .CK(clk), .D(wdata[145]), .Q(n414), .QN( ));
Q_FDP0 U113 ( .CK(clk), .D(wdata[144]), .Q(n413), .QN( ));
Q_FDP0 U114 ( .CK(clk), .D(wdata[143]), .Q(n412), .QN( ));
Q_FDP0 U115 ( .CK(clk), .D(wdata[142]), .Q(n411), .QN( ));
Q_FDP0 U116 ( .CK(clk), .D(wdata[141]), .Q(n410), .QN( ));
Q_FDP0 U117 ( .CK(clk), .D(wdata[140]), .Q(n409), .QN( ));
Q_FDP0 U118 ( .CK(clk), .D(wdata[139]), .Q(n408), .QN( ));
Q_FDP0 U119 ( .CK(clk), .D(wdata[138]), .Q(n407), .QN( ));
Q_FDP0 U120 ( .CK(clk), .D(wdata[137]), .Q(n406), .QN( ));
Q_FDP0 U121 ( .CK(clk), .D(wdata[136]), .Q(n405), .QN( ));
Q_FDP0 U122 ( .CK(clk), .D(wdata[135]), .Q(n404), .QN( ));
Q_FDP0 U123 ( .CK(clk), .D(wdata[134]), .Q(n403), .QN( ));
Q_FDP0 U124 ( .CK(clk), .D(wdata[133]), .Q(n402), .QN( ));
Q_FDP0 U125 ( .CK(clk), .D(wdata[132]), .Q(n401), .QN( ));
Q_FDP0 U126 ( .CK(clk), .D(wdata[131]), .Q(n400), .QN( ));
Q_FDP0 U127 ( .CK(clk), .D(wdata[130]), .Q(n399), .QN( ));
Q_FDP0 U128 ( .CK(clk), .D(wdata[129]), .Q(n398), .QN( ));
Q_FDP0 U129 ( .CK(clk), .D(wdata[128]), .Q(n397), .QN( ));
Q_FDP0 U130 ( .CK(clk), .D(wdata[127]), .Q(n396), .QN( ));
Q_FDP0 U131 ( .CK(clk), .D(wdata[126]), .Q(n395), .QN( ));
Q_FDP0 U132 ( .CK(clk), .D(wdata[125]), .Q(n394), .QN( ));
Q_FDP0 U133 ( .CK(clk), .D(wdata[124]), .Q(n393), .QN( ));
Q_FDP0 U134 ( .CK(clk), .D(wdata[123]), .Q(n392), .QN( ));
Q_FDP0 U135 ( .CK(clk), .D(wdata[122]), .Q(n391), .QN( ));
Q_FDP0 U136 ( .CK(clk), .D(wdata[121]), .Q(n390), .QN( ));
Q_FDP0 U137 ( .CK(clk), .D(wdata[120]), .Q(n389), .QN( ));
Q_FDP0 U138 ( .CK(clk), .D(wdata[119]), .Q(n388), .QN( ));
Q_FDP0 U139 ( .CK(clk), .D(wdata[118]), .Q(n387), .QN( ));
Q_FDP0 U140 ( .CK(clk), .D(wdata[117]), .Q(n386), .QN( ));
Q_FDP0 U141 ( .CK(clk), .D(wdata[116]), .Q(n385), .QN( ));
Q_FDP0 U142 ( .CK(clk), .D(wdata[115]), .Q(n384), .QN( ));
Q_FDP0 U143 ( .CK(clk), .D(wdata[114]), .Q(n383), .QN( ));
Q_FDP0 U144 ( .CK(clk), .D(wdata[113]), .Q(n382), .QN( ));
Q_FDP0 U145 ( .CK(clk), .D(wdata[112]), .Q(n381), .QN( ));
Q_FDP0 U146 ( .CK(clk), .D(wdata[111]), .Q(n380), .QN( ));
Q_FDP0 U147 ( .CK(clk), .D(wdata[110]), .Q(n379), .QN( ));
Q_FDP0 U148 ( .CK(clk), .D(wdata[109]), .Q(n378), .QN( ));
Q_FDP0 U149 ( .CK(clk), .D(wdata[108]), .Q(n377), .QN( ));
Q_FDP0 U150 ( .CK(clk), .D(wdata[107]), .Q(n376), .QN( ));
Q_FDP0 U151 ( .CK(clk), .D(wdata[106]), .Q(n375), .QN( ));
Q_FDP0 U152 ( .CK(clk), .D(wdata[105]), .Q(n374), .QN( ));
Q_FDP0 U153 ( .CK(clk), .D(wdata[104]), .Q(n373), .QN( ));
Q_FDP0 U154 ( .CK(clk), .D(wdata[103]), .Q(n372), .QN( ));
Q_FDP0 U155 ( .CK(clk), .D(wdata[102]), .Q(n371), .QN( ));
Q_FDP0 U156 ( .CK(clk), .D(wdata[101]), .Q(n370), .QN( ));
Q_FDP0 U157 ( .CK(clk), .D(wdata[100]), .Q(n369), .QN( ));
Q_FDP0 U158 ( .CK(clk), .D(wdata[99]), .Q(n368), .QN( ));
Q_FDP0 U159 ( .CK(clk), .D(wdata[98]), .Q(n367), .QN( ));
Q_FDP0 U160 ( .CK(clk), .D(wdata[97]), .Q(n366), .QN( ));
Q_FDP0 U161 ( .CK(clk), .D(wdata[96]), .Q(n365), .QN( ));
Q_FDP0 U162 ( .CK(clk), .D(wdata[95]), .Q(n364), .QN( ));
Q_FDP0 U163 ( .CK(clk), .D(wdata[94]), .Q(n363), .QN( ));
Q_FDP0 U164 ( .CK(clk), .D(wdata[93]), .Q(n362), .QN( ));
Q_FDP0 U165 ( .CK(clk), .D(wdata[92]), .Q(n361), .QN( ));
Q_FDP0 U166 ( .CK(clk), .D(wdata[91]), .Q(n360), .QN( ));
Q_FDP0 U167 ( .CK(clk), .D(wdata[90]), .Q(n359), .QN( ));
Q_FDP0 U168 ( .CK(clk), .D(wdata[89]), .Q(n358), .QN( ));
Q_FDP0 U169 ( .CK(clk), .D(wdata[88]), .Q(n357), .QN( ));
Q_FDP0 U170 ( .CK(clk), .D(wdata[87]), .Q(n356), .QN( ));
Q_FDP0 U171 ( .CK(clk), .D(wdata[86]), .Q(n355), .QN( ));
Q_FDP0 U172 ( .CK(clk), .D(wdata[85]), .Q(n354), .QN( ));
Q_FDP0 U173 ( .CK(clk), .D(wdata[84]), .Q(n353), .QN( ));
Q_FDP0 U174 ( .CK(clk), .D(wdata[83]), .Q(n352), .QN( ));
Q_FDP0 U175 ( .CK(clk), .D(wdata[82]), .Q(n351), .QN( ));
Q_FDP0 U176 ( .CK(clk), .D(wdata[81]), .Q(n350), .QN( ));
Q_FDP0 U177 ( .CK(clk), .D(wdata[80]), .Q(n349), .QN( ));
Q_FDP0 U178 ( .CK(clk), .D(wdata[79]), .Q(n348), .QN( ));
Q_FDP0 U179 ( .CK(clk), .D(wdata[78]), .Q(n347), .QN( ));
Q_FDP0 U180 ( .CK(clk), .D(wdata[77]), .Q(n346), .QN( ));
Q_FDP0 U181 ( .CK(clk), .D(wdata[76]), .Q(n345), .QN( ));
Q_FDP0 U182 ( .CK(clk), .D(wdata[75]), .Q(n344), .QN( ));
Q_FDP0 U183 ( .CK(clk), .D(wdata[74]), .Q(n343), .QN( ));
Q_FDP0 U184 ( .CK(clk), .D(wdata[73]), .Q(n342), .QN( ));
Q_FDP0 U185 ( .CK(clk), .D(wdata[72]), .Q(n341), .QN( ));
Q_FDP0 U186 ( .CK(clk), .D(wdata[71]), .Q(n340), .QN( ));
Q_FDP0 U187 ( .CK(clk), .D(wdata[70]), .Q(n339), .QN( ));
Q_FDP0 U188 ( .CK(clk), .D(wdata[69]), .Q(n338), .QN( ));
Q_FDP0 U189 ( .CK(clk), .D(wdata[68]), .Q(n337), .QN( ));
Q_FDP0 U190 ( .CK(clk), .D(wdata[67]), .Q(n336), .QN( ));
Q_FDP0 U191 ( .CK(clk), .D(wdata[66]), .Q(n335), .QN( ));
Q_FDP0 U192 ( .CK(clk), .D(wdata[65]), .Q(n334), .QN( ));
Q_FDP0 U193 ( .CK(clk), .D(wdata[64]), .Q(n333), .QN( ));
Q_FDP0 U194 ( .CK(clk), .D(wdata[63]), .Q(n332), .QN( ));
Q_FDP0 U195 ( .CK(clk), .D(wdata[62]), .Q(n331), .QN( ));
Q_FDP0 U196 ( .CK(clk), .D(wdata[61]), .Q(n330), .QN( ));
Q_FDP0 U197 ( .CK(clk), .D(wdata[60]), .Q(n329), .QN( ));
Q_FDP0 U198 ( .CK(clk), .D(wdata[59]), .Q(n328), .QN( ));
Q_FDP0 U199 ( .CK(clk), .D(wdata[58]), .Q(n327), .QN( ));
Q_FDP0 U200 ( .CK(clk), .D(wdata[57]), .Q(n326), .QN( ));
Q_FDP0 U201 ( .CK(clk), .D(wdata[56]), .Q(n325), .QN( ));
Q_FDP0 U202 ( .CK(clk), .D(wdata[55]), .Q(n324), .QN( ));
Q_FDP0 U203 ( .CK(clk), .D(wdata[54]), .Q(n323), .QN( ));
Q_FDP0 U204 ( .CK(clk), .D(wdata[53]), .Q(n322), .QN( ));
Q_FDP0 U205 ( .CK(clk), .D(wdata[52]), .Q(n321), .QN( ));
Q_FDP0 U206 ( .CK(clk), .D(wdata[51]), .Q(n320), .QN( ));
Q_FDP0 U207 ( .CK(clk), .D(wdata[50]), .Q(n319), .QN( ));
Q_FDP0 U208 ( .CK(clk), .D(wdata[49]), .Q(n318), .QN( ));
Q_FDP0 U209 ( .CK(clk), .D(wdata[48]), .Q(n317), .QN( ));
Q_FDP0 U210 ( .CK(clk), .D(wdata[47]), .Q(n316), .QN( ));
Q_FDP0 U211 ( .CK(clk), .D(wdata[46]), .Q(n315), .QN( ));
Q_FDP0 U212 ( .CK(clk), .D(wdata[45]), .Q(n314), .QN( ));
Q_FDP0 U213 ( .CK(clk), .D(wdata[44]), .Q(n313), .QN( ));
Q_FDP0 U214 ( .CK(clk), .D(wdata[43]), .Q(n312), .QN( ));
Q_FDP0 U215 ( .CK(clk), .D(wdata[42]), .Q(n311), .QN( ));
Q_FDP0 U216 ( .CK(clk), .D(wdata[41]), .Q(n310), .QN( ));
Q_FDP0 U217 ( .CK(clk), .D(wdata[40]), .Q(n309), .QN( ));
Q_FDP0 U218 ( .CK(clk), .D(wdata[39]), .Q(n308), .QN( ));
Q_FDP0 U219 ( .CK(clk), .D(wdata[38]), .Q(n307), .QN( ));
Q_FDP0 U220 ( .CK(clk), .D(wdata[37]), .Q(n306), .QN( ));
Q_FDP0 U221 ( .CK(clk), .D(wdata[36]), .Q(n305), .QN( ));
Q_FDP0 U222 ( .CK(clk), .D(wdata[35]), .Q(n304), .QN( ));
Q_FDP0 U223 ( .CK(clk), .D(wdata[34]), .Q(n303), .QN( ));
Q_FDP0 U224 ( .CK(clk), .D(wdata[33]), .Q(n302), .QN( ));
Q_FDP0 U225 ( .CK(clk), .D(wdata[32]), .Q(n301), .QN( ));
Q_FDP0 U226 ( .CK(clk), .D(wdata[31]), .Q(n300), .QN( ));
Q_FDP0 U227 ( .CK(clk), .D(wdata[30]), .Q(n299), .QN( ));
Q_FDP0 U228 ( .CK(clk), .D(wdata[29]), .Q(n298), .QN( ));
Q_FDP0 U229 ( .CK(clk), .D(wdata[28]), .Q(n297), .QN( ));
Q_FDP0 U230 ( .CK(clk), .D(wdata[27]), .Q(n296), .QN( ));
Q_FDP0 U231 ( .CK(clk), .D(wdata[26]), .Q(n295), .QN( ));
Q_FDP0 U232 ( .CK(clk), .D(wdata[25]), .Q(n294), .QN( ));
Q_FDP0 U233 ( .CK(clk), .D(wdata[24]), .Q(n293), .QN( ));
Q_FDP0 U234 ( .CK(clk), .D(wdata[23]), .Q(n292), .QN( ));
Q_FDP0 U235 ( .CK(clk), .D(wdata[22]), .Q(n291), .QN( ));
Q_FDP0 U236 ( .CK(clk), .D(wdata[21]), .Q(n290), .QN( ));
Q_FDP0 U237 ( .CK(clk), .D(wdata[20]), .Q(n289), .QN( ));
Q_FDP0 U238 ( .CK(clk), .D(wdata[19]), .Q(n288), .QN( ));
Q_FDP0 U239 ( .CK(clk), .D(wdata[18]), .Q(n287), .QN( ));
Q_FDP0 U240 ( .CK(clk), .D(wdata[17]), .Q(n286), .QN( ));
Q_FDP0 U241 ( .CK(clk), .D(wdata[16]), .Q(n285), .QN( ));
Q_FDP0 U242 ( .CK(clk), .D(wdata[15]), .Q(n284), .QN( ));
Q_FDP0 U243 ( .CK(clk), .D(wdata[14]), .Q(n283), .QN( ));
Q_FDP0 U244 ( .CK(clk), .D(wdata[13]), .Q(n282), .QN( ));
Q_FDP0 U245 ( .CK(clk), .D(wdata[12]), .Q(n281), .QN( ));
Q_FDP0 U246 ( .CK(clk), .D(wdata[11]), .Q(n280), .QN( ));
Q_FDP0 U247 ( .CK(clk), .D(wdata[10]), .Q(n279), .QN( ));
Q_FDP0 U248 ( .CK(clk), .D(wdata[9]), .Q(n278), .QN( ));
Q_FDP0 U249 ( .CK(clk), .D(wdata[8]), .Q(n277), .QN( ));
Q_FDP0 U250 ( .CK(clk), .D(wdata[7]), .Q(n276), .QN( ));
Q_FDP0 U251 ( .CK(clk), .D(wdata[6]), .Q(n275), .QN( ));
Q_FDP0 U252 ( .CK(clk), .D(wdata[5]), .Q(n274), .QN( ));
Q_FDP0 U253 ( .CK(clk), .D(wdata[4]), .Q(n273), .QN( ));
Q_FDP0 U254 ( .CK(clk), .D(wdata[3]), .Q(n272), .QN( ));
Q_FDP0 U255 ( .CK(clk), .D(wdata[2]), .Q(n271), .QN( ));
Q_FDP0 U256 ( .CK(clk), .D(wdata[1]), .Q(n270), .QN( ));
Q_FDP0 U257 ( .CK(clk), .D(wdata[0]), .Q(n269), .QN( ));
Q_FDP0 U258 ( .CK(clk), .D(\depth_n.wptr [1]), .Q(n268), .QN( ));
Q_FDP0 U259 ( .CK(clk), .D(\depth_n.wptr [0]), .Q(n267), .QN( ));
Q_AN02 U260 ( .A0(n262), .A1(n265), .Z(n266));
Q_XOR2 U261 ( .A0(n261), .A1(n264), .Z(n265));
// pragma CVAINTPROP NET n261 _2_state_ 1
// pragma CVAINTPROP INSTANCE U261 NOBREAKS 1
Q_FDP0B U262 ( .D(n261), .QTFCLK( ), .Q(n264));
Q_FDP0 U263 ( .CK(clk), .D(n3), .Q(n262), .QN( ));
Q_FDP0 U264 ( .CK(clk), .D(n263), .Q(n261), .QN(n263));
Q_INV U265 ( .A(empty), .Z(n260));
Q_AN02 U266 ( .A0(n260), .A1(n4), .Z(rdata[255]));
Q_AN02 U267 ( .A0(n260), .A1(n5), .Z(rdata[254]));
Q_AN02 U268 ( .A0(n260), .A1(n6), .Z(rdata[253]));
Q_AN02 U269 ( .A0(n260), .A1(n7), .Z(rdata[252]));
Q_AN02 U270 ( .A0(n260), .A1(n8), .Z(rdata[251]));
Q_AN02 U271 ( .A0(n260), .A1(n9), .Z(rdata[250]));
Q_AN02 U272 ( .A0(n260), .A1(n10), .Z(rdata[249]));
Q_AN02 U273 ( .A0(n260), .A1(n11), .Z(rdata[248]));
Q_AN02 U274 ( .A0(n260), .A1(n12), .Z(rdata[247]));
Q_AN02 U275 ( .A0(n260), .A1(n13), .Z(rdata[246]));
Q_AN02 U276 ( .A0(n260), .A1(n14), .Z(rdata[245]));
Q_AN02 U277 ( .A0(n260), .A1(n15), .Z(rdata[244]));
Q_AN02 U278 ( .A0(n260), .A1(n16), .Z(rdata[243]));
Q_AN02 U279 ( .A0(n260), .A1(n17), .Z(rdata[242]));
Q_AN02 U280 ( .A0(n260), .A1(n18), .Z(rdata[241]));
Q_AN02 U281 ( .A0(n260), .A1(n19), .Z(rdata[240]));
Q_AN02 U282 ( .A0(n260), .A1(n20), .Z(rdata[239]));
Q_AN02 U283 ( .A0(n260), .A1(n21), .Z(rdata[238]));
Q_AN02 U284 ( .A0(n260), .A1(n22), .Z(rdata[237]));
Q_AN02 U285 ( .A0(n260), .A1(n23), .Z(rdata[236]));
Q_AN02 U286 ( .A0(n260), .A1(n24), .Z(rdata[235]));
Q_AN02 U287 ( .A0(n260), .A1(n25), .Z(rdata[234]));
Q_AN02 U288 ( .A0(n260), .A1(n26), .Z(rdata[233]));
Q_AN02 U289 ( .A0(n260), .A1(n27), .Z(rdata[232]));
Q_AN02 U290 ( .A0(n260), .A1(n28), .Z(rdata[231]));
Q_AN02 U291 ( .A0(n260), .A1(n29), .Z(rdata[230]));
Q_AN02 U292 ( .A0(n260), .A1(n30), .Z(rdata[229]));
Q_AN02 U293 ( .A0(n260), .A1(n31), .Z(rdata[228]));
Q_AN02 U294 ( .A0(n260), .A1(n32), .Z(rdata[227]));
Q_AN02 U295 ( .A0(n260), .A1(n33), .Z(rdata[226]));
Q_AN02 U296 ( .A0(n260), .A1(n34), .Z(rdata[225]));
Q_AN02 U297 ( .A0(n260), .A1(n35), .Z(rdata[224]));
Q_AN02 U298 ( .A0(n260), .A1(n36), .Z(rdata[223]));
Q_AN02 U299 ( .A0(n260), .A1(n37), .Z(rdata[222]));
Q_AN02 U300 ( .A0(n260), .A1(n38), .Z(rdata[221]));
Q_AN02 U301 ( .A0(n260), .A1(n39), .Z(rdata[220]));
Q_AN02 U302 ( .A0(n260), .A1(n40), .Z(rdata[219]));
Q_AN02 U303 ( .A0(n260), .A1(n41), .Z(rdata[218]));
Q_AN02 U304 ( .A0(n260), .A1(n42), .Z(rdata[217]));
Q_AN02 U305 ( .A0(n260), .A1(n43), .Z(rdata[216]));
Q_AN02 U306 ( .A0(n260), .A1(n44), .Z(rdata[215]));
Q_AN02 U307 ( .A0(n260), .A1(n45), .Z(rdata[214]));
Q_AN02 U308 ( .A0(n260), .A1(n46), .Z(rdata[213]));
Q_AN02 U309 ( .A0(n260), .A1(n47), .Z(rdata[212]));
Q_AN02 U310 ( .A0(n260), .A1(n48), .Z(rdata[211]));
Q_AN02 U311 ( .A0(n260), .A1(n49), .Z(rdata[210]));
Q_AN02 U312 ( .A0(n260), .A1(n50), .Z(rdata[209]));
Q_AN02 U313 ( .A0(n260), .A1(n51), .Z(rdata[208]));
Q_AN02 U314 ( .A0(n260), .A1(n52), .Z(rdata[207]));
Q_AN02 U315 ( .A0(n260), .A1(n53), .Z(rdata[206]));
Q_AN02 U316 ( .A0(n260), .A1(n54), .Z(rdata[205]));
Q_AN02 U317 ( .A0(n260), .A1(n55), .Z(rdata[204]));
Q_AN02 U318 ( .A0(n260), .A1(n56), .Z(rdata[203]));
Q_AN02 U319 ( .A0(n260), .A1(n57), .Z(rdata[202]));
Q_AN02 U320 ( .A0(n260), .A1(n58), .Z(rdata[201]));
Q_AN02 U321 ( .A0(n260), .A1(n59), .Z(rdata[200]));
Q_AN02 U322 ( .A0(n260), .A1(n60), .Z(rdata[199]));
Q_AN02 U323 ( .A0(n260), .A1(n61), .Z(rdata[198]));
Q_AN02 U324 ( .A0(n260), .A1(n62), .Z(rdata[197]));
Q_AN02 U325 ( .A0(n260), .A1(n63), .Z(rdata[196]));
Q_AN02 U326 ( .A0(n260), .A1(n64), .Z(rdata[195]));
Q_AN02 U327 ( .A0(n260), .A1(n65), .Z(rdata[194]));
Q_AN02 U328 ( .A0(n260), .A1(n66), .Z(rdata[193]));
Q_AN02 U329 ( .A0(n260), .A1(n67), .Z(rdata[192]));
Q_AN02 U330 ( .A0(n260), .A1(n68), .Z(rdata[191]));
Q_AN02 U331 ( .A0(n260), .A1(n69), .Z(rdata[190]));
Q_AN02 U332 ( .A0(n260), .A1(n70), .Z(rdata[189]));
Q_AN02 U333 ( .A0(n260), .A1(n71), .Z(rdata[188]));
Q_AN02 U334 ( .A0(n260), .A1(n72), .Z(rdata[187]));
Q_AN02 U335 ( .A0(n260), .A1(n73), .Z(rdata[186]));
Q_AN02 U336 ( .A0(n260), .A1(n74), .Z(rdata[185]));
Q_AN02 U337 ( .A0(n260), .A1(n75), .Z(rdata[184]));
Q_AN02 U338 ( .A0(n260), .A1(n76), .Z(rdata[183]));
Q_AN02 U339 ( .A0(n260), .A1(n77), .Z(rdata[182]));
Q_AN02 U340 ( .A0(n260), .A1(n78), .Z(rdata[181]));
Q_AN02 U341 ( .A0(n260), .A1(n79), .Z(rdata[180]));
Q_AN02 U342 ( .A0(n260), .A1(n80), .Z(rdata[179]));
Q_AN02 U343 ( .A0(n260), .A1(n81), .Z(rdata[178]));
Q_AN02 U344 ( .A0(n260), .A1(n82), .Z(rdata[177]));
Q_AN02 U345 ( .A0(n260), .A1(n83), .Z(rdata[176]));
Q_AN02 U346 ( .A0(n260), .A1(n84), .Z(rdata[175]));
Q_AN02 U347 ( .A0(n260), .A1(n85), .Z(rdata[174]));
Q_AN02 U348 ( .A0(n260), .A1(n86), .Z(rdata[173]));
Q_AN02 U349 ( .A0(n260), .A1(n87), .Z(rdata[172]));
Q_AN02 U350 ( .A0(n260), .A1(n88), .Z(rdata[171]));
Q_AN02 U351 ( .A0(n260), .A1(n89), .Z(rdata[170]));
Q_AN02 U352 ( .A0(n260), .A1(n90), .Z(rdata[169]));
Q_AN02 U353 ( .A0(n260), .A1(n91), .Z(rdata[168]));
Q_AN02 U354 ( .A0(n260), .A1(n92), .Z(rdata[167]));
Q_AN02 U355 ( .A0(n260), .A1(n93), .Z(rdata[166]));
Q_AN02 U356 ( .A0(n260), .A1(n94), .Z(rdata[165]));
Q_AN02 U357 ( .A0(n260), .A1(n95), .Z(rdata[164]));
Q_AN02 U358 ( .A0(n260), .A1(n96), .Z(rdata[163]));
Q_AN02 U359 ( .A0(n260), .A1(n97), .Z(rdata[162]));
Q_AN02 U360 ( .A0(n260), .A1(n98), .Z(rdata[161]));
Q_AN02 U361 ( .A0(n260), .A1(n99), .Z(rdata[160]));
Q_AN02 U362 ( .A0(n260), .A1(n100), .Z(rdata[159]));
Q_AN02 U363 ( .A0(n260), .A1(n101), .Z(rdata[158]));
Q_AN02 U364 ( .A0(n260), .A1(n102), .Z(rdata[157]));
Q_AN02 U365 ( .A0(n260), .A1(n103), .Z(rdata[156]));
Q_AN02 U366 ( .A0(n260), .A1(n104), .Z(rdata[155]));
Q_AN02 U367 ( .A0(n260), .A1(n105), .Z(rdata[154]));
Q_AN02 U368 ( .A0(n260), .A1(n106), .Z(rdata[153]));
Q_AN02 U369 ( .A0(n260), .A1(n107), .Z(rdata[152]));
Q_AN02 U370 ( .A0(n260), .A1(n108), .Z(rdata[151]));
Q_AN02 U371 ( .A0(n260), .A1(n109), .Z(rdata[150]));
Q_AN02 U372 ( .A0(n260), .A1(n110), .Z(rdata[149]));
Q_AN02 U373 ( .A0(n260), .A1(n111), .Z(rdata[148]));
Q_AN02 U374 ( .A0(n260), .A1(n112), .Z(rdata[147]));
Q_AN02 U375 ( .A0(n260), .A1(n113), .Z(rdata[146]));
Q_AN02 U376 ( .A0(n260), .A1(n114), .Z(rdata[145]));
Q_AN02 U377 ( .A0(n260), .A1(n115), .Z(rdata[144]));
Q_AN02 U378 ( .A0(n260), .A1(n116), .Z(rdata[143]));
Q_AN02 U379 ( .A0(n260), .A1(n117), .Z(rdata[142]));
Q_AN02 U380 ( .A0(n260), .A1(n118), .Z(rdata[141]));
Q_AN02 U381 ( .A0(n260), .A1(n119), .Z(rdata[140]));
Q_AN02 U382 ( .A0(n260), .A1(n120), .Z(rdata[139]));
Q_AN02 U383 ( .A0(n260), .A1(n121), .Z(rdata[138]));
Q_AN02 U384 ( .A0(n260), .A1(n122), .Z(rdata[137]));
Q_AN02 U385 ( .A0(n260), .A1(n123), .Z(rdata[136]));
Q_AN02 U386 ( .A0(n260), .A1(n124), .Z(rdata[135]));
Q_AN02 U387 ( .A0(n260), .A1(n125), .Z(rdata[134]));
Q_AN02 U388 ( .A0(n260), .A1(n126), .Z(rdata[133]));
Q_AN02 U389 ( .A0(n260), .A1(n127), .Z(rdata[132]));
Q_AN02 U390 ( .A0(n260), .A1(n128), .Z(rdata[131]));
Q_AN02 U391 ( .A0(n260), .A1(n129), .Z(rdata[130]));
Q_AN02 U392 ( .A0(n260), .A1(n130), .Z(rdata[129]));
Q_AN02 U393 ( .A0(n260), .A1(n131), .Z(rdata[128]));
Q_AN02 U394 ( .A0(n260), .A1(n132), .Z(rdata[127]));
Q_AN02 U395 ( .A0(n260), .A1(n133), .Z(rdata[126]));
Q_AN02 U396 ( .A0(n260), .A1(n134), .Z(rdata[125]));
Q_AN02 U397 ( .A0(n260), .A1(n135), .Z(rdata[124]));
Q_AN02 U398 ( .A0(n260), .A1(n136), .Z(rdata[123]));
Q_AN02 U399 ( .A0(n260), .A1(n137), .Z(rdata[122]));
Q_AN02 U400 ( .A0(n260), .A1(n138), .Z(rdata[121]));
Q_AN02 U401 ( .A0(n260), .A1(n139), .Z(rdata[120]));
Q_AN02 U402 ( .A0(n260), .A1(n140), .Z(rdata[119]));
Q_AN02 U403 ( .A0(n260), .A1(n141), .Z(rdata[118]));
Q_AN02 U404 ( .A0(n260), .A1(n142), .Z(rdata[117]));
Q_AN02 U405 ( .A0(n260), .A1(n143), .Z(rdata[116]));
Q_AN02 U406 ( .A0(n260), .A1(n144), .Z(rdata[115]));
Q_AN02 U407 ( .A0(n260), .A1(n145), .Z(rdata[114]));
Q_AN02 U408 ( .A0(n260), .A1(n146), .Z(rdata[113]));
Q_AN02 U409 ( .A0(n260), .A1(n147), .Z(rdata[112]));
Q_AN02 U410 ( .A0(n260), .A1(n148), .Z(rdata[111]));
Q_AN02 U411 ( .A0(n260), .A1(n149), .Z(rdata[110]));
Q_AN02 U412 ( .A0(n260), .A1(n150), .Z(rdata[109]));
Q_AN02 U413 ( .A0(n260), .A1(n151), .Z(rdata[108]));
Q_AN02 U414 ( .A0(n260), .A1(n152), .Z(rdata[107]));
Q_AN02 U415 ( .A0(n260), .A1(n153), .Z(rdata[106]));
Q_AN02 U416 ( .A0(n260), .A1(n154), .Z(rdata[105]));
Q_AN02 U417 ( .A0(n260), .A1(n155), .Z(rdata[104]));
Q_AN02 U418 ( .A0(n260), .A1(n156), .Z(rdata[103]));
Q_AN02 U419 ( .A0(n260), .A1(n157), .Z(rdata[102]));
Q_AN02 U420 ( .A0(n260), .A1(n158), .Z(rdata[101]));
Q_AN02 U421 ( .A0(n260), .A1(n159), .Z(rdata[100]));
Q_AN02 U422 ( .A0(n260), .A1(n160), .Z(rdata[99]));
Q_AN02 U423 ( .A0(n260), .A1(n161), .Z(rdata[98]));
Q_AN02 U424 ( .A0(n260), .A1(n162), .Z(rdata[97]));
Q_AN02 U425 ( .A0(n260), .A1(n163), .Z(rdata[96]));
Q_AN02 U426 ( .A0(n260), .A1(n164), .Z(rdata[95]));
Q_AN02 U427 ( .A0(n260), .A1(n165), .Z(rdata[94]));
Q_AN02 U428 ( .A0(n260), .A1(n166), .Z(rdata[93]));
Q_AN02 U429 ( .A0(n260), .A1(n167), .Z(rdata[92]));
Q_AN02 U430 ( .A0(n260), .A1(n168), .Z(rdata[91]));
Q_AN02 U431 ( .A0(n260), .A1(n169), .Z(rdata[90]));
Q_AN02 U432 ( .A0(n260), .A1(n170), .Z(rdata[89]));
Q_AN02 U433 ( .A0(n260), .A1(n171), .Z(rdata[88]));
Q_AN02 U434 ( .A0(n260), .A1(n172), .Z(rdata[87]));
Q_AN02 U435 ( .A0(n260), .A1(n173), .Z(rdata[86]));
Q_AN02 U436 ( .A0(n260), .A1(n174), .Z(rdata[85]));
Q_AN02 U437 ( .A0(n260), .A1(n175), .Z(rdata[84]));
Q_AN02 U438 ( .A0(n260), .A1(n176), .Z(rdata[83]));
Q_AN02 U439 ( .A0(n260), .A1(n177), .Z(rdata[82]));
Q_AN02 U440 ( .A0(n260), .A1(n178), .Z(rdata[81]));
Q_AN02 U441 ( .A0(n260), .A1(n179), .Z(rdata[80]));
Q_AN02 U442 ( .A0(n260), .A1(n180), .Z(rdata[79]));
Q_AN02 U443 ( .A0(n260), .A1(n181), .Z(rdata[78]));
Q_AN02 U444 ( .A0(n260), .A1(n182), .Z(rdata[77]));
Q_AN02 U445 ( .A0(n260), .A1(n183), .Z(rdata[76]));
Q_AN02 U446 ( .A0(n260), .A1(n184), .Z(rdata[75]));
Q_AN02 U447 ( .A0(n260), .A1(n185), .Z(rdata[74]));
Q_AN02 U448 ( .A0(n260), .A1(n186), .Z(rdata[73]));
Q_AN02 U449 ( .A0(n260), .A1(n187), .Z(rdata[72]));
Q_AN02 U450 ( .A0(n260), .A1(n188), .Z(rdata[71]));
Q_AN02 U451 ( .A0(n260), .A1(n189), .Z(rdata[70]));
Q_AN02 U452 ( .A0(n260), .A1(n190), .Z(rdata[69]));
Q_AN02 U453 ( .A0(n260), .A1(n191), .Z(rdata[68]));
Q_AN02 U454 ( .A0(n260), .A1(n192), .Z(rdata[67]));
Q_AN02 U455 ( .A0(n260), .A1(n193), .Z(rdata[66]));
Q_AN02 U456 ( .A0(n260), .A1(n194), .Z(rdata[65]));
Q_AN02 U457 ( .A0(n260), .A1(n195), .Z(rdata[64]));
Q_AN02 U458 ( .A0(n260), .A1(n196), .Z(rdata[63]));
Q_AN02 U459 ( .A0(n260), .A1(n197), .Z(rdata[62]));
Q_AN02 U460 ( .A0(n260), .A1(n198), .Z(rdata[61]));
Q_AN02 U461 ( .A0(n260), .A1(n199), .Z(rdata[60]));
Q_AN02 U462 ( .A0(n260), .A1(n200), .Z(rdata[59]));
Q_AN02 U463 ( .A0(n260), .A1(n201), .Z(rdata[58]));
Q_AN02 U464 ( .A0(n260), .A1(n202), .Z(rdata[57]));
Q_AN02 U465 ( .A0(n260), .A1(n203), .Z(rdata[56]));
Q_AN02 U466 ( .A0(n260), .A1(n204), .Z(rdata[55]));
Q_AN02 U467 ( .A0(n260), .A1(n205), .Z(rdata[54]));
Q_AN02 U468 ( .A0(n260), .A1(n206), .Z(rdata[53]));
Q_AN02 U469 ( .A0(n260), .A1(n207), .Z(rdata[52]));
Q_AN02 U470 ( .A0(n260), .A1(n208), .Z(rdata[51]));
Q_AN02 U471 ( .A0(n260), .A1(n209), .Z(rdata[50]));
Q_AN02 U472 ( .A0(n260), .A1(n210), .Z(rdata[49]));
Q_AN02 U473 ( .A0(n260), .A1(n211), .Z(rdata[48]));
Q_AN02 U474 ( .A0(n260), .A1(n212), .Z(rdata[47]));
Q_AN02 U475 ( .A0(n260), .A1(n213), .Z(rdata[46]));
Q_AN02 U476 ( .A0(n260), .A1(n214), .Z(rdata[45]));
Q_AN02 U477 ( .A0(n260), .A1(n215), .Z(rdata[44]));
Q_AN02 U478 ( .A0(n260), .A1(n216), .Z(rdata[43]));
Q_AN02 U479 ( .A0(n260), .A1(n217), .Z(rdata[42]));
Q_AN02 U480 ( .A0(n260), .A1(n218), .Z(rdata[41]));
Q_AN02 U481 ( .A0(n260), .A1(n219), .Z(rdata[40]));
Q_AN02 U482 ( .A0(n260), .A1(n220), .Z(rdata[39]));
Q_AN02 U483 ( .A0(n260), .A1(n221), .Z(rdata[38]));
Q_AN02 U484 ( .A0(n260), .A1(n222), .Z(rdata[37]));
Q_AN02 U485 ( .A0(n260), .A1(n223), .Z(rdata[36]));
Q_AN02 U486 ( .A0(n260), .A1(n224), .Z(rdata[35]));
Q_AN02 U487 ( .A0(n260), .A1(n225), .Z(rdata[34]));
Q_AN02 U488 ( .A0(n260), .A1(n226), .Z(rdata[33]));
Q_AN02 U489 ( .A0(n260), .A1(n227), .Z(rdata[32]));
Q_AN02 U490 ( .A0(n260), .A1(n228), .Z(rdata[31]));
Q_AN02 U491 ( .A0(n260), .A1(n229), .Z(rdata[30]));
Q_AN02 U492 ( .A0(n260), .A1(n230), .Z(rdata[29]));
Q_AN02 U493 ( .A0(n260), .A1(n231), .Z(rdata[28]));
Q_AN02 U494 ( .A0(n260), .A1(n232), .Z(rdata[27]));
Q_AN02 U495 ( .A0(n260), .A1(n233), .Z(rdata[26]));
Q_AN02 U496 ( .A0(n260), .A1(n234), .Z(rdata[25]));
Q_AN02 U497 ( .A0(n260), .A1(n235), .Z(rdata[24]));
Q_AN02 U498 ( .A0(n260), .A1(n236), .Z(rdata[23]));
Q_AN02 U499 ( .A0(n260), .A1(n237), .Z(rdata[22]));
Q_AN02 U500 ( .A0(n260), .A1(n238), .Z(rdata[21]));
Q_AN02 U501 ( .A0(n260), .A1(n239), .Z(rdata[20]));
Q_AN02 U502 ( .A0(n260), .A1(n240), .Z(rdata[19]));
Q_AN02 U503 ( .A0(n260), .A1(n241), .Z(rdata[18]));
Q_AN02 U504 ( .A0(n260), .A1(n242), .Z(rdata[17]));
Q_AN02 U505 ( .A0(n260), .A1(n243), .Z(rdata[16]));
Q_AN02 U506 ( .A0(n260), .A1(n244), .Z(rdata[15]));
Q_AN02 U507 ( .A0(n260), .A1(n245), .Z(rdata[14]));
Q_AN02 U508 ( .A0(n260), .A1(n246), .Z(rdata[13]));
Q_AN02 U509 ( .A0(n260), .A1(n247), .Z(rdata[12]));
Q_AN02 U510 ( .A0(n260), .A1(n248), .Z(rdata[11]));
Q_AN02 U511 ( .A0(n260), .A1(n249), .Z(rdata[10]));
Q_AN02 U512 ( .A0(n260), .A1(n250), .Z(rdata[9]));
Q_AN02 U513 ( .A0(n260), .A1(n251), .Z(rdata[8]));
Q_AN02 U514 ( .A0(n260), .A1(n252), .Z(rdata[7]));
Q_AN02 U515 ( .A0(n260), .A1(n253), .Z(rdata[6]));
Q_AN02 U516 ( .A0(n260), .A1(n254), .Z(rdata[5]));
Q_AN02 U517 ( .A0(n260), .A1(n255), .Z(rdata[4]));
Q_AN02 U518 ( .A0(n260), .A1(n256), .Z(rdata[3]));
Q_AN02 U519 ( .A0(n260), .A1(n257), .Z(rdata[2]));
Q_AN02 U520 ( .A0(n260), .A1(n258), .Z(rdata[1]));
Q_AN02 U521 ( .A0(n260), .A1(n259), .Z(rdata[0]));
Q_INV U522 ( .A(full), .Z(n2));
Q_AN02 U523 ( .A0(wen), .A1(n2), .Z(n3));
nx_fifo_ctrl_xcm36 \depth_n.fifo_ctrl ( .empty( empty), .full( full), 
	.used_slots( used_slots[2:0]), .free_slots( free_slots[2:0]), 
	.rptr( \depth_n.rptr [1:0]), .wptr( \depth_n.wptr [1:0]), 
	.underflow( \depth_n._zy_simnet_underflow_2_w$ ), .overflow( 
	\depth_n._zy_simnet_overflow_3_w$ ), .clk( clk), .rst_n( rst_n), 
	.wen( wen), .ren( ren), .clear( clear));
ixc_assign \depth_n._zz_strnp_1 ( overflow, 
	\depth_n._zy_simnet_overflow_3_w$ );
ixc_assign \depth_n._zz_strnp_0 ( underflow, 
	\depth_n._zy_simnet_underflow_2_w$ );
`ifdef CBV

reg [255:0] \depth_n.r_data  [3:0];
initial begin: U527
  integer i;
  for (i=3; i>=0; i=i-1) \depth_n.r_data [i] =
`ifdef CBV_MEM_INIT1
  {256{1'b1}};
`else
  256'b0;
`endif
end
reg [255:0] n526;
assign {n4, n5, n6, n7, n8, n9, n10,
n11, n12, n13, n14, n15, n16, n17, n18,
n19, n20, n21, n22, n23, n24, n25, n26,
n27, n28, n29, n30, n31, n32, n33, n34,
n35, n36, n37, n38, n39, n40, n41, n42,
n43, n44, n45, n46, n47, n48, n49, n50,
n51, n52, n53, n54, n55, n56, n57, n58,
n59, n60, n61, n62, n63, n64, n65, n66,
n67, n68, n69, n70, n71, n72, n73, n74,
n75, n76, n77, n78, n79, n80, n81, n82,
n83, n84, n85, n86, n87, n88, n89, n90,
n91, n92, n93, n94, n95, n96, n97, n98,
n99, n100, n101, n102, n103, n104, n105, n106,
n107, n108, n109, n110, n111, n112, n113, n114,
n115, n116, n117, n118, n119, n120, n121, n122,
n123, n124, n125, n126, n127, n128, n129, n130,
n131, n132, n133, n134, n135, n136, n137, n138,
n139, n140, n141, n142, n143, n144, n145, n146,
n147, n148, n149, n150, n151, n152, n153, n154,
n155, n156, n157, n158, n159, n160, n161, n162,
n163, n164, n165, n166, n167, n168, n169, n170,
n171, n172, n173, n174, n175, n176, n177, n178,
n179, n180, n181, n182, n183, n184, n185, n186,
n187, n188, n189, n190, n191, n192, n193, n194,
n195, n196, n197, n198, n199, n200, n201, n202,
n203, n204, n205, n206, n207, n208, n209, n210,
n211, n212, n213, n214, n215, n216, n217, n218,
n219, n220, n221, n222, n223, n224, n225, n226,
n227, n228, n229, n230, n231, n232, n233, n234,
n235, n236, n237, n238, n239, n240, n241, n242,
n243, n244, n245, n246, n247, n248, n249, n250,
n251, n252, n253, n254, n255, n256, n257, n258,
n259} = n526; 
always @(n268 or n267 or n524 or n523 or n522
 or n521 or n520 or n519 or n518 or n517 or n516 or n515 or n514
 or n513 or n512 or n511 or n510 or n509 or n508 or n507 or n506
 or n505 or n504 or n503 or n502 or n501 or n500 or n499 or n498
 or n497 or n496 or n495 or n494 or n493 or n492 or n491 or n490
 or n489 or n488 or n487 or n486 or n485 or n484 or n483 or n482
 or n481 or n480 or n479 or n478 or n477 or n476 or n475 or n474
 or n473 or n472 or n471 or n470 or n469 or n468 or n467 or n466
 or n465 or n464 or n463 or n462 or n461 or n460 or n459 or n458
 or n457 or n456 or n455 or n454 or n453 or n452 or n451 or n450
 or n449 or n448 or n447 or n446 or n445 or n444 or n443 or n442
 or n441 or n440 or n439 or n438 or n437 or n436 or n435 or n434
 or n433 or n432 or n431 or n430 or n429 or n428 or n427 or n426
 or n425 or n424 or n423 or n422 or n421 or n420 or n419 or n418
 or n417 or n416 or n415 or n414 or n413 or n412 or n411 or n410
 or n409 or n408 or n407 or n406 or n405 or n404 or n403 or n402
 or n401 or n400 or n399 or n398 or n397 or n396 or n395 or n394
 or n393 or n392 or n391 or n390 or n389 or n388 or n387 or n386
 or n385 or n384 or n383 or n382 or n381 or n380 or n379 or n378
 or n377 or n376 or n375 or n374 or n373 or n372 or n371 or n370
 or n369 or n368 or n367 or n366 or n365 or n364 or n363 or n362
 or n361 or n360 or n359 or n358 or n357 or n356 or n355 or n354
 or n353 or n352 or n351 or n350 or n349 or n348 or n347 or n346
 or n345 or n344 or n343 or n342 or n341 or n340 or n339 or n338
 or n337 or n336 or n335 or n334 or n333 or n332 or n331 or n330
 or n329 or n328 or n327 or n326 or n325 or n324 or n323 or n322
 or n321 or n320 or n319 or n318 or n317 or n316 or n315 or n314
 or n313 or n312 or n311 or n310 or n309 or n308 or n307 or n306
 or n305 or n304 or n303 or n302 or n301 or n300 or n299 or n298
 or n297 or n296 or n295 or n294 or n293 or n292 or n291 or n290
 or n289 or n288 or n287 or n286 or n285 or n284 or n283 or n282
 or n281 or n280 or n279 or n278 or n277 or n276 or n275 or n274
 or n273 or n272 or n271 or n270 or n269 or n266 or \depth_n.rptr [1] or \depth_n.rptr [0])
#0 begin
if (n266)
\depth_n.r_data [{n268, n267}] =
{n524, n523, n522, n521, n520,
 n519, n518, n517, n516, n515, n514, n513, n512,
 n511, n510, n509, n508, n507, n506, n505, n504,
 n503, n502, n501, n500, n499, n498, n497, n496,
 n495, n494, n493, n492, n491, n490, n489, n488,
 n487, n486, n485, n484, n483, n482, n481, n480,
 n479, n478, n477, n476, n475, n474, n473, n472,
 n471, n470, n469, n468, n467, n466, n465, n464,
 n463, n462, n461, n460, n459, n458, n457, n456,
 n455, n454, n453, n452, n451, n450, n449, n448,
 n447, n446, n445, n444, n443, n442, n441, n440,
 n439, n438, n437, n436, n435, n434, n433, n432,
 n431, n430, n429, n428, n427, n426, n425, n424,
 n423, n422, n421, n420, n419, n418, n417, n416,
 n415, n414, n413, n412, n411, n410, n409, n408,
 n407, n406, n405, n404, n403, n402, n401, n400,
 n399, n398, n397, n396, n395, n394, n393, n392,
 n391, n390, n389, n388, n387, n386, n385, n384,
 n383, n382, n381, n380, n379, n378, n377, n376,
 n375, n374, n373, n372, n371, n370, n369, n368,
 n367, n366, n365, n364, n363, n362, n361, n360,
 n359, n358, n357, n356, n355, n354, n353, n352,
 n351, n350, n349, n348, n347, n346, n345, n344,
 n343, n342, n341, n340, n339, n338, n337, n336,
 n335, n334, n333, n332, n331, n330, n329, n328,
 n327, n326, n325, n324, n323, n322, n321, n320,
 n319, n318, n317, n316, n315, n314, n313, n312,
 n311, n310, n309, n308, n307, n306, n305, n304,
 n303, n302, n301, n300, n299, n298, n297, n296,
 n295, n294, n293, n292, n291, n290, n289, n288,
 n287, n286, n285, n284, n283, n282, n281, n280,
 n279, n278, n277, n276, n275, n274, n273, n272,
 n271, n270, n269};
n526 = \depth_n.r_data [{\depth_n.rptr [1], \depth_n.rptr [0]}];
end
`else

MPW4X256 \depth_n.r_data  ( .A1(n268), .A0(n267), .DI255(n524), .DI254(n523), .DI253(n522), .DI252(n521),
 .DI251(n520), .DI250(n519), .DI249(n518), .DI248(n517), .DI247(n516), .DI246(n515), .DI245(n514), .DI244(n513),
 .DI243(n512), .DI242(n511), .DI241(n510), .DI240(n509), .DI239(n508), .DI238(n507), .DI237(n506), .DI236(n505),
 .DI235(n504), .DI234(n503), .DI233(n502), .DI232(n501), .DI231(n500), .DI230(n499), .DI229(n498), .DI228(n497),
 .DI227(n496), .DI226(n495), .DI225(n494), .DI224(n493), .DI223(n492), .DI222(n491), .DI221(n490), .DI220(n489),
 .DI219(n488), .DI218(n487), .DI217(n486), .DI216(n485), .DI215(n484), .DI214(n483), .DI213(n482), .DI212(n481),
 .DI211(n480), .DI210(n479), .DI209(n478), .DI208(n477), .DI207(n476), .DI206(n475), .DI205(n474), .DI204(n473),
 .DI203(n472), .DI202(n471), .DI201(n470), .DI200(n469), .DI199(n468), .DI198(n467), .DI197(n466), .DI196(n465),
 .DI195(n464), .DI194(n463), .DI193(n462), .DI192(n461), .DI191(n460), .DI190(n459), .DI189(n458), .DI188(n457),
 .DI187(n456), .DI186(n455), .DI185(n454), .DI184(n453), .DI183(n452), .DI182(n451), .DI181(n450), .DI180(n449),
 .DI179(n448), .DI178(n447), .DI177(n446), .DI176(n445), .DI175(n444), .DI174(n443), .DI173(n442), .DI172(n441),
 .DI171(n440), .DI170(n439), .DI169(n438), .DI168(n437), .DI167(n436), .DI166(n435), .DI165(n434), .DI164(n433),
 .DI163(n432), .DI162(n431), .DI161(n430), .DI160(n429), .DI159(n428), .DI158(n427), .DI157(n426), .DI156(n425),
 .DI155(n424), .DI154(n423), .DI153(n422), .DI152(n421), .DI151(n420), .DI150(n419), .DI149(n418), .DI148(n417),
 .DI147(n416), .DI146(n415), .DI145(n414), .DI144(n413), .DI143(n412), .DI142(n411), .DI141(n410), .DI140(n409),
 .DI139(n408), .DI138(n407), .DI137(n406), .DI136(n405), .DI135(n404), .DI134(n403), .DI133(n402), .DI132(n401),
 .DI131(n400), .DI130(n399), .DI129(n398), .DI128(n397), .DI127(n396), .DI126(n395), .DI125(n394), .DI124(n393),
 .DI123(n392), .DI122(n391), .DI121(n390), .DI120(n389), .DI119(n388), .DI118(n387), .DI117(n386), .DI116(n385),
 .DI115(n384), .DI114(n383), .DI113(n382), .DI112(n381), .DI111(n380), .DI110(n379), .DI109(n378), .DI108(n377),
 .DI107(n376), .DI106(n375), .DI105(n374), .DI104(n373), .DI103(n372), .DI102(n371), .DI101(n370), .DI100(n369),
 .DI99(n368), .DI98(n367), .DI97(n366), .DI96(n365), .DI95(n364), .DI94(n363), .DI93(n362), .DI92(n361),
 .DI91(n360), .DI90(n359), .DI89(n358), .DI88(n357), .DI87(n356), .DI86(n355), .DI85(n354), .DI84(n353),
 .DI83(n352), .DI82(n351), .DI81(n350), .DI80(n349), .DI79(n348), .DI78(n347), .DI77(n346), .DI76(n345),
 .DI75(n344), .DI74(n343), .DI73(n342), .DI72(n341), .DI71(n340), .DI70(n339), .DI69(n338), .DI68(n337),
 .DI67(n336), .DI66(n335), .DI65(n334), .DI64(n333), .DI63(n332), .DI62(n331), .DI61(n330), .DI60(n329),
 .DI59(n328), .DI58(n327), .DI57(n326), .DI56(n325), .DI55(n324), .DI54(n323), .DI53(n322), .DI52(n321),
 .DI51(n320), .DI50(n319), .DI49(n318), .DI48(n317), .DI47(n316), .DI46(n315), .DI45(n314), .DI44(n313),
 .DI43(n312), .DI42(n311), .DI41(n310), .DI40(n309), .DI39(n308), .DI38(n307), .DI37(n306), .DI36(n305),
 .DI35(n304), .DI34(n303), .DI33(n302), .DI32(n301), .DI31(n300), .DI30(n299), .DI29(n298), .DI28(n297),
 .DI27(n296), .DI26(n295), .DI25(n294), .DI24(n293), .DI23(n292), .DI22(n291), .DI21(n290), .DI20(n289),
 .DI19(n288), .DI18(n287), .DI17(n286), .DI16(n285), .DI15(n284), .DI14(n283), .DI13(n282), .DI12(n281),
 .DI11(n280), .DI10(n279), .DI9(n278), .DI8(n277), .DI7(n276), .DI6(n275), .DI5(n274), .DI4(n273),
 .DI3(n272), .DI2(n271), .DI1(n270), .DI0(n269), .WE(n266), .SYNC_IN(n525), .SYNC_OUT(n526));
// pragma CVASTRPROP INSTANCE "\depth_n.r_data " HDL_MEMORY_DECL "1 255 0 3 0"
MPR4X256 U528 ( .A1(\depth_n.rptr [1]), .A0(\depth_n.rptr [0]), .SYNC_IN(n526), .DO255(n4), .DO254(n5), .DO253(n6),
 .DO252(n7), .DO251(n8), .DO250(n9), .DO249(n10), .DO248(n11), .DO247(n12), .DO246(n13), .DO245(n14),
 .DO244(n15), .DO243(n16), .DO242(n17), .DO241(n18), .DO240(n19), .DO239(n20), .DO238(n21), .DO237(n22),
 .DO236(n23), .DO235(n24), .DO234(n25), .DO233(n26), .DO232(n27), .DO231(n28), .DO230(n29), .DO229(n30),
 .DO228(n31), .DO227(n32), .DO226(n33), .DO225(n34), .DO224(n35), .DO223(n36), .DO222(n37), .DO221(n38),
 .DO220(n39), .DO219(n40), .DO218(n41), .DO217(n42), .DO216(n43), .DO215(n44), .DO214(n45), .DO213(n46),
 .DO212(n47), .DO211(n48), .DO210(n49), .DO209(n50), .DO208(n51), .DO207(n52), .DO206(n53), .DO205(n54),
 .DO204(n55), .DO203(n56), .DO202(n57), .DO201(n58), .DO200(n59), .DO199(n60), .DO198(n61), .DO197(n62),
 .DO196(n63), .DO195(n64), .DO194(n65), .DO193(n66), .DO192(n67), .DO191(n68), .DO190(n69), .DO189(n70),
 .DO188(n71), .DO187(n72), .DO186(n73), .DO185(n74), .DO184(n75), .DO183(n76), .DO182(n77), .DO181(n78),
 .DO180(n79), .DO179(n80), .DO178(n81), .DO177(n82), .DO176(n83), .DO175(n84), .DO174(n85), .DO173(n86),
 .DO172(n87), .DO171(n88), .DO170(n89), .DO169(n90), .DO168(n91), .DO167(n92), .DO166(n93), .DO165(n94),
 .DO164(n95), .DO163(n96), .DO162(n97), .DO161(n98), .DO160(n99), .DO159(n100), .DO158(n101), .DO157(n102),
 .DO156(n103), .DO155(n104), .DO154(n105), .DO153(n106), .DO152(n107), .DO151(n108), .DO150(n109), .DO149(n110),
 .DO148(n111), .DO147(n112), .DO146(n113), .DO145(n114), .DO144(n115), .DO143(n116), .DO142(n117), .DO141(n118),
 .DO140(n119), .DO139(n120), .DO138(n121), .DO137(n122), .DO136(n123), .DO135(n124), .DO134(n125), .DO133(n126),
 .DO132(n127), .DO131(n128), .DO130(n129), .DO129(n130), .DO128(n131), .DO127(n132), .DO126(n133), .DO125(n134),
 .DO124(n135), .DO123(n136), .DO122(n137), .DO121(n138), .DO120(n139), .DO119(n140), .DO118(n141), .DO117(n142),
 .DO116(n143), .DO115(n144), .DO114(n145), .DO113(n146), .DO112(n147), .DO111(n148), .DO110(n149), .DO109(n150),
 .DO108(n151), .DO107(n152), .DO106(n153), .DO105(n154), .DO104(n155), .DO103(n156), .DO102(n157), .DO101(n158),
 .DO100(n159), .DO99(n160), .DO98(n161), .DO97(n162), .DO96(n163), .DO95(n164), .DO94(n165), .DO93(n166),
 .DO92(n167), .DO91(n168), .DO90(n169), .DO89(n170), .DO88(n171), .DO87(n172), .DO86(n173), .DO85(n174),
 .DO84(n175), .DO83(n176), .DO82(n177), .DO81(n178), .DO80(n179), .DO79(n180), .DO78(n181), .DO77(n182),
 .DO76(n183), .DO75(n184), .DO74(n185), .DO73(n186), .DO72(n187), .DO71(n188), .DO70(n189), .DO69(n190),
 .DO68(n191), .DO67(n192), .DO66(n193), .DO65(n194), .DO64(n195), .DO63(n196), .DO62(n197), .DO61(n198),
 .DO60(n199), .DO59(n200), .DO58(n201), .DO57(n202), .DO56(n203), .DO55(n204), .DO54(n205), .DO53(n206),
 .DO52(n207), .DO51(n208), .DO50(n209), .DO49(n210), .DO48(n211), .DO47(n212), .DO46(n213), .DO45(n214),
 .DO44(n215), .DO43(n216), .DO42(n217), .DO41(n218), .DO40(n219), .DO39(n220), .DO38(n221), .DO37(n222),
 .DO36(n223), .DO35(n224), .DO34(n225), .DO33(n226), .DO32(n227), .DO31(n228), .DO30(n229), .DO29(n230),
 .DO28(n231), .DO27(n232), .DO26(n233), .DO25(n234), .DO24(n235), .DO23(n236), .DO22(n237), .DO21(n238),
 .DO20(n239), .DO19(n240), .DO18(n241), .DO17(n242), .DO16(n243), .DO15(n244), .DO14(n245), .DO13(n246),
 .DO12(n247), .DO11(n248), .DO10(n249), .DO9(n250), .DO8(n251), .DO7(n252), .DO6(n253), .DO5(n254),
 .DO4(n255), .DO3(n256), .DO2(n257), .DO1(n258), .DO0(n259), .SYNC_OUT( ));
`endif
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "\depth_n.r_data  1 255 0 3 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "1"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_1 "0 genblk1  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_0 "-1 depth_n  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "depth_n.genblk1"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "depth_n"
endmodule
`ifdef CBV
`else
`ifdef MPW4X256_MPR4X256
`else
module MPW4X256( A1, A0, DI255, DI254, DI253, DI252, DI251,
 DI250, DI249, DI248, DI247, DI246, DI245, DI244, DI243,
 DI242, DI241, DI240, DI239, DI238, DI237, DI236, DI235,
 DI234, DI233, DI232, DI231, DI230, DI229, DI228, DI227,
 DI226, DI225, DI224, DI223, DI222, DI221, DI220, DI219,
 DI218, DI217, DI216, DI215, DI214, DI213, DI212, DI211,
 DI210, DI209, DI208, DI207, DI206, DI205, DI204, DI203,
 DI202, DI201, DI200, DI199, DI198, DI197, DI196, DI195,
 DI194, DI193, DI192, DI191, DI190, DI189, DI188, DI187,
 DI186, DI185, DI184, DI183, DI182, DI181, DI180, DI179,
 DI178, DI177, DI176, DI175, DI174, DI173, DI172, DI171,
 DI170, DI169, DI168, DI167, DI166, DI165, DI164, DI163,
 DI162, DI161, DI160, DI159, DI158, DI157, DI156, DI155,
 DI154, DI153, DI152, DI151, DI150, DI149, DI148, DI147,
 DI146, DI145, DI144, DI143, DI142, DI141, DI140, DI139,
 DI138, DI137, DI136, DI135, DI134, DI133, DI132, DI131,
 DI130, DI129, DI128, DI127, DI126, DI125, DI124, DI123,
 DI122, DI121, DI120, DI119, DI118, DI117, DI116, DI115,
 DI114, DI113, DI112, DI111, DI110, DI109, DI108, DI107,
 DI106, DI105, DI104, DI103, DI102, DI101, DI100, DI99,
 DI98, DI97, DI96, DI95, DI94, DI93, DI92, DI91,
 DI90, DI89, DI88, DI87, DI86, DI85, DI84, DI83,
 DI82, DI81, DI80, DI79, DI78, DI77, DI76, DI75,
 DI74, DI73, DI72, DI71, DI70, DI69, DI68, DI67,
 DI66, DI65, DI64, DI63, DI62, DI61, DI60, DI59,
 DI58, DI57, DI56, DI55, DI54, DI53, DI52, DI51,
 DI50, DI49, DI48, DI47, DI46, DI45, DI44, DI43,
 DI42, DI41, DI40, DI39, DI38, DI37, DI36, DI35,
 DI34, DI33, DI32, DI31, DI30, DI29, DI28, DI27,
 DI26, DI25, DI24, DI23, DI22, DI21, DI20, DI19,
 DI18, DI17, DI16, DI15, DI14, DI13, DI12, DI11,
 DI10, DI9, DI8, DI7, DI6, DI5, DI4, DI3,
 DI2, DI1, DI0, WE, SYNC_IN, SYNC_OUT);
input  A1, A0, DI255, DI254, DI253, DI252, DI251, DI250,
 DI249, DI248, DI247, DI246, DI245, DI244, DI243, DI242, DI241, DI240,
 DI239, DI238, DI237, DI236, DI235, DI234, DI233, DI232, DI231, DI230,
 DI229, DI228, DI227, DI226, DI225, DI224, DI223, DI222, DI221, DI220,
 DI219, DI218, DI217, DI216, DI215, DI214, DI213, DI212, DI211, DI210,
 DI209, DI208, DI207, DI206, DI205, DI204, DI203, DI202, DI201, DI200,
 DI199, DI198, DI197, DI196, DI195, DI194, DI193, DI192, DI191, DI190,
 DI189, DI188, DI187, DI186, DI185, DI184, DI183, DI182, DI181, DI180,
 DI179, DI178, DI177, DI176, DI175, DI174, DI173, DI172, DI171, DI170,
 DI169, DI168, DI167, DI166, DI165, DI164, DI163, DI162, DI161, DI160,
 DI159, DI158, DI157, DI156, DI155, DI154, DI153, DI152, DI151, DI150,
 DI149, DI148, DI147, DI146, DI145, DI144, DI143, DI142, DI141, DI140,
 DI139, DI138, DI137, DI136, DI135, DI134, DI133, DI132, DI131, DI130,
 DI129, DI128, DI127, DI126, DI125, DI124, DI123, DI122, DI121, DI120,
 DI119, DI118, DI117, DI116, DI115, DI114, DI113, DI112, DI111, DI110,
 DI109, DI108, DI107, DI106, DI105, DI104, DI103, DI102, DI101, DI100,
 DI99, DI98, DI97, DI96, DI95, DI94, DI93, DI92, DI91, DI90,
 DI89, DI88, DI87, DI86, DI85, DI84, DI83, DI82, DI81, DI80,
 DI79, DI78, DI77, DI76, DI75, DI74, DI73, DI72, DI71, DI70,
 DI69, DI68, DI67, DI66, DI65, DI64, DI63, DI62, DI61, DI60,
 DI59, DI58, DI57, DI56, DI55, DI54, DI53, DI52, DI51, DI50,
 DI49, DI48, DI47, DI46, DI45, DI44, DI43, DI42, DI41, DI40,
 DI39, DI38, DI37, DI36, DI35, DI34, DI33, DI32, DI31, DI30,
 DI29, DI28, DI27, DI26, DI25, DI24, DI23, DI22, DI21, DI20,
 DI19, DI18, DI17, DI16, DI15, DI14, DI13, DI12, DI11, DI10,
 DI9, DI8, DI7, DI6, DI5, DI4, DI3, DI2, DI1, DI0,
 WE, SYNC_IN;
output  SYNC_OUT;
endmodule
`ifdef _MPR4X256_
`else
module MPR4X256( A1, A0, SYNC_IN, DO255, DO254, DO253, DO252,
 DO251, DO250, DO249, DO248, DO247, DO246, DO245, DO244,
 DO243, DO242, DO241, DO240, DO239, DO238, DO237, DO236,
 DO235, DO234, DO233, DO232, DO231, DO230, DO229, DO228,
 DO227, DO226, DO225, DO224, DO223, DO222, DO221, DO220,
 DO219, DO218, DO217, DO216, DO215, DO214, DO213, DO212,
 DO211, DO210, DO209, DO208, DO207, DO206, DO205, DO204,
 DO203, DO202, DO201, DO200, DO199, DO198, DO197, DO196,
 DO195, DO194, DO193, DO192, DO191, DO190, DO189, DO188,
 DO187, DO186, DO185, DO184, DO183, DO182, DO181, DO180,
 DO179, DO178, DO177, DO176, DO175, DO174, DO173, DO172,
 DO171, DO170, DO169, DO168, DO167, DO166, DO165, DO164,
 DO163, DO162, DO161, DO160, DO159, DO158, DO157, DO156,
 DO155, DO154, DO153, DO152, DO151, DO150, DO149, DO148,
 DO147, DO146, DO145, DO144, DO143, DO142, DO141, DO140,
 DO139, DO138, DO137, DO136, DO135, DO134, DO133, DO132,
 DO131, DO130, DO129, DO128, DO127, DO126, DO125, DO124,
 DO123, DO122, DO121, DO120, DO119, DO118, DO117, DO116,
 DO115, DO114, DO113, DO112, DO111, DO110, DO109, DO108,
 DO107, DO106, DO105, DO104, DO103, DO102, DO101, DO100,
 DO99, DO98, DO97, DO96, DO95, DO94, DO93, DO92,
 DO91, DO90, DO89, DO88, DO87, DO86, DO85, DO84,
 DO83, DO82, DO81, DO80, DO79, DO78, DO77, DO76,
 DO75, DO74, DO73, DO72, DO71, DO70, DO69, DO68,
 DO67, DO66, DO65, DO64, DO63, DO62, DO61, DO60,
 DO59, DO58, DO57, DO56, DO55, DO54, DO53, DO52,
 DO51, DO50, DO49, DO48, DO47, DO46, DO45, DO44,
 DO43, DO42, DO41, DO40, DO39, DO38, DO37, DO36,
 DO35, DO34, DO33, DO32, DO31, DO30, DO29, DO28,
 DO27, DO26, DO25, DO24, DO23, DO22, DO21, DO20,
 DO19, DO18, DO17, DO16, DO15, DO14, DO13, DO12,
 DO11, DO10, DO9, DO8, DO7, DO6, DO5, DO4,
 DO3, DO2, DO1, DO0, SYNC_OUT);
input  A1, A0, SYNC_IN;
output  DO255, DO254, DO253, DO252, DO251, DO250, DO249, DO248,
 DO247, DO246, DO245, DO244, DO243, DO242, DO241, DO240, DO239, DO238,
 DO237, DO236, DO235, DO234, DO233, DO232, DO231, DO230, DO229, DO228,
 DO227, DO226, DO225, DO224, DO223, DO222, DO221, DO220, DO219, DO218,
 DO217, DO216, DO215, DO214, DO213, DO212, DO211, DO210, DO209, DO208,
 DO207, DO206, DO205, DO204, DO203, DO202, DO201, DO200, DO199, DO198,
 DO197, DO196, DO195, DO194, DO193, DO192, DO191, DO190, DO189, DO188,
 DO187, DO186, DO185, DO184, DO183, DO182, DO181, DO180, DO179, DO178,
 DO177, DO176, DO175, DO174, DO173, DO172, DO171, DO170, DO169, DO168,
 DO167, DO166, DO165, DO164, DO163, DO162, DO161, DO160, DO159, DO158,
 DO157, DO156, DO155, DO154, DO153, DO152, DO151, DO150, DO149, DO148,
 DO147, DO146, DO145, DO144, DO143, DO142, DO141, DO140, DO139, DO138,
 DO137, DO136, DO135, DO134, DO133, DO132, DO131, DO130, DO129, DO128,
 DO127, DO126, DO125, DO124, DO123, DO122, DO121, DO120, DO119, DO118,
 DO117, DO116, DO115, DO114, DO113, DO112, DO111, DO110, DO109, DO108,
 DO107, DO106, DO105, DO104, DO103, DO102, DO101, DO100, DO99, DO98,
 DO97, DO96, DO95, DO94, DO93, DO92, DO91, DO90, DO89, DO88,
 DO87, DO86, DO85, DO84, DO83, DO82, DO81, DO80, DO79, DO78,
 DO77, DO76, DO75, DO74, DO73, DO72, DO71, DO70, DO69, DO68,
 DO67, DO66, DO65, DO64, DO63, DO62, DO61, DO60, DO59, DO58,
 DO57, DO56, DO55, DO54, DO53, DO52, DO51, DO50, DO49, DO48,
 DO47, DO46, DO45, DO44, DO43, DO42, DO41, DO40, DO39, DO38,
 DO37, DO36, DO35, DO34, DO33, DO32, DO31, DO30, DO29, DO28,
 DO27, DO26, DO25, DO24, DO23, DO22, DO21, DO20, DO19, DO18,
 DO17, DO16, DO15, DO14, DO13, DO12, DO11, DO10, DO9, DO8,
 DO7, DO6, DO5, DO4, DO3, DO2, DO1, DO0, SYNC_OUT;
endmodule
`define _MPR4X256_
`endif
`define MPW4X256_MPR4X256
`endif
`endif
