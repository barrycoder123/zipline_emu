
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
`_2_ (* upf_always_on = 1 *) 
module xc_top_1 ;
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
wire fclk;
wire _ET3_COMPILER_RESERVED_NAME_DUTPI_APPLY_;
wire _ET3_COMPILER_RESERVED_NAME_LBRKER_ON_;
wire [63:0] _ET3_COMPILER_RESERVED_NAME_QT_CURR_EMUL_CYCLE_;
wire xc1xEcm;
wire callEmuPI;
wire [63:0] evalStepPI;
wire ckgHoldPI;
wire tbcHoldPI;
wire noOutputPI;
wire stopEmuPI;
wire oneStepPI;
wire stop1;
wire stop2;
wire stop4;
wire GFReset;
wire GFbusy;
wire svGFbusy;
wire otbGFbusy;
wire asyncCall;
wire svAsyncCall;
wire otbAsyncCall;
wire isfWait;
wire osfWait;
wire gfifoWait;
wire ecmHoldBusy;
wire sdlStop;
wire cpfStop;
wire eClk;
wire hasSFIFO;
wire hasGFIFO1;
wire hasGFIFO2;
wire hasPTX;
wire bpWait;
wire bWait;
wire eClkHold;
wire xpHold;
wire mpEnable;
wire ixcHoldClk;
wire oneFclkEval;
wire cakeCcEnable;
wire ptxBusy;
wire holdEcm;
wire bpHalt;
wire acHalt;
wire lockTrace;
wire [63:0] mioPOW_0;
wire [63:0] mioPOW_2;
wire mioPICnt;
wire [63:0] evalStepPIi;
wire callEmuPIi;
wire ckgHoldPIi;
wire stopEmuPIi;
wire oneStepPIi;
wire callEmuEv;
wire eventOn;
wire APPLY_PI;
wire lbrOnAll;
wire anyStop;
wire GFLock1;
wire GFLBfull;
wire GFGBfull;
wire GFBw;
wire GFGBfullBw;
wire GFAck;
wire [4:0] GF2LevelMask;
wire bClk;
wire sampleXpChg;
wire bClkRH;
wire bClkHold;
wire it_endBuf;
wire it_newBuf;
wire _zz_xmr0;
wire dummyW;
wire syncEn;
wire ecmOn;
wire ecmSync;
wire ecmNotSync;
wire holdEcmTb;
wire ptxHoldEcm;
wire [31:0] mcDelta;
wire mcp;
wire uClk;
`_2_ wire _ET3_COMPILER_RESERVED_NAME_ORION_INTERRUPT_;
`_2_ wire _ET3_COMPILER_RESERVED_NAME_DBI_APPLY_;
`_2_ wire _ET3_COMPILER_RESERVED_NAME_DBO_SAMPLE_;
`_2_ wire hotSwapOnPI;
`_2_ wire hssReset;
`_2_ wire sendPO;
`_2_ wire tbcPO;
`_2_ wire tbcPOd;
`_2_ wire stop1PO;
`_2_ wire stop1POd;
`_2_ wire stop2PO;
`_2_ wire stop2POd;
`_2_ wire stop4PO;
`_2_ wire stop4POd;
`_2_ wire stop3PO;
`_2_ wire stop3POd;
`_2_ wire it_newBufPO;
`_2_ wire stopSDLPO;
`_2_ wire stopEmuPO;
`_2_ wire stopCPFPO;
`_2_ wire [63:0] remStepPO;
`_2_ wire stop3;
`_2_ wire stop1R;
`_2_ wire stop2R;
`_2_ wire stop4R;
`_2_ wire stopSDL;
`_2_ wire sdlStopRply;
`_2_ wire sdlStopRplyD;
`_2_ wire sdlEnable;
`_2_ wire sdlHaltHwClk;
`_2_ wire GFbusyW;
`_2_ wire FTcallW;
`_2_ wire FvSimple2;
`_2_ wire [7:0] DccFrameCycle;
`_2_ wire [7:0] DccFrameMark;
`_2_ wire [7:0] dccFrameFill;
`_2_ wire noHoldOn;
`_2_ wire tbcEnable;
`_2_ wire hwClkEnable;
`_2_ wire hwClkDbgEn;
`_2_ wire hwClkDbg;
`_2_ wire hwClkDbgOn;
`_2_ wire hwClkDbgTime;
`_2_ wire [63:0] hwSimTime;
`_2_ wire [63:0] ixcSimTime;
`_2_ wire [31:0] hwClkDelay;
`_2_ wire bpOn;
`_2_ wire bpOnD;
`_2_ wire mpOn;
`_2_ wire ecmOne;
`_2_ wire [7:0] fclkPerEval;
`_2_ wire tbcHold;
`_2_ wire stopT;
`_2_ wire stopTL;
`_2_ wire stopTLd;
`_2_ wire clockMC;
`_2_ wire clockMCInit;
`_2_ wire evalOn;
`_2_ wire evalOnOrig;
`_2_ wire sfifoSyncMode;
`_2_ wire syncOtbChannels;
`_2_ wire [7:0] gfPushDly;
`_2_ wire [3:0] gfPushFill;
`_2_ wire bWaitExtend;
`_2_ wire lastDelta;
`_2_ wire callEmuR;
`_2_ wire evalOnC;
`_2_ wire evalOnD;
`_2_ wire [2:0] fcnt;
`_2_ wire eClkR;
`_2_ wire [7:0] evalOnDExt;
`_2_ wire [7:0] evalOnDCtl;
`_2_ wire simTimeOn;
`_2_ wire callEmu;
`_2_ wire nextTime;
`_2_ wire active;
`_2_ wire syncBp;
`_2_ wire [63:0] eCount;
`_2_ wire [63:0] bCount;
`_2_ wire [63:0] bpCount;
`_2_ wire [63:0] nbaCount;
`_2_ wire [63:0] evfCount;
`_2_ wire [31:0] aCount;
`_2_ wire [63:0] ixcHoldClkCnt;
`_2_ wire [63:0] ixcHoldSyncCnt;
`_2_ wire [63:0] ixcHoldEcmCnt;
`_2_ wire [63:0] fvSCount;
`_2_ wire [63:0] simTime;
`_2_ wire simTimeEnable;
`_2_ wire cakeUcEnable;
`_2_ wire initClock;
`_2_ wire holdEcmC;
`_2_ wire holdEcmD;
`_2_ wire xcReplayOn;
`_2_ wire xcRecordOn;
`_2_ wire evalOnSync;
`_2_ wire evalOnInt;
`_2_ wire evalOnIntD;
`_2_ wire [1:0] evalOnIntR;
`_2_ wire forceAbort;
`_2_ wire [15:0] bHaltCnt;
`_2_ wire [15:0] maxBpCycle;
`_2_ wire [15:0] aHaltCnt;
`_2_ wire [15:0] maxAcCycle;
`_2_ wire [3:0] lockTraceC;
`_2_ wire lockTraceOn;
`_2_ wire [63:0] lockTraceTime;
`_2_ wire xc_mioOn;
`_2_ wire mioPOCnt;
`_2_ wire tbcPOmio;
`_2_ wire [63:0] mioPIW_0;
`_2_ wire [63:0] mioPIW_1;
`_2_ wire mioPICntd;
`_2_ wire [63:0] evalStepPImio;
`_2_ wire callEmuPImio;
`_2_ wire ckgHoldPImio;
`_2_ wire oneStepPImio;
`_2_ wire [63:0] nextDutTimeS;
`_2_ wire callEmuWaitC;
`_2_ wire callEmuWait;
`_2_ wire callEmuWaitN;
`_2_ wire callEmuPre;
`_2_ wire applyPiR;
`_2_ wire dbiEvent;
`_2_ wire FvUseOnly;
`_2_ wire FvUseOnlyR;
`_2_ wire eventOnR;
`_2_ wire mpSampleOv;
`_2_ wire lbrOn;
`_2_ wire gfifoOff;
`_2_ wire gfifoAsyncOff;
`_2_ wire GFLock2;
`_2_ wire GFGBfullBwD;
`_2_ wire GFLBfullD;
`_2_ wire tbcPOReg;
`_2_ wire GFLock2R;
`_2_ wire SFIFOLock;
`_2_ wire [7:0] gfifoAckWait;
`_2_ wire asyncBusy;
`_2_ wire GFbusyD;
`_2_ wire GFbusyD2;
`_2_ wire [4:0] tbcPODly;
`_2_ wire tbcPORdy;
`_2_ wire [1:0] tbcPOState;
`_2_ wire [1:0] tbcPOStateN;
`_2_ wire SFIFOLock2;
`_2_ wire bClkR;
`_2_ wire sampleXpV;
`_2_ wire [1:0] bpSt;
`_2_ wire bClkHoldD;
`_2_ wire ixcHoldClkR;
`_2_ wire intr;
`_2_ wire it_capture;
`_2_ wire it_replay;
`_2_ wire dummyR;
`_2_ wire hwClkHalt;
`_2_ wire sdlHaltHwClkR;
`_2_ wire [63:0] gfifoGBfullCnt;
`_2_ wire [63:0] gfifoLBfullCnt;
`_2_ wire [63:0] gfifoTBsyncCnt;
`_2_ wire [15:0] maxFck2Sync;
`_2_ wire [15:0] maxGfifo2Sync;
`_2_ wire [15:0] Fck2Sync;
`_2_ wire [15:0] Gfifo2Sync;
`_2_ wire ptxStop;
`_2_ wire ecmOnD;
`_2_ wire ecmNotSyncD;
`_2_ wire holdEcmPtxOn;
`_2_ wire holdEcmSync;
`_2_ wire uClkT;
`_2_ wire dccState;
`_2_ wire [63:0] nextDutTimeP;
`_2_ wire [63:0] fclkCntr;
`_2_ wire [63:0] uClkCntr;
`_2_ wire [63:0] uClkErrTime;
supply1 n3552;
supply0 n4029;
supply1 n4030;
supply0 n4031;
supply1 n4032;
Q_BUF U0 ( .A(n4029), .Z(xc1xEcm));
Q_BUF U1 ( .A(n3552), .Z(_ET3_COMPILER_RESERVED_NAME_DUTPI_APPLY_));
Q_BUF U2 ( .A(n4029), .Z(mioPOW_2[63]));
Q_BUF U3 ( .A(n4029), .Z(mioPOW_2[62]));
Q_BUF U4 ( .A(n4029), .Z(mioPOW_2[61]));
Q_BUF U5 ( .A(n4029), .Z(mioPOW_2[60]));
Q_BUF U6 ( .A(n4029), .Z(mioPOW_2[59]));
Q_BUF U7 ( .A(n4029), .Z(mioPOW_2[58]));
Q_BUF U8 ( .A(n4029), .Z(mioPOW_2[57]));
Q_BUF U9 ( .A(n4029), .Z(mioPOW_2[56]));
Q_BUF U10 ( .A(n4029), .Z(mioPOW_2[55]));
Q_BUF U11 ( .A(n4029), .Z(mioPOW_2[54]));
Q_BUF U12 ( .A(n4029), .Z(mioPOW_2[53]));
Q_BUF U13 ( .A(n4029), .Z(mioPOW_2[52]));
Q_BUF U14 ( .A(n4029), .Z(mioPOW_2[51]));
Q_BUF U15 ( .A(n4029), .Z(mioPOW_2[50]));
Q_BUF U16 ( .A(n4029), .Z(mioPOW_2[49]));
Q_BUF U17 ( .A(n4029), .Z(mioPOW_2[48]));
Q_BUF U18 ( .A(n4029), .Z(mioPOW_2[47]));
Q_BUF U19 ( .A(n4029), .Z(mioPOW_2[46]));
Q_BUF U20 ( .A(n4029), .Z(mioPOW_2[45]));
Q_BUF U21 ( .A(n4029), .Z(mioPOW_2[44]));
Q_BUF U22 ( .A(n4029), .Z(mioPOW_2[43]));
Q_BUF U23 ( .A(n4029), .Z(mioPOW_2[42]));
Q_BUF U24 ( .A(n4029), .Z(mioPOW_2[41]));
Q_BUF U25 ( .A(n4029), .Z(mioPOW_2[40]));
Q_BUF U26 ( .A(n4029), .Z(mioPOW_2[39]));
Q_BUF U27 ( .A(n4029), .Z(mioPOW_2[38]));
Q_BUF U28 ( .A(n4029), .Z(mioPOW_2[37]));
Q_BUF U29 ( .A(n4029), .Z(mioPOW_2[36]));
Q_BUF U30 ( .A(n4029), .Z(mioPOW_2[35]));
Q_BUF U31 ( .A(n4029), .Z(mioPOW_2[34]));
Q_BUF U32 ( .A(n4029), .Z(mioPOW_2[33]));
Q_BUF U33 ( .A(n4029), .Z(mioPOW_2[32]));
Q_BUF U34 ( .A(n4029), .Z(mioPOW_2[31]));
Q_BUF U35 ( .A(n4029), .Z(mioPOW_2[30]));
Q_BUF U36 ( .A(n4029), .Z(mioPOW_2[29]));
Q_BUF U37 ( .A(n4029), .Z(mioPOW_2[28]));
Q_BUF U38 ( .A(n4029), .Z(mioPOW_2[27]));
Q_BUF U39 ( .A(n4029), .Z(mioPOW_2[26]));
Q_BUF U40 ( .A(n4029), .Z(mioPOW_2[25]));
Q_BUF U41 ( .A(n4029), .Z(mioPOW_2[24]));
Q_BUF U42 ( .A(n4029), .Z(mioPOW_2[23]));
Q_BUF U43 ( .A(n4029), .Z(mioPOW_2[22]));
Q_BUF U44 ( .A(n4029), .Z(mioPOW_2[21]));
Q_BUF U45 ( .A(n4029), .Z(mioPOW_2[20]));
Q_BUF U46 ( .A(n4029), .Z(mioPOW_2[19]));
Q_BUF U47 ( .A(n4029), .Z(mioPOW_2[18]));
Q_BUF U48 ( .A(n4029), .Z(mioPOW_2[17]));
Q_BUF U49 ( .A(n4029), .Z(mioPOW_2[16]));
Q_BUF U50 ( .A(n4029), .Z(mioPOW_2[15]));
Q_BUF U51 ( .A(n4029), .Z(mioPOW_2[14]));
Q_BUF U52 ( .A(n4029), .Z(mioPOW_2[13]));
Q_BUF U53 ( .A(n4029), .Z(mioPOW_2[12]));
Q_BUF U54 ( .A(n4029), .Z(mioPOW_2[11]));
Q_BUF U55 ( .A(n4029), .Z(mioPOW_2[10]));
Q_BUF U56 ( .A(n4029), .Z(mioPOW_2[9]));
Q_BUF U57 ( .A(lockTraceC[3]), .Z(lockTrace));
Q_BUF U58 ( .A(mioPOCnt), .Z(mioPOW_0[63]));
Q_BUF U59 ( .A(evalStepPIi[63]), .Z(ixc_time.nextTbTime[63]));
Q_BUF U60 ( .A(evalStepPIi[62]), .Z(ixc_time.nextTbTime[62]));
Q_BUF U61 ( .A(evalStepPIi[61]), .Z(ixc_time.nextTbTime[61]));
Q_BUF U62 ( .A(evalStepPIi[60]), .Z(ixc_time.nextTbTime[60]));
Q_BUF U63 ( .A(evalStepPIi[59]), .Z(ixc_time.nextTbTime[59]));
Q_BUF U64 ( .A(evalStepPIi[58]), .Z(ixc_time.nextTbTime[58]));
Q_BUF U65 ( .A(evalStepPIi[57]), .Z(ixc_time.nextTbTime[57]));
Q_BUF U66 ( .A(evalStepPIi[56]), .Z(ixc_time.nextTbTime[56]));
Q_BUF U67 ( .A(evalStepPIi[55]), .Z(ixc_time.nextTbTime[55]));
Q_BUF U68 ( .A(evalStepPIi[54]), .Z(ixc_time.nextTbTime[54]));
Q_BUF U69 ( .A(evalStepPIi[53]), .Z(ixc_time.nextTbTime[53]));
Q_BUF U70 ( .A(evalStepPIi[52]), .Z(ixc_time.nextTbTime[52]));
Q_BUF U71 ( .A(evalStepPIi[51]), .Z(ixc_time.nextTbTime[51]));
Q_BUF U72 ( .A(evalStepPIi[50]), .Z(ixc_time.nextTbTime[50]));
Q_BUF U73 ( .A(evalStepPIi[49]), .Z(ixc_time.nextTbTime[49]));
Q_BUF U74 ( .A(evalStepPIi[48]), .Z(ixc_time.nextTbTime[48]));
Q_BUF U75 ( .A(evalStepPIi[47]), .Z(ixc_time.nextTbTime[47]));
Q_BUF U76 ( .A(evalStepPIi[46]), .Z(ixc_time.nextTbTime[46]));
Q_BUF U77 ( .A(evalStepPIi[45]), .Z(ixc_time.nextTbTime[45]));
Q_BUF U78 ( .A(evalStepPIi[44]), .Z(ixc_time.nextTbTime[44]));
Q_BUF U79 ( .A(evalStepPIi[43]), .Z(ixc_time.nextTbTime[43]));
Q_BUF U80 ( .A(evalStepPIi[42]), .Z(ixc_time.nextTbTime[42]));
Q_BUF U81 ( .A(evalStepPIi[41]), .Z(ixc_time.nextTbTime[41]));
Q_BUF U82 ( .A(evalStepPIi[40]), .Z(ixc_time.nextTbTime[40]));
Q_BUF U83 ( .A(evalStepPIi[39]), .Z(ixc_time.nextTbTime[39]));
Q_BUF U84 ( .A(evalStepPIi[38]), .Z(ixc_time.nextTbTime[38]));
Q_BUF U85 ( .A(evalStepPIi[37]), .Z(ixc_time.nextTbTime[37]));
Q_BUF U86 ( .A(evalStepPIi[36]), .Z(ixc_time.nextTbTime[36]));
Q_BUF U87 ( .A(evalStepPIi[35]), .Z(ixc_time.nextTbTime[35]));
Q_BUF U88 ( .A(evalStepPIi[34]), .Z(ixc_time.nextTbTime[34]));
Q_BUF U89 ( .A(evalStepPIi[33]), .Z(ixc_time.nextTbTime[33]));
Q_BUF U90 ( .A(evalStepPIi[32]), .Z(ixc_time.nextTbTime[32]));
Q_BUF U91 ( .A(evalStepPIi[31]), .Z(ixc_time.nextTbTime[31]));
Q_BUF U92 ( .A(evalStepPIi[30]), .Z(ixc_time.nextTbTime[30]));
Q_BUF U93 ( .A(evalStepPIi[29]), .Z(ixc_time.nextTbTime[29]));
Q_BUF U94 ( .A(evalStepPIi[28]), .Z(ixc_time.nextTbTime[28]));
Q_BUF U95 ( .A(evalStepPIi[27]), .Z(ixc_time.nextTbTime[27]));
Q_BUF U96 ( .A(evalStepPIi[26]), .Z(ixc_time.nextTbTime[26]));
Q_BUF U97 ( .A(evalStepPIi[25]), .Z(ixc_time.nextTbTime[25]));
Q_BUF U98 ( .A(evalStepPIi[24]), .Z(ixc_time.nextTbTime[24]));
Q_BUF U99 ( .A(evalStepPIi[23]), .Z(ixc_time.nextTbTime[23]));
Q_BUF U100 ( .A(evalStepPIi[22]), .Z(ixc_time.nextTbTime[22]));
Q_BUF U101 ( .A(evalStepPIi[21]), .Z(ixc_time.nextTbTime[21]));
Q_BUF U102 ( .A(evalStepPIi[20]), .Z(ixc_time.nextTbTime[20]));
Q_BUF U103 ( .A(evalStepPIi[19]), .Z(ixc_time.nextTbTime[19]));
Q_BUF U104 ( .A(evalStepPIi[18]), .Z(ixc_time.nextTbTime[18]));
Q_BUF U105 ( .A(evalStepPIi[17]), .Z(ixc_time.nextTbTime[17]));
Q_BUF U106 ( .A(evalStepPIi[16]), .Z(ixc_time.nextTbTime[16]));
Q_BUF U107 ( .A(evalStepPIi[15]), .Z(ixc_time.nextTbTime[15]));
Q_BUF U108 ( .A(evalStepPIi[14]), .Z(ixc_time.nextTbTime[14]));
Q_BUF U109 ( .A(evalStepPIi[13]), .Z(ixc_time.nextTbTime[13]));
Q_BUF U110 ( .A(evalStepPIi[12]), .Z(ixc_time.nextTbTime[12]));
Q_BUF U111 ( .A(evalStepPIi[11]), .Z(ixc_time.nextTbTime[11]));
Q_BUF U112 ( .A(evalStepPIi[10]), .Z(ixc_time.nextTbTime[10]));
Q_BUF U113 ( .A(evalStepPIi[9]), .Z(ixc_time.nextTbTime[9]));
Q_BUF U114 ( .A(evalStepPIi[8]), .Z(ixc_time.nextTbTime[8]));
Q_BUF U115 ( .A(evalStepPIi[7]), .Z(ixc_time.nextTbTime[7]));
Q_BUF U116 ( .A(evalStepPIi[6]), .Z(ixc_time.nextTbTime[6]));
Q_BUF U117 ( .A(evalStepPIi[5]), .Z(ixc_time.nextTbTime[5]));
Q_BUF U118 ( .A(evalStepPIi[4]), .Z(ixc_time.nextTbTime[4]));
Q_BUF U119 ( .A(evalStepPIi[3]), .Z(ixc_time.nextTbTime[3]));
Q_BUF U120 ( .A(evalStepPIi[2]), .Z(ixc_time.nextTbTime[2]));
Q_BUF U121 ( .A(evalStepPIi[1]), .Z(ixc_time.nextTbTime[1]));
Q_BUF U122 ( .A(evalStepPIi[0]), .Z(ixc_time.nextTbTime[0]));
Q_BUF U123 ( .A(sendPO), .Z(mioPOW_2[0]));
Q_ASSIGN U124 ( .B(GFBw), .A(bClkHold));
Q_BUF U125 ( .A(stopSDLPO), .Z(mioPOW_2[7]));
Q_BUF U126 ( .A(stopCPFPO), .Z(mioPOW_2[8]));
Q_BUF U127 ( .A(eventOnR), .Z(eventOn));
Q_BUF U128 ( .A(stop1PO), .Z(mioPOW_2[2]));
Q_BUF U129 ( .A(stop2PO), .Z(mioPOW_2[3]));
Q_BUF U130 ( .A(stop4PO), .Z(mioPOW_2[5]));
Q_BUF U131 ( .A(stop3PO), .Z(mioPOW_2[4]));
Q_BUF U132 ( .A(stopEmuPIi), .Z(stopEmuPO));
Q_BUF U133 ( .A(remStepPO[62]), .Z(mioPOW_0[62]));
Q_BUF U134 ( .A(remStepPO[61]), .Z(mioPOW_0[61]));
Q_BUF U135 ( .A(remStepPO[60]), .Z(mioPOW_0[60]));
Q_BUF U136 ( .A(remStepPO[59]), .Z(mioPOW_0[59]));
Q_BUF U137 ( .A(remStepPO[58]), .Z(mioPOW_0[58]));
Q_BUF U138 ( .A(remStepPO[57]), .Z(mioPOW_0[57]));
Q_BUF U139 ( .A(remStepPO[56]), .Z(mioPOW_0[56]));
Q_BUF U140 ( .A(remStepPO[55]), .Z(mioPOW_0[55]));
Q_BUF U141 ( .A(remStepPO[54]), .Z(mioPOW_0[54]));
Q_BUF U142 ( .A(remStepPO[53]), .Z(mioPOW_0[53]));
Q_BUF U143 ( .A(remStepPO[52]), .Z(mioPOW_0[52]));
Q_BUF U144 ( .A(remStepPO[51]), .Z(mioPOW_0[51]));
Q_BUF U145 ( .A(remStepPO[50]), .Z(mioPOW_0[50]));
Q_BUF U146 ( .A(remStepPO[49]), .Z(mioPOW_0[49]));
Q_BUF U147 ( .A(remStepPO[48]), .Z(mioPOW_0[48]));
Q_BUF U148 ( .A(remStepPO[47]), .Z(mioPOW_0[47]));
Q_BUF U149 ( .A(remStepPO[46]), .Z(mioPOW_0[46]));
Q_BUF U150 ( .A(remStepPO[45]), .Z(mioPOW_0[45]));
Q_BUF U151 ( .A(remStepPO[44]), .Z(mioPOW_0[44]));
Q_BUF U152 ( .A(remStepPO[43]), .Z(mioPOW_0[43]));
Q_BUF U153 ( .A(remStepPO[42]), .Z(mioPOW_0[42]));
Q_BUF U154 ( .A(remStepPO[41]), .Z(mioPOW_0[41]));
Q_BUF U155 ( .A(remStepPO[40]), .Z(mioPOW_0[40]));
Q_BUF U156 ( .A(remStepPO[39]), .Z(mioPOW_0[39]));
Q_BUF U157 ( .A(remStepPO[38]), .Z(mioPOW_0[38]));
Q_BUF U158 ( .A(remStepPO[37]), .Z(mioPOW_0[37]));
Q_BUF U159 ( .A(remStepPO[36]), .Z(mioPOW_0[36]));
Q_BUF U160 ( .A(remStepPO[35]), .Z(mioPOW_0[35]));
Q_BUF U161 ( .A(remStepPO[34]), .Z(mioPOW_0[34]));
Q_BUF U162 ( .A(remStepPO[33]), .Z(mioPOW_0[33]));
Q_BUF U163 ( .A(remStepPO[32]), .Z(mioPOW_0[32]));
Q_BUF U164 ( .A(remStepPO[31]), .Z(mioPOW_0[31]));
Q_BUF U165 ( .A(remStepPO[30]), .Z(mioPOW_0[30]));
Q_BUF U166 ( .A(remStepPO[29]), .Z(mioPOW_0[29]));
Q_BUF U167 ( .A(remStepPO[28]), .Z(mioPOW_0[28]));
Q_BUF U168 ( .A(remStepPO[27]), .Z(mioPOW_0[27]));
Q_BUF U169 ( .A(remStepPO[26]), .Z(mioPOW_0[26]));
Q_BUF U170 ( .A(remStepPO[25]), .Z(mioPOW_0[25]));
Q_BUF U171 ( .A(remStepPO[24]), .Z(mioPOW_0[24]));
Q_BUF U172 ( .A(remStepPO[23]), .Z(mioPOW_0[23]));
Q_BUF U173 ( .A(remStepPO[22]), .Z(mioPOW_0[22]));
Q_BUF U174 ( .A(remStepPO[21]), .Z(mioPOW_0[21]));
Q_BUF U175 ( .A(remStepPO[20]), .Z(mioPOW_0[20]));
Q_BUF U176 ( .A(remStepPO[19]), .Z(mioPOW_0[19]));
Q_BUF U177 ( .A(remStepPO[18]), .Z(mioPOW_0[18]));
Q_BUF U178 ( .A(remStepPO[17]), .Z(mioPOW_0[17]));
Q_BUF U179 ( .A(remStepPO[16]), .Z(mioPOW_0[16]));
Q_BUF U180 ( .A(remStepPO[15]), .Z(mioPOW_0[15]));
Q_BUF U181 ( .A(remStepPO[14]), .Z(mioPOW_0[14]));
Q_BUF U182 ( .A(remStepPO[13]), .Z(mioPOW_0[13]));
Q_BUF U183 ( .A(remStepPO[12]), .Z(mioPOW_0[12]));
Q_BUF U184 ( .A(remStepPO[11]), .Z(mioPOW_0[11]));
Q_BUF U185 ( .A(remStepPO[10]), .Z(mioPOW_0[10]));
Q_BUF U186 ( .A(remStepPO[9]), .Z(mioPOW_0[9]));
Q_BUF U187 ( .A(remStepPO[8]), .Z(mioPOW_0[8]));
Q_BUF U188 ( .A(remStepPO[7]), .Z(mioPOW_0[7]));
Q_BUF U189 ( .A(remStepPO[6]), .Z(mioPOW_0[6]));
Q_BUF U190 ( .A(remStepPO[5]), .Z(mioPOW_0[5]));
Q_BUF U191 ( .A(remStepPO[4]), .Z(mioPOW_0[4]));
Q_BUF U192 ( .A(remStepPO[3]), .Z(mioPOW_0[3]));
Q_BUF U193 ( .A(remStepPO[2]), .Z(mioPOW_0[2]));
Q_BUF U194 ( .A(remStepPO[1]), .Z(mioPOW_0[1]));
Q_BUF U195 ( .A(remStepPO[0]), .Z(mioPOW_0[0]));
Q_BUF U196 ( .A(tbcPO), .Z(mioPOW_2[1]));
Q_BUF U197 ( .A(SFIFOLock), .Z(SFIFOLock2));
Q_BUF U198 ( .A(it_newBufPO), .Z(mioPOW_2[6]));
Q_ASSIGN U199 ( .B(mioPIW_1[0]), .A(mioPICnt));
Q_BUF U200 ( .A(callEmu), .Z(callEmuPre));
Q_BUF U201 ( .A(n4029), .Z(n1));
Q_AN02 U202 ( .A0(n3551), .A1(initClock), .Z(n2));
Q_AN02 U203 ( .A0(n2783), .A1(n2530), .Z(n3));
Q_AN02 U204 ( .A0(n2659), .A1(evalOn), .Z(n4));
Q_AN02 U205 ( .A0(n2406), .A1(n1958), .Z(n5));
Q_AN02 U206 ( .A0(n2282), .A1(n1957), .Z(n6));
Q_AN02 U207 ( .A0(n2158), .A1(n1956), .Z(n7));
Q_AN02 U208 ( .A0(n1832), .A1(n1766), .Z(n8));
Q_AN02 U209 ( .A0(n1706), .A1(n1671), .Z(n9));
Q_AN02 U210 ( .A0(n1508), .A1(hwClkDbgOn), .Z(n10));
Q_AN02 U211 ( .A0(n908), .A1(n646), .Z(n11));
Q_AN02 U212 ( .A0(n1280), .A1(n645), .Z(n12));
Q_AN02 U213 ( .A0(n1156), .A1(n644), .Z(n13));
Q_AN02 U214 ( .A0(n1032), .A1(n643), .Z(n14));
Q_AN02 U215 ( .A0(n81), .A1(initClock), .Z(n15));
Q_XNR3 U216 ( .A0(n3981), .A1(ixc_time.nextDutTime[31]), .A2(nextDutTimeP[31]), .Z(mcDelta[31]));
Q_XOR2 U217 ( .A0(initClock), .A1(fclkCntr[0]), .Z(n17));
Q_FDP0UA U218 ( .D(n17), .QTFCLK( ), .Q(fclkCntr[0]));
Q_MX02 U219 ( .S(initClock), .A0(fclkCntr[1]), .A1(n204), .Z(n18));
Q_FDP0UA U220 ( .D(n18), .QTFCLK( ), .Q(fclkCntr[1]));
Q_MX02 U221 ( .S(initClock), .A0(fclkCntr[2]), .A1(n202), .Z(n19));
Q_FDP0UA U222 ( .D(n19), .QTFCLK( ), .Q(fclkCntr[2]));
Q_MX02 U223 ( .S(initClock), .A0(fclkCntr[3]), .A1(n200), .Z(n20));
Q_FDP0UA U224 ( .D(n20), .QTFCLK( ), .Q(fclkCntr[3]));
Q_MX02 U225 ( .S(initClock), .A0(fclkCntr[4]), .A1(n198), .Z(n21));
Q_FDP0UA U226 ( .D(n21), .QTFCLK( ), .Q(fclkCntr[4]));
Q_MX02 U227 ( .S(initClock), .A0(fclkCntr[5]), .A1(n196), .Z(n22));
Q_FDP0UA U228 ( .D(n22), .QTFCLK( ), .Q(fclkCntr[5]));
Q_MX02 U229 ( .S(initClock), .A0(fclkCntr[6]), .A1(n194), .Z(n23));
Q_FDP0UA U230 ( .D(n23), .QTFCLK( ), .Q(fclkCntr[6]));
Q_MX02 U231 ( .S(initClock), .A0(fclkCntr[7]), .A1(n192), .Z(n24));
Q_FDP0UA U232 ( .D(n24), .QTFCLK( ), .Q(fclkCntr[7]));
Q_MX02 U233 ( .S(initClock), .A0(fclkCntr[8]), .A1(n190), .Z(n25));
Q_FDP0UA U234 ( .D(n25), .QTFCLK( ), .Q(fclkCntr[8]));
Q_MX02 U235 ( .S(initClock), .A0(fclkCntr[9]), .A1(n188), .Z(n26));
Q_FDP0UA U236 ( .D(n26), .QTFCLK( ), .Q(fclkCntr[9]));
Q_MX02 U237 ( .S(initClock), .A0(fclkCntr[10]), .A1(n186), .Z(n27));
Q_FDP0UA U238 ( .D(n27), .QTFCLK( ), .Q(fclkCntr[10]));
Q_MX02 U239 ( .S(initClock), .A0(fclkCntr[11]), .A1(n184), .Z(n28));
Q_FDP0UA U240 ( .D(n28), .QTFCLK( ), .Q(fclkCntr[11]));
Q_MX02 U241 ( .S(initClock), .A0(fclkCntr[12]), .A1(n182), .Z(n29));
Q_FDP0UA U242 ( .D(n29), .QTFCLK( ), .Q(fclkCntr[12]));
Q_MX02 U243 ( .S(initClock), .A0(fclkCntr[13]), .A1(n180), .Z(n30));
Q_FDP0UA U244 ( .D(n30), .QTFCLK( ), .Q(fclkCntr[13]));
Q_MX02 U245 ( .S(initClock), .A0(fclkCntr[14]), .A1(n178), .Z(n31));
Q_FDP0UA U246 ( .D(n31), .QTFCLK( ), .Q(fclkCntr[14]));
Q_MX02 U247 ( .S(initClock), .A0(fclkCntr[15]), .A1(n176), .Z(n32));
Q_FDP0UA U248 ( .D(n32), .QTFCLK( ), .Q(fclkCntr[15]));
Q_MX02 U249 ( .S(initClock), .A0(fclkCntr[16]), .A1(n174), .Z(n33));
Q_FDP0UA U250 ( .D(n33), .QTFCLK( ), .Q(fclkCntr[16]));
Q_MX02 U251 ( .S(initClock), .A0(fclkCntr[17]), .A1(n172), .Z(n34));
Q_FDP0UA U252 ( .D(n34), .QTFCLK( ), .Q(fclkCntr[17]));
Q_MX02 U253 ( .S(initClock), .A0(fclkCntr[18]), .A1(n170), .Z(n35));
Q_FDP0UA U254 ( .D(n35), .QTFCLK( ), .Q(fclkCntr[18]));
Q_MX02 U255 ( .S(initClock), .A0(fclkCntr[19]), .A1(n168), .Z(n36));
Q_FDP0UA U256 ( .D(n36), .QTFCLK( ), .Q(fclkCntr[19]));
Q_MX02 U257 ( .S(initClock), .A0(fclkCntr[20]), .A1(n166), .Z(n37));
Q_FDP0UA U258 ( .D(n37), .QTFCLK( ), .Q(fclkCntr[20]));
Q_MX02 U259 ( .S(initClock), .A0(fclkCntr[21]), .A1(n164), .Z(n38));
Q_FDP0UA U260 ( .D(n38), .QTFCLK( ), .Q(fclkCntr[21]));
Q_MX02 U261 ( .S(initClock), .A0(fclkCntr[22]), .A1(n162), .Z(n39));
Q_FDP0UA U262 ( .D(n39), .QTFCLK( ), .Q(fclkCntr[22]));
Q_MX02 U263 ( .S(initClock), .A0(fclkCntr[23]), .A1(n160), .Z(n40));
Q_FDP0UA U264 ( .D(n40), .QTFCLK( ), .Q(fclkCntr[23]));
Q_MX02 U265 ( .S(initClock), .A0(fclkCntr[24]), .A1(n158), .Z(n41));
Q_FDP0UA U266 ( .D(n41), .QTFCLK( ), .Q(fclkCntr[24]));
Q_MX02 U267 ( .S(initClock), .A0(fclkCntr[25]), .A1(n156), .Z(n42));
Q_FDP0UA U268 ( .D(n42), .QTFCLK( ), .Q(fclkCntr[25]));
Q_MX02 U269 ( .S(initClock), .A0(fclkCntr[26]), .A1(n154), .Z(n43));
Q_FDP0UA U270 ( .D(n43), .QTFCLK( ), .Q(fclkCntr[26]));
Q_MX02 U271 ( .S(initClock), .A0(fclkCntr[27]), .A1(n152), .Z(n44));
Q_FDP0UA U272 ( .D(n44), .QTFCLK( ), .Q(fclkCntr[27]));
Q_MX02 U273 ( .S(initClock), .A0(fclkCntr[28]), .A1(n150), .Z(n45));
Q_FDP0UA U274 ( .D(n45), .QTFCLK( ), .Q(fclkCntr[28]));
Q_MX02 U275 ( .S(initClock), .A0(fclkCntr[29]), .A1(n148), .Z(n46));
Q_FDP0UA U276 ( .D(n46), .QTFCLK( ), .Q(fclkCntr[29]));
Q_MX02 U277 ( .S(initClock), .A0(fclkCntr[30]), .A1(n146), .Z(n47));
Q_FDP0UA U278 ( .D(n47), .QTFCLK( ), .Q(fclkCntr[30]));
Q_MX02 U279 ( .S(initClock), .A0(fclkCntr[31]), .A1(n144), .Z(n48));
Q_FDP0UA U280 ( .D(n48), .QTFCLK( ), .Q(fclkCntr[31]));
Q_MX02 U281 ( .S(initClock), .A0(fclkCntr[32]), .A1(n142), .Z(n49));
Q_FDP0UA U282 ( .D(n49), .QTFCLK( ), .Q(fclkCntr[32]));
Q_MX02 U283 ( .S(initClock), .A0(fclkCntr[33]), .A1(n140), .Z(n50));
Q_FDP0UA U284 ( .D(n50), .QTFCLK( ), .Q(fclkCntr[33]));
Q_MX02 U285 ( .S(initClock), .A0(fclkCntr[34]), .A1(n138), .Z(n51));
Q_FDP0UA U286 ( .D(n51), .QTFCLK( ), .Q(fclkCntr[34]));
Q_MX02 U287 ( .S(initClock), .A0(fclkCntr[35]), .A1(n136), .Z(n52));
Q_FDP0UA U288 ( .D(n52), .QTFCLK( ), .Q(fclkCntr[35]));
Q_MX02 U289 ( .S(initClock), .A0(fclkCntr[36]), .A1(n134), .Z(n53));
Q_FDP0UA U290 ( .D(n53), .QTFCLK( ), .Q(fclkCntr[36]));
Q_MX02 U291 ( .S(initClock), .A0(fclkCntr[37]), .A1(n132), .Z(n54));
Q_FDP0UA U292 ( .D(n54), .QTFCLK( ), .Q(fclkCntr[37]));
Q_MX02 U293 ( .S(initClock), .A0(fclkCntr[38]), .A1(n130), .Z(n55));
Q_FDP0UA U294 ( .D(n55), .QTFCLK( ), .Q(fclkCntr[38]));
Q_MX02 U295 ( .S(initClock), .A0(fclkCntr[39]), .A1(n128), .Z(n56));
Q_FDP0UA U296 ( .D(n56), .QTFCLK( ), .Q(fclkCntr[39]));
Q_MX02 U297 ( .S(initClock), .A0(fclkCntr[40]), .A1(n126), .Z(n57));
Q_FDP0UA U298 ( .D(n57), .QTFCLK( ), .Q(fclkCntr[40]));
Q_MX02 U299 ( .S(initClock), .A0(fclkCntr[41]), .A1(n124), .Z(n58));
Q_FDP0UA U300 ( .D(n58), .QTFCLK( ), .Q(fclkCntr[41]));
Q_MX02 U301 ( .S(initClock), .A0(fclkCntr[42]), .A1(n122), .Z(n59));
Q_FDP0UA U302 ( .D(n59), .QTFCLK( ), .Q(fclkCntr[42]));
Q_MX02 U303 ( .S(initClock), .A0(fclkCntr[43]), .A1(n120), .Z(n60));
Q_FDP0UA U304 ( .D(n60), .QTFCLK( ), .Q(fclkCntr[43]));
Q_MX02 U305 ( .S(initClock), .A0(fclkCntr[44]), .A1(n118), .Z(n61));
Q_FDP0UA U306 ( .D(n61), .QTFCLK( ), .Q(fclkCntr[44]));
Q_MX02 U307 ( .S(initClock), .A0(fclkCntr[45]), .A1(n116), .Z(n62));
Q_FDP0UA U308 ( .D(n62), .QTFCLK( ), .Q(fclkCntr[45]));
Q_MX02 U309 ( .S(initClock), .A0(fclkCntr[46]), .A1(n114), .Z(n63));
Q_FDP0UA U310 ( .D(n63), .QTFCLK( ), .Q(fclkCntr[46]));
Q_MX02 U311 ( .S(initClock), .A0(fclkCntr[47]), .A1(n112), .Z(n64));
Q_FDP0UA U312 ( .D(n64), .QTFCLK( ), .Q(fclkCntr[47]));
Q_MX02 U313 ( .S(initClock), .A0(fclkCntr[48]), .A1(n110), .Z(n65));
Q_FDP0UA U314 ( .D(n65), .QTFCLK( ), .Q(fclkCntr[48]));
Q_MX02 U315 ( .S(initClock), .A0(fclkCntr[49]), .A1(n108), .Z(n66));
Q_FDP0UA U316 ( .D(n66), .QTFCLK( ), .Q(fclkCntr[49]));
Q_MX02 U317 ( .S(initClock), .A0(fclkCntr[50]), .A1(n106), .Z(n67));
Q_FDP0UA U318 ( .D(n67), .QTFCLK( ), .Q(fclkCntr[50]));
Q_MX02 U319 ( .S(initClock), .A0(fclkCntr[51]), .A1(n104), .Z(n68));
Q_FDP0UA U320 ( .D(n68), .QTFCLK( ), .Q(fclkCntr[51]));
Q_MX02 U321 ( .S(initClock), .A0(fclkCntr[52]), .A1(n102), .Z(n69));
Q_FDP0UA U322 ( .D(n69), .QTFCLK( ), .Q(fclkCntr[52]));
Q_MX02 U323 ( .S(initClock), .A0(fclkCntr[53]), .A1(n100), .Z(n70));
Q_FDP0UA U324 ( .D(n70), .QTFCLK( ), .Q(fclkCntr[53]));
Q_MX02 U325 ( .S(initClock), .A0(fclkCntr[54]), .A1(n98), .Z(n71));
Q_FDP0UA U326 ( .D(n71), .QTFCLK( ), .Q(fclkCntr[54]));
Q_MX02 U327 ( .S(initClock), .A0(fclkCntr[55]), .A1(n96), .Z(n72));
Q_FDP0UA U328 ( .D(n72), .QTFCLK( ), .Q(fclkCntr[55]));
Q_MX02 U329 ( .S(initClock), .A0(fclkCntr[56]), .A1(n94), .Z(n73));
Q_FDP0UA U330 ( .D(n73), .QTFCLK( ), .Q(fclkCntr[56]));
Q_MX02 U331 ( .S(initClock), .A0(fclkCntr[57]), .A1(n92), .Z(n74));
Q_FDP0UA U332 ( .D(n74), .QTFCLK( ), .Q(fclkCntr[57]));
Q_MX02 U333 ( .S(initClock), .A0(fclkCntr[58]), .A1(n90), .Z(n75));
Q_FDP0UA U334 ( .D(n75), .QTFCLK( ), .Q(fclkCntr[58]));
Q_MX02 U335 ( .S(initClock), .A0(fclkCntr[59]), .A1(n88), .Z(n76));
Q_FDP0UA U336 ( .D(n76), .QTFCLK( ), .Q(fclkCntr[59]));
Q_MX02 U337 ( .S(initClock), .A0(fclkCntr[60]), .A1(n86), .Z(n77));
Q_FDP0UA U338 ( .D(n77), .QTFCLK( ), .Q(fclkCntr[60]));
Q_MX02 U339 ( .S(initClock), .A0(fclkCntr[61]), .A1(n84), .Z(n78));
Q_FDP0UA U340 ( .D(n78), .QTFCLK( ), .Q(fclkCntr[61]));
Q_MX02 U341 ( .S(initClock), .A0(fclkCntr[62]), .A1(n82), .Z(n79));
Q_FDP0UA U342 ( .D(n79), .QTFCLK( ), .Q(fclkCntr[62]));
Q_FDP0UA U343 ( .D(n80), .QTFCLK( ), .Q(fclkCntr[63]));
Q_XOR2 U344 ( .A0(fclkCntr[63]), .A1(n15), .Z(n80));
Q_AD01HF U345 ( .A0(fclkCntr[62]), .B0(n83), .S(n82), .CO(n81));
Q_AD01HF U346 ( .A0(fclkCntr[61]), .B0(n85), .S(n84), .CO(n83));
Q_AD01HF U347 ( .A0(fclkCntr[60]), .B0(n87), .S(n86), .CO(n85));
Q_AD01HF U348 ( .A0(fclkCntr[59]), .B0(n89), .S(n88), .CO(n87));
Q_AD01HF U349 ( .A0(fclkCntr[58]), .B0(n91), .S(n90), .CO(n89));
Q_AD01HF U350 ( .A0(fclkCntr[57]), .B0(n93), .S(n92), .CO(n91));
Q_AD01HF U351 ( .A0(fclkCntr[56]), .B0(n95), .S(n94), .CO(n93));
Q_AD01HF U352 ( .A0(fclkCntr[55]), .B0(n97), .S(n96), .CO(n95));
Q_AD01HF U353 ( .A0(fclkCntr[54]), .B0(n99), .S(n98), .CO(n97));
Q_AD01HF U354 ( .A0(fclkCntr[53]), .B0(n101), .S(n100), .CO(n99));
Q_AD01HF U355 ( .A0(fclkCntr[52]), .B0(n103), .S(n102), .CO(n101));
Q_AD01HF U356 ( .A0(fclkCntr[51]), .B0(n105), .S(n104), .CO(n103));
Q_AD01HF U357 ( .A0(fclkCntr[50]), .B0(n107), .S(n106), .CO(n105));
Q_AD01HF U358 ( .A0(fclkCntr[49]), .B0(n109), .S(n108), .CO(n107));
Q_AD01HF U359 ( .A0(fclkCntr[48]), .B0(n111), .S(n110), .CO(n109));
Q_AD01HF U360 ( .A0(fclkCntr[47]), .B0(n113), .S(n112), .CO(n111));
Q_AD01HF U361 ( .A0(fclkCntr[46]), .B0(n115), .S(n114), .CO(n113));
Q_AD01HF U362 ( .A0(fclkCntr[45]), .B0(n117), .S(n116), .CO(n115));
Q_AD01HF U363 ( .A0(fclkCntr[44]), .B0(n119), .S(n118), .CO(n117));
Q_AD01HF U364 ( .A0(fclkCntr[43]), .B0(n121), .S(n120), .CO(n119));
Q_AD01HF U365 ( .A0(fclkCntr[42]), .B0(n123), .S(n122), .CO(n121));
Q_AD01HF U366 ( .A0(fclkCntr[41]), .B0(n125), .S(n124), .CO(n123));
Q_AD01HF U367 ( .A0(fclkCntr[40]), .B0(n127), .S(n126), .CO(n125));
Q_AD01HF U368 ( .A0(fclkCntr[39]), .B0(n129), .S(n128), .CO(n127));
Q_AD01HF U369 ( .A0(fclkCntr[38]), .B0(n131), .S(n130), .CO(n129));
Q_AD01HF U370 ( .A0(fclkCntr[37]), .B0(n133), .S(n132), .CO(n131));
Q_AD01HF U371 ( .A0(fclkCntr[36]), .B0(n135), .S(n134), .CO(n133));
Q_AD01HF U372 ( .A0(fclkCntr[35]), .B0(n137), .S(n136), .CO(n135));
Q_AD01HF U373 ( .A0(fclkCntr[34]), .B0(n139), .S(n138), .CO(n137));
Q_AD01HF U374 ( .A0(fclkCntr[33]), .B0(n141), .S(n140), .CO(n139));
Q_AD01HF U375 ( .A0(fclkCntr[32]), .B0(n143), .S(n142), .CO(n141));
Q_AD01HF U376 ( .A0(fclkCntr[31]), .B0(n145), .S(n144), .CO(n143));
Q_AD01HF U377 ( .A0(fclkCntr[30]), .B0(n147), .S(n146), .CO(n145));
Q_AD01HF U378 ( .A0(fclkCntr[29]), .B0(n149), .S(n148), .CO(n147));
Q_AD01HF U379 ( .A0(fclkCntr[28]), .B0(n151), .S(n150), .CO(n149));
Q_AD01HF U380 ( .A0(fclkCntr[27]), .B0(n153), .S(n152), .CO(n151));
Q_AD01HF U381 ( .A0(fclkCntr[26]), .B0(n155), .S(n154), .CO(n153));
Q_AD01HF U382 ( .A0(fclkCntr[25]), .B0(n157), .S(n156), .CO(n155));
Q_AD01HF U383 ( .A0(fclkCntr[24]), .B0(n159), .S(n158), .CO(n157));
Q_AD01HF U384 ( .A0(fclkCntr[23]), .B0(n161), .S(n160), .CO(n159));
Q_AD01HF U385 ( .A0(fclkCntr[22]), .B0(n163), .S(n162), .CO(n161));
Q_AD01HF U386 ( .A0(fclkCntr[21]), .B0(n165), .S(n164), .CO(n163));
Q_AD01HF U387 ( .A0(fclkCntr[20]), .B0(n167), .S(n166), .CO(n165));
Q_AD01HF U388 ( .A0(fclkCntr[19]), .B0(n169), .S(n168), .CO(n167));
Q_AD01HF U389 ( .A0(fclkCntr[18]), .B0(n171), .S(n170), .CO(n169));
Q_AD01HF U390 ( .A0(fclkCntr[17]), .B0(n173), .S(n172), .CO(n171));
Q_AD01HF U391 ( .A0(fclkCntr[16]), .B0(n175), .S(n174), .CO(n173));
Q_AD01HF U392 ( .A0(fclkCntr[15]), .B0(n177), .S(n176), .CO(n175));
Q_AD01HF U393 ( .A0(fclkCntr[14]), .B0(n179), .S(n178), .CO(n177));
Q_AD01HF U394 ( .A0(fclkCntr[13]), .B0(n181), .S(n180), .CO(n179));
Q_AD01HF U395 ( .A0(fclkCntr[12]), .B0(n183), .S(n182), .CO(n181));
Q_AD01HF U396 ( .A0(fclkCntr[11]), .B0(n185), .S(n184), .CO(n183));
Q_AD01HF U397 ( .A0(fclkCntr[10]), .B0(n187), .S(n186), .CO(n185));
Q_AD01HF U398 ( .A0(fclkCntr[9]), .B0(n189), .S(n188), .CO(n187));
Q_AD01HF U399 ( .A0(fclkCntr[8]), .B0(n191), .S(n190), .CO(n189));
Q_AD01HF U400 ( .A0(fclkCntr[7]), .B0(n193), .S(n192), .CO(n191));
Q_AD01HF U401 ( .A0(fclkCntr[6]), .B0(n195), .S(n194), .CO(n193));
Q_AD01HF U402 ( .A0(fclkCntr[5]), .B0(n197), .S(n196), .CO(n195));
Q_AD01HF U403 ( .A0(fclkCntr[4]), .B0(n199), .S(n198), .CO(n197));
Q_AD01HF U404 ( .A0(fclkCntr[3]), .B0(n201), .S(n200), .CO(n199));
Q_AD01HF U405 ( .A0(fclkCntr[2]), .B0(n203), .S(n202), .CO(n201));
Q_AD01HF U406 ( .A0(fclkCntr[1]), .B0(fclkCntr[0]), .S(n204), .CO(n203));
Q_NR02 U407 ( .A0(n301), .A1(n205), .Z(n16));
Q_AN02 U408 ( .A0(n207), .A1(n206), .Z(n205));
Q_AN03 U409 ( .A0(n210), .A1(n209), .A2(n208), .Z(n206));
Q_AN03 U410 ( .A0(n213), .A1(n212), .A2(n211), .Z(n207));
Q_AN03 U411 ( .A0(n216), .A1(n215), .A2(n214), .Z(n208));
Q_AN03 U412 ( .A0(n219), .A1(n218), .A2(n217), .Z(n209));
Q_AN03 U413 ( .A0(n222), .A1(n221), .A2(n220), .Z(n210));
Q_AN03 U414 ( .A0(n225), .A1(n224), .A2(n223), .Z(n211));
Q_AN03 U415 ( .A0(n228), .A1(n227), .A2(n226), .Z(n212));
Q_AN03 U416 ( .A0(n231), .A1(n230), .A2(n229), .Z(n213));
Q_AN03 U417 ( .A0(n234), .A1(n233), .A2(n232), .Z(n214));
Q_AN03 U418 ( .A0(n300), .A1(n236), .A2(n235), .Z(n215));
Q_AN03 U419 ( .A0(n297), .A1(n298), .A2(n299), .Z(n216));
Q_AN03 U420 ( .A0(n294), .A1(n295), .A2(n296), .Z(n217));
Q_AN03 U421 ( .A0(n291), .A1(n292), .A2(n293), .Z(n218));
Q_AN03 U422 ( .A0(n288), .A1(n289), .A2(n290), .Z(n219));
Q_AN03 U423 ( .A0(n285), .A1(n286), .A2(n287), .Z(n220));
Q_AN03 U424 ( .A0(n282), .A1(n283), .A2(n284), .Z(n221));
Q_AN03 U425 ( .A0(n279), .A1(n280), .A2(n281), .Z(n222));
Q_AN03 U426 ( .A0(n276), .A1(n277), .A2(n278), .Z(n223));
Q_AN03 U427 ( .A0(n273), .A1(n274), .A2(n275), .Z(n224));
Q_AN03 U428 ( .A0(n270), .A1(n271), .A2(n272), .Z(n225));
Q_AN03 U429 ( .A0(n267), .A1(n268), .A2(n269), .Z(n226));
Q_AN03 U430 ( .A0(n264), .A1(n265), .A2(n266), .Z(n227));
Q_AN03 U431 ( .A0(n261), .A1(n262), .A2(n263), .Z(n228));
Q_AN03 U432 ( .A0(n258), .A1(n259), .A2(n260), .Z(n229));
Q_AN03 U433 ( .A0(n255), .A1(n256), .A2(n257), .Z(n230));
Q_AN03 U434 ( .A0(n252), .A1(n253), .A2(n254), .Z(n231));
Q_AN03 U435 ( .A0(n249), .A1(n250), .A2(n251), .Z(n232));
Q_AN03 U436 ( .A0(n246), .A1(n247), .A2(n248), .Z(n233));
Q_AN03 U437 ( .A0(n243), .A1(n244), .A2(n245), .Z(n234));
Q_AN03 U438 ( .A0(n240), .A1(n241), .A2(n242), .Z(n235));
Q_AN03 U439 ( .A0(n237), .A1(n238), .A2(n239), .Z(n236));
Q_XNR2 U440 ( .A0(fclkCntr[63]), .A1(uClkCntr[63]), .Z(n237));
Q_XNR2 U441 ( .A0(fclkCntr[62]), .A1(uClkCntr[62]), .Z(n238));
Q_XNR2 U442 ( .A0(fclkCntr[61]), .A1(uClkCntr[61]), .Z(n239));
Q_XNR2 U443 ( .A0(fclkCntr[60]), .A1(uClkCntr[60]), .Z(n240));
Q_XNR2 U444 ( .A0(fclkCntr[59]), .A1(uClkCntr[59]), .Z(n241));
Q_XNR2 U445 ( .A0(fclkCntr[58]), .A1(uClkCntr[58]), .Z(n242));
Q_XNR2 U446 ( .A0(fclkCntr[57]), .A1(uClkCntr[57]), .Z(n243));
Q_XNR2 U447 ( .A0(fclkCntr[56]), .A1(uClkCntr[56]), .Z(n244));
Q_XNR2 U448 ( .A0(fclkCntr[55]), .A1(uClkCntr[55]), .Z(n245));
Q_XNR2 U449 ( .A0(fclkCntr[54]), .A1(uClkCntr[54]), .Z(n246));
Q_XNR2 U450 ( .A0(fclkCntr[53]), .A1(uClkCntr[53]), .Z(n247));
Q_XNR2 U451 ( .A0(fclkCntr[52]), .A1(uClkCntr[52]), .Z(n248));
Q_XNR2 U452 ( .A0(fclkCntr[51]), .A1(uClkCntr[51]), .Z(n249));
Q_XNR2 U453 ( .A0(fclkCntr[50]), .A1(uClkCntr[50]), .Z(n250));
Q_XNR2 U454 ( .A0(fclkCntr[49]), .A1(uClkCntr[49]), .Z(n251));
Q_XNR2 U455 ( .A0(fclkCntr[48]), .A1(uClkCntr[48]), .Z(n252));
Q_XNR2 U456 ( .A0(fclkCntr[47]), .A1(uClkCntr[47]), .Z(n253));
Q_XNR2 U457 ( .A0(fclkCntr[46]), .A1(uClkCntr[46]), .Z(n254));
Q_XNR2 U458 ( .A0(fclkCntr[45]), .A1(uClkCntr[45]), .Z(n255));
Q_XNR2 U459 ( .A0(fclkCntr[44]), .A1(uClkCntr[44]), .Z(n256));
Q_XNR2 U460 ( .A0(fclkCntr[43]), .A1(uClkCntr[43]), .Z(n257));
Q_XNR2 U461 ( .A0(fclkCntr[42]), .A1(uClkCntr[42]), .Z(n258));
Q_XNR2 U462 ( .A0(fclkCntr[41]), .A1(uClkCntr[41]), .Z(n259));
Q_XNR2 U463 ( .A0(fclkCntr[40]), .A1(uClkCntr[40]), .Z(n260));
Q_XNR2 U464 ( .A0(fclkCntr[39]), .A1(uClkCntr[39]), .Z(n261));
Q_XNR2 U465 ( .A0(fclkCntr[38]), .A1(uClkCntr[38]), .Z(n262));
Q_XNR2 U466 ( .A0(fclkCntr[37]), .A1(uClkCntr[37]), .Z(n263));
Q_XNR2 U467 ( .A0(fclkCntr[36]), .A1(uClkCntr[36]), .Z(n264));
Q_XNR2 U468 ( .A0(fclkCntr[35]), .A1(uClkCntr[35]), .Z(n265));
Q_XNR2 U469 ( .A0(fclkCntr[34]), .A1(uClkCntr[34]), .Z(n266));
Q_XNR2 U470 ( .A0(fclkCntr[33]), .A1(uClkCntr[33]), .Z(n267));
Q_XNR2 U471 ( .A0(fclkCntr[32]), .A1(uClkCntr[32]), .Z(n268));
Q_XNR2 U472 ( .A0(fclkCntr[31]), .A1(uClkCntr[31]), .Z(n269));
Q_XNR2 U473 ( .A0(fclkCntr[30]), .A1(uClkCntr[30]), .Z(n270));
Q_XNR2 U474 ( .A0(fclkCntr[29]), .A1(uClkCntr[29]), .Z(n271));
Q_XNR2 U475 ( .A0(fclkCntr[28]), .A1(uClkCntr[28]), .Z(n272));
Q_XNR2 U476 ( .A0(fclkCntr[27]), .A1(uClkCntr[27]), .Z(n273));
Q_XNR2 U477 ( .A0(fclkCntr[26]), .A1(uClkCntr[26]), .Z(n274));
Q_XNR2 U478 ( .A0(fclkCntr[25]), .A1(uClkCntr[25]), .Z(n275));
Q_XNR2 U479 ( .A0(fclkCntr[24]), .A1(uClkCntr[24]), .Z(n276));
Q_XNR2 U480 ( .A0(fclkCntr[23]), .A1(uClkCntr[23]), .Z(n277));
Q_XNR2 U481 ( .A0(fclkCntr[22]), .A1(uClkCntr[22]), .Z(n278));
Q_XNR2 U482 ( .A0(fclkCntr[21]), .A1(uClkCntr[21]), .Z(n279));
Q_XNR2 U483 ( .A0(fclkCntr[20]), .A1(uClkCntr[20]), .Z(n280));
Q_XNR2 U484 ( .A0(fclkCntr[19]), .A1(uClkCntr[19]), .Z(n281));
Q_XNR2 U485 ( .A0(fclkCntr[18]), .A1(uClkCntr[18]), .Z(n282));
Q_XNR2 U486 ( .A0(fclkCntr[17]), .A1(uClkCntr[17]), .Z(n283));
Q_XNR2 U487 ( .A0(fclkCntr[16]), .A1(uClkCntr[16]), .Z(n284));
Q_XNR2 U488 ( .A0(fclkCntr[15]), .A1(uClkCntr[15]), .Z(n285));
Q_XNR2 U489 ( .A0(fclkCntr[14]), .A1(uClkCntr[14]), .Z(n286));
Q_XNR2 U490 ( .A0(fclkCntr[13]), .A1(uClkCntr[13]), .Z(n287));
Q_XNR2 U491 ( .A0(fclkCntr[12]), .A1(uClkCntr[12]), .Z(n288));
Q_XNR2 U492 ( .A0(fclkCntr[11]), .A1(uClkCntr[11]), .Z(n289));
Q_XNR2 U493 ( .A0(fclkCntr[10]), .A1(uClkCntr[10]), .Z(n290));
Q_XNR2 U494 ( .A0(fclkCntr[9]), .A1(uClkCntr[9]), .Z(n291));
Q_XNR2 U495 ( .A0(fclkCntr[8]), .A1(uClkCntr[8]), .Z(n292));
Q_XNR2 U496 ( .A0(fclkCntr[7]), .A1(uClkCntr[7]), .Z(n293));
Q_XNR2 U497 ( .A0(fclkCntr[6]), .A1(uClkCntr[6]), .Z(n294));
Q_XNR2 U498 ( .A0(fclkCntr[5]), .A1(uClkCntr[5]), .Z(n295));
Q_XNR2 U499 ( .A0(fclkCntr[4]), .A1(uClkCntr[4]), .Z(n296));
Q_XNR2 U500 ( .A0(fclkCntr[3]), .A1(uClkCntr[3]), .Z(n297));
Q_XNR2 U501 ( .A0(fclkCntr[2]), .A1(uClkCntr[2]), .Z(n298));
Q_XNR2 U502 ( .A0(fclkCntr[1]), .A1(uClkCntr[1]), .Z(n299));
Q_XNR2 U503 ( .A0(fclkCntr[0]), .A1(uClkCntr[0]), .Z(n300));
Q_OR02 U504 ( .A0(n303), .A1(n302), .Z(n301));
Q_OR03 U505 ( .A0(n306), .A1(n305), .A2(n304), .Z(n302));
Q_OR03 U506 ( .A0(n309), .A1(n308), .A2(n307), .Z(n303));
Q_OR03 U507 ( .A0(n312), .A1(n311), .A2(n310), .Z(n304));
Q_OR03 U508 ( .A0(n315), .A1(n314), .A2(n313), .Z(n305));
Q_OR03 U509 ( .A0(n318), .A1(n317), .A2(n316), .Z(n306));
Q_OR03 U510 ( .A0(n321), .A1(n320), .A2(n319), .Z(n307));
Q_OR03 U511 ( .A0(n324), .A1(n323), .A2(n322), .Z(n308));
Q_OR03 U512 ( .A0(n327), .A1(n326), .A2(n325), .Z(n309));
Q_OR03 U513 ( .A0(n330), .A1(n329), .A2(n328), .Z(n310));
Q_OR03 U514 ( .A0(uClkErrTime[0]), .A1(n332), .A2(n331), .Z(n311));
Q_OR03 U515 ( .A0(uClkErrTime[3]), .A1(uClkErrTime[2]), .A2(uClkErrTime[1]), .Z(n312));
Q_OR03 U516 ( .A0(uClkErrTime[6]), .A1(uClkErrTime[5]), .A2(uClkErrTime[4]), .Z(n313));
Q_OR03 U517 ( .A0(uClkErrTime[9]), .A1(uClkErrTime[8]), .A2(uClkErrTime[7]), .Z(n314));
Q_OR03 U518 ( .A0(uClkErrTime[12]), .A1(uClkErrTime[11]), .A2(uClkErrTime[10]), .Z(n315));
Q_OR03 U519 ( .A0(uClkErrTime[15]), .A1(uClkErrTime[14]), .A2(uClkErrTime[13]), .Z(n316));
Q_OR03 U520 ( .A0(uClkErrTime[18]), .A1(uClkErrTime[17]), .A2(uClkErrTime[16]), .Z(n317));
Q_OR03 U521 ( .A0(uClkErrTime[21]), .A1(uClkErrTime[20]), .A2(uClkErrTime[19]), .Z(n318));
Q_OR03 U522 ( .A0(uClkErrTime[24]), .A1(uClkErrTime[23]), .A2(uClkErrTime[22]), .Z(n319));
Q_OR03 U523 ( .A0(uClkErrTime[27]), .A1(uClkErrTime[26]), .A2(uClkErrTime[25]), .Z(n320));
Q_OR03 U524 ( .A0(uClkErrTime[30]), .A1(uClkErrTime[29]), .A2(uClkErrTime[28]), .Z(n321));
Q_OR03 U525 ( .A0(uClkErrTime[33]), .A1(uClkErrTime[32]), .A2(uClkErrTime[31]), .Z(n322));
Q_OR03 U526 ( .A0(uClkErrTime[36]), .A1(uClkErrTime[35]), .A2(uClkErrTime[34]), .Z(n323));
Q_OR03 U527 ( .A0(uClkErrTime[39]), .A1(uClkErrTime[38]), .A2(uClkErrTime[37]), .Z(n324));
Q_OR03 U528 ( .A0(uClkErrTime[42]), .A1(uClkErrTime[41]), .A2(uClkErrTime[40]), .Z(n325));
Q_OR03 U529 ( .A0(uClkErrTime[45]), .A1(uClkErrTime[44]), .A2(uClkErrTime[43]), .Z(n326));
Q_OR03 U530 ( .A0(uClkErrTime[48]), .A1(uClkErrTime[47]), .A2(uClkErrTime[46]), .Z(n327));
Q_OR03 U531 ( .A0(uClkErrTime[51]), .A1(uClkErrTime[50]), .A2(uClkErrTime[49]), .Z(n328));
Q_OR03 U532 ( .A0(uClkErrTime[54]), .A1(uClkErrTime[53]), .A2(uClkErrTime[52]), .Z(n329));
Q_OR03 U533 ( .A0(uClkErrTime[57]), .A1(uClkErrTime[56]), .A2(uClkErrTime[55]), .Z(n330));
Q_OR03 U534 ( .A0(uClkErrTime[60]), .A1(uClkErrTime[59]), .A2(uClkErrTime[58]), .Z(n331));
Q_OR03 U535 ( .A0(uClkErrTime[63]), .A1(uClkErrTime[62]), .A2(uClkErrTime[61]), .Z(n332));
Q_MX02 U536 ( .S(n16), .A0(uClkErrTime[0]), .A1(simTime[0]), .Z(n333));
Q_FDP0UA U537 ( .D(n333), .QTFCLK( ), .Q(uClkErrTime[0]));
Q_MX02 U538 ( .S(n16), .A0(uClkErrTime[1]), .A1(simTime[1]), .Z(n334));
Q_FDP0UA U539 ( .D(n334), .QTFCLK( ), .Q(uClkErrTime[1]));
Q_MX02 U540 ( .S(n16), .A0(uClkErrTime[2]), .A1(simTime[2]), .Z(n335));
Q_FDP0UA U541 ( .D(n335), .QTFCLK( ), .Q(uClkErrTime[2]));
Q_MX02 U542 ( .S(n16), .A0(uClkErrTime[3]), .A1(simTime[3]), .Z(n336));
Q_FDP0UA U543 ( .D(n336), .QTFCLK( ), .Q(uClkErrTime[3]));
Q_MX02 U544 ( .S(n16), .A0(uClkErrTime[4]), .A1(simTime[4]), .Z(n337));
Q_FDP0UA U545 ( .D(n337), .QTFCLK( ), .Q(uClkErrTime[4]));
Q_MX02 U546 ( .S(n16), .A0(uClkErrTime[5]), .A1(simTime[5]), .Z(n338));
Q_FDP0UA U547 ( .D(n338), .QTFCLK( ), .Q(uClkErrTime[5]));
Q_MX02 U548 ( .S(n16), .A0(uClkErrTime[6]), .A1(simTime[6]), .Z(n339));
Q_FDP0UA U549 ( .D(n339), .QTFCLK( ), .Q(uClkErrTime[6]));
Q_MX02 U550 ( .S(n16), .A0(uClkErrTime[7]), .A1(simTime[7]), .Z(n340));
Q_FDP0UA U551 ( .D(n340), .QTFCLK( ), .Q(uClkErrTime[7]));
Q_MX02 U552 ( .S(n16), .A0(uClkErrTime[8]), .A1(simTime[8]), .Z(n341));
Q_FDP0UA U553 ( .D(n341), .QTFCLK( ), .Q(uClkErrTime[8]));
Q_MX02 U554 ( .S(n16), .A0(uClkErrTime[9]), .A1(simTime[9]), .Z(n342));
Q_FDP0UA U555 ( .D(n342), .QTFCLK( ), .Q(uClkErrTime[9]));
Q_MX02 U556 ( .S(n16), .A0(uClkErrTime[10]), .A1(simTime[10]), .Z(n343));
Q_FDP0UA U557 ( .D(n343), .QTFCLK( ), .Q(uClkErrTime[10]));
Q_MX02 U558 ( .S(n16), .A0(uClkErrTime[11]), .A1(simTime[11]), .Z(n344));
Q_FDP0UA U559 ( .D(n344), .QTFCLK( ), .Q(uClkErrTime[11]));
Q_MX02 U560 ( .S(n16), .A0(uClkErrTime[12]), .A1(simTime[12]), .Z(n345));
Q_FDP0UA U561 ( .D(n345), .QTFCLK( ), .Q(uClkErrTime[12]));
Q_MX02 U562 ( .S(n16), .A0(uClkErrTime[13]), .A1(simTime[13]), .Z(n346));
Q_FDP0UA U563 ( .D(n346), .QTFCLK( ), .Q(uClkErrTime[13]));
Q_MX02 U564 ( .S(n16), .A0(uClkErrTime[14]), .A1(simTime[14]), .Z(n347));
Q_FDP0UA U565 ( .D(n347), .QTFCLK( ), .Q(uClkErrTime[14]));
Q_MX02 U566 ( .S(n16), .A0(uClkErrTime[15]), .A1(simTime[15]), .Z(n348));
Q_FDP0UA U567 ( .D(n348), .QTFCLK( ), .Q(uClkErrTime[15]));
Q_MX02 U568 ( .S(n16), .A0(uClkErrTime[16]), .A1(simTime[16]), .Z(n349));
Q_FDP0UA U569 ( .D(n349), .QTFCLK( ), .Q(uClkErrTime[16]));
Q_MX02 U570 ( .S(n16), .A0(uClkErrTime[17]), .A1(simTime[17]), .Z(n350));
Q_FDP0UA U571 ( .D(n350), .QTFCLK( ), .Q(uClkErrTime[17]));
Q_MX02 U572 ( .S(n16), .A0(uClkErrTime[18]), .A1(simTime[18]), .Z(n351));
Q_FDP0UA U573 ( .D(n351), .QTFCLK( ), .Q(uClkErrTime[18]));
Q_MX02 U574 ( .S(n16), .A0(uClkErrTime[19]), .A1(simTime[19]), .Z(n352));
Q_FDP0UA U575 ( .D(n352), .QTFCLK( ), .Q(uClkErrTime[19]));
Q_MX02 U576 ( .S(n16), .A0(uClkErrTime[20]), .A1(simTime[20]), .Z(n353));
Q_FDP0UA U577 ( .D(n353), .QTFCLK( ), .Q(uClkErrTime[20]));
Q_MX02 U578 ( .S(n16), .A0(uClkErrTime[21]), .A1(simTime[21]), .Z(n354));
Q_FDP0UA U579 ( .D(n354), .QTFCLK( ), .Q(uClkErrTime[21]));
Q_MX02 U580 ( .S(n16), .A0(uClkErrTime[22]), .A1(simTime[22]), .Z(n355));
Q_FDP0UA U581 ( .D(n355), .QTFCLK( ), .Q(uClkErrTime[22]));
Q_MX02 U582 ( .S(n16), .A0(uClkErrTime[23]), .A1(simTime[23]), .Z(n356));
Q_FDP0UA U583 ( .D(n356), .QTFCLK( ), .Q(uClkErrTime[23]));
Q_MX02 U584 ( .S(n16), .A0(uClkErrTime[24]), .A1(simTime[24]), .Z(n357));
Q_FDP0UA U585 ( .D(n357), .QTFCLK( ), .Q(uClkErrTime[24]));
Q_MX02 U586 ( .S(n16), .A0(uClkErrTime[25]), .A1(simTime[25]), .Z(n358));
Q_FDP0UA U587 ( .D(n358), .QTFCLK( ), .Q(uClkErrTime[25]));
Q_MX02 U588 ( .S(n16), .A0(uClkErrTime[26]), .A1(simTime[26]), .Z(n359));
Q_FDP0UA U589 ( .D(n359), .QTFCLK( ), .Q(uClkErrTime[26]));
Q_MX02 U590 ( .S(n16), .A0(uClkErrTime[27]), .A1(simTime[27]), .Z(n360));
Q_FDP0UA U591 ( .D(n360), .QTFCLK( ), .Q(uClkErrTime[27]));
Q_MX02 U592 ( .S(n16), .A0(uClkErrTime[28]), .A1(simTime[28]), .Z(n361));
Q_FDP0UA U593 ( .D(n361), .QTFCLK( ), .Q(uClkErrTime[28]));
Q_MX02 U594 ( .S(n16), .A0(uClkErrTime[29]), .A1(simTime[29]), .Z(n362));
Q_FDP0UA U595 ( .D(n362), .QTFCLK( ), .Q(uClkErrTime[29]));
Q_MX02 U596 ( .S(n16), .A0(uClkErrTime[30]), .A1(simTime[30]), .Z(n363));
Q_FDP0UA U597 ( .D(n363), .QTFCLK( ), .Q(uClkErrTime[30]));
Q_MX02 U598 ( .S(n16), .A0(uClkErrTime[31]), .A1(simTime[31]), .Z(n364));
Q_FDP0UA U599 ( .D(n364), .QTFCLK( ), .Q(uClkErrTime[31]));
Q_MX02 U600 ( .S(n16), .A0(uClkErrTime[32]), .A1(simTime[32]), .Z(n365));
Q_FDP0UA U601 ( .D(n365), .QTFCLK( ), .Q(uClkErrTime[32]));
Q_MX02 U602 ( .S(n16), .A0(uClkErrTime[33]), .A1(simTime[33]), .Z(n366));
Q_FDP0UA U603 ( .D(n366), .QTFCLK( ), .Q(uClkErrTime[33]));
Q_MX02 U604 ( .S(n16), .A0(uClkErrTime[34]), .A1(simTime[34]), .Z(n367));
Q_FDP0UA U605 ( .D(n367), .QTFCLK( ), .Q(uClkErrTime[34]));
Q_MX02 U606 ( .S(n16), .A0(uClkErrTime[35]), .A1(simTime[35]), .Z(n368));
Q_FDP0UA U607 ( .D(n368), .QTFCLK( ), .Q(uClkErrTime[35]));
Q_MX02 U608 ( .S(n16), .A0(uClkErrTime[36]), .A1(simTime[36]), .Z(n369));
Q_FDP0UA U609 ( .D(n369), .QTFCLK( ), .Q(uClkErrTime[36]));
Q_MX02 U610 ( .S(n16), .A0(uClkErrTime[37]), .A1(simTime[37]), .Z(n370));
Q_FDP0UA U611 ( .D(n370), .QTFCLK( ), .Q(uClkErrTime[37]));
Q_MX02 U612 ( .S(n16), .A0(uClkErrTime[38]), .A1(simTime[38]), .Z(n371));
Q_FDP0UA U613 ( .D(n371), .QTFCLK( ), .Q(uClkErrTime[38]));
Q_MX02 U614 ( .S(n16), .A0(uClkErrTime[39]), .A1(simTime[39]), .Z(n372));
Q_FDP0UA U615 ( .D(n372), .QTFCLK( ), .Q(uClkErrTime[39]));
Q_MX02 U616 ( .S(n16), .A0(uClkErrTime[40]), .A1(simTime[40]), .Z(n373));
Q_FDP0UA U617 ( .D(n373), .QTFCLK( ), .Q(uClkErrTime[40]));
Q_MX02 U618 ( .S(n16), .A0(uClkErrTime[41]), .A1(simTime[41]), .Z(n374));
Q_FDP0UA U619 ( .D(n374), .QTFCLK( ), .Q(uClkErrTime[41]));
Q_MX02 U620 ( .S(n16), .A0(uClkErrTime[42]), .A1(simTime[42]), .Z(n375));
Q_FDP0UA U621 ( .D(n375), .QTFCLK( ), .Q(uClkErrTime[42]));
Q_MX02 U622 ( .S(n16), .A0(uClkErrTime[43]), .A1(simTime[43]), .Z(n376));
Q_FDP0UA U623 ( .D(n376), .QTFCLK( ), .Q(uClkErrTime[43]));
Q_MX02 U624 ( .S(n16), .A0(uClkErrTime[44]), .A1(simTime[44]), .Z(n377));
Q_FDP0UA U625 ( .D(n377), .QTFCLK( ), .Q(uClkErrTime[44]));
Q_MX02 U626 ( .S(n16), .A0(uClkErrTime[45]), .A1(simTime[45]), .Z(n378));
Q_FDP0UA U627 ( .D(n378), .QTFCLK( ), .Q(uClkErrTime[45]));
Q_MX02 U628 ( .S(n16), .A0(uClkErrTime[46]), .A1(simTime[46]), .Z(n379));
Q_FDP0UA U629 ( .D(n379), .QTFCLK( ), .Q(uClkErrTime[46]));
Q_MX02 U630 ( .S(n16), .A0(uClkErrTime[47]), .A1(simTime[47]), .Z(n380));
Q_FDP0UA U631 ( .D(n380), .QTFCLK( ), .Q(uClkErrTime[47]));
Q_MX02 U632 ( .S(n16), .A0(uClkErrTime[48]), .A1(simTime[48]), .Z(n381));
Q_FDP0UA U633 ( .D(n381), .QTFCLK( ), .Q(uClkErrTime[48]));
Q_MX02 U634 ( .S(n16), .A0(uClkErrTime[49]), .A1(simTime[49]), .Z(n382));
Q_FDP0UA U635 ( .D(n382), .QTFCLK( ), .Q(uClkErrTime[49]));
Q_MX02 U636 ( .S(n16), .A0(uClkErrTime[50]), .A1(simTime[50]), .Z(n383));
Q_FDP0UA U637 ( .D(n383), .QTFCLK( ), .Q(uClkErrTime[50]));
Q_MX02 U638 ( .S(n16), .A0(uClkErrTime[51]), .A1(simTime[51]), .Z(n384));
Q_FDP0UA U639 ( .D(n384), .QTFCLK( ), .Q(uClkErrTime[51]));
Q_MX02 U640 ( .S(n16), .A0(uClkErrTime[52]), .A1(simTime[52]), .Z(n385));
Q_FDP0UA U641 ( .D(n385), .QTFCLK( ), .Q(uClkErrTime[52]));
Q_MX02 U642 ( .S(n16), .A0(uClkErrTime[53]), .A1(simTime[53]), .Z(n386));
Q_FDP0UA U643 ( .D(n386), .QTFCLK( ), .Q(uClkErrTime[53]));
Q_MX02 U644 ( .S(n16), .A0(uClkErrTime[54]), .A1(simTime[54]), .Z(n387));
Q_FDP0UA U645 ( .D(n387), .QTFCLK( ), .Q(uClkErrTime[54]));
Q_MX02 U646 ( .S(n16), .A0(uClkErrTime[55]), .A1(simTime[55]), .Z(n388));
Q_FDP0UA U647 ( .D(n388), .QTFCLK( ), .Q(uClkErrTime[55]));
Q_MX02 U648 ( .S(n16), .A0(uClkErrTime[56]), .A1(simTime[56]), .Z(n389));
Q_FDP0UA U649 ( .D(n389), .QTFCLK( ), .Q(uClkErrTime[56]));
Q_MX02 U650 ( .S(n16), .A0(uClkErrTime[57]), .A1(simTime[57]), .Z(n390));
Q_FDP0UA U651 ( .D(n390), .QTFCLK( ), .Q(uClkErrTime[57]));
Q_MX02 U652 ( .S(n16), .A0(uClkErrTime[58]), .A1(simTime[58]), .Z(n391));
Q_FDP0UA U653 ( .D(n391), .QTFCLK( ), .Q(uClkErrTime[58]));
Q_MX02 U654 ( .S(n16), .A0(uClkErrTime[59]), .A1(simTime[59]), .Z(n392));
Q_FDP0UA U655 ( .D(n392), .QTFCLK( ), .Q(uClkErrTime[59]));
Q_MX02 U656 ( .S(n16), .A0(uClkErrTime[60]), .A1(simTime[60]), .Z(n393));
Q_FDP0UA U657 ( .D(n393), .QTFCLK( ), .Q(uClkErrTime[60]));
Q_MX02 U658 ( .S(n16), .A0(uClkErrTime[61]), .A1(simTime[61]), .Z(n394));
Q_FDP0UA U659 ( .D(n394), .QTFCLK( ), .Q(uClkErrTime[61]));
Q_MX02 U660 ( .S(n16), .A0(uClkErrTime[62]), .A1(simTime[62]), .Z(n395));
Q_FDP0UA U661 ( .D(n395), .QTFCLK( ), .Q(uClkErrTime[62]));
Q_MX02 U662 ( .S(n16), .A0(uClkErrTime[63]), .A1(simTime[63]), .Z(n396));
Q_FDP0UA U663 ( .D(n396), .QTFCLK( ), .Q(uClkErrTime[63]));
Q_OR02 U664 ( .A0(bpWait), .A1(xpHold), .Z(n401));
Q_AO21 U665 ( .A0(n457), .A1(n401), .B0(lbrOn), .Z(n402));
Q_AO21 U666 ( .A0(n402), .A1(dccState), .B0(n403), .Z(n404));
Q_INV U667 ( .A(n407), .Z(n403));
Q_INV U668 ( .A(n398), .Z(n405));
Q_OR02 U669 ( .A0(n405), .A1(n404), .Z(n406));
Q_OR02 U670 ( .A0(dccState), .A1(lbrOn), .Z(n407));
Q_AN02 U671 ( .A0(n398), .A1(n407), .Z(n399));
Q_INV U672 ( .A(n397), .Z(n400));
Q_MX02 U673 ( .S(n406), .A0(lbrOn), .A1(dccState), .Z(n408));
Q_FDP0UA U674 ( .D(n408), .QTFCLK( ), .Q(dccState));
Q_MX02 U675 ( .S(n399), .A0(dccFrameFill[0]), .A1(n425), .Z(n409));
Q_FDP0UA U676 ( .D(n409), .QTFCLK( ), .Q(dccFrameFill[0]));
Q_MX02 U677 ( .S(n399), .A0(dccFrameFill[1]), .A1(n424), .Z(n410));
Q_FDP0UA U678 ( .D(n410), .QTFCLK( ), .Q(dccFrameFill[1]));
Q_MX02 U679 ( .S(n399), .A0(dccFrameFill[2]), .A1(n423), .Z(n411));
Q_FDP0UA U680 ( .D(n411), .QTFCLK( ), .Q(dccFrameFill[2]));
Q_MX02 U681 ( .S(n399), .A0(dccFrameFill[3]), .A1(n422), .Z(n412));
Q_FDP0UA U682 ( .D(n412), .QTFCLK( ), .Q(dccFrameFill[3]));
Q_MX02 U683 ( .S(n399), .A0(dccFrameFill[4]), .A1(n421), .Z(n413));
Q_FDP0UA U684 ( .D(n413), .QTFCLK( ), .Q(dccFrameFill[4]));
Q_MX02 U685 ( .S(n399), .A0(dccFrameFill[5]), .A1(n420), .Z(n414));
Q_FDP0UA U686 ( .D(n414), .QTFCLK( ), .Q(dccFrameFill[5]));
Q_MX02 U687 ( .S(n399), .A0(dccFrameFill[6]), .A1(n419), .Z(n415));
Q_FDP0UA U688 ( .D(n415), .QTFCLK( ), .Q(dccFrameFill[6]));
Q_MX02 U689 ( .S(n399), .A0(dccFrameFill[7]), .A1(n418), .Z(n416));
Q_FDP0UA U690 ( .D(n416), .QTFCLK( ), .Q(dccFrameFill[7]));
Q_MX02 U691 ( .S(n398), .A0(bWaitExtend), .A1(n427), .Z(n417));
Q_FDP0UA U692 ( .D(n417), .QTFCLK( ), .Q(bWaitExtend));
Q_AN02 U693 ( .A0(dccState), .A1(n461), .Z(n418));
Q_AN02 U694 ( .A0(dccState), .A1(n462), .Z(n419));
Q_AN02 U695 ( .A0(dccState), .A1(n463), .Z(n420));
Q_AN02 U696 ( .A0(dccState), .A1(n464), .Z(n421));
Q_AN02 U697 ( .A0(dccState), .A1(n465), .Z(n422));
Q_AN02 U698 ( .A0(dccState), .A1(n466), .Z(n423));
Q_AN02 U699 ( .A0(dccState), .A1(n467), .Z(n424));
Q_OR02 U700 ( .A0(n426), .A1(n468), .Z(n425));
Q_INV U701 ( .A(dccState), .Z(n426));
Q_AN03 U702 ( .A0(n401), .A1(n428), .A2(dccState), .Z(n427));
Q_AO21 U703 ( .A0(n443), .A1(n429), .B0(n444), .Z(n428));
Q_OR03 U704 ( .A0(n441), .A1(n430), .A2(n431), .Z(n429));
Q_AO21 U705 ( .A0(n433), .A1(n437), .B0(n432), .Z(n431));
Q_AN03 U706 ( .A0(n433), .A1(n436), .A2(n434), .Z(n432));
Q_AN02 U707 ( .A0(n468), .A1(n435), .Z(n434));
Q_INV U708 ( .A(DccFrameMark[0]), .Z(n435));
Q_OR02 U709 ( .A0(n467), .A1(n438), .Z(n436));
Q_AN02 U710 ( .A0(n467), .A1(n438), .Z(n437));
Q_INV U711 ( .A(DccFrameMark[1]), .Z(n438));
Q_OA21 U712 ( .A0(n466), .A1(n439), .B0(n440), .Z(n433));
Q_AN03 U713 ( .A0(n466), .A1(n439), .A2(n440), .Z(n430));
Q_INV U714 ( .A(DccFrameMark[2]), .Z(n439));
Q_OR02 U715 ( .A0(n465), .A1(n442), .Z(n440));
Q_AN02 U716 ( .A0(n465), .A1(n442), .Z(n441));
Q_INV U717 ( .A(DccFrameMark[3]), .Z(n442));
Q_OR03 U718 ( .A0(n455), .A1(n445), .A2(n446), .Z(n444));
Q_AO21 U719 ( .A0(n449), .A1(n451), .B0(n447), .Z(n446));
Q_OA21 U720 ( .A0(n464), .A1(n450), .B0(n448), .Z(n443));
Q_AN03 U721 ( .A0(n464), .A1(n450), .A2(n448), .Z(n447));
Q_INV U722 ( .A(DccFrameMark[4]), .Z(n450));
Q_OA21 U723 ( .A0(n463), .A1(n452), .B0(n449), .Z(n448));
Q_AN02 U724 ( .A0(n463), .A1(n452), .Z(n451));
Q_INV U725 ( .A(DccFrameMark[5]), .Z(n452));
Q_OA21 U726 ( .A0(n462), .A1(n453), .B0(n454), .Z(n449));
Q_AN03 U727 ( .A0(n462), .A1(n453), .A2(n454), .Z(n445));
Q_INV U728 ( .A(DccFrameMark[6]), .Z(n453));
Q_OR02 U729 ( .A0(n461), .A1(n456), .Z(n454));
Q_AN02 U730 ( .A0(n461), .A1(n456), .Z(n455));
Q_INV U731 ( .A(DccFrameMark[7]), .Z(n456));
Q_OR02 U732 ( .A0(n459), .A1(n458), .Z(n457));
Q_OR03 U733 ( .A0(n462), .A1(n461), .A2(n460), .Z(n458));
Q_OR03 U734 ( .A0(n465), .A1(n464), .A2(n463), .Z(n459));
Q_OR03 U735 ( .A0(n468), .A1(n467), .A2(n466), .Z(n460));
Q_AN02 U736 ( .A0(n400), .A1(n480), .Z(n461));
Q_AN02 U737 ( .A0(n400), .A1(n482), .Z(n462));
Q_AN02 U738 ( .A0(n400), .A1(n484), .Z(n463));
Q_AN02 U739 ( .A0(n400), .A1(n486), .Z(n464));
Q_AN02 U740 ( .A0(n400), .A1(n488), .Z(n465));
Q_AN02 U741 ( .A0(n400), .A1(n490), .Z(n466));
Q_AN02 U742 ( .A0(n400), .A1(n492), .Z(n467));
Q_NR02 U743 ( .A0(n397), .A1(dccFrameFill[0]), .Z(n468));
Q_AN02 U744 ( .A0(n470), .A1(n469), .Z(n397));
Q_AN03 U745 ( .A0(n473), .A1(n472), .A2(n471), .Z(n469));
Q_AN03 U746 ( .A0(n476), .A1(n475), .A2(n474), .Z(n470));
Q_AN03 U747 ( .A0(n479), .A1(n478), .A2(n477), .Z(n471));
Q_XNR2 U748 ( .A0(n480), .A1(DccFrameCycle[7]), .Z(n472));
Q_XNR2 U749 ( .A0(n482), .A1(DccFrameCycle[6]), .Z(n473));
Q_XNR2 U750 ( .A0(n484), .A1(DccFrameCycle[5]), .Z(n474));
Q_XNR2 U751 ( .A0(n486), .A1(DccFrameCycle[4]), .Z(n475));
Q_XNR2 U752 ( .A0(n488), .A1(DccFrameCycle[3]), .Z(n476));
Q_XNR2 U753 ( .A0(n490), .A1(DccFrameCycle[2]), .Z(n477));
Q_XNR2 U754 ( .A0(n492), .A1(DccFrameCycle[1]), .Z(n478));
Q_XOR2 U755 ( .A0(dccFrameFill[0]), .A1(DccFrameCycle[0]), .Z(n479));
Q_XOR2 U756 ( .A0(dccFrameFill[7]), .A1(n481), .Z(n480));
Q_AD01HF U757 ( .A0(dccFrameFill[6]), .B0(n483), .S(n482), .CO(n481));
Q_AD01HF U758 ( .A0(dccFrameFill[5]), .B0(n485), .S(n484), .CO(n483));
Q_AD01HF U759 ( .A0(dccFrameFill[4]), .B0(n487), .S(n486), .CO(n485));
Q_AD01HF U760 ( .A0(dccFrameFill[3]), .B0(n489), .S(n488), .CO(n487));
Q_AD01HF U761 ( .A0(dccFrameFill[2]), .B0(n491), .S(n490), .CO(n489));
Q_AD01HF U762 ( .A0(dccFrameFill[1]), .B0(dccFrameFill[0]), .S(n492), .CO(n491));
Q_OR02 U763 ( .A0(n494), .A1(n493), .Z(n398));
Q_OR03 U764 ( .A0(DccFrameCycle[1]), .A1(DccFrameCycle[0]), .A2(n495), .Z(n493));
Q_OR03 U765 ( .A0(DccFrameCycle[4]), .A1(DccFrameCycle[3]), .A2(DccFrameCycle[2]), .Z(n494));
Q_OR03 U766 ( .A0(DccFrameCycle[7]), .A1(DccFrameCycle[6]), .A2(DccFrameCycle[5]), .Z(n495));
Q_INV U767 ( .A(uClkT), .Z(n496));
Q_FDP0UA U768 ( .D(n496), .QTFCLK( ), .Q(uClkT));
Q_INV U769 ( .A(holdEcmTb), .Z(n497));
Q_AN02 U770 ( .A0(n497), .A1(n3979), .Z(n498));
Q_MX02 U771 ( .S(n498), .A0(holdEcmTb), .A1(holdEcmSync), .Z(n499));
Q_FDP0UA U772 ( .D(n499), .QTFCLK( ), .Q(holdEcmSync));
Q_AN02 U773 ( .A0(ptxHoldEcm), .A1(xcRecordOn), .Z(n500));
Q_FDP0UA U774 ( .D(n500), .QTFCLK( ), .Q(holdEcmPtxOn));
Q_FDP0UA U775 ( .D(ecmNotSync), .QTFCLK( ), .Q(ecmNotSyncD));
Q_FDP0UA U776 ( .D(ecmOn), .QTFCLK( ), .Q(ecmOnD));
Q_FDP0UA U777 ( .D(anyStop), .QTFCLK( ), .Q(ptxStop));
Q_INV U778 ( .A(evalOnC), .Z(n503));
Q_OR02 U779 ( .A0(GFbusy), .A1(n503), .Z(n504));
Q_MX02 U780 ( .S(n501), .A0(Gfifo2Sync[0]), .A1(n568), .Z(n505));
Q_FDP0UA U781 ( .D(n505), .QTFCLK( ), .Q(Gfifo2Sync[0]));
Q_MX02 U782 ( .S(n501), .A0(Gfifo2Sync[1]), .A1(n567), .Z(n506));
Q_FDP0UA U783 ( .D(n506), .QTFCLK( ), .Q(Gfifo2Sync[1]));
Q_MX02 U784 ( .S(n501), .A0(Gfifo2Sync[2]), .A1(n566), .Z(n507));
Q_FDP0UA U785 ( .D(n507), .QTFCLK( ), .Q(Gfifo2Sync[2]));
Q_MX02 U786 ( .S(n501), .A0(Gfifo2Sync[3]), .A1(n565), .Z(n508));
Q_FDP0UA U787 ( .D(n508), .QTFCLK( ), .Q(Gfifo2Sync[3]));
Q_MX02 U788 ( .S(n501), .A0(Gfifo2Sync[4]), .A1(n564), .Z(n509));
Q_FDP0UA U789 ( .D(n509), .QTFCLK( ), .Q(Gfifo2Sync[4]));
Q_MX02 U790 ( .S(n501), .A0(Gfifo2Sync[5]), .A1(n563), .Z(n510));
Q_FDP0UA U791 ( .D(n510), .QTFCLK( ), .Q(Gfifo2Sync[5]));
Q_MX02 U792 ( .S(n501), .A0(Gfifo2Sync[6]), .A1(n562), .Z(n511));
Q_FDP0UA U793 ( .D(n511), .QTFCLK( ), .Q(Gfifo2Sync[6]));
Q_MX02 U794 ( .S(n501), .A0(Gfifo2Sync[7]), .A1(n561), .Z(n512));
Q_FDP0UA U795 ( .D(n512), .QTFCLK( ), .Q(Gfifo2Sync[7]));
Q_MX02 U796 ( .S(n501), .A0(Gfifo2Sync[8]), .A1(n560), .Z(n513));
Q_FDP0UA U797 ( .D(n513), .QTFCLK( ), .Q(Gfifo2Sync[8]));
Q_MX02 U798 ( .S(n501), .A0(Gfifo2Sync[9]), .A1(n559), .Z(n514));
Q_FDP0UA U799 ( .D(n514), .QTFCLK( ), .Q(Gfifo2Sync[9]));
Q_MX02 U800 ( .S(n501), .A0(Gfifo2Sync[10]), .A1(n558), .Z(n515));
Q_FDP0UA U801 ( .D(n515), .QTFCLK( ), .Q(Gfifo2Sync[10]));
Q_MX02 U802 ( .S(n501), .A0(Gfifo2Sync[11]), .A1(n557), .Z(n516));
Q_FDP0UA U803 ( .D(n516), .QTFCLK( ), .Q(Gfifo2Sync[11]));
Q_MX02 U804 ( .S(n501), .A0(Gfifo2Sync[12]), .A1(n556), .Z(n517));
Q_FDP0UA U805 ( .D(n517), .QTFCLK( ), .Q(Gfifo2Sync[12]));
Q_MX02 U806 ( .S(n501), .A0(Gfifo2Sync[13]), .A1(n555), .Z(n518));
Q_FDP0UA U807 ( .D(n518), .QTFCLK( ), .Q(Gfifo2Sync[13]));
Q_MX02 U808 ( .S(n501), .A0(Gfifo2Sync[14]), .A1(n554), .Z(n519));
Q_FDP0UA U809 ( .D(n519), .QTFCLK( ), .Q(Gfifo2Sync[14]));
Q_MX02 U810 ( .S(n501), .A0(Gfifo2Sync[15]), .A1(n553), .Z(n520));
Q_FDP0UA U811 ( .D(n520), .QTFCLK( ), .Q(Gfifo2Sync[15]));
Q_MX02 U812 ( .S(n502), .A0(Fck2Sync[0]), .A1(n552), .Z(n521));
Q_FDP0UA U813 ( .D(n521), .QTFCLK( ), .Q(Fck2Sync[0]));
Q_MX02 U814 ( .S(n502), .A0(Fck2Sync[1]), .A1(n551), .Z(n522));
Q_FDP0UA U815 ( .D(n522), .QTFCLK( ), .Q(Fck2Sync[1]));
Q_MX02 U816 ( .S(n502), .A0(Fck2Sync[2]), .A1(n550), .Z(n523));
Q_FDP0UA U817 ( .D(n523), .QTFCLK( ), .Q(Fck2Sync[2]));
Q_MX02 U818 ( .S(n502), .A0(Fck2Sync[3]), .A1(n549), .Z(n524));
Q_FDP0UA U819 ( .D(n524), .QTFCLK( ), .Q(Fck2Sync[3]));
Q_MX02 U820 ( .S(n502), .A0(Fck2Sync[4]), .A1(n548), .Z(n525));
Q_FDP0UA U821 ( .D(n525), .QTFCLK( ), .Q(Fck2Sync[4]));
Q_MX02 U822 ( .S(n502), .A0(Fck2Sync[5]), .A1(n547), .Z(n526));
Q_FDP0UA U823 ( .D(n526), .QTFCLK( ), .Q(Fck2Sync[5]));
Q_MX02 U824 ( .S(n502), .A0(Fck2Sync[6]), .A1(n546), .Z(n527));
Q_FDP0UA U825 ( .D(n527), .QTFCLK( ), .Q(Fck2Sync[6]));
Q_MX02 U826 ( .S(n502), .A0(Fck2Sync[7]), .A1(n545), .Z(n528));
Q_FDP0UA U827 ( .D(n528), .QTFCLK( ), .Q(Fck2Sync[7]));
Q_MX02 U828 ( .S(n502), .A0(Fck2Sync[8]), .A1(n544), .Z(n529));
Q_FDP0UA U829 ( .D(n529), .QTFCLK( ), .Q(Fck2Sync[8]));
Q_MX02 U830 ( .S(n502), .A0(Fck2Sync[9]), .A1(n543), .Z(n530));
Q_FDP0UA U831 ( .D(n530), .QTFCLK( ), .Q(Fck2Sync[9]));
Q_MX02 U832 ( .S(n502), .A0(Fck2Sync[10]), .A1(n542), .Z(n531));
Q_FDP0UA U833 ( .D(n531), .QTFCLK( ), .Q(Fck2Sync[10]));
Q_MX02 U834 ( .S(n502), .A0(Fck2Sync[11]), .A1(n541), .Z(n532));
Q_FDP0UA U835 ( .D(n532), .QTFCLK( ), .Q(Fck2Sync[11]));
Q_MX02 U836 ( .S(n502), .A0(Fck2Sync[12]), .A1(n540), .Z(n533));
Q_FDP0UA U837 ( .D(n533), .QTFCLK( ), .Q(Fck2Sync[12]));
Q_MX02 U838 ( .S(n502), .A0(Fck2Sync[13]), .A1(n539), .Z(n534));
Q_FDP0UA U839 ( .D(n534), .QTFCLK( ), .Q(Fck2Sync[13]));
Q_MX02 U840 ( .S(n502), .A0(Fck2Sync[14]), .A1(n538), .Z(n535));
Q_FDP0UA U841 ( .D(n535), .QTFCLK( ), .Q(Fck2Sync[14]));
Q_MX02 U842 ( .S(n502), .A0(Fck2Sync[15]), .A1(n537), .Z(n536));
Q_FDP0UA U843 ( .D(n536), .QTFCLK( ), .Q(Fck2Sync[15]));
Q_MX02 U844 ( .S(evalOnC), .A0(maxFck2Sync[15]), .A1(n599), .Z(n537));
Q_MX02 U845 ( .S(evalOnC), .A0(maxFck2Sync[14]), .A1(n601), .Z(n538));
Q_MX02 U846 ( .S(evalOnC), .A0(maxFck2Sync[13]), .A1(n603), .Z(n539));
Q_MX02 U847 ( .S(evalOnC), .A0(maxFck2Sync[12]), .A1(n605), .Z(n540));
Q_MX02 U848 ( .S(evalOnC), .A0(maxFck2Sync[11]), .A1(n607), .Z(n541));
Q_MX02 U849 ( .S(evalOnC), .A0(maxFck2Sync[10]), .A1(n609), .Z(n542));
Q_MX02 U850 ( .S(evalOnC), .A0(maxFck2Sync[9]), .A1(n611), .Z(n543));
Q_MX02 U851 ( .S(evalOnC), .A0(maxFck2Sync[8]), .A1(n613), .Z(n544));
Q_MX02 U852 ( .S(evalOnC), .A0(maxFck2Sync[7]), .A1(n615), .Z(n545));
Q_MX02 U853 ( .S(evalOnC), .A0(maxFck2Sync[6]), .A1(n617), .Z(n546));
Q_MX02 U854 ( .S(evalOnC), .A0(maxFck2Sync[5]), .A1(n619), .Z(n547));
Q_MX02 U855 ( .S(evalOnC), .A0(maxFck2Sync[4]), .A1(n621), .Z(n548));
Q_MX02 U856 ( .S(evalOnC), .A0(maxFck2Sync[3]), .A1(n623), .Z(n549));
Q_MX02 U857 ( .S(evalOnC), .A0(maxFck2Sync[2]), .A1(n625), .Z(n550));
Q_MX02 U858 ( .S(evalOnC), .A0(maxFck2Sync[1]), .A1(n627), .Z(n551));
Q_MX02 U859 ( .S(evalOnC), .A0(maxFck2Sync[0]), .A1(n628), .Z(n552));
Q_MX02 U860 ( .S(n504), .A0(n569), .A1(maxGfifo2Sync[15]), .Z(n553));
Q_MX02 U861 ( .S(n504), .A0(n571), .A1(maxGfifo2Sync[14]), .Z(n554));
Q_MX02 U862 ( .S(n504), .A0(n573), .A1(maxGfifo2Sync[13]), .Z(n555));
Q_MX02 U863 ( .S(n504), .A0(n575), .A1(maxGfifo2Sync[12]), .Z(n556));
Q_MX02 U864 ( .S(n504), .A0(n577), .A1(maxGfifo2Sync[11]), .Z(n557));
Q_MX02 U865 ( .S(n504), .A0(n579), .A1(maxGfifo2Sync[10]), .Z(n558));
Q_MX02 U866 ( .S(n504), .A0(n581), .A1(maxGfifo2Sync[9]), .Z(n559));
Q_MX02 U867 ( .S(n504), .A0(n583), .A1(maxGfifo2Sync[8]), .Z(n560));
Q_MX02 U868 ( .S(n504), .A0(n585), .A1(maxGfifo2Sync[7]), .Z(n561));
Q_MX02 U869 ( .S(n504), .A0(n587), .A1(maxGfifo2Sync[6]), .Z(n562));
Q_MX02 U870 ( .S(n504), .A0(n589), .A1(maxGfifo2Sync[5]), .Z(n563));
Q_MX02 U871 ( .S(n504), .A0(n591), .A1(maxGfifo2Sync[4]), .Z(n564));
Q_MX02 U872 ( .S(n504), .A0(n593), .A1(maxGfifo2Sync[3]), .Z(n565));
Q_MX02 U873 ( .S(n504), .A0(n595), .A1(maxGfifo2Sync[2]), .Z(n566));
Q_MX02 U874 ( .S(n504), .A0(n597), .A1(maxGfifo2Sync[1]), .Z(n567));
Q_MX02 U875 ( .S(n504), .A0(n598), .A1(maxGfifo2Sync[0]), .Z(n568));
Q_XNR2 U876 ( .A0(Gfifo2Sync[15]), .A1(n570), .Z(n569));
Q_OR02 U877 ( .A0(Gfifo2Sync[14]), .A1(n572), .Z(n570));
Q_XNR2 U878 ( .A0(Gfifo2Sync[14]), .A1(n572), .Z(n571));
Q_OR02 U879 ( .A0(Gfifo2Sync[13]), .A1(n574), .Z(n572));
Q_XNR2 U880 ( .A0(Gfifo2Sync[13]), .A1(n574), .Z(n573));
Q_OR02 U881 ( .A0(Gfifo2Sync[12]), .A1(n576), .Z(n574));
Q_XNR2 U882 ( .A0(Gfifo2Sync[12]), .A1(n576), .Z(n575));
Q_OR02 U883 ( .A0(Gfifo2Sync[11]), .A1(n578), .Z(n576));
Q_XNR2 U884 ( .A0(Gfifo2Sync[11]), .A1(n578), .Z(n577));
Q_OR02 U885 ( .A0(Gfifo2Sync[10]), .A1(n580), .Z(n578));
Q_XNR2 U886 ( .A0(Gfifo2Sync[10]), .A1(n580), .Z(n579));
Q_OR02 U887 ( .A0(Gfifo2Sync[9]), .A1(n582), .Z(n580));
Q_XNR2 U888 ( .A0(Gfifo2Sync[9]), .A1(n582), .Z(n581));
Q_OR02 U889 ( .A0(Gfifo2Sync[8]), .A1(n584), .Z(n582));
Q_XNR2 U890 ( .A0(Gfifo2Sync[8]), .A1(n584), .Z(n583));
Q_OR02 U891 ( .A0(Gfifo2Sync[7]), .A1(n586), .Z(n584));
Q_XNR2 U892 ( .A0(Gfifo2Sync[7]), .A1(n586), .Z(n585));
Q_OR02 U893 ( .A0(Gfifo2Sync[6]), .A1(n588), .Z(n586));
Q_XNR2 U894 ( .A0(Gfifo2Sync[6]), .A1(n588), .Z(n587));
Q_OR02 U895 ( .A0(Gfifo2Sync[5]), .A1(n590), .Z(n588));
Q_XNR2 U896 ( .A0(Gfifo2Sync[5]), .A1(n590), .Z(n589));
Q_OR02 U897 ( .A0(Gfifo2Sync[4]), .A1(n592), .Z(n590));
Q_XNR2 U898 ( .A0(Gfifo2Sync[4]), .A1(n592), .Z(n591));
Q_OR02 U899 ( .A0(Gfifo2Sync[3]), .A1(n594), .Z(n592));
Q_XNR2 U900 ( .A0(Gfifo2Sync[3]), .A1(n594), .Z(n593));
Q_OR02 U901 ( .A0(Gfifo2Sync[2]), .A1(n596), .Z(n594));
Q_XNR2 U902 ( .A0(Gfifo2Sync[2]), .A1(n596), .Z(n595));
Q_OR02 U903 ( .A0(Gfifo2Sync[1]), .A1(Gfifo2Sync[0]), .Z(n596));
Q_XNR2 U904 ( .A0(Gfifo2Sync[1]), .A1(Gfifo2Sync[0]), .Z(n597));
Q_INV U905 ( .A(Gfifo2Sync[0]), .Z(n598));
Q_XNR2 U906 ( .A0(Fck2Sync[15]), .A1(n600), .Z(n599));
Q_OR02 U907 ( .A0(Fck2Sync[14]), .A1(n602), .Z(n600));
Q_XNR2 U908 ( .A0(Fck2Sync[14]), .A1(n602), .Z(n601));
Q_OR02 U909 ( .A0(Fck2Sync[13]), .A1(n604), .Z(n602));
Q_XNR2 U910 ( .A0(Fck2Sync[13]), .A1(n604), .Z(n603));
Q_OR02 U911 ( .A0(Fck2Sync[12]), .A1(n606), .Z(n604));
Q_XNR2 U912 ( .A0(Fck2Sync[12]), .A1(n606), .Z(n605));
Q_OR02 U913 ( .A0(Fck2Sync[11]), .A1(n608), .Z(n606));
Q_XNR2 U914 ( .A0(Fck2Sync[11]), .A1(n608), .Z(n607));
Q_OR02 U915 ( .A0(Fck2Sync[10]), .A1(n610), .Z(n608));
Q_XNR2 U916 ( .A0(Fck2Sync[10]), .A1(n610), .Z(n609));
Q_OR02 U917 ( .A0(Fck2Sync[9]), .A1(n612), .Z(n610));
Q_XNR2 U918 ( .A0(Fck2Sync[9]), .A1(n612), .Z(n611));
Q_OR02 U919 ( .A0(Fck2Sync[8]), .A1(n614), .Z(n612));
Q_XNR2 U920 ( .A0(Fck2Sync[8]), .A1(n614), .Z(n613));
Q_OR02 U921 ( .A0(Fck2Sync[7]), .A1(n616), .Z(n614));
Q_XNR2 U922 ( .A0(Fck2Sync[7]), .A1(n616), .Z(n615));
Q_OR02 U923 ( .A0(Fck2Sync[6]), .A1(n618), .Z(n616));
Q_XNR2 U924 ( .A0(Fck2Sync[6]), .A1(n618), .Z(n617));
Q_OR02 U925 ( .A0(Fck2Sync[5]), .A1(n620), .Z(n618));
Q_XNR2 U926 ( .A0(Fck2Sync[5]), .A1(n620), .Z(n619));
Q_OR02 U927 ( .A0(Fck2Sync[4]), .A1(n622), .Z(n620));
Q_XNR2 U928 ( .A0(Fck2Sync[4]), .A1(n622), .Z(n621));
Q_OR02 U929 ( .A0(Fck2Sync[3]), .A1(n624), .Z(n622));
Q_XNR2 U930 ( .A0(Fck2Sync[3]), .A1(n624), .Z(n623));
Q_OR02 U931 ( .A0(Fck2Sync[2]), .A1(n626), .Z(n624));
Q_XNR2 U932 ( .A0(Fck2Sync[2]), .A1(n626), .Z(n625));
Q_OR02 U933 ( .A0(Fck2Sync[1]), .A1(Fck2Sync[0]), .Z(n626));
Q_XNR2 U934 ( .A0(Fck2Sync[1]), .A1(Fck2Sync[0]), .Z(n627));
Q_INV U935 ( .A(Fck2Sync[0]), .Z(n628));
Q_OR03 U936 ( .A0(n630), .A1(n629), .A2(n504), .Z(n501));
Q_OR03 U937 ( .A0(n633), .A1(n632), .A2(n631), .Z(n629));
Q_OR03 U938 ( .A0(Gfifo2Sync[0]), .A1(n635), .A2(n634), .Z(n630));
Q_OR03 U939 ( .A0(Gfifo2Sync[3]), .A1(Gfifo2Sync[2]), .A2(Gfifo2Sync[1]), .Z(n631));
Q_OR03 U940 ( .A0(Gfifo2Sync[6]), .A1(Gfifo2Sync[5]), .A2(Gfifo2Sync[4]), .Z(n632));
Q_OR03 U941 ( .A0(Gfifo2Sync[9]), .A1(Gfifo2Sync[8]), .A2(Gfifo2Sync[7]), .Z(n633));
Q_OR03 U942 ( .A0(Gfifo2Sync[12]), .A1(Gfifo2Sync[11]), .A2(Gfifo2Sync[10]), .Z(n634));
Q_OR03 U943 ( .A0(Gfifo2Sync[15]), .A1(Gfifo2Sync[14]), .A2(Gfifo2Sync[13]), .Z(n635));
Q_OR03 U944 ( .A0(n637), .A1(n636), .A2(n503), .Z(n502));
Q_OR03 U945 ( .A0(n640), .A1(n639), .A2(n638), .Z(n636));
Q_OR03 U946 ( .A0(Fck2Sync[0]), .A1(n642), .A2(n641), .Z(n637));
Q_OR03 U947 ( .A0(Fck2Sync[3]), .A1(Fck2Sync[2]), .A2(Fck2Sync[1]), .Z(n638));
Q_OR03 U948 ( .A0(Fck2Sync[6]), .A1(Fck2Sync[5]), .A2(Fck2Sync[4]), .Z(n639));
Q_OR03 U949 ( .A0(Fck2Sync[9]), .A1(Fck2Sync[8]), .A2(Fck2Sync[7]), .Z(n640));
Q_OR03 U950 ( .A0(Fck2Sync[12]), .A1(Fck2Sync[11]), .A2(Fck2Sync[10]), .Z(n641));
Q_OR03 U951 ( .A0(Fck2Sync[15]), .A1(Fck2Sync[14]), .A2(Fck2Sync[13]), .Z(n642));
Q_FDP0UA U952 ( .D(maxFck2Sync[15]), .QTFCLK( ), .Q(maxFck2Sync[15]));
Q_FDP0UA U953 ( .D(maxFck2Sync[14]), .QTFCLK( ), .Q(maxFck2Sync[14]));
Q_FDP0UA U954 ( .D(maxFck2Sync[13]), .QTFCLK( ), .Q(maxFck2Sync[13]));
Q_FDP0UA U955 ( .D(maxFck2Sync[12]), .QTFCLK( ), .Q(maxFck2Sync[12]));
Q_FDP0UA U956 ( .D(maxFck2Sync[11]), .QTFCLK( ), .Q(maxFck2Sync[11]));
Q_FDP0UA U957 ( .D(maxFck2Sync[10]), .QTFCLK( ), .Q(maxFck2Sync[10]));
Q_FDP0UA U958 ( .D(maxFck2Sync[9]), .QTFCLK( ), .Q(maxFck2Sync[9]));
Q_FDP0UA U959 ( .D(maxFck2Sync[8]), .QTFCLK( ), .Q(maxFck2Sync[8]));
Q_FDP0UA U960 ( .D(maxFck2Sync[7]), .QTFCLK( ), .Q(maxFck2Sync[7]));
Q_FDP0UA U961 ( .D(maxFck2Sync[6]), .QTFCLK( ), .Q(maxFck2Sync[6]));
Q_FDP0UA U962 ( .D(maxFck2Sync[5]), .QTFCLK( ), .Q(maxFck2Sync[5]));
Q_FDP0UA U963 ( .D(maxFck2Sync[4]), .QTFCLK( ), .Q(maxFck2Sync[4]));
Q_FDP0UA U964 ( .D(maxFck2Sync[3]), .QTFCLK( ), .Q(maxFck2Sync[3]));
Q_FDP0UA U965 ( .D(maxFck2Sync[2]), .QTFCLK( ), .Q(maxFck2Sync[2]));
Q_FDP0UA U966 ( .D(maxFck2Sync[1]), .QTFCLK( ), .Q(maxFck2Sync[1]));
Q_FDP0UA U967 ( .D(maxFck2Sync[0]), .QTFCLK( ), .Q(maxFck2Sync[0]));
Q_FDP0UA U968 ( .D(maxGfifo2Sync[15]), .QTFCLK( ), .Q(maxGfifo2Sync[15]));
Q_FDP0UA U969 ( .D(maxGfifo2Sync[14]), .QTFCLK( ), .Q(maxGfifo2Sync[14]));
Q_FDP0UA U970 ( .D(maxGfifo2Sync[13]), .QTFCLK( ), .Q(maxGfifo2Sync[13]));
Q_FDP0UA U971 ( .D(maxGfifo2Sync[12]), .QTFCLK( ), .Q(maxGfifo2Sync[12]));
Q_FDP0UA U972 ( .D(maxGfifo2Sync[11]), .QTFCLK( ), .Q(maxGfifo2Sync[11]));
Q_FDP0UA U973 ( .D(maxGfifo2Sync[10]), .QTFCLK( ), .Q(maxGfifo2Sync[10]));
Q_FDP0UA U974 ( .D(maxGfifo2Sync[9]), .QTFCLK( ), .Q(maxGfifo2Sync[9]));
Q_FDP0UA U975 ( .D(maxGfifo2Sync[8]), .QTFCLK( ), .Q(maxGfifo2Sync[8]));
Q_FDP0UA U976 ( .D(maxGfifo2Sync[7]), .QTFCLK( ), .Q(maxGfifo2Sync[7]));
Q_FDP0UA U977 ( .D(maxGfifo2Sync[6]), .QTFCLK( ), .Q(maxGfifo2Sync[6]));
Q_FDP0UA U978 ( .D(maxGfifo2Sync[5]), .QTFCLK( ), .Q(maxGfifo2Sync[5]));
Q_FDP0UA U979 ( .D(maxGfifo2Sync[4]), .QTFCLK( ), .Q(maxGfifo2Sync[4]));
Q_FDP0UA U980 ( .D(maxGfifo2Sync[3]), .QTFCLK( ), .Q(maxGfifo2Sync[3]));
Q_FDP0UA U981 ( .D(maxGfifo2Sync[2]), .QTFCLK( ), .Q(maxGfifo2Sync[2]));
Q_FDP0UA U982 ( .D(maxGfifo2Sync[1]), .QTFCLK( ), .Q(maxGfifo2Sync[1]));
Q_FDP0UA U983 ( .D(maxGfifo2Sync[0]), .QTFCLK( ), .Q(maxGfifo2Sync[0]));
Q_NR02 U984 ( .A0(GFGBfullBw), .A1(GFGBfullBwD), .Z(n650));
Q_NR02 U985 ( .A0(GFLBfull), .A1(GFLBfullD), .Z(n648));
Q_AN02 U986 ( .A0(n650), .A1(n648), .Z(n647));
Q_AN03 U987 ( .A0(GFbusy), .A1(n503), .A2(n647), .Z(n643));
Q_INV U988 ( .A(n648), .Z(n649));
Q_AN02 U989 ( .A0(n650), .A1(n649), .Z(n644));
Q_INV U990 ( .A(n650), .Z(n645));
Q_NR02 U991 ( .A0(holdEcm), .A1(holdEcmD), .Z(n651));
Q_INV U992 ( .A(n651), .Z(n646));
Q_XOR2 U993 ( .A0(n643), .A1(gfifoTBsyncCnt[0]), .Z(n652));
Q_FDP0UA U994 ( .D(n652), .QTFCLK( ), .Q(gfifoTBsyncCnt[0]));
Q_MX02 U995 ( .S(n643), .A0(gfifoTBsyncCnt[1]), .A1(n1155), .Z(n653));
Q_FDP0UA U996 ( .D(n653), .QTFCLK( ), .Q(gfifoTBsyncCnt[1]));
Q_MX02 U997 ( .S(n643), .A0(gfifoTBsyncCnt[2]), .A1(n1153), .Z(n654));
Q_FDP0UA U998 ( .D(n654), .QTFCLK( ), .Q(gfifoTBsyncCnt[2]));
Q_MX02 U999 ( .S(n643), .A0(gfifoTBsyncCnt[3]), .A1(n1151), .Z(n655));
Q_FDP0UA U1000 ( .D(n655), .QTFCLK( ), .Q(gfifoTBsyncCnt[3]));
Q_MX02 U1001 ( .S(n643), .A0(gfifoTBsyncCnt[4]), .A1(n1149), .Z(n656));
Q_FDP0UA U1002 ( .D(n656), .QTFCLK( ), .Q(gfifoTBsyncCnt[4]));
Q_MX02 U1003 ( .S(n643), .A0(gfifoTBsyncCnt[5]), .A1(n1147), .Z(n657));
Q_FDP0UA U1004 ( .D(n657), .QTFCLK( ), .Q(gfifoTBsyncCnt[5]));
Q_MX02 U1005 ( .S(n643), .A0(gfifoTBsyncCnt[6]), .A1(n1145), .Z(n658));
Q_FDP0UA U1006 ( .D(n658), .QTFCLK( ), .Q(gfifoTBsyncCnt[6]));
Q_MX02 U1007 ( .S(n643), .A0(gfifoTBsyncCnt[7]), .A1(n1143), .Z(n659));
Q_FDP0UA U1008 ( .D(n659), .QTFCLK( ), .Q(gfifoTBsyncCnt[7]));
Q_MX02 U1009 ( .S(n643), .A0(gfifoTBsyncCnt[8]), .A1(n1141), .Z(n660));
Q_FDP0UA U1010 ( .D(n660), .QTFCLK( ), .Q(gfifoTBsyncCnt[8]));
Q_MX02 U1011 ( .S(n643), .A0(gfifoTBsyncCnt[9]), .A1(n1139), .Z(n661));
Q_FDP0UA U1012 ( .D(n661), .QTFCLK( ), .Q(gfifoTBsyncCnt[9]));
Q_MX02 U1013 ( .S(n643), .A0(gfifoTBsyncCnt[10]), .A1(n1137), .Z(n662));
Q_FDP0UA U1014 ( .D(n662), .QTFCLK( ), .Q(gfifoTBsyncCnt[10]));
Q_MX02 U1015 ( .S(n643), .A0(gfifoTBsyncCnt[11]), .A1(n1135), .Z(n663));
Q_FDP0UA U1016 ( .D(n663), .QTFCLK( ), .Q(gfifoTBsyncCnt[11]));
Q_MX02 U1017 ( .S(n643), .A0(gfifoTBsyncCnt[12]), .A1(n1133), .Z(n664));
Q_FDP0UA U1018 ( .D(n664), .QTFCLK( ), .Q(gfifoTBsyncCnt[12]));
Q_MX02 U1019 ( .S(n643), .A0(gfifoTBsyncCnt[13]), .A1(n1131), .Z(n665));
Q_FDP0UA U1020 ( .D(n665), .QTFCLK( ), .Q(gfifoTBsyncCnt[13]));
Q_MX02 U1021 ( .S(n643), .A0(gfifoTBsyncCnt[14]), .A1(n1129), .Z(n666));
Q_FDP0UA U1022 ( .D(n666), .QTFCLK( ), .Q(gfifoTBsyncCnt[14]));
Q_MX02 U1023 ( .S(n643), .A0(gfifoTBsyncCnt[15]), .A1(n1127), .Z(n667));
Q_FDP0UA U1024 ( .D(n667), .QTFCLK( ), .Q(gfifoTBsyncCnt[15]));
Q_MX02 U1025 ( .S(n643), .A0(gfifoTBsyncCnt[16]), .A1(n1125), .Z(n668));
Q_FDP0UA U1026 ( .D(n668), .QTFCLK( ), .Q(gfifoTBsyncCnt[16]));
Q_MX02 U1027 ( .S(n643), .A0(gfifoTBsyncCnt[17]), .A1(n1123), .Z(n669));
Q_FDP0UA U1028 ( .D(n669), .QTFCLK( ), .Q(gfifoTBsyncCnt[17]));
Q_MX02 U1029 ( .S(n643), .A0(gfifoTBsyncCnt[18]), .A1(n1121), .Z(n670));
Q_FDP0UA U1030 ( .D(n670), .QTFCLK( ), .Q(gfifoTBsyncCnt[18]));
Q_MX02 U1031 ( .S(n643), .A0(gfifoTBsyncCnt[19]), .A1(n1119), .Z(n671));
Q_FDP0UA U1032 ( .D(n671), .QTFCLK( ), .Q(gfifoTBsyncCnt[19]));
Q_MX02 U1033 ( .S(n643), .A0(gfifoTBsyncCnt[20]), .A1(n1117), .Z(n672));
Q_FDP0UA U1034 ( .D(n672), .QTFCLK( ), .Q(gfifoTBsyncCnt[20]));
Q_MX02 U1035 ( .S(n643), .A0(gfifoTBsyncCnt[21]), .A1(n1115), .Z(n673));
Q_FDP0UA U1036 ( .D(n673), .QTFCLK( ), .Q(gfifoTBsyncCnt[21]));
Q_MX02 U1037 ( .S(n643), .A0(gfifoTBsyncCnt[22]), .A1(n1113), .Z(n674));
Q_FDP0UA U1038 ( .D(n674), .QTFCLK( ), .Q(gfifoTBsyncCnt[22]));
Q_MX02 U1039 ( .S(n643), .A0(gfifoTBsyncCnt[23]), .A1(n1111), .Z(n675));
Q_FDP0UA U1040 ( .D(n675), .QTFCLK( ), .Q(gfifoTBsyncCnt[23]));
Q_MX02 U1041 ( .S(n643), .A0(gfifoTBsyncCnt[24]), .A1(n1109), .Z(n676));
Q_FDP0UA U1042 ( .D(n676), .QTFCLK( ), .Q(gfifoTBsyncCnt[24]));
Q_MX02 U1043 ( .S(n643), .A0(gfifoTBsyncCnt[25]), .A1(n1107), .Z(n677));
Q_FDP0UA U1044 ( .D(n677), .QTFCLK( ), .Q(gfifoTBsyncCnt[25]));
Q_MX02 U1045 ( .S(n643), .A0(gfifoTBsyncCnt[26]), .A1(n1105), .Z(n678));
Q_FDP0UA U1046 ( .D(n678), .QTFCLK( ), .Q(gfifoTBsyncCnt[26]));
Q_MX02 U1047 ( .S(n643), .A0(gfifoTBsyncCnt[27]), .A1(n1103), .Z(n679));
Q_FDP0UA U1048 ( .D(n679), .QTFCLK( ), .Q(gfifoTBsyncCnt[27]));
Q_MX02 U1049 ( .S(n643), .A0(gfifoTBsyncCnt[28]), .A1(n1101), .Z(n680));
Q_FDP0UA U1050 ( .D(n680), .QTFCLK( ), .Q(gfifoTBsyncCnt[28]));
Q_MX02 U1051 ( .S(n643), .A0(gfifoTBsyncCnt[29]), .A1(n1099), .Z(n681));
Q_FDP0UA U1052 ( .D(n681), .QTFCLK( ), .Q(gfifoTBsyncCnt[29]));
Q_MX02 U1053 ( .S(n643), .A0(gfifoTBsyncCnt[30]), .A1(n1097), .Z(n682));
Q_FDP0UA U1054 ( .D(n682), .QTFCLK( ), .Q(gfifoTBsyncCnt[30]));
Q_MX02 U1055 ( .S(n643), .A0(gfifoTBsyncCnt[31]), .A1(n1095), .Z(n683));
Q_FDP0UA U1056 ( .D(n683), .QTFCLK( ), .Q(gfifoTBsyncCnt[31]));
Q_MX02 U1057 ( .S(n643), .A0(gfifoTBsyncCnt[32]), .A1(n1093), .Z(n684));
Q_FDP0UA U1058 ( .D(n684), .QTFCLK( ), .Q(gfifoTBsyncCnt[32]));
Q_MX02 U1059 ( .S(n643), .A0(gfifoTBsyncCnt[33]), .A1(n1091), .Z(n685));
Q_FDP0UA U1060 ( .D(n685), .QTFCLK( ), .Q(gfifoTBsyncCnt[33]));
Q_MX02 U1061 ( .S(n643), .A0(gfifoTBsyncCnt[34]), .A1(n1089), .Z(n686));
Q_FDP0UA U1062 ( .D(n686), .QTFCLK( ), .Q(gfifoTBsyncCnt[34]));
Q_MX02 U1063 ( .S(n643), .A0(gfifoTBsyncCnt[35]), .A1(n1087), .Z(n687));
Q_FDP0UA U1064 ( .D(n687), .QTFCLK( ), .Q(gfifoTBsyncCnt[35]));
Q_MX02 U1065 ( .S(n643), .A0(gfifoTBsyncCnt[36]), .A1(n1085), .Z(n688));
Q_FDP0UA U1066 ( .D(n688), .QTFCLK( ), .Q(gfifoTBsyncCnt[36]));
Q_MX02 U1067 ( .S(n643), .A0(gfifoTBsyncCnt[37]), .A1(n1083), .Z(n689));
Q_FDP0UA U1068 ( .D(n689), .QTFCLK( ), .Q(gfifoTBsyncCnt[37]));
Q_MX02 U1069 ( .S(n643), .A0(gfifoTBsyncCnt[38]), .A1(n1081), .Z(n690));
Q_FDP0UA U1070 ( .D(n690), .QTFCLK( ), .Q(gfifoTBsyncCnt[38]));
Q_MX02 U1071 ( .S(n643), .A0(gfifoTBsyncCnt[39]), .A1(n1079), .Z(n691));
Q_FDP0UA U1072 ( .D(n691), .QTFCLK( ), .Q(gfifoTBsyncCnt[39]));
Q_MX02 U1073 ( .S(n643), .A0(gfifoTBsyncCnt[40]), .A1(n1077), .Z(n692));
Q_FDP0UA U1074 ( .D(n692), .QTFCLK( ), .Q(gfifoTBsyncCnt[40]));
Q_MX02 U1075 ( .S(n643), .A0(gfifoTBsyncCnt[41]), .A1(n1075), .Z(n693));
Q_FDP0UA U1076 ( .D(n693), .QTFCLK( ), .Q(gfifoTBsyncCnt[41]));
Q_MX02 U1077 ( .S(n643), .A0(gfifoTBsyncCnt[42]), .A1(n1073), .Z(n694));
Q_FDP0UA U1078 ( .D(n694), .QTFCLK( ), .Q(gfifoTBsyncCnt[42]));
Q_MX02 U1079 ( .S(n643), .A0(gfifoTBsyncCnt[43]), .A1(n1071), .Z(n695));
Q_FDP0UA U1080 ( .D(n695), .QTFCLK( ), .Q(gfifoTBsyncCnt[43]));
Q_MX02 U1081 ( .S(n643), .A0(gfifoTBsyncCnt[44]), .A1(n1069), .Z(n696));
Q_FDP0UA U1082 ( .D(n696), .QTFCLK( ), .Q(gfifoTBsyncCnt[44]));
Q_MX02 U1083 ( .S(n643), .A0(gfifoTBsyncCnt[45]), .A1(n1067), .Z(n697));
Q_FDP0UA U1084 ( .D(n697), .QTFCLK( ), .Q(gfifoTBsyncCnt[45]));
Q_MX02 U1085 ( .S(n643), .A0(gfifoTBsyncCnt[46]), .A1(n1065), .Z(n698));
Q_FDP0UA U1086 ( .D(n698), .QTFCLK( ), .Q(gfifoTBsyncCnt[46]));
Q_MX02 U1087 ( .S(n643), .A0(gfifoTBsyncCnt[47]), .A1(n1063), .Z(n699));
Q_FDP0UA U1088 ( .D(n699), .QTFCLK( ), .Q(gfifoTBsyncCnt[47]));
Q_MX02 U1089 ( .S(n643), .A0(gfifoTBsyncCnt[48]), .A1(n1061), .Z(n700));
Q_FDP0UA U1090 ( .D(n700), .QTFCLK( ), .Q(gfifoTBsyncCnt[48]));
Q_MX02 U1091 ( .S(n643), .A0(gfifoTBsyncCnt[49]), .A1(n1059), .Z(n701));
Q_FDP0UA U1092 ( .D(n701), .QTFCLK( ), .Q(gfifoTBsyncCnt[49]));
Q_MX02 U1093 ( .S(n643), .A0(gfifoTBsyncCnt[50]), .A1(n1057), .Z(n702));
Q_FDP0UA U1094 ( .D(n702), .QTFCLK( ), .Q(gfifoTBsyncCnt[50]));
Q_MX02 U1095 ( .S(n643), .A0(gfifoTBsyncCnt[51]), .A1(n1055), .Z(n703));
Q_FDP0UA U1096 ( .D(n703), .QTFCLK( ), .Q(gfifoTBsyncCnt[51]));
Q_MX02 U1097 ( .S(n643), .A0(gfifoTBsyncCnt[52]), .A1(n1053), .Z(n704));
Q_FDP0UA U1098 ( .D(n704), .QTFCLK( ), .Q(gfifoTBsyncCnt[52]));
Q_MX02 U1099 ( .S(n643), .A0(gfifoTBsyncCnt[53]), .A1(n1051), .Z(n705));
Q_FDP0UA U1100 ( .D(n705), .QTFCLK( ), .Q(gfifoTBsyncCnt[53]));
Q_MX02 U1101 ( .S(n643), .A0(gfifoTBsyncCnt[54]), .A1(n1049), .Z(n706));
Q_FDP0UA U1102 ( .D(n706), .QTFCLK( ), .Q(gfifoTBsyncCnt[54]));
Q_MX02 U1103 ( .S(n643), .A0(gfifoTBsyncCnt[55]), .A1(n1047), .Z(n707));
Q_FDP0UA U1104 ( .D(n707), .QTFCLK( ), .Q(gfifoTBsyncCnt[55]));
Q_MX02 U1105 ( .S(n643), .A0(gfifoTBsyncCnt[56]), .A1(n1045), .Z(n708));
Q_FDP0UA U1106 ( .D(n708), .QTFCLK( ), .Q(gfifoTBsyncCnt[56]));
Q_MX02 U1107 ( .S(n643), .A0(gfifoTBsyncCnt[57]), .A1(n1043), .Z(n709));
Q_FDP0UA U1108 ( .D(n709), .QTFCLK( ), .Q(gfifoTBsyncCnt[57]));
Q_MX02 U1109 ( .S(n643), .A0(gfifoTBsyncCnt[58]), .A1(n1041), .Z(n710));
Q_FDP0UA U1110 ( .D(n710), .QTFCLK( ), .Q(gfifoTBsyncCnt[58]));
Q_MX02 U1111 ( .S(n643), .A0(gfifoTBsyncCnt[59]), .A1(n1039), .Z(n711));
Q_FDP0UA U1112 ( .D(n711), .QTFCLK( ), .Q(gfifoTBsyncCnt[59]));
Q_MX02 U1113 ( .S(n643), .A0(gfifoTBsyncCnt[60]), .A1(n1037), .Z(n712));
Q_FDP0UA U1114 ( .D(n712), .QTFCLK( ), .Q(gfifoTBsyncCnt[60]));
Q_MX02 U1115 ( .S(n643), .A0(gfifoTBsyncCnt[61]), .A1(n1035), .Z(n713));
Q_FDP0UA U1116 ( .D(n713), .QTFCLK( ), .Q(gfifoTBsyncCnt[61]));
Q_MX02 U1117 ( .S(n643), .A0(gfifoTBsyncCnt[62]), .A1(n1033), .Z(n714));
Q_FDP0UA U1118 ( .D(n714), .QTFCLK( ), .Q(gfifoTBsyncCnt[62]));
Q_FDP0UA U1119 ( .D(n715), .QTFCLK( ), .Q(gfifoTBsyncCnt[63]));
Q_XOR2 U1120 ( .A0(n644), .A1(gfifoLBfullCnt[0]), .Z(n716));
Q_FDP0UA U1121 ( .D(n716), .QTFCLK( ), .Q(gfifoLBfullCnt[0]));
Q_MX02 U1122 ( .S(n644), .A0(gfifoLBfullCnt[1]), .A1(n1279), .Z(n717));
Q_FDP0UA U1123 ( .D(n717), .QTFCLK( ), .Q(gfifoLBfullCnt[1]));
Q_MX02 U1124 ( .S(n644), .A0(gfifoLBfullCnt[2]), .A1(n1277), .Z(n718));
Q_FDP0UA U1125 ( .D(n718), .QTFCLK( ), .Q(gfifoLBfullCnt[2]));
Q_MX02 U1126 ( .S(n644), .A0(gfifoLBfullCnt[3]), .A1(n1275), .Z(n719));
Q_FDP0UA U1127 ( .D(n719), .QTFCLK( ), .Q(gfifoLBfullCnt[3]));
Q_MX02 U1128 ( .S(n644), .A0(gfifoLBfullCnt[4]), .A1(n1273), .Z(n720));
Q_FDP0UA U1129 ( .D(n720), .QTFCLK( ), .Q(gfifoLBfullCnt[4]));
Q_MX02 U1130 ( .S(n644), .A0(gfifoLBfullCnt[5]), .A1(n1271), .Z(n721));
Q_FDP0UA U1131 ( .D(n721), .QTFCLK( ), .Q(gfifoLBfullCnt[5]));
Q_MX02 U1132 ( .S(n644), .A0(gfifoLBfullCnt[6]), .A1(n1269), .Z(n722));
Q_FDP0UA U1133 ( .D(n722), .QTFCLK( ), .Q(gfifoLBfullCnt[6]));
Q_MX02 U1134 ( .S(n644), .A0(gfifoLBfullCnt[7]), .A1(n1267), .Z(n723));
Q_FDP0UA U1135 ( .D(n723), .QTFCLK( ), .Q(gfifoLBfullCnt[7]));
Q_MX02 U1136 ( .S(n644), .A0(gfifoLBfullCnt[8]), .A1(n1265), .Z(n724));
Q_FDP0UA U1137 ( .D(n724), .QTFCLK( ), .Q(gfifoLBfullCnt[8]));
Q_MX02 U1138 ( .S(n644), .A0(gfifoLBfullCnt[9]), .A1(n1263), .Z(n725));
Q_FDP0UA U1139 ( .D(n725), .QTFCLK( ), .Q(gfifoLBfullCnt[9]));
Q_MX02 U1140 ( .S(n644), .A0(gfifoLBfullCnt[10]), .A1(n1261), .Z(n726));
Q_FDP0UA U1141 ( .D(n726), .QTFCLK( ), .Q(gfifoLBfullCnt[10]));
Q_MX02 U1142 ( .S(n644), .A0(gfifoLBfullCnt[11]), .A1(n1259), .Z(n727));
Q_FDP0UA U1143 ( .D(n727), .QTFCLK( ), .Q(gfifoLBfullCnt[11]));
Q_MX02 U1144 ( .S(n644), .A0(gfifoLBfullCnt[12]), .A1(n1257), .Z(n728));
Q_FDP0UA U1145 ( .D(n728), .QTFCLK( ), .Q(gfifoLBfullCnt[12]));
Q_MX02 U1146 ( .S(n644), .A0(gfifoLBfullCnt[13]), .A1(n1255), .Z(n729));
Q_FDP0UA U1147 ( .D(n729), .QTFCLK( ), .Q(gfifoLBfullCnt[13]));
Q_MX02 U1148 ( .S(n644), .A0(gfifoLBfullCnt[14]), .A1(n1253), .Z(n730));
Q_FDP0UA U1149 ( .D(n730), .QTFCLK( ), .Q(gfifoLBfullCnt[14]));
Q_MX02 U1150 ( .S(n644), .A0(gfifoLBfullCnt[15]), .A1(n1251), .Z(n731));
Q_FDP0UA U1151 ( .D(n731), .QTFCLK( ), .Q(gfifoLBfullCnt[15]));
Q_MX02 U1152 ( .S(n644), .A0(gfifoLBfullCnt[16]), .A1(n1249), .Z(n732));
Q_FDP0UA U1153 ( .D(n732), .QTFCLK( ), .Q(gfifoLBfullCnt[16]));
Q_MX02 U1154 ( .S(n644), .A0(gfifoLBfullCnt[17]), .A1(n1247), .Z(n733));
Q_FDP0UA U1155 ( .D(n733), .QTFCLK( ), .Q(gfifoLBfullCnt[17]));
Q_MX02 U1156 ( .S(n644), .A0(gfifoLBfullCnt[18]), .A1(n1245), .Z(n734));
Q_FDP0UA U1157 ( .D(n734), .QTFCLK( ), .Q(gfifoLBfullCnt[18]));
Q_MX02 U1158 ( .S(n644), .A0(gfifoLBfullCnt[19]), .A1(n1243), .Z(n735));
Q_FDP0UA U1159 ( .D(n735), .QTFCLK( ), .Q(gfifoLBfullCnt[19]));
Q_MX02 U1160 ( .S(n644), .A0(gfifoLBfullCnt[20]), .A1(n1241), .Z(n736));
Q_FDP0UA U1161 ( .D(n736), .QTFCLK( ), .Q(gfifoLBfullCnt[20]));
Q_MX02 U1162 ( .S(n644), .A0(gfifoLBfullCnt[21]), .A1(n1239), .Z(n737));
Q_FDP0UA U1163 ( .D(n737), .QTFCLK( ), .Q(gfifoLBfullCnt[21]));
Q_MX02 U1164 ( .S(n644), .A0(gfifoLBfullCnt[22]), .A1(n1237), .Z(n738));
Q_FDP0UA U1165 ( .D(n738), .QTFCLK( ), .Q(gfifoLBfullCnt[22]));
Q_MX02 U1166 ( .S(n644), .A0(gfifoLBfullCnt[23]), .A1(n1235), .Z(n739));
Q_FDP0UA U1167 ( .D(n739), .QTFCLK( ), .Q(gfifoLBfullCnt[23]));
Q_MX02 U1168 ( .S(n644), .A0(gfifoLBfullCnt[24]), .A1(n1233), .Z(n740));
Q_FDP0UA U1169 ( .D(n740), .QTFCLK( ), .Q(gfifoLBfullCnt[24]));
Q_MX02 U1170 ( .S(n644), .A0(gfifoLBfullCnt[25]), .A1(n1231), .Z(n741));
Q_FDP0UA U1171 ( .D(n741), .QTFCLK( ), .Q(gfifoLBfullCnt[25]));
Q_MX02 U1172 ( .S(n644), .A0(gfifoLBfullCnt[26]), .A1(n1229), .Z(n742));
Q_FDP0UA U1173 ( .D(n742), .QTFCLK( ), .Q(gfifoLBfullCnt[26]));
Q_MX02 U1174 ( .S(n644), .A0(gfifoLBfullCnt[27]), .A1(n1227), .Z(n743));
Q_FDP0UA U1175 ( .D(n743), .QTFCLK( ), .Q(gfifoLBfullCnt[27]));
Q_MX02 U1176 ( .S(n644), .A0(gfifoLBfullCnt[28]), .A1(n1225), .Z(n744));
Q_FDP0UA U1177 ( .D(n744), .QTFCLK( ), .Q(gfifoLBfullCnt[28]));
Q_MX02 U1178 ( .S(n644), .A0(gfifoLBfullCnt[29]), .A1(n1223), .Z(n745));
Q_FDP0UA U1179 ( .D(n745), .QTFCLK( ), .Q(gfifoLBfullCnt[29]));
Q_MX02 U1180 ( .S(n644), .A0(gfifoLBfullCnt[30]), .A1(n1221), .Z(n746));
Q_FDP0UA U1181 ( .D(n746), .QTFCLK( ), .Q(gfifoLBfullCnt[30]));
Q_MX02 U1182 ( .S(n644), .A0(gfifoLBfullCnt[31]), .A1(n1219), .Z(n747));
Q_FDP0UA U1183 ( .D(n747), .QTFCLK( ), .Q(gfifoLBfullCnt[31]));
Q_MX02 U1184 ( .S(n644), .A0(gfifoLBfullCnt[32]), .A1(n1217), .Z(n748));
Q_FDP0UA U1185 ( .D(n748), .QTFCLK( ), .Q(gfifoLBfullCnt[32]));
Q_MX02 U1186 ( .S(n644), .A0(gfifoLBfullCnt[33]), .A1(n1215), .Z(n749));
Q_FDP0UA U1187 ( .D(n749), .QTFCLK( ), .Q(gfifoLBfullCnt[33]));
Q_MX02 U1188 ( .S(n644), .A0(gfifoLBfullCnt[34]), .A1(n1213), .Z(n750));
Q_FDP0UA U1189 ( .D(n750), .QTFCLK( ), .Q(gfifoLBfullCnt[34]));
Q_MX02 U1190 ( .S(n644), .A0(gfifoLBfullCnt[35]), .A1(n1211), .Z(n751));
Q_FDP0UA U1191 ( .D(n751), .QTFCLK( ), .Q(gfifoLBfullCnt[35]));
Q_MX02 U1192 ( .S(n644), .A0(gfifoLBfullCnt[36]), .A1(n1209), .Z(n752));
Q_FDP0UA U1193 ( .D(n752), .QTFCLK( ), .Q(gfifoLBfullCnt[36]));
Q_MX02 U1194 ( .S(n644), .A0(gfifoLBfullCnt[37]), .A1(n1207), .Z(n753));
Q_FDP0UA U1195 ( .D(n753), .QTFCLK( ), .Q(gfifoLBfullCnt[37]));
Q_MX02 U1196 ( .S(n644), .A0(gfifoLBfullCnt[38]), .A1(n1205), .Z(n754));
Q_FDP0UA U1197 ( .D(n754), .QTFCLK( ), .Q(gfifoLBfullCnt[38]));
Q_MX02 U1198 ( .S(n644), .A0(gfifoLBfullCnt[39]), .A1(n1203), .Z(n755));
Q_FDP0UA U1199 ( .D(n755), .QTFCLK( ), .Q(gfifoLBfullCnt[39]));
Q_MX02 U1200 ( .S(n644), .A0(gfifoLBfullCnt[40]), .A1(n1201), .Z(n756));
Q_FDP0UA U1201 ( .D(n756), .QTFCLK( ), .Q(gfifoLBfullCnt[40]));
Q_MX02 U1202 ( .S(n644), .A0(gfifoLBfullCnt[41]), .A1(n1199), .Z(n757));
Q_FDP0UA U1203 ( .D(n757), .QTFCLK( ), .Q(gfifoLBfullCnt[41]));
Q_MX02 U1204 ( .S(n644), .A0(gfifoLBfullCnt[42]), .A1(n1197), .Z(n758));
Q_FDP0UA U1205 ( .D(n758), .QTFCLK( ), .Q(gfifoLBfullCnt[42]));
Q_MX02 U1206 ( .S(n644), .A0(gfifoLBfullCnt[43]), .A1(n1195), .Z(n759));
Q_FDP0UA U1207 ( .D(n759), .QTFCLK( ), .Q(gfifoLBfullCnt[43]));
Q_MX02 U1208 ( .S(n644), .A0(gfifoLBfullCnt[44]), .A1(n1193), .Z(n760));
Q_FDP0UA U1209 ( .D(n760), .QTFCLK( ), .Q(gfifoLBfullCnt[44]));
Q_MX02 U1210 ( .S(n644), .A0(gfifoLBfullCnt[45]), .A1(n1191), .Z(n761));
Q_FDP0UA U1211 ( .D(n761), .QTFCLK( ), .Q(gfifoLBfullCnt[45]));
Q_MX02 U1212 ( .S(n644), .A0(gfifoLBfullCnt[46]), .A1(n1189), .Z(n762));
Q_FDP0UA U1213 ( .D(n762), .QTFCLK( ), .Q(gfifoLBfullCnt[46]));
Q_MX02 U1214 ( .S(n644), .A0(gfifoLBfullCnt[47]), .A1(n1187), .Z(n763));
Q_FDP0UA U1215 ( .D(n763), .QTFCLK( ), .Q(gfifoLBfullCnt[47]));
Q_MX02 U1216 ( .S(n644), .A0(gfifoLBfullCnt[48]), .A1(n1185), .Z(n764));
Q_FDP0UA U1217 ( .D(n764), .QTFCLK( ), .Q(gfifoLBfullCnt[48]));
Q_MX02 U1218 ( .S(n644), .A0(gfifoLBfullCnt[49]), .A1(n1183), .Z(n765));
Q_FDP0UA U1219 ( .D(n765), .QTFCLK( ), .Q(gfifoLBfullCnt[49]));
Q_MX02 U1220 ( .S(n644), .A0(gfifoLBfullCnt[50]), .A1(n1181), .Z(n766));
Q_FDP0UA U1221 ( .D(n766), .QTFCLK( ), .Q(gfifoLBfullCnt[50]));
Q_MX02 U1222 ( .S(n644), .A0(gfifoLBfullCnt[51]), .A1(n1179), .Z(n767));
Q_FDP0UA U1223 ( .D(n767), .QTFCLK( ), .Q(gfifoLBfullCnt[51]));
Q_MX02 U1224 ( .S(n644), .A0(gfifoLBfullCnt[52]), .A1(n1177), .Z(n768));
Q_FDP0UA U1225 ( .D(n768), .QTFCLK( ), .Q(gfifoLBfullCnt[52]));
Q_MX02 U1226 ( .S(n644), .A0(gfifoLBfullCnt[53]), .A1(n1175), .Z(n769));
Q_FDP0UA U1227 ( .D(n769), .QTFCLK( ), .Q(gfifoLBfullCnt[53]));
Q_MX02 U1228 ( .S(n644), .A0(gfifoLBfullCnt[54]), .A1(n1173), .Z(n770));
Q_FDP0UA U1229 ( .D(n770), .QTFCLK( ), .Q(gfifoLBfullCnt[54]));
Q_MX02 U1230 ( .S(n644), .A0(gfifoLBfullCnt[55]), .A1(n1171), .Z(n771));
Q_FDP0UA U1231 ( .D(n771), .QTFCLK( ), .Q(gfifoLBfullCnt[55]));
Q_MX02 U1232 ( .S(n644), .A0(gfifoLBfullCnt[56]), .A1(n1169), .Z(n772));
Q_FDP0UA U1233 ( .D(n772), .QTFCLK( ), .Q(gfifoLBfullCnt[56]));
Q_MX02 U1234 ( .S(n644), .A0(gfifoLBfullCnt[57]), .A1(n1167), .Z(n773));
Q_FDP0UA U1235 ( .D(n773), .QTFCLK( ), .Q(gfifoLBfullCnt[57]));
Q_MX02 U1236 ( .S(n644), .A0(gfifoLBfullCnt[58]), .A1(n1165), .Z(n774));
Q_FDP0UA U1237 ( .D(n774), .QTFCLK( ), .Q(gfifoLBfullCnt[58]));
Q_MX02 U1238 ( .S(n644), .A0(gfifoLBfullCnt[59]), .A1(n1163), .Z(n775));
Q_FDP0UA U1239 ( .D(n775), .QTFCLK( ), .Q(gfifoLBfullCnt[59]));
Q_MX02 U1240 ( .S(n644), .A0(gfifoLBfullCnt[60]), .A1(n1161), .Z(n776));
Q_FDP0UA U1241 ( .D(n776), .QTFCLK( ), .Q(gfifoLBfullCnt[60]));
Q_MX02 U1242 ( .S(n644), .A0(gfifoLBfullCnt[61]), .A1(n1159), .Z(n777));
Q_FDP0UA U1243 ( .D(n777), .QTFCLK( ), .Q(gfifoLBfullCnt[61]));
Q_MX02 U1244 ( .S(n644), .A0(gfifoLBfullCnt[62]), .A1(n1157), .Z(n778));
Q_FDP0UA U1245 ( .D(n778), .QTFCLK( ), .Q(gfifoLBfullCnt[62]));
Q_FDP0UA U1246 ( .D(n779), .QTFCLK( ), .Q(gfifoLBfullCnt[63]));
Q_XOR2 U1247 ( .A0(n645), .A1(gfifoGBfullCnt[0]), .Z(n780));
Q_FDP0UA U1248 ( .D(n780), .QTFCLK( ), .Q(gfifoGBfullCnt[0]));
Q_MX02 U1249 ( .S(n650), .A0(n1403), .A1(gfifoGBfullCnt[1]), .Z(n781));
Q_FDP0UA U1250 ( .D(n781), .QTFCLK( ), .Q(gfifoGBfullCnt[1]));
Q_MX02 U1251 ( .S(n650), .A0(n1401), .A1(gfifoGBfullCnt[2]), .Z(n782));
Q_FDP0UA U1252 ( .D(n782), .QTFCLK( ), .Q(gfifoGBfullCnt[2]));
Q_MX02 U1253 ( .S(n650), .A0(n1399), .A1(gfifoGBfullCnt[3]), .Z(n783));
Q_FDP0UA U1254 ( .D(n783), .QTFCLK( ), .Q(gfifoGBfullCnt[3]));
Q_MX02 U1255 ( .S(n650), .A0(n1397), .A1(gfifoGBfullCnt[4]), .Z(n784));
Q_FDP0UA U1256 ( .D(n784), .QTFCLK( ), .Q(gfifoGBfullCnt[4]));
Q_MX02 U1257 ( .S(n650), .A0(n1395), .A1(gfifoGBfullCnt[5]), .Z(n785));
Q_FDP0UA U1258 ( .D(n785), .QTFCLK( ), .Q(gfifoGBfullCnt[5]));
Q_MX02 U1259 ( .S(n650), .A0(n1393), .A1(gfifoGBfullCnt[6]), .Z(n786));
Q_FDP0UA U1260 ( .D(n786), .QTFCLK( ), .Q(gfifoGBfullCnt[6]));
Q_MX02 U1261 ( .S(n650), .A0(n1391), .A1(gfifoGBfullCnt[7]), .Z(n787));
Q_FDP0UA U1262 ( .D(n787), .QTFCLK( ), .Q(gfifoGBfullCnt[7]));
Q_MX02 U1263 ( .S(n650), .A0(n1389), .A1(gfifoGBfullCnt[8]), .Z(n788));
Q_FDP0UA U1264 ( .D(n788), .QTFCLK( ), .Q(gfifoGBfullCnt[8]));
Q_MX02 U1265 ( .S(n650), .A0(n1387), .A1(gfifoGBfullCnt[9]), .Z(n789));
Q_FDP0UA U1266 ( .D(n789), .QTFCLK( ), .Q(gfifoGBfullCnt[9]));
Q_MX02 U1267 ( .S(n650), .A0(n1385), .A1(gfifoGBfullCnt[10]), .Z(n790));
Q_FDP0UA U1268 ( .D(n790), .QTFCLK( ), .Q(gfifoGBfullCnt[10]));
Q_MX02 U1269 ( .S(n650), .A0(n1383), .A1(gfifoGBfullCnt[11]), .Z(n791));
Q_FDP0UA U1270 ( .D(n791), .QTFCLK( ), .Q(gfifoGBfullCnt[11]));
Q_MX02 U1271 ( .S(n650), .A0(n1381), .A1(gfifoGBfullCnt[12]), .Z(n792));
Q_FDP0UA U1272 ( .D(n792), .QTFCLK( ), .Q(gfifoGBfullCnt[12]));
Q_MX02 U1273 ( .S(n650), .A0(n1379), .A1(gfifoGBfullCnt[13]), .Z(n793));
Q_FDP0UA U1274 ( .D(n793), .QTFCLK( ), .Q(gfifoGBfullCnt[13]));
Q_MX02 U1275 ( .S(n650), .A0(n1377), .A1(gfifoGBfullCnt[14]), .Z(n794));
Q_FDP0UA U1276 ( .D(n794), .QTFCLK( ), .Q(gfifoGBfullCnt[14]));
Q_MX02 U1277 ( .S(n650), .A0(n1375), .A1(gfifoGBfullCnt[15]), .Z(n795));
Q_FDP0UA U1278 ( .D(n795), .QTFCLK( ), .Q(gfifoGBfullCnt[15]));
Q_MX02 U1279 ( .S(n650), .A0(n1373), .A1(gfifoGBfullCnt[16]), .Z(n796));
Q_FDP0UA U1280 ( .D(n796), .QTFCLK( ), .Q(gfifoGBfullCnt[16]));
Q_MX02 U1281 ( .S(n650), .A0(n1371), .A1(gfifoGBfullCnt[17]), .Z(n797));
Q_FDP0UA U1282 ( .D(n797), .QTFCLK( ), .Q(gfifoGBfullCnt[17]));
Q_MX02 U1283 ( .S(n650), .A0(n1369), .A1(gfifoGBfullCnt[18]), .Z(n798));
Q_FDP0UA U1284 ( .D(n798), .QTFCLK( ), .Q(gfifoGBfullCnt[18]));
Q_MX02 U1285 ( .S(n650), .A0(n1367), .A1(gfifoGBfullCnt[19]), .Z(n799));
Q_FDP0UA U1286 ( .D(n799), .QTFCLK( ), .Q(gfifoGBfullCnt[19]));
Q_MX02 U1287 ( .S(n650), .A0(n1365), .A1(gfifoGBfullCnt[20]), .Z(n800));
Q_FDP0UA U1288 ( .D(n800), .QTFCLK( ), .Q(gfifoGBfullCnt[20]));
Q_MX02 U1289 ( .S(n650), .A0(n1363), .A1(gfifoGBfullCnt[21]), .Z(n801));
Q_FDP0UA U1290 ( .D(n801), .QTFCLK( ), .Q(gfifoGBfullCnt[21]));
Q_MX02 U1291 ( .S(n650), .A0(n1361), .A1(gfifoGBfullCnt[22]), .Z(n802));
Q_FDP0UA U1292 ( .D(n802), .QTFCLK( ), .Q(gfifoGBfullCnt[22]));
Q_MX02 U1293 ( .S(n650), .A0(n1359), .A1(gfifoGBfullCnt[23]), .Z(n803));
Q_FDP0UA U1294 ( .D(n803), .QTFCLK( ), .Q(gfifoGBfullCnt[23]));
Q_MX02 U1295 ( .S(n650), .A0(n1357), .A1(gfifoGBfullCnt[24]), .Z(n804));
Q_FDP0UA U1296 ( .D(n804), .QTFCLK( ), .Q(gfifoGBfullCnt[24]));
Q_MX02 U1297 ( .S(n650), .A0(n1355), .A1(gfifoGBfullCnt[25]), .Z(n805));
Q_FDP0UA U1298 ( .D(n805), .QTFCLK( ), .Q(gfifoGBfullCnt[25]));
Q_MX02 U1299 ( .S(n650), .A0(n1353), .A1(gfifoGBfullCnt[26]), .Z(n806));
Q_FDP0UA U1300 ( .D(n806), .QTFCLK( ), .Q(gfifoGBfullCnt[26]));
Q_MX02 U1301 ( .S(n650), .A0(n1351), .A1(gfifoGBfullCnt[27]), .Z(n807));
Q_FDP0UA U1302 ( .D(n807), .QTFCLK( ), .Q(gfifoGBfullCnt[27]));
Q_MX02 U1303 ( .S(n650), .A0(n1349), .A1(gfifoGBfullCnt[28]), .Z(n808));
Q_FDP0UA U1304 ( .D(n808), .QTFCLK( ), .Q(gfifoGBfullCnt[28]));
Q_MX02 U1305 ( .S(n650), .A0(n1347), .A1(gfifoGBfullCnt[29]), .Z(n809));
Q_FDP0UA U1306 ( .D(n809), .QTFCLK( ), .Q(gfifoGBfullCnt[29]));
Q_MX02 U1307 ( .S(n650), .A0(n1345), .A1(gfifoGBfullCnt[30]), .Z(n810));
Q_FDP0UA U1308 ( .D(n810), .QTFCLK( ), .Q(gfifoGBfullCnt[30]));
Q_MX02 U1309 ( .S(n650), .A0(n1343), .A1(gfifoGBfullCnt[31]), .Z(n811));
Q_FDP0UA U1310 ( .D(n811), .QTFCLK( ), .Q(gfifoGBfullCnt[31]));
Q_MX02 U1311 ( .S(n650), .A0(n1341), .A1(gfifoGBfullCnt[32]), .Z(n812));
Q_FDP0UA U1312 ( .D(n812), .QTFCLK( ), .Q(gfifoGBfullCnt[32]));
Q_MX02 U1313 ( .S(n650), .A0(n1339), .A1(gfifoGBfullCnt[33]), .Z(n813));
Q_FDP0UA U1314 ( .D(n813), .QTFCLK( ), .Q(gfifoGBfullCnt[33]));
Q_MX02 U1315 ( .S(n650), .A0(n1337), .A1(gfifoGBfullCnt[34]), .Z(n814));
Q_FDP0UA U1316 ( .D(n814), .QTFCLK( ), .Q(gfifoGBfullCnt[34]));
Q_MX02 U1317 ( .S(n650), .A0(n1335), .A1(gfifoGBfullCnt[35]), .Z(n815));
Q_FDP0UA U1318 ( .D(n815), .QTFCLK( ), .Q(gfifoGBfullCnt[35]));
Q_MX02 U1319 ( .S(n650), .A0(n1333), .A1(gfifoGBfullCnt[36]), .Z(n816));
Q_FDP0UA U1320 ( .D(n816), .QTFCLK( ), .Q(gfifoGBfullCnt[36]));
Q_MX02 U1321 ( .S(n650), .A0(n1331), .A1(gfifoGBfullCnt[37]), .Z(n817));
Q_FDP0UA U1322 ( .D(n817), .QTFCLK( ), .Q(gfifoGBfullCnt[37]));
Q_MX02 U1323 ( .S(n650), .A0(n1329), .A1(gfifoGBfullCnt[38]), .Z(n818));
Q_FDP0UA U1324 ( .D(n818), .QTFCLK( ), .Q(gfifoGBfullCnt[38]));
Q_MX02 U1325 ( .S(n650), .A0(n1327), .A1(gfifoGBfullCnt[39]), .Z(n819));
Q_FDP0UA U1326 ( .D(n819), .QTFCLK( ), .Q(gfifoGBfullCnt[39]));
Q_MX02 U1327 ( .S(n650), .A0(n1325), .A1(gfifoGBfullCnt[40]), .Z(n820));
Q_FDP0UA U1328 ( .D(n820), .QTFCLK( ), .Q(gfifoGBfullCnt[40]));
Q_MX02 U1329 ( .S(n650), .A0(n1323), .A1(gfifoGBfullCnt[41]), .Z(n821));
Q_FDP0UA U1330 ( .D(n821), .QTFCLK( ), .Q(gfifoGBfullCnt[41]));
Q_MX02 U1331 ( .S(n650), .A0(n1321), .A1(gfifoGBfullCnt[42]), .Z(n822));
Q_FDP0UA U1332 ( .D(n822), .QTFCLK( ), .Q(gfifoGBfullCnt[42]));
Q_MX02 U1333 ( .S(n650), .A0(n1319), .A1(gfifoGBfullCnt[43]), .Z(n823));
Q_FDP0UA U1334 ( .D(n823), .QTFCLK( ), .Q(gfifoGBfullCnt[43]));
Q_MX02 U1335 ( .S(n650), .A0(n1317), .A1(gfifoGBfullCnt[44]), .Z(n824));
Q_FDP0UA U1336 ( .D(n824), .QTFCLK( ), .Q(gfifoGBfullCnt[44]));
Q_MX02 U1337 ( .S(n650), .A0(n1315), .A1(gfifoGBfullCnt[45]), .Z(n825));
Q_FDP0UA U1338 ( .D(n825), .QTFCLK( ), .Q(gfifoGBfullCnt[45]));
Q_MX02 U1339 ( .S(n650), .A0(n1313), .A1(gfifoGBfullCnt[46]), .Z(n826));
Q_FDP0UA U1340 ( .D(n826), .QTFCLK( ), .Q(gfifoGBfullCnt[46]));
Q_MX02 U1341 ( .S(n650), .A0(n1311), .A1(gfifoGBfullCnt[47]), .Z(n827));
Q_FDP0UA U1342 ( .D(n827), .QTFCLK( ), .Q(gfifoGBfullCnt[47]));
Q_MX02 U1343 ( .S(n650), .A0(n1309), .A1(gfifoGBfullCnt[48]), .Z(n828));
Q_FDP0UA U1344 ( .D(n828), .QTFCLK( ), .Q(gfifoGBfullCnt[48]));
Q_MX02 U1345 ( .S(n650), .A0(n1307), .A1(gfifoGBfullCnt[49]), .Z(n829));
Q_FDP0UA U1346 ( .D(n829), .QTFCLK( ), .Q(gfifoGBfullCnt[49]));
Q_MX02 U1347 ( .S(n650), .A0(n1305), .A1(gfifoGBfullCnt[50]), .Z(n830));
Q_FDP0UA U1348 ( .D(n830), .QTFCLK( ), .Q(gfifoGBfullCnt[50]));
Q_MX02 U1349 ( .S(n650), .A0(n1303), .A1(gfifoGBfullCnt[51]), .Z(n831));
Q_FDP0UA U1350 ( .D(n831), .QTFCLK( ), .Q(gfifoGBfullCnt[51]));
Q_MX02 U1351 ( .S(n650), .A0(n1301), .A1(gfifoGBfullCnt[52]), .Z(n832));
Q_FDP0UA U1352 ( .D(n832), .QTFCLK( ), .Q(gfifoGBfullCnt[52]));
Q_MX02 U1353 ( .S(n650), .A0(n1299), .A1(gfifoGBfullCnt[53]), .Z(n833));
Q_FDP0UA U1354 ( .D(n833), .QTFCLK( ), .Q(gfifoGBfullCnt[53]));
Q_MX02 U1355 ( .S(n650), .A0(n1297), .A1(gfifoGBfullCnt[54]), .Z(n834));
Q_FDP0UA U1356 ( .D(n834), .QTFCLK( ), .Q(gfifoGBfullCnt[54]));
Q_MX02 U1357 ( .S(n650), .A0(n1295), .A1(gfifoGBfullCnt[55]), .Z(n835));
Q_FDP0UA U1358 ( .D(n835), .QTFCLK( ), .Q(gfifoGBfullCnt[55]));
Q_MX02 U1359 ( .S(n650), .A0(n1293), .A1(gfifoGBfullCnt[56]), .Z(n836));
Q_FDP0UA U1360 ( .D(n836), .QTFCLK( ), .Q(gfifoGBfullCnt[56]));
Q_MX02 U1361 ( .S(n650), .A0(n1291), .A1(gfifoGBfullCnt[57]), .Z(n837));
Q_FDP0UA U1362 ( .D(n837), .QTFCLK( ), .Q(gfifoGBfullCnt[57]));
Q_MX02 U1363 ( .S(n650), .A0(n1289), .A1(gfifoGBfullCnt[58]), .Z(n838));
Q_FDP0UA U1364 ( .D(n838), .QTFCLK( ), .Q(gfifoGBfullCnt[58]));
Q_MX02 U1365 ( .S(n650), .A0(n1287), .A1(gfifoGBfullCnt[59]), .Z(n839));
Q_FDP0UA U1366 ( .D(n839), .QTFCLK( ), .Q(gfifoGBfullCnt[59]));
Q_MX02 U1367 ( .S(n650), .A0(n1285), .A1(gfifoGBfullCnt[60]), .Z(n840));
Q_FDP0UA U1368 ( .D(n840), .QTFCLK( ), .Q(gfifoGBfullCnt[60]));
Q_MX02 U1369 ( .S(n650), .A0(n1283), .A1(gfifoGBfullCnt[61]), .Z(n841));
Q_FDP0UA U1370 ( .D(n841), .QTFCLK( ), .Q(gfifoGBfullCnt[61]));
Q_MX02 U1371 ( .S(n650), .A0(n1281), .A1(gfifoGBfullCnt[62]), .Z(n842));
Q_FDP0UA U1372 ( .D(n842), .QTFCLK( ), .Q(gfifoGBfullCnt[62]));
Q_FDP0UA U1373 ( .D(n843), .QTFCLK( ), .Q(gfifoGBfullCnt[63]));
Q_XOR2 U1374 ( .A0(n646), .A1(ixcHoldEcmCnt[0]), .Z(n844));
Q_FDP0UA U1375 ( .D(n844), .QTFCLK( ), .Q(ixcHoldEcmCnt[0]));
Q_MX02 U1376 ( .S(n651), .A0(n1031), .A1(ixcHoldEcmCnt[1]), .Z(n845));
Q_FDP0UA U1377 ( .D(n845), .QTFCLK( ), .Q(ixcHoldEcmCnt[1]));
Q_MX02 U1378 ( .S(n651), .A0(n1029), .A1(ixcHoldEcmCnt[2]), .Z(n846));
Q_FDP0UA U1379 ( .D(n846), .QTFCLK( ), .Q(ixcHoldEcmCnt[2]));
Q_MX02 U1380 ( .S(n651), .A0(n1027), .A1(ixcHoldEcmCnt[3]), .Z(n847));
Q_FDP0UA U1381 ( .D(n847), .QTFCLK( ), .Q(ixcHoldEcmCnt[3]));
Q_MX02 U1382 ( .S(n651), .A0(n1025), .A1(ixcHoldEcmCnt[4]), .Z(n848));
Q_FDP0UA U1383 ( .D(n848), .QTFCLK( ), .Q(ixcHoldEcmCnt[4]));
Q_MX02 U1384 ( .S(n651), .A0(n1023), .A1(ixcHoldEcmCnt[5]), .Z(n849));
Q_FDP0UA U1385 ( .D(n849), .QTFCLK( ), .Q(ixcHoldEcmCnt[5]));
Q_MX02 U1386 ( .S(n651), .A0(n1021), .A1(ixcHoldEcmCnt[6]), .Z(n850));
Q_FDP0UA U1387 ( .D(n850), .QTFCLK( ), .Q(ixcHoldEcmCnt[6]));
Q_MX02 U1388 ( .S(n651), .A0(n1019), .A1(ixcHoldEcmCnt[7]), .Z(n851));
Q_FDP0UA U1389 ( .D(n851), .QTFCLK( ), .Q(ixcHoldEcmCnt[7]));
Q_MX02 U1390 ( .S(n651), .A0(n1017), .A1(ixcHoldEcmCnt[8]), .Z(n852));
Q_FDP0UA U1391 ( .D(n852), .QTFCLK( ), .Q(ixcHoldEcmCnt[8]));
Q_MX02 U1392 ( .S(n651), .A0(n1015), .A1(ixcHoldEcmCnt[9]), .Z(n853));
Q_FDP0UA U1393 ( .D(n853), .QTFCLK( ), .Q(ixcHoldEcmCnt[9]));
Q_MX02 U1394 ( .S(n651), .A0(n1013), .A1(ixcHoldEcmCnt[10]), .Z(n854));
Q_FDP0UA U1395 ( .D(n854), .QTFCLK( ), .Q(ixcHoldEcmCnt[10]));
Q_MX02 U1396 ( .S(n651), .A0(n1011), .A1(ixcHoldEcmCnt[11]), .Z(n855));
Q_FDP0UA U1397 ( .D(n855), .QTFCLK( ), .Q(ixcHoldEcmCnt[11]));
Q_MX02 U1398 ( .S(n651), .A0(n1009), .A1(ixcHoldEcmCnt[12]), .Z(n856));
Q_FDP0UA U1399 ( .D(n856), .QTFCLK( ), .Q(ixcHoldEcmCnt[12]));
Q_MX02 U1400 ( .S(n651), .A0(n1007), .A1(ixcHoldEcmCnt[13]), .Z(n857));
Q_FDP0UA U1401 ( .D(n857), .QTFCLK( ), .Q(ixcHoldEcmCnt[13]));
Q_MX02 U1402 ( .S(n651), .A0(n1005), .A1(ixcHoldEcmCnt[14]), .Z(n858));
Q_FDP0UA U1403 ( .D(n858), .QTFCLK( ), .Q(ixcHoldEcmCnt[14]));
Q_MX02 U1404 ( .S(n651), .A0(n1003), .A1(ixcHoldEcmCnt[15]), .Z(n859));
Q_FDP0UA U1405 ( .D(n859), .QTFCLK( ), .Q(ixcHoldEcmCnt[15]));
Q_MX02 U1406 ( .S(n651), .A0(n1001), .A1(ixcHoldEcmCnt[16]), .Z(n860));
Q_FDP0UA U1407 ( .D(n860), .QTFCLK( ), .Q(ixcHoldEcmCnt[16]));
Q_MX02 U1408 ( .S(n651), .A0(n999), .A1(ixcHoldEcmCnt[17]), .Z(n861));
Q_FDP0UA U1409 ( .D(n861), .QTFCLK( ), .Q(ixcHoldEcmCnt[17]));
Q_MX02 U1410 ( .S(n651), .A0(n997), .A1(ixcHoldEcmCnt[18]), .Z(n862));
Q_FDP0UA U1411 ( .D(n862), .QTFCLK( ), .Q(ixcHoldEcmCnt[18]));
Q_MX02 U1412 ( .S(n651), .A0(n995), .A1(ixcHoldEcmCnt[19]), .Z(n863));
Q_FDP0UA U1413 ( .D(n863), .QTFCLK( ), .Q(ixcHoldEcmCnt[19]));
Q_MX02 U1414 ( .S(n651), .A0(n993), .A1(ixcHoldEcmCnt[20]), .Z(n864));
Q_FDP0UA U1415 ( .D(n864), .QTFCLK( ), .Q(ixcHoldEcmCnt[20]));
Q_MX02 U1416 ( .S(n651), .A0(n991), .A1(ixcHoldEcmCnt[21]), .Z(n865));
Q_FDP0UA U1417 ( .D(n865), .QTFCLK( ), .Q(ixcHoldEcmCnt[21]));
Q_MX02 U1418 ( .S(n651), .A0(n989), .A1(ixcHoldEcmCnt[22]), .Z(n866));
Q_FDP0UA U1419 ( .D(n866), .QTFCLK( ), .Q(ixcHoldEcmCnt[22]));
Q_MX02 U1420 ( .S(n651), .A0(n987), .A1(ixcHoldEcmCnt[23]), .Z(n867));
Q_FDP0UA U1421 ( .D(n867), .QTFCLK( ), .Q(ixcHoldEcmCnt[23]));
Q_MX02 U1422 ( .S(n651), .A0(n985), .A1(ixcHoldEcmCnt[24]), .Z(n868));
Q_FDP0UA U1423 ( .D(n868), .QTFCLK( ), .Q(ixcHoldEcmCnt[24]));
Q_MX02 U1424 ( .S(n651), .A0(n983), .A1(ixcHoldEcmCnt[25]), .Z(n869));
Q_FDP0UA U1425 ( .D(n869), .QTFCLK( ), .Q(ixcHoldEcmCnt[25]));
Q_MX02 U1426 ( .S(n651), .A0(n981), .A1(ixcHoldEcmCnt[26]), .Z(n870));
Q_FDP0UA U1427 ( .D(n870), .QTFCLK( ), .Q(ixcHoldEcmCnt[26]));
Q_MX02 U1428 ( .S(n651), .A0(n979), .A1(ixcHoldEcmCnt[27]), .Z(n871));
Q_FDP0UA U1429 ( .D(n871), .QTFCLK( ), .Q(ixcHoldEcmCnt[27]));
Q_MX02 U1430 ( .S(n651), .A0(n977), .A1(ixcHoldEcmCnt[28]), .Z(n872));
Q_FDP0UA U1431 ( .D(n872), .QTFCLK( ), .Q(ixcHoldEcmCnt[28]));
Q_MX02 U1432 ( .S(n651), .A0(n975), .A1(ixcHoldEcmCnt[29]), .Z(n873));
Q_FDP0UA U1433 ( .D(n873), .QTFCLK( ), .Q(ixcHoldEcmCnt[29]));
Q_MX02 U1434 ( .S(n651), .A0(n973), .A1(ixcHoldEcmCnt[30]), .Z(n874));
Q_FDP0UA U1435 ( .D(n874), .QTFCLK( ), .Q(ixcHoldEcmCnt[30]));
Q_MX02 U1436 ( .S(n651), .A0(n971), .A1(ixcHoldEcmCnt[31]), .Z(n875));
Q_FDP0UA U1437 ( .D(n875), .QTFCLK( ), .Q(ixcHoldEcmCnt[31]));
Q_MX02 U1438 ( .S(n651), .A0(n969), .A1(ixcHoldEcmCnt[32]), .Z(n876));
Q_FDP0UA U1439 ( .D(n876), .QTFCLK( ), .Q(ixcHoldEcmCnt[32]));
Q_MX02 U1440 ( .S(n651), .A0(n967), .A1(ixcHoldEcmCnt[33]), .Z(n877));
Q_FDP0UA U1441 ( .D(n877), .QTFCLK( ), .Q(ixcHoldEcmCnt[33]));
Q_MX02 U1442 ( .S(n651), .A0(n965), .A1(ixcHoldEcmCnt[34]), .Z(n878));
Q_FDP0UA U1443 ( .D(n878), .QTFCLK( ), .Q(ixcHoldEcmCnt[34]));
Q_MX02 U1444 ( .S(n651), .A0(n963), .A1(ixcHoldEcmCnt[35]), .Z(n879));
Q_FDP0UA U1445 ( .D(n879), .QTFCLK( ), .Q(ixcHoldEcmCnt[35]));
Q_MX02 U1446 ( .S(n651), .A0(n961), .A1(ixcHoldEcmCnt[36]), .Z(n880));
Q_FDP0UA U1447 ( .D(n880), .QTFCLK( ), .Q(ixcHoldEcmCnt[36]));
Q_MX02 U1448 ( .S(n651), .A0(n959), .A1(ixcHoldEcmCnt[37]), .Z(n881));
Q_FDP0UA U1449 ( .D(n881), .QTFCLK( ), .Q(ixcHoldEcmCnt[37]));
Q_MX02 U1450 ( .S(n651), .A0(n957), .A1(ixcHoldEcmCnt[38]), .Z(n882));
Q_FDP0UA U1451 ( .D(n882), .QTFCLK( ), .Q(ixcHoldEcmCnt[38]));
Q_MX02 U1452 ( .S(n651), .A0(n955), .A1(ixcHoldEcmCnt[39]), .Z(n883));
Q_FDP0UA U1453 ( .D(n883), .QTFCLK( ), .Q(ixcHoldEcmCnt[39]));
Q_MX02 U1454 ( .S(n651), .A0(n953), .A1(ixcHoldEcmCnt[40]), .Z(n884));
Q_FDP0UA U1455 ( .D(n884), .QTFCLK( ), .Q(ixcHoldEcmCnt[40]));
Q_MX02 U1456 ( .S(n651), .A0(n951), .A1(ixcHoldEcmCnt[41]), .Z(n885));
Q_FDP0UA U1457 ( .D(n885), .QTFCLK( ), .Q(ixcHoldEcmCnt[41]));
Q_MX02 U1458 ( .S(n651), .A0(n949), .A1(ixcHoldEcmCnt[42]), .Z(n886));
Q_FDP0UA U1459 ( .D(n886), .QTFCLK( ), .Q(ixcHoldEcmCnt[42]));
Q_MX02 U1460 ( .S(n651), .A0(n947), .A1(ixcHoldEcmCnt[43]), .Z(n887));
Q_FDP0UA U1461 ( .D(n887), .QTFCLK( ), .Q(ixcHoldEcmCnt[43]));
Q_MX02 U1462 ( .S(n651), .A0(n945), .A1(ixcHoldEcmCnt[44]), .Z(n888));
Q_FDP0UA U1463 ( .D(n888), .QTFCLK( ), .Q(ixcHoldEcmCnt[44]));
Q_MX02 U1464 ( .S(n651), .A0(n943), .A1(ixcHoldEcmCnt[45]), .Z(n889));
Q_FDP0UA U1465 ( .D(n889), .QTFCLK( ), .Q(ixcHoldEcmCnt[45]));
Q_MX02 U1466 ( .S(n651), .A0(n941), .A1(ixcHoldEcmCnt[46]), .Z(n890));
Q_FDP0UA U1467 ( .D(n890), .QTFCLK( ), .Q(ixcHoldEcmCnt[46]));
Q_MX02 U1468 ( .S(n651), .A0(n939), .A1(ixcHoldEcmCnt[47]), .Z(n891));
Q_FDP0UA U1469 ( .D(n891), .QTFCLK( ), .Q(ixcHoldEcmCnt[47]));
Q_MX02 U1470 ( .S(n651), .A0(n937), .A1(ixcHoldEcmCnt[48]), .Z(n892));
Q_FDP0UA U1471 ( .D(n892), .QTFCLK( ), .Q(ixcHoldEcmCnt[48]));
Q_MX02 U1472 ( .S(n651), .A0(n935), .A1(ixcHoldEcmCnt[49]), .Z(n893));
Q_FDP0UA U1473 ( .D(n893), .QTFCLK( ), .Q(ixcHoldEcmCnt[49]));
Q_MX02 U1474 ( .S(n651), .A0(n933), .A1(ixcHoldEcmCnt[50]), .Z(n894));
Q_FDP0UA U1475 ( .D(n894), .QTFCLK( ), .Q(ixcHoldEcmCnt[50]));
Q_MX02 U1476 ( .S(n651), .A0(n931), .A1(ixcHoldEcmCnt[51]), .Z(n895));
Q_FDP0UA U1477 ( .D(n895), .QTFCLK( ), .Q(ixcHoldEcmCnt[51]));
Q_MX02 U1478 ( .S(n651), .A0(n929), .A1(ixcHoldEcmCnt[52]), .Z(n896));
Q_FDP0UA U1479 ( .D(n896), .QTFCLK( ), .Q(ixcHoldEcmCnt[52]));
Q_MX02 U1480 ( .S(n651), .A0(n927), .A1(ixcHoldEcmCnt[53]), .Z(n897));
Q_FDP0UA U1481 ( .D(n897), .QTFCLK( ), .Q(ixcHoldEcmCnt[53]));
Q_MX02 U1482 ( .S(n651), .A0(n925), .A1(ixcHoldEcmCnt[54]), .Z(n898));
Q_FDP0UA U1483 ( .D(n898), .QTFCLK( ), .Q(ixcHoldEcmCnt[54]));
Q_MX02 U1484 ( .S(n651), .A0(n923), .A1(ixcHoldEcmCnt[55]), .Z(n899));
Q_FDP0UA U1485 ( .D(n899), .QTFCLK( ), .Q(ixcHoldEcmCnt[55]));
Q_MX02 U1486 ( .S(n651), .A0(n921), .A1(ixcHoldEcmCnt[56]), .Z(n900));
Q_FDP0UA U1487 ( .D(n900), .QTFCLK( ), .Q(ixcHoldEcmCnt[56]));
Q_MX02 U1488 ( .S(n651), .A0(n919), .A1(ixcHoldEcmCnt[57]), .Z(n901));
Q_FDP0UA U1489 ( .D(n901), .QTFCLK( ), .Q(ixcHoldEcmCnt[57]));
Q_MX02 U1490 ( .S(n651), .A0(n917), .A1(ixcHoldEcmCnt[58]), .Z(n902));
Q_FDP0UA U1491 ( .D(n902), .QTFCLK( ), .Q(ixcHoldEcmCnt[58]));
Q_MX02 U1492 ( .S(n651), .A0(n915), .A1(ixcHoldEcmCnt[59]), .Z(n903));
Q_FDP0UA U1493 ( .D(n903), .QTFCLK( ), .Q(ixcHoldEcmCnt[59]));
Q_MX02 U1494 ( .S(n651), .A0(n913), .A1(ixcHoldEcmCnt[60]), .Z(n904));
Q_FDP0UA U1495 ( .D(n904), .QTFCLK( ), .Q(ixcHoldEcmCnt[60]));
Q_MX02 U1496 ( .S(n651), .A0(n911), .A1(ixcHoldEcmCnt[61]), .Z(n905));
Q_FDP0UA U1497 ( .D(n905), .QTFCLK( ), .Q(ixcHoldEcmCnt[61]));
Q_MX02 U1498 ( .S(n651), .A0(n909), .A1(ixcHoldEcmCnt[62]), .Z(n906));
Q_FDP0UA U1499 ( .D(n906), .QTFCLK( ), .Q(ixcHoldEcmCnt[62]));
Q_FDP0UA U1500 ( .D(n907), .QTFCLK( ), .Q(ixcHoldEcmCnt[63]));
Q_XOR2 U1501 ( .A0(ixcHoldEcmCnt[63]), .A1(n11), .Z(n907));
Q_AD01HF U1502 ( .A0(ixcHoldEcmCnt[62]), .B0(n910), .S(n909), .CO(n908));
Q_AD01HF U1503 ( .A0(ixcHoldEcmCnt[61]), .B0(n912), .S(n911), .CO(n910));
Q_AD01HF U1504 ( .A0(ixcHoldEcmCnt[60]), .B0(n914), .S(n913), .CO(n912));
Q_AD01HF U1505 ( .A0(ixcHoldEcmCnt[59]), .B0(n916), .S(n915), .CO(n914));
Q_AD01HF U1506 ( .A0(ixcHoldEcmCnt[58]), .B0(n918), .S(n917), .CO(n916));
Q_AD01HF U1507 ( .A0(ixcHoldEcmCnt[57]), .B0(n920), .S(n919), .CO(n918));
Q_AD01HF U1508 ( .A0(ixcHoldEcmCnt[56]), .B0(n922), .S(n921), .CO(n920));
Q_AD01HF U1509 ( .A0(ixcHoldEcmCnt[55]), .B0(n924), .S(n923), .CO(n922));
Q_AD01HF U1510 ( .A0(ixcHoldEcmCnt[54]), .B0(n926), .S(n925), .CO(n924));
Q_AD01HF U1511 ( .A0(ixcHoldEcmCnt[53]), .B0(n928), .S(n927), .CO(n926));
Q_AD01HF U1512 ( .A0(ixcHoldEcmCnt[52]), .B0(n930), .S(n929), .CO(n928));
Q_AD01HF U1513 ( .A0(ixcHoldEcmCnt[51]), .B0(n932), .S(n931), .CO(n930));
Q_AD01HF U1514 ( .A0(ixcHoldEcmCnt[50]), .B0(n934), .S(n933), .CO(n932));
Q_AD01HF U1515 ( .A0(ixcHoldEcmCnt[49]), .B0(n936), .S(n935), .CO(n934));
Q_AD01HF U1516 ( .A0(ixcHoldEcmCnt[48]), .B0(n938), .S(n937), .CO(n936));
Q_AD01HF U1517 ( .A0(ixcHoldEcmCnt[47]), .B0(n940), .S(n939), .CO(n938));
Q_AD01HF U1518 ( .A0(ixcHoldEcmCnt[46]), .B0(n942), .S(n941), .CO(n940));
Q_AD01HF U1519 ( .A0(ixcHoldEcmCnt[45]), .B0(n944), .S(n943), .CO(n942));
Q_AD01HF U1520 ( .A0(ixcHoldEcmCnt[44]), .B0(n946), .S(n945), .CO(n944));
Q_AD01HF U1521 ( .A0(ixcHoldEcmCnt[43]), .B0(n948), .S(n947), .CO(n946));
Q_AD01HF U1522 ( .A0(ixcHoldEcmCnt[42]), .B0(n950), .S(n949), .CO(n948));
Q_AD01HF U1523 ( .A0(ixcHoldEcmCnt[41]), .B0(n952), .S(n951), .CO(n950));
Q_AD01HF U1524 ( .A0(ixcHoldEcmCnt[40]), .B0(n954), .S(n953), .CO(n952));
Q_AD01HF U1525 ( .A0(ixcHoldEcmCnt[39]), .B0(n956), .S(n955), .CO(n954));
Q_AD01HF U1526 ( .A0(ixcHoldEcmCnt[38]), .B0(n958), .S(n957), .CO(n956));
Q_AD01HF U1527 ( .A0(ixcHoldEcmCnt[37]), .B0(n960), .S(n959), .CO(n958));
Q_AD01HF U1528 ( .A0(ixcHoldEcmCnt[36]), .B0(n962), .S(n961), .CO(n960));
Q_AD01HF U1529 ( .A0(ixcHoldEcmCnt[35]), .B0(n964), .S(n963), .CO(n962));
Q_AD01HF U1530 ( .A0(ixcHoldEcmCnt[34]), .B0(n966), .S(n965), .CO(n964));
Q_AD01HF U1531 ( .A0(ixcHoldEcmCnt[33]), .B0(n968), .S(n967), .CO(n966));
Q_AD01HF U1532 ( .A0(ixcHoldEcmCnt[32]), .B0(n970), .S(n969), .CO(n968));
Q_AD01HF U1533 ( .A0(ixcHoldEcmCnt[31]), .B0(n972), .S(n971), .CO(n970));
Q_AD01HF U1534 ( .A0(ixcHoldEcmCnt[30]), .B0(n974), .S(n973), .CO(n972));
Q_AD01HF U1535 ( .A0(ixcHoldEcmCnt[29]), .B0(n976), .S(n975), .CO(n974));
Q_AD01HF U1536 ( .A0(ixcHoldEcmCnt[28]), .B0(n978), .S(n977), .CO(n976));
Q_AD01HF U1537 ( .A0(ixcHoldEcmCnt[27]), .B0(n980), .S(n979), .CO(n978));
Q_AD01HF U1538 ( .A0(ixcHoldEcmCnt[26]), .B0(n982), .S(n981), .CO(n980));
Q_AD01HF U1539 ( .A0(ixcHoldEcmCnt[25]), .B0(n984), .S(n983), .CO(n982));
Q_AD01HF U1540 ( .A0(ixcHoldEcmCnt[24]), .B0(n986), .S(n985), .CO(n984));
Q_AD01HF U1541 ( .A0(ixcHoldEcmCnt[23]), .B0(n988), .S(n987), .CO(n986));
Q_AD01HF U1542 ( .A0(ixcHoldEcmCnt[22]), .B0(n990), .S(n989), .CO(n988));
Q_AD01HF U1543 ( .A0(ixcHoldEcmCnt[21]), .B0(n992), .S(n991), .CO(n990));
Q_AD01HF U1544 ( .A0(ixcHoldEcmCnt[20]), .B0(n994), .S(n993), .CO(n992));
Q_AD01HF U1545 ( .A0(ixcHoldEcmCnt[19]), .B0(n996), .S(n995), .CO(n994));
Q_AD01HF U1546 ( .A0(ixcHoldEcmCnt[18]), .B0(n998), .S(n997), .CO(n996));
Q_AD01HF U1547 ( .A0(ixcHoldEcmCnt[17]), .B0(n1000), .S(n999), .CO(n998));
Q_AD01HF U1548 ( .A0(ixcHoldEcmCnt[16]), .B0(n1002), .S(n1001), .CO(n1000));
Q_AD01HF U1549 ( .A0(ixcHoldEcmCnt[15]), .B0(n1004), .S(n1003), .CO(n1002));
Q_AD01HF U1550 ( .A0(ixcHoldEcmCnt[14]), .B0(n1006), .S(n1005), .CO(n1004));
Q_AD01HF U1551 ( .A0(ixcHoldEcmCnt[13]), .B0(n1008), .S(n1007), .CO(n1006));
Q_AD01HF U1552 ( .A0(ixcHoldEcmCnt[12]), .B0(n1010), .S(n1009), .CO(n1008));
Q_AD01HF U1553 ( .A0(ixcHoldEcmCnt[11]), .B0(n1012), .S(n1011), .CO(n1010));
Q_AD01HF U1554 ( .A0(ixcHoldEcmCnt[10]), .B0(n1014), .S(n1013), .CO(n1012));
Q_AD01HF U1555 ( .A0(ixcHoldEcmCnt[9]), .B0(n1016), .S(n1015), .CO(n1014));
Q_AD01HF U1556 ( .A0(ixcHoldEcmCnt[8]), .B0(n1018), .S(n1017), .CO(n1016));
Q_AD01HF U1557 ( .A0(ixcHoldEcmCnt[7]), .B0(n1020), .S(n1019), .CO(n1018));
Q_AD01HF U1558 ( .A0(ixcHoldEcmCnt[6]), .B0(n1022), .S(n1021), .CO(n1020));
Q_AD01HF U1559 ( .A0(ixcHoldEcmCnt[5]), .B0(n1024), .S(n1023), .CO(n1022));
Q_AD01HF U1560 ( .A0(ixcHoldEcmCnt[4]), .B0(n1026), .S(n1025), .CO(n1024));
Q_AD01HF U1561 ( .A0(ixcHoldEcmCnt[3]), .B0(n1028), .S(n1027), .CO(n1026));
Q_AD01HF U1562 ( .A0(ixcHoldEcmCnt[2]), .B0(n1030), .S(n1029), .CO(n1028));
Q_AD01HF U1563 ( .A0(ixcHoldEcmCnt[1]), .B0(ixcHoldEcmCnt[0]), .S(n1031), .CO(n1030));
Q_XOR2 U1564 ( .A0(gfifoTBsyncCnt[63]), .A1(n14), .Z(n715));
Q_AD01HF U1565 ( .A0(gfifoTBsyncCnt[62]), .B0(n1034), .S(n1033), .CO(n1032));
Q_AD01HF U1566 ( .A0(gfifoTBsyncCnt[61]), .B0(n1036), .S(n1035), .CO(n1034));
Q_AD01HF U1567 ( .A0(gfifoTBsyncCnt[60]), .B0(n1038), .S(n1037), .CO(n1036));
Q_AD01HF U1568 ( .A0(gfifoTBsyncCnt[59]), .B0(n1040), .S(n1039), .CO(n1038));
Q_AD01HF U1569 ( .A0(gfifoTBsyncCnt[58]), .B0(n1042), .S(n1041), .CO(n1040));
Q_AD01HF U1570 ( .A0(gfifoTBsyncCnt[57]), .B0(n1044), .S(n1043), .CO(n1042));
Q_AD01HF U1571 ( .A0(gfifoTBsyncCnt[56]), .B0(n1046), .S(n1045), .CO(n1044));
Q_AD01HF U1572 ( .A0(gfifoTBsyncCnt[55]), .B0(n1048), .S(n1047), .CO(n1046));
Q_AD01HF U1573 ( .A0(gfifoTBsyncCnt[54]), .B0(n1050), .S(n1049), .CO(n1048));
Q_AD01HF U1574 ( .A0(gfifoTBsyncCnt[53]), .B0(n1052), .S(n1051), .CO(n1050));
Q_AD01HF U1575 ( .A0(gfifoTBsyncCnt[52]), .B0(n1054), .S(n1053), .CO(n1052));
Q_AD01HF U1576 ( .A0(gfifoTBsyncCnt[51]), .B0(n1056), .S(n1055), .CO(n1054));
Q_AD01HF U1577 ( .A0(gfifoTBsyncCnt[50]), .B0(n1058), .S(n1057), .CO(n1056));
Q_AD01HF U1578 ( .A0(gfifoTBsyncCnt[49]), .B0(n1060), .S(n1059), .CO(n1058));
Q_AD01HF U1579 ( .A0(gfifoTBsyncCnt[48]), .B0(n1062), .S(n1061), .CO(n1060));
Q_AD01HF U1580 ( .A0(gfifoTBsyncCnt[47]), .B0(n1064), .S(n1063), .CO(n1062));
Q_AD01HF U1581 ( .A0(gfifoTBsyncCnt[46]), .B0(n1066), .S(n1065), .CO(n1064));
Q_AD01HF U1582 ( .A0(gfifoTBsyncCnt[45]), .B0(n1068), .S(n1067), .CO(n1066));
Q_AD01HF U1583 ( .A0(gfifoTBsyncCnt[44]), .B0(n1070), .S(n1069), .CO(n1068));
Q_AD01HF U1584 ( .A0(gfifoTBsyncCnt[43]), .B0(n1072), .S(n1071), .CO(n1070));
Q_AD01HF U1585 ( .A0(gfifoTBsyncCnt[42]), .B0(n1074), .S(n1073), .CO(n1072));
Q_AD01HF U1586 ( .A0(gfifoTBsyncCnt[41]), .B0(n1076), .S(n1075), .CO(n1074));
Q_AD01HF U1587 ( .A0(gfifoTBsyncCnt[40]), .B0(n1078), .S(n1077), .CO(n1076));
Q_AD01HF U1588 ( .A0(gfifoTBsyncCnt[39]), .B0(n1080), .S(n1079), .CO(n1078));
Q_AD01HF U1589 ( .A0(gfifoTBsyncCnt[38]), .B0(n1082), .S(n1081), .CO(n1080));
Q_AD01HF U1590 ( .A0(gfifoTBsyncCnt[37]), .B0(n1084), .S(n1083), .CO(n1082));
Q_AD01HF U1591 ( .A0(gfifoTBsyncCnt[36]), .B0(n1086), .S(n1085), .CO(n1084));
Q_AD01HF U1592 ( .A0(gfifoTBsyncCnt[35]), .B0(n1088), .S(n1087), .CO(n1086));
Q_AD01HF U1593 ( .A0(gfifoTBsyncCnt[34]), .B0(n1090), .S(n1089), .CO(n1088));
Q_AD01HF U1594 ( .A0(gfifoTBsyncCnt[33]), .B0(n1092), .S(n1091), .CO(n1090));
Q_AD01HF U1595 ( .A0(gfifoTBsyncCnt[32]), .B0(n1094), .S(n1093), .CO(n1092));
Q_AD01HF U1596 ( .A0(gfifoTBsyncCnt[31]), .B0(n1096), .S(n1095), .CO(n1094));
Q_AD01HF U1597 ( .A0(gfifoTBsyncCnt[30]), .B0(n1098), .S(n1097), .CO(n1096));
Q_AD01HF U1598 ( .A0(gfifoTBsyncCnt[29]), .B0(n1100), .S(n1099), .CO(n1098));
Q_AD01HF U1599 ( .A0(gfifoTBsyncCnt[28]), .B0(n1102), .S(n1101), .CO(n1100));
Q_AD01HF U1600 ( .A0(gfifoTBsyncCnt[27]), .B0(n1104), .S(n1103), .CO(n1102));
Q_AD01HF U1601 ( .A0(gfifoTBsyncCnt[26]), .B0(n1106), .S(n1105), .CO(n1104));
Q_AD01HF U1602 ( .A0(gfifoTBsyncCnt[25]), .B0(n1108), .S(n1107), .CO(n1106));
Q_AD01HF U1603 ( .A0(gfifoTBsyncCnt[24]), .B0(n1110), .S(n1109), .CO(n1108));
Q_AD01HF U1604 ( .A0(gfifoTBsyncCnt[23]), .B0(n1112), .S(n1111), .CO(n1110));
Q_AD01HF U1605 ( .A0(gfifoTBsyncCnt[22]), .B0(n1114), .S(n1113), .CO(n1112));
Q_AD01HF U1606 ( .A0(gfifoTBsyncCnt[21]), .B0(n1116), .S(n1115), .CO(n1114));
Q_AD01HF U1607 ( .A0(gfifoTBsyncCnt[20]), .B0(n1118), .S(n1117), .CO(n1116));
Q_AD01HF U1608 ( .A0(gfifoTBsyncCnt[19]), .B0(n1120), .S(n1119), .CO(n1118));
Q_AD01HF U1609 ( .A0(gfifoTBsyncCnt[18]), .B0(n1122), .S(n1121), .CO(n1120));
Q_AD01HF U1610 ( .A0(gfifoTBsyncCnt[17]), .B0(n1124), .S(n1123), .CO(n1122));
Q_AD01HF U1611 ( .A0(gfifoTBsyncCnt[16]), .B0(n1126), .S(n1125), .CO(n1124));
Q_AD01HF U1612 ( .A0(gfifoTBsyncCnt[15]), .B0(n1128), .S(n1127), .CO(n1126));
Q_AD01HF U1613 ( .A0(gfifoTBsyncCnt[14]), .B0(n1130), .S(n1129), .CO(n1128));
Q_AD01HF U1614 ( .A0(gfifoTBsyncCnt[13]), .B0(n1132), .S(n1131), .CO(n1130));
Q_AD01HF U1615 ( .A0(gfifoTBsyncCnt[12]), .B0(n1134), .S(n1133), .CO(n1132));
Q_AD01HF U1616 ( .A0(gfifoTBsyncCnt[11]), .B0(n1136), .S(n1135), .CO(n1134));
Q_AD01HF U1617 ( .A0(gfifoTBsyncCnt[10]), .B0(n1138), .S(n1137), .CO(n1136));
Q_AD01HF U1618 ( .A0(gfifoTBsyncCnt[9]), .B0(n1140), .S(n1139), .CO(n1138));
Q_AD01HF U1619 ( .A0(gfifoTBsyncCnt[8]), .B0(n1142), .S(n1141), .CO(n1140));
Q_AD01HF U1620 ( .A0(gfifoTBsyncCnt[7]), .B0(n1144), .S(n1143), .CO(n1142));
Q_AD01HF U1621 ( .A0(gfifoTBsyncCnt[6]), .B0(n1146), .S(n1145), .CO(n1144));
Q_AD01HF U1622 ( .A0(gfifoTBsyncCnt[5]), .B0(n1148), .S(n1147), .CO(n1146));
Q_AD01HF U1623 ( .A0(gfifoTBsyncCnt[4]), .B0(n1150), .S(n1149), .CO(n1148));
Q_AD01HF U1624 ( .A0(gfifoTBsyncCnt[3]), .B0(n1152), .S(n1151), .CO(n1150));
Q_AD01HF U1625 ( .A0(gfifoTBsyncCnt[2]), .B0(n1154), .S(n1153), .CO(n1152));
Q_AD01HF U1626 ( .A0(gfifoTBsyncCnt[1]), .B0(gfifoTBsyncCnt[0]), .S(n1155), .CO(n1154));
Q_XOR2 U1627 ( .A0(gfifoLBfullCnt[63]), .A1(n13), .Z(n779));
Q_AD01HF U1628 ( .A0(gfifoLBfullCnt[62]), .B0(n1158), .S(n1157), .CO(n1156));
Q_AD01HF U1629 ( .A0(gfifoLBfullCnt[61]), .B0(n1160), .S(n1159), .CO(n1158));
Q_AD01HF U1630 ( .A0(gfifoLBfullCnt[60]), .B0(n1162), .S(n1161), .CO(n1160));
Q_AD01HF U1631 ( .A0(gfifoLBfullCnt[59]), .B0(n1164), .S(n1163), .CO(n1162));
Q_AD01HF U1632 ( .A0(gfifoLBfullCnt[58]), .B0(n1166), .S(n1165), .CO(n1164));
Q_AD01HF U1633 ( .A0(gfifoLBfullCnt[57]), .B0(n1168), .S(n1167), .CO(n1166));
Q_AD01HF U1634 ( .A0(gfifoLBfullCnt[56]), .B0(n1170), .S(n1169), .CO(n1168));
Q_AD01HF U1635 ( .A0(gfifoLBfullCnt[55]), .B0(n1172), .S(n1171), .CO(n1170));
Q_AD01HF U1636 ( .A0(gfifoLBfullCnt[54]), .B0(n1174), .S(n1173), .CO(n1172));
Q_AD01HF U1637 ( .A0(gfifoLBfullCnt[53]), .B0(n1176), .S(n1175), .CO(n1174));
Q_AD01HF U1638 ( .A0(gfifoLBfullCnt[52]), .B0(n1178), .S(n1177), .CO(n1176));
Q_AD01HF U1639 ( .A0(gfifoLBfullCnt[51]), .B0(n1180), .S(n1179), .CO(n1178));
Q_AD01HF U1640 ( .A0(gfifoLBfullCnt[50]), .B0(n1182), .S(n1181), .CO(n1180));
Q_AD01HF U1641 ( .A0(gfifoLBfullCnt[49]), .B0(n1184), .S(n1183), .CO(n1182));
Q_AD01HF U1642 ( .A0(gfifoLBfullCnt[48]), .B0(n1186), .S(n1185), .CO(n1184));
Q_AD01HF U1643 ( .A0(gfifoLBfullCnt[47]), .B0(n1188), .S(n1187), .CO(n1186));
Q_AD01HF U1644 ( .A0(gfifoLBfullCnt[46]), .B0(n1190), .S(n1189), .CO(n1188));
Q_AD01HF U1645 ( .A0(gfifoLBfullCnt[45]), .B0(n1192), .S(n1191), .CO(n1190));
Q_AD01HF U1646 ( .A0(gfifoLBfullCnt[44]), .B0(n1194), .S(n1193), .CO(n1192));
Q_AD01HF U1647 ( .A0(gfifoLBfullCnt[43]), .B0(n1196), .S(n1195), .CO(n1194));
Q_AD01HF U1648 ( .A0(gfifoLBfullCnt[42]), .B0(n1198), .S(n1197), .CO(n1196));
Q_AD01HF U1649 ( .A0(gfifoLBfullCnt[41]), .B0(n1200), .S(n1199), .CO(n1198));
Q_AD01HF U1650 ( .A0(gfifoLBfullCnt[40]), .B0(n1202), .S(n1201), .CO(n1200));
Q_AD01HF U1651 ( .A0(gfifoLBfullCnt[39]), .B0(n1204), .S(n1203), .CO(n1202));
Q_AD01HF U1652 ( .A0(gfifoLBfullCnt[38]), .B0(n1206), .S(n1205), .CO(n1204));
Q_AD01HF U1653 ( .A0(gfifoLBfullCnt[37]), .B0(n1208), .S(n1207), .CO(n1206));
Q_AD01HF U1654 ( .A0(gfifoLBfullCnt[36]), .B0(n1210), .S(n1209), .CO(n1208));
Q_AD01HF U1655 ( .A0(gfifoLBfullCnt[35]), .B0(n1212), .S(n1211), .CO(n1210));
Q_AD01HF U1656 ( .A0(gfifoLBfullCnt[34]), .B0(n1214), .S(n1213), .CO(n1212));
Q_AD01HF U1657 ( .A0(gfifoLBfullCnt[33]), .B0(n1216), .S(n1215), .CO(n1214));
Q_AD01HF U1658 ( .A0(gfifoLBfullCnt[32]), .B0(n1218), .S(n1217), .CO(n1216));
Q_AD01HF U1659 ( .A0(gfifoLBfullCnt[31]), .B0(n1220), .S(n1219), .CO(n1218));
Q_AD01HF U1660 ( .A0(gfifoLBfullCnt[30]), .B0(n1222), .S(n1221), .CO(n1220));
Q_AD01HF U1661 ( .A0(gfifoLBfullCnt[29]), .B0(n1224), .S(n1223), .CO(n1222));
Q_AD01HF U1662 ( .A0(gfifoLBfullCnt[28]), .B0(n1226), .S(n1225), .CO(n1224));
Q_AD01HF U1663 ( .A0(gfifoLBfullCnt[27]), .B0(n1228), .S(n1227), .CO(n1226));
Q_AD01HF U1664 ( .A0(gfifoLBfullCnt[26]), .B0(n1230), .S(n1229), .CO(n1228));
Q_AD01HF U1665 ( .A0(gfifoLBfullCnt[25]), .B0(n1232), .S(n1231), .CO(n1230));
Q_AD01HF U1666 ( .A0(gfifoLBfullCnt[24]), .B0(n1234), .S(n1233), .CO(n1232));
Q_AD01HF U1667 ( .A0(gfifoLBfullCnt[23]), .B0(n1236), .S(n1235), .CO(n1234));
Q_AD01HF U1668 ( .A0(gfifoLBfullCnt[22]), .B0(n1238), .S(n1237), .CO(n1236));
Q_AD01HF U1669 ( .A0(gfifoLBfullCnt[21]), .B0(n1240), .S(n1239), .CO(n1238));
Q_AD01HF U1670 ( .A0(gfifoLBfullCnt[20]), .B0(n1242), .S(n1241), .CO(n1240));
Q_AD01HF U1671 ( .A0(gfifoLBfullCnt[19]), .B0(n1244), .S(n1243), .CO(n1242));
Q_AD01HF U1672 ( .A0(gfifoLBfullCnt[18]), .B0(n1246), .S(n1245), .CO(n1244));
Q_AD01HF U1673 ( .A0(gfifoLBfullCnt[17]), .B0(n1248), .S(n1247), .CO(n1246));
Q_AD01HF U1674 ( .A0(gfifoLBfullCnt[16]), .B0(n1250), .S(n1249), .CO(n1248));
Q_AD01HF U1675 ( .A0(gfifoLBfullCnt[15]), .B0(n1252), .S(n1251), .CO(n1250));
Q_AD01HF U1676 ( .A0(gfifoLBfullCnt[14]), .B0(n1254), .S(n1253), .CO(n1252));
Q_AD01HF U1677 ( .A0(gfifoLBfullCnt[13]), .B0(n1256), .S(n1255), .CO(n1254));
Q_AD01HF U1678 ( .A0(gfifoLBfullCnt[12]), .B0(n1258), .S(n1257), .CO(n1256));
Q_AD01HF U1679 ( .A0(gfifoLBfullCnt[11]), .B0(n1260), .S(n1259), .CO(n1258));
Q_AD01HF U1680 ( .A0(gfifoLBfullCnt[10]), .B0(n1262), .S(n1261), .CO(n1260));
Q_AD01HF U1681 ( .A0(gfifoLBfullCnt[9]), .B0(n1264), .S(n1263), .CO(n1262));
Q_AD01HF U1682 ( .A0(gfifoLBfullCnt[8]), .B0(n1266), .S(n1265), .CO(n1264));
Q_AD01HF U1683 ( .A0(gfifoLBfullCnt[7]), .B0(n1268), .S(n1267), .CO(n1266));
Q_AD01HF U1684 ( .A0(gfifoLBfullCnt[6]), .B0(n1270), .S(n1269), .CO(n1268));
Q_AD01HF U1685 ( .A0(gfifoLBfullCnt[5]), .B0(n1272), .S(n1271), .CO(n1270));
Q_AD01HF U1686 ( .A0(gfifoLBfullCnt[4]), .B0(n1274), .S(n1273), .CO(n1272));
Q_AD01HF U1687 ( .A0(gfifoLBfullCnt[3]), .B0(n1276), .S(n1275), .CO(n1274));
Q_AD01HF U1688 ( .A0(gfifoLBfullCnt[2]), .B0(n1278), .S(n1277), .CO(n1276));
Q_AD01HF U1689 ( .A0(gfifoLBfullCnt[1]), .B0(gfifoLBfullCnt[0]), .S(n1279), .CO(n1278));
Q_XOR2 U1690 ( .A0(gfifoGBfullCnt[63]), .A1(n12), .Z(n843));
Q_AD01HF U1691 ( .A0(gfifoGBfullCnt[62]), .B0(n1282), .S(n1281), .CO(n1280));
Q_AD01HF U1692 ( .A0(gfifoGBfullCnt[61]), .B0(n1284), .S(n1283), .CO(n1282));
Q_AD01HF U1693 ( .A0(gfifoGBfullCnt[60]), .B0(n1286), .S(n1285), .CO(n1284));
Q_AD01HF U1694 ( .A0(gfifoGBfullCnt[59]), .B0(n1288), .S(n1287), .CO(n1286));
Q_AD01HF U1695 ( .A0(gfifoGBfullCnt[58]), .B0(n1290), .S(n1289), .CO(n1288));
Q_AD01HF U1696 ( .A0(gfifoGBfullCnt[57]), .B0(n1292), .S(n1291), .CO(n1290));
Q_AD01HF U1697 ( .A0(gfifoGBfullCnt[56]), .B0(n1294), .S(n1293), .CO(n1292));
Q_AD01HF U1698 ( .A0(gfifoGBfullCnt[55]), .B0(n1296), .S(n1295), .CO(n1294));
Q_AD01HF U1699 ( .A0(gfifoGBfullCnt[54]), .B0(n1298), .S(n1297), .CO(n1296));
Q_AD01HF U1700 ( .A0(gfifoGBfullCnt[53]), .B0(n1300), .S(n1299), .CO(n1298));
Q_AD01HF U1701 ( .A0(gfifoGBfullCnt[52]), .B0(n1302), .S(n1301), .CO(n1300));
Q_AD01HF U1702 ( .A0(gfifoGBfullCnt[51]), .B0(n1304), .S(n1303), .CO(n1302));
Q_AD01HF U1703 ( .A0(gfifoGBfullCnt[50]), .B0(n1306), .S(n1305), .CO(n1304));
Q_AD01HF U1704 ( .A0(gfifoGBfullCnt[49]), .B0(n1308), .S(n1307), .CO(n1306));
Q_AD01HF U1705 ( .A0(gfifoGBfullCnt[48]), .B0(n1310), .S(n1309), .CO(n1308));
Q_AD01HF U1706 ( .A0(gfifoGBfullCnt[47]), .B0(n1312), .S(n1311), .CO(n1310));
Q_AD01HF U1707 ( .A0(gfifoGBfullCnt[46]), .B0(n1314), .S(n1313), .CO(n1312));
Q_AD01HF U1708 ( .A0(gfifoGBfullCnt[45]), .B0(n1316), .S(n1315), .CO(n1314));
Q_AD01HF U1709 ( .A0(gfifoGBfullCnt[44]), .B0(n1318), .S(n1317), .CO(n1316));
Q_AD01HF U1710 ( .A0(gfifoGBfullCnt[43]), .B0(n1320), .S(n1319), .CO(n1318));
Q_AD01HF U1711 ( .A0(gfifoGBfullCnt[42]), .B0(n1322), .S(n1321), .CO(n1320));
Q_AD01HF U1712 ( .A0(gfifoGBfullCnt[41]), .B0(n1324), .S(n1323), .CO(n1322));
Q_AD01HF U1713 ( .A0(gfifoGBfullCnt[40]), .B0(n1326), .S(n1325), .CO(n1324));
Q_AD01HF U1714 ( .A0(gfifoGBfullCnt[39]), .B0(n1328), .S(n1327), .CO(n1326));
Q_AD01HF U1715 ( .A0(gfifoGBfullCnt[38]), .B0(n1330), .S(n1329), .CO(n1328));
Q_AD01HF U1716 ( .A0(gfifoGBfullCnt[37]), .B0(n1332), .S(n1331), .CO(n1330));
Q_AD01HF U1717 ( .A0(gfifoGBfullCnt[36]), .B0(n1334), .S(n1333), .CO(n1332));
Q_AD01HF U1718 ( .A0(gfifoGBfullCnt[35]), .B0(n1336), .S(n1335), .CO(n1334));
Q_AD01HF U1719 ( .A0(gfifoGBfullCnt[34]), .B0(n1338), .S(n1337), .CO(n1336));
Q_AD01HF U1720 ( .A0(gfifoGBfullCnt[33]), .B0(n1340), .S(n1339), .CO(n1338));
Q_AD01HF U1721 ( .A0(gfifoGBfullCnt[32]), .B0(n1342), .S(n1341), .CO(n1340));
Q_AD01HF U1722 ( .A0(gfifoGBfullCnt[31]), .B0(n1344), .S(n1343), .CO(n1342));
Q_AD01HF U1723 ( .A0(gfifoGBfullCnt[30]), .B0(n1346), .S(n1345), .CO(n1344));
Q_AD01HF U1724 ( .A0(gfifoGBfullCnt[29]), .B0(n1348), .S(n1347), .CO(n1346));
Q_AD01HF U1725 ( .A0(gfifoGBfullCnt[28]), .B0(n1350), .S(n1349), .CO(n1348));
Q_AD01HF U1726 ( .A0(gfifoGBfullCnt[27]), .B0(n1352), .S(n1351), .CO(n1350));
Q_AD01HF U1727 ( .A0(gfifoGBfullCnt[26]), .B0(n1354), .S(n1353), .CO(n1352));
Q_AD01HF U1728 ( .A0(gfifoGBfullCnt[25]), .B0(n1356), .S(n1355), .CO(n1354));
Q_AD01HF U1729 ( .A0(gfifoGBfullCnt[24]), .B0(n1358), .S(n1357), .CO(n1356));
Q_AD01HF U1730 ( .A0(gfifoGBfullCnt[23]), .B0(n1360), .S(n1359), .CO(n1358));
Q_AD01HF U1731 ( .A0(gfifoGBfullCnt[22]), .B0(n1362), .S(n1361), .CO(n1360));
Q_AD01HF U1732 ( .A0(gfifoGBfullCnt[21]), .B0(n1364), .S(n1363), .CO(n1362));
Q_AD01HF U1733 ( .A0(gfifoGBfullCnt[20]), .B0(n1366), .S(n1365), .CO(n1364));
Q_AD01HF U1734 ( .A0(gfifoGBfullCnt[19]), .B0(n1368), .S(n1367), .CO(n1366));
Q_AD01HF U1735 ( .A0(gfifoGBfullCnt[18]), .B0(n1370), .S(n1369), .CO(n1368));
Q_AD01HF U1736 ( .A0(gfifoGBfullCnt[17]), .B0(n1372), .S(n1371), .CO(n1370));
Q_AD01HF U1737 ( .A0(gfifoGBfullCnt[16]), .B0(n1374), .S(n1373), .CO(n1372));
Q_AD01HF U1738 ( .A0(gfifoGBfullCnt[15]), .B0(n1376), .S(n1375), .CO(n1374));
Q_AD01HF U1739 ( .A0(gfifoGBfullCnt[14]), .B0(n1378), .S(n1377), .CO(n1376));
Q_AD01HF U1740 ( .A0(gfifoGBfullCnt[13]), .B0(n1380), .S(n1379), .CO(n1378));
Q_AD01HF U1741 ( .A0(gfifoGBfullCnt[12]), .B0(n1382), .S(n1381), .CO(n1380));
Q_AD01HF U1742 ( .A0(gfifoGBfullCnt[11]), .B0(n1384), .S(n1383), .CO(n1382));
Q_AD01HF U1743 ( .A0(gfifoGBfullCnt[10]), .B0(n1386), .S(n1385), .CO(n1384));
Q_AD01HF U1744 ( .A0(gfifoGBfullCnt[9]), .B0(n1388), .S(n1387), .CO(n1386));
Q_AD01HF U1745 ( .A0(gfifoGBfullCnt[8]), .B0(n1390), .S(n1389), .CO(n1388));
Q_AD01HF U1746 ( .A0(gfifoGBfullCnt[7]), .B0(n1392), .S(n1391), .CO(n1390));
Q_AD01HF U1747 ( .A0(gfifoGBfullCnt[6]), .B0(n1394), .S(n1393), .CO(n1392));
Q_AD01HF U1748 ( .A0(gfifoGBfullCnt[5]), .B0(n1396), .S(n1395), .CO(n1394));
Q_AD01HF U1749 ( .A0(gfifoGBfullCnt[4]), .B0(n1398), .S(n1397), .CO(n1396));
Q_AD01HF U1750 ( .A0(gfifoGBfullCnt[3]), .B0(n1400), .S(n1399), .CO(n1398));
Q_AD01HF U1751 ( .A0(gfifoGBfullCnt[2]), .B0(n1402), .S(n1401), .CO(n1400));
Q_AD01HF U1752 ( .A0(gfifoGBfullCnt[1]), .B0(gfifoGBfullCnt[0]), .S(n1403), .CO(n1402));
Q_INV U1753 ( .A(sdlHaltHwClk), .Z(n1405));
Q_INV U1754 ( .A(sdlStop), .Z(n1404));
Q_AO21 U1755 ( .A0(sdlHaltHwClkR), .A1(n1404), .B0(n1405), .Z(n1407));
Q_INV U1756 ( .A(callEmuPre), .Z(n1406));
Q_NR02 U1757 ( .A0(callEmuPre), .A1(evalOnC), .Z(n1409));
Q_AN02 U1758 ( .A0(n1409), .A1(n1407), .Z(n1408));
Q_MX02 U1759 ( .S(n1408), .A0(n1411), .A1(hwClkHalt), .Z(n1410));
Q_FDP0UA U1760 ( .D(n1410), .QTFCLK( ), .Q(hwClkHalt));
Q_AO21 U1761 ( .A0(sdlStop), .A1(sdlHaltHwClk), .B0(n1409), .Z(n1411));
Q_FDP0UA U1762 ( .D(sdlHaltHwClk), .QTFCLK( ), .Q(sdlHaltHwClkR));
Q_MX02 U1763 ( .S(hwClkDbgOn), .A0(hwClkDelay[0]), .A1(n1650), .Z(n1412));
Q_FDP0UA U1764 ( .D(n1412), .QTFCLK( ), .Q(hwClkDelay[0]));
Q_MX02 U1765 ( .S(hwClkDbgOn), .A0(hwClkDelay[1]), .A1(n1649), .Z(n1413));
Q_FDP0UA U1766 ( .D(n1413), .QTFCLK( ), .Q(hwClkDelay[1]));
Q_MX02 U1767 ( .S(hwClkDbgOn), .A0(hwClkDelay[2]), .A1(n1648), .Z(n1414));
Q_FDP0UA U1768 ( .D(n1414), .QTFCLK( ), .Q(hwClkDelay[2]));
Q_MX02 U1769 ( .S(hwClkDbgOn), .A0(hwClkDelay[3]), .A1(n1647), .Z(n1415));
Q_FDP0UA U1770 ( .D(n1415), .QTFCLK( ), .Q(hwClkDelay[3]));
Q_MX02 U1771 ( .S(hwClkDbgOn), .A0(hwClkDelay[4]), .A1(n1646), .Z(n1416));
Q_FDP0UA U1772 ( .D(n1416), .QTFCLK( ), .Q(hwClkDelay[4]));
Q_MX02 U1773 ( .S(hwClkDbgOn), .A0(hwClkDelay[5]), .A1(n1645), .Z(n1417));
Q_FDP0UA U1774 ( .D(n1417), .QTFCLK( ), .Q(hwClkDelay[5]));
Q_MX02 U1775 ( .S(hwClkDbgOn), .A0(hwClkDelay[6]), .A1(n1644), .Z(n1418));
Q_FDP0UA U1776 ( .D(n1418), .QTFCLK( ), .Q(hwClkDelay[6]));
Q_MX02 U1777 ( .S(hwClkDbgOn), .A0(hwClkDelay[7]), .A1(n1643), .Z(n1419));
Q_FDP0UA U1778 ( .D(n1419), .QTFCLK( ), .Q(hwClkDelay[7]));
Q_MX02 U1779 ( .S(hwClkDbgOn), .A0(hwClkDelay[8]), .A1(n1642), .Z(n1420));
Q_FDP0UA U1780 ( .D(n1420), .QTFCLK( ), .Q(hwClkDelay[8]));
Q_MX02 U1781 ( .S(hwClkDbgOn), .A0(hwClkDelay[9]), .A1(n1641), .Z(n1421));
Q_FDP0UA U1782 ( .D(n1421), .QTFCLK( ), .Q(hwClkDelay[9]));
Q_MX02 U1783 ( .S(hwClkDbgOn), .A0(hwClkDelay[10]), .A1(n1640), .Z(n1422));
Q_FDP0UA U1784 ( .D(n1422), .QTFCLK( ), .Q(hwClkDelay[10]));
Q_MX02 U1785 ( .S(hwClkDbgOn), .A0(hwClkDelay[11]), .A1(n1639), .Z(n1423));
Q_FDP0UA U1786 ( .D(n1423), .QTFCLK( ), .Q(hwClkDelay[11]));
Q_MX02 U1787 ( .S(hwClkDbgOn), .A0(hwClkDelay[12]), .A1(n1638), .Z(n1424));
Q_FDP0UA U1788 ( .D(n1424), .QTFCLK( ), .Q(hwClkDelay[12]));
Q_MX02 U1789 ( .S(hwClkDbgOn), .A0(hwClkDelay[13]), .A1(n1637), .Z(n1425));
Q_FDP0UA U1790 ( .D(n1425), .QTFCLK( ), .Q(hwClkDelay[13]));
Q_MX02 U1791 ( .S(hwClkDbgOn), .A0(hwClkDelay[14]), .A1(n1636), .Z(n1426));
Q_FDP0UA U1792 ( .D(n1426), .QTFCLK( ), .Q(hwClkDelay[14]));
Q_MX02 U1793 ( .S(hwClkDbgOn), .A0(hwClkDelay[15]), .A1(n1635), .Z(n1427));
Q_FDP0UA U1794 ( .D(n1427), .QTFCLK( ), .Q(hwClkDelay[15]));
Q_MX02 U1795 ( .S(hwClkDbgOn), .A0(hwClkDelay[16]), .A1(n1634), .Z(n1428));
Q_FDP0UA U1796 ( .D(n1428), .QTFCLK( ), .Q(hwClkDelay[16]));
Q_MX02 U1797 ( .S(hwClkDbgOn), .A0(hwClkDelay[17]), .A1(n1633), .Z(n1429));
Q_FDP0UA U1798 ( .D(n1429), .QTFCLK( ), .Q(hwClkDelay[17]));
Q_MX02 U1799 ( .S(hwClkDbgOn), .A0(hwClkDelay[18]), .A1(n1632), .Z(n1430));
Q_FDP0UA U1800 ( .D(n1430), .QTFCLK( ), .Q(hwClkDelay[18]));
Q_MX02 U1801 ( .S(hwClkDbgOn), .A0(hwClkDelay[19]), .A1(n1631), .Z(n1431));
Q_FDP0UA U1802 ( .D(n1431), .QTFCLK( ), .Q(hwClkDelay[19]));
Q_MX02 U1803 ( .S(hwClkDbgOn), .A0(hwClkDelay[20]), .A1(n1630), .Z(n1432));
Q_FDP0UA U1804 ( .D(n1432), .QTFCLK( ), .Q(hwClkDelay[20]));
Q_MX02 U1805 ( .S(hwClkDbgOn), .A0(hwClkDelay[21]), .A1(n1629), .Z(n1433));
Q_FDP0UA U1806 ( .D(n1433), .QTFCLK( ), .Q(hwClkDelay[21]));
Q_MX02 U1807 ( .S(hwClkDbgOn), .A0(hwClkDelay[22]), .A1(n1628), .Z(n1434));
Q_FDP0UA U1808 ( .D(n1434), .QTFCLK( ), .Q(hwClkDelay[22]));
Q_MX02 U1809 ( .S(hwClkDbgOn), .A0(hwClkDelay[23]), .A1(n1627), .Z(n1435));
Q_FDP0UA U1810 ( .D(n1435), .QTFCLK( ), .Q(hwClkDelay[23]));
Q_MX02 U1811 ( .S(hwClkDbgOn), .A0(hwClkDelay[24]), .A1(n1626), .Z(n1436));
Q_FDP0UA U1812 ( .D(n1436), .QTFCLK( ), .Q(hwClkDelay[24]));
Q_MX02 U1813 ( .S(hwClkDbgOn), .A0(hwClkDelay[25]), .A1(n1625), .Z(n1437));
Q_FDP0UA U1814 ( .D(n1437), .QTFCLK( ), .Q(hwClkDelay[25]));
Q_MX02 U1815 ( .S(hwClkDbgOn), .A0(hwClkDelay[26]), .A1(n1624), .Z(n1438));
Q_FDP0UA U1816 ( .D(n1438), .QTFCLK( ), .Q(hwClkDelay[26]));
Q_MX02 U1817 ( .S(hwClkDbgOn), .A0(hwClkDelay[27]), .A1(n1623), .Z(n1439));
Q_FDP0UA U1818 ( .D(n1439), .QTFCLK( ), .Q(hwClkDelay[27]));
Q_MX02 U1819 ( .S(hwClkDbgOn), .A0(hwClkDelay[28]), .A1(n1622), .Z(n1440));
Q_FDP0UA U1820 ( .D(n1440), .QTFCLK( ), .Q(hwClkDelay[28]));
Q_MX02 U1821 ( .S(hwClkDbgOn), .A0(hwClkDelay[29]), .A1(n1621), .Z(n1441));
Q_FDP0UA U1822 ( .D(n1441), .QTFCLK( ), .Q(hwClkDelay[29]));
Q_MX02 U1823 ( .S(hwClkDbgOn), .A0(hwClkDelay[30]), .A1(n1620), .Z(n1442));
Q_FDP0UA U1824 ( .D(n1442), .QTFCLK( ), .Q(hwClkDelay[30]));
Q_MX02 U1825 ( .S(hwClkDbgOn), .A0(hwClkDelay[31]), .A1(n1619), .Z(n1443));
Q_FDP0UA U1826 ( .D(n1443), .QTFCLK( ), .Q(hwClkDelay[31]));
Q_MX02 U1827 ( .S(hwClkDbgOn), .A0(hwSimTime[0]), .A1(n1618), .Z(n1444));
Q_FDP0UA U1828 ( .D(n1444), .QTFCLK( ), .Q(hwSimTime[0]));
Q_MX02 U1829 ( .S(hwClkDbgOn), .A0(hwSimTime[1]), .A1(n1616), .Z(n1445));
Q_FDP0UA U1830 ( .D(n1445), .QTFCLK( ), .Q(hwSimTime[1]));
Q_MX02 U1831 ( .S(hwClkDbgOn), .A0(hwSimTime[2]), .A1(n1614), .Z(n1446));
Q_FDP0UA U1832 ( .D(n1446), .QTFCLK( ), .Q(hwSimTime[2]));
Q_MX02 U1833 ( .S(hwClkDbgOn), .A0(hwSimTime[3]), .A1(n1613), .Z(n1447));
Q_FDP0UA U1834 ( .D(n1447), .QTFCLK( ), .Q(hwSimTime[3]));
Q_MX02 U1835 ( .S(hwClkDbgOn), .A0(hwSimTime[4]), .A1(n1611), .Z(n1448));
Q_FDP0UA U1836 ( .D(n1448), .QTFCLK( ), .Q(hwSimTime[4]));
Q_MX02 U1837 ( .S(hwClkDbgOn), .A0(hwSimTime[5]), .A1(n1610), .Z(n1449));
Q_FDP0UA U1838 ( .D(n1449), .QTFCLK( ), .Q(hwSimTime[5]));
Q_MX02 U1839 ( .S(hwClkDbgOn), .A0(hwSimTime[6]), .A1(n1608), .Z(n1450));
Q_FDP0UA U1840 ( .D(n1450), .QTFCLK( ), .Q(hwSimTime[6]));
Q_MX02 U1841 ( .S(hwClkDbgOn), .A0(hwSimTime[7]), .A1(n1607), .Z(n1451));
Q_FDP0UA U1842 ( .D(n1451), .QTFCLK( ), .Q(hwSimTime[7]));
Q_MX02 U1843 ( .S(hwClkDbgOn), .A0(hwSimTime[8]), .A1(n1605), .Z(n1452));
Q_FDP0UA U1844 ( .D(n1452), .QTFCLK( ), .Q(hwSimTime[8]));
Q_MX02 U1845 ( .S(hwClkDbgOn), .A0(hwSimTime[9]), .A1(n1604), .Z(n1453));
Q_FDP0UA U1846 ( .D(n1453), .QTFCLK( ), .Q(hwSimTime[9]));
Q_MX02 U1847 ( .S(hwClkDbgOn), .A0(hwSimTime[10]), .A1(n1602), .Z(n1454));
Q_FDP0UA U1848 ( .D(n1454), .QTFCLK( ), .Q(hwSimTime[10]));
Q_MX02 U1849 ( .S(hwClkDbgOn), .A0(hwSimTime[11]), .A1(n1601), .Z(n1455));
Q_FDP0UA U1850 ( .D(n1455), .QTFCLK( ), .Q(hwSimTime[11]));
Q_MX02 U1851 ( .S(hwClkDbgOn), .A0(hwSimTime[12]), .A1(n1599), .Z(n1456));
Q_FDP0UA U1852 ( .D(n1456), .QTFCLK( ), .Q(hwSimTime[12]));
Q_MX02 U1853 ( .S(hwClkDbgOn), .A0(hwSimTime[13]), .A1(n1598), .Z(n1457));
Q_FDP0UA U1854 ( .D(n1457), .QTFCLK( ), .Q(hwSimTime[13]));
Q_MX02 U1855 ( .S(hwClkDbgOn), .A0(hwSimTime[14]), .A1(n1596), .Z(n1458));
Q_FDP0UA U1856 ( .D(n1458), .QTFCLK( ), .Q(hwSimTime[14]));
Q_MX02 U1857 ( .S(hwClkDbgOn), .A0(hwSimTime[15]), .A1(n1595), .Z(n1459));
Q_FDP0UA U1858 ( .D(n1459), .QTFCLK( ), .Q(hwSimTime[15]));
Q_MX02 U1859 ( .S(hwClkDbgOn), .A0(hwSimTime[16]), .A1(n1593), .Z(n1460));
Q_FDP0UA U1860 ( .D(n1460), .QTFCLK( ), .Q(hwSimTime[16]));
Q_MX02 U1861 ( .S(hwClkDbgOn), .A0(hwSimTime[17]), .A1(n1592), .Z(n1461));
Q_FDP0UA U1862 ( .D(n1461), .QTFCLK( ), .Q(hwSimTime[17]));
Q_MX02 U1863 ( .S(hwClkDbgOn), .A0(hwSimTime[18]), .A1(n1590), .Z(n1462));
Q_FDP0UA U1864 ( .D(n1462), .QTFCLK( ), .Q(hwSimTime[18]));
Q_MX02 U1865 ( .S(hwClkDbgOn), .A0(hwSimTime[19]), .A1(n1589), .Z(n1463));
Q_FDP0UA U1866 ( .D(n1463), .QTFCLK( ), .Q(hwSimTime[19]));
Q_MX02 U1867 ( .S(hwClkDbgOn), .A0(hwSimTime[20]), .A1(n1587), .Z(n1464));
Q_FDP0UA U1868 ( .D(n1464), .QTFCLK( ), .Q(hwSimTime[20]));
Q_MX02 U1869 ( .S(hwClkDbgOn), .A0(hwSimTime[21]), .A1(n1586), .Z(n1465));
Q_FDP0UA U1870 ( .D(n1465), .QTFCLK( ), .Q(hwSimTime[21]));
Q_MX02 U1871 ( .S(hwClkDbgOn), .A0(hwSimTime[22]), .A1(n1584), .Z(n1466));
Q_FDP0UA U1872 ( .D(n1466), .QTFCLK( ), .Q(hwSimTime[22]));
Q_MX02 U1873 ( .S(hwClkDbgOn), .A0(hwSimTime[23]), .A1(n1583), .Z(n1467));
Q_FDP0UA U1874 ( .D(n1467), .QTFCLK( ), .Q(hwSimTime[23]));
Q_MX02 U1875 ( .S(hwClkDbgOn), .A0(hwSimTime[24]), .A1(n1581), .Z(n1468));
Q_FDP0UA U1876 ( .D(n1468), .QTFCLK( ), .Q(hwSimTime[24]));
Q_MX02 U1877 ( .S(hwClkDbgOn), .A0(hwSimTime[25]), .A1(n1580), .Z(n1469));
Q_FDP0UA U1878 ( .D(n1469), .QTFCLK( ), .Q(hwSimTime[25]));
Q_MX02 U1879 ( .S(hwClkDbgOn), .A0(hwSimTime[26]), .A1(n1578), .Z(n1470));
Q_FDP0UA U1880 ( .D(n1470), .QTFCLK( ), .Q(hwSimTime[26]));
Q_MX02 U1881 ( .S(hwClkDbgOn), .A0(hwSimTime[27]), .A1(n1577), .Z(n1471));
Q_FDP0UA U1882 ( .D(n1471), .QTFCLK( ), .Q(hwSimTime[27]));
Q_MX02 U1883 ( .S(hwClkDbgOn), .A0(hwSimTime[28]), .A1(n1575), .Z(n1472));
Q_FDP0UA U1884 ( .D(n1472), .QTFCLK( ), .Q(hwSimTime[28]));
Q_MX02 U1885 ( .S(hwClkDbgOn), .A0(hwSimTime[29]), .A1(n1574), .Z(n1473));
Q_FDP0UA U1886 ( .D(n1473), .QTFCLK( ), .Q(hwSimTime[29]));
Q_MX02 U1887 ( .S(hwClkDbgOn), .A0(hwSimTime[30]), .A1(n1572), .Z(n1474));
Q_FDP0UA U1888 ( .D(n1474), .QTFCLK( ), .Q(hwSimTime[30]));
Q_MX02 U1889 ( .S(hwClkDbgOn), .A0(hwSimTime[31]), .A1(n1571), .Z(n1475));
Q_FDP0UA U1890 ( .D(n1475), .QTFCLK( ), .Q(hwSimTime[31]));
Q_MX02 U1891 ( .S(hwClkDbgOn), .A0(hwSimTime[32]), .A1(n1569), .Z(n1476));
Q_FDP0UA U1892 ( .D(n1476), .QTFCLK( ), .Q(hwSimTime[32]));
Q_MX02 U1893 ( .S(hwClkDbgOn), .A0(hwSimTime[33]), .A1(n1567), .Z(n1477));
Q_FDP0UA U1894 ( .D(n1477), .QTFCLK( ), .Q(hwSimTime[33]));
Q_MX02 U1895 ( .S(hwClkDbgOn), .A0(hwSimTime[34]), .A1(n1565), .Z(n1478));
Q_FDP0UA U1896 ( .D(n1478), .QTFCLK( ), .Q(hwSimTime[34]));
Q_MX02 U1897 ( .S(hwClkDbgOn), .A0(hwSimTime[35]), .A1(n1563), .Z(n1479));
Q_FDP0UA U1898 ( .D(n1479), .QTFCLK( ), .Q(hwSimTime[35]));
Q_MX02 U1899 ( .S(hwClkDbgOn), .A0(hwSimTime[36]), .A1(n1561), .Z(n1480));
Q_FDP0UA U1900 ( .D(n1480), .QTFCLK( ), .Q(hwSimTime[36]));
Q_MX02 U1901 ( .S(hwClkDbgOn), .A0(hwSimTime[37]), .A1(n1559), .Z(n1481));
Q_FDP0UA U1902 ( .D(n1481), .QTFCLK( ), .Q(hwSimTime[37]));
Q_MX02 U1903 ( .S(hwClkDbgOn), .A0(hwSimTime[38]), .A1(n1557), .Z(n1482));
Q_FDP0UA U1904 ( .D(n1482), .QTFCLK( ), .Q(hwSimTime[38]));
Q_MX02 U1905 ( .S(hwClkDbgOn), .A0(hwSimTime[39]), .A1(n1555), .Z(n1483));
Q_FDP0UA U1906 ( .D(n1483), .QTFCLK( ), .Q(hwSimTime[39]));
Q_MX02 U1907 ( .S(hwClkDbgOn), .A0(hwSimTime[40]), .A1(n1553), .Z(n1484));
Q_FDP0UA U1908 ( .D(n1484), .QTFCLK( ), .Q(hwSimTime[40]));
Q_MX02 U1909 ( .S(hwClkDbgOn), .A0(hwSimTime[41]), .A1(n1551), .Z(n1485));
Q_FDP0UA U1910 ( .D(n1485), .QTFCLK( ), .Q(hwSimTime[41]));
Q_MX02 U1911 ( .S(hwClkDbgOn), .A0(hwSimTime[42]), .A1(n1549), .Z(n1486));
Q_FDP0UA U1912 ( .D(n1486), .QTFCLK( ), .Q(hwSimTime[42]));
Q_MX02 U1913 ( .S(hwClkDbgOn), .A0(hwSimTime[43]), .A1(n1547), .Z(n1487));
Q_FDP0UA U1914 ( .D(n1487), .QTFCLK( ), .Q(hwSimTime[43]));
Q_MX02 U1915 ( .S(hwClkDbgOn), .A0(hwSimTime[44]), .A1(n1545), .Z(n1488));
Q_FDP0UA U1916 ( .D(n1488), .QTFCLK( ), .Q(hwSimTime[44]));
Q_MX02 U1917 ( .S(hwClkDbgOn), .A0(hwSimTime[45]), .A1(n1543), .Z(n1489));
Q_FDP0UA U1918 ( .D(n1489), .QTFCLK( ), .Q(hwSimTime[45]));
Q_MX02 U1919 ( .S(hwClkDbgOn), .A0(hwSimTime[46]), .A1(n1541), .Z(n1490));
Q_FDP0UA U1920 ( .D(n1490), .QTFCLK( ), .Q(hwSimTime[46]));
Q_MX02 U1921 ( .S(hwClkDbgOn), .A0(hwSimTime[47]), .A1(n1539), .Z(n1491));
Q_FDP0UA U1922 ( .D(n1491), .QTFCLK( ), .Q(hwSimTime[47]));
Q_MX02 U1923 ( .S(hwClkDbgOn), .A0(hwSimTime[48]), .A1(n1537), .Z(n1492));
Q_FDP0UA U1924 ( .D(n1492), .QTFCLK( ), .Q(hwSimTime[48]));
Q_MX02 U1925 ( .S(hwClkDbgOn), .A0(hwSimTime[49]), .A1(n1535), .Z(n1493));
Q_FDP0UA U1926 ( .D(n1493), .QTFCLK( ), .Q(hwSimTime[49]));
Q_MX02 U1927 ( .S(hwClkDbgOn), .A0(hwSimTime[50]), .A1(n1533), .Z(n1494));
Q_FDP0UA U1928 ( .D(n1494), .QTFCLK( ), .Q(hwSimTime[50]));
Q_MX02 U1929 ( .S(hwClkDbgOn), .A0(hwSimTime[51]), .A1(n1531), .Z(n1495));
Q_FDP0UA U1930 ( .D(n1495), .QTFCLK( ), .Q(hwSimTime[51]));
Q_MX02 U1931 ( .S(hwClkDbgOn), .A0(hwSimTime[52]), .A1(n1529), .Z(n1496));
Q_FDP0UA U1932 ( .D(n1496), .QTFCLK( ), .Q(hwSimTime[52]));
Q_MX02 U1933 ( .S(hwClkDbgOn), .A0(hwSimTime[53]), .A1(n1527), .Z(n1497));
Q_FDP0UA U1934 ( .D(n1497), .QTFCLK( ), .Q(hwSimTime[53]));
Q_MX02 U1935 ( .S(hwClkDbgOn), .A0(hwSimTime[54]), .A1(n1525), .Z(n1498));
Q_FDP0UA U1936 ( .D(n1498), .QTFCLK( ), .Q(hwSimTime[54]));
Q_MX02 U1937 ( .S(hwClkDbgOn), .A0(hwSimTime[55]), .A1(n1523), .Z(n1499));
Q_FDP0UA U1938 ( .D(n1499), .QTFCLK( ), .Q(hwSimTime[55]));
Q_MX02 U1939 ( .S(hwClkDbgOn), .A0(hwSimTime[56]), .A1(n1521), .Z(n1500));
Q_FDP0UA U1940 ( .D(n1500), .QTFCLK( ), .Q(hwSimTime[56]));
Q_MX02 U1941 ( .S(hwClkDbgOn), .A0(hwSimTime[57]), .A1(n1519), .Z(n1501));
Q_FDP0UA U1942 ( .D(n1501), .QTFCLK( ), .Q(hwSimTime[57]));
Q_MX02 U1943 ( .S(hwClkDbgOn), .A0(hwSimTime[58]), .A1(n1517), .Z(n1502));
Q_FDP0UA U1944 ( .D(n1502), .QTFCLK( ), .Q(hwSimTime[58]));
Q_MX02 U1945 ( .S(hwClkDbgOn), .A0(hwSimTime[59]), .A1(n1515), .Z(n1503));
Q_FDP0UA U1946 ( .D(n1503), .QTFCLK( ), .Q(hwSimTime[59]));
Q_MX02 U1947 ( .S(hwClkDbgOn), .A0(hwSimTime[60]), .A1(n1513), .Z(n1504));
Q_FDP0UA U1948 ( .D(n1504), .QTFCLK( ), .Q(hwSimTime[60]));
Q_MX02 U1949 ( .S(hwClkDbgOn), .A0(hwSimTime[61]), .A1(n1511), .Z(n1505));
Q_FDP0UA U1950 ( .D(n1505), .QTFCLK( ), .Q(hwSimTime[61]));
Q_MX02 U1951 ( .S(hwClkDbgOn), .A0(hwSimTime[62]), .A1(n1509), .Z(n1506));
Q_FDP0UA U1952 ( .D(n1506), .QTFCLK( ), .Q(hwSimTime[62]));
Q_FDP0UA U1953 ( .D(n1507), .QTFCLK( ), .Q(hwSimTime[63]));
Q_XOR2 U1954 ( .A0(hwSimTime[63]), .A1(n10), .Z(n1507));
Q_AD01HF U1955 ( .A0(hwSimTime[62]), .B0(n1510), .S(n1509), .CO(n1508));
Q_AD01HF U1956 ( .A0(hwSimTime[61]), .B0(n1512), .S(n1511), .CO(n1510));
Q_AD01HF U1957 ( .A0(hwSimTime[60]), .B0(n1514), .S(n1513), .CO(n1512));
Q_AD01HF U1958 ( .A0(hwSimTime[59]), .B0(n1516), .S(n1515), .CO(n1514));
Q_AD01HF U1959 ( .A0(hwSimTime[58]), .B0(n1518), .S(n1517), .CO(n1516));
Q_AD01HF U1960 ( .A0(hwSimTime[57]), .B0(n1520), .S(n1519), .CO(n1518));
Q_AD01HF U1961 ( .A0(hwSimTime[56]), .B0(n1522), .S(n1521), .CO(n1520));
Q_AD01HF U1962 ( .A0(hwSimTime[55]), .B0(n1524), .S(n1523), .CO(n1522));
Q_AD01HF U1963 ( .A0(hwSimTime[54]), .B0(n1526), .S(n1525), .CO(n1524));
Q_AD01HF U1964 ( .A0(hwSimTime[53]), .B0(n1528), .S(n1527), .CO(n1526));
Q_AD01HF U1965 ( .A0(hwSimTime[52]), .B0(n1530), .S(n1529), .CO(n1528));
Q_AD01HF U1966 ( .A0(hwSimTime[51]), .B0(n1532), .S(n1531), .CO(n1530));
Q_AD01HF U1967 ( .A0(hwSimTime[50]), .B0(n1534), .S(n1533), .CO(n1532));
Q_AD01HF U1968 ( .A0(hwSimTime[49]), .B0(n1536), .S(n1535), .CO(n1534));
Q_AD01HF U1969 ( .A0(hwSimTime[48]), .B0(n1538), .S(n1537), .CO(n1536));
Q_AD01HF U1970 ( .A0(hwSimTime[47]), .B0(n1540), .S(n1539), .CO(n1538));
Q_AD01HF U1971 ( .A0(hwSimTime[46]), .B0(n1542), .S(n1541), .CO(n1540));
Q_AD01HF U1972 ( .A0(hwSimTime[45]), .B0(n1544), .S(n1543), .CO(n1542));
Q_AD01HF U1973 ( .A0(hwSimTime[44]), .B0(n1546), .S(n1545), .CO(n1544));
Q_AD01HF U1974 ( .A0(hwSimTime[43]), .B0(n1548), .S(n1547), .CO(n1546));
Q_AD01HF U1975 ( .A0(hwSimTime[42]), .B0(n1550), .S(n1549), .CO(n1548));
Q_AD01HF U1976 ( .A0(hwSimTime[41]), .B0(n1552), .S(n1551), .CO(n1550));
Q_AD01HF U1977 ( .A0(hwSimTime[40]), .B0(n1554), .S(n1553), .CO(n1552));
Q_AD01HF U1978 ( .A0(hwSimTime[39]), .B0(n1556), .S(n1555), .CO(n1554));
Q_AD01HF U1979 ( .A0(hwSimTime[38]), .B0(n1558), .S(n1557), .CO(n1556));
Q_AD01HF U1980 ( .A0(hwSimTime[37]), .B0(n1560), .S(n1559), .CO(n1558));
Q_AD01HF U1981 ( .A0(hwSimTime[36]), .B0(n1562), .S(n1561), .CO(n1560));
Q_AD01HF U1982 ( .A0(hwSimTime[35]), .B0(n1564), .S(n1563), .CO(n1562));
Q_AD01HF U1983 ( .A0(hwSimTime[34]), .B0(n1566), .S(n1565), .CO(n1564));
Q_AD01HF U1984 ( .A0(hwSimTime[33]), .B0(n1568), .S(n1567), .CO(n1566));
Q_AD01HF U1985 ( .A0(hwSimTime[32]), .B0(n1570), .S(n1569), .CO(n1568));
Q_AD02 U1986 ( .CI(n1573), .A0(hwSimTime[30]), .A1(hwSimTime[31]), .B0(n1620), .B1(n1619), .S0(n1572), .S1(n1571), .CO(n1570));
Q_AD02 U1987 ( .CI(n1576), .A0(hwSimTime[28]), .A1(hwSimTime[29]), .B0(n1622), .B1(n1621), .S0(n1575), .S1(n1574), .CO(n1573));
Q_AD02 U1988 ( .CI(n1579), .A0(hwSimTime[26]), .A1(hwSimTime[27]), .B0(n1624), .B1(n1623), .S0(n1578), .S1(n1577), .CO(n1576));
Q_AD02 U1989 ( .CI(n1582), .A0(hwSimTime[24]), .A1(hwSimTime[25]), .B0(n1626), .B1(n1625), .S0(n1581), .S1(n1580), .CO(n1579));
Q_AD02 U1990 ( .CI(n1585), .A0(hwSimTime[22]), .A1(hwSimTime[23]), .B0(n1628), .B1(n1627), .S0(n1584), .S1(n1583), .CO(n1582));
Q_AD02 U1991 ( .CI(n1588), .A0(hwSimTime[20]), .A1(hwSimTime[21]), .B0(n1630), .B1(n1629), .S0(n1587), .S1(n1586), .CO(n1585));
Q_AD02 U1992 ( .CI(n1591), .A0(hwSimTime[18]), .A1(hwSimTime[19]), .B0(n1632), .B1(n1631), .S0(n1590), .S1(n1589), .CO(n1588));
Q_AD02 U1993 ( .CI(n1594), .A0(hwSimTime[16]), .A1(hwSimTime[17]), .B0(n1634), .B1(n1633), .S0(n1593), .S1(n1592), .CO(n1591));
Q_AD02 U1994 ( .CI(n1597), .A0(hwSimTime[14]), .A1(hwSimTime[15]), .B0(n1636), .B1(n1635), .S0(n1596), .S1(n1595), .CO(n1594));
Q_AD02 U1995 ( .CI(n1600), .A0(hwSimTime[12]), .A1(hwSimTime[13]), .B0(n1638), .B1(n1637), .S0(n1599), .S1(n1598), .CO(n1597));
Q_AD02 U1996 ( .CI(n1603), .A0(hwSimTime[10]), .A1(hwSimTime[11]), .B0(n1640), .B1(n1639), .S0(n1602), .S1(n1601), .CO(n1600));
Q_AD02 U1997 ( .CI(n1606), .A0(hwSimTime[8]), .A1(hwSimTime[9]), .B0(n1642), .B1(n1641), .S0(n1605), .S1(n1604), .CO(n1603));
Q_AD02 U1998 ( .CI(n1609), .A0(hwSimTime[6]), .A1(hwSimTime[7]), .B0(n1644), .B1(n1643), .S0(n1608), .S1(n1607), .CO(n1606));
Q_AD02 U1999 ( .CI(n1612), .A0(hwSimTime[4]), .A1(hwSimTime[5]), .B0(n1646), .B1(n1645), .S0(n1611), .S1(n1610), .CO(n1609));
Q_AD02 U2000 ( .CI(n1615), .A0(hwSimTime[2]), .A1(hwSimTime[3]), .B0(n1648), .B1(n1647), .S0(n1614), .S1(n1613), .CO(n1612));
Q_AD01 U2001 ( .CI(n1649), .A0(hwSimTime[1]), .B0(n1617), .S(n1616), .CO(n1615));
Q_AD01HF U2002 ( .A0(hwSimTime[0]), .B0(n1650), .S(n1618), .CO(n1617));
Q_AN02 U2003 ( .A0(n1652), .A1(hwClkDelay[31]), .Z(n1619));
Q_AN02 U2004 ( .A0(n1652), .A1(hwClkDelay[30]), .Z(n1620));
Q_AN02 U2005 ( .A0(n1652), .A1(hwClkDelay[29]), .Z(n1621));
Q_AN02 U2006 ( .A0(n1652), .A1(hwClkDelay[28]), .Z(n1622));
Q_AN02 U2007 ( .A0(n1652), .A1(hwClkDelay[27]), .Z(n1623));
Q_AN02 U2008 ( .A0(n1652), .A1(hwClkDelay[26]), .Z(n1624));
Q_AN02 U2009 ( .A0(n1652), .A1(hwClkDelay[25]), .Z(n1625));
Q_AN02 U2010 ( .A0(n1652), .A1(hwClkDelay[24]), .Z(n1626));
Q_AN02 U2011 ( .A0(n1652), .A1(hwClkDelay[23]), .Z(n1627));
Q_AN02 U2012 ( .A0(n1652), .A1(hwClkDelay[22]), .Z(n1628));
Q_AN02 U2013 ( .A0(n1652), .A1(hwClkDelay[21]), .Z(n1629));
Q_AN02 U2014 ( .A0(n1652), .A1(hwClkDelay[20]), .Z(n1630));
Q_AN02 U2015 ( .A0(n1652), .A1(hwClkDelay[19]), .Z(n1631));
Q_AN02 U2016 ( .A0(n1652), .A1(hwClkDelay[18]), .Z(n1632));
Q_AN02 U2017 ( .A0(n1652), .A1(hwClkDelay[17]), .Z(n1633));
Q_AN02 U2018 ( .A0(n1652), .A1(hwClkDelay[16]), .Z(n1634));
Q_AN02 U2019 ( .A0(n1652), .A1(hwClkDelay[15]), .Z(n1635));
Q_AN02 U2020 ( .A0(n1652), .A1(hwClkDelay[14]), .Z(n1636));
Q_AN02 U2021 ( .A0(n1652), .A1(hwClkDelay[13]), .Z(n1637));
Q_AN02 U2022 ( .A0(n1652), .A1(hwClkDelay[12]), .Z(n1638));
Q_AN02 U2023 ( .A0(n1652), .A1(hwClkDelay[11]), .Z(n1639));
Q_AN02 U2024 ( .A0(n1652), .A1(hwClkDelay[10]), .Z(n1640));
Q_AN02 U2025 ( .A0(n1652), .A1(hwClkDelay[9]), .Z(n1641));
Q_AN02 U2026 ( .A0(n1652), .A1(hwClkDelay[8]), .Z(n1642));
Q_AN02 U2027 ( .A0(n1652), .A1(hwClkDelay[7]), .Z(n1643));
Q_AN02 U2028 ( .A0(n1652), .A1(hwClkDelay[6]), .Z(n1644));
Q_AN02 U2029 ( .A0(n1652), .A1(hwClkDelay[5]), .Z(n1645));
Q_AN02 U2030 ( .A0(n1652), .A1(hwClkDelay[4]), .Z(n1646));
Q_AN02 U2031 ( .A0(n1652), .A1(hwClkDelay[3]), .Z(n1647));
Q_AN02 U2032 ( .A0(n1652), .A1(hwClkDelay[2]), .Z(n1648));
Q_AN02 U2033 ( .A0(n1652), .A1(hwClkDelay[1]), .Z(n1649));
Q_OR02 U2034 ( .A0(n1651), .A1(hwClkDelay[0]), .Z(n1650));
Q_INV U2035 ( .A(n1652), .Z(n1651));
Q_OR02 U2036 ( .A0(n1654), .A1(n1653), .Z(n1652));
Q_OR03 U2037 ( .A0(n1657), .A1(n1656), .A2(n1655), .Z(n1653));
Q_OR03 U2038 ( .A0(n1660), .A1(n1659), .A2(n1658), .Z(n1654));
Q_OR03 U2039 ( .A0(n1663), .A1(n1662), .A2(n1661), .Z(n1655));
Q_OR03 U2040 ( .A0(n1666), .A1(n1665), .A2(n1664), .Z(n1656));
Q_OR03 U2041 ( .A0(hwClkDelay[1]), .A1(hwClkDelay[0]), .A2(n1667), .Z(n1657));
Q_OR03 U2042 ( .A0(hwClkDelay[4]), .A1(hwClkDelay[3]), .A2(hwClkDelay[2]), .Z(n1658));
Q_OR03 U2043 ( .A0(hwClkDelay[7]), .A1(hwClkDelay[6]), .A2(hwClkDelay[5]), .Z(n1659));
Q_OR03 U2044 ( .A0(hwClkDelay[10]), .A1(hwClkDelay[9]), .A2(hwClkDelay[8]), .Z(n1660));
Q_OR03 U2045 ( .A0(hwClkDelay[13]), .A1(hwClkDelay[12]), .A2(hwClkDelay[11]), .Z(n1661));
Q_OR03 U2046 ( .A0(hwClkDelay[16]), .A1(hwClkDelay[15]), .A2(hwClkDelay[14]), .Z(n1662));
Q_OR03 U2047 ( .A0(hwClkDelay[19]), .A1(hwClkDelay[18]), .A2(hwClkDelay[17]), .Z(n1663));
Q_OR03 U2048 ( .A0(hwClkDelay[22]), .A1(hwClkDelay[21]), .A2(hwClkDelay[20]), .Z(n1664));
Q_OR03 U2049 ( .A0(hwClkDelay[25]), .A1(hwClkDelay[24]), .A2(hwClkDelay[23]), .Z(n1665));
Q_OR03 U2050 ( .A0(hwClkDelay[28]), .A1(hwClkDelay[27]), .A2(hwClkDelay[26]), .Z(n1666));
Q_OR03 U2051 ( .A0(hwClkDelay[31]), .A1(hwClkDelay[30]), .A2(hwClkDelay[29]), .Z(n1667));
Q_AO21 U2052 ( .A0(ckgHoldPIi), .A1(oneStepPIi), .B0(n1406), .Z(n1669));
Q_INV U2053 ( .A(n1669), .Z(n1668));
Q_OR02 U2054 ( .A0(n1668), .A1(hwClkEnable), .Z(n1670));
Q_FDP0UA U2055 ( .D(n1670), .QTFCLK( ), .Q(hwClkEnable));
Q_FDP0UA U2056 ( .D(dummyW), .QTFCLK( ), .Q(dummyR));
Q_FDP0UA U2057 ( .D(it_capture), .QTFCLK( ), .Q(it_capture));
Q_FDP0UA U2058 ( .D(it_replay), .QTFCLK( ), .Q(it_replay));
Q_INV U2059 ( .A(acHalt), .Z(n1672));
Q_AN02 U2060 ( .A0(asyncCall), .A1(n1672), .Z(n1673));
Q_AN02 U2061 ( .A0(n1673), .A1(n503), .Z(n1671));
Q_XOR2 U2062 ( .A0(n1671), .A1(aCount[0]), .Z(n1674));
Q_FDP0UA U2063 ( .D(n1674), .QTFCLK( ), .Q(aCount[0]));
Q_MX02 U2064 ( .S(n1671), .A0(aCount[1]), .A1(n1765), .Z(n1675));
Q_FDP0UA U2065 ( .D(n1675), .QTFCLK( ), .Q(aCount[1]));
Q_MX02 U2066 ( .S(n1671), .A0(aCount[2]), .A1(n1763), .Z(n1676));
Q_FDP0UA U2067 ( .D(n1676), .QTFCLK( ), .Q(aCount[2]));
Q_MX02 U2068 ( .S(n1671), .A0(aCount[3]), .A1(n1761), .Z(n1677));
Q_FDP0UA U2069 ( .D(n1677), .QTFCLK( ), .Q(aCount[3]));
Q_MX02 U2070 ( .S(n1671), .A0(aCount[4]), .A1(n1759), .Z(n1678));
Q_FDP0UA U2071 ( .D(n1678), .QTFCLK( ), .Q(aCount[4]));
Q_MX02 U2072 ( .S(n1671), .A0(aCount[5]), .A1(n1757), .Z(n1679));
Q_FDP0UA U2073 ( .D(n1679), .QTFCLK( ), .Q(aCount[5]));
Q_MX02 U2074 ( .S(n1671), .A0(aCount[6]), .A1(n1755), .Z(n1680));
Q_FDP0UA U2075 ( .D(n1680), .QTFCLK( ), .Q(aCount[6]));
Q_MX02 U2076 ( .S(n1671), .A0(aCount[7]), .A1(n1753), .Z(n1681));
Q_FDP0UA U2077 ( .D(n1681), .QTFCLK( ), .Q(aCount[7]));
Q_MX02 U2078 ( .S(n1671), .A0(aCount[8]), .A1(n1751), .Z(n1682));
Q_FDP0UA U2079 ( .D(n1682), .QTFCLK( ), .Q(aCount[8]));
Q_MX02 U2080 ( .S(n1671), .A0(aCount[9]), .A1(n1749), .Z(n1683));
Q_FDP0UA U2081 ( .D(n1683), .QTFCLK( ), .Q(aCount[9]));
Q_MX02 U2082 ( .S(n1671), .A0(aCount[10]), .A1(n1747), .Z(n1684));
Q_FDP0UA U2083 ( .D(n1684), .QTFCLK( ), .Q(aCount[10]));
Q_MX02 U2084 ( .S(n1671), .A0(aCount[11]), .A1(n1745), .Z(n1685));
Q_FDP0UA U2085 ( .D(n1685), .QTFCLK( ), .Q(aCount[11]));
Q_MX02 U2086 ( .S(n1671), .A0(aCount[12]), .A1(n1743), .Z(n1686));
Q_FDP0UA U2087 ( .D(n1686), .QTFCLK( ), .Q(aCount[12]));
Q_MX02 U2088 ( .S(n1671), .A0(aCount[13]), .A1(n1741), .Z(n1687));
Q_FDP0UA U2089 ( .D(n1687), .QTFCLK( ), .Q(aCount[13]));
Q_MX02 U2090 ( .S(n1671), .A0(aCount[14]), .A1(n1739), .Z(n1688));
Q_FDP0UA U2091 ( .D(n1688), .QTFCLK( ), .Q(aCount[14]));
Q_MX02 U2092 ( .S(n1671), .A0(aCount[15]), .A1(n1737), .Z(n1689));
Q_FDP0UA U2093 ( .D(n1689), .QTFCLK( ), .Q(aCount[15]));
Q_MX02 U2094 ( .S(n1671), .A0(aCount[16]), .A1(n1735), .Z(n1690));
Q_FDP0UA U2095 ( .D(n1690), .QTFCLK( ), .Q(aCount[16]));
Q_MX02 U2096 ( .S(n1671), .A0(aCount[17]), .A1(n1733), .Z(n1691));
Q_FDP0UA U2097 ( .D(n1691), .QTFCLK( ), .Q(aCount[17]));
Q_MX02 U2098 ( .S(n1671), .A0(aCount[18]), .A1(n1731), .Z(n1692));
Q_FDP0UA U2099 ( .D(n1692), .QTFCLK( ), .Q(aCount[18]));
Q_MX02 U2100 ( .S(n1671), .A0(aCount[19]), .A1(n1729), .Z(n1693));
Q_FDP0UA U2101 ( .D(n1693), .QTFCLK( ), .Q(aCount[19]));
Q_MX02 U2102 ( .S(n1671), .A0(aCount[20]), .A1(n1727), .Z(n1694));
Q_FDP0UA U2103 ( .D(n1694), .QTFCLK( ), .Q(aCount[20]));
Q_MX02 U2104 ( .S(n1671), .A0(aCount[21]), .A1(n1725), .Z(n1695));
Q_FDP0UA U2105 ( .D(n1695), .QTFCLK( ), .Q(aCount[21]));
Q_MX02 U2106 ( .S(n1671), .A0(aCount[22]), .A1(n1723), .Z(n1696));
Q_FDP0UA U2107 ( .D(n1696), .QTFCLK( ), .Q(aCount[22]));
Q_MX02 U2108 ( .S(n1671), .A0(aCount[23]), .A1(n1721), .Z(n1697));
Q_FDP0UA U2109 ( .D(n1697), .QTFCLK( ), .Q(aCount[23]));
Q_MX02 U2110 ( .S(n1671), .A0(aCount[24]), .A1(n1719), .Z(n1698));
Q_FDP0UA U2111 ( .D(n1698), .QTFCLK( ), .Q(aCount[24]));
Q_MX02 U2112 ( .S(n1671), .A0(aCount[25]), .A1(n1717), .Z(n1699));
Q_FDP0UA U2113 ( .D(n1699), .QTFCLK( ), .Q(aCount[25]));
Q_MX02 U2114 ( .S(n1671), .A0(aCount[26]), .A1(n1715), .Z(n1700));
Q_FDP0UA U2115 ( .D(n1700), .QTFCLK( ), .Q(aCount[26]));
Q_MX02 U2116 ( .S(n1671), .A0(aCount[27]), .A1(n1713), .Z(n1701));
Q_FDP0UA U2117 ( .D(n1701), .QTFCLK( ), .Q(aCount[27]));
Q_MX02 U2118 ( .S(n1671), .A0(aCount[28]), .A1(n1711), .Z(n1702));
Q_FDP0UA U2119 ( .D(n1702), .QTFCLK( ), .Q(aCount[28]));
Q_MX02 U2120 ( .S(n1671), .A0(aCount[29]), .A1(n1709), .Z(n1703));
Q_FDP0UA U2121 ( .D(n1703), .QTFCLK( ), .Q(aCount[29]));
Q_MX02 U2122 ( .S(n1671), .A0(aCount[30]), .A1(n1707), .Z(n1704));
Q_FDP0UA U2123 ( .D(n1704), .QTFCLK( ), .Q(aCount[30]));
Q_FDP0UA U2124 ( .D(n1705), .QTFCLK( ), .Q(aCount[31]));
Q_XOR2 U2125 ( .A0(aCount[31]), .A1(n9), .Z(n1705));
Q_AD01HF U2126 ( .A0(aCount[30]), .B0(n1708), .S(n1707), .CO(n1706));
Q_AD01HF U2127 ( .A0(aCount[29]), .B0(n1710), .S(n1709), .CO(n1708));
Q_AD01HF U2128 ( .A0(aCount[28]), .B0(n1712), .S(n1711), .CO(n1710));
Q_AD01HF U2129 ( .A0(aCount[27]), .B0(n1714), .S(n1713), .CO(n1712));
Q_AD01HF U2130 ( .A0(aCount[26]), .B0(n1716), .S(n1715), .CO(n1714));
Q_AD01HF U2131 ( .A0(aCount[25]), .B0(n1718), .S(n1717), .CO(n1716));
Q_AD01HF U2132 ( .A0(aCount[24]), .B0(n1720), .S(n1719), .CO(n1718));
Q_AD01HF U2133 ( .A0(aCount[23]), .B0(n1722), .S(n1721), .CO(n1720));
Q_AD01HF U2134 ( .A0(aCount[22]), .B0(n1724), .S(n1723), .CO(n1722));
Q_AD01HF U2135 ( .A0(aCount[21]), .B0(n1726), .S(n1725), .CO(n1724));
Q_AD01HF U2136 ( .A0(aCount[20]), .B0(n1728), .S(n1727), .CO(n1726));
Q_AD01HF U2137 ( .A0(aCount[19]), .B0(n1730), .S(n1729), .CO(n1728));
Q_AD01HF U2138 ( .A0(aCount[18]), .B0(n1732), .S(n1731), .CO(n1730));
Q_AD01HF U2139 ( .A0(aCount[17]), .B0(n1734), .S(n1733), .CO(n1732));
Q_AD01HF U2140 ( .A0(aCount[16]), .B0(n1736), .S(n1735), .CO(n1734));
Q_AD01HF U2141 ( .A0(aCount[15]), .B0(n1738), .S(n1737), .CO(n1736));
Q_AD01HF U2142 ( .A0(aCount[14]), .B0(n1740), .S(n1739), .CO(n1738));
Q_AD01HF U2143 ( .A0(aCount[13]), .B0(n1742), .S(n1741), .CO(n1740));
Q_AD01HF U2144 ( .A0(aCount[12]), .B0(n1744), .S(n1743), .CO(n1742));
Q_AD01HF U2145 ( .A0(aCount[11]), .B0(n1746), .S(n1745), .CO(n1744));
Q_AD01HF U2146 ( .A0(aCount[10]), .B0(n1748), .S(n1747), .CO(n1746));
Q_AD01HF U2147 ( .A0(aCount[9]), .B0(n1750), .S(n1749), .CO(n1748));
Q_AD01HF U2148 ( .A0(aCount[8]), .B0(n1752), .S(n1751), .CO(n1750));
Q_AD01HF U2149 ( .A0(aCount[7]), .B0(n1754), .S(n1753), .CO(n1752));
Q_AD01HF U2150 ( .A0(aCount[6]), .B0(n1756), .S(n1755), .CO(n1754));
Q_AD01HF U2151 ( .A0(aCount[5]), .B0(n1758), .S(n1757), .CO(n1756));
Q_AD01HF U2152 ( .A0(aCount[4]), .B0(n1760), .S(n1759), .CO(n1758));
Q_AD01HF U2153 ( .A0(aCount[3]), .B0(n1762), .S(n1761), .CO(n1760));
Q_AD01HF U2154 ( .A0(aCount[2]), .B0(n1764), .S(n1763), .CO(n1762));
Q_AD01HF U2155 ( .A0(aCount[1]), .B0(aCount[0]), .S(n1765), .CO(n1764));
Q_INV U2156 ( .A(ixcHoldClkR), .Z(n1767));
Q_AN02 U2157 ( .A0(ixcHoldClk), .A1(n1767), .Z(n1766));
Q_XOR2 U2158 ( .A0(n1766), .A1(ixcHoldSyncCnt[0]), .Z(n1768));
Q_FDP0UA U2159 ( .D(n1768), .QTFCLK( ), .Q(ixcHoldSyncCnt[0]));
Q_MX02 U2160 ( .S(n1766), .A0(ixcHoldSyncCnt[1]), .A1(n1955), .Z(n1769));
Q_FDP0UA U2161 ( .D(n1769), .QTFCLK( ), .Q(ixcHoldSyncCnt[1]));
Q_MX02 U2162 ( .S(n1766), .A0(ixcHoldSyncCnt[2]), .A1(n1953), .Z(n1770));
Q_FDP0UA U2163 ( .D(n1770), .QTFCLK( ), .Q(ixcHoldSyncCnt[2]));
Q_MX02 U2164 ( .S(n1766), .A0(ixcHoldSyncCnt[3]), .A1(n1951), .Z(n1771));
Q_FDP0UA U2165 ( .D(n1771), .QTFCLK( ), .Q(ixcHoldSyncCnt[3]));
Q_MX02 U2166 ( .S(n1766), .A0(ixcHoldSyncCnt[4]), .A1(n1949), .Z(n1772));
Q_FDP0UA U2167 ( .D(n1772), .QTFCLK( ), .Q(ixcHoldSyncCnt[4]));
Q_MX02 U2168 ( .S(n1766), .A0(ixcHoldSyncCnt[5]), .A1(n1947), .Z(n1773));
Q_FDP0UA U2169 ( .D(n1773), .QTFCLK( ), .Q(ixcHoldSyncCnt[5]));
Q_MX02 U2170 ( .S(n1766), .A0(ixcHoldSyncCnt[6]), .A1(n1945), .Z(n1774));
Q_FDP0UA U2171 ( .D(n1774), .QTFCLK( ), .Q(ixcHoldSyncCnt[6]));
Q_MX02 U2172 ( .S(n1766), .A0(ixcHoldSyncCnt[7]), .A1(n1943), .Z(n1775));
Q_FDP0UA U2173 ( .D(n1775), .QTFCLK( ), .Q(ixcHoldSyncCnt[7]));
Q_MX02 U2174 ( .S(n1766), .A0(ixcHoldSyncCnt[8]), .A1(n1941), .Z(n1776));
Q_FDP0UA U2175 ( .D(n1776), .QTFCLK( ), .Q(ixcHoldSyncCnt[8]));
Q_MX02 U2176 ( .S(n1766), .A0(ixcHoldSyncCnt[9]), .A1(n1939), .Z(n1777));
Q_FDP0UA U2177 ( .D(n1777), .QTFCLK( ), .Q(ixcHoldSyncCnt[9]));
Q_MX02 U2178 ( .S(n1766), .A0(ixcHoldSyncCnt[10]), .A1(n1937), .Z(n1778));
Q_FDP0UA U2179 ( .D(n1778), .QTFCLK( ), .Q(ixcHoldSyncCnt[10]));
Q_MX02 U2180 ( .S(n1766), .A0(ixcHoldSyncCnt[11]), .A1(n1935), .Z(n1779));
Q_FDP0UA U2181 ( .D(n1779), .QTFCLK( ), .Q(ixcHoldSyncCnt[11]));
Q_MX02 U2182 ( .S(n1766), .A0(ixcHoldSyncCnt[12]), .A1(n1933), .Z(n1780));
Q_FDP0UA U2183 ( .D(n1780), .QTFCLK( ), .Q(ixcHoldSyncCnt[12]));
Q_MX02 U2184 ( .S(n1766), .A0(ixcHoldSyncCnt[13]), .A1(n1931), .Z(n1781));
Q_FDP0UA U2185 ( .D(n1781), .QTFCLK( ), .Q(ixcHoldSyncCnt[13]));
Q_MX02 U2186 ( .S(n1766), .A0(ixcHoldSyncCnt[14]), .A1(n1929), .Z(n1782));
Q_FDP0UA U2187 ( .D(n1782), .QTFCLK( ), .Q(ixcHoldSyncCnt[14]));
Q_MX02 U2188 ( .S(n1766), .A0(ixcHoldSyncCnt[15]), .A1(n1927), .Z(n1783));
Q_FDP0UA U2189 ( .D(n1783), .QTFCLK( ), .Q(ixcHoldSyncCnt[15]));
Q_MX02 U2190 ( .S(n1766), .A0(ixcHoldSyncCnt[16]), .A1(n1925), .Z(n1784));
Q_FDP0UA U2191 ( .D(n1784), .QTFCLK( ), .Q(ixcHoldSyncCnt[16]));
Q_MX02 U2192 ( .S(n1766), .A0(ixcHoldSyncCnt[17]), .A1(n1923), .Z(n1785));
Q_FDP0UA U2193 ( .D(n1785), .QTFCLK( ), .Q(ixcHoldSyncCnt[17]));
Q_MX02 U2194 ( .S(n1766), .A0(ixcHoldSyncCnt[18]), .A1(n1921), .Z(n1786));
Q_FDP0UA U2195 ( .D(n1786), .QTFCLK( ), .Q(ixcHoldSyncCnt[18]));
Q_MX02 U2196 ( .S(n1766), .A0(ixcHoldSyncCnt[19]), .A1(n1919), .Z(n1787));
Q_FDP0UA U2197 ( .D(n1787), .QTFCLK( ), .Q(ixcHoldSyncCnt[19]));
Q_MX02 U2198 ( .S(n1766), .A0(ixcHoldSyncCnt[20]), .A1(n1917), .Z(n1788));
Q_FDP0UA U2199 ( .D(n1788), .QTFCLK( ), .Q(ixcHoldSyncCnt[20]));
Q_MX02 U2200 ( .S(n1766), .A0(ixcHoldSyncCnt[21]), .A1(n1915), .Z(n1789));
Q_FDP0UA U2201 ( .D(n1789), .QTFCLK( ), .Q(ixcHoldSyncCnt[21]));
Q_MX02 U2202 ( .S(n1766), .A0(ixcHoldSyncCnt[22]), .A1(n1913), .Z(n1790));
Q_FDP0UA U2203 ( .D(n1790), .QTFCLK( ), .Q(ixcHoldSyncCnt[22]));
Q_MX02 U2204 ( .S(n1766), .A0(ixcHoldSyncCnt[23]), .A1(n1911), .Z(n1791));
Q_FDP0UA U2205 ( .D(n1791), .QTFCLK( ), .Q(ixcHoldSyncCnt[23]));
Q_MX02 U2206 ( .S(n1766), .A0(ixcHoldSyncCnt[24]), .A1(n1909), .Z(n1792));
Q_FDP0UA U2207 ( .D(n1792), .QTFCLK( ), .Q(ixcHoldSyncCnt[24]));
Q_MX02 U2208 ( .S(n1766), .A0(ixcHoldSyncCnt[25]), .A1(n1907), .Z(n1793));
Q_FDP0UA U2209 ( .D(n1793), .QTFCLK( ), .Q(ixcHoldSyncCnt[25]));
Q_MX02 U2210 ( .S(n1766), .A0(ixcHoldSyncCnt[26]), .A1(n1905), .Z(n1794));
Q_FDP0UA U2211 ( .D(n1794), .QTFCLK( ), .Q(ixcHoldSyncCnt[26]));
Q_MX02 U2212 ( .S(n1766), .A0(ixcHoldSyncCnt[27]), .A1(n1903), .Z(n1795));
Q_FDP0UA U2213 ( .D(n1795), .QTFCLK( ), .Q(ixcHoldSyncCnt[27]));
Q_MX02 U2214 ( .S(n1766), .A0(ixcHoldSyncCnt[28]), .A1(n1901), .Z(n1796));
Q_FDP0UA U2215 ( .D(n1796), .QTFCLK( ), .Q(ixcHoldSyncCnt[28]));
Q_MX02 U2216 ( .S(n1766), .A0(ixcHoldSyncCnt[29]), .A1(n1899), .Z(n1797));
Q_FDP0UA U2217 ( .D(n1797), .QTFCLK( ), .Q(ixcHoldSyncCnt[29]));
Q_MX02 U2218 ( .S(n1766), .A0(ixcHoldSyncCnt[30]), .A1(n1897), .Z(n1798));
Q_FDP0UA U2219 ( .D(n1798), .QTFCLK( ), .Q(ixcHoldSyncCnt[30]));
Q_MX02 U2220 ( .S(n1766), .A0(ixcHoldSyncCnt[31]), .A1(n1895), .Z(n1799));
Q_FDP0UA U2221 ( .D(n1799), .QTFCLK( ), .Q(ixcHoldSyncCnt[31]));
Q_MX02 U2222 ( .S(n1766), .A0(ixcHoldSyncCnt[32]), .A1(n1893), .Z(n1800));
Q_FDP0UA U2223 ( .D(n1800), .QTFCLK( ), .Q(ixcHoldSyncCnt[32]));
Q_MX02 U2224 ( .S(n1766), .A0(ixcHoldSyncCnt[33]), .A1(n1891), .Z(n1801));
Q_FDP0UA U2225 ( .D(n1801), .QTFCLK( ), .Q(ixcHoldSyncCnt[33]));
Q_MX02 U2226 ( .S(n1766), .A0(ixcHoldSyncCnt[34]), .A1(n1889), .Z(n1802));
Q_FDP0UA U2227 ( .D(n1802), .QTFCLK( ), .Q(ixcHoldSyncCnt[34]));
Q_MX02 U2228 ( .S(n1766), .A0(ixcHoldSyncCnt[35]), .A1(n1887), .Z(n1803));
Q_FDP0UA U2229 ( .D(n1803), .QTFCLK( ), .Q(ixcHoldSyncCnt[35]));
Q_MX02 U2230 ( .S(n1766), .A0(ixcHoldSyncCnt[36]), .A1(n1885), .Z(n1804));
Q_FDP0UA U2231 ( .D(n1804), .QTFCLK( ), .Q(ixcHoldSyncCnt[36]));
Q_MX02 U2232 ( .S(n1766), .A0(ixcHoldSyncCnt[37]), .A1(n1883), .Z(n1805));
Q_FDP0UA U2233 ( .D(n1805), .QTFCLK( ), .Q(ixcHoldSyncCnt[37]));
Q_MX02 U2234 ( .S(n1766), .A0(ixcHoldSyncCnt[38]), .A1(n1881), .Z(n1806));
Q_FDP0UA U2235 ( .D(n1806), .QTFCLK( ), .Q(ixcHoldSyncCnt[38]));
Q_MX02 U2236 ( .S(n1766), .A0(ixcHoldSyncCnt[39]), .A1(n1879), .Z(n1807));
Q_FDP0UA U2237 ( .D(n1807), .QTFCLK( ), .Q(ixcHoldSyncCnt[39]));
Q_MX02 U2238 ( .S(n1766), .A0(ixcHoldSyncCnt[40]), .A1(n1877), .Z(n1808));
Q_FDP0UA U2239 ( .D(n1808), .QTFCLK( ), .Q(ixcHoldSyncCnt[40]));
Q_MX02 U2240 ( .S(n1766), .A0(ixcHoldSyncCnt[41]), .A1(n1875), .Z(n1809));
Q_FDP0UA U2241 ( .D(n1809), .QTFCLK( ), .Q(ixcHoldSyncCnt[41]));
Q_MX02 U2242 ( .S(n1766), .A0(ixcHoldSyncCnt[42]), .A1(n1873), .Z(n1810));
Q_FDP0UA U2243 ( .D(n1810), .QTFCLK( ), .Q(ixcHoldSyncCnt[42]));
Q_MX02 U2244 ( .S(n1766), .A0(ixcHoldSyncCnt[43]), .A1(n1871), .Z(n1811));
Q_FDP0UA U2245 ( .D(n1811), .QTFCLK( ), .Q(ixcHoldSyncCnt[43]));
Q_MX02 U2246 ( .S(n1766), .A0(ixcHoldSyncCnt[44]), .A1(n1869), .Z(n1812));
Q_FDP0UA U2247 ( .D(n1812), .QTFCLK( ), .Q(ixcHoldSyncCnt[44]));
Q_MX02 U2248 ( .S(n1766), .A0(ixcHoldSyncCnt[45]), .A1(n1867), .Z(n1813));
Q_FDP0UA U2249 ( .D(n1813), .QTFCLK( ), .Q(ixcHoldSyncCnt[45]));
Q_MX02 U2250 ( .S(n1766), .A0(ixcHoldSyncCnt[46]), .A1(n1865), .Z(n1814));
Q_FDP0UA U2251 ( .D(n1814), .QTFCLK( ), .Q(ixcHoldSyncCnt[46]));
Q_MX02 U2252 ( .S(n1766), .A0(ixcHoldSyncCnt[47]), .A1(n1863), .Z(n1815));
Q_FDP0UA U2253 ( .D(n1815), .QTFCLK( ), .Q(ixcHoldSyncCnt[47]));
Q_MX02 U2254 ( .S(n1766), .A0(ixcHoldSyncCnt[48]), .A1(n1861), .Z(n1816));
Q_FDP0UA U2255 ( .D(n1816), .QTFCLK( ), .Q(ixcHoldSyncCnt[48]));
Q_MX02 U2256 ( .S(n1766), .A0(ixcHoldSyncCnt[49]), .A1(n1859), .Z(n1817));
Q_FDP0UA U2257 ( .D(n1817), .QTFCLK( ), .Q(ixcHoldSyncCnt[49]));
Q_MX02 U2258 ( .S(n1766), .A0(ixcHoldSyncCnt[50]), .A1(n1857), .Z(n1818));
Q_FDP0UA U2259 ( .D(n1818), .QTFCLK( ), .Q(ixcHoldSyncCnt[50]));
Q_MX02 U2260 ( .S(n1766), .A0(ixcHoldSyncCnt[51]), .A1(n1855), .Z(n1819));
Q_FDP0UA U2261 ( .D(n1819), .QTFCLK( ), .Q(ixcHoldSyncCnt[51]));
Q_MX02 U2262 ( .S(n1766), .A0(ixcHoldSyncCnt[52]), .A1(n1853), .Z(n1820));
Q_FDP0UA U2263 ( .D(n1820), .QTFCLK( ), .Q(ixcHoldSyncCnt[52]));
Q_MX02 U2264 ( .S(n1766), .A0(ixcHoldSyncCnt[53]), .A1(n1851), .Z(n1821));
Q_FDP0UA U2265 ( .D(n1821), .QTFCLK( ), .Q(ixcHoldSyncCnt[53]));
Q_MX02 U2266 ( .S(n1766), .A0(ixcHoldSyncCnt[54]), .A1(n1849), .Z(n1822));
Q_FDP0UA U2267 ( .D(n1822), .QTFCLK( ), .Q(ixcHoldSyncCnt[54]));
Q_MX02 U2268 ( .S(n1766), .A0(ixcHoldSyncCnt[55]), .A1(n1847), .Z(n1823));
Q_FDP0UA U2269 ( .D(n1823), .QTFCLK( ), .Q(ixcHoldSyncCnt[55]));
Q_MX02 U2270 ( .S(n1766), .A0(ixcHoldSyncCnt[56]), .A1(n1845), .Z(n1824));
Q_FDP0UA U2271 ( .D(n1824), .QTFCLK( ), .Q(ixcHoldSyncCnt[56]));
Q_MX02 U2272 ( .S(n1766), .A0(ixcHoldSyncCnt[57]), .A1(n1843), .Z(n1825));
Q_FDP0UA U2273 ( .D(n1825), .QTFCLK( ), .Q(ixcHoldSyncCnt[57]));
Q_MX02 U2274 ( .S(n1766), .A0(ixcHoldSyncCnt[58]), .A1(n1841), .Z(n1826));
Q_FDP0UA U2275 ( .D(n1826), .QTFCLK( ), .Q(ixcHoldSyncCnt[58]));
Q_MX02 U2276 ( .S(n1766), .A0(ixcHoldSyncCnt[59]), .A1(n1839), .Z(n1827));
Q_FDP0UA U2277 ( .D(n1827), .QTFCLK( ), .Q(ixcHoldSyncCnt[59]));
Q_MX02 U2278 ( .S(n1766), .A0(ixcHoldSyncCnt[60]), .A1(n1837), .Z(n1828));
Q_FDP0UA U2279 ( .D(n1828), .QTFCLK( ), .Q(ixcHoldSyncCnt[60]));
Q_MX02 U2280 ( .S(n1766), .A0(ixcHoldSyncCnt[61]), .A1(n1835), .Z(n1829));
Q_FDP0UA U2281 ( .D(n1829), .QTFCLK( ), .Q(ixcHoldSyncCnt[61]));
Q_MX02 U2282 ( .S(n1766), .A0(ixcHoldSyncCnt[62]), .A1(n1833), .Z(n1830));
Q_FDP0UA U2283 ( .D(n1830), .QTFCLK( ), .Q(ixcHoldSyncCnt[62]));
Q_FDP0UA U2284 ( .D(n1831), .QTFCLK( ), .Q(ixcHoldSyncCnt[63]));
Q_XOR2 U2285 ( .A0(ixcHoldSyncCnt[63]), .A1(n8), .Z(n1831));
Q_AD01HF U2286 ( .A0(ixcHoldSyncCnt[62]), .B0(n1834), .S(n1833), .CO(n1832));
Q_AD01HF U2287 ( .A0(ixcHoldSyncCnt[61]), .B0(n1836), .S(n1835), .CO(n1834));
Q_AD01HF U2288 ( .A0(ixcHoldSyncCnt[60]), .B0(n1838), .S(n1837), .CO(n1836));
Q_AD01HF U2289 ( .A0(ixcHoldSyncCnt[59]), .B0(n1840), .S(n1839), .CO(n1838));
Q_AD01HF U2290 ( .A0(ixcHoldSyncCnt[58]), .B0(n1842), .S(n1841), .CO(n1840));
Q_AD01HF U2291 ( .A0(ixcHoldSyncCnt[57]), .B0(n1844), .S(n1843), .CO(n1842));
Q_AD01HF U2292 ( .A0(ixcHoldSyncCnt[56]), .B0(n1846), .S(n1845), .CO(n1844));
Q_AD01HF U2293 ( .A0(ixcHoldSyncCnt[55]), .B0(n1848), .S(n1847), .CO(n1846));
Q_AD01HF U2294 ( .A0(ixcHoldSyncCnt[54]), .B0(n1850), .S(n1849), .CO(n1848));
Q_AD01HF U2295 ( .A0(ixcHoldSyncCnt[53]), .B0(n1852), .S(n1851), .CO(n1850));
Q_AD01HF U2296 ( .A0(ixcHoldSyncCnt[52]), .B0(n1854), .S(n1853), .CO(n1852));
Q_AD01HF U2297 ( .A0(ixcHoldSyncCnt[51]), .B0(n1856), .S(n1855), .CO(n1854));
Q_AD01HF U2298 ( .A0(ixcHoldSyncCnt[50]), .B0(n1858), .S(n1857), .CO(n1856));
Q_AD01HF U2299 ( .A0(ixcHoldSyncCnt[49]), .B0(n1860), .S(n1859), .CO(n1858));
Q_AD01HF U2300 ( .A0(ixcHoldSyncCnt[48]), .B0(n1862), .S(n1861), .CO(n1860));
Q_AD01HF U2301 ( .A0(ixcHoldSyncCnt[47]), .B0(n1864), .S(n1863), .CO(n1862));
Q_AD01HF U2302 ( .A0(ixcHoldSyncCnt[46]), .B0(n1866), .S(n1865), .CO(n1864));
Q_AD01HF U2303 ( .A0(ixcHoldSyncCnt[45]), .B0(n1868), .S(n1867), .CO(n1866));
Q_AD01HF U2304 ( .A0(ixcHoldSyncCnt[44]), .B0(n1870), .S(n1869), .CO(n1868));
Q_AD01HF U2305 ( .A0(ixcHoldSyncCnt[43]), .B0(n1872), .S(n1871), .CO(n1870));
Q_AD01HF U2306 ( .A0(ixcHoldSyncCnt[42]), .B0(n1874), .S(n1873), .CO(n1872));
Q_AD01HF U2307 ( .A0(ixcHoldSyncCnt[41]), .B0(n1876), .S(n1875), .CO(n1874));
Q_AD01HF U2308 ( .A0(ixcHoldSyncCnt[40]), .B0(n1878), .S(n1877), .CO(n1876));
Q_AD01HF U2309 ( .A0(ixcHoldSyncCnt[39]), .B0(n1880), .S(n1879), .CO(n1878));
Q_AD01HF U2310 ( .A0(ixcHoldSyncCnt[38]), .B0(n1882), .S(n1881), .CO(n1880));
Q_AD01HF U2311 ( .A0(ixcHoldSyncCnt[37]), .B0(n1884), .S(n1883), .CO(n1882));
Q_AD01HF U2312 ( .A0(ixcHoldSyncCnt[36]), .B0(n1886), .S(n1885), .CO(n1884));
Q_AD01HF U2313 ( .A0(ixcHoldSyncCnt[35]), .B0(n1888), .S(n1887), .CO(n1886));
Q_AD01HF U2314 ( .A0(ixcHoldSyncCnt[34]), .B0(n1890), .S(n1889), .CO(n1888));
Q_AD01HF U2315 ( .A0(ixcHoldSyncCnt[33]), .B0(n1892), .S(n1891), .CO(n1890));
Q_AD01HF U2316 ( .A0(ixcHoldSyncCnt[32]), .B0(n1894), .S(n1893), .CO(n1892));
Q_AD01HF U2317 ( .A0(ixcHoldSyncCnt[31]), .B0(n1896), .S(n1895), .CO(n1894));
Q_AD01HF U2318 ( .A0(ixcHoldSyncCnt[30]), .B0(n1898), .S(n1897), .CO(n1896));
Q_AD01HF U2319 ( .A0(ixcHoldSyncCnt[29]), .B0(n1900), .S(n1899), .CO(n1898));
Q_AD01HF U2320 ( .A0(ixcHoldSyncCnt[28]), .B0(n1902), .S(n1901), .CO(n1900));
Q_AD01HF U2321 ( .A0(ixcHoldSyncCnt[27]), .B0(n1904), .S(n1903), .CO(n1902));
Q_AD01HF U2322 ( .A0(ixcHoldSyncCnt[26]), .B0(n1906), .S(n1905), .CO(n1904));
Q_AD01HF U2323 ( .A0(ixcHoldSyncCnt[25]), .B0(n1908), .S(n1907), .CO(n1906));
Q_AD01HF U2324 ( .A0(ixcHoldSyncCnt[24]), .B0(n1910), .S(n1909), .CO(n1908));
Q_AD01HF U2325 ( .A0(ixcHoldSyncCnt[23]), .B0(n1912), .S(n1911), .CO(n1910));
Q_AD01HF U2326 ( .A0(ixcHoldSyncCnt[22]), .B0(n1914), .S(n1913), .CO(n1912));
Q_AD01HF U2327 ( .A0(ixcHoldSyncCnt[21]), .B0(n1916), .S(n1915), .CO(n1914));
Q_AD01HF U2328 ( .A0(ixcHoldSyncCnt[20]), .B0(n1918), .S(n1917), .CO(n1916));
Q_AD01HF U2329 ( .A0(ixcHoldSyncCnt[19]), .B0(n1920), .S(n1919), .CO(n1918));
Q_AD01HF U2330 ( .A0(ixcHoldSyncCnt[18]), .B0(n1922), .S(n1921), .CO(n1920));
Q_AD01HF U2331 ( .A0(ixcHoldSyncCnt[17]), .B0(n1924), .S(n1923), .CO(n1922));
Q_AD01HF U2332 ( .A0(ixcHoldSyncCnt[16]), .B0(n1926), .S(n1925), .CO(n1924));
Q_AD01HF U2333 ( .A0(ixcHoldSyncCnt[15]), .B0(n1928), .S(n1927), .CO(n1926));
Q_AD01HF U2334 ( .A0(ixcHoldSyncCnt[14]), .B0(n1930), .S(n1929), .CO(n1928));
Q_AD01HF U2335 ( .A0(ixcHoldSyncCnt[13]), .B0(n1932), .S(n1931), .CO(n1930));
Q_AD01HF U2336 ( .A0(ixcHoldSyncCnt[12]), .B0(n1934), .S(n1933), .CO(n1932));
Q_AD01HF U2337 ( .A0(ixcHoldSyncCnt[11]), .B0(n1936), .S(n1935), .CO(n1934));
Q_AD01HF U2338 ( .A0(ixcHoldSyncCnt[10]), .B0(n1938), .S(n1937), .CO(n1936));
Q_AD01HF U2339 ( .A0(ixcHoldSyncCnt[9]), .B0(n1940), .S(n1939), .CO(n1938));
Q_AD01HF U2340 ( .A0(ixcHoldSyncCnt[8]), .B0(n1942), .S(n1941), .CO(n1940));
Q_AD01HF U2341 ( .A0(ixcHoldSyncCnt[7]), .B0(n1944), .S(n1943), .CO(n1942));
Q_AD01HF U2342 ( .A0(ixcHoldSyncCnt[6]), .B0(n1946), .S(n1945), .CO(n1944));
Q_AD01HF U2343 ( .A0(ixcHoldSyncCnt[5]), .B0(n1948), .S(n1947), .CO(n1946));
Q_AD01HF U2344 ( .A0(ixcHoldSyncCnt[4]), .B0(n1950), .S(n1949), .CO(n1948));
Q_AD01HF U2345 ( .A0(ixcHoldSyncCnt[3]), .B0(n1952), .S(n1951), .CO(n1950));
Q_AD01HF U2346 ( .A0(ixcHoldSyncCnt[2]), .B0(n1954), .S(n1953), .CO(n1952));
Q_AD01HF U2347 ( .A0(ixcHoldSyncCnt[1]), .B0(ixcHoldSyncCnt[0]), .S(n1955), .CO(n1954));
Q_FDP0UA U2348 ( .D(ixcHoldClk), .QTFCLK( ), .Q(ixcHoldClkR));
Q_NR02 U2349 ( .A0(sampleXpChg), .A1(n401), .Z(n1959));
Q_OR02 U2350 ( .A0(GFBw), .A1(n1959), .Z(n1965));
Q_INV U2351 ( .A(ixcHoldClk), .Z(n1960));
Q_OR02 U2352 ( .A0(n1960), .A1(n1965), .Z(n1961));
Q_INV U2353 ( .A(n1961), .Z(n1956));
Q_INV U2354 ( .A(sampleXpChg), .Z(n1962));
Q_OR02 U2355 ( .A0(n1962), .A1(bpWait), .Z(n1963));
Q_OR02 U2356 ( .A0(GFBw), .A1(n1963), .Z(n1964));
Q_INV U2357 ( .A(n1964), .Z(n1957));
Q_INV U2358 ( .A(n1965), .Z(n1958));
Q_XOR2 U2359 ( .A0(n1956), .A1(ixcHoldClkCnt[0]), .Z(n1966));
Q_FDP0UA U2360 ( .D(n1966), .QTFCLK( ), .Q(ixcHoldClkCnt[0]));
Q_MX02 U2361 ( .S(n1961), .A0(n2281), .A1(ixcHoldClkCnt[1]), .Z(n1967));
Q_FDP0UA U2362 ( .D(n1967), .QTFCLK( ), .Q(ixcHoldClkCnt[1]));
Q_MX02 U2363 ( .S(n1961), .A0(n2279), .A1(ixcHoldClkCnt[2]), .Z(n1968));
Q_FDP0UA U2364 ( .D(n1968), .QTFCLK( ), .Q(ixcHoldClkCnt[2]));
Q_MX02 U2365 ( .S(n1961), .A0(n2277), .A1(ixcHoldClkCnt[3]), .Z(n1969));
Q_FDP0UA U2366 ( .D(n1969), .QTFCLK( ), .Q(ixcHoldClkCnt[3]));
Q_MX02 U2367 ( .S(n1961), .A0(n2275), .A1(ixcHoldClkCnt[4]), .Z(n1970));
Q_FDP0UA U2368 ( .D(n1970), .QTFCLK( ), .Q(ixcHoldClkCnt[4]));
Q_MX02 U2369 ( .S(n1961), .A0(n2273), .A1(ixcHoldClkCnt[5]), .Z(n1971));
Q_FDP0UA U2370 ( .D(n1971), .QTFCLK( ), .Q(ixcHoldClkCnt[5]));
Q_MX02 U2371 ( .S(n1961), .A0(n2271), .A1(ixcHoldClkCnt[6]), .Z(n1972));
Q_FDP0UA U2372 ( .D(n1972), .QTFCLK( ), .Q(ixcHoldClkCnt[6]));
Q_MX02 U2373 ( .S(n1961), .A0(n2269), .A1(ixcHoldClkCnt[7]), .Z(n1973));
Q_FDP0UA U2374 ( .D(n1973), .QTFCLK( ), .Q(ixcHoldClkCnt[7]));
Q_MX02 U2375 ( .S(n1961), .A0(n2267), .A1(ixcHoldClkCnt[8]), .Z(n1974));
Q_FDP0UA U2376 ( .D(n1974), .QTFCLK( ), .Q(ixcHoldClkCnt[8]));
Q_MX02 U2377 ( .S(n1961), .A0(n2265), .A1(ixcHoldClkCnt[9]), .Z(n1975));
Q_FDP0UA U2378 ( .D(n1975), .QTFCLK( ), .Q(ixcHoldClkCnt[9]));
Q_MX02 U2379 ( .S(n1961), .A0(n2263), .A1(ixcHoldClkCnt[10]), .Z(n1976));
Q_FDP0UA U2380 ( .D(n1976), .QTFCLK( ), .Q(ixcHoldClkCnt[10]));
Q_MX02 U2381 ( .S(n1961), .A0(n2261), .A1(ixcHoldClkCnt[11]), .Z(n1977));
Q_FDP0UA U2382 ( .D(n1977), .QTFCLK( ), .Q(ixcHoldClkCnt[11]));
Q_MX02 U2383 ( .S(n1961), .A0(n2259), .A1(ixcHoldClkCnt[12]), .Z(n1978));
Q_FDP0UA U2384 ( .D(n1978), .QTFCLK( ), .Q(ixcHoldClkCnt[12]));
Q_MX02 U2385 ( .S(n1961), .A0(n2257), .A1(ixcHoldClkCnt[13]), .Z(n1979));
Q_FDP0UA U2386 ( .D(n1979), .QTFCLK( ), .Q(ixcHoldClkCnt[13]));
Q_MX02 U2387 ( .S(n1961), .A0(n2255), .A1(ixcHoldClkCnt[14]), .Z(n1980));
Q_FDP0UA U2388 ( .D(n1980), .QTFCLK( ), .Q(ixcHoldClkCnt[14]));
Q_MX02 U2389 ( .S(n1961), .A0(n2253), .A1(ixcHoldClkCnt[15]), .Z(n1981));
Q_FDP0UA U2390 ( .D(n1981), .QTFCLK( ), .Q(ixcHoldClkCnt[15]));
Q_MX02 U2391 ( .S(n1961), .A0(n2251), .A1(ixcHoldClkCnt[16]), .Z(n1982));
Q_FDP0UA U2392 ( .D(n1982), .QTFCLK( ), .Q(ixcHoldClkCnt[16]));
Q_MX02 U2393 ( .S(n1961), .A0(n2249), .A1(ixcHoldClkCnt[17]), .Z(n1983));
Q_FDP0UA U2394 ( .D(n1983), .QTFCLK( ), .Q(ixcHoldClkCnt[17]));
Q_MX02 U2395 ( .S(n1961), .A0(n2247), .A1(ixcHoldClkCnt[18]), .Z(n1984));
Q_FDP0UA U2396 ( .D(n1984), .QTFCLK( ), .Q(ixcHoldClkCnt[18]));
Q_MX02 U2397 ( .S(n1961), .A0(n2245), .A1(ixcHoldClkCnt[19]), .Z(n1985));
Q_FDP0UA U2398 ( .D(n1985), .QTFCLK( ), .Q(ixcHoldClkCnt[19]));
Q_MX02 U2399 ( .S(n1961), .A0(n2243), .A1(ixcHoldClkCnt[20]), .Z(n1986));
Q_FDP0UA U2400 ( .D(n1986), .QTFCLK( ), .Q(ixcHoldClkCnt[20]));
Q_MX02 U2401 ( .S(n1961), .A0(n2241), .A1(ixcHoldClkCnt[21]), .Z(n1987));
Q_FDP0UA U2402 ( .D(n1987), .QTFCLK( ), .Q(ixcHoldClkCnt[21]));
Q_MX02 U2403 ( .S(n1961), .A0(n2239), .A1(ixcHoldClkCnt[22]), .Z(n1988));
Q_FDP0UA U2404 ( .D(n1988), .QTFCLK( ), .Q(ixcHoldClkCnt[22]));
Q_MX02 U2405 ( .S(n1961), .A0(n2237), .A1(ixcHoldClkCnt[23]), .Z(n1989));
Q_FDP0UA U2406 ( .D(n1989), .QTFCLK( ), .Q(ixcHoldClkCnt[23]));
Q_MX02 U2407 ( .S(n1961), .A0(n2235), .A1(ixcHoldClkCnt[24]), .Z(n1990));
Q_FDP0UA U2408 ( .D(n1990), .QTFCLK( ), .Q(ixcHoldClkCnt[24]));
Q_MX02 U2409 ( .S(n1961), .A0(n2233), .A1(ixcHoldClkCnt[25]), .Z(n1991));
Q_FDP0UA U2410 ( .D(n1991), .QTFCLK( ), .Q(ixcHoldClkCnt[25]));
Q_MX02 U2411 ( .S(n1961), .A0(n2231), .A1(ixcHoldClkCnt[26]), .Z(n1992));
Q_FDP0UA U2412 ( .D(n1992), .QTFCLK( ), .Q(ixcHoldClkCnt[26]));
Q_MX02 U2413 ( .S(n1961), .A0(n2229), .A1(ixcHoldClkCnt[27]), .Z(n1993));
Q_FDP0UA U2414 ( .D(n1993), .QTFCLK( ), .Q(ixcHoldClkCnt[27]));
Q_MX02 U2415 ( .S(n1961), .A0(n2227), .A1(ixcHoldClkCnt[28]), .Z(n1994));
Q_FDP0UA U2416 ( .D(n1994), .QTFCLK( ), .Q(ixcHoldClkCnt[28]));
Q_MX02 U2417 ( .S(n1961), .A0(n2225), .A1(ixcHoldClkCnt[29]), .Z(n1995));
Q_FDP0UA U2418 ( .D(n1995), .QTFCLK( ), .Q(ixcHoldClkCnt[29]));
Q_MX02 U2419 ( .S(n1961), .A0(n2223), .A1(ixcHoldClkCnt[30]), .Z(n1996));
Q_FDP0UA U2420 ( .D(n1996), .QTFCLK( ), .Q(ixcHoldClkCnt[30]));
Q_MX02 U2421 ( .S(n1961), .A0(n2221), .A1(ixcHoldClkCnt[31]), .Z(n1997));
Q_FDP0UA U2422 ( .D(n1997), .QTFCLK( ), .Q(ixcHoldClkCnt[31]));
Q_MX02 U2423 ( .S(n1961), .A0(n2219), .A1(ixcHoldClkCnt[32]), .Z(n1998));
Q_FDP0UA U2424 ( .D(n1998), .QTFCLK( ), .Q(ixcHoldClkCnt[32]));
Q_MX02 U2425 ( .S(n1961), .A0(n2217), .A1(ixcHoldClkCnt[33]), .Z(n1999));
Q_FDP0UA U2426 ( .D(n1999), .QTFCLK( ), .Q(ixcHoldClkCnt[33]));
Q_MX02 U2427 ( .S(n1961), .A0(n2215), .A1(ixcHoldClkCnt[34]), .Z(n2000));
Q_FDP0UA U2428 ( .D(n2000), .QTFCLK( ), .Q(ixcHoldClkCnt[34]));
Q_MX02 U2429 ( .S(n1961), .A0(n2213), .A1(ixcHoldClkCnt[35]), .Z(n2001));
Q_FDP0UA U2430 ( .D(n2001), .QTFCLK( ), .Q(ixcHoldClkCnt[35]));
Q_MX02 U2431 ( .S(n1961), .A0(n2211), .A1(ixcHoldClkCnt[36]), .Z(n2002));
Q_FDP0UA U2432 ( .D(n2002), .QTFCLK( ), .Q(ixcHoldClkCnt[36]));
Q_MX02 U2433 ( .S(n1961), .A0(n2209), .A1(ixcHoldClkCnt[37]), .Z(n2003));
Q_FDP0UA U2434 ( .D(n2003), .QTFCLK( ), .Q(ixcHoldClkCnt[37]));
Q_MX02 U2435 ( .S(n1961), .A0(n2207), .A1(ixcHoldClkCnt[38]), .Z(n2004));
Q_FDP0UA U2436 ( .D(n2004), .QTFCLK( ), .Q(ixcHoldClkCnt[38]));
Q_MX02 U2437 ( .S(n1961), .A0(n2205), .A1(ixcHoldClkCnt[39]), .Z(n2005));
Q_FDP0UA U2438 ( .D(n2005), .QTFCLK( ), .Q(ixcHoldClkCnt[39]));
Q_MX02 U2439 ( .S(n1961), .A0(n2203), .A1(ixcHoldClkCnt[40]), .Z(n2006));
Q_FDP0UA U2440 ( .D(n2006), .QTFCLK( ), .Q(ixcHoldClkCnt[40]));
Q_MX02 U2441 ( .S(n1961), .A0(n2201), .A1(ixcHoldClkCnt[41]), .Z(n2007));
Q_FDP0UA U2442 ( .D(n2007), .QTFCLK( ), .Q(ixcHoldClkCnt[41]));
Q_MX02 U2443 ( .S(n1961), .A0(n2199), .A1(ixcHoldClkCnt[42]), .Z(n2008));
Q_FDP0UA U2444 ( .D(n2008), .QTFCLK( ), .Q(ixcHoldClkCnt[42]));
Q_MX02 U2445 ( .S(n1961), .A0(n2197), .A1(ixcHoldClkCnt[43]), .Z(n2009));
Q_FDP0UA U2446 ( .D(n2009), .QTFCLK( ), .Q(ixcHoldClkCnt[43]));
Q_MX02 U2447 ( .S(n1961), .A0(n2195), .A1(ixcHoldClkCnt[44]), .Z(n2010));
Q_FDP0UA U2448 ( .D(n2010), .QTFCLK( ), .Q(ixcHoldClkCnt[44]));
Q_MX02 U2449 ( .S(n1961), .A0(n2193), .A1(ixcHoldClkCnt[45]), .Z(n2011));
Q_FDP0UA U2450 ( .D(n2011), .QTFCLK( ), .Q(ixcHoldClkCnt[45]));
Q_MX02 U2451 ( .S(n1961), .A0(n2191), .A1(ixcHoldClkCnt[46]), .Z(n2012));
Q_FDP0UA U2452 ( .D(n2012), .QTFCLK( ), .Q(ixcHoldClkCnt[46]));
Q_MX02 U2453 ( .S(n1961), .A0(n2189), .A1(ixcHoldClkCnt[47]), .Z(n2013));
Q_FDP0UA U2454 ( .D(n2013), .QTFCLK( ), .Q(ixcHoldClkCnt[47]));
Q_MX02 U2455 ( .S(n1961), .A0(n2187), .A1(ixcHoldClkCnt[48]), .Z(n2014));
Q_FDP0UA U2456 ( .D(n2014), .QTFCLK( ), .Q(ixcHoldClkCnt[48]));
Q_MX02 U2457 ( .S(n1961), .A0(n2185), .A1(ixcHoldClkCnt[49]), .Z(n2015));
Q_FDP0UA U2458 ( .D(n2015), .QTFCLK( ), .Q(ixcHoldClkCnt[49]));
Q_MX02 U2459 ( .S(n1961), .A0(n2183), .A1(ixcHoldClkCnt[50]), .Z(n2016));
Q_FDP0UA U2460 ( .D(n2016), .QTFCLK( ), .Q(ixcHoldClkCnt[50]));
Q_MX02 U2461 ( .S(n1961), .A0(n2181), .A1(ixcHoldClkCnt[51]), .Z(n2017));
Q_FDP0UA U2462 ( .D(n2017), .QTFCLK( ), .Q(ixcHoldClkCnt[51]));
Q_MX02 U2463 ( .S(n1961), .A0(n2179), .A1(ixcHoldClkCnt[52]), .Z(n2018));
Q_FDP0UA U2464 ( .D(n2018), .QTFCLK( ), .Q(ixcHoldClkCnt[52]));
Q_MX02 U2465 ( .S(n1961), .A0(n2177), .A1(ixcHoldClkCnt[53]), .Z(n2019));
Q_FDP0UA U2466 ( .D(n2019), .QTFCLK( ), .Q(ixcHoldClkCnt[53]));
Q_MX02 U2467 ( .S(n1961), .A0(n2175), .A1(ixcHoldClkCnt[54]), .Z(n2020));
Q_FDP0UA U2468 ( .D(n2020), .QTFCLK( ), .Q(ixcHoldClkCnt[54]));
Q_MX02 U2469 ( .S(n1961), .A0(n2173), .A1(ixcHoldClkCnt[55]), .Z(n2021));
Q_FDP0UA U2470 ( .D(n2021), .QTFCLK( ), .Q(ixcHoldClkCnt[55]));
Q_MX02 U2471 ( .S(n1961), .A0(n2171), .A1(ixcHoldClkCnt[56]), .Z(n2022));
Q_FDP0UA U2472 ( .D(n2022), .QTFCLK( ), .Q(ixcHoldClkCnt[56]));
Q_MX02 U2473 ( .S(n1961), .A0(n2169), .A1(ixcHoldClkCnt[57]), .Z(n2023));
Q_FDP0UA U2474 ( .D(n2023), .QTFCLK( ), .Q(ixcHoldClkCnt[57]));
Q_MX02 U2475 ( .S(n1961), .A0(n2167), .A1(ixcHoldClkCnt[58]), .Z(n2024));
Q_FDP0UA U2476 ( .D(n2024), .QTFCLK( ), .Q(ixcHoldClkCnt[58]));
Q_MX02 U2477 ( .S(n1961), .A0(n2165), .A1(ixcHoldClkCnt[59]), .Z(n2025));
Q_FDP0UA U2478 ( .D(n2025), .QTFCLK( ), .Q(ixcHoldClkCnt[59]));
Q_MX02 U2479 ( .S(n1961), .A0(n2163), .A1(ixcHoldClkCnt[60]), .Z(n2026));
Q_FDP0UA U2480 ( .D(n2026), .QTFCLK( ), .Q(ixcHoldClkCnt[60]));
Q_MX02 U2481 ( .S(n1961), .A0(n2161), .A1(ixcHoldClkCnt[61]), .Z(n2027));
Q_FDP0UA U2482 ( .D(n2027), .QTFCLK( ), .Q(ixcHoldClkCnt[61]));
Q_MX02 U2483 ( .S(n1961), .A0(n2159), .A1(ixcHoldClkCnt[62]), .Z(n2028));
Q_FDP0UA U2484 ( .D(n2028), .QTFCLK( ), .Q(ixcHoldClkCnt[62]));
Q_FDP0UA U2485 ( .D(n2029), .QTFCLK( ), .Q(ixcHoldClkCnt[63]));
Q_XOR2 U2486 ( .A0(n1957), .A1(nbaCount[0]), .Z(n2030));
Q_FDP0UA U2487 ( .D(n2030), .QTFCLK( ), .Q(nbaCount[0]));
Q_MX02 U2488 ( .S(n1964), .A0(n2405), .A1(nbaCount[1]), .Z(n2031));
Q_FDP0UA U2489 ( .D(n2031), .QTFCLK( ), .Q(nbaCount[1]));
Q_MX02 U2490 ( .S(n1964), .A0(n2403), .A1(nbaCount[2]), .Z(n2032));
Q_FDP0UA U2491 ( .D(n2032), .QTFCLK( ), .Q(nbaCount[2]));
Q_MX02 U2492 ( .S(n1964), .A0(n2401), .A1(nbaCount[3]), .Z(n2033));
Q_FDP0UA U2493 ( .D(n2033), .QTFCLK( ), .Q(nbaCount[3]));
Q_MX02 U2494 ( .S(n1964), .A0(n2399), .A1(nbaCount[4]), .Z(n2034));
Q_FDP0UA U2495 ( .D(n2034), .QTFCLK( ), .Q(nbaCount[4]));
Q_MX02 U2496 ( .S(n1964), .A0(n2397), .A1(nbaCount[5]), .Z(n2035));
Q_FDP0UA U2497 ( .D(n2035), .QTFCLK( ), .Q(nbaCount[5]));
Q_MX02 U2498 ( .S(n1964), .A0(n2395), .A1(nbaCount[6]), .Z(n2036));
Q_FDP0UA U2499 ( .D(n2036), .QTFCLK( ), .Q(nbaCount[6]));
Q_MX02 U2500 ( .S(n1964), .A0(n2393), .A1(nbaCount[7]), .Z(n2037));
Q_FDP0UA U2501 ( .D(n2037), .QTFCLK( ), .Q(nbaCount[7]));
Q_MX02 U2502 ( .S(n1964), .A0(n2391), .A1(nbaCount[8]), .Z(n2038));
Q_FDP0UA U2503 ( .D(n2038), .QTFCLK( ), .Q(nbaCount[8]));
Q_MX02 U2504 ( .S(n1964), .A0(n2389), .A1(nbaCount[9]), .Z(n2039));
Q_FDP0UA U2505 ( .D(n2039), .QTFCLK( ), .Q(nbaCount[9]));
Q_MX02 U2506 ( .S(n1964), .A0(n2387), .A1(nbaCount[10]), .Z(n2040));
Q_FDP0UA U2507 ( .D(n2040), .QTFCLK( ), .Q(nbaCount[10]));
Q_MX02 U2508 ( .S(n1964), .A0(n2385), .A1(nbaCount[11]), .Z(n2041));
Q_FDP0UA U2509 ( .D(n2041), .QTFCLK( ), .Q(nbaCount[11]));
Q_MX02 U2510 ( .S(n1964), .A0(n2383), .A1(nbaCount[12]), .Z(n2042));
Q_FDP0UA U2511 ( .D(n2042), .QTFCLK( ), .Q(nbaCount[12]));
Q_MX02 U2512 ( .S(n1964), .A0(n2381), .A1(nbaCount[13]), .Z(n2043));
Q_FDP0UA U2513 ( .D(n2043), .QTFCLK( ), .Q(nbaCount[13]));
Q_MX02 U2514 ( .S(n1964), .A0(n2379), .A1(nbaCount[14]), .Z(n2044));
Q_FDP0UA U2515 ( .D(n2044), .QTFCLK( ), .Q(nbaCount[14]));
Q_MX02 U2516 ( .S(n1964), .A0(n2377), .A1(nbaCount[15]), .Z(n2045));
Q_FDP0UA U2517 ( .D(n2045), .QTFCLK( ), .Q(nbaCount[15]));
Q_MX02 U2518 ( .S(n1964), .A0(n2375), .A1(nbaCount[16]), .Z(n2046));
Q_FDP0UA U2519 ( .D(n2046), .QTFCLK( ), .Q(nbaCount[16]));
Q_MX02 U2520 ( .S(n1964), .A0(n2373), .A1(nbaCount[17]), .Z(n2047));
Q_FDP0UA U2521 ( .D(n2047), .QTFCLK( ), .Q(nbaCount[17]));
Q_MX02 U2522 ( .S(n1964), .A0(n2371), .A1(nbaCount[18]), .Z(n2048));
Q_FDP0UA U2523 ( .D(n2048), .QTFCLK( ), .Q(nbaCount[18]));
Q_MX02 U2524 ( .S(n1964), .A0(n2369), .A1(nbaCount[19]), .Z(n2049));
Q_FDP0UA U2525 ( .D(n2049), .QTFCLK( ), .Q(nbaCount[19]));
Q_MX02 U2526 ( .S(n1964), .A0(n2367), .A1(nbaCount[20]), .Z(n2050));
Q_FDP0UA U2527 ( .D(n2050), .QTFCLK( ), .Q(nbaCount[20]));
Q_MX02 U2528 ( .S(n1964), .A0(n2365), .A1(nbaCount[21]), .Z(n2051));
Q_FDP0UA U2529 ( .D(n2051), .QTFCLK( ), .Q(nbaCount[21]));
Q_MX02 U2530 ( .S(n1964), .A0(n2363), .A1(nbaCount[22]), .Z(n2052));
Q_FDP0UA U2531 ( .D(n2052), .QTFCLK( ), .Q(nbaCount[22]));
Q_MX02 U2532 ( .S(n1964), .A0(n2361), .A1(nbaCount[23]), .Z(n2053));
Q_FDP0UA U2533 ( .D(n2053), .QTFCLK( ), .Q(nbaCount[23]));
Q_MX02 U2534 ( .S(n1964), .A0(n2359), .A1(nbaCount[24]), .Z(n2054));
Q_FDP0UA U2535 ( .D(n2054), .QTFCLK( ), .Q(nbaCount[24]));
Q_MX02 U2536 ( .S(n1964), .A0(n2357), .A1(nbaCount[25]), .Z(n2055));
Q_FDP0UA U2537 ( .D(n2055), .QTFCLK( ), .Q(nbaCount[25]));
Q_MX02 U2538 ( .S(n1964), .A0(n2355), .A1(nbaCount[26]), .Z(n2056));
Q_FDP0UA U2539 ( .D(n2056), .QTFCLK( ), .Q(nbaCount[26]));
Q_MX02 U2540 ( .S(n1964), .A0(n2353), .A1(nbaCount[27]), .Z(n2057));
Q_FDP0UA U2541 ( .D(n2057), .QTFCLK( ), .Q(nbaCount[27]));
Q_MX02 U2542 ( .S(n1964), .A0(n2351), .A1(nbaCount[28]), .Z(n2058));
Q_FDP0UA U2543 ( .D(n2058), .QTFCLK( ), .Q(nbaCount[28]));
Q_MX02 U2544 ( .S(n1964), .A0(n2349), .A1(nbaCount[29]), .Z(n2059));
Q_FDP0UA U2545 ( .D(n2059), .QTFCLK( ), .Q(nbaCount[29]));
Q_MX02 U2546 ( .S(n1964), .A0(n2347), .A1(nbaCount[30]), .Z(n2060));
Q_FDP0UA U2547 ( .D(n2060), .QTFCLK( ), .Q(nbaCount[30]));
Q_MX02 U2548 ( .S(n1964), .A0(n2345), .A1(nbaCount[31]), .Z(n2061));
Q_FDP0UA U2549 ( .D(n2061), .QTFCLK( ), .Q(nbaCount[31]));
Q_MX02 U2550 ( .S(n1964), .A0(n2343), .A1(nbaCount[32]), .Z(n2062));
Q_FDP0UA U2551 ( .D(n2062), .QTFCLK( ), .Q(nbaCount[32]));
Q_MX02 U2552 ( .S(n1964), .A0(n2341), .A1(nbaCount[33]), .Z(n2063));
Q_FDP0UA U2553 ( .D(n2063), .QTFCLK( ), .Q(nbaCount[33]));
Q_MX02 U2554 ( .S(n1964), .A0(n2339), .A1(nbaCount[34]), .Z(n2064));
Q_FDP0UA U2555 ( .D(n2064), .QTFCLK( ), .Q(nbaCount[34]));
Q_MX02 U2556 ( .S(n1964), .A0(n2337), .A1(nbaCount[35]), .Z(n2065));
Q_FDP0UA U2557 ( .D(n2065), .QTFCLK( ), .Q(nbaCount[35]));
Q_MX02 U2558 ( .S(n1964), .A0(n2335), .A1(nbaCount[36]), .Z(n2066));
Q_FDP0UA U2559 ( .D(n2066), .QTFCLK( ), .Q(nbaCount[36]));
Q_MX02 U2560 ( .S(n1964), .A0(n2333), .A1(nbaCount[37]), .Z(n2067));
Q_FDP0UA U2561 ( .D(n2067), .QTFCLK( ), .Q(nbaCount[37]));
Q_MX02 U2562 ( .S(n1964), .A0(n2331), .A1(nbaCount[38]), .Z(n2068));
Q_FDP0UA U2563 ( .D(n2068), .QTFCLK( ), .Q(nbaCount[38]));
Q_MX02 U2564 ( .S(n1964), .A0(n2329), .A1(nbaCount[39]), .Z(n2069));
Q_FDP0UA U2565 ( .D(n2069), .QTFCLK( ), .Q(nbaCount[39]));
Q_MX02 U2566 ( .S(n1964), .A0(n2327), .A1(nbaCount[40]), .Z(n2070));
Q_FDP0UA U2567 ( .D(n2070), .QTFCLK( ), .Q(nbaCount[40]));
Q_MX02 U2568 ( .S(n1964), .A0(n2325), .A1(nbaCount[41]), .Z(n2071));
Q_FDP0UA U2569 ( .D(n2071), .QTFCLK( ), .Q(nbaCount[41]));
Q_MX02 U2570 ( .S(n1964), .A0(n2323), .A1(nbaCount[42]), .Z(n2072));
Q_FDP0UA U2571 ( .D(n2072), .QTFCLK( ), .Q(nbaCount[42]));
Q_MX02 U2572 ( .S(n1964), .A0(n2321), .A1(nbaCount[43]), .Z(n2073));
Q_FDP0UA U2573 ( .D(n2073), .QTFCLK( ), .Q(nbaCount[43]));
Q_MX02 U2574 ( .S(n1964), .A0(n2319), .A1(nbaCount[44]), .Z(n2074));
Q_FDP0UA U2575 ( .D(n2074), .QTFCLK( ), .Q(nbaCount[44]));
Q_MX02 U2576 ( .S(n1964), .A0(n2317), .A1(nbaCount[45]), .Z(n2075));
Q_FDP0UA U2577 ( .D(n2075), .QTFCLK( ), .Q(nbaCount[45]));
Q_MX02 U2578 ( .S(n1964), .A0(n2315), .A1(nbaCount[46]), .Z(n2076));
Q_FDP0UA U2579 ( .D(n2076), .QTFCLK( ), .Q(nbaCount[46]));
Q_MX02 U2580 ( .S(n1964), .A0(n2313), .A1(nbaCount[47]), .Z(n2077));
Q_FDP0UA U2581 ( .D(n2077), .QTFCLK( ), .Q(nbaCount[47]));
Q_MX02 U2582 ( .S(n1964), .A0(n2311), .A1(nbaCount[48]), .Z(n2078));
Q_FDP0UA U2583 ( .D(n2078), .QTFCLK( ), .Q(nbaCount[48]));
Q_MX02 U2584 ( .S(n1964), .A0(n2309), .A1(nbaCount[49]), .Z(n2079));
Q_FDP0UA U2585 ( .D(n2079), .QTFCLK( ), .Q(nbaCount[49]));
Q_MX02 U2586 ( .S(n1964), .A0(n2307), .A1(nbaCount[50]), .Z(n2080));
Q_FDP0UA U2587 ( .D(n2080), .QTFCLK( ), .Q(nbaCount[50]));
Q_MX02 U2588 ( .S(n1964), .A0(n2305), .A1(nbaCount[51]), .Z(n2081));
Q_FDP0UA U2589 ( .D(n2081), .QTFCLK( ), .Q(nbaCount[51]));
Q_MX02 U2590 ( .S(n1964), .A0(n2303), .A1(nbaCount[52]), .Z(n2082));
Q_FDP0UA U2591 ( .D(n2082), .QTFCLK( ), .Q(nbaCount[52]));
Q_MX02 U2592 ( .S(n1964), .A0(n2301), .A1(nbaCount[53]), .Z(n2083));
Q_FDP0UA U2593 ( .D(n2083), .QTFCLK( ), .Q(nbaCount[53]));
Q_MX02 U2594 ( .S(n1964), .A0(n2299), .A1(nbaCount[54]), .Z(n2084));
Q_FDP0UA U2595 ( .D(n2084), .QTFCLK( ), .Q(nbaCount[54]));
Q_MX02 U2596 ( .S(n1964), .A0(n2297), .A1(nbaCount[55]), .Z(n2085));
Q_FDP0UA U2597 ( .D(n2085), .QTFCLK( ), .Q(nbaCount[55]));
Q_MX02 U2598 ( .S(n1964), .A0(n2295), .A1(nbaCount[56]), .Z(n2086));
Q_FDP0UA U2599 ( .D(n2086), .QTFCLK( ), .Q(nbaCount[56]));
Q_MX02 U2600 ( .S(n1964), .A0(n2293), .A1(nbaCount[57]), .Z(n2087));
Q_FDP0UA U2601 ( .D(n2087), .QTFCLK( ), .Q(nbaCount[57]));
Q_MX02 U2602 ( .S(n1964), .A0(n2291), .A1(nbaCount[58]), .Z(n2088));
Q_FDP0UA U2603 ( .D(n2088), .QTFCLK( ), .Q(nbaCount[58]));
Q_MX02 U2604 ( .S(n1964), .A0(n2289), .A1(nbaCount[59]), .Z(n2089));
Q_FDP0UA U2605 ( .D(n2089), .QTFCLK( ), .Q(nbaCount[59]));
Q_MX02 U2606 ( .S(n1964), .A0(n2287), .A1(nbaCount[60]), .Z(n2090));
Q_FDP0UA U2607 ( .D(n2090), .QTFCLK( ), .Q(nbaCount[60]));
Q_MX02 U2608 ( .S(n1964), .A0(n2285), .A1(nbaCount[61]), .Z(n2091));
Q_FDP0UA U2609 ( .D(n2091), .QTFCLK( ), .Q(nbaCount[61]));
Q_MX02 U2610 ( .S(n1964), .A0(n2283), .A1(nbaCount[62]), .Z(n2092));
Q_FDP0UA U2611 ( .D(n2092), .QTFCLK( ), .Q(nbaCount[62]));
Q_FDP0UA U2612 ( .D(n2093), .QTFCLK( ), .Q(nbaCount[63]));
Q_XOR2 U2613 ( .A0(n1958), .A1(bCount[0]), .Z(n2094));
Q_FDP0UA U2614 ( .D(n2094), .QTFCLK( ), .Q(bCount[0]));
Q_MX02 U2615 ( .S(n1965), .A0(n2529), .A1(bCount[1]), .Z(n2095));
Q_FDP0UA U2616 ( .D(n2095), .QTFCLK( ), .Q(bCount[1]));
Q_MX02 U2617 ( .S(n1965), .A0(n2527), .A1(bCount[2]), .Z(n2096));
Q_FDP0UA U2618 ( .D(n2096), .QTFCLK( ), .Q(bCount[2]));
Q_MX02 U2619 ( .S(n1965), .A0(n2525), .A1(bCount[3]), .Z(n2097));
Q_FDP0UA U2620 ( .D(n2097), .QTFCLK( ), .Q(bCount[3]));
Q_MX02 U2621 ( .S(n1965), .A0(n2523), .A1(bCount[4]), .Z(n2098));
Q_FDP0UA U2622 ( .D(n2098), .QTFCLK( ), .Q(bCount[4]));
Q_MX02 U2623 ( .S(n1965), .A0(n2521), .A1(bCount[5]), .Z(n2099));
Q_FDP0UA U2624 ( .D(n2099), .QTFCLK( ), .Q(bCount[5]));
Q_MX02 U2625 ( .S(n1965), .A0(n2519), .A1(bCount[6]), .Z(n2100));
Q_FDP0UA U2626 ( .D(n2100), .QTFCLK( ), .Q(bCount[6]));
Q_MX02 U2627 ( .S(n1965), .A0(n2517), .A1(bCount[7]), .Z(n2101));
Q_FDP0UA U2628 ( .D(n2101), .QTFCLK( ), .Q(bCount[7]));
Q_MX02 U2629 ( .S(n1965), .A0(n2515), .A1(bCount[8]), .Z(n2102));
Q_FDP0UA U2630 ( .D(n2102), .QTFCLK( ), .Q(bCount[8]));
Q_MX02 U2631 ( .S(n1965), .A0(n2513), .A1(bCount[9]), .Z(n2103));
Q_FDP0UA U2632 ( .D(n2103), .QTFCLK( ), .Q(bCount[9]));
Q_MX02 U2633 ( .S(n1965), .A0(n2511), .A1(bCount[10]), .Z(n2104));
Q_FDP0UA U2634 ( .D(n2104), .QTFCLK( ), .Q(bCount[10]));
Q_MX02 U2635 ( .S(n1965), .A0(n2509), .A1(bCount[11]), .Z(n2105));
Q_FDP0UA U2636 ( .D(n2105), .QTFCLK( ), .Q(bCount[11]));
Q_MX02 U2637 ( .S(n1965), .A0(n2507), .A1(bCount[12]), .Z(n2106));
Q_FDP0UA U2638 ( .D(n2106), .QTFCLK( ), .Q(bCount[12]));
Q_MX02 U2639 ( .S(n1965), .A0(n2505), .A1(bCount[13]), .Z(n2107));
Q_FDP0UA U2640 ( .D(n2107), .QTFCLK( ), .Q(bCount[13]));
Q_MX02 U2641 ( .S(n1965), .A0(n2503), .A1(bCount[14]), .Z(n2108));
Q_FDP0UA U2642 ( .D(n2108), .QTFCLK( ), .Q(bCount[14]));
Q_MX02 U2643 ( .S(n1965), .A0(n2501), .A1(bCount[15]), .Z(n2109));
Q_FDP0UA U2644 ( .D(n2109), .QTFCLK( ), .Q(bCount[15]));
Q_MX02 U2645 ( .S(n1965), .A0(n2499), .A1(bCount[16]), .Z(n2110));
Q_FDP0UA U2646 ( .D(n2110), .QTFCLK( ), .Q(bCount[16]));
Q_MX02 U2647 ( .S(n1965), .A0(n2497), .A1(bCount[17]), .Z(n2111));
Q_FDP0UA U2648 ( .D(n2111), .QTFCLK( ), .Q(bCount[17]));
Q_MX02 U2649 ( .S(n1965), .A0(n2495), .A1(bCount[18]), .Z(n2112));
Q_FDP0UA U2650 ( .D(n2112), .QTFCLK( ), .Q(bCount[18]));
Q_MX02 U2651 ( .S(n1965), .A0(n2493), .A1(bCount[19]), .Z(n2113));
Q_FDP0UA U2652 ( .D(n2113), .QTFCLK( ), .Q(bCount[19]));
Q_MX02 U2653 ( .S(n1965), .A0(n2491), .A1(bCount[20]), .Z(n2114));
Q_FDP0UA U2654 ( .D(n2114), .QTFCLK( ), .Q(bCount[20]));
Q_MX02 U2655 ( .S(n1965), .A0(n2489), .A1(bCount[21]), .Z(n2115));
Q_FDP0UA U2656 ( .D(n2115), .QTFCLK( ), .Q(bCount[21]));
Q_MX02 U2657 ( .S(n1965), .A0(n2487), .A1(bCount[22]), .Z(n2116));
Q_FDP0UA U2658 ( .D(n2116), .QTFCLK( ), .Q(bCount[22]));
Q_MX02 U2659 ( .S(n1965), .A0(n2485), .A1(bCount[23]), .Z(n2117));
Q_FDP0UA U2660 ( .D(n2117), .QTFCLK( ), .Q(bCount[23]));
Q_MX02 U2661 ( .S(n1965), .A0(n2483), .A1(bCount[24]), .Z(n2118));
Q_FDP0UA U2662 ( .D(n2118), .QTFCLK( ), .Q(bCount[24]));
Q_MX02 U2663 ( .S(n1965), .A0(n2481), .A1(bCount[25]), .Z(n2119));
Q_FDP0UA U2664 ( .D(n2119), .QTFCLK( ), .Q(bCount[25]));
Q_MX02 U2665 ( .S(n1965), .A0(n2479), .A1(bCount[26]), .Z(n2120));
Q_FDP0UA U2666 ( .D(n2120), .QTFCLK( ), .Q(bCount[26]));
Q_MX02 U2667 ( .S(n1965), .A0(n2477), .A1(bCount[27]), .Z(n2121));
Q_FDP0UA U2668 ( .D(n2121), .QTFCLK( ), .Q(bCount[27]));
Q_MX02 U2669 ( .S(n1965), .A0(n2475), .A1(bCount[28]), .Z(n2122));
Q_FDP0UA U2670 ( .D(n2122), .QTFCLK( ), .Q(bCount[28]));
Q_MX02 U2671 ( .S(n1965), .A0(n2473), .A1(bCount[29]), .Z(n2123));
Q_FDP0UA U2672 ( .D(n2123), .QTFCLK( ), .Q(bCount[29]));
Q_MX02 U2673 ( .S(n1965), .A0(n2471), .A1(bCount[30]), .Z(n2124));
Q_FDP0UA U2674 ( .D(n2124), .QTFCLK( ), .Q(bCount[30]));
Q_MX02 U2675 ( .S(n1965), .A0(n2469), .A1(bCount[31]), .Z(n2125));
Q_FDP0UA U2676 ( .D(n2125), .QTFCLK( ), .Q(bCount[31]));
Q_MX02 U2677 ( .S(n1965), .A0(n2467), .A1(bCount[32]), .Z(n2126));
Q_FDP0UA U2678 ( .D(n2126), .QTFCLK( ), .Q(bCount[32]));
Q_MX02 U2679 ( .S(n1965), .A0(n2465), .A1(bCount[33]), .Z(n2127));
Q_FDP0UA U2680 ( .D(n2127), .QTFCLK( ), .Q(bCount[33]));
Q_MX02 U2681 ( .S(n1965), .A0(n2463), .A1(bCount[34]), .Z(n2128));
Q_FDP0UA U2682 ( .D(n2128), .QTFCLK( ), .Q(bCount[34]));
Q_MX02 U2683 ( .S(n1965), .A0(n2461), .A1(bCount[35]), .Z(n2129));
Q_FDP0UA U2684 ( .D(n2129), .QTFCLK( ), .Q(bCount[35]));
Q_MX02 U2685 ( .S(n1965), .A0(n2459), .A1(bCount[36]), .Z(n2130));
Q_FDP0UA U2686 ( .D(n2130), .QTFCLK( ), .Q(bCount[36]));
Q_MX02 U2687 ( .S(n1965), .A0(n2457), .A1(bCount[37]), .Z(n2131));
Q_FDP0UA U2688 ( .D(n2131), .QTFCLK( ), .Q(bCount[37]));
Q_MX02 U2689 ( .S(n1965), .A0(n2455), .A1(bCount[38]), .Z(n2132));
Q_FDP0UA U2690 ( .D(n2132), .QTFCLK( ), .Q(bCount[38]));
Q_MX02 U2691 ( .S(n1965), .A0(n2453), .A1(bCount[39]), .Z(n2133));
Q_FDP0UA U2692 ( .D(n2133), .QTFCLK( ), .Q(bCount[39]));
Q_MX02 U2693 ( .S(n1965), .A0(n2451), .A1(bCount[40]), .Z(n2134));
Q_FDP0UA U2694 ( .D(n2134), .QTFCLK( ), .Q(bCount[40]));
Q_MX02 U2695 ( .S(n1965), .A0(n2449), .A1(bCount[41]), .Z(n2135));
Q_FDP0UA U2696 ( .D(n2135), .QTFCLK( ), .Q(bCount[41]));
Q_MX02 U2697 ( .S(n1965), .A0(n2447), .A1(bCount[42]), .Z(n2136));
Q_FDP0UA U2698 ( .D(n2136), .QTFCLK( ), .Q(bCount[42]));
Q_MX02 U2699 ( .S(n1965), .A0(n2445), .A1(bCount[43]), .Z(n2137));
Q_FDP0UA U2700 ( .D(n2137), .QTFCLK( ), .Q(bCount[43]));
Q_MX02 U2701 ( .S(n1965), .A0(n2443), .A1(bCount[44]), .Z(n2138));
Q_FDP0UA U2702 ( .D(n2138), .QTFCLK( ), .Q(bCount[44]));
Q_MX02 U2703 ( .S(n1965), .A0(n2441), .A1(bCount[45]), .Z(n2139));
Q_FDP0UA U2704 ( .D(n2139), .QTFCLK( ), .Q(bCount[45]));
Q_MX02 U2705 ( .S(n1965), .A0(n2439), .A1(bCount[46]), .Z(n2140));
Q_FDP0UA U2706 ( .D(n2140), .QTFCLK( ), .Q(bCount[46]));
Q_MX02 U2707 ( .S(n1965), .A0(n2437), .A1(bCount[47]), .Z(n2141));
Q_FDP0UA U2708 ( .D(n2141), .QTFCLK( ), .Q(bCount[47]));
Q_MX02 U2709 ( .S(n1965), .A0(n2435), .A1(bCount[48]), .Z(n2142));
Q_FDP0UA U2710 ( .D(n2142), .QTFCLK( ), .Q(bCount[48]));
Q_MX02 U2711 ( .S(n1965), .A0(n2433), .A1(bCount[49]), .Z(n2143));
Q_FDP0UA U2712 ( .D(n2143), .QTFCLK( ), .Q(bCount[49]));
Q_MX02 U2713 ( .S(n1965), .A0(n2431), .A1(bCount[50]), .Z(n2144));
Q_FDP0UA U2714 ( .D(n2144), .QTFCLK( ), .Q(bCount[50]));
Q_MX02 U2715 ( .S(n1965), .A0(n2429), .A1(bCount[51]), .Z(n2145));
Q_FDP0UA U2716 ( .D(n2145), .QTFCLK( ), .Q(bCount[51]));
Q_MX02 U2717 ( .S(n1965), .A0(n2427), .A1(bCount[52]), .Z(n2146));
Q_FDP0UA U2718 ( .D(n2146), .QTFCLK( ), .Q(bCount[52]));
Q_MX02 U2719 ( .S(n1965), .A0(n2425), .A1(bCount[53]), .Z(n2147));
Q_FDP0UA U2720 ( .D(n2147), .QTFCLK( ), .Q(bCount[53]));
Q_MX02 U2721 ( .S(n1965), .A0(n2423), .A1(bCount[54]), .Z(n2148));
Q_FDP0UA U2722 ( .D(n2148), .QTFCLK( ), .Q(bCount[54]));
Q_MX02 U2723 ( .S(n1965), .A0(n2421), .A1(bCount[55]), .Z(n2149));
Q_FDP0UA U2724 ( .D(n2149), .QTFCLK( ), .Q(bCount[55]));
Q_MX02 U2725 ( .S(n1965), .A0(n2419), .A1(bCount[56]), .Z(n2150));
Q_FDP0UA U2726 ( .D(n2150), .QTFCLK( ), .Q(bCount[56]));
Q_MX02 U2727 ( .S(n1965), .A0(n2417), .A1(bCount[57]), .Z(n2151));
Q_FDP0UA U2728 ( .D(n2151), .QTFCLK( ), .Q(bCount[57]));
Q_MX02 U2729 ( .S(n1965), .A0(n2415), .A1(bCount[58]), .Z(n2152));
Q_FDP0UA U2730 ( .D(n2152), .QTFCLK( ), .Q(bCount[58]));
Q_MX02 U2731 ( .S(n1965), .A0(n2413), .A1(bCount[59]), .Z(n2153));
Q_FDP0UA U2732 ( .D(n2153), .QTFCLK( ), .Q(bCount[59]));
Q_MX02 U2733 ( .S(n1965), .A0(n2411), .A1(bCount[60]), .Z(n2154));
Q_FDP0UA U2734 ( .D(n2154), .QTFCLK( ), .Q(bCount[60]));
Q_MX02 U2735 ( .S(n1965), .A0(n2409), .A1(bCount[61]), .Z(n2155));
Q_FDP0UA U2736 ( .D(n2155), .QTFCLK( ), .Q(bCount[61]));
Q_MX02 U2737 ( .S(n1965), .A0(n2407), .A1(bCount[62]), .Z(n2156));
Q_FDP0UA U2738 ( .D(n2156), .QTFCLK( ), .Q(bCount[62]));
Q_FDP0UA U2739 ( .D(n2157), .QTFCLK( ), .Q(bCount[63]));
Q_XOR2 U2740 ( .A0(ixcHoldClkCnt[63]), .A1(n7), .Z(n2029));
Q_AD01HF U2741 ( .A0(ixcHoldClkCnt[62]), .B0(n2160), .S(n2159), .CO(n2158));
Q_AD01HF U2742 ( .A0(ixcHoldClkCnt[61]), .B0(n2162), .S(n2161), .CO(n2160));
Q_AD01HF U2743 ( .A0(ixcHoldClkCnt[60]), .B0(n2164), .S(n2163), .CO(n2162));
Q_AD01HF U2744 ( .A0(ixcHoldClkCnt[59]), .B0(n2166), .S(n2165), .CO(n2164));
Q_AD01HF U2745 ( .A0(ixcHoldClkCnt[58]), .B0(n2168), .S(n2167), .CO(n2166));
Q_AD01HF U2746 ( .A0(ixcHoldClkCnt[57]), .B0(n2170), .S(n2169), .CO(n2168));
Q_AD01HF U2747 ( .A0(ixcHoldClkCnt[56]), .B0(n2172), .S(n2171), .CO(n2170));
Q_AD01HF U2748 ( .A0(ixcHoldClkCnt[55]), .B0(n2174), .S(n2173), .CO(n2172));
Q_AD01HF U2749 ( .A0(ixcHoldClkCnt[54]), .B0(n2176), .S(n2175), .CO(n2174));
Q_AD01HF U2750 ( .A0(ixcHoldClkCnt[53]), .B0(n2178), .S(n2177), .CO(n2176));
Q_AD01HF U2751 ( .A0(ixcHoldClkCnt[52]), .B0(n2180), .S(n2179), .CO(n2178));
Q_AD01HF U2752 ( .A0(ixcHoldClkCnt[51]), .B0(n2182), .S(n2181), .CO(n2180));
Q_AD01HF U2753 ( .A0(ixcHoldClkCnt[50]), .B0(n2184), .S(n2183), .CO(n2182));
Q_AD01HF U2754 ( .A0(ixcHoldClkCnt[49]), .B0(n2186), .S(n2185), .CO(n2184));
Q_AD01HF U2755 ( .A0(ixcHoldClkCnt[48]), .B0(n2188), .S(n2187), .CO(n2186));
Q_AD01HF U2756 ( .A0(ixcHoldClkCnt[47]), .B0(n2190), .S(n2189), .CO(n2188));
Q_AD01HF U2757 ( .A0(ixcHoldClkCnt[46]), .B0(n2192), .S(n2191), .CO(n2190));
Q_AD01HF U2758 ( .A0(ixcHoldClkCnt[45]), .B0(n2194), .S(n2193), .CO(n2192));
Q_AD01HF U2759 ( .A0(ixcHoldClkCnt[44]), .B0(n2196), .S(n2195), .CO(n2194));
Q_AD01HF U2760 ( .A0(ixcHoldClkCnt[43]), .B0(n2198), .S(n2197), .CO(n2196));
Q_AD01HF U2761 ( .A0(ixcHoldClkCnt[42]), .B0(n2200), .S(n2199), .CO(n2198));
Q_AD01HF U2762 ( .A0(ixcHoldClkCnt[41]), .B0(n2202), .S(n2201), .CO(n2200));
Q_AD01HF U2763 ( .A0(ixcHoldClkCnt[40]), .B0(n2204), .S(n2203), .CO(n2202));
Q_AD01HF U2764 ( .A0(ixcHoldClkCnt[39]), .B0(n2206), .S(n2205), .CO(n2204));
Q_AD01HF U2765 ( .A0(ixcHoldClkCnt[38]), .B0(n2208), .S(n2207), .CO(n2206));
Q_AD01HF U2766 ( .A0(ixcHoldClkCnt[37]), .B0(n2210), .S(n2209), .CO(n2208));
Q_AD01HF U2767 ( .A0(ixcHoldClkCnt[36]), .B0(n2212), .S(n2211), .CO(n2210));
Q_AD01HF U2768 ( .A0(ixcHoldClkCnt[35]), .B0(n2214), .S(n2213), .CO(n2212));
Q_AD01HF U2769 ( .A0(ixcHoldClkCnt[34]), .B0(n2216), .S(n2215), .CO(n2214));
Q_AD01HF U2770 ( .A0(ixcHoldClkCnt[33]), .B0(n2218), .S(n2217), .CO(n2216));
Q_AD01HF U2771 ( .A0(ixcHoldClkCnt[32]), .B0(n2220), .S(n2219), .CO(n2218));
Q_AD01HF U2772 ( .A0(ixcHoldClkCnt[31]), .B0(n2222), .S(n2221), .CO(n2220));
Q_AD01HF U2773 ( .A0(ixcHoldClkCnt[30]), .B0(n2224), .S(n2223), .CO(n2222));
Q_AD01HF U2774 ( .A0(ixcHoldClkCnt[29]), .B0(n2226), .S(n2225), .CO(n2224));
Q_AD01HF U2775 ( .A0(ixcHoldClkCnt[28]), .B0(n2228), .S(n2227), .CO(n2226));
Q_AD01HF U2776 ( .A0(ixcHoldClkCnt[27]), .B0(n2230), .S(n2229), .CO(n2228));
Q_AD01HF U2777 ( .A0(ixcHoldClkCnt[26]), .B0(n2232), .S(n2231), .CO(n2230));
Q_AD01HF U2778 ( .A0(ixcHoldClkCnt[25]), .B0(n2234), .S(n2233), .CO(n2232));
Q_AD01HF U2779 ( .A0(ixcHoldClkCnt[24]), .B0(n2236), .S(n2235), .CO(n2234));
Q_AD01HF U2780 ( .A0(ixcHoldClkCnt[23]), .B0(n2238), .S(n2237), .CO(n2236));
Q_AD01HF U2781 ( .A0(ixcHoldClkCnt[22]), .B0(n2240), .S(n2239), .CO(n2238));
Q_AD01HF U2782 ( .A0(ixcHoldClkCnt[21]), .B0(n2242), .S(n2241), .CO(n2240));
Q_AD01HF U2783 ( .A0(ixcHoldClkCnt[20]), .B0(n2244), .S(n2243), .CO(n2242));
Q_AD01HF U2784 ( .A0(ixcHoldClkCnt[19]), .B0(n2246), .S(n2245), .CO(n2244));
Q_AD01HF U2785 ( .A0(ixcHoldClkCnt[18]), .B0(n2248), .S(n2247), .CO(n2246));
Q_AD01HF U2786 ( .A0(ixcHoldClkCnt[17]), .B0(n2250), .S(n2249), .CO(n2248));
Q_AD01HF U2787 ( .A0(ixcHoldClkCnt[16]), .B0(n2252), .S(n2251), .CO(n2250));
Q_AD01HF U2788 ( .A0(ixcHoldClkCnt[15]), .B0(n2254), .S(n2253), .CO(n2252));
Q_AD01HF U2789 ( .A0(ixcHoldClkCnt[14]), .B0(n2256), .S(n2255), .CO(n2254));
Q_AD01HF U2790 ( .A0(ixcHoldClkCnt[13]), .B0(n2258), .S(n2257), .CO(n2256));
Q_AD01HF U2791 ( .A0(ixcHoldClkCnt[12]), .B0(n2260), .S(n2259), .CO(n2258));
Q_AD01HF U2792 ( .A0(ixcHoldClkCnt[11]), .B0(n2262), .S(n2261), .CO(n2260));
Q_AD01HF U2793 ( .A0(ixcHoldClkCnt[10]), .B0(n2264), .S(n2263), .CO(n2262));
Q_AD01HF U2794 ( .A0(ixcHoldClkCnt[9]), .B0(n2266), .S(n2265), .CO(n2264));
Q_AD01HF U2795 ( .A0(ixcHoldClkCnt[8]), .B0(n2268), .S(n2267), .CO(n2266));
Q_AD01HF U2796 ( .A0(ixcHoldClkCnt[7]), .B0(n2270), .S(n2269), .CO(n2268));
Q_AD01HF U2797 ( .A0(ixcHoldClkCnt[6]), .B0(n2272), .S(n2271), .CO(n2270));
Q_AD01HF U2798 ( .A0(ixcHoldClkCnt[5]), .B0(n2274), .S(n2273), .CO(n2272));
Q_AD01HF U2799 ( .A0(ixcHoldClkCnt[4]), .B0(n2276), .S(n2275), .CO(n2274));
Q_AD01HF U2800 ( .A0(ixcHoldClkCnt[3]), .B0(n2278), .S(n2277), .CO(n2276));
Q_AD01HF U2801 ( .A0(ixcHoldClkCnt[2]), .B0(n2280), .S(n2279), .CO(n2278));
Q_AD01HF U2802 ( .A0(ixcHoldClkCnt[1]), .B0(ixcHoldClkCnt[0]), .S(n2281), .CO(n2280));
Q_XOR2 U2803 ( .A0(nbaCount[63]), .A1(n6), .Z(n2093));
Q_AD01HF U2804 ( .A0(nbaCount[62]), .B0(n2284), .S(n2283), .CO(n2282));
Q_AD01HF U2805 ( .A0(nbaCount[61]), .B0(n2286), .S(n2285), .CO(n2284));
Q_AD01HF U2806 ( .A0(nbaCount[60]), .B0(n2288), .S(n2287), .CO(n2286));
Q_AD01HF U2807 ( .A0(nbaCount[59]), .B0(n2290), .S(n2289), .CO(n2288));
Q_AD01HF U2808 ( .A0(nbaCount[58]), .B0(n2292), .S(n2291), .CO(n2290));
Q_AD01HF U2809 ( .A0(nbaCount[57]), .B0(n2294), .S(n2293), .CO(n2292));
Q_AD01HF U2810 ( .A0(nbaCount[56]), .B0(n2296), .S(n2295), .CO(n2294));
Q_AD01HF U2811 ( .A0(nbaCount[55]), .B0(n2298), .S(n2297), .CO(n2296));
Q_AD01HF U2812 ( .A0(nbaCount[54]), .B0(n2300), .S(n2299), .CO(n2298));
Q_AD01HF U2813 ( .A0(nbaCount[53]), .B0(n2302), .S(n2301), .CO(n2300));
Q_AD01HF U2814 ( .A0(nbaCount[52]), .B0(n2304), .S(n2303), .CO(n2302));
Q_AD01HF U2815 ( .A0(nbaCount[51]), .B0(n2306), .S(n2305), .CO(n2304));
Q_AD01HF U2816 ( .A0(nbaCount[50]), .B0(n2308), .S(n2307), .CO(n2306));
Q_AD01HF U2817 ( .A0(nbaCount[49]), .B0(n2310), .S(n2309), .CO(n2308));
Q_AD01HF U2818 ( .A0(nbaCount[48]), .B0(n2312), .S(n2311), .CO(n2310));
Q_AD01HF U2819 ( .A0(nbaCount[47]), .B0(n2314), .S(n2313), .CO(n2312));
Q_AD01HF U2820 ( .A0(nbaCount[46]), .B0(n2316), .S(n2315), .CO(n2314));
Q_AD01HF U2821 ( .A0(nbaCount[45]), .B0(n2318), .S(n2317), .CO(n2316));
Q_AD01HF U2822 ( .A0(nbaCount[44]), .B0(n2320), .S(n2319), .CO(n2318));
Q_AD01HF U2823 ( .A0(nbaCount[43]), .B0(n2322), .S(n2321), .CO(n2320));
Q_AD01HF U2824 ( .A0(nbaCount[42]), .B0(n2324), .S(n2323), .CO(n2322));
Q_AD01HF U2825 ( .A0(nbaCount[41]), .B0(n2326), .S(n2325), .CO(n2324));
Q_AD01HF U2826 ( .A0(nbaCount[40]), .B0(n2328), .S(n2327), .CO(n2326));
Q_AD01HF U2827 ( .A0(nbaCount[39]), .B0(n2330), .S(n2329), .CO(n2328));
Q_AD01HF U2828 ( .A0(nbaCount[38]), .B0(n2332), .S(n2331), .CO(n2330));
Q_AD01HF U2829 ( .A0(nbaCount[37]), .B0(n2334), .S(n2333), .CO(n2332));
Q_AD01HF U2830 ( .A0(nbaCount[36]), .B0(n2336), .S(n2335), .CO(n2334));
Q_AD01HF U2831 ( .A0(nbaCount[35]), .B0(n2338), .S(n2337), .CO(n2336));
Q_AD01HF U2832 ( .A0(nbaCount[34]), .B0(n2340), .S(n2339), .CO(n2338));
Q_AD01HF U2833 ( .A0(nbaCount[33]), .B0(n2342), .S(n2341), .CO(n2340));
Q_AD01HF U2834 ( .A0(nbaCount[32]), .B0(n2344), .S(n2343), .CO(n2342));
Q_AD01HF U2835 ( .A0(nbaCount[31]), .B0(n2346), .S(n2345), .CO(n2344));
Q_AD01HF U2836 ( .A0(nbaCount[30]), .B0(n2348), .S(n2347), .CO(n2346));
Q_AD01HF U2837 ( .A0(nbaCount[29]), .B0(n2350), .S(n2349), .CO(n2348));
Q_AD01HF U2838 ( .A0(nbaCount[28]), .B0(n2352), .S(n2351), .CO(n2350));
Q_AD01HF U2839 ( .A0(nbaCount[27]), .B0(n2354), .S(n2353), .CO(n2352));
Q_AD01HF U2840 ( .A0(nbaCount[26]), .B0(n2356), .S(n2355), .CO(n2354));
Q_AD01HF U2841 ( .A0(nbaCount[25]), .B0(n2358), .S(n2357), .CO(n2356));
Q_AD01HF U2842 ( .A0(nbaCount[24]), .B0(n2360), .S(n2359), .CO(n2358));
Q_AD01HF U2843 ( .A0(nbaCount[23]), .B0(n2362), .S(n2361), .CO(n2360));
Q_AD01HF U2844 ( .A0(nbaCount[22]), .B0(n2364), .S(n2363), .CO(n2362));
Q_AD01HF U2845 ( .A0(nbaCount[21]), .B0(n2366), .S(n2365), .CO(n2364));
Q_AD01HF U2846 ( .A0(nbaCount[20]), .B0(n2368), .S(n2367), .CO(n2366));
Q_AD01HF U2847 ( .A0(nbaCount[19]), .B0(n2370), .S(n2369), .CO(n2368));
Q_AD01HF U2848 ( .A0(nbaCount[18]), .B0(n2372), .S(n2371), .CO(n2370));
Q_AD01HF U2849 ( .A0(nbaCount[17]), .B0(n2374), .S(n2373), .CO(n2372));
Q_AD01HF U2850 ( .A0(nbaCount[16]), .B0(n2376), .S(n2375), .CO(n2374));
Q_AD01HF U2851 ( .A0(nbaCount[15]), .B0(n2378), .S(n2377), .CO(n2376));
Q_AD01HF U2852 ( .A0(nbaCount[14]), .B0(n2380), .S(n2379), .CO(n2378));
Q_AD01HF U2853 ( .A0(nbaCount[13]), .B0(n2382), .S(n2381), .CO(n2380));
Q_AD01HF U2854 ( .A0(nbaCount[12]), .B0(n2384), .S(n2383), .CO(n2382));
Q_AD01HF U2855 ( .A0(nbaCount[11]), .B0(n2386), .S(n2385), .CO(n2384));
Q_AD01HF U2856 ( .A0(nbaCount[10]), .B0(n2388), .S(n2387), .CO(n2386));
Q_AD01HF U2857 ( .A0(nbaCount[9]), .B0(n2390), .S(n2389), .CO(n2388));
Q_AD01HF U2858 ( .A0(nbaCount[8]), .B0(n2392), .S(n2391), .CO(n2390));
Q_AD01HF U2859 ( .A0(nbaCount[7]), .B0(n2394), .S(n2393), .CO(n2392));
Q_AD01HF U2860 ( .A0(nbaCount[6]), .B0(n2396), .S(n2395), .CO(n2394));
Q_AD01HF U2861 ( .A0(nbaCount[5]), .B0(n2398), .S(n2397), .CO(n2396));
Q_AD01HF U2862 ( .A0(nbaCount[4]), .B0(n2400), .S(n2399), .CO(n2398));
Q_AD01HF U2863 ( .A0(nbaCount[3]), .B0(n2402), .S(n2401), .CO(n2400));
Q_AD01HF U2864 ( .A0(nbaCount[2]), .B0(n2404), .S(n2403), .CO(n2402));
Q_AD01HF U2865 ( .A0(nbaCount[1]), .B0(nbaCount[0]), .S(n2405), .CO(n2404));
Q_XOR2 U2866 ( .A0(bCount[63]), .A1(n5), .Z(n2157));
Q_AD01HF U2867 ( .A0(bCount[62]), .B0(n2408), .S(n2407), .CO(n2406));
Q_AD01HF U2868 ( .A0(bCount[61]), .B0(n2410), .S(n2409), .CO(n2408));
Q_AD01HF U2869 ( .A0(bCount[60]), .B0(n2412), .S(n2411), .CO(n2410));
Q_AD01HF U2870 ( .A0(bCount[59]), .B0(n2414), .S(n2413), .CO(n2412));
Q_AD01HF U2871 ( .A0(bCount[58]), .B0(n2416), .S(n2415), .CO(n2414));
Q_AD01HF U2872 ( .A0(bCount[57]), .B0(n2418), .S(n2417), .CO(n2416));
Q_AD01HF U2873 ( .A0(bCount[56]), .B0(n2420), .S(n2419), .CO(n2418));
Q_AD01HF U2874 ( .A0(bCount[55]), .B0(n2422), .S(n2421), .CO(n2420));
Q_AD01HF U2875 ( .A0(bCount[54]), .B0(n2424), .S(n2423), .CO(n2422));
Q_AD01HF U2876 ( .A0(bCount[53]), .B0(n2426), .S(n2425), .CO(n2424));
Q_AD01HF U2877 ( .A0(bCount[52]), .B0(n2428), .S(n2427), .CO(n2426));
Q_AD01HF U2878 ( .A0(bCount[51]), .B0(n2430), .S(n2429), .CO(n2428));
Q_AD01HF U2879 ( .A0(bCount[50]), .B0(n2432), .S(n2431), .CO(n2430));
Q_AD01HF U2880 ( .A0(bCount[49]), .B0(n2434), .S(n2433), .CO(n2432));
Q_AD01HF U2881 ( .A0(bCount[48]), .B0(n2436), .S(n2435), .CO(n2434));
Q_AD01HF U2882 ( .A0(bCount[47]), .B0(n2438), .S(n2437), .CO(n2436));
Q_AD01HF U2883 ( .A0(bCount[46]), .B0(n2440), .S(n2439), .CO(n2438));
Q_AD01HF U2884 ( .A0(bCount[45]), .B0(n2442), .S(n2441), .CO(n2440));
Q_AD01HF U2885 ( .A0(bCount[44]), .B0(n2444), .S(n2443), .CO(n2442));
Q_AD01HF U2886 ( .A0(bCount[43]), .B0(n2446), .S(n2445), .CO(n2444));
Q_AD01HF U2887 ( .A0(bCount[42]), .B0(n2448), .S(n2447), .CO(n2446));
Q_AD01HF U2888 ( .A0(bCount[41]), .B0(n2450), .S(n2449), .CO(n2448));
Q_AD01HF U2889 ( .A0(bCount[40]), .B0(n2452), .S(n2451), .CO(n2450));
Q_AD01HF U2890 ( .A0(bCount[39]), .B0(n2454), .S(n2453), .CO(n2452));
Q_AD01HF U2891 ( .A0(bCount[38]), .B0(n2456), .S(n2455), .CO(n2454));
Q_AD01HF U2892 ( .A0(bCount[37]), .B0(n2458), .S(n2457), .CO(n2456));
Q_AD01HF U2893 ( .A0(bCount[36]), .B0(n2460), .S(n2459), .CO(n2458));
Q_AD01HF U2894 ( .A0(bCount[35]), .B0(n2462), .S(n2461), .CO(n2460));
Q_AD01HF U2895 ( .A0(bCount[34]), .B0(n2464), .S(n2463), .CO(n2462));
Q_AD01HF U2896 ( .A0(bCount[33]), .B0(n2466), .S(n2465), .CO(n2464));
Q_AD01HF U2897 ( .A0(bCount[32]), .B0(n2468), .S(n2467), .CO(n2466));
Q_AD01HF U2898 ( .A0(bCount[31]), .B0(n2470), .S(n2469), .CO(n2468));
Q_AD01HF U2899 ( .A0(bCount[30]), .B0(n2472), .S(n2471), .CO(n2470));
Q_AD01HF U2900 ( .A0(bCount[29]), .B0(n2474), .S(n2473), .CO(n2472));
Q_AD01HF U2901 ( .A0(bCount[28]), .B0(n2476), .S(n2475), .CO(n2474));
Q_AD01HF U2902 ( .A0(bCount[27]), .B0(n2478), .S(n2477), .CO(n2476));
Q_AD01HF U2903 ( .A0(bCount[26]), .B0(n2480), .S(n2479), .CO(n2478));
Q_AD01HF U2904 ( .A0(bCount[25]), .B0(n2482), .S(n2481), .CO(n2480));
Q_AD01HF U2905 ( .A0(bCount[24]), .B0(n2484), .S(n2483), .CO(n2482));
Q_AD01HF U2906 ( .A0(bCount[23]), .B0(n2486), .S(n2485), .CO(n2484));
Q_AD01HF U2907 ( .A0(bCount[22]), .B0(n2488), .S(n2487), .CO(n2486));
Q_AD01HF U2908 ( .A0(bCount[21]), .B0(n2490), .S(n2489), .CO(n2488));
Q_AD01HF U2909 ( .A0(bCount[20]), .B0(n2492), .S(n2491), .CO(n2490));
Q_AD01HF U2910 ( .A0(bCount[19]), .B0(n2494), .S(n2493), .CO(n2492));
Q_AD01HF U2911 ( .A0(bCount[18]), .B0(n2496), .S(n2495), .CO(n2494));
Q_AD01HF U2912 ( .A0(bCount[17]), .B0(n2498), .S(n2497), .CO(n2496));
Q_AD01HF U2913 ( .A0(bCount[16]), .B0(n2500), .S(n2499), .CO(n2498));
Q_AD01HF U2914 ( .A0(bCount[15]), .B0(n2502), .S(n2501), .CO(n2500));
Q_AD01HF U2915 ( .A0(bCount[14]), .B0(n2504), .S(n2503), .CO(n2502));
Q_AD01HF U2916 ( .A0(bCount[13]), .B0(n2506), .S(n2505), .CO(n2504));
Q_AD01HF U2917 ( .A0(bCount[12]), .B0(n2508), .S(n2507), .CO(n2506));
Q_AD01HF U2918 ( .A0(bCount[11]), .B0(n2510), .S(n2509), .CO(n2508));
Q_AD01HF U2919 ( .A0(bCount[10]), .B0(n2512), .S(n2511), .CO(n2510));
Q_AD01HF U2920 ( .A0(bCount[9]), .B0(n2514), .S(n2513), .CO(n2512));
Q_AD01HF U2921 ( .A0(bCount[8]), .B0(n2516), .S(n2515), .CO(n2514));
Q_AD01HF U2922 ( .A0(bCount[7]), .B0(n2518), .S(n2517), .CO(n2516));
Q_AD01HF U2923 ( .A0(bCount[6]), .B0(n2520), .S(n2519), .CO(n2518));
Q_AD01HF U2924 ( .A0(bCount[5]), .B0(n2522), .S(n2521), .CO(n2520));
Q_AD01HF U2925 ( .A0(bCount[4]), .B0(n2524), .S(n2523), .CO(n2522));
Q_AD01HF U2926 ( .A0(bCount[3]), .B0(n2526), .S(n2525), .CO(n2524));
Q_AD01HF U2927 ( .A0(bCount[2]), .B0(n2528), .S(n2527), .CO(n2526));
Q_AD01HF U2928 ( .A0(bCount[1]), .B0(bCount[0]), .S(n2529), .CO(n2528));
Q_INV U2929 ( .A(n1409), .Z(n2530));
Q_XOR2 U2930 ( .A0(evalOn), .A1(fvSCount[0]), .Z(n2531));
Q_FDP0UA U2931 ( .D(n2531), .QTFCLK( ), .Q(fvSCount[0]));
Q_MX02 U2932 ( .S(evalOn), .A0(fvSCount[1]), .A1(n2782), .Z(n2532));
Q_FDP0UA U2933 ( .D(n2532), .QTFCLK( ), .Q(fvSCount[1]));
Q_MX02 U2934 ( .S(evalOn), .A0(fvSCount[2]), .A1(n2780), .Z(n2533));
Q_FDP0UA U2935 ( .D(n2533), .QTFCLK( ), .Q(fvSCount[2]));
Q_MX02 U2936 ( .S(evalOn), .A0(fvSCount[3]), .A1(n2778), .Z(n2534));
Q_FDP0UA U2937 ( .D(n2534), .QTFCLK( ), .Q(fvSCount[3]));
Q_MX02 U2938 ( .S(evalOn), .A0(fvSCount[4]), .A1(n2776), .Z(n2535));
Q_FDP0UA U2939 ( .D(n2535), .QTFCLK( ), .Q(fvSCount[4]));
Q_MX02 U2940 ( .S(evalOn), .A0(fvSCount[5]), .A1(n2774), .Z(n2536));
Q_FDP0UA U2941 ( .D(n2536), .QTFCLK( ), .Q(fvSCount[5]));
Q_MX02 U2942 ( .S(evalOn), .A0(fvSCount[6]), .A1(n2772), .Z(n2537));
Q_FDP0UA U2943 ( .D(n2537), .QTFCLK( ), .Q(fvSCount[6]));
Q_MX02 U2944 ( .S(evalOn), .A0(fvSCount[7]), .A1(n2770), .Z(n2538));
Q_FDP0UA U2945 ( .D(n2538), .QTFCLK( ), .Q(fvSCount[7]));
Q_MX02 U2946 ( .S(evalOn), .A0(fvSCount[8]), .A1(n2768), .Z(n2539));
Q_FDP0UA U2947 ( .D(n2539), .QTFCLK( ), .Q(fvSCount[8]));
Q_MX02 U2948 ( .S(evalOn), .A0(fvSCount[9]), .A1(n2766), .Z(n2540));
Q_FDP0UA U2949 ( .D(n2540), .QTFCLK( ), .Q(fvSCount[9]));
Q_MX02 U2950 ( .S(evalOn), .A0(fvSCount[10]), .A1(n2764), .Z(n2541));
Q_FDP0UA U2951 ( .D(n2541), .QTFCLK( ), .Q(fvSCount[10]));
Q_MX02 U2952 ( .S(evalOn), .A0(fvSCount[11]), .A1(n2762), .Z(n2542));
Q_FDP0UA U2953 ( .D(n2542), .QTFCLK( ), .Q(fvSCount[11]));
Q_MX02 U2954 ( .S(evalOn), .A0(fvSCount[12]), .A1(n2760), .Z(n2543));
Q_FDP0UA U2955 ( .D(n2543), .QTFCLK( ), .Q(fvSCount[12]));
Q_MX02 U2956 ( .S(evalOn), .A0(fvSCount[13]), .A1(n2758), .Z(n2544));
Q_FDP0UA U2957 ( .D(n2544), .QTFCLK( ), .Q(fvSCount[13]));
Q_MX02 U2958 ( .S(evalOn), .A0(fvSCount[14]), .A1(n2756), .Z(n2545));
Q_FDP0UA U2959 ( .D(n2545), .QTFCLK( ), .Q(fvSCount[14]));
Q_MX02 U2960 ( .S(evalOn), .A0(fvSCount[15]), .A1(n2754), .Z(n2546));
Q_FDP0UA U2961 ( .D(n2546), .QTFCLK( ), .Q(fvSCount[15]));
Q_MX02 U2962 ( .S(evalOn), .A0(fvSCount[16]), .A1(n2752), .Z(n2547));
Q_FDP0UA U2963 ( .D(n2547), .QTFCLK( ), .Q(fvSCount[16]));
Q_MX02 U2964 ( .S(evalOn), .A0(fvSCount[17]), .A1(n2750), .Z(n2548));
Q_FDP0UA U2965 ( .D(n2548), .QTFCLK( ), .Q(fvSCount[17]));
Q_MX02 U2966 ( .S(evalOn), .A0(fvSCount[18]), .A1(n2748), .Z(n2549));
Q_FDP0UA U2967 ( .D(n2549), .QTFCLK( ), .Q(fvSCount[18]));
Q_MX02 U2968 ( .S(evalOn), .A0(fvSCount[19]), .A1(n2746), .Z(n2550));
Q_FDP0UA U2969 ( .D(n2550), .QTFCLK( ), .Q(fvSCount[19]));
Q_MX02 U2970 ( .S(evalOn), .A0(fvSCount[20]), .A1(n2744), .Z(n2551));
Q_FDP0UA U2971 ( .D(n2551), .QTFCLK( ), .Q(fvSCount[20]));
Q_MX02 U2972 ( .S(evalOn), .A0(fvSCount[21]), .A1(n2742), .Z(n2552));
Q_FDP0UA U2973 ( .D(n2552), .QTFCLK( ), .Q(fvSCount[21]));
Q_MX02 U2974 ( .S(evalOn), .A0(fvSCount[22]), .A1(n2740), .Z(n2553));
Q_FDP0UA U2975 ( .D(n2553), .QTFCLK( ), .Q(fvSCount[22]));
Q_MX02 U2976 ( .S(evalOn), .A0(fvSCount[23]), .A1(n2738), .Z(n2554));
Q_FDP0UA U2977 ( .D(n2554), .QTFCLK( ), .Q(fvSCount[23]));
Q_MX02 U2978 ( .S(evalOn), .A0(fvSCount[24]), .A1(n2736), .Z(n2555));
Q_FDP0UA U2979 ( .D(n2555), .QTFCLK( ), .Q(fvSCount[24]));
Q_MX02 U2980 ( .S(evalOn), .A0(fvSCount[25]), .A1(n2734), .Z(n2556));
Q_FDP0UA U2981 ( .D(n2556), .QTFCLK( ), .Q(fvSCount[25]));
Q_MX02 U2982 ( .S(evalOn), .A0(fvSCount[26]), .A1(n2732), .Z(n2557));
Q_FDP0UA U2983 ( .D(n2557), .QTFCLK( ), .Q(fvSCount[26]));
Q_MX02 U2984 ( .S(evalOn), .A0(fvSCount[27]), .A1(n2730), .Z(n2558));
Q_FDP0UA U2985 ( .D(n2558), .QTFCLK( ), .Q(fvSCount[27]));
Q_MX02 U2986 ( .S(evalOn), .A0(fvSCount[28]), .A1(n2728), .Z(n2559));
Q_FDP0UA U2987 ( .D(n2559), .QTFCLK( ), .Q(fvSCount[28]));
Q_MX02 U2988 ( .S(evalOn), .A0(fvSCount[29]), .A1(n2726), .Z(n2560));
Q_FDP0UA U2989 ( .D(n2560), .QTFCLK( ), .Q(fvSCount[29]));
Q_MX02 U2990 ( .S(evalOn), .A0(fvSCount[30]), .A1(n2724), .Z(n2561));
Q_FDP0UA U2991 ( .D(n2561), .QTFCLK( ), .Q(fvSCount[30]));
Q_MX02 U2992 ( .S(evalOn), .A0(fvSCount[31]), .A1(n2722), .Z(n2562));
Q_FDP0UA U2993 ( .D(n2562), .QTFCLK( ), .Q(fvSCount[31]));
Q_MX02 U2994 ( .S(evalOn), .A0(fvSCount[32]), .A1(n2720), .Z(n2563));
Q_FDP0UA U2995 ( .D(n2563), .QTFCLK( ), .Q(fvSCount[32]));
Q_MX02 U2996 ( .S(evalOn), .A0(fvSCount[33]), .A1(n2718), .Z(n2564));
Q_FDP0UA U2997 ( .D(n2564), .QTFCLK( ), .Q(fvSCount[33]));
Q_MX02 U2998 ( .S(evalOn), .A0(fvSCount[34]), .A1(n2716), .Z(n2565));
Q_FDP0UA U2999 ( .D(n2565), .QTFCLK( ), .Q(fvSCount[34]));
Q_MX02 U3000 ( .S(evalOn), .A0(fvSCount[35]), .A1(n2714), .Z(n2566));
Q_FDP0UA U3001 ( .D(n2566), .QTFCLK( ), .Q(fvSCount[35]));
Q_MX02 U3002 ( .S(evalOn), .A0(fvSCount[36]), .A1(n2712), .Z(n2567));
Q_FDP0UA U3003 ( .D(n2567), .QTFCLK( ), .Q(fvSCount[36]));
Q_MX02 U3004 ( .S(evalOn), .A0(fvSCount[37]), .A1(n2710), .Z(n2568));
Q_FDP0UA U3005 ( .D(n2568), .QTFCLK( ), .Q(fvSCount[37]));
Q_MX02 U3006 ( .S(evalOn), .A0(fvSCount[38]), .A1(n2708), .Z(n2569));
Q_FDP0UA U3007 ( .D(n2569), .QTFCLK( ), .Q(fvSCount[38]));
Q_MX02 U3008 ( .S(evalOn), .A0(fvSCount[39]), .A1(n2706), .Z(n2570));
Q_FDP0UA U3009 ( .D(n2570), .QTFCLK( ), .Q(fvSCount[39]));
Q_MX02 U3010 ( .S(evalOn), .A0(fvSCount[40]), .A1(n2704), .Z(n2571));
Q_FDP0UA U3011 ( .D(n2571), .QTFCLK( ), .Q(fvSCount[40]));
Q_MX02 U3012 ( .S(evalOn), .A0(fvSCount[41]), .A1(n2702), .Z(n2572));
Q_FDP0UA U3013 ( .D(n2572), .QTFCLK( ), .Q(fvSCount[41]));
Q_MX02 U3014 ( .S(evalOn), .A0(fvSCount[42]), .A1(n2700), .Z(n2573));
Q_FDP0UA U3015 ( .D(n2573), .QTFCLK( ), .Q(fvSCount[42]));
Q_MX02 U3016 ( .S(evalOn), .A0(fvSCount[43]), .A1(n2698), .Z(n2574));
Q_FDP0UA U3017 ( .D(n2574), .QTFCLK( ), .Q(fvSCount[43]));
Q_MX02 U3018 ( .S(evalOn), .A0(fvSCount[44]), .A1(n2696), .Z(n2575));
Q_FDP0UA U3019 ( .D(n2575), .QTFCLK( ), .Q(fvSCount[44]));
Q_MX02 U3020 ( .S(evalOn), .A0(fvSCount[45]), .A1(n2694), .Z(n2576));
Q_FDP0UA U3021 ( .D(n2576), .QTFCLK( ), .Q(fvSCount[45]));
Q_MX02 U3022 ( .S(evalOn), .A0(fvSCount[46]), .A1(n2692), .Z(n2577));
Q_FDP0UA U3023 ( .D(n2577), .QTFCLK( ), .Q(fvSCount[46]));
Q_MX02 U3024 ( .S(evalOn), .A0(fvSCount[47]), .A1(n2690), .Z(n2578));
Q_FDP0UA U3025 ( .D(n2578), .QTFCLK( ), .Q(fvSCount[47]));
Q_MX02 U3026 ( .S(evalOn), .A0(fvSCount[48]), .A1(n2688), .Z(n2579));
Q_FDP0UA U3027 ( .D(n2579), .QTFCLK( ), .Q(fvSCount[48]));
Q_MX02 U3028 ( .S(evalOn), .A0(fvSCount[49]), .A1(n2686), .Z(n2580));
Q_FDP0UA U3029 ( .D(n2580), .QTFCLK( ), .Q(fvSCount[49]));
Q_MX02 U3030 ( .S(evalOn), .A0(fvSCount[50]), .A1(n2684), .Z(n2581));
Q_FDP0UA U3031 ( .D(n2581), .QTFCLK( ), .Q(fvSCount[50]));
Q_MX02 U3032 ( .S(evalOn), .A0(fvSCount[51]), .A1(n2682), .Z(n2582));
Q_FDP0UA U3033 ( .D(n2582), .QTFCLK( ), .Q(fvSCount[51]));
Q_MX02 U3034 ( .S(evalOn), .A0(fvSCount[52]), .A1(n2680), .Z(n2583));
Q_FDP0UA U3035 ( .D(n2583), .QTFCLK( ), .Q(fvSCount[52]));
Q_MX02 U3036 ( .S(evalOn), .A0(fvSCount[53]), .A1(n2678), .Z(n2584));
Q_FDP0UA U3037 ( .D(n2584), .QTFCLK( ), .Q(fvSCount[53]));
Q_MX02 U3038 ( .S(evalOn), .A0(fvSCount[54]), .A1(n2676), .Z(n2585));
Q_FDP0UA U3039 ( .D(n2585), .QTFCLK( ), .Q(fvSCount[54]));
Q_MX02 U3040 ( .S(evalOn), .A0(fvSCount[55]), .A1(n2674), .Z(n2586));
Q_FDP0UA U3041 ( .D(n2586), .QTFCLK( ), .Q(fvSCount[55]));
Q_MX02 U3042 ( .S(evalOn), .A0(fvSCount[56]), .A1(n2672), .Z(n2587));
Q_FDP0UA U3043 ( .D(n2587), .QTFCLK( ), .Q(fvSCount[56]));
Q_MX02 U3044 ( .S(evalOn), .A0(fvSCount[57]), .A1(n2670), .Z(n2588));
Q_FDP0UA U3045 ( .D(n2588), .QTFCLK( ), .Q(fvSCount[57]));
Q_MX02 U3046 ( .S(evalOn), .A0(fvSCount[58]), .A1(n2668), .Z(n2589));
Q_FDP0UA U3047 ( .D(n2589), .QTFCLK( ), .Q(fvSCount[58]));
Q_MX02 U3048 ( .S(evalOn), .A0(fvSCount[59]), .A1(n2666), .Z(n2590));
Q_FDP0UA U3049 ( .D(n2590), .QTFCLK( ), .Q(fvSCount[59]));
Q_MX02 U3050 ( .S(evalOn), .A0(fvSCount[60]), .A1(n2664), .Z(n2591));
Q_FDP0UA U3051 ( .D(n2591), .QTFCLK( ), .Q(fvSCount[60]));
Q_MX02 U3052 ( .S(evalOn), .A0(fvSCount[61]), .A1(n2662), .Z(n2592));
Q_FDP0UA U3053 ( .D(n2592), .QTFCLK( ), .Q(fvSCount[61]));
Q_MX02 U3054 ( .S(evalOn), .A0(fvSCount[62]), .A1(n2660), .Z(n2593));
Q_FDP0UA U3055 ( .D(n2593), .QTFCLK( ), .Q(fvSCount[62]));
Q_FDP0UA U3056 ( .D(n2594), .QTFCLK( ), .Q(fvSCount[63]));
Q_XOR2 U3057 ( .A0(n2530), .A1(evfCount[0]), .Z(n2595));
Q_FDP0UA U3058 ( .D(n2595), .QTFCLK( ), .Q(evfCount[0]));
Q_MX02 U3059 ( .S(n1409), .A0(n2906), .A1(evfCount[1]), .Z(n2596));
Q_FDP0UA U3060 ( .D(n2596), .QTFCLK( ), .Q(evfCount[1]));
Q_MX02 U3061 ( .S(n1409), .A0(n2904), .A1(evfCount[2]), .Z(n2597));
Q_FDP0UA U3062 ( .D(n2597), .QTFCLK( ), .Q(evfCount[2]));
Q_MX02 U3063 ( .S(n1409), .A0(n2902), .A1(evfCount[3]), .Z(n2598));
Q_FDP0UA U3064 ( .D(n2598), .QTFCLK( ), .Q(evfCount[3]));
Q_MX02 U3065 ( .S(n1409), .A0(n2900), .A1(evfCount[4]), .Z(n2599));
Q_FDP0UA U3066 ( .D(n2599), .QTFCLK( ), .Q(evfCount[4]));
Q_MX02 U3067 ( .S(n1409), .A0(n2898), .A1(evfCount[5]), .Z(n2600));
Q_FDP0UA U3068 ( .D(n2600), .QTFCLK( ), .Q(evfCount[5]));
Q_MX02 U3069 ( .S(n1409), .A0(n2896), .A1(evfCount[6]), .Z(n2601));
Q_FDP0UA U3070 ( .D(n2601), .QTFCLK( ), .Q(evfCount[6]));
Q_MX02 U3071 ( .S(n1409), .A0(n2894), .A1(evfCount[7]), .Z(n2602));
Q_FDP0UA U3072 ( .D(n2602), .QTFCLK( ), .Q(evfCount[7]));
Q_MX02 U3073 ( .S(n1409), .A0(n2892), .A1(evfCount[8]), .Z(n2603));
Q_FDP0UA U3074 ( .D(n2603), .QTFCLK( ), .Q(evfCount[8]));
Q_MX02 U3075 ( .S(n1409), .A0(n2890), .A1(evfCount[9]), .Z(n2604));
Q_FDP0UA U3076 ( .D(n2604), .QTFCLK( ), .Q(evfCount[9]));
Q_MX02 U3077 ( .S(n1409), .A0(n2888), .A1(evfCount[10]), .Z(n2605));
Q_FDP0UA U3078 ( .D(n2605), .QTFCLK( ), .Q(evfCount[10]));
Q_MX02 U3079 ( .S(n1409), .A0(n2886), .A1(evfCount[11]), .Z(n2606));
Q_FDP0UA U3080 ( .D(n2606), .QTFCLK( ), .Q(evfCount[11]));
Q_MX02 U3081 ( .S(n1409), .A0(n2884), .A1(evfCount[12]), .Z(n2607));
Q_FDP0UA U3082 ( .D(n2607), .QTFCLK( ), .Q(evfCount[12]));
Q_MX02 U3083 ( .S(n1409), .A0(n2882), .A1(evfCount[13]), .Z(n2608));
Q_FDP0UA U3084 ( .D(n2608), .QTFCLK( ), .Q(evfCount[13]));
Q_MX02 U3085 ( .S(n1409), .A0(n2880), .A1(evfCount[14]), .Z(n2609));
Q_FDP0UA U3086 ( .D(n2609), .QTFCLK( ), .Q(evfCount[14]));
Q_MX02 U3087 ( .S(n1409), .A0(n2878), .A1(evfCount[15]), .Z(n2610));
Q_FDP0UA U3088 ( .D(n2610), .QTFCLK( ), .Q(evfCount[15]));
Q_MX02 U3089 ( .S(n1409), .A0(n2876), .A1(evfCount[16]), .Z(n2611));
Q_FDP0UA U3090 ( .D(n2611), .QTFCLK( ), .Q(evfCount[16]));
Q_MX02 U3091 ( .S(n1409), .A0(n2874), .A1(evfCount[17]), .Z(n2612));
Q_FDP0UA U3092 ( .D(n2612), .QTFCLK( ), .Q(evfCount[17]));
Q_MX02 U3093 ( .S(n1409), .A0(n2872), .A1(evfCount[18]), .Z(n2613));
Q_FDP0UA U3094 ( .D(n2613), .QTFCLK( ), .Q(evfCount[18]));
Q_MX02 U3095 ( .S(n1409), .A0(n2870), .A1(evfCount[19]), .Z(n2614));
Q_FDP0UA U3096 ( .D(n2614), .QTFCLK( ), .Q(evfCount[19]));
Q_MX02 U3097 ( .S(n1409), .A0(n2868), .A1(evfCount[20]), .Z(n2615));
Q_FDP0UA U3098 ( .D(n2615), .QTFCLK( ), .Q(evfCount[20]));
Q_MX02 U3099 ( .S(n1409), .A0(n2866), .A1(evfCount[21]), .Z(n2616));
Q_FDP0UA U3100 ( .D(n2616), .QTFCLK( ), .Q(evfCount[21]));
Q_MX02 U3101 ( .S(n1409), .A0(n2864), .A1(evfCount[22]), .Z(n2617));
Q_FDP0UA U3102 ( .D(n2617), .QTFCLK( ), .Q(evfCount[22]));
Q_MX02 U3103 ( .S(n1409), .A0(n2862), .A1(evfCount[23]), .Z(n2618));
Q_FDP0UA U3104 ( .D(n2618), .QTFCLK( ), .Q(evfCount[23]));
Q_MX02 U3105 ( .S(n1409), .A0(n2860), .A1(evfCount[24]), .Z(n2619));
Q_FDP0UA U3106 ( .D(n2619), .QTFCLK( ), .Q(evfCount[24]));
Q_MX02 U3107 ( .S(n1409), .A0(n2858), .A1(evfCount[25]), .Z(n2620));
Q_FDP0UA U3108 ( .D(n2620), .QTFCLK( ), .Q(evfCount[25]));
Q_MX02 U3109 ( .S(n1409), .A0(n2856), .A1(evfCount[26]), .Z(n2621));
Q_FDP0UA U3110 ( .D(n2621), .QTFCLK( ), .Q(evfCount[26]));
Q_MX02 U3111 ( .S(n1409), .A0(n2854), .A1(evfCount[27]), .Z(n2622));
Q_FDP0UA U3112 ( .D(n2622), .QTFCLK( ), .Q(evfCount[27]));
Q_MX02 U3113 ( .S(n1409), .A0(n2852), .A1(evfCount[28]), .Z(n2623));
Q_FDP0UA U3114 ( .D(n2623), .QTFCLK( ), .Q(evfCount[28]));
Q_MX02 U3115 ( .S(n1409), .A0(n2850), .A1(evfCount[29]), .Z(n2624));
Q_FDP0UA U3116 ( .D(n2624), .QTFCLK( ), .Q(evfCount[29]));
Q_MX02 U3117 ( .S(n1409), .A0(n2848), .A1(evfCount[30]), .Z(n2625));
Q_FDP0UA U3118 ( .D(n2625), .QTFCLK( ), .Q(evfCount[30]));
Q_MX02 U3119 ( .S(n1409), .A0(n2846), .A1(evfCount[31]), .Z(n2626));
Q_FDP0UA U3120 ( .D(n2626), .QTFCLK( ), .Q(evfCount[31]));
Q_MX02 U3121 ( .S(n1409), .A0(n2844), .A1(evfCount[32]), .Z(n2627));
Q_FDP0UA U3122 ( .D(n2627), .QTFCLK( ), .Q(evfCount[32]));
Q_MX02 U3123 ( .S(n1409), .A0(n2842), .A1(evfCount[33]), .Z(n2628));
Q_FDP0UA U3124 ( .D(n2628), .QTFCLK( ), .Q(evfCount[33]));
Q_MX02 U3125 ( .S(n1409), .A0(n2840), .A1(evfCount[34]), .Z(n2629));
Q_FDP0UA U3126 ( .D(n2629), .QTFCLK( ), .Q(evfCount[34]));
Q_MX02 U3127 ( .S(n1409), .A0(n2838), .A1(evfCount[35]), .Z(n2630));
Q_FDP0UA U3128 ( .D(n2630), .QTFCLK( ), .Q(evfCount[35]));
Q_MX02 U3129 ( .S(n1409), .A0(n2836), .A1(evfCount[36]), .Z(n2631));
Q_FDP0UA U3130 ( .D(n2631), .QTFCLK( ), .Q(evfCount[36]));
Q_MX02 U3131 ( .S(n1409), .A0(n2834), .A1(evfCount[37]), .Z(n2632));
Q_FDP0UA U3132 ( .D(n2632), .QTFCLK( ), .Q(evfCount[37]));
Q_MX02 U3133 ( .S(n1409), .A0(n2832), .A1(evfCount[38]), .Z(n2633));
Q_FDP0UA U3134 ( .D(n2633), .QTFCLK( ), .Q(evfCount[38]));
Q_MX02 U3135 ( .S(n1409), .A0(n2830), .A1(evfCount[39]), .Z(n2634));
Q_FDP0UA U3136 ( .D(n2634), .QTFCLK( ), .Q(evfCount[39]));
Q_MX02 U3137 ( .S(n1409), .A0(n2828), .A1(evfCount[40]), .Z(n2635));
Q_FDP0UA U3138 ( .D(n2635), .QTFCLK( ), .Q(evfCount[40]));
Q_MX02 U3139 ( .S(n1409), .A0(n2826), .A1(evfCount[41]), .Z(n2636));
Q_FDP0UA U3140 ( .D(n2636), .QTFCLK( ), .Q(evfCount[41]));
Q_MX02 U3141 ( .S(n1409), .A0(n2824), .A1(evfCount[42]), .Z(n2637));
Q_FDP0UA U3142 ( .D(n2637), .QTFCLK( ), .Q(evfCount[42]));
Q_MX02 U3143 ( .S(n1409), .A0(n2822), .A1(evfCount[43]), .Z(n2638));
Q_FDP0UA U3144 ( .D(n2638), .QTFCLK( ), .Q(evfCount[43]));
Q_MX02 U3145 ( .S(n1409), .A0(n2820), .A1(evfCount[44]), .Z(n2639));
Q_FDP0UA U3146 ( .D(n2639), .QTFCLK( ), .Q(evfCount[44]));
Q_MX02 U3147 ( .S(n1409), .A0(n2818), .A1(evfCount[45]), .Z(n2640));
Q_FDP0UA U3148 ( .D(n2640), .QTFCLK( ), .Q(evfCount[45]));
Q_MX02 U3149 ( .S(n1409), .A0(n2816), .A1(evfCount[46]), .Z(n2641));
Q_FDP0UA U3150 ( .D(n2641), .QTFCLK( ), .Q(evfCount[46]));
Q_MX02 U3151 ( .S(n1409), .A0(n2814), .A1(evfCount[47]), .Z(n2642));
Q_FDP0UA U3152 ( .D(n2642), .QTFCLK( ), .Q(evfCount[47]));
Q_MX02 U3153 ( .S(n1409), .A0(n2812), .A1(evfCount[48]), .Z(n2643));
Q_FDP0UA U3154 ( .D(n2643), .QTFCLK( ), .Q(evfCount[48]));
Q_MX02 U3155 ( .S(n1409), .A0(n2810), .A1(evfCount[49]), .Z(n2644));
Q_FDP0UA U3156 ( .D(n2644), .QTFCLK( ), .Q(evfCount[49]));
Q_MX02 U3157 ( .S(n1409), .A0(n2808), .A1(evfCount[50]), .Z(n2645));
Q_FDP0UA U3158 ( .D(n2645), .QTFCLK( ), .Q(evfCount[50]));
Q_MX02 U3159 ( .S(n1409), .A0(n2806), .A1(evfCount[51]), .Z(n2646));
Q_FDP0UA U3160 ( .D(n2646), .QTFCLK( ), .Q(evfCount[51]));
Q_MX02 U3161 ( .S(n1409), .A0(n2804), .A1(evfCount[52]), .Z(n2647));
Q_FDP0UA U3162 ( .D(n2647), .QTFCLK( ), .Q(evfCount[52]));
Q_MX02 U3163 ( .S(n1409), .A0(n2802), .A1(evfCount[53]), .Z(n2648));
Q_FDP0UA U3164 ( .D(n2648), .QTFCLK( ), .Q(evfCount[53]));
Q_MX02 U3165 ( .S(n1409), .A0(n2800), .A1(evfCount[54]), .Z(n2649));
Q_FDP0UA U3166 ( .D(n2649), .QTFCLK( ), .Q(evfCount[54]));
Q_MX02 U3167 ( .S(n1409), .A0(n2798), .A1(evfCount[55]), .Z(n2650));
Q_FDP0UA U3168 ( .D(n2650), .QTFCLK( ), .Q(evfCount[55]));
Q_MX02 U3169 ( .S(n1409), .A0(n2796), .A1(evfCount[56]), .Z(n2651));
Q_FDP0UA U3170 ( .D(n2651), .QTFCLK( ), .Q(evfCount[56]));
Q_MX02 U3171 ( .S(n1409), .A0(n2794), .A1(evfCount[57]), .Z(n2652));
Q_FDP0UA U3172 ( .D(n2652), .QTFCLK( ), .Q(evfCount[57]));
Q_MX02 U3173 ( .S(n1409), .A0(n2792), .A1(evfCount[58]), .Z(n2653));
Q_FDP0UA U3174 ( .D(n2653), .QTFCLK( ), .Q(evfCount[58]));
Q_MX02 U3175 ( .S(n1409), .A0(n2790), .A1(evfCount[59]), .Z(n2654));
Q_FDP0UA U3176 ( .D(n2654), .QTFCLK( ), .Q(evfCount[59]));
Q_MX02 U3177 ( .S(n1409), .A0(n2788), .A1(evfCount[60]), .Z(n2655));
Q_FDP0UA U3178 ( .D(n2655), .QTFCLK( ), .Q(evfCount[60]));
Q_MX02 U3179 ( .S(n1409), .A0(n2786), .A1(evfCount[61]), .Z(n2656));
Q_FDP0UA U3180 ( .D(n2656), .QTFCLK( ), .Q(evfCount[61]));
Q_MX02 U3181 ( .S(n1409), .A0(n2784), .A1(evfCount[62]), .Z(n2657));
Q_FDP0UA U3182 ( .D(n2657), .QTFCLK( ), .Q(evfCount[62]));
Q_FDP0UA U3183 ( .D(n2658), .QTFCLK( ), .Q(evfCount[63]));
Q_XOR2 U3184 ( .A0(fvSCount[63]), .A1(n4), .Z(n2594));
Q_AD01HF U3185 ( .A0(fvSCount[62]), .B0(n2661), .S(n2660), .CO(n2659));
Q_AD01HF U3186 ( .A0(fvSCount[61]), .B0(n2663), .S(n2662), .CO(n2661));
Q_AD01HF U3187 ( .A0(fvSCount[60]), .B0(n2665), .S(n2664), .CO(n2663));
Q_AD01HF U3188 ( .A0(fvSCount[59]), .B0(n2667), .S(n2666), .CO(n2665));
Q_AD01HF U3189 ( .A0(fvSCount[58]), .B0(n2669), .S(n2668), .CO(n2667));
Q_AD01HF U3190 ( .A0(fvSCount[57]), .B0(n2671), .S(n2670), .CO(n2669));
Q_AD01HF U3191 ( .A0(fvSCount[56]), .B0(n2673), .S(n2672), .CO(n2671));
Q_AD01HF U3192 ( .A0(fvSCount[55]), .B0(n2675), .S(n2674), .CO(n2673));
Q_AD01HF U3193 ( .A0(fvSCount[54]), .B0(n2677), .S(n2676), .CO(n2675));
Q_AD01HF U3194 ( .A0(fvSCount[53]), .B0(n2679), .S(n2678), .CO(n2677));
Q_AD01HF U3195 ( .A0(fvSCount[52]), .B0(n2681), .S(n2680), .CO(n2679));
Q_AD01HF U3196 ( .A0(fvSCount[51]), .B0(n2683), .S(n2682), .CO(n2681));
Q_AD01HF U3197 ( .A0(fvSCount[50]), .B0(n2685), .S(n2684), .CO(n2683));
Q_AD01HF U3198 ( .A0(fvSCount[49]), .B0(n2687), .S(n2686), .CO(n2685));
Q_AD01HF U3199 ( .A0(fvSCount[48]), .B0(n2689), .S(n2688), .CO(n2687));
Q_AD01HF U3200 ( .A0(fvSCount[47]), .B0(n2691), .S(n2690), .CO(n2689));
Q_AD01HF U3201 ( .A0(fvSCount[46]), .B0(n2693), .S(n2692), .CO(n2691));
Q_AD01HF U3202 ( .A0(fvSCount[45]), .B0(n2695), .S(n2694), .CO(n2693));
Q_AD01HF U3203 ( .A0(fvSCount[44]), .B0(n2697), .S(n2696), .CO(n2695));
Q_AD01HF U3204 ( .A0(fvSCount[43]), .B0(n2699), .S(n2698), .CO(n2697));
Q_AD01HF U3205 ( .A0(fvSCount[42]), .B0(n2701), .S(n2700), .CO(n2699));
Q_AD01HF U3206 ( .A0(fvSCount[41]), .B0(n2703), .S(n2702), .CO(n2701));
Q_AD01HF U3207 ( .A0(fvSCount[40]), .B0(n2705), .S(n2704), .CO(n2703));
Q_AD01HF U3208 ( .A0(fvSCount[39]), .B0(n2707), .S(n2706), .CO(n2705));
Q_AD01HF U3209 ( .A0(fvSCount[38]), .B0(n2709), .S(n2708), .CO(n2707));
Q_AD01HF U3210 ( .A0(fvSCount[37]), .B0(n2711), .S(n2710), .CO(n2709));
Q_AD01HF U3211 ( .A0(fvSCount[36]), .B0(n2713), .S(n2712), .CO(n2711));
Q_AD01HF U3212 ( .A0(fvSCount[35]), .B0(n2715), .S(n2714), .CO(n2713));
Q_AD01HF U3213 ( .A0(fvSCount[34]), .B0(n2717), .S(n2716), .CO(n2715));
Q_AD01HF U3214 ( .A0(fvSCount[33]), .B0(n2719), .S(n2718), .CO(n2717));
Q_AD01HF U3215 ( .A0(fvSCount[32]), .B0(n2721), .S(n2720), .CO(n2719));
Q_AD01HF U3216 ( .A0(fvSCount[31]), .B0(n2723), .S(n2722), .CO(n2721));
Q_AD01HF U3217 ( .A0(fvSCount[30]), .B0(n2725), .S(n2724), .CO(n2723));
Q_AD01HF U3218 ( .A0(fvSCount[29]), .B0(n2727), .S(n2726), .CO(n2725));
Q_AD01HF U3219 ( .A0(fvSCount[28]), .B0(n2729), .S(n2728), .CO(n2727));
Q_AD01HF U3220 ( .A0(fvSCount[27]), .B0(n2731), .S(n2730), .CO(n2729));
Q_AD01HF U3221 ( .A0(fvSCount[26]), .B0(n2733), .S(n2732), .CO(n2731));
Q_AD01HF U3222 ( .A0(fvSCount[25]), .B0(n2735), .S(n2734), .CO(n2733));
Q_AD01HF U3223 ( .A0(fvSCount[24]), .B0(n2737), .S(n2736), .CO(n2735));
Q_AD01HF U3224 ( .A0(fvSCount[23]), .B0(n2739), .S(n2738), .CO(n2737));
Q_AD01HF U3225 ( .A0(fvSCount[22]), .B0(n2741), .S(n2740), .CO(n2739));
Q_AD01HF U3226 ( .A0(fvSCount[21]), .B0(n2743), .S(n2742), .CO(n2741));
Q_AD01HF U3227 ( .A0(fvSCount[20]), .B0(n2745), .S(n2744), .CO(n2743));
Q_AD01HF U3228 ( .A0(fvSCount[19]), .B0(n2747), .S(n2746), .CO(n2745));
Q_AD01HF U3229 ( .A0(fvSCount[18]), .B0(n2749), .S(n2748), .CO(n2747));
Q_AD01HF U3230 ( .A0(fvSCount[17]), .B0(n2751), .S(n2750), .CO(n2749));
Q_AD01HF U3231 ( .A0(fvSCount[16]), .B0(n2753), .S(n2752), .CO(n2751));
Q_AD01HF U3232 ( .A0(fvSCount[15]), .B0(n2755), .S(n2754), .CO(n2753));
Q_AD01HF U3233 ( .A0(fvSCount[14]), .B0(n2757), .S(n2756), .CO(n2755));
Q_AD01HF U3234 ( .A0(fvSCount[13]), .B0(n2759), .S(n2758), .CO(n2757));
Q_AD01HF U3235 ( .A0(fvSCount[12]), .B0(n2761), .S(n2760), .CO(n2759));
Q_AD01HF U3236 ( .A0(fvSCount[11]), .B0(n2763), .S(n2762), .CO(n2761));
Q_AD01HF U3237 ( .A0(fvSCount[10]), .B0(n2765), .S(n2764), .CO(n2763));
Q_AD01HF U3238 ( .A0(fvSCount[9]), .B0(n2767), .S(n2766), .CO(n2765));
Q_AD01HF U3239 ( .A0(fvSCount[8]), .B0(n2769), .S(n2768), .CO(n2767));
Q_AD01HF U3240 ( .A0(fvSCount[7]), .B0(n2771), .S(n2770), .CO(n2769));
Q_AD01HF U3241 ( .A0(fvSCount[6]), .B0(n2773), .S(n2772), .CO(n2771));
Q_AD01HF U3242 ( .A0(fvSCount[5]), .B0(n2775), .S(n2774), .CO(n2773));
Q_AD01HF U3243 ( .A0(fvSCount[4]), .B0(n2777), .S(n2776), .CO(n2775));
Q_AD01HF U3244 ( .A0(fvSCount[3]), .B0(n2779), .S(n2778), .CO(n2777));
Q_AD01HF U3245 ( .A0(fvSCount[2]), .B0(n2781), .S(n2780), .CO(n2779));
Q_AD01HF U3246 ( .A0(fvSCount[1]), .B0(fvSCount[0]), .S(n2782), .CO(n2781));
Q_XOR2 U3247 ( .A0(evfCount[63]), .A1(n3), .Z(n2658));
Q_AD01HF U3248 ( .A0(evfCount[62]), .B0(n2785), .S(n2784), .CO(n2783));
Q_AD01HF U3249 ( .A0(evfCount[61]), .B0(n2787), .S(n2786), .CO(n2785));
Q_AD01HF U3250 ( .A0(evfCount[60]), .B0(n2789), .S(n2788), .CO(n2787));
Q_AD01HF U3251 ( .A0(evfCount[59]), .B0(n2791), .S(n2790), .CO(n2789));
Q_AD01HF U3252 ( .A0(evfCount[58]), .B0(n2793), .S(n2792), .CO(n2791));
Q_AD01HF U3253 ( .A0(evfCount[57]), .B0(n2795), .S(n2794), .CO(n2793));
Q_AD01HF U3254 ( .A0(evfCount[56]), .B0(n2797), .S(n2796), .CO(n2795));
Q_AD01HF U3255 ( .A0(evfCount[55]), .B0(n2799), .S(n2798), .CO(n2797));
Q_AD01HF U3256 ( .A0(evfCount[54]), .B0(n2801), .S(n2800), .CO(n2799));
Q_AD01HF U3257 ( .A0(evfCount[53]), .B0(n2803), .S(n2802), .CO(n2801));
Q_AD01HF U3258 ( .A0(evfCount[52]), .B0(n2805), .S(n2804), .CO(n2803));
Q_AD01HF U3259 ( .A0(evfCount[51]), .B0(n2807), .S(n2806), .CO(n2805));
Q_AD01HF U3260 ( .A0(evfCount[50]), .B0(n2809), .S(n2808), .CO(n2807));
Q_AD01HF U3261 ( .A0(evfCount[49]), .B0(n2811), .S(n2810), .CO(n2809));
Q_AD01HF U3262 ( .A0(evfCount[48]), .B0(n2813), .S(n2812), .CO(n2811));
Q_AD01HF U3263 ( .A0(evfCount[47]), .B0(n2815), .S(n2814), .CO(n2813));
Q_AD01HF U3264 ( .A0(evfCount[46]), .B0(n2817), .S(n2816), .CO(n2815));
Q_AD01HF U3265 ( .A0(evfCount[45]), .B0(n2819), .S(n2818), .CO(n2817));
Q_AD01HF U3266 ( .A0(evfCount[44]), .B0(n2821), .S(n2820), .CO(n2819));
Q_AD01HF U3267 ( .A0(evfCount[43]), .B0(n2823), .S(n2822), .CO(n2821));
Q_AD01HF U3268 ( .A0(evfCount[42]), .B0(n2825), .S(n2824), .CO(n2823));
Q_AD01HF U3269 ( .A0(evfCount[41]), .B0(n2827), .S(n2826), .CO(n2825));
Q_AD01HF U3270 ( .A0(evfCount[40]), .B0(n2829), .S(n2828), .CO(n2827));
Q_AD01HF U3271 ( .A0(evfCount[39]), .B0(n2831), .S(n2830), .CO(n2829));
Q_AD01HF U3272 ( .A0(evfCount[38]), .B0(n2833), .S(n2832), .CO(n2831));
Q_AD01HF U3273 ( .A0(evfCount[37]), .B0(n2835), .S(n2834), .CO(n2833));
Q_AD01HF U3274 ( .A0(evfCount[36]), .B0(n2837), .S(n2836), .CO(n2835));
Q_AD01HF U3275 ( .A0(evfCount[35]), .B0(n2839), .S(n2838), .CO(n2837));
Q_AD01HF U3276 ( .A0(evfCount[34]), .B0(n2841), .S(n2840), .CO(n2839));
Q_AD01HF U3277 ( .A0(evfCount[33]), .B0(n2843), .S(n2842), .CO(n2841));
Q_AD01HF U3278 ( .A0(evfCount[32]), .B0(n2845), .S(n2844), .CO(n2843));
Q_AD01HF U3279 ( .A0(evfCount[31]), .B0(n2847), .S(n2846), .CO(n2845));
Q_AD01HF U3280 ( .A0(evfCount[30]), .B0(n2849), .S(n2848), .CO(n2847));
Q_AD01HF U3281 ( .A0(evfCount[29]), .B0(n2851), .S(n2850), .CO(n2849));
Q_AD01HF U3282 ( .A0(evfCount[28]), .B0(n2853), .S(n2852), .CO(n2851));
Q_AD01HF U3283 ( .A0(evfCount[27]), .B0(n2855), .S(n2854), .CO(n2853));
Q_AD01HF U3284 ( .A0(evfCount[26]), .B0(n2857), .S(n2856), .CO(n2855));
Q_AD01HF U3285 ( .A0(evfCount[25]), .B0(n2859), .S(n2858), .CO(n2857));
Q_AD01HF U3286 ( .A0(evfCount[24]), .B0(n2861), .S(n2860), .CO(n2859));
Q_AD01HF U3287 ( .A0(evfCount[23]), .B0(n2863), .S(n2862), .CO(n2861));
Q_AD01HF U3288 ( .A0(evfCount[22]), .B0(n2865), .S(n2864), .CO(n2863));
Q_AD01HF U3289 ( .A0(evfCount[21]), .B0(n2867), .S(n2866), .CO(n2865));
Q_AD01HF U3290 ( .A0(evfCount[20]), .B0(n2869), .S(n2868), .CO(n2867));
Q_AD01HF U3291 ( .A0(evfCount[19]), .B0(n2871), .S(n2870), .CO(n2869));
Q_AD01HF U3292 ( .A0(evfCount[18]), .B0(n2873), .S(n2872), .CO(n2871));
Q_AD01HF U3293 ( .A0(evfCount[17]), .B0(n2875), .S(n2874), .CO(n2873));
Q_AD01HF U3294 ( .A0(evfCount[16]), .B0(n2877), .S(n2876), .CO(n2875));
Q_AD01HF U3295 ( .A0(evfCount[15]), .B0(n2879), .S(n2878), .CO(n2877));
Q_AD01HF U3296 ( .A0(evfCount[14]), .B0(n2881), .S(n2880), .CO(n2879));
Q_AD01HF U3297 ( .A0(evfCount[13]), .B0(n2883), .S(n2882), .CO(n2881));
Q_AD01HF U3298 ( .A0(evfCount[12]), .B0(n2885), .S(n2884), .CO(n2883));
Q_AD01HF U3299 ( .A0(evfCount[11]), .B0(n2887), .S(n2886), .CO(n2885));
Q_AD01HF U3300 ( .A0(evfCount[10]), .B0(n2889), .S(n2888), .CO(n2887));
Q_AD01HF U3301 ( .A0(evfCount[9]), .B0(n2891), .S(n2890), .CO(n2889));
Q_AD01HF U3302 ( .A0(evfCount[8]), .B0(n2893), .S(n2892), .CO(n2891));
Q_AD01HF U3303 ( .A0(evfCount[7]), .B0(n2895), .S(n2894), .CO(n2893));
Q_AD01HF U3304 ( .A0(evfCount[6]), .B0(n2897), .S(n2896), .CO(n2895));
Q_AD01HF U3305 ( .A0(evfCount[5]), .B0(n2899), .S(n2898), .CO(n2897));
Q_AD01HF U3306 ( .A0(evfCount[4]), .B0(n2901), .S(n2900), .CO(n2899));
Q_AD01HF U3307 ( .A0(evfCount[3]), .B0(n2903), .S(n2902), .CO(n2901));
Q_AD01HF U3308 ( .A0(evfCount[2]), .B0(n2905), .S(n2904), .CO(n2903));
Q_AD01HF U3309 ( .A0(evfCount[1]), .B0(evfCount[0]), .S(n2906), .CO(n2905));
Q_INV U3310 ( .A(bpSt[0]), .Z(n2921));
Q_AN03 U3311 ( .A0(n2921), .A1(sampleXpChg), .A2(mpOn), .Z(n2910));
Q_INV U3312 ( .A(bpWait), .Z(n2922));
Q_AO21 U3313 ( .A0(bpSt[0]), .A1(n2922), .B0(n2910), .Z(n2912));
Q_OA21 U3314 ( .A0(bpSt[1]), .A1(mpOn), .B0(bpWait), .Z(n2911));
Q_AO21 U3315 ( .A0(bpSt[1]), .A1(n1962), .B0(n2911), .Z(n2913));
Q_INV U3316 ( .A(bpSt[1]), .Z(n2923));
Q_AN02 U3317 ( .A0(n2912), .A1(n2923), .Z(n2914));
Q_AO21 U3318 ( .A0(n2913), .A1(n2921), .B0(n2914), .Z(n2907));
Q_NR02 U3319 ( .A0(bpSt[1]), .A1(bpSt[0]), .Z(n2916));
Q_INV U3320 ( .A(mpOn), .Z(n2915));
Q_AO21 U3321 ( .A0(n2916), .A1(n2915), .B0(n2919), .Z(n2920));
Q_NR02 U3322 ( .A0(bpWait), .A1(sampleXpChg), .Z(n2917));
Q_AN02 U3323 ( .A0(bpSt[1]), .A1(bpSt[0]), .Z(n2918));
Q_OR03 U3324 ( .A0(GFBw), .A1(n2918), .A2(n2917), .Z(n2919));
Q_AN02 U3325 ( .A0(n2921), .A1(bpWait), .Z(n2908));
Q_NR02 U3326 ( .A0(bpSt[1]), .A1(n1963), .Z(n2909));
Q_MX02 U3327 ( .S(n2907), .A0(bpSt[0]), .A1(n2908), .Z(n2924));
Q_FDP0UA U3328 ( .D(n2924), .QTFCLK( ), .Q(bpSt[0]));
Q_MX02 U3329 ( .S(n2907), .A0(bpSt[1]), .A1(n2909), .Z(n2925));
Q_FDP0UA U3330 ( .D(n2925), .QTFCLK( ), .Q(bpSt[1]));
Q_XNR2 U3331 ( .A0(n2920), .A1(bClkR), .Z(n2926));
Q_FDP0UA U3332 ( .D(n2926), .QTFCLK( ), .Q(bClkR));
Q_FDP0UA U3333 ( .D(GFBw), .QTFCLK( ), .Q(bClkHoldD));
Q_FDP0UA U3334 ( .D(holdEcm), .QTFCLK( ), .Q(holdEcmD));
Q_FDP0UA U3335 ( .D(tbcPOStateN[1]), .QTFCLK( ), .Q(tbcPOState[1]));
Q_FDP0UA U3336 ( .D(tbcPOStateN[0]), .QTFCLK( ), .Q(tbcPOState[0]));
Q_INV U3337 ( .A(GF2LevelMask[0]), .Z(n2927));
Q_INV U3338 ( .A(GF2LevelMask[1]), .Z(n2928));
Q_INV U3339 ( .A(GF2LevelMask[2]), .Z(n2929));
Q_INV U3340 ( .A(GF2LevelMask[3]), .Z(n2930));
Q_INV U3341 ( .A(GF2LevelMask[4]), .Z(n2931));
Q_OR02 U3342 ( .A0(tbcPOd), .A1(n2927), .Z(n2932));
Q_OR02 U3343 ( .A0(tbcPODly[0]), .A1(n2928), .Z(n2933));
Q_OR02 U3344 ( .A0(tbcPODly[1]), .A1(n2929), .Z(n2934));
Q_OR02 U3345 ( .A0(tbcPODly[2]), .A1(n2930), .Z(n2935));
Q_OR02 U3346 ( .A0(tbcPODly[3]), .A1(n2931), .Z(n2936));
Q_FDP0UA U3347 ( .D(n2936), .QTFCLK( ), .Q(tbcPODly[4]));
Q_FDP0UA U3348 ( .D(n2935), .QTFCLK( ), .Q(tbcPODly[3]));
Q_FDP0UA U3349 ( .D(n2934), .QTFCLK( ), .Q(tbcPODly[2]));
Q_FDP0UA U3350 ( .D(n2933), .QTFCLK( ), .Q(tbcPODly[1]));
Q_FDP0UA U3351 ( .D(n2932), .QTFCLK( ), .Q(tbcPODly[0]));
Q_FDP0UA U3352 ( .D(GFbusyD), .QTFCLK( ), .Q(GFbusyD2));
Q_FDP0UA U3353 ( .D(GFbusy), .QTFCLK( ), .Q(GFbusyD));
Q_INV U3354 ( .A(active), .Z(n2937));
Q_NR02 U3355 ( .A0(active), .A1(asyncBusy), .Z(n2938));
Q_MX02 U3356 ( .S(n2938), .A0(n1673), .A1(asyncBusy), .Z(n2939));
Q_FDP0UA U3357 ( .D(n2939), .QTFCLK( ), .Q(asyncBusy));
Q_INV U3358 ( .A(gfifoOff), .Z(n2950));
Q_AO21 U3359 ( .A0(callEmuPre), .A1(n2950), .B0(initClock), .Z(n3002));
Q_OR02 U3360 ( .A0(mpEnable), .A1(bpHalt), .Z(n2958));
Q_INV U3361 ( .A(bpHalt), .Z(n2951));
Q_AN02 U3362 ( .A0(mpEnable), .A1(n2951), .Z(n2952));
Q_AO21 U3363 ( .A0(n2958), .A1(stopEmuPO), .B0(n2952), .Z(n2953));
Q_AN02 U3364 ( .A0(n2937), .A1(syncBp), .Z(n2959));
Q_AN02 U3365 ( .A0(n2953), .A1(n2959), .Z(n2965));
Q_AN02 U3366 ( .A0(active), .A1(n2940), .Z(n2966));
Q_AN02 U3367 ( .A0(n2966), .A1(n2941), .Z(n2962));
Q_OA21 U3368 ( .A0(n2965), .A1(n2962), .B0(n1406), .Z(n2942));
Q_OR02 U3369 ( .A0(n2962), .A1(callEmuPre), .Z(n2943));
Q_INV U3370 ( .A(n2941), .Z(n2972));
Q_AN02 U3371 ( .A0(n2972), .A1(mpEnable), .Z(n2956));
Q_AO21 U3372 ( .A0(n2966), .A1(n2956), .B0(n2959), .Z(n2954));
Q_AO21 U3373 ( .A0(n2954), .A1(n1406), .B0(n2976), .Z(n2944));
Q_INV U3374 ( .A(ckgHoldPIi), .Z(n2955));
Q_AN02 U3375 ( .A0(callEmuPre), .A1(n2955), .Z(n2976));
Q_INV U3376 ( .A(mpEnable), .Z(n2971));
Q_NR02 U3377 ( .A0(n2956), .A1(n3001), .Z(n2973));
Q_OA21 U3378 ( .A0(n2937), .A1(n2973), .B0(n1406), .Z(n2957));
Q_ND02 U3379 ( .A0(n2958), .A1(n2959), .Z(n2960));
Q_AN02 U3380 ( .A0(n1406), .A1(n2960), .Z(n2961));
Q_OR02 U3381 ( .A0(callEmuPre), .A1(n2966), .Z(n2946));
Q_NR02 U3382 ( .A0(active), .A1(syncBp), .Z(n2963));
Q_OA21 U3383 ( .A0(n2963), .A1(n2962), .B0(n1406), .Z(n2964));
Q_OR02 U3384 ( .A0(n2965), .A1(callEmuPre), .Z(n2945));
Q_AO21 U3385 ( .A0(n2966), .A1(n2971), .B0(n2937), .Z(n2967));
Q_AN02 U3386 ( .A0(n1406), .A1(n2967), .Z(n2968));
Q_AN02 U3387 ( .A0(n1406), .A1(n3001), .Z(n2947));
Q_OR02 U3388 ( .A0(callEmuPre), .A1(active), .Z(n2969));
Q_AN02 U3389 ( .A0(n1406), .A1(active), .Z(n2974));
Q_AN03 U3390 ( .A0(n2940), .A1(n2970), .A2(n2974), .Z(n2948));
Q_NR02 U3391 ( .A0(n2941), .A1(mpEnable), .Z(n2970));
Q_INV U3392 ( .A(n2973), .Z(n2975));
Q_AO21 U3393 ( .A0(n2975), .A1(n2974), .B0(n2976), .Z(n2949));
Q_MX02 U3394 ( .S(n2942), .A0(syncBp), .A1(active), .Z(n2977));
Q_FDP0UA U3395 ( .D(n2977), .QTFCLK( ), .Q(syncBp));
Q_MX02 U3396 ( .S(n2943), .A0(active), .A1(callEmuPre), .Z(n2978));
Q_FDP0UA U3397 ( .D(n2978), .QTFCLK( ), .Q(active));
Q_MX02 U3398 ( .S(n2944), .A0(simTimeOn), .A1(n2969), .Z(n2979));
Q_FDP0UA U3399 ( .D(n2979), .QTFCLK( ), .Q(simTimeOn));
Q_MX02 U3400 ( .S(n2961), .A0(callEmuPre), .A1(evalOnC), .Z(n2980));
Q_FDP0UA U3401 ( .D(n2980), .QTFCLK( ), .Q(evalOnC));
Q_MX02 U3402 ( .S(n2945), .A0(tbcPOd), .A1(n1406), .Z(n2981));
Q_FDP0UA U3403 ( .D(n2981), .QTFCLK( ), .Q(tbcPOd));
Q_FDP0UA U3404 ( .D(n2994), .QTFCLK( ), .Q(lbrOn));
Q_MX02 U3405 ( .S(n2957), .A0(n2993), .A1(fcnt[0]), .Z(n2982));
Q_FDP0UA U3406 ( .D(n2982), .QTFCLK( ), .Q(fcnt[0]));
Q_MX02 U3407 ( .S(n2957), .A0(n2992), .A1(fcnt[1]), .Z(n2983));
Q_FDP0UA U3408 ( .D(n2983), .QTFCLK( ), .Q(fcnt[1]));
Q_MX02 U3409 ( .S(n2957), .A0(n2991), .A1(fcnt[2]), .Z(n2984));
Q_FDP0UA U3410 ( .D(n2984), .QTFCLK( ), .Q(fcnt[2]));
Q_MX02 U3411 ( .S(n2946), .A0(tbcHold), .A1(n2990), .Z(n2985));
Q_FDP0UA U3412 ( .D(n2985), .QTFCLK( ), .Q(tbcHold));
Q_MX02 U3413 ( .S(n2964), .A0(n2987), .A1(mpOn), .Z(n2986));
Q_FDP0UA U3414 ( .D(n2986), .QTFCLK( ), .Q(mpOn));
Q_MX02 U3415 ( .S(n2946), .A0(n2988), .A1(n2989), .Z(n2987));
Q_NR02 U3416 ( .A0(n2968), .A1(n2998), .Z(n2988));
Q_MX02 U3417 ( .S(n2968), .A0(oneFclkEval), .A1(eClkHold), .Z(n2989));
Q_AN02 U3418 ( .A0(callEmuPre), .A1(tbcHoldPI), .Z(n2990));
Q_MX02 U3419 ( .S(n2947), .A0(fclkPerEval[2]), .A1(n2995), .Z(n2991));
Q_MX02 U3420 ( .S(n2947), .A0(fclkPerEval[1]), .A1(n2997), .Z(n2992));
Q_MX02 U3421 ( .S(n2947), .A0(fclkPerEval[0]), .A1(n2999), .Z(n2993));
Q_MX02 U3422 ( .S(n2948), .A0(n2949), .A1(eClkHold), .Z(n2994));
Q_XNR2 U3423 ( .A0(fcnt[2]), .A1(n2996), .Z(n2995));
Q_OR02 U3424 ( .A0(fcnt[1]), .A1(fcnt[0]), .Z(n2996));
Q_XNR2 U3425 ( .A0(fcnt[1]), .A1(fcnt[0]), .Z(n2997));
Q_OR03 U3426 ( .A0(n2999), .A1(fcnt[1]), .A2(fcnt[2]), .Z(n2998));
Q_INV U3427 ( .A(fcnt[0]), .Z(n2999));
Q_OR03 U3428 ( .A0(mioPOW_2[3]), .A1(mioPOW_2[2]), .A2(n3000), .Z(n2941));
Q_OR03 U3429 ( .A0(stop3), .A1(stopT), .A2(mioPOW_2[5]), .Z(n3000));
Q_INV U3430 ( .A(n3001), .Z(n2940));
Q_OR03 U3431 ( .A0(fcnt[0]), .A1(fcnt[1]), .A2(fcnt[2]), .Z(n3001));
Q_FDP0UA U3432 ( .D(n3002), .QTFCLK( ), .Q(initClock));
Q_FDP0UA U3433 ( .D(n3003), .QTFCLK( ), .Q(eClkR));
Q_XOR2 U3434 ( .A0(simTimeEnable), .A1(eClkR), .Z(n3003));
Q_INV U3435 ( .A(hotSwapOnPI), .Z(n3004));
Q_NR02 U3436 ( .A0(hotSwapOnPI), .A1(cakeCcEnable), .Z(n3005));
Q_MX02 U3437 ( .S(n3005), .A0(n3007), .A1(clockMC), .Z(n3006));
Q_FDP0UA U3438 ( .D(n3006), .QTFCLK( ), .Q(clockMC));
Q_MX02 U3439 ( .S(hotSwapOnPI), .A0(n3008), .A1(clockMCInit), .Z(n3007));
Q_INV U3440 ( .A(clockMC), .Z(n3008));
Q_NR02 U3441 ( .A0(n3010), .A1(n3009), .Z(n3011));
Q_FDP0UA U3442 ( .D(evalOnInt), .QTFCLK( ), .Q(evalOnIntR[0]));
Q_FDP0UA U3443 ( .D(evalOnIntR[0]), .QTFCLK( ), .Q(evalOnIntR[1]));
Q_FDP0UA U3444 ( .D(n3010), .QTFCLK( ), .Q(evalOnIntD));
Q_MX02 U3445 ( .S(n3011), .A0(n3027), .A1(evalOnDExt[0]), .Z(n3012));
Q_FDP0UA U3446 ( .D(n3012), .QTFCLK( ), .Q(evalOnDExt[0]));
Q_MX02 U3447 ( .S(n3011), .A0(n3026), .A1(evalOnDExt[1]), .Z(n3013));
Q_FDP0UA U3448 ( .D(n3013), .QTFCLK( ), .Q(evalOnDExt[1]));
Q_MX02 U3449 ( .S(n3011), .A0(n3025), .A1(evalOnDExt[2]), .Z(n3014));
Q_FDP0UA U3450 ( .D(n3014), .QTFCLK( ), .Q(evalOnDExt[2]));
Q_MX02 U3451 ( .S(n3011), .A0(n3024), .A1(evalOnDExt[3]), .Z(n3015));
Q_FDP0UA U3452 ( .D(n3015), .QTFCLK( ), .Q(evalOnDExt[3]));
Q_MX02 U3453 ( .S(n3011), .A0(n3023), .A1(evalOnDExt[4]), .Z(n3016));
Q_FDP0UA U3454 ( .D(n3016), .QTFCLK( ), .Q(evalOnDExt[4]));
Q_MX02 U3455 ( .S(n3011), .A0(n3022), .A1(evalOnDExt[5]), .Z(n3017));
Q_FDP0UA U3456 ( .D(n3017), .QTFCLK( ), .Q(evalOnDExt[5]));
Q_MX02 U3457 ( .S(n3011), .A0(n3021), .A1(evalOnDExt[6]), .Z(n3018));
Q_FDP0UA U3458 ( .D(n3018), .QTFCLK( ), .Q(evalOnDExt[6]));
Q_MX02 U3459 ( .S(n3011), .A0(n3020), .A1(evalOnDExt[7]), .Z(n3019));
Q_FDP0UA U3460 ( .D(n3019), .QTFCLK( ), .Q(evalOnDExt[7]));
Q_MX02 U3461 ( .S(n3010), .A0(n3028), .A1(evalOnDCtl[7]), .Z(n3020));
Q_MX02 U3462 ( .S(n3010), .A0(n3030), .A1(evalOnDCtl[6]), .Z(n3021));
Q_MX02 U3463 ( .S(n3010), .A0(n3032), .A1(evalOnDCtl[5]), .Z(n3022));
Q_MX02 U3464 ( .S(n3010), .A0(n3034), .A1(evalOnDCtl[4]), .Z(n3023));
Q_MX02 U3465 ( .S(n3010), .A0(n3036), .A1(evalOnDCtl[3]), .Z(n3024));
Q_MX02 U3466 ( .S(n3010), .A0(n3038), .A1(evalOnDCtl[2]), .Z(n3025));
Q_MX02 U3467 ( .S(n3010), .A0(n3040), .A1(evalOnDCtl[1]), .Z(n3026));
Q_MX02 U3468 ( .S(n3010), .A0(n3041), .A1(evalOnDCtl[0]), .Z(n3027));
Q_XNR2 U3469 ( .A0(evalOnDExt[7]), .A1(n3029), .Z(n3028));
Q_OR02 U3470 ( .A0(evalOnDExt[6]), .A1(n3031), .Z(n3029));
Q_XNR2 U3471 ( .A0(evalOnDExt[6]), .A1(n3031), .Z(n3030));
Q_OR02 U3472 ( .A0(evalOnDExt[5]), .A1(n3033), .Z(n3031));
Q_XNR2 U3473 ( .A0(evalOnDExt[5]), .A1(n3033), .Z(n3032));
Q_OR02 U3474 ( .A0(evalOnDExt[4]), .A1(n3035), .Z(n3033));
Q_XNR2 U3475 ( .A0(evalOnDExt[4]), .A1(n3035), .Z(n3034));
Q_OR02 U3476 ( .A0(evalOnDExt[3]), .A1(n3037), .Z(n3035));
Q_XNR2 U3477 ( .A0(evalOnDExt[3]), .A1(n3037), .Z(n3036));
Q_OR02 U3478 ( .A0(evalOnDExt[2]), .A1(n3039), .Z(n3037));
Q_XNR2 U3479 ( .A0(evalOnDExt[2]), .A1(n3039), .Z(n3038));
Q_OR02 U3480 ( .A0(evalOnDExt[1]), .A1(evalOnDExt[0]), .Z(n3039));
Q_XNR2 U3481 ( .A0(evalOnDExt[1]), .A1(evalOnDExt[0]), .Z(n3040));
Q_INV U3482 ( .A(evalOnDExt[0]), .Z(n3041));
Q_OR02 U3483 ( .A0(evalOnInt), .A1(evalOnIntR[0]), .Z(n3010));
Q_OR02 U3484 ( .A0(n3043), .A1(n3042), .Z(n3009));
Q_OR03 U3485 ( .A0(evalOnDExt[1]), .A1(evalOnDExt[0]), .A2(n3044), .Z(n3042));
Q_OR03 U3486 ( .A0(evalOnDExt[4]), .A1(evalOnDExt[3]), .A2(evalOnDExt[2]), .Z(n3043));
Q_OR03 U3487 ( .A0(evalOnDExt[7]), .A1(evalOnDExt[6]), .A2(evalOnDExt[5]), .Z(n3044));
Q_FDP0UA U3488 ( .D(evalOnC), .QTFCLK( ), .Q(evalOnD));
Q_FDP0UA U3489 ( .D(stopTL), .QTFCLK( ), .Q(stopTLd));
Q_FDP0UA U3490 ( .D(mioPOW_2[4]), .QTFCLK( ), .Q(stop3POd));
Q_FDP0UA U3491 ( .D(mioPOW_2[5]), .QTFCLK( ), .Q(stop4POd));
Q_FDP0UA U3492 ( .D(mioPOW_2[3]), .QTFCLK( ), .Q(stop2POd));
Q_FDP0UA U3493 ( .D(mioPOW_2[2]), .QTFCLK( ), .Q(stop1POd));
Q_FDP0UA U3494 ( .D(sdlStopRply), .QTFCLK( ), .Q(sdlStopRplyD));
Q_INV U3495 ( .A(hasGFIFO2), .Z(n3046));
Q_NR02 U3496 ( .A0(hasGFIFO1), .A1(hasGFIFO2), .Z(n3047));
Q_INV U3497 ( .A(n3047), .Z(n3045));
Q_MX02 U3498 ( .S(n3047), .A0(GFAck), .A1(gfifoAckWait[0]), .Z(n3048));
Q_FDP0UA U3499 ( .D(n3048), .QTFCLK( ), .Q(gfifoAckWait[0]));
Q_MX02 U3500 ( .S(n3047), .A0(gfifoAckWait[0]), .A1(gfifoAckWait[1]), .Z(n3049));
Q_FDP0UA U3501 ( .D(n3049), .QTFCLK( ), .Q(gfifoAckWait[1]));
Q_MX02 U3502 ( .S(n3047), .A0(gfifoAckWait[1]), .A1(gfifoAckWait[2]), .Z(n3050));
Q_FDP0UA U3503 ( .D(n3050), .QTFCLK( ), .Q(gfifoAckWait[2]));
Q_MX02 U3504 ( .S(n3047), .A0(n3060), .A1(gfifoAckWait[3]), .Z(n3051));
Q_FDP0UA U3505 ( .D(n3051), .QTFCLK( ), .Q(gfifoAckWait[3]));
Q_MX02 U3506 ( .S(n3047), .A0(n3059), .A1(gfifoAckWait[4]), .Z(n3052));
Q_FDP0UA U3507 ( .D(n3052), .QTFCLK( ), .Q(gfifoAckWait[4]));
Q_MX02 U3508 ( .S(n3047), .A0(n3058), .A1(gfifoAckWait[5]), .Z(n3053));
Q_FDP0UA U3509 ( .D(n3053), .QTFCLK( ), .Q(gfifoAckWait[5]));
Q_MX02 U3510 ( .S(n3047), .A0(n3057), .A1(gfifoAckWait[6]), .Z(n3054));
Q_FDP0UA U3511 ( .D(n3054), .QTFCLK( ), .Q(gfifoAckWait[6]));
Q_MX02 U3512 ( .S(n3047), .A0(n3056), .A1(gfifoAckWait[7]), .Z(n3055));
Q_FDP0UA U3513 ( .D(n3055), .QTFCLK( ), .Q(gfifoAckWait[7]));
Q_AN02 U3514 ( .A0(hasGFIFO1), .A1(gfifoAckWait[6]), .Z(n3056));
Q_AN02 U3515 ( .A0(hasGFIFO1), .A1(gfifoAckWait[5]), .Z(n3057));
Q_AN02 U3516 ( .A0(hasGFIFO1), .A1(gfifoAckWait[4]), .Z(n3058));
Q_AN02 U3517 ( .A0(hasGFIFO1), .A1(gfifoAckWait[3]), .Z(n3059));
Q_AN02 U3518 ( .A0(hasGFIFO1), .A1(gfifoAckWait[2]), .Z(n3060));
Q_FDP0UA U3519 ( .D(SFIFOLock2), .QTFCLK( ), .Q(SFIFOLock));
Q_FDP0UA U3520 ( .D(mioPOW_2[1]), .QTFCLK( ), .Q(tbcPOReg));
Q_FDP0UA U3521 ( .D(GFLBfull), .QTFCLK( ), .Q(GFLBfullD));
Q_FDP0UA U3522 ( .D(GFGBfullBw), .QTFCLK( ), .Q(GFGBfullBwD));
Q_FDP0UA U3523 ( .D(gfifoOff), .QTFCLK( ), .Q(gfifoOff));
Q_FDP0UA U3524 ( .D(gfifoAsyncOff), .QTFCLK( ), .Q(gfifoAsyncOff));
Q_FDP0UA U3525 ( .D(APPLY_PI), .QTFCLK( ), .Q(applyPiR));
Q_FDP0UA U3526 ( .D(FvUseOnly), .QTFCLK( ), .Q(FvUseOnlyR));
Q_FDP0UA U3527 ( .D(callEmuPIi), .QTFCLK( ), .Q(sendPO));
Q_FDP0UA U3528 ( .D(callEmuWaitN), .QTFCLK( ), .Q(callEmuWait));
Q_AO21 U3529 ( .A0(asyncCall), .A1(sfifoSyncMode), .B0(n3061), .Z(n3062));
Q_OR03 U3530 ( .A0(holdEcm), .A1(ptxBusy), .A2(isfWait), .Z(n3061));
Q_FDP0UA U3531 ( .D(n3062), .QTFCLK( ), .Q(callEmuWaitC));
Q_FDP0UA U3532 ( .D(sfifoSyncMode), .QTFCLK( ), .Q(sfifoSyncMode));
Q_FDP0UA U3533 ( .D(syncOtbChannels), .QTFCLK( ), .Q(syncOtbChannels));
Q_OR02 U3534 ( .A0(hotSwapOnPI), .A1(callEmuPre), .Z(n3063));
Q_FDP0UA U3535 ( .D(xc_mioOn), .QTFCLK( ), .Q(xc_mioOn));
Q_FDP0UA U3536 ( .D(maxAcCycle[0]), .QTFCLK( ), .Q(maxAcCycle[0]));
Q_FDP0UA U3537 ( .D(maxAcCycle[1]), .QTFCLK( ), .Q(maxAcCycle[1]));
Q_FDP0UA U3538 ( .D(maxAcCycle[2]), .QTFCLK( ), .Q(maxAcCycle[2]));
Q_FDP0UA U3539 ( .D(maxAcCycle[3]), .QTFCLK( ), .Q(maxAcCycle[3]));
Q_FDP0UA U3540 ( .D(maxAcCycle[4]), .QTFCLK( ), .Q(maxAcCycle[4]));
Q_FDP0UA U3541 ( .D(maxAcCycle[5]), .QTFCLK( ), .Q(maxAcCycle[5]));
Q_FDP0UA U3542 ( .D(maxAcCycle[6]), .QTFCLK( ), .Q(maxAcCycle[6]));
Q_FDP0UA U3543 ( .D(maxAcCycle[7]), .QTFCLK( ), .Q(maxAcCycle[7]));
Q_FDP0UA U3544 ( .D(maxAcCycle[8]), .QTFCLK( ), .Q(maxAcCycle[8]));
Q_FDP0UA U3545 ( .D(maxAcCycle[9]), .QTFCLK( ), .Q(maxAcCycle[9]));
Q_FDP0UA U3546 ( .D(maxAcCycle[10]), .QTFCLK( ), .Q(maxAcCycle[10]));
Q_FDP0UA U3547 ( .D(maxAcCycle[11]), .QTFCLK( ), .Q(maxAcCycle[11]));
Q_FDP0UA U3548 ( .D(maxAcCycle[12]), .QTFCLK( ), .Q(maxAcCycle[12]));
Q_FDP0UA U3549 ( .D(maxAcCycle[13]), .QTFCLK( ), .Q(maxAcCycle[13]));
Q_FDP0UA U3550 ( .D(maxAcCycle[14]), .QTFCLK( ), .Q(maxAcCycle[14]));
Q_FDP0UA U3551 ( .D(maxAcCycle[15]), .QTFCLK( ), .Q(maxAcCycle[15]));
Q_FDP0UA U3552 ( .D(maxBpCycle[0]), .QTFCLK( ), .Q(maxBpCycle[0]));
Q_FDP0UA U3553 ( .D(maxBpCycle[1]), .QTFCLK( ), .Q(maxBpCycle[1]));
Q_FDP0UA U3554 ( .D(maxBpCycle[2]), .QTFCLK( ), .Q(maxBpCycle[2]));
Q_FDP0UA U3555 ( .D(maxBpCycle[3]), .QTFCLK( ), .Q(maxBpCycle[3]));
Q_FDP0UA U3556 ( .D(maxBpCycle[4]), .QTFCLK( ), .Q(maxBpCycle[4]));
Q_FDP0UA U3557 ( .D(maxBpCycle[5]), .QTFCLK( ), .Q(maxBpCycle[5]));
Q_FDP0UA U3558 ( .D(maxBpCycle[6]), .QTFCLK( ), .Q(maxBpCycle[6]));
Q_FDP0UA U3559 ( .D(maxBpCycle[7]), .QTFCLK( ), .Q(maxBpCycle[7]));
Q_FDP0UA U3560 ( .D(maxBpCycle[8]), .QTFCLK( ), .Q(maxBpCycle[8]));
Q_FDP0UA U3561 ( .D(maxBpCycle[9]), .QTFCLK( ), .Q(maxBpCycle[9]));
Q_FDP0UA U3562 ( .D(maxBpCycle[10]), .QTFCLK( ), .Q(maxBpCycle[10]));
Q_FDP0UA U3563 ( .D(maxBpCycle[11]), .QTFCLK( ), .Q(maxBpCycle[11]));
Q_FDP0UA U3564 ( .D(maxBpCycle[12]), .QTFCLK( ), .Q(maxBpCycle[12]));
Q_FDP0UA U3565 ( .D(maxBpCycle[13]), .QTFCLK( ), .Q(maxBpCycle[13]));
Q_FDP0UA U3566 ( .D(maxBpCycle[14]), .QTFCLK( ), .Q(maxBpCycle[14]));
Q_FDP0UA U3567 ( .D(maxBpCycle[15]), .QTFCLK( ), .Q(maxBpCycle[15]));
Q_FDP0UA U3568 ( .D(forceAbort), .QTFCLK( ), .Q(forceAbort));
Q_FDP0UA U3569 ( .D(xcRecordOn), .QTFCLK( ), .Q(xcRecordOn));
Q_FDP0UA U3570 ( .D(xcReplayOn), .QTFCLK( ), .Q(xcReplayOn));
Q_FDP0UA U3571 ( .D(evalOnDCtl[0]), .QTFCLK( ), .Q(evalOnDCtl[0]));
Q_FDP0UA U3572 ( .D(evalOnDCtl[1]), .QTFCLK( ), .Q(evalOnDCtl[1]));
Q_FDP0UA U3573 ( .D(evalOnDCtl[2]), .QTFCLK( ), .Q(evalOnDCtl[2]));
Q_FDP0UA U3574 ( .D(evalOnDCtl[3]), .QTFCLK( ), .Q(evalOnDCtl[3]));
Q_FDP0UA U3575 ( .D(evalOnDCtl[4]), .QTFCLK( ), .Q(evalOnDCtl[4]));
Q_FDP0UA U3576 ( .D(evalOnDCtl[5]), .QTFCLK( ), .Q(evalOnDCtl[5]));
Q_FDP0UA U3577 ( .D(evalOnDCtl[6]), .QTFCLK( ), .Q(evalOnDCtl[6]));
Q_FDP0UA U3578 ( .D(evalOnDCtl[7]), .QTFCLK( ), .Q(evalOnDCtl[7]));
Q_FDP0UA U3579 ( .D(gfPushFill[0]), .QTFCLK( ), .Q(gfPushFill[0]));
Q_FDP0UA U3580 ( .D(gfPushFill[1]), .QTFCLK( ), .Q(gfPushFill[1]));
Q_FDP0UA U3581 ( .D(gfPushFill[2]), .QTFCLK( ), .Q(gfPushFill[2]));
Q_FDP0UA U3582 ( .D(gfPushFill[3]), .QTFCLK( ), .Q(gfPushFill[3]));
Q_FDP0UA U3583 ( .D(gfPushDly[0]), .QTFCLK( ), .Q(gfPushDly[0]));
Q_FDP0UA U3584 ( .D(gfPushDly[1]), .QTFCLK( ), .Q(gfPushDly[1]));
Q_FDP0UA U3585 ( .D(gfPushDly[2]), .QTFCLK( ), .Q(gfPushDly[2]));
Q_FDP0UA U3586 ( .D(gfPushDly[3]), .QTFCLK( ), .Q(gfPushDly[3]));
Q_FDP0UA U3587 ( .D(gfPushDly[4]), .QTFCLK( ), .Q(gfPushDly[4]));
Q_FDP0UA U3588 ( .D(gfPushDly[5]), .QTFCLK( ), .Q(gfPushDly[5]));
Q_FDP0UA U3589 ( .D(gfPushDly[6]), .QTFCLK( ), .Q(gfPushDly[6]));
Q_FDP0UA U3590 ( .D(gfPushDly[7]), .QTFCLK( ), .Q(gfPushDly[7]));
Q_FDP0UA U3591 ( .D(fclkPerEval[0]), .QTFCLK( ), .Q(fclkPerEval[0]));
Q_FDP0UA U3592 ( .D(fclkPerEval[1]), .QTFCLK( ), .Q(fclkPerEval[1]));
Q_FDP0UA U3593 ( .D(fclkPerEval[2]), .QTFCLK( ), .Q(fclkPerEval[2]));
Q_FDP0UA U3594 ( .D(fclkPerEval[3]), .QTFCLK( ), .Q(fclkPerEval[3]));
Q_FDP0UA U3595 ( .D(fclkPerEval[4]), .QTFCLK( ), .Q(fclkPerEval[4]));
Q_FDP0UA U3596 ( .D(fclkPerEval[5]), .QTFCLK( ), .Q(fclkPerEval[5]));
Q_FDP0UA U3597 ( .D(fclkPerEval[6]), .QTFCLK( ), .Q(fclkPerEval[6]));
Q_FDP0UA U3598 ( .D(fclkPerEval[7]), .QTFCLK( ), .Q(fclkPerEval[7]));
Q_OR02 U3599 ( .A0(n3063), .A1(ecmOne), .Z(n3064));
Q_FDP0UA U3600 ( .D(n3064), .QTFCLK( ), .Q(ecmOne));
Q_FDP0UA U3601 ( .D(hwClkDbgTime), .QTFCLK( ), .Q(hwClkDbgTime));
Q_FDP0UA U3602 ( .D(hwClkDbg), .QTFCLK( ), .Q(hwClkDbg));
Q_FDP0UA U3603 ( .D(tbcEnable), .QTFCLK( ), .Q(tbcEnable));
Q_FDP0UA U3604 ( .D(DccFrameMark[0]), .QTFCLK( ), .Q(DccFrameMark[0]));
Q_FDP0UA U3605 ( .D(DccFrameMark[1]), .QTFCLK( ), .Q(DccFrameMark[1]));
Q_FDP0UA U3606 ( .D(DccFrameMark[2]), .QTFCLK( ), .Q(DccFrameMark[2]));
Q_FDP0UA U3607 ( .D(DccFrameMark[3]), .QTFCLK( ), .Q(DccFrameMark[3]));
Q_FDP0UA U3608 ( .D(DccFrameMark[4]), .QTFCLK( ), .Q(DccFrameMark[4]));
Q_FDP0UA U3609 ( .D(DccFrameMark[5]), .QTFCLK( ), .Q(DccFrameMark[5]));
Q_FDP0UA U3610 ( .D(DccFrameMark[6]), .QTFCLK( ), .Q(DccFrameMark[6]));
Q_FDP0UA U3611 ( .D(DccFrameMark[7]), .QTFCLK( ), .Q(DccFrameMark[7]));
Q_FDP0UA U3612 ( .D(DccFrameCycle[0]), .QTFCLK( ), .Q(DccFrameCycle[0]));
Q_FDP0UA U3613 ( .D(DccFrameCycle[1]), .QTFCLK( ), .Q(DccFrameCycle[1]));
Q_FDP0UA U3614 ( .D(DccFrameCycle[2]), .QTFCLK( ), .Q(DccFrameCycle[2]));
Q_FDP0UA U3615 ( .D(DccFrameCycle[3]), .QTFCLK( ), .Q(DccFrameCycle[3]));
Q_FDP0UA U3616 ( .D(DccFrameCycle[4]), .QTFCLK( ), .Q(DccFrameCycle[4]));
Q_FDP0UA U3617 ( .D(DccFrameCycle[5]), .QTFCLK( ), .Q(DccFrameCycle[5]));
Q_FDP0UA U3618 ( .D(DccFrameCycle[6]), .QTFCLK( ), .Q(DccFrameCycle[6]));
Q_FDP0UA U3619 ( .D(DccFrameCycle[7]), .QTFCLK( ), .Q(DccFrameCycle[7]));
Q_FDP0UA U3620 ( .D(FvSimple2), .QTFCLK( ), .Q(FvSimple2));
Q_FDP0UA U3621 ( .D(sdlHaltHwClk), .QTFCLK( ), .Q(sdlHaltHwClk));
Q_FDP0UA U3622 ( .D(sdlEnable), .QTFCLK( ), .Q(sdlEnable));
Q_FDP0UA U3623 ( .D(hssReset), .QTFCLK( ), .Q(hssReset));
Q_FDP0UA U3624 ( .D(callEmuPIi), .QTFCLK( ), .Q(callEmuR));
Q_FDP0UA U3625 ( .D(ixc_time.nextDutTime[63]), .QTFCLK( ), .Q(nextDutTimeS[63]));
Q_FDP0UA U3626 ( .D(ixc_time.nextDutTime[62]), .QTFCLK( ), .Q(nextDutTimeS[62]));
Q_FDP0UA U3627 ( .D(ixc_time.nextDutTime[61]), .QTFCLK( ), .Q(nextDutTimeS[61]));
Q_FDP0UA U3628 ( .D(ixc_time.nextDutTime[60]), .QTFCLK( ), .Q(nextDutTimeS[60]));
Q_FDP0UA U3629 ( .D(ixc_time.nextDutTime[59]), .QTFCLK( ), .Q(nextDutTimeS[59]));
Q_FDP0UA U3630 ( .D(ixc_time.nextDutTime[58]), .QTFCLK( ), .Q(nextDutTimeS[58]));
Q_FDP0UA U3631 ( .D(ixc_time.nextDutTime[57]), .QTFCLK( ), .Q(nextDutTimeS[57]));
Q_FDP0UA U3632 ( .D(ixc_time.nextDutTime[56]), .QTFCLK( ), .Q(nextDutTimeS[56]));
Q_FDP0UA U3633 ( .D(ixc_time.nextDutTime[55]), .QTFCLK( ), .Q(nextDutTimeS[55]));
Q_FDP0UA U3634 ( .D(ixc_time.nextDutTime[54]), .QTFCLK( ), .Q(nextDutTimeS[54]));
Q_FDP0UA U3635 ( .D(ixc_time.nextDutTime[53]), .QTFCLK( ), .Q(nextDutTimeS[53]));
Q_FDP0UA U3636 ( .D(ixc_time.nextDutTime[52]), .QTFCLK( ), .Q(nextDutTimeS[52]));
Q_FDP0UA U3637 ( .D(ixc_time.nextDutTime[51]), .QTFCLK( ), .Q(nextDutTimeS[51]));
Q_FDP0UA U3638 ( .D(ixc_time.nextDutTime[50]), .QTFCLK( ), .Q(nextDutTimeS[50]));
Q_FDP0UA U3639 ( .D(ixc_time.nextDutTime[49]), .QTFCLK( ), .Q(nextDutTimeS[49]));
Q_FDP0UA U3640 ( .D(ixc_time.nextDutTime[48]), .QTFCLK( ), .Q(nextDutTimeS[48]));
Q_FDP0UA U3641 ( .D(ixc_time.nextDutTime[47]), .QTFCLK( ), .Q(nextDutTimeS[47]));
Q_FDP0UA U3642 ( .D(ixc_time.nextDutTime[46]), .QTFCLK( ), .Q(nextDutTimeS[46]));
Q_FDP0UA U3643 ( .D(ixc_time.nextDutTime[45]), .QTFCLK( ), .Q(nextDutTimeS[45]));
Q_FDP0UA U3644 ( .D(ixc_time.nextDutTime[44]), .QTFCLK( ), .Q(nextDutTimeS[44]));
Q_FDP0UA U3645 ( .D(ixc_time.nextDutTime[43]), .QTFCLK( ), .Q(nextDutTimeS[43]));
Q_FDP0UA U3646 ( .D(ixc_time.nextDutTime[42]), .QTFCLK( ), .Q(nextDutTimeS[42]));
Q_FDP0UA U3647 ( .D(ixc_time.nextDutTime[41]), .QTFCLK( ), .Q(nextDutTimeS[41]));
Q_FDP0UA U3648 ( .D(ixc_time.nextDutTime[40]), .QTFCLK( ), .Q(nextDutTimeS[40]));
Q_FDP0UA U3649 ( .D(ixc_time.nextDutTime[39]), .QTFCLK( ), .Q(nextDutTimeS[39]));
Q_FDP0UA U3650 ( .D(ixc_time.nextDutTime[38]), .QTFCLK( ), .Q(nextDutTimeS[38]));
Q_FDP0UA U3651 ( .D(ixc_time.nextDutTime[37]), .QTFCLK( ), .Q(nextDutTimeS[37]));
Q_FDP0UA U3652 ( .D(ixc_time.nextDutTime[36]), .QTFCLK( ), .Q(nextDutTimeS[36]));
Q_FDP0UA U3653 ( .D(ixc_time.nextDutTime[35]), .QTFCLK( ), .Q(nextDutTimeS[35]));
Q_FDP0UA U3654 ( .D(ixc_time.nextDutTime[34]), .QTFCLK( ), .Q(nextDutTimeS[34]));
Q_FDP0UA U3655 ( .D(ixc_time.nextDutTime[33]), .QTFCLK( ), .Q(nextDutTimeS[33]));
Q_FDP0UA U3656 ( .D(ixc_time.nextDutTime[32]), .QTFCLK( ), .Q(nextDutTimeS[32]));
Q_FDP0UA U3657 ( .D(ixc_time.nextDutTime[31]), .QTFCLK( ), .Q(nextDutTimeS[31]));
Q_FDP0UA U3658 ( .D(ixc_time.nextDutTime[30]), .QTFCLK( ), .Q(nextDutTimeS[30]));
Q_FDP0UA U3659 ( .D(ixc_time.nextDutTime[29]), .QTFCLK( ), .Q(nextDutTimeS[29]));
Q_FDP0UA U3660 ( .D(ixc_time.nextDutTime[28]), .QTFCLK( ), .Q(nextDutTimeS[28]));
Q_FDP0UA U3661 ( .D(ixc_time.nextDutTime[27]), .QTFCLK( ), .Q(nextDutTimeS[27]));
Q_FDP0UA U3662 ( .D(ixc_time.nextDutTime[26]), .QTFCLK( ), .Q(nextDutTimeS[26]));
Q_FDP0UA U3663 ( .D(ixc_time.nextDutTime[25]), .QTFCLK( ), .Q(nextDutTimeS[25]));
Q_FDP0UA U3664 ( .D(ixc_time.nextDutTime[24]), .QTFCLK( ), .Q(nextDutTimeS[24]));
Q_FDP0UA U3665 ( .D(ixc_time.nextDutTime[23]), .QTFCLK( ), .Q(nextDutTimeS[23]));
Q_FDP0UA U3666 ( .D(ixc_time.nextDutTime[22]), .QTFCLK( ), .Q(nextDutTimeS[22]));
Q_FDP0UA U3667 ( .D(ixc_time.nextDutTime[21]), .QTFCLK( ), .Q(nextDutTimeS[21]));
Q_FDP0UA U3668 ( .D(ixc_time.nextDutTime[20]), .QTFCLK( ), .Q(nextDutTimeS[20]));
Q_FDP0UA U3669 ( .D(ixc_time.nextDutTime[19]), .QTFCLK( ), .Q(nextDutTimeS[19]));
Q_FDP0UA U3670 ( .D(ixc_time.nextDutTime[18]), .QTFCLK( ), .Q(nextDutTimeS[18]));
Q_FDP0UA U3671 ( .D(ixc_time.nextDutTime[17]), .QTFCLK( ), .Q(nextDutTimeS[17]));
Q_FDP0UA U3672 ( .D(ixc_time.nextDutTime[16]), .QTFCLK( ), .Q(nextDutTimeS[16]));
Q_FDP0UA U3673 ( .D(ixc_time.nextDutTime[15]), .QTFCLK( ), .Q(nextDutTimeS[15]));
Q_FDP0UA U3674 ( .D(ixc_time.nextDutTime[14]), .QTFCLK( ), .Q(nextDutTimeS[14]));
Q_FDP0UA U3675 ( .D(ixc_time.nextDutTime[13]), .QTFCLK( ), .Q(nextDutTimeS[13]));
Q_FDP0UA U3676 ( .D(ixc_time.nextDutTime[12]), .QTFCLK( ), .Q(nextDutTimeS[12]));
Q_FDP0UA U3677 ( .D(ixc_time.nextDutTime[11]), .QTFCLK( ), .Q(nextDutTimeS[11]));
Q_FDP0UA U3678 ( .D(ixc_time.nextDutTime[10]), .QTFCLK( ), .Q(nextDutTimeS[10]));
Q_FDP0UA U3679 ( .D(ixc_time.nextDutTime[9]), .QTFCLK( ), .Q(nextDutTimeS[9]));
Q_FDP0UA U3680 ( .D(ixc_time.nextDutTime[8]), .QTFCLK( ), .Q(nextDutTimeS[8]));
Q_FDP0UA U3681 ( .D(ixc_time.nextDutTime[7]), .QTFCLK( ), .Q(nextDutTimeS[7]));
Q_FDP0UA U3682 ( .D(ixc_time.nextDutTime[6]), .QTFCLK( ), .Q(nextDutTimeS[6]));
Q_FDP0UA U3683 ( .D(ixc_time.nextDutTime[5]), .QTFCLK( ), .Q(nextDutTimeS[5]));
Q_FDP0UA U3684 ( .D(ixc_time.nextDutTime[4]), .QTFCLK( ), .Q(nextDutTimeS[4]));
Q_FDP0UA U3685 ( .D(ixc_time.nextDutTime[3]), .QTFCLK( ), .Q(nextDutTimeS[3]));
Q_FDP0UA U3686 ( .D(ixc_time.nextDutTime[2]), .QTFCLK( ), .Q(nextDutTimeS[2]));
Q_FDP0UA U3687 ( .D(ixc_time.nextDutTime[1]), .QTFCLK( ), .Q(nextDutTimeS[1]));
Q_FDP0UA U3688 ( .D(ixc_time.nextDutTime[0]), .QTFCLK( ), .Q(nextDutTimeS[0]));
Q_FDP0UA U3689 ( .D(n3065), .QTFCLK( ), .Q(mioPICntd));
Q_MX02 U3690 ( .S(xc_mioOn), .A0(mioPICntd), .A1(mioPICnt), .Z(n3065));
Q_INV U3691 ( .A(tbcPOmio), .Z(n3067));
Q_AN03 U3692 ( .A0(xc_mioOn), .A1(n3067), .A2(mioPOW_2[1]), .Z(n3066));
Q_XOR2 U3693 ( .A0(n3066), .A1(mioPOW_0[63]), .Z(n3068));
Q_FDP0UA U3694 ( .D(n3068), .QTFCLK( ), .Q(mioPOCnt));
Q_FDP0UA U3695 ( .D(mioPOW_2[1]), .QTFCLK( ), .Q(tbcPOmio));
Q_OR03 U3696 ( .A0(bpHalt), .A1(acHalt), .A2(forceAbort), .Z(n3075));
Q_INV U3697 ( .A(lockTrace), .Z(n3071));
Q_NR02 U3698 ( .A0(lockTrace), .A1(lockTraceC[2]), .Z(n3074));
Q_INV U3699 ( .A(lockTraceC[0]), .Z(n3072));
Q_NR02 U3700 ( .A0(lockTraceC[1]), .A1(lockTraceC[0]), .Z(n3073));
Q_AN02 U3701 ( .A0(n3074), .A1(n3073), .Z(n3077));
Q_AN02 U3702 ( .A0(n3077), .A1(n3075), .Z(n3069));
Q_INV U3703 ( .A(n3077), .Z(n3070));
Q_INV U3704 ( .A(n3075), .Z(n3076));
Q_MX02 U3705 ( .S(n3077), .A0(lockTrace), .A1(n3076), .Z(n3078));
Q_MX02 U3706 ( .S(n3069), .A0(lockTraceTime[0]), .A1(simTime[0]), .Z(n3079));
Q_FDP0UA U3707 ( .D(n3079), .QTFCLK( ), .Q(lockTraceTime[0]));
Q_MX02 U3708 ( .S(n3069), .A0(lockTraceTime[1]), .A1(simTime[1]), .Z(n3080));
Q_FDP0UA U3709 ( .D(n3080), .QTFCLK( ), .Q(lockTraceTime[1]));
Q_MX02 U3710 ( .S(n3069), .A0(lockTraceTime[2]), .A1(n3277), .Z(n3081));
Q_FDP0UA U3711 ( .D(n3081), .QTFCLK( ), .Q(lockTraceTime[2]));
Q_MX02 U3712 ( .S(n3069), .A0(lockTraceTime[3]), .A1(n3276), .Z(n3082));
Q_FDP0UA U3713 ( .D(n3082), .QTFCLK( ), .Q(lockTraceTime[3]));
Q_MX02 U3714 ( .S(n3069), .A0(lockTraceTime[4]), .A1(n3274), .Z(n3083));
Q_FDP0UA U3715 ( .D(n3083), .QTFCLK( ), .Q(lockTraceTime[4]));
Q_MX02 U3716 ( .S(n3069), .A0(lockTraceTime[5]), .A1(n3272), .Z(n3084));
Q_FDP0UA U3717 ( .D(n3084), .QTFCLK( ), .Q(lockTraceTime[5]));
Q_MX02 U3718 ( .S(n3069), .A0(lockTraceTime[6]), .A1(n3270), .Z(n3085));
Q_FDP0UA U3719 ( .D(n3085), .QTFCLK( ), .Q(lockTraceTime[6]));
Q_MX02 U3720 ( .S(n3069), .A0(lockTraceTime[7]), .A1(n3268), .Z(n3086));
Q_FDP0UA U3721 ( .D(n3086), .QTFCLK( ), .Q(lockTraceTime[7]));
Q_MX02 U3722 ( .S(n3069), .A0(lockTraceTime[8]), .A1(n3266), .Z(n3087));
Q_FDP0UA U3723 ( .D(n3087), .QTFCLK( ), .Q(lockTraceTime[8]));
Q_MX02 U3724 ( .S(n3069), .A0(lockTraceTime[9]), .A1(n3264), .Z(n3088));
Q_FDP0UA U3725 ( .D(n3088), .QTFCLK( ), .Q(lockTraceTime[9]));
Q_MX02 U3726 ( .S(n3069), .A0(lockTraceTime[10]), .A1(n3262), .Z(n3089));
Q_FDP0UA U3727 ( .D(n3089), .QTFCLK( ), .Q(lockTraceTime[10]));
Q_MX02 U3728 ( .S(n3069), .A0(lockTraceTime[11]), .A1(n3260), .Z(n3090));
Q_FDP0UA U3729 ( .D(n3090), .QTFCLK( ), .Q(lockTraceTime[11]));
Q_MX02 U3730 ( .S(n3069), .A0(lockTraceTime[12]), .A1(n3258), .Z(n3091));
Q_FDP0UA U3731 ( .D(n3091), .QTFCLK( ), .Q(lockTraceTime[12]));
Q_MX02 U3732 ( .S(n3069), .A0(lockTraceTime[13]), .A1(n3256), .Z(n3092));
Q_FDP0UA U3733 ( .D(n3092), .QTFCLK( ), .Q(lockTraceTime[13]));
Q_MX02 U3734 ( .S(n3069), .A0(lockTraceTime[14]), .A1(n3254), .Z(n3093));
Q_FDP0UA U3735 ( .D(n3093), .QTFCLK( ), .Q(lockTraceTime[14]));
Q_MX02 U3736 ( .S(n3069), .A0(lockTraceTime[15]), .A1(n3252), .Z(n3094));
Q_FDP0UA U3737 ( .D(n3094), .QTFCLK( ), .Q(lockTraceTime[15]));
Q_MX02 U3738 ( .S(n3069), .A0(lockTraceTime[16]), .A1(n3250), .Z(n3095));
Q_FDP0UA U3739 ( .D(n3095), .QTFCLK( ), .Q(lockTraceTime[16]));
Q_MX02 U3740 ( .S(n3069), .A0(lockTraceTime[17]), .A1(n3248), .Z(n3096));
Q_FDP0UA U3741 ( .D(n3096), .QTFCLK( ), .Q(lockTraceTime[17]));
Q_MX02 U3742 ( .S(n3069), .A0(lockTraceTime[18]), .A1(n3246), .Z(n3097));
Q_FDP0UA U3743 ( .D(n3097), .QTFCLK( ), .Q(lockTraceTime[18]));
Q_MX02 U3744 ( .S(n3069), .A0(lockTraceTime[19]), .A1(n3244), .Z(n3098));
Q_FDP0UA U3745 ( .D(n3098), .QTFCLK( ), .Q(lockTraceTime[19]));
Q_MX02 U3746 ( .S(n3069), .A0(lockTraceTime[20]), .A1(n3242), .Z(n3099));
Q_FDP0UA U3747 ( .D(n3099), .QTFCLK( ), .Q(lockTraceTime[20]));
Q_MX02 U3748 ( .S(n3069), .A0(lockTraceTime[21]), .A1(n3240), .Z(n3100));
Q_FDP0UA U3749 ( .D(n3100), .QTFCLK( ), .Q(lockTraceTime[21]));
Q_MX02 U3750 ( .S(n3069), .A0(lockTraceTime[22]), .A1(n3238), .Z(n3101));
Q_FDP0UA U3751 ( .D(n3101), .QTFCLK( ), .Q(lockTraceTime[22]));
Q_MX02 U3752 ( .S(n3069), .A0(lockTraceTime[23]), .A1(n3236), .Z(n3102));
Q_FDP0UA U3753 ( .D(n3102), .QTFCLK( ), .Q(lockTraceTime[23]));
Q_MX02 U3754 ( .S(n3069), .A0(lockTraceTime[24]), .A1(n3234), .Z(n3103));
Q_FDP0UA U3755 ( .D(n3103), .QTFCLK( ), .Q(lockTraceTime[24]));
Q_MX02 U3756 ( .S(n3069), .A0(lockTraceTime[25]), .A1(n3232), .Z(n3104));
Q_FDP0UA U3757 ( .D(n3104), .QTFCLK( ), .Q(lockTraceTime[25]));
Q_MX02 U3758 ( .S(n3069), .A0(lockTraceTime[26]), .A1(n3230), .Z(n3105));
Q_FDP0UA U3759 ( .D(n3105), .QTFCLK( ), .Q(lockTraceTime[26]));
Q_MX02 U3760 ( .S(n3069), .A0(lockTraceTime[27]), .A1(n3228), .Z(n3106));
Q_FDP0UA U3761 ( .D(n3106), .QTFCLK( ), .Q(lockTraceTime[27]));
Q_MX02 U3762 ( .S(n3069), .A0(lockTraceTime[28]), .A1(n3226), .Z(n3107));
Q_FDP0UA U3763 ( .D(n3107), .QTFCLK( ), .Q(lockTraceTime[28]));
Q_MX02 U3764 ( .S(n3069), .A0(lockTraceTime[29]), .A1(n3224), .Z(n3108));
Q_FDP0UA U3765 ( .D(n3108), .QTFCLK( ), .Q(lockTraceTime[29]));
Q_MX02 U3766 ( .S(n3069), .A0(lockTraceTime[30]), .A1(n3222), .Z(n3109));
Q_FDP0UA U3767 ( .D(n3109), .QTFCLK( ), .Q(lockTraceTime[30]));
Q_MX02 U3768 ( .S(n3069), .A0(lockTraceTime[31]), .A1(n3220), .Z(n3110));
Q_FDP0UA U3769 ( .D(n3110), .QTFCLK( ), .Q(lockTraceTime[31]));
Q_MX02 U3770 ( .S(n3069), .A0(lockTraceTime[32]), .A1(n3218), .Z(n3111));
Q_FDP0UA U3771 ( .D(n3111), .QTFCLK( ), .Q(lockTraceTime[32]));
Q_MX02 U3772 ( .S(n3069), .A0(lockTraceTime[33]), .A1(n3216), .Z(n3112));
Q_FDP0UA U3773 ( .D(n3112), .QTFCLK( ), .Q(lockTraceTime[33]));
Q_MX02 U3774 ( .S(n3069), .A0(lockTraceTime[34]), .A1(n3214), .Z(n3113));
Q_FDP0UA U3775 ( .D(n3113), .QTFCLK( ), .Q(lockTraceTime[34]));
Q_MX02 U3776 ( .S(n3069), .A0(lockTraceTime[35]), .A1(n3212), .Z(n3114));
Q_FDP0UA U3777 ( .D(n3114), .QTFCLK( ), .Q(lockTraceTime[35]));
Q_MX02 U3778 ( .S(n3069), .A0(lockTraceTime[36]), .A1(n3210), .Z(n3115));
Q_FDP0UA U3779 ( .D(n3115), .QTFCLK( ), .Q(lockTraceTime[36]));
Q_MX02 U3780 ( .S(n3069), .A0(lockTraceTime[37]), .A1(n3208), .Z(n3116));
Q_FDP0UA U3781 ( .D(n3116), .QTFCLK( ), .Q(lockTraceTime[37]));
Q_MX02 U3782 ( .S(n3069), .A0(lockTraceTime[38]), .A1(n3206), .Z(n3117));
Q_FDP0UA U3783 ( .D(n3117), .QTFCLK( ), .Q(lockTraceTime[38]));
Q_MX02 U3784 ( .S(n3069), .A0(lockTraceTime[39]), .A1(n3204), .Z(n3118));
Q_FDP0UA U3785 ( .D(n3118), .QTFCLK( ), .Q(lockTraceTime[39]));
Q_MX02 U3786 ( .S(n3069), .A0(lockTraceTime[40]), .A1(n3202), .Z(n3119));
Q_FDP0UA U3787 ( .D(n3119), .QTFCLK( ), .Q(lockTraceTime[40]));
Q_MX02 U3788 ( .S(n3069), .A0(lockTraceTime[41]), .A1(n3200), .Z(n3120));
Q_FDP0UA U3789 ( .D(n3120), .QTFCLK( ), .Q(lockTraceTime[41]));
Q_MX02 U3790 ( .S(n3069), .A0(lockTraceTime[42]), .A1(n3198), .Z(n3121));
Q_FDP0UA U3791 ( .D(n3121), .QTFCLK( ), .Q(lockTraceTime[42]));
Q_MX02 U3792 ( .S(n3069), .A0(lockTraceTime[43]), .A1(n3196), .Z(n3122));
Q_FDP0UA U3793 ( .D(n3122), .QTFCLK( ), .Q(lockTraceTime[43]));
Q_MX02 U3794 ( .S(n3069), .A0(lockTraceTime[44]), .A1(n3194), .Z(n3123));
Q_FDP0UA U3795 ( .D(n3123), .QTFCLK( ), .Q(lockTraceTime[44]));
Q_MX02 U3796 ( .S(n3069), .A0(lockTraceTime[45]), .A1(n3192), .Z(n3124));
Q_FDP0UA U3797 ( .D(n3124), .QTFCLK( ), .Q(lockTraceTime[45]));
Q_MX02 U3798 ( .S(n3069), .A0(lockTraceTime[46]), .A1(n3190), .Z(n3125));
Q_FDP0UA U3799 ( .D(n3125), .QTFCLK( ), .Q(lockTraceTime[46]));
Q_MX02 U3800 ( .S(n3069), .A0(lockTraceTime[47]), .A1(n3188), .Z(n3126));
Q_FDP0UA U3801 ( .D(n3126), .QTFCLK( ), .Q(lockTraceTime[47]));
Q_MX02 U3802 ( .S(n3069), .A0(lockTraceTime[48]), .A1(n3186), .Z(n3127));
Q_FDP0UA U3803 ( .D(n3127), .QTFCLK( ), .Q(lockTraceTime[48]));
Q_MX02 U3804 ( .S(n3069), .A0(lockTraceTime[49]), .A1(n3184), .Z(n3128));
Q_FDP0UA U3805 ( .D(n3128), .QTFCLK( ), .Q(lockTraceTime[49]));
Q_MX02 U3806 ( .S(n3069), .A0(lockTraceTime[50]), .A1(n3182), .Z(n3129));
Q_FDP0UA U3807 ( .D(n3129), .QTFCLK( ), .Q(lockTraceTime[50]));
Q_MX02 U3808 ( .S(n3069), .A0(lockTraceTime[51]), .A1(n3180), .Z(n3130));
Q_FDP0UA U3809 ( .D(n3130), .QTFCLK( ), .Q(lockTraceTime[51]));
Q_MX02 U3810 ( .S(n3069), .A0(lockTraceTime[52]), .A1(n3178), .Z(n3131));
Q_FDP0UA U3811 ( .D(n3131), .QTFCLK( ), .Q(lockTraceTime[52]));
Q_MX02 U3812 ( .S(n3069), .A0(lockTraceTime[53]), .A1(n3176), .Z(n3132));
Q_FDP0UA U3813 ( .D(n3132), .QTFCLK( ), .Q(lockTraceTime[53]));
Q_MX02 U3814 ( .S(n3069), .A0(lockTraceTime[54]), .A1(n3174), .Z(n3133));
Q_FDP0UA U3815 ( .D(n3133), .QTFCLK( ), .Q(lockTraceTime[54]));
Q_MX02 U3816 ( .S(n3069), .A0(lockTraceTime[55]), .A1(n3172), .Z(n3134));
Q_FDP0UA U3817 ( .D(n3134), .QTFCLK( ), .Q(lockTraceTime[55]));
Q_MX02 U3818 ( .S(n3069), .A0(lockTraceTime[56]), .A1(n3170), .Z(n3135));
Q_FDP0UA U3819 ( .D(n3135), .QTFCLK( ), .Q(lockTraceTime[56]));
Q_MX02 U3820 ( .S(n3069), .A0(lockTraceTime[57]), .A1(n3168), .Z(n3136));
Q_FDP0UA U3821 ( .D(n3136), .QTFCLK( ), .Q(lockTraceTime[57]));
Q_MX02 U3822 ( .S(n3069), .A0(lockTraceTime[58]), .A1(n3166), .Z(n3137));
Q_FDP0UA U3823 ( .D(n3137), .QTFCLK( ), .Q(lockTraceTime[58]));
Q_MX02 U3824 ( .S(n3069), .A0(lockTraceTime[59]), .A1(n3164), .Z(n3138));
Q_FDP0UA U3825 ( .D(n3138), .QTFCLK( ), .Q(lockTraceTime[59]));
Q_MX02 U3826 ( .S(n3069), .A0(lockTraceTime[60]), .A1(n3162), .Z(n3139));
Q_FDP0UA U3827 ( .D(n3139), .QTFCLK( ), .Q(lockTraceTime[60]));
Q_MX02 U3828 ( .S(n3069), .A0(lockTraceTime[61]), .A1(n3160), .Z(n3140));
Q_FDP0UA U3829 ( .D(n3140), .QTFCLK( ), .Q(lockTraceTime[61]));
Q_MX02 U3830 ( .S(n3069), .A0(lockTraceTime[62]), .A1(n3158), .Z(n3141));
Q_FDP0UA U3831 ( .D(n3141), .QTFCLK( ), .Q(lockTraceTime[62]));
Q_MX02 U3832 ( .S(n3069), .A0(lockTraceTime[63]), .A1(n3156), .Z(n3142));
Q_FDP0UA U3833 ( .D(n3142), .QTFCLK( ), .Q(lockTraceTime[63]));
Q_MX02 U3834 ( .S(n3078), .A0(n3150), .A1(lockTraceC[0]), .Z(n3143));
Q_FDP0UA U3835 ( .D(n3143), .QTFCLK( ), .Q(lockTraceC[0]));
Q_MX02 U3836 ( .S(n3078), .A0(n3149), .A1(lockTraceC[1]), .Z(n3144));
Q_FDP0UA U3837 ( .D(n3144), .QTFCLK( ), .Q(lockTraceC[1]));
Q_MX02 U3838 ( .S(n3078), .A0(n3148), .A1(lockTraceC[2]), .Z(n3145));
Q_FDP0UA U3839 ( .D(n3145), .QTFCLK( ), .Q(lockTraceC[2]));
Q_MX02 U3840 ( .S(n3078), .A0(n3147), .A1(lockTrace), .Z(n3146));
Q_FDP0UA U3841 ( .D(n3146), .QTFCLK( ), .Q(lockTraceC[3]));
Q_AN02 U3842 ( .A0(n3070), .A1(n3151), .Z(n3147));
Q_AN02 U3843 ( .A0(n3070), .A1(n3153), .Z(n3148));
Q_AN02 U3844 ( .A0(n3070), .A1(n3155), .Z(n3149));
Q_OR02 U3845 ( .A0(n3077), .A1(n3072), .Z(n3150));
Q_XOR2 U3846 ( .A0(lockTrace), .A1(n3152), .Z(n3151));
Q_AD01HF U3847 ( .A0(lockTraceC[2]), .B0(n3154), .S(n3153), .CO(n3152));
Q_AD01HF U3848 ( .A0(lockTraceC[1]), .B0(lockTraceC[0]), .S(n3155), .CO(n3154));
Q_XOR2 U3849 ( .A0(simTime[63]), .A1(n3157), .Z(n3156));
Q_AD01HF U3850 ( .A0(simTime[62]), .B0(n3159), .S(n3158), .CO(n3157));
Q_AD01HF U3851 ( .A0(simTime[61]), .B0(n3161), .S(n3160), .CO(n3159));
Q_AD01HF U3852 ( .A0(simTime[60]), .B0(n3163), .S(n3162), .CO(n3161));
Q_AD01HF U3853 ( .A0(simTime[59]), .B0(n3165), .S(n3164), .CO(n3163));
Q_AD01HF U3854 ( .A0(simTime[58]), .B0(n3167), .S(n3166), .CO(n3165));
Q_AD01HF U3855 ( .A0(simTime[57]), .B0(n3169), .S(n3168), .CO(n3167));
Q_AD01HF U3856 ( .A0(simTime[56]), .B0(n3171), .S(n3170), .CO(n3169));
Q_AD01HF U3857 ( .A0(simTime[55]), .B0(n3173), .S(n3172), .CO(n3171));
Q_AD01HF U3858 ( .A0(simTime[54]), .B0(n3175), .S(n3174), .CO(n3173));
Q_AD01HF U3859 ( .A0(simTime[53]), .B0(n3177), .S(n3176), .CO(n3175));
Q_AD01HF U3860 ( .A0(simTime[52]), .B0(n3179), .S(n3178), .CO(n3177));
Q_AD01HF U3861 ( .A0(simTime[51]), .B0(n3181), .S(n3180), .CO(n3179));
Q_AD01HF U3862 ( .A0(simTime[50]), .B0(n3183), .S(n3182), .CO(n3181));
Q_AD01HF U3863 ( .A0(simTime[49]), .B0(n3185), .S(n3184), .CO(n3183));
Q_AD01HF U3864 ( .A0(simTime[48]), .B0(n3187), .S(n3186), .CO(n3185));
Q_AD01HF U3865 ( .A0(simTime[47]), .B0(n3189), .S(n3188), .CO(n3187));
Q_AD01HF U3866 ( .A0(simTime[46]), .B0(n3191), .S(n3190), .CO(n3189));
Q_AD01HF U3867 ( .A0(simTime[45]), .B0(n3193), .S(n3192), .CO(n3191));
Q_AD01HF U3868 ( .A0(simTime[44]), .B0(n3195), .S(n3194), .CO(n3193));
Q_AD01HF U3869 ( .A0(simTime[43]), .B0(n3197), .S(n3196), .CO(n3195));
Q_AD01HF U3870 ( .A0(simTime[42]), .B0(n3199), .S(n3198), .CO(n3197));
Q_AD01HF U3871 ( .A0(simTime[41]), .B0(n3201), .S(n3200), .CO(n3199));
Q_AD01HF U3872 ( .A0(simTime[40]), .B0(n3203), .S(n3202), .CO(n3201));
Q_AD01HF U3873 ( .A0(simTime[39]), .B0(n3205), .S(n3204), .CO(n3203));
Q_AD01HF U3874 ( .A0(simTime[38]), .B0(n3207), .S(n3206), .CO(n3205));
Q_AD01HF U3875 ( .A0(simTime[37]), .B0(n3209), .S(n3208), .CO(n3207));
Q_AD01HF U3876 ( .A0(simTime[36]), .B0(n3211), .S(n3210), .CO(n3209));
Q_AD01HF U3877 ( .A0(simTime[35]), .B0(n3213), .S(n3212), .CO(n3211));
Q_AD01HF U3878 ( .A0(simTime[34]), .B0(n3215), .S(n3214), .CO(n3213));
Q_AD01HF U3879 ( .A0(simTime[33]), .B0(n3217), .S(n3216), .CO(n3215));
Q_AD01HF U3880 ( .A0(simTime[32]), .B0(n3219), .S(n3218), .CO(n3217));
Q_AD01HF U3881 ( .A0(simTime[31]), .B0(n3221), .S(n3220), .CO(n3219));
Q_AD01HF U3882 ( .A0(simTime[30]), .B0(n3223), .S(n3222), .CO(n3221));
Q_AD01HF U3883 ( .A0(simTime[29]), .B0(n3225), .S(n3224), .CO(n3223));
Q_AD01HF U3884 ( .A0(simTime[28]), .B0(n3227), .S(n3226), .CO(n3225));
Q_AD01HF U3885 ( .A0(simTime[27]), .B0(n3229), .S(n3228), .CO(n3227));
Q_AD01HF U3886 ( .A0(simTime[26]), .B0(n3231), .S(n3230), .CO(n3229));
Q_AD01HF U3887 ( .A0(simTime[25]), .B0(n3233), .S(n3232), .CO(n3231));
Q_AD01HF U3888 ( .A0(simTime[24]), .B0(n3235), .S(n3234), .CO(n3233));
Q_AD01HF U3889 ( .A0(simTime[23]), .B0(n3237), .S(n3236), .CO(n3235));
Q_AD01HF U3890 ( .A0(simTime[22]), .B0(n3239), .S(n3238), .CO(n3237));
Q_AD01HF U3891 ( .A0(simTime[21]), .B0(n3241), .S(n3240), .CO(n3239));
Q_AD01HF U3892 ( .A0(simTime[20]), .B0(n3243), .S(n3242), .CO(n3241));
Q_AD01HF U3893 ( .A0(simTime[19]), .B0(n3245), .S(n3244), .CO(n3243));
Q_AD01HF U3894 ( .A0(simTime[18]), .B0(n3247), .S(n3246), .CO(n3245));
Q_AD01HF U3895 ( .A0(simTime[17]), .B0(n3249), .S(n3248), .CO(n3247));
Q_AD01HF U3896 ( .A0(simTime[16]), .B0(n3251), .S(n3250), .CO(n3249));
Q_AD01HF U3897 ( .A0(simTime[15]), .B0(n3253), .S(n3252), .CO(n3251));
Q_AD01HF U3898 ( .A0(simTime[14]), .B0(n3255), .S(n3254), .CO(n3253));
Q_AD01HF U3899 ( .A0(simTime[13]), .B0(n3257), .S(n3256), .CO(n3255));
Q_AD01HF U3900 ( .A0(simTime[12]), .B0(n3259), .S(n3258), .CO(n3257));
Q_AD01HF U3901 ( .A0(simTime[11]), .B0(n3261), .S(n3260), .CO(n3259));
Q_AD01HF U3902 ( .A0(simTime[10]), .B0(n3263), .S(n3262), .CO(n3261));
Q_AD01HF U3903 ( .A0(simTime[9]), .B0(n3265), .S(n3264), .CO(n3263));
Q_AD01HF U3904 ( .A0(simTime[8]), .B0(n3267), .S(n3266), .CO(n3265));
Q_AD01HF U3905 ( .A0(simTime[7]), .B0(n3269), .S(n3268), .CO(n3267));
Q_AD01HF U3906 ( .A0(simTime[6]), .B0(n3271), .S(n3270), .CO(n3269));
Q_AD01HF U3907 ( .A0(simTime[5]), .B0(n3273), .S(n3272), .CO(n3271));
Q_AD01HF U3908 ( .A0(simTime[4]), .B0(n3275), .S(n3274), .CO(n3273));
Q_AD01HF U3909 ( .A0(simTime[3]), .B0(simTime[2]), .S(n3276), .CO(n3275));
Q_OR02 U3910 ( .A0(n3069), .A1(lockTraceOn), .Z(n3278));
Q_FDP0UA U3911 ( .D(n3278), .QTFCLK( ), .Q(lockTraceOn));
Q_AN02 U3912 ( .A0(asyncCall), .A1(acHalt), .Z(n3279));
Q_MX02 U3913 ( .S(n3279), .A0(n3311), .A1(aHaltCnt[0]), .Z(n3280));
Q_FDP0UA U3914 ( .D(n3280), .QTFCLK( ), .Q(aHaltCnt[0]));
Q_MX02 U3915 ( .S(n3279), .A0(n3310), .A1(aHaltCnt[1]), .Z(n3281));
Q_FDP0UA U3916 ( .D(n3281), .QTFCLK( ), .Q(aHaltCnt[1]));
Q_MX02 U3917 ( .S(n3279), .A0(n3309), .A1(aHaltCnt[2]), .Z(n3282));
Q_FDP0UA U3918 ( .D(n3282), .QTFCLK( ), .Q(aHaltCnt[2]));
Q_MX02 U3919 ( .S(n3279), .A0(n3308), .A1(aHaltCnt[3]), .Z(n3283));
Q_FDP0UA U3920 ( .D(n3283), .QTFCLK( ), .Q(aHaltCnt[3]));
Q_MX02 U3921 ( .S(n3279), .A0(n3307), .A1(aHaltCnt[4]), .Z(n3284));
Q_FDP0UA U3922 ( .D(n3284), .QTFCLK( ), .Q(aHaltCnt[4]));
Q_MX02 U3923 ( .S(n3279), .A0(n3306), .A1(aHaltCnt[5]), .Z(n3285));
Q_FDP0UA U3924 ( .D(n3285), .QTFCLK( ), .Q(aHaltCnt[5]));
Q_MX02 U3925 ( .S(n3279), .A0(n3305), .A1(aHaltCnt[6]), .Z(n3286));
Q_FDP0UA U3926 ( .D(n3286), .QTFCLK( ), .Q(aHaltCnt[6]));
Q_MX02 U3927 ( .S(n3279), .A0(n3304), .A1(aHaltCnt[7]), .Z(n3287));
Q_FDP0UA U3928 ( .D(n3287), .QTFCLK( ), .Q(aHaltCnt[7]));
Q_MX02 U3929 ( .S(n3279), .A0(n3303), .A1(aHaltCnt[8]), .Z(n3288));
Q_FDP0UA U3930 ( .D(n3288), .QTFCLK( ), .Q(aHaltCnt[8]));
Q_MX02 U3931 ( .S(n3279), .A0(n3302), .A1(aHaltCnt[9]), .Z(n3289));
Q_FDP0UA U3932 ( .D(n3289), .QTFCLK( ), .Q(aHaltCnt[9]));
Q_MX02 U3933 ( .S(n3279), .A0(n3301), .A1(aHaltCnt[10]), .Z(n3290));
Q_FDP0UA U3934 ( .D(n3290), .QTFCLK( ), .Q(aHaltCnt[10]));
Q_MX02 U3935 ( .S(n3279), .A0(n3300), .A1(aHaltCnt[11]), .Z(n3291));
Q_FDP0UA U3936 ( .D(n3291), .QTFCLK( ), .Q(aHaltCnt[11]));
Q_MX02 U3937 ( .S(n3279), .A0(n3299), .A1(aHaltCnt[12]), .Z(n3292));
Q_FDP0UA U3938 ( .D(n3292), .QTFCLK( ), .Q(aHaltCnt[12]));
Q_MX02 U3939 ( .S(n3279), .A0(n3298), .A1(aHaltCnt[13]), .Z(n3293));
Q_FDP0UA U3940 ( .D(n3293), .QTFCLK( ), .Q(aHaltCnt[13]));
Q_MX02 U3941 ( .S(n3279), .A0(n3297), .A1(aHaltCnt[14]), .Z(n3294));
Q_FDP0UA U3942 ( .D(n3294), .QTFCLK( ), .Q(aHaltCnt[14]));
Q_MX02 U3943 ( .S(n3279), .A0(n3296), .A1(aHaltCnt[15]), .Z(n3295));
Q_FDP0UA U3944 ( .D(n3295), .QTFCLK( ), .Q(aHaltCnt[15]));
Q_AN02 U3945 ( .A0(asyncCall), .A1(n3312), .Z(n3296));
Q_AN02 U3946 ( .A0(asyncCall), .A1(n3314), .Z(n3297));
Q_AN02 U3947 ( .A0(asyncCall), .A1(n3316), .Z(n3298));
Q_AN02 U3948 ( .A0(asyncCall), .A1(n3318), .Z(n3299));
Q_AN02 U3949 ( .A0(asyncCall), .A1(n3320), .Z(n3300));
Q_AN02 U3950 ( .A0(asyncCall), .A1(n3322), .Z(n3301));
Q_AN02 U3951 ( .A0(asyncCall), .A1(n3324), .Z(n3302));
Q_AN02 U3952 ( .A0(asyncCall), .A1(n3326), .Z(n3303));
Q_AN02 U3953 ( .A0(asyncCall), .A1(n3328), .Z(n3304));
Q_AN02 U3954 ( .A0(asyncCall), .A1(n3330), .Z(n3305));
Q_AN02 U3955 ( .A0(asyncCall), .A1(n3332), .Z(n3306));
Q_AN02 U3956 ( .A0(asyncCall), .A1(n3334), .Z(n3307));
Q_AN02 U3957 ( .A0(asyncCall), .A1(n3336), .Z(n3308));
Q_AN02 U3958 ( .A0(asyncCall), .A1(n3338), .Z(n3309));
Q_AN02 U3959 ( .A0(asyncCall), .A1(n3340), .Z(n3310));
Q_AN02 U3960 ( .A0(asyncCall), .A1(n3341), .Z(n3311));
Q_XOR2 U3961 ( .A0(aHaltCnt[15]), .A1(n3313), .Z(n3312));
Q_AD01HF U3962 ( .A0(aHaltCnt[14]), .B0(n3315), .S(n3314), .CO(n3313));
Q_AD01HF U3963 ( .A0(aHaltCnt[13]), .B0(n3317), .S(n3316), .CO(n3315));
Q_AD01HF U3964 ( .A0(aHaltCnt[12]), .B0(n3319), .S(n3318), .CO(n3317));
Q_AD01HF U3965 ( .A0(aHaltCnt[11]), .B0(n3321), .S(n3320), .CO(n3319));
Q_AD01HF U3966 ( .A0(aHaltCnt[10]), .B0(n3323), .S(n3322), .CO(n3321));
Q_AD01HF U3967 ( .A0(aHaltCnt[9]), .B0(n3325), .S(n3324), .CO(n3323));
Q_AD01HF U3968 ( .A0(aHaltCnt[8]), .B0(n3327), .S(n3326), .CO(n3325));
Q_AD01HF U3969 ( .A0(aHaltCnt[7]), .B0(n3329), .S(n3328), .CO(n3327));
Q_AD01HF U3970 ( .A0(aHaltCnt[6]), .B0(n3331), .S(n3330), .CO(n3329));
Q_AD01HF U3971 ( .A0(aHaltCnt[5]), .B0(n3333), .S(n3332), .CO(n3331));
Q_AD01HF U3972 ( .A0(aHaltCnt[4]), .B0(n3335), .S(n3334), .CO(n3333));
Q_AD01HF U3973 ( .A0(aHaltCnt[3]), .B0(n3337), .S(n3336), .CO(n3335));
Q_AD01HF U3974 ( .A0(aHaltCnt[2]), .B0(n3339), .S(n3338), .CO(n3337));
Q_AD01HF U3975 ( .A0(aHaltCnt[1]), .B0(aHaltCnt[0]), .S(n3340), .CO(n3339));
Q_INV U3976 ( .A(aHaltCnt[0]), .Z(n3341));
Q_INV U3977 ( .A(evalOnInt), .Z(n3342));
Q_OA21 U3978 ( .A0(n3342), .A1(bpHalt), .B0(n2915), .Z(n3343));
Q_MX02 U3979 ( .S(n3343), .A0(n3375), .A1(bHaltCnt[0]), .Z(n3344));
Q_FDP0UA U3980 ( .D(n3344), .QTFCLK( ), .Q(bHaltCnt[0]));
Q_MX02 U3981 ( .S(n3343), .A0(n3374), .A1(bHaltCnt[1]), .Z(n3345));
Q_FDP0UA U3982 ( .D(n3345), .QTFCLK( ), .Q(bHaltCnt[1]));
Q_MX02 U3983 ( .S(n3343), .A0(n3373), .A1(bHaltCnt[2]), .Z(n3346));
Q_FDP0UA U3984 ( .D(n3346), .QTFCLK( ), .Q(bHaltCnt[2]));
Q_MX02 U3985 ( .S(n3343), .A0(n3372), .A1(bHaltCnt[3]), .Z(n3347));
Q_FDP0UA U3986 ( .D(n3347), .QTFCLK( ), .Q(bHaltCnt[3]));
Q_MX02 U3987 ( .S(n3343), .A0(n3371), .A1(bHaltCnt[4]), .Z(n3348));
Q_FDP0UA U3988 ( .D(n3348), .QTFCLK( ), .Q(bHaltCnt[4]));
Q_MX02 U3989 ( .S(n3343), .A0(n3370), .A1(bHaltCnt[5]), .Z(n3349));
Q_FDP0UA U3990 ( .D(n3349), .QTFCLK( ), .Q(bHaltCnt[5]));
Q_MX02 U3991 ( .S(n3343), .A0(n3369), .A1(bHaltCnt[6]), .Z(n3350));
Q_FDP0UA U3992 ( .D(n3350), .QTFCLK( ), .Q(bHaltCnt[6]));
Q_MX02 U3993 ( .S(n3343), .A0(n3368), .A1(bHaltCnt[7]), .Z(n3351));
Q_FDP0UA U3994 ( .D(n3351), .QTFCLK( ), .Q(bHaltCnt[7]));
Q_MX02 U3995 ( .S(n3343), .A0(n3367), .A1(bHaltCnt[8]), .Z(n3352));
Q_FDP0UA U3996 ( .D(n3352), .QTFCLK( ), .Q(bHaltCnt[8]));
Q_MX02 U3997 ( .S(n3343), .A0(n3366), .A1(bHaltCnt[9]), .Z(n3353));
Q_FDP0UA U3998 ( .D(n3353), .QTFCLK( ), .Q(bHaltCnt[9]));
Q_MX02 U3999 ( .S(n3343), .A0(n3365), .A1(bHaltCnt[10]), .Z(n3354));
Q_FDP0UA U4000 ( .D(n3354), .QTFCLK( ), .Q(bHaltCnt[10]));
Q_MX02 U4001 ( .S(n3343), .A0(n3364), .A1(bHaltCnt[11]), .Z(n3355));
Q_FDP0UA U4002 ( .D(n3355), .QTFCLK( ), .Q(bHaltCnt[11]));
Q_MX02 U4003 ( .S(n3343), .A0(n3363), .A1(bHaltCnt[12]), .Z(n3356));
Q_FDP0UA U4004 ( .D(n3356), .QTFCLK( ), .Q(bHaltCnt[12]));
Q_MX02 U4005 ( .S(n3343), .A0(n3362), .A1(bHaltCnt[13]), .Z(n3357));
Q_FDP0UA U4006 ( .D(n3357), .QTFCLK( ), .Q(bHaltCnt[13]));
Q_MX02 U4007 ( .S(n3343), .A0(n3361), .A1(bHaltCnt[14]), .Z(n3358));
Q_FDP0UA U4008 ( .D(n3358), .QTFCLK( ), .Q(bHaltCnt[14]));
Q_MX02 U4009 ( .S(n3343), .A0(n3360), .A1(bHaltCnt[15]), .Z(n3359));
Q_FDP0UA U4010 ( .D(n3359), .QTFCLK( ), .Q(bHaltCnt[15]));
Q_AN02 U4011 ( .A0(n2915), .A1(n3376), .Z(n3360));
Q_AN02 U4012 ( .A0(n2915), .A1(n3378), .Z(n3361));
Q_AN02 U4013 ( .A0(n2915), .A1(n3380), .Z(n3362));
Q_AN02 U4014 ( .A0(n2915), .A1(n3382), .Z(n3363));
Q_AN02 U4015 ( .A0(n2915), .A1(n3384), .Z(n3364));
Q_AN02 U4016 ( .A0(n2915), .A1(n3386), .Z(n3365));
Q_AN02 U4017 ( .A0(n2915), .A1(n3388), .Z(n3366));
Q_AN02 U4018 ( .A0(n2915), .A1(n3390), .Z(n3367));
Q_AN02 U4019 ( .A0(n2915), .A1(n3392), .Z(n3368));
Q_AN02 U4020 ( .A0(n2915), .A1(n3394), .Z(n3369));
Q_AN02 U4021 ( .A0(n2915), .A1(n3396), .Z(n3370));
Q_AN02 U4022 ( .A0(n2915), .A1(n3398), .Z(n3371));
Q_AN02 U4023 ( .A0(n2915), .A1(n3400), .Z(n3372));
Q_AN02 U4024 ( .A0(n2915), .A1(n3402), .Z(n3373));
Q_AN02 U4025 ( .A0(n2915), .A1(n3404), .Z(n3374));
Q_NR02 U4026 ( .A0(mpOn), .A1(bHaltCnt[0]), .Z(n3375));
Q_XOR2 U4027 ( .A0(bHaltCnt[15]), .A1(n3377), .Z(n3376));
Q_AD01HF U4028 ( .A0(bHaltCnt[14]), .B0(n3379), .S(n3378), .CO(n3377));
Q_AD01HF U4029 ( .A0(bHaltCnt[13]), .B0(n3381), .S(n3380), .CO(n3379));
Q_AD01HF U4030 ( .A0(bHaltCnt[12]), .B0(n3383), .S(n3382), .CO(n3381));
Q_AD01HF U4031 ( .A0(bHaltCnt[11]), .B0(n3385), .S(n3384), .CO(n3383));
Q_AD01HF U4032 ( .A0(bHaltCnt[10]), .B0(n3387), .S(n3386), .CO(n3385));
Q_AD01HF U4033 ( .A0(bHaltCnt[9]), .B0(n3389), .S(n3388), .CO(n3387));
Q_AD01HF U4034 ( .A0(bHaltCnt[8]), .B0(n3391), .S(n3390), .CO(n3389));
Q_AD01HF U4035 ( .A0(bHaltCnt[7]), .B0(n3393), .S(n3392), .CO(n3391));
Q_AD01HF U4036 ( .A0(bHaltCnt[6]), .B0(n3395), .S(n3394), .CO(n3393));
Q_AD01HF U4037 ( .A0(bHaltCnt[5]), .B0(n3397), .S(n3396), .CO(n3395));
Q_AD01HF U4038 ( .A0(bHaltCnt[4]), .B0(n3399), .S(n3398), .CO(n3397));
Q_AD01HF U4039 ( .A0(bHaltCnt[3]), .B0(n3401), .S(n3400), .CO(n3399));
Q_AD01HF U4040 ( .A0(bHaltCnt[2]), .B0(n3403), .S(n3402), .CO(n3401));
Q_AD01HF U4041 ( .A0(bHaltCnt[1]), .B0(bHaltCnt[0]), .S(n3404), .CO(n3403));
Q_FDP0UA U4042 ( .D(n3406), .QTFCLK( ), .Q(cakeUcEnable));
Q_OR02 U4043 ( .A0(simTimeEnable), .A1(cakeUcEnable), .Z(n3406));
Q_AN02 U4044 ( .A0(active), .A1(holdEcm), .Z(holdEcmC));
Q_NR02 U4045 ( .A0(n3001), .A1(n2941), .Z(n3407));
Q_AN03 U4046 ( .A0(n2974), .A1(n3407), .A2(mpEnable), .Z(n3408));
Q_MX02 U4047 ( .S(callEmuPre), .A0(n3408), .A1(n2955), .Z(simTimeEnable));
Q_OR02 U4048 ( .A0(callEmuPre), .A1(stopSDL), .Z(n3409));
Q_INV U4049 ( .A(cpfStop), .Z(n3410));
Q_LSN01 U4050 ( .S(n3410), .R(n1406), .Q(stopCPFPO), .QN( ));
Q_OR03 U4051 ( .A0(mioPOW_2[7]), .A1(stopEmuPO), .A2(n3411), .Z(stop3));
Q_OR03 U4052 ( .A0(bpHalt), .A1(mioPOW_2[6]), .A2(mioPOW_2[8]), .Z(n3411));
Q_LDP0 stopSDLPO_REG  ( .G(n3409), .D(stopSDL), .Q(stopSDLPO), .QN( ));
Q_MX02 U4054 ( .S(oneStepPIi), .A0(ixc_time.stopEcm), .A1(mpOn), .Z(stopT));
Q_AO21 U4055 ( .A0(lastDelta), .A1(evalOnC), .B0(hotSwapOnPI), .Z(mpSampleOv));
Q_OR02 U4056 ( .A0(evalOnC), .A1(hotSwapOnPI), .Z(eventOnR));
Q_AN02 U4057 ( .A0(dbiEvent), .A1(n3555), .Z(FvUseOnly));
Q_OR03 U4058 ( .A0(evalOnInt), .A1(n3412), .A2(n3009), .Z(evalOn));
Q_AN02 U4059 ( .A0(evalOnIntD), .A1(n3427), .Z(n3412));
Q_AN03 U4060 ( .A0(sdlEnable), .A1(sdlStop), .A2(xcReplayOn), .Z(sdlStopRply));
Q_AN03 U4061 ( .A0(sdlEnable), .A1(sdlStop), .A2(n3413), .Z(stopSDL));
Q_INV U4062 ( .A(xcReplayOn), .Z(n3413));
Q_AN02 U4063 ( .A0(stop4), .A1(tbcEnable), .Z(stop4R));
Q_AN02 U4064 ( .A0(stop2), .A1(tbcEnable), .Z(stop2R));
Q_AN02 U4065 ( .A0(stop1), .A1(tbcEnable), .Z(stop1R));
Q_AN02 U4066 ( .A0(n3071), .A1(n3414), .Z(evalOnInt));
Q_OR03 U4067 ( .A0(FTcallW), .A1(evalOnSync), .A2(lockTraceOn), .Z(n3414));
Q_INV U4068 ( .A(sdlStopRplyD), .Z(n3415));
Q_OA21 U4069 ( .A0(evalOnOrig), .A1(GFbusyW), .B0(n3415), .Z(evalOnSync));
Q_OR03 U4070 ( .A0(hwClkDbgOn), .A1(evalOnC), .A2(callEmuPre), .Z(n3416));
Q_AO21 U4071 ( .A0(tbcPOd), .A1(n3417), .B0(n3416), .Z(evalOnOrig));
Q_INV U4072 ( .A(mioPOW_2[1]), .Z(n3417));
Q_AN02 U4073 ( .A0(n3418), .A1(n3427), .Z(GFbusyW));
Q_OR03 U4074 ( .A0(dbiEvent), .A1(n3420), .A2(n3419), .Z(n3418));
Q_OR03 U4075 ( .A0(isfWait), .A1(gfifoWait), .A2(ptxBusy), .Z(n3419));
Q_OR03 U4076 ( .A0(callEmuWait), .A1(callEmuEv), .A2(osfWait), .Z(n3420));
Q_AN03 U4077 ( .A0(n3421), .A1(APPLY_PI), .A2(n3004), .Z(dbiEvent));
Q_INV U4078 ( .A(applyPiR), .Z(n3421));
Q_OR03 U4079 ( .A0(svAsyncCall), .A1(n3422), .A2(n3423), .Z(FTcallW));
Q_OR03 U4080 ( .A0(ecmHoldBusy), .A1(GFAck), .A2(otbAsyncCall), .Z(n3422));
Q_OR02 U4081 ( .A0(n3425), .A1(n3424), .Z(n3423));
Q_OR03 U4082 ( .A0(gfifoAckWait[1]), .A1(gfifoAckWait[0]), .A2(n3426), .Z(n3424));
Q_OR03 U4083 ( .A0(gfifoAckWait[4]), .A1(gfifoAckWait[3]), .A2(gfifoAckWait[2]), .Z(n3425));
Q_OR03 U4084 ( .A0(gfifoAckWait[7]), .A1(gfifoAckWait[6]), .A2(gfifoAckWait[5]), .Z(n3426));
Q_INV U4085 ( .A(FvSimple2), .Z(n3427));
Q_AD01HF U4086 ( .A0(uClkCntr[1]), .B0(uClkCntr[0]), .S(n3428), .CO(n3429));
Q_AD01HF U4087 ( .A0(uClkCntr[2]), .B0(n3429), .S(n3430), .CO(n3431));
Q_AD01HF U4088 ( .A0(uClkCntr[3]), .B0(n3431), .S(n3432), .CO(n3433));
Q_AD01HF U4089 ( .A0(uClkCntr[4]), .B0(n3433), .S(n3434), .CO(n3435));
Q_AD01HF U4090 ( .A0(uClkCntr[5]), .B0(n3435), .S(n3436), .CO(n3437));
Q_AD01HF U4091 ( .A0(uClkCntr[6]), .B0(n3437), .S(n3438), .CO(n3439));
Q_AD01HF U4092 ( .A0(uClkCntr[7]), .B0(n3439), .S(n3440), .CO(n3441));
Q_AD01HF U4093 ( .A0(uClkCntr[8]), .B0(n3441), .S(n3442), .CO(n3443));
Q_AD01HF U4094 ( .A0(uClkCntr[9]), .B0(n3443), .S(n3444), .CO(n3445));
Q_AD01HF U4095 ( .A0(uClkCntr[10]), .B0(n3445), .S(n3446), .CO(n3447));
Q_AD01HF U4096 ( .A0(uClkCntr[11]), .B0(n3447), .S(n3448), .CO(n3449));
Q_AD01HF U4097 ( .A0(uClkCntr[12]), .B0(n3449), .S(n3450), .CO(n3451));
Q_AD01HF U4098 ( .A0(uClkCntr[13]), .B0(n3451), .S(n3452), .CO(n3453));
Q_AD01HF U4099 ( .A0(uClkCntr[14]), .B0(n3453), .S(n3454), .CO(n3455));
Q_AD01HF U4100 ( .A0(uClkCntr[15]), .B0(n3455), .S(n3456), .CO(n3457));
Q_AD01HF U4101 ( .A0(uClkCntr[16]), .B0(n3457), .S(n3458), .CO(n3459));
Q_AD01HF U4102 ( .A0(uClkCntr[17]), .B0(n3459), .S(n3460), .CO(n3461));
Q_AD01HF U4103 ( .A0(uClkCntr[18]), .B0(n3461), .S(n3462), .CO(n3463));
Q_AD01HF U4104 ( .A0(uClkCntr[19]), .B0(n3463), .S(n3464), .CO(n3465));
Q_AD01HF U4105 ( .A0(uClkCntr[20]), .B0(n3465), .S(n3466), .CO(n3467));
Q_AD01HF U4106 ( .A0(uClkCntr[21]), .B0(n3467), .S(n3468), .CO(n3469));
Q_AD01HF U4107 ( .A0(uClkCntr[22]), .B0(n3469), .S(n3470), .CO(n3471));
Q_AD01HF U4108 ( .A0(uClkCntr[23]), .B0(n3471), .S(n3472), .CO(n3473));
Q_AD01HF U4109 ( .A0(uClkCntr[24]), .B0(n3473), .S(n3474), .CO(n3475));
Q_AD01HF U4110 ( .A0(uClkCntr[25]), .B0(n3475), .S(n3476), .CO(n3477));
Q_AD01HF U4111 ( .A0(uClkCntr[26]), .B0(n3477), .S(n3478), .CO(n3479));
Q_AD01HF U4112 ( .A0(uClkCntr[27]), .B0(n3479), .S(n3480), .CO(n3481));
Q_AD01HF U4113 ( .A0(uClkCntr[28]), .B0(n3481), .S(n3482), .CO(n3483));
Q_AD01HF U4114 ( .A0(uClkCntr[29]), .B0(n3483), .S(n3484), .CO(n3485));
Q_AD01HF U4115 ( .A0(uClkCntr[30]), .B0(n3485), .S(n3486), .CO(n3487));
Q_AD01HF U4116 ( .A0(uClkCntr[31]), .B0(n3487), .S(n3488), .CO(n3489));
Q_AD01HF U4117 ( .A0(uClkCntr[32]), .B0(n3489), .S(n3490), .CO(n3491));
Q_AD01HF U4118 ( .A0(uClkCntr[33]), .B0(n3491), .S(n3492), .CO(n3493));
Q_AD01HF U4119 ( .A0(uClkCntr[34]), .B0(n3493), .S(n3494), .CO(n3495));
Q_AD01HF U4120 ( .A0(uClkCntr[35]), .B0(n3495), .S(n3496), .CO(n3497));
Q_AD01HF U4121 ( .A0(uClkCntr[36]), .B0(n3497), .S(n3498), .CO(n3499));
Q_AD01HF U4122 ( .A0(uClkCntr[37]), .B0(n3499), .S(n3500), .CO(n3501));
Q_AD01HF U4123 ( .A0(uClkCntr[38]), .B0(n3501), .S(n3502), .CO(n3503));
Q_AD01HF U4124 ( .A0(uClkCntr[39]), .B0(n3503), .S(n3504), .CO(n3505));
Q_AD01HF U4125 ( .A0(uClkCntr[40]), .B0(n3505), .S(n3506), .CO(n3507));
Q_AD01HF U4126 ( .A0(uClkCntr[41]), .B0(n3507), .S(n3508), .CO(n3509));
Q_AD01HF U4127 ( .A0(uClkCntr[42]), .B0(n3509), .S(n3510), .CO(n3511));
Q_AD01HF U4128 ( .A0(uClkCntr[43]), .B0(n3511), .S(n3512), .CO(n3513));
Q_AD01HF U4129 ( .A0(uClkCntr[44]), .B0(n3513), .S(n3514), .CO(n3515));
Q_AD01HF U4130 ( .A0(uClkCntr[45]), .B0(n3515), .S(n3516), .CO(n3517));
Q_AD01HF U4131 ( .A0(uClkCntr[46]), .B0(n3517), .S(n3518), .CO(n3519));
Q_AD01HF U4132 ( .A0(uClkCntr[47]), .B0(n3519), .S(n3520), .CO(n3521));
Q_AD01HF U4133 ( .A0(uClkCntr[48]), .B0(n3521), .S(n3522), .CO(n3523));
Q_AD01HF U4134 ( .A0(uClkCntr[49]), .B0(n3523), .S(n3524), .CO(n3525));
Q_AD01HF U4135 ( .A0(uClkCntr[50]), .B0(n3525), .S(n3526), .CO(n3527));
Q_AD01HF U4136 ( .A0(uClkCntr[51]), .B0(n3527), .S(n3528), .CO(n3529));
Q_AD01HF U4137 ( .A0(uClkCntr[52]), .B0(n3529), .S(n3530), .CO(n3531));
Q_AD01HF U4138 ( .A0(uClkCntr[53]), .B0(n3531), .S(n3532), .CO(n3533));
Q_AD01HF U4139 ( .A0(uClkCntr[54]), .B0(n3533), .S(n3534), .CO(n3535));
Q_AD01HF U4140 ( .A0(uClkCntr[55]), .B0(n3535), .S(n3536), .CO(n3537));
Q_AD01HF U4141 ( .A0(uClkCntr[56]), .B0(n3537), .S(n3538), .CO(n3539));
Q_AD01HF U4142 ( .A0(uClkCntr[57]), .B0(n3539), .S(n3540), .CO(n3541));
Q_AD01HF U4143 ( .A0(uClkCntr[58]), .B0(n3541), .S(n3542), .CO(n3543));
Q_AD01HF U4144 ( .A0(uClkCntr[59]), .B0(n3543), .S(n3544), .CO(n3545));
Q_AD01HF U4145 ( .A0(uClkCntr[60]), .B0(n3545), .S(n3546), .CO(n3547));
Q_AD01HF U4146 ( .A0(uClkCntr[61]), .B0(n3547), .S(n3548), .CO(n3549));
Q_AD01HF U4147 ( .A0(uClkCntr[62]), .B0(n3549), .S(n3550), .CO(n3551));
Q_FDP0 \nextDutTimeP_REG[63] ( .CK(mcp), .D(ixc_time.nextDutTime[63]), .Q(nextDutTimeP[63]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[62] ( .CK(mcp), .D(ixc_time.nextDutTime[62]), .Q(nextDutTimeP[62]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[61] ( .CK(mcp), .D(ixc_time.nextDutTime[61]), .Q(nextDutTimeP[61]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[60] ( .CK(mcp), .D(ixc_time.nextDutTime[60]), .Q(nextDutTimeP[60]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[59] ( .CK(mcp), .D(ixc_time.nextDutTime[59]), .Q(nextDutTimeP[59]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[58] ( .CK(mcp), .D(ixc_time.nextDutTime[58]), .Q(nextDutTimeP[58]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[57] ( .CK(mcp), .D(ixc_time.nextDutTime[57]), .Q(nextDutTimeP[57]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[56] ( .CK(mcp), .D(ixc_time.nextDutTime[56]), .Q(nextDutTimeP[56]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[55] ( .CK(mcp), .D(ixc_time.nextDutTime[55]), .Q(nextDutTimeP[55]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[54] ( .CK(mcp), .D(ixc_time.nextDutTime[54]), .Q(nextDutTimeP[54]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[53] ( .CK(mcp), .D(ixc_time.nextDutTime[53]), .Q(nextDutTimeP[53]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[52] ( .CK(mcp), .D(ixc_time.nextDutTime[52]), .Q(nextDutTimeP[52]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[51] ( .CK(mcp), .D(ixc_time.nextDutTime[51]), .Q(nextDutTimeP[51]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[50] ( .CK(mcp), .D(ixc_time.nextDutTime[50]), .Q(nextDutTimeP[50]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[49] ( .CK(mcp), .D(ixc_time.nextDutTime[49]), .Q(nextDutTimeP[49]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[48] ( .CK(mcp), .D(ixc_time.nextDutTime[48]), .Q(nextDutTimeP[48]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[47] ( .CK(mcp), .D(ixc_time.nextDutTime[47]), .Q(nextDutTimeP[47]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[46] ( .CK(mcp), .D(ixc_time.nextDutTime[46]), .Q(nextDutTimeP[46]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[45] ( .CK(mcp), .D(ixc_time.nextDutTime[45]), .Q(nextDutTimeP[45]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[44] ( .CK(mcp), .D(ixc_time.nextDutTime[44]), .Q(nextDutTimeP[44]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[43] ( .CK(mcp), .D(ixc_time.nextDutTime[43]), .Q(nextDutTimeP[43]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[42] ( .CK(mcp), .D(ixc_time.nextDutTime[42]), .Q(nextDutTimeP[42]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[41] ( .CK(mcp), .D(ixc_time.nextDutTime[41]), .Q(nextDutTimeP[41]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[40] ( .CK(mcp), .D(ixc_time.nextDutTime[40]), .Q(nextDutTimeP[40]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[39] ( .CK(mcp), .D(ixc_time.nextDutTime[39]), .Q(nextDutTimeP[39]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[38] ( .CK(mcp), .D(ixc_time.nextDutTime[38]), .Q(nextDutTimeP[38]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[37] ( .CK(mcp), .D(ixc_time.nextDutTime[37]), .Q(nextDutTimeP[37]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[36] ( .CK(mcp), .D(ixc_time.nextDutTime[36]), .Q(nextDutTimeP[36]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[35] ( .CK(mcp), .D(ixc_time.nextDutTime[35]), .Q(nextDutTimeP[35]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[34] ( .CK(mcp), .D(ixc_time.nextDutTime[34]), .Q(nextDutTimeP[34]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[33] ( .CK(mcp), .D(ixc_time.nextDutTime[33]), .Q(nextDutTimeP[33]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[32] ( .CK(mcp), .D(ixc_time.nextDutTime[32]), .Q(nextDutTimeP[32]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[31] ( .CK(mcp), .D(ixc_time.nextDutTime[31]), .Q(nextDutTimeP[31]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[30] ( .CK(mcp), .D(ixc_time.nextDutTime[30]), .Q(nextDutTimeP[30]), .QN(n3997));
Q_FDP0 \nextDutTimeP_REG[29] ( .CK(mcp), .D(ixc_time.nextDutTime[29]), .Q(nextDutTimeP[29]), .QN(n3998));
Q_FDP0 \nextDutTimeP_REG[28] ( .CK(mcp), .D(ixc_time.nextDutTime[28]), .Q(nextDutTimeP[28]), .QN(n3999));
Q_FDP0 \nextDutTimeP_REG[27] ( .CK(mcp), .D(ixc_time.nextDutTime[27]), .Q(nextDutTimeP[27]), .QN(n4000));
Q_FDP0 \nextDutTimeP_REG[26] ( .CK(mcp), .D(ixc_time.nextDutTime[26]), .Q(nextDutTimeP[26]), .QN(n4001));
Q_FDP0 \nextDutTimeP_REG[25] ( .CK(mcp), .D(ixc_time.nextDutTime[25]), .Q(nextDutTimeP[25]), .QN(n4002));
Q_FDP0 \nextDutTimeP_REG[24] ( .CK(mcp), .D(ixc_time.nextDutTime[24]), .Q(nextDutTimeP[24]), .QN(n4003));
Q_FDP0 \nextDutTimeP_REG[23] ( .CK(mcp), .D(ixc_time.nextDutTime[23]), .Q(nextDutTimeP[23]), .QN(n4004));
Q_FDP0 \nextDutTimeP_REG[22] ( .CK(mcp), .D(ixc_time.nextDutTime[22]), .Q(nextDutTimeP[22]), .QN(n4005));
Q_FDP0 \nextDutTimeP_REG[21] ( .CK(mcp), .D(ixc_time.nextDutTime[21]), .Q(nextDutTimeP[21]), .QN(n4006));
Q_FDP0 \nextDutTimeP_REG[20] ( .CK(mcp), .D(ixc_time.nextDutTime[20]), .Q(nextDutTimeP[20]), .QN(n4007));
Q_FDP0 \nextDutTimeP_REG[19] ( .CK(mcp), .D(ixc_time.nextDutTime[19]), .Q(nextDutTimeP[19]), .QN(n4008));
Q_FDP0 \nextDutTimeP_REG[18] ( .CK(mcp), .D(ixc_time.nextDutTime[18]), .Q(nextDutTimeP[18]), .QN(n4009));
Q_FDP0 \nextDutTimeP_REG[17] ( .CK(mcp), .D(ixc_time.nextDutTime[17]), .Q(nextDutTimeP[17]), .QN(n4010));
Q_FDP0 \nextDutTimeP_REG[16] ( .CK(mcp), .D(ixc_time.nextDutTime[16]), .Q(nextDutTimeP[16]), .QN(n4011));
Q_FDP0 \nextDutTimeP_REG[15] ( .CK(mcp), .D(ixc_time.nextDutTime[15]), .Q(nextDutTimeP[15]), .QN(n4012));
Q_FDP0 \nextDutTimeP_REG[14] ( .CK(mcp), .D(ixc_time.nextDutTime[14]), .Q(nextDutTimeP[14]), .QN(n4013));
Q_FDP0 \nextDutTimeP_REG[13] ( .CK(mcp), .D(ixc_time.nextDutTime[13]), .Q(nextDutTimeP[13]), .QN(n4014));
Q_FDP0 \nextDutTimeP_REG[12] ( .CK(mcp), .D(ixc_time.nextDutTime[12]), .Q(nextDutTimeP[12]), .QN(n4015));
Q_FDP0 \nextDutTimeP_REG[11] ( .CK(mcp), .D(ixc_time.nextDutTime[11]), .Q(nextDutTimeP[11]), .QN(n4016));
Q_FDP0 \nextDutTimeP_REG[10] ( .CK(mcp), .D(ixc_time.nextDutTime[10]), .Q(nextDutTimeP[10]), .QN(n4017));
Q_FDP0 \nextDutTimeP_REG[9] ( .CK(mcp), .D(ixc_time.nextDutTime[9]), .Q(nextDutTimeP[9]), .QN(n4018));
Q_FDP0 \nextDutTimeP_REG[8] ( .CK(mcp), .D(ixc_time.nextDutTime[8]), .Q(nextDutTimeP[8]), .QN(n4019));
Q_FDP0 \nextDutTimeP_REG[7] ( .CK(mcp), .D(ixc_time.nextDutTime[7]), .Q(nextDutTimeP[7]), .QN(n4020));
Q_FDP0 \nextDutTimeP_REG[6] ( .CK(mcp), .D(ixc_time.nextDutTime[6]), .Q(nextDutTimeP[6]), .QN(n4021));
Q_FDP0 \nextDutTimeP_REG[5] ( .CK(mcp), .D(ixc_time.nextDutTime[5]), .Q(nextDutTimeP[5]), .QN(n4022));
Q_FDP0 \nextDutTimeP_REG[4] ( .CK(mcp), .D(ixc_time.nextDutTime[4]), .Q(nextDutTimeP[4]), .QN(n4023));
Q_FDP0 \nextDutTimeP_REG[3] ( .CK(mcp), .D(ixc_time.nextDutTime[3]), .Q(nextDutTimeP[3]), .QN(n4024));
Q_FDP0 \nextDutTimeP_REG[2] ( .CK(mcp), .D(ixc_time.nextDutTime[2]), .Q(nextDutTimeP[2]), .QN(n4025));
Q_FDP0 \nextDutTimeP_REG[1] ( .CK(mcp), .D(ixc_time.nextDutTime[1]), .Q(nextDutTimeP[1]), .QN(n4026));
Q_FDP0 \nextDutTimeP_REG[0] ( .CK(mcp), .D(ixc_time.nextDutTime[0]), .Q(nextDutTimeP[0]), .QN(n4027));
Q_BUFZP U4212 ( .OE(syncEn), .A(n3552), .Z(stop1));
Q_OA21 U4213 ( .A0(hwClkDbgEn), .A1(cakeUcEnable), .B0(hwClkDbg), .Z(hwClkDbgOn));
Q_OR02 U4214 ( .A0(callEmuPre), .A1(it_newBuf), .Z(n3553));
Q_LDP0 it_newBufPO_REG  ( .G(n3553), .D(it_newBuf), .Q(it_newBufPO), .QN( ));
Q_INV U4216 ( .A(callEmuEv), .Z(n3555));
Q_NR02 U4217 ( .A0(callEmuEv), .A1(hasGFIFO1), .Z(n3557));
Q_NR02 U4218 ( .A0(hasGFIFO2), .A1(hasSFIFO), .Z(n3558));
Q_INV U4219 ( .A(hasPTX), .Z(n3556));
Q_AN03 U4220 ( .A0(n3557), .A1(n3556), .A2(n3558), .Z(n3554));
Q_NR02 U4221 ( .A0(n3554), .A1(callEmuEv), .Z(n3559));
Q_MX02 U4222 ( .S(n3554), .A0(n3559), .A1(mioPOW_2[1]), .Z(intr));
Q_AD01HF U4223 ( .A0(bpCount[1]), .B0(bpCount[0]), .S(n3561), .CO(n3562));
Q_AD01HF U4224 ( .A0(bpCount[2]), .B0(n3562), .S(n3563), .CO(n3564));
Q_AD01HF U4225 ( .A0(bpCount[3]), .B0(n3564), .S(n3565), .CO(n3566));
Q_AD01HF U4226 ( .A0(bpCount[4]), .B0(n3566), .S(n3567), .CO(n3568));
Q_AD01HF U4227 ( .A0(bpCount[5]), .B0(n3568), .S(n3569), .CO(n3570));
Q_AD01HF U4228 ( .A0(bpCount[6]), .B0(n3570), .S(n3571), .CO(n3572));
Q_AD01HF U4229 ( .A0(bpCount[7]), .B0(n3572), .S(n3573), .CO(n3574));
Q_AD01HF U4230 ( .A0(bpCount[8]), .B0(n3574), .S(n3575), .CO(n3576));
Q_AD01HF U4231 ( .A0(bpCount[9]), .B0(n3576), .S(n3577), .CO(n3578));
Q_AD01HF U4232 ( .A0(bpCount[10]), .B0(n3578), .S(n3579), .CO(n3580));
Q_AD01HF U4233 ( .A0(bpCount[11]), .B0(n3580), .S(n3581), .CO(n3582));
Q_AD01HF U4234 ( .A0(bpCount[12]), .B0(n3582), .S(n3583), .CO(n3584));
Q_AD01HF U4235 ( .A0(bpCount[13]), .B0(n3584), .S(n3585), .CO(n3586));
Q_AD01HF U4236 ( .A0(bpCount[14]), .B0(n3586), .S(n3587), .CO(n3588));
Q_AD01HF U4237 ( .A0(bpCount[15]), .B0(n3588), .S(n3589), .CO(n3590));
Q_AD01HF U4238 ( .A0(bpCount[16]), .B0(n3590), .S(n3591), .CO(n3592));
Q_AD01HF U4239 ( .A0(bpCount[17]), .B0(n3592), .S(n3593), .CO(n3594));
Q_AD01HF U4240 ( .A0(bpCount[18]), .B0(n3594), .S(n3595), .CO(n3596));
Q_AD01HF U4241 ( .A0(bpCount[19]), .B0(n3596), .S(n3597), .CO(n3598));
Q_AD01HF U4242 ( .A0(bpCount[20]), .B0(n3598), .S(n3599), .CO(n3600));
Q_AD01HF U4243 ( .A0(bpCount[21]), .B0(n3600), .S(n3601), .CO(n3602));
Q_AD01HF U4244 ( .A0(bpCount[22]), .B0(n3602), .S(n3603), .CO(n3604));
Q_AD01HF U4245 ( .A0(bpCount[23]), .B0(n3604), .S(n3605), .CO(n3606));
Q_AD01HF U4246 ( .A0(bpCount[24]), .B0(n3606), .S(n3607), .CO(n3608));
Q_AD01HF U4247 ( .A0(bpCount[25]), .B0(n3608), .S(n3609), .CO(n3610));
Q_AD01HF U4248 ( .A0(bpCount[26]), .B0(n3610), .S(n3611), .CO(n3612));
Q_AD01HF U4249 ( .A0(bpCount[27]), .B0(n3612), .S(n3613), .CO(n3614));
Q_AD01HF U4250 ( .A0(bpCount[28]), .B0(n3614), .S(n3615), .CO(n3616));
Q_AD01HF U4251 ( .A0(bpCount[29]), .B0(n3616), .S(n3617), .CO(n3618));
Q_AD01HF U4252 ( .A0(bpCount[30]), .B0(n3618), .S(n3619), .CO(n3620));
Q_AD01HF U4253 ( .A0(bpCount[31]), .B0(n3620), .S(n3621), .CO(n3622));
Q_AD01HF U4254 ( .A0(bpCount[32]), .B0(n3622), .S(n3623), .CO(n3624));
Q_AD01HF U4255 ( .A0(bpCount[33]), .B0(n3624), .S(n3625), .CO(n3626));
Q_AD01HF U4256 ( .A0(bpCount[34]), .B0(n3626), .S(n3627), .CO(n3628));
Q_AD01HF U4257 ( .A0(bpCount[35]), .B0(n3628), .S(n3629), .CO(n3630));
Q_AD01HF U4258 ( .A0(bpCount[36]), .B0(n3630), .S(n3631), .CO(n3632));
Q_AD01HF U4259 ( .A0(bpCount[37]), .B0(n3632), .S(n3633), .CO(n3634));
Q_AD01HF U4260 ( .A0(bpCount[38]), .B0(n3634), .S(n3635), .CO(n3636));
Q_AD01HF U4261 ( .A0(bpCount[39]), .B0(n3636), .S(n3637), .CO(n3638));
Q_AD01HF U4262 ( .A0(bpCount[40]), .B0(n3638), .S(n3639), .CO(n3640));
Q_AD01HF U4263 ( .A0(bpCount[41]), .B0(n3640), .S(n3641), .CO(n3642));
Q_AD01HF U4264 ( .A0(bpCount[42]), .B0(n3642), .S(n3643), .CO(n3644));
Q_AD01HF U4265 ( .A0(bpCount[43]), .B0(n3644), .S(n3645), .CO(n3646));
Q_AD01HF U4266 ( .A0(bpCount[44]), .B0(n3646), .S(n3647), .CO(n3648));
Q_AD01HF U4267 ( .A0(bpCount[45]), .B0(n3648), .S(n3649), .CO(n3650));
Q_AD01HF U4268 ( .A0(bpCount[46]), .B0(n3650), .S(n3651), .CO(n3652));
Q_AD01HF U4269 ( .A0(bpCount[47]), .B0(n3652), .S(n3653), .CO(n3654));
Q_AD01HF U4270 ( .A0(bpCount[48]), .B0(n3654), .S(n3655), .CO(n3656));
Q_AD01HF U4271 ( .A0(bpCount[49]), .B0(n3656), .S(n3657), .CO(n3658));
Q_AD01HF U4272 ( .A0(bpCount[50]), .B0(n3658), .S(n3659), .CO(n3660));
Q_AD01HF U4273 ( .A0(bpCount[51]), .B0(n3660), .S(n3661), .CO(n3662));
Q_AD01HF U4274 ( .A0(bpCount[52]), .B0(n3662), .S(n3663), .CO(n3664));
Q_AD01HF U4275 ( .A0(bpCount[53]), .B0(n3664), .S(n3665), .CO(n3666));
Q_AD01HF U4276 ( .A0(bpCount[54]), .B0(n3666), .S(n3667), .CO(n3668));
Q_AD01HF U4277 ( .A0(bpCount[55]), .B0(n3668), .S(n3669), .CO(n3670));
Q_AD01HF U4278 ( .A0(bpCount[56]), .B0(n3670), .S(n3671), .CO(n3672));
Q_AD01HF U4279 ( .A0(bpCount[57]), .B0(n3672), .S(n3673), .CO(n3674));
Q_AD01HF U4280 ( .A0(bpCount[58]), .B0(n3674), .S(n3675), .CO(n3676));
Q_AD01HF U4281 ( .A0(bpCount[59]), .B0(n3676), .S(n3677), .CO(n3678));
Q_AD01HF U4282 ( .A0(bpCount[60]), .B0(n3678), .S(n3679), .CO(n3680));
Q_AD01HF U4283 ( .A0(bpCount[61]), .B0(n3680), .S(n3681), .CO(n3682));
Q_AD01HF U4284 ( .A0(bpCount[62]), .B0(n3682), .S(n3683), .CO(n3684));
Q_FDP0 \bpCount_REG[62] ( .CK(bClk), .D(n3683), .Q(bpCount[62]), .QN( ));
Q_FDP0 \bpCount_REG[61] ( .CK(bClk), .D(n3681), .Q(bpCount[61]), .QN( ));
Q_FDP0 \bpCount_REG[60] ( .CK(bClk), .D(n3679), .Q(bpCount[60]), .QN( ));
Q_FDP0 \bpCount_REG[59] ( .CK(bClk), .D(n3677), .Q(bpCount[59]), .QN( ));
Q_FDP0 \bpCount_REG[58] ( .CK(bClk), .D(n3675), .Q(bpCount[58]), .QN( ));
Q_FDP0 \bpCount_REG[57] ( .CK(bClk), .D(n3673), .Q(bpCount[57]), .QN( ));
Q_FDP0 \bpCount_REG[56] ( .CK(bClk), .D(n3671), .Q(bpCount[56]), .QN( ));
Q_FDP0 \bpCount_REG[55] ( .CK(bClk), .D(n3669), .Q(bpCount[55]), .QN( ));
Q_FDP0 \bpCount_REG[54] ( .CK(bClk), .D(n3667), .Q(bpCount[54]), .QN( ));
Q_FDP0 \bpCount_REG[53] ( .CK(bClk), .D(n3665), .Q(bpCount[53]), .QN( ));
Q_FDP0 \bpCount_REG[52] ( .CK(bClk), .D(n3663), .Q(bpCount[52]), .QN( ));
Q_FDP0 \bpCount_REG[51] ( .CK(bClk), .D(n3661), .Q(bpCount[51]), .QN( ));
Q_FDP0 \bpCount_REG[50] ( .CK(bClk), .D(n3659), .Q(bpCount[50]), .QN( ));
Q_FDP0 \bpCount_REG[49] ( .CK(bClk), .D(n3657), .Q(bpCount[49]), .QN( ));
Q_FDP0 \bpCount_REG[48] ( .CK(bClk), .D(n3655), .Q(bpCount[48]), .QN( ));
Q_FDP0 \bpCount_REG[47] ( .CK(bClk), .D(n3653), .Q(bpCount[47]), .QN( ));
Q_FDP0 \bpCount_REG[46] ( .CK(bClk), .D(n3651), .Q(bpCount[46]), .QN( ));
Q_FDP0 \bpCount_REG[45] ( .CK(bClk), .D(n3649), .Q(bpCount[45]), .QN( ));
Q_FDP0 \bpCount_REG[44] ( .CK(bClk), .D(n3647), .Q(bpCount[44]), .QN( ));
Q_FDP0 \bpCount_REG[43] ( .CK(bClk), .D(n3645), .Q(bpCount[43]), .QN( ));
Q_FDP0 \bpCount_REG[42] ( .CK(bClk), .D(n3643), .Q(bpCount[42]), .QN( ));
Q_FDP0 \bpCount_REG[41] ( .CK(bClk), .D(n3641), .Q(bpCount[41]), .QN( ));
Q_FDP0 \bpCount_REG[40] ( .CK(bClk), .D(n3639), .Q(bpCount[40]), .QN( ));
Q_FDP0 \bpCount_REG[39] ( .CK(bClk), .D(n3637), .Q(bpCount[39]), .QN( ));
Q_FDP0 \bpCount_REG[38] ( .CK(bClk), .D(n3635), .Q(bpCount[38]), .QN( ));
Q_FDP0 \bpCount_REG[37] ( .CK(bClk), .D(n3633), .Q(bpCount[37]), .QN( ));
Q_FDP0 \bpCount_REG[36] ( .CK(bClk), .D(n3631), .Q(bpCount[36]), .QN( ));
Q_FDP0 \bpCount_REG[35] ( .CK(bClk), .D(n3629), .Q(bpCount[35]), .QN( ));
Q_FDP0 \bpCount_REG[34] ( .CK(bClk), .D(n3627), .Q(bpCount[34]), .QN( ));
Q_FDP0 \bpCount_REG[33] ( .CK(bClk), .D(n3625), .Q(bpCount[33]), .QN( ));
Q_FDP0 \bpCount_REG[32] ( .CK(bClk), .D(n3623), .Q(bpCount[32]), .QN( ));
Q_FDP0 \bpCount_REG[31] ( .CK(bClk), .D(n3621), .Q(bpCount[31]), .QN( ));
Q_FDP0 \bpCount_REG[30] ( .CK(bClk), .D(n3619), .Q(bpCount[30]), .QN( ));
Q_FDP0 \bpCount_REG[29] ( .CK(bClk), .D(n3617), .Q(bpCount[29]), .QN( ));
Q_FDP0 \bpCount_REG[28] ( .CK(bClk), .D(n3615), .Q(bpCount[28]), .QN( ));
Q_FDP0 \bpCount_REG[27] ( .CK(bClk), .D(n3613), .Q(bpCount[27]), .QN( ));
Q_FDP0 \bpCount_REG[26] ( .CK(bClk), .D(n3611), .Q(bpCount[26]), .QN( ));
Q_FDP0 \bpCount_REG[25] ( .CK(bClk), .D(n3609), .Q(bpCount[25]), .QN( ));
Q_FDP0 \bpCount_REG[24] ( .CK(bClk), .D(n3607), .Q(bpCount[24]), .QN( ));
Q_FDP0 \bpCount_REG[23] ( .CK(bClk), .D(n3605), .Q(bpCount[23]), .QN( ));
Q_FDP0 \bpCount_REG[22] ( .CK(bClk), .D(n3603), .Q(bpCount[22]), .QN( ));
Q_FDP0 \bpCount_REG[21] ( .CK(bClk), .D(n3601), .Q(bpCount[21]), .QN( ));
Q_FDP0 \bpCount_REG[20] ( .CK(bClk), .D(n3599), .Q(bpCount[20]), .QN( ));
Q_FDP0 \bpCount_REG[19] ( .CK(bClk), .D(n3597), .Q(bpCount[19]), .QN( ));
Q_FDP0 \bpCount_REG[18] ( .CK(bClk), .D(n3595), .Q(bpCount[18]), .QN( ));
Q_FDP0 \bpCount_REG[17] ( .CK(bClk), .D(n3593), .Q(bpCount[17]), .QN( ));
Q_FDP0 \bpCount_REG[16] ( .CK(bClk), .D(n3591), .Q(bpCount[16]), .QN( ));
Q_FDP0 \bpCount_REG[15] ( .CK(bClk), .D(n3589), .Q(bpCount[15]), .QN( ));
Q_FDP0 \bpCount_REG[14] ( .CK(bClk), .D(n3587), .Q(bpCount[14]), .QN( ));
Q_FDP0 \bpCount_REG[13] ( .CK(bClk), .D(n3585), .Q(bpCount[13]), .QN( ));
Q_FDP0 \bpCount_REG[12] ( .CK(bClk), .D(n3583), .Q(bpCount[12]), .QN( ));
Q_FDP0 \bpCount_REG[11] ( .CK(bClk), .D(n3581), .Q(bpCount[11]), .QN( ));
Q_FDP0 \bpCount_REG[10] ( .CK(bClk), .D(n3579), .Q(bpCount[10]), .QN( ));
Q_FDP0 \bpCount_REG[9] ( .CK(bClk), .D(n3577), .Q(bpCount[9]), .QN( ));
Q_FDP0 \bpCount_REG[8] ( .CK(bClk), .D(n3575), .Q(bpCount[8]), .QN( ));
Q_FDP0 \bpCount_REG[7] ( .CK(bClk), .D(n3573), .Q(bpCount[7]), .QN( ));
Q_FDP0 \bpCount_REG[6] ( .CK(bClk), .D(n3571), .Q(bpCount[6]), .QN( ));
Q_FDP0 \bpCount_REG[5] ( .CK(bClk), .D(n3569), .Q(bpCount[5]), .QN( ));
Q_FDP0 \bpCount_REG[4] ( .CK(bClk), .D(n3567), .Q(bpCount[4]), .QN( ));
Q_FDP0 \bpCount_REG[3] ( .CK(bClk), .D(n3565), .Q(bpCount[3]), .QN( ));
Q_FDP0 \bpCount_REG[2] ( .CK(bClk), .D(n3563), .Q(bpCount[2]), .QN( ));
Q_FDP0 \bpCount_REG[1] ( .CK(bClk), .D(n3561), .Q(bpCount[1]), .QN( ));
Q_FDP0 \bpCount_REG[0] ( .CK(bClk), .D(n3560), .Q(bpCount[0]), .QN(n3560));
Q_AD01HF U4348 ( .A0(eCount[1]), .B0(eCount[0]), .S(n3686), .CO(n3687));
Q_AD01HF U4349 ( .A0(eCount[2]), .B0(n3687), .S(n3688), .CO(n3689));
Q_AD01HF U4350 ( .A0(eCount[3]), .B0(n3689), .S(n3690), .CO(n3691));
Q_AD01HF U4351 ( .A0(eCount[4]), .B0(n3691), .S(n3692), .CO(n3693));
Q_AD01HF U4352 ( .A0(eCount[5]), .B0(n3693), .S(n3694), .CO(n3695));
Q_AD01HF U4353 ( .A0(eCount[6]), .B0(n3695), .S(n3696), .CO(n3697));
Q_AD01HF U4354 ( .A0(eCount[7]), .B0(n3697), .S(n3698), .CO(n3699));
Q_AD01HF U4355 ( .A0(eCount[8]), .B0(n3699), .S(n3700), .CO(n3701));
Q_AD01HF U4356 ( .A0(eCount[9]), .B0(n3701), .S(n3702), .CO(n3703));
Q_AD01HF U4357 ( .A0(eCount[10]), .B0(n3703), .S(n3704), .CO(n3705));
Q_AD01HF U4358 ( .A0(eCount[11]), .B0(n3705), .S(n3706), .CO(n3707));
Q_AD01HF U4359 ( .A0(eCount[12]), .B0(n3707), .S(n3708), .CO(n3709));
Q_AD01HF U4360 ( .A0(eCount[13]), .B0(n3709), .S(n3710), .CO(n3711));
Q_AD01HF U4361 ( .A0(eCount[14]), .B0(n3711), .S(n3712), .CO(n3713));
Q_AD01HF U4362 ( .A0(eCount[15]), .B0(n3713), .S(n3714), .CO(n3715));
Q_AD01HF U4363 ( .A0(eCount[16]), .B0(n3715), .S(n3716), .CO(n3717));
Q_AD01HF U4364 ( .A0(eCount[17]), .B0(n3717), .S(n3718), .CO(n3719));
Q_AD01HF U4365 ( .A0(eCount[18]), .B0(n3719), .S(n3720), .CO(n3721));
Q_AD01HF U4366 ( .A0(eCount[19]), .B0(n3721), .S(n3722), .CO(n3723));
Q_AD01HF U4367 ( .A0(eCount[20]), .B0(n3723), .S(n3724), .CO(n3725));
Q_AD01HF U4368 ( .A0(eCount[21]), .B0(n3725), .S(n3726), .CO(n3727));
Q_AD01HF U4369 ( .A0(eCount[22]), .B0(n3727), .S(n3728), .CO(n3729));
Q_AD01HF U4370 ( .A0(eCount[23]), .B0(n3729), .S(n3730), .CO(n3731));
Q_AD01HF U4371 ( .A0(eCount[24]), .B0(n3731), .S(n3732), .CO(n3733));
Q_AD01HF U4372 ( .A0(eCount[25]), .B0(n3733), .S(n3734), .CO(n3735));
Q_AD01HF U4373 ( .A0(eCount[26]), .B0(n3735), .S(n3736), .CO(n3737));
Q_AD01HF U4374 ( .A0(eCount[27]), .B0(n3737), .S(n3738), .CO(n3739));
Q_AD01HF U4375 ( .A0(eCount[28]), .B0(n3739), .S(n3740), .CO(n3741));
Q_AD01HF U4376 ( .A0(eCount[29]), .B0(n3741), .S(n3742), .CO(n3743));
Q_AD01HF U4377 ( .A0(eCount[30]), .B0(n3743), .S(n3744), .CO(n3745));
Q_AD01HF U4378 ( .A0(eCount[31]), .B0(n3745), .S(n3746), .CO(n3747));
Q_AD01HF U4379 ( .A0(eCount[32]), .B0(n3747), .S(n3748), .CO(n3749));
Q_AD01HF U4380 ( .A0(eCount[33]), .B0(n3749), .S(n3750), .CO(n3751));
Q_AD01HF U4381 ( .A0(eCount[34]), .B0(n3751), .S(n3752), .CO(n3753));
Q_AD01HF U4382 ( .A0(eCount[35]), .B0(n3753), .S(n3754), .CO(n3755));
Q_AD01HF U4383 ( .A0(eCount[36]), .B0(n3755), .S(n3756), .CO(n3757));
Q_AD01HF U4384 ( .A0(eCount[37]), .B0(n3757), .S(n3758), .CO(n3759));
Q_AD01HF U4385 ( .A0(eCount[38]), .B0(n3759), .S(n3760), .CO(n3761));
Q_AD01HF U4386 ( .A0(eCount[39]), .B0(n3761), .S(n3762), .CO(n3763));
Q_AD01HF U4387 ( .A0(eCount[40]), .B0(n3763), .S(n3764), .CO(n3765));
Q_AD01HF U4388 ( .A0(eCount[41]), .B0(n3765), .S(n3766), .CO(n3767));
Q_AD01HF U4389 ( .A0(eCount[42]), .B0(n3767), .S(n3768), .CO(n3769));
Q_AD01HF U4390 ( .A0(eCount[43]), .B0(n3769), .S(n3770), .CO(n3771));
Q_AD01HF U4391 ( .A0(eCount[44]), .B0(n3771), .S(n3772), .CO(n3773));
Q_AD01HF U4392 ( .A0(eCount[45]), .B0(n3773), .S(n3774), .CO(n3775));
Q_AD01HF U4393 ( .A0(eCount[46]), .B0(n3775), .S(n3776), .CO(n3777));
Q_AD01HF U4394 ( .A0(eCount[47]), .B0(n3777), .S(n3778), .CO(n3779));
Q_AD01HF U4395 ( .A0(eCount[48]), .B0(n3779), .S(n3780), .CO(n3781));
Q_AD01HF U4396 ( .A0(eCount[49]), .B0(n3781), .S(n3782), .CO(n3783));
Q_AD01HF U4397 ( .A0(eCount[50]), .B0(n3783), .S(n3784), .CO(n3785));
Q_AD01HF U4398 ( .A0(eCount[51]), .B0(n3785), .S(n3786), .CO(n3787));
Q_AD01HF U4399 ( .A0(eCount[52]), .B0(n3787), .S(n3788), .CO(n3789));
Q_AD01HF U4400 ( .A0(eCount[53]), .B0(n3789), .S(n3790), .CO(n3791));
Q_AD01HF U4401 ( .A0(eCount[54]), .B0(n3791), .S(n3792), .CO(n3793));
Q_AD01HF U4402 ( .A0(eCount[55]), .B0(n3793), .S(n3794), .CO(n3795));
Q_AD01HF U4403 ( .A0(eCount[56]), .B0(n3795), .S(n3796), .CO(n3797));
Q_AD01HF U4404 ( .A0(eCount[57]), .B0(n3797), .S(n3798), .CO(n3799));
Q_AD01HF U4405 ( .A0(eCount[58]), .B0(n3799), .S(n3800), .CO(n3801));
Q_AD01HF U4406 ( .A0(eCount[59]), .B0(n3801), .S(n3802), .CO(n3803));
Q_AD01HF U4407 ( .A0(eCount[60]), .B0(n3803), .S(n3804), .CO(n3805));
Q_AD01HF U4408 ( .A0(eCount[61]), .B0(n3805), .S(n3806), .CO(n3807));
Q_AD01HF U4409 ( .A0(eCount[62]), .B0(n3807), .S(n3808), .CO(n3809));
Q_FDP0 \eCount_REG[62] ( .CK(eClk), .D(n3808), .Q(eCount[62]), .QN( ));
Q_FDP0 \eCount_REG[61] ( .CK(eClk), .D(n3806), .Q(eCount[61]), .QN( ));
Q_FDP0 \eCount_REG[60] ( .CK(eClk), .D(n3804), .Q(eCount[60]), .QN( ));
Q_FDP0 \eCount_REG[59] ( .CK(eClk), .D(n3802), .Q(eCount[59]), .QN( ));
Q_FDP0 \eCount_REG[58] ( .CK(eClk), .D(n3800), .Q(eCount[58]), .QN( ));
Q_FDP0 \eCount_REG[57] ( .CK(eClk), .D(n3798), .Q(eCount[57]), .QN( ));
Q_FDP0 \eCount_REG[56] ( .CK(eClk), .D(n3796), .Q(eCount[56]), .QN( ));
Q_FDP0 \eCount_REG[55] ( .CK(eClk), .D(n3794), .Q(eCount[55]), .QN( ));
Q_FDP0 \eCount_REG[54] ( .CK(eClk), .D(n3792), .Q(eCount[54]), .QN( ));
Q_FDP0 \eCount_REG[53] ( .CK(eClk), .D(n3790), .Q(eCount[53]), .QN( ));
Q_FDP0 \eCount_REG[52] ( .CK(eClk), .D(n3788), .Q(eCount[52]), .QN( ));
Q_FDP0 \eCount_REG[51] ( .CK(eClk), .D(n3786), .Q(eCount[51]), .QN( ));
Q_FDP0 \eCount_REG[50] ( .CK(eClk), .D(n3784), .Q(eCount[50]), .QN( ));
Q_FDP0 \eCount_REG[49] ( .CK(eClk), .D(n3782), .Q(eCount[49]), .QN( ));
Q_FDP0 \eCount_REG[48] ( .CK(eClk), .D(n3780), .Q(eCount[48]), .QN( ));
Q_FDP0 \eCount_REG[47] ( .CK(eClk), .D(n3778), .Q(eCount[47]), .QN( ));
Q_FDP0 \eCount_REG[46] ( .CK(eClk), .D(n3776), .Q(eCount[46]), .QN( ));
Q_FDP0 \eCount_REG[45] ( .CK(eClk), .D(n3774), .Q(eCount[45]), .QN( ));
Q_FDP0 \eCount_REG[44] ( .CK(eClk), .D(n3772), .Q(eCount[44]), .QN( ));
Q_FDP0 \eCount_REG[43] ( .CK(eClk), .D(n3770), .Q(eCount[43]), .QN( ));
Q_FDP0 \eCount_REG[42] ( .CK(eClk), .D(n3768), .Q(eCount[42]), .QN( ));
Q_FDP0 \eCount_REG[41] ( .CK(eClk), .D(n3766), .Q(eCount[41]), .QN( ));
Q_FDP0 \eCount_REG[40] ( .CK(eClk), .D(n3764), .Q(eCount[40]), .QN( ));
Q_FDP0 \eCount_REG[39] ( .CK(eClk), .D(n3762), .Q(eCount[39]), .QN( ));
Q_FDP0 \eCount_REG[38] ( .CK(eClk), .D(n3760), .Q(eCount[38]), .QN( ));
Q_FDP0 \eCount_REG[37] ( .CK(eClk), .D(n3758), .Q(eCount[37]), .QN( ));
Q_FDP0 \eCount_REG[36] ( .CK(eClk), .D(n3756), .Q(eCount[36]), .QN( ));
Q_FDP0 \eCount_REG[35] ( .CK(eClk), .D(n3754), .Q(eCount[35]), .QN( ));
Q_FDP0 \eCount_REG[34] ( .CK(eClk), .D(n3752), .Q(eCount[34]), .QN( ));
Q_FDP0 \eCount_REG[33] ( .CK(eClk), .D(n3750), .Q(eCount[33]), .QN( ));
Q_FDP0 \eCount_REG[32] ( .CK(eClk), .D(n3748), .Q(eCount[32]), .QN( ));
Q_FDP0 \eCount_REG[31] ( .CK(eClk), .D(n3746), .Q(eCount[31]), .QN( ));
Q_FDP0 \eCount_REG[30] ( .CK(eClk), .D(n3744), .Q(eCount[30]), .QN( ));
Q_FDP0 \eCount_REG[29] ( .CK(eClk), .D(n3742), .Q(eCount[29]), .QN( ));
Q_FDP0 \eCount_REG[28] ( .CK(eClk), .D(n3740), .Q(eCount[28]), .QN( ));
Q_FDP0 \eCount_REG[27] ( .CK(eClk), .D(n3738), .Q(eCount[27]), .QN( ));
Q_FDP0 \eCount_REG[26] ( .CK(eClk), .D(n3736), .Q(eCount[26]), .QN( ));
Q_FDP0 \eCount_REG[25] ( .CK(eClk), .D(n3734), .Q(eCount[25]), .QN( ));
Q_FDP0 \eCount_REG[24] ( .CK(eClk), .D(n3732), .Q(eCount[24]), .QN( ));
Q_FDP0 \eCount_REG[23] ( .CK(eClk), .D(n3730), .Q(eCount[23]), .QN( ));
Q_FDP0 \eCount_REG[22] ( .CK(eClk), .D(n3728), .Q(eCount[22]), .QN( ));
Q_FDP0 \eCount_REG[21] ( .CK(eClk), .D(n3726), .Q(eCount[21]), .QN( ));
Q_FDP0 \eCount_REG[20] ( .CK(eClk), .D(n3724), .Q(eCount[20]), .QN( ));
Q_FDP0 \eCount_REG[19] ( .CK(eClk), .D(n3722), .Q(eCount[19]), .QN( ));
Q_FDP0 \eCount_REG[18] ( .CK(eClk), .D(n3720), .Q(eCount[18]), .QN( ));
Q_FDP0 \eCount_REG[17] ( .CK(eClk), .D(n3718), .Q(eCount[17]), .QN( ));
Q_FDP0 \eCount_REG[16] ( .CK(eClk), .D(n3716), .Q(eCount[16]), .QN( ));
Q_FDP0 \eCount_REG[15] ( .CK(eClk), .D(n3714), .Q(eCount[15]), .QN( ));
Q_FDP0 \eCount_REG[14] ( .CK(eClk), .D(n3712), .Q(eCount[14]), .QN( ));
Q_FDP0 \eCount_REG[13] ( .CK(eClk), .D(n3710), .Q(eCount[13]), .QN( ));
Q_FDP0 \eCount_REG[12] ( .CK(eClk), .D(n3708), .Q(eCount[12]), .QN( ));
Q_FDP0 \eCount_REG[11] ( .CK(eClk), .D(n3706), .Q(eCount[11]), .QN( ));
Q_FDP0 \eCount_REG[10] ( .CK(eClk), .D(n3704), .Q(eCount[10]), .QN( ));
Q_FDP0 \eCount_REG[9] ( .CK(eClk), .D(n3702), .Q(eCount[9]), .QN( ));
Q_FDP0 \eCount_REG[8] ( .CK(eClk), .D(n3700), .Q(eCount[8]), .QN( ));
Q_FDP0 \eCount_REG[7] ( .CK(eClk), .D(n3698), .Q(eCount[7]), .QN( ));
Q_FDP0 \eCount_REG[6] ( .CK(eClk), .D(n3696), .Q(eCount[6]), .QN( ));
Q_FDP0 \eCount_REG[5] ( .CK(eClk), .D(n3694), .Q(eCount[5]), .QN( ));
Q_FDP0 \eCount_REG[4] ( .CK(eClk), .D(n3692), .Q(eCount[4]), .QN( ));
Q_FDP0 \eCount_REG[3] ( .CK(eClk), .D(n3690), .Q(eCount[3]), .QN( ));
Q_FDP0 \eCount_REG[2] ( .CK(eClk), .D(n3688), .Q(eCount[2]), .QN( ));
Q_FDP0 \eCount_REG[1] ( .CK(eClk), .D(n3686), .Q(eCount[1]), .QN( ));
Q_FDP0 \eCount_REG[0] ( .CK(eClk), .D(n3685), .Q(eCount[0]), .QN(n3685));
Q_OA21 U4473 ( .A0(n2917), .A1(n2915), .B0(n2916), .Z(n3810));
Q_INV U4474 ( .A(n2916), .Z(n3811));
Q_MX02 U4475 ( .S(n3810), .A0(n3812), .A1(n3813), .Z(lastDelta));
Q_AN02 U4476 ( .A0(n3811), .A1(n2917), .Z(n3812));
Q_NR03 U4477 ( .A0(n2916), .A1(bpHalt), .A2(bClkHoldD), .Z(bpOn));
Q_OR02 U4478 ( .A0(hotSwapOnPI), .A1(n3814), .Z(n3813));
Q_NR02 U4479 ( .A0(n3001), .A1(eClkHold), .Z(n3814));
Q_AO21 U4480 ( .A0(callEmuEv), .A1(tbcPOState[0]), .B0(n3821), .Z(n3816));
Q_AO21 U4481 ( .A0(tbcPOd), .A1(tbcPORdy), .B0(tbcPOState[0]), .Z(n3820));
Q_OR02 U4482 ( .A0(tbcPOState[1]), .A1(n3816), .Z(n3823));
Q_INV U4483 ( .A(n3823), .Z(n3817));
Q_OR02 U4484 ( .A0(forceAbort), .A1(n3817), .Z(tbcPO));
Q_INV U4485 ( .A(tbcPOd), .Z(n3818));
Q_OR02 U4486 ( .A0(tbcPOState[0]), .A1(n3818), .Z(n3819));
Q_INV U4487 ( .A(n3820), .Z(n3821));
Q_MX02 U4488 ( .S(tbcPOState[1]), .A0(n3821), .A1(n3819), .Z(n3822));
Q_OR02 U4489 ( .A0(forceAbort), .A1(n3822), .Z(n3815));
Q_OR02 U4490 ( .A0(forceAbort), .A1(n3823), .Z(n3824));
Q_INV U4491 ( .A(n3824), .Z(tbcPOStateN[0]));
Q_XOR2 U4492 ( .A0(n3824), .A1(n3815), .Z(tbcPOStateN[1]));
Q_AN03 U4493 ( .A0(tbcPODly[4]), .A1(tbcPODly[3]), .A2(tbcPODly[2]), .Z(n3825));
Q_AN03 U4494 ( .A0(tbcPODly[1]), .A1(tbcPODly[0]), .A2(n3825), .Z(n3826));
Q_OR02 U4495 ( .A0(n3826), .A1(n3046), .Z(n3827));
Q_INV U4496 ( .A(gfifoWait), .Z(n3828));
Q_NR03 U4497 ( .A0(osfWait), .A1(asyncBusy), .A2(ptxBusy), .Z(n3829));
Q_AN03 U4498 ( .A0(n3828), .A1(n3829), .A2(n3827), .Z(tbcPORdy));
Q_NR02 U4499 ( .A0(callEmuPre), .A1(stop3), .Z(n3830));
Q_AN02 U4500 ( .A0(n1406), .A1(stop3), .Z(n3831));
Q_NR02 U4501 ( .A0(callEmuPre), .A1(stopT), .Z(n3832));
Q_AN02 U4502 ( .A0(n1406), .A1(stopT), .Z(n3833));
Q_MX02 U4503 ( .S(n3830), .A0(n3831), .A1(stop3POd), .Z(stop3PO));
Q_MX02 U4504 ( .S(oneStepPIi), .A0(ixcSimTime[63]), .A1(evfCount[63]), .Z(remStepPO[63]));
Q_MX02 U4505 ( .S(oneStepPIi), .A0(ixcSimTime[62]), .A1(evfCount[62]), .Z(remStepPO[62]));
Q_MX02 U4506 ( .S(oneStepPIi), .A0(ixcSimTime[61]), .A1(evfCount[61]), .Z(remStepPO[61]));
Q_MX02 U4507 ( .S(oneStepPIi), .A0(ixcSimTime[60]), .A1(evfCount[60]), .Z(remStepPO[60]));
Q_MX02 U4508 ( .S(oneStepPIi), .A0(ixcSimTime[59]), .A1(evfCount[59]), .Z(remStepPO[59]));
Q_MX02 U4509 ( .S(oneStepPIi), .A0(ixcSimTime[58]), .A1(evfCount[58]), .Z(remStepPO[58]));
Q_MX02 U4510 ( .S(oneStepPIi), .A0(ixcSimTime[57]), .A1(evfCount[57]), .Z(remStepPO[57]));
Q_MX02 U4511 ( .S(oneStepPIi), .A0(ixcSimTime[56]), .A1(evfCount[56]), .Z(remStepPO[56]));
Q_MX02 U4512 ( .S(oneStepPIi), .A0(ixcSimTime[55]), .A1(evfCount[55]), .Z(remStepPO[55]));
Q_MX02 U4513 ( .S(oneStepPIi), .A0(ixcSimTime[54]), .A1(evfCount[54]), .Z(remStepPO[54]));
Q_MX02 U4514 ( .S(oneStepPIi), .A0(ixcSimTime[53]), .A1(evfCount[53]), .Z(remStepPO[53]));
Q_MX02 U4515 ( .S(oneStepPIi), .A0(ixcSimTime[52]), .A1(evfCount[52]), .Z(remStepPO[52]));
Q_MX02 U4516 ( .S(oneStepPIi), .A0(ixcSimTime[51]), .A1(evfCount[51]), .Z(remStepPO[51]));
Q_MX02 U4517 ( .S(oneStepPIi), .A0(ixcSimTime[50]), .A1(evfCount[50]), .Z(remStepPO[50]));
Q_MX02 U4518 ( .S(oneStepPIi), .A0(ixcSimTime[49]), .A1(evfCount[49]), .Z(remStepPO[49]));
Q_MX02 U4519 ( .S(oneStepPIi), .A0(ixcSimTime[48]), .A1(evfCount[48]), .Z(remStepPO[48]));
Q_MX02 U4520 ( .S(oneStepPIi), .A0(ixcSimTime[47]), .A1(evfCount[47]), .Z(remStepPO[47]));
Q_MX02 U4521 ( .S(oneStepPIi), .A0(ixcSimTime[46]), .A1(evfCount[46]), .Z(remStepPO[46]));
Q_MX02 U4522 ( .S(oneStepPIi), .A0(ixcSimTime[45]), .A1(evfCount[45]), .Z(remStepPO[45]));
Q_MX02 U4523 ( .S(oneStepPIi), .A0(ixcSimTime[44]), .A1(evfCount[44]), .Z(remStepPO[44]));
Q_MX02 U4524 ( .S(oneStepPIi), .A0(ixcSimTime[43]), .A1(evfCount[43]), .Z(remStepPO[43]));
Q_MX02 U4525 ( .S(oneStepPIi), .A0(ixcSimTime[42]), .A1(evfCount[42]), .Z(remStepPO[42]));
Q_MX02 U4526 ( .S(oneStepPIi), .A0(ixcSimTime[41]), .A1(evfCount[41]), .Z(remStepPO[41]));
Q_MX02 U4527 ( .S(oneStepPIi), .A0(ixcSimTime[40]), .A1(evfCount[40]), .Z(remStepPO[40]));
Q_MX02 U4528 ( .S(oneStepPIi), .A0(ixcSimTime[39]), .A1(evfCount[39]), .Z(remStepPO[39]));
Q_MX02 U4529 ( .S(oneStepPIi), .A0(ixcSimTime[38]), .A1(evfCount[38]), .Z(remStepPO[38]));
Q_MX02 U4530 ( .S(oneStepPIi), .A0(ixcSimTime[37]), .A1(evfCount[37]), .Z(remStepPO[37]));
Q_MX02 U4531 ( .S(oneStepPIi), .A0(ixcSimTime[36]), .A1(evfCount[36]), .Z(remStepPO[36]));
Q_MX02 U4532 ( .S(oneStepPIi), .A0(ixcSimTime[35]), .A1(evfCount[35]), .Z(remStepPO[35]));
Q_MX02 U4533 ( .S(oneStepPIi), .A0(ixcSimTime[34]), .A1(evfCount[34]), .Z(remStepPO[34]));
Q_MX02 U4534 ( .S(oneStepPIi), .A0(ixcSimTime[33]), .A1(evfCount[33]), .Z(remStepPO[33]));
Q_MX02 U4535 ( .S(oneStepPIi), .A0(ixcSimTime[32]), .A1(evfCount[32]), .Z(remStepPO[32]));
Q_MX02 U4536 ( .S(oneStepPIi), .A0(ixcSimTime[31]), .A1(evfCount[31]), .Z(remStepPO[31]));
Q_MX02 U4537 ( .S(oneStepPIi), .A0(ixcSimTime[30]), .A1(evfCount[30]), .Z(remStepPO[30]));
Q_MX02 U4538 ( .S(oneStepPIi), .A0(ixcSimTime[29]), .A1(evfCount[29]), .Z(remStepPO[29]));
Q_MX02 U4539 ( .S(oneStepPIi), .A0(ixcSimTime[28]), .A1(evfCount[28]), .Z(remStepPO[28]));
Q_MX02 U4540 ( .S(oneStepPIi), .A0(ixcSimTime[27]), .A1(evfCount[27]), .Z(remStepPO[27]));
Q_MX02 U4541 ( .S(oneStepPIi), .A0(ixcSimTime[26]), .A1(evfCount[26]), .Z(remStepPO[26]));
Q_MX02 U4542 ( .S(oneStepPIi), .A0(ixcSimTime[25]), .A1(evfCount[25]), .Z(remStepPO[25]));
Q_MX02 U4543 ( .S(oneStepPIi), .A0(ixcSimTime[24]), .A1(evfCount[24]), .Z(remStepPO[24]));
Q_MX02 U4544 ( .S(oneStepPIi), .A0(ixcSimTime[23]), .A1(evfCount[23]), .Z(remStepPO[23]));
Q_MX02 U4545 ( .S(oneStepPIi), .A0(ixcSimTime[22]), .A1(evfCount[22]), .Z(remStepPO[22]));
Q_MX02 U4546 ( .S(oneStepPIi), .A0(ixcSimTime[21]), .A1(evfCount[21]), .Z(remStepPO[21]));
Q_MX02 U4547 ( .S(oneStepPIi), .A0(ixcSimTime[20]), .A1(evfCount[20]), .Z(remStepPO[20]));
Q_MX02 U4548 ( .S(oneStepPIi), .A0(ixcSimTime[19]), .A1(evfCount[19]), .Z(remStepPO[19]));
Q_MX02 U4549 ( .S(oneStepPIi), .A0(ixcSimTime[18]), .A1(evfCount[18]), .Z(remStepPO[18]));
Q_MX02 U4550 ( .S(oneStepPIi), .A0(ixcSimTime[17]), .A1(evfCount[17]), .Z(remStepPO[17]));
Q_MX02 U4551 ( .S(oneStepPIi), .A0(ixcSimTime[16]), .A1(evfCount[16]), .Z(remStepPO[16]));
Q_MX02 U4552 ( .S(oneStepPIi), .A0(ixcSimTime[15]), .A1(evfCount[15]), .Z(remStepPO[15]));
Q_MX02 U4553 ( .S(oneStepPIi), .A0(ixcSimTime[14]), .A1(evfCount[14]), .Z(remStepPO[14]));
Q_MX02 U4554 ( .S(oneStepPIi), .A0(ixcSimTime[13]), .A1(evfCount[13]), .Z(remStepPO[13]));
Q_MX02 U4555 ( .S(oneStepPIi), .A0(ixcSimTime[12]), .A1(evfCount[12]), .Z(remStepPO[12]));
Q_MX02 U4556 ( .S(oneStepPIi), .A0(ixcSimTime[11]), .A1(evfCount[11]), .Z(remStepPO[11]));
Q_MX02 U4557 ( .S(oneStepPIi), .A0(ixcSimTime[10]), .A1(evfCount[10]), .Z(remStepPO[10]));
Q_MX02 U4558 ( .S(oneStepPIi), .A0(ixcSimTime[9]), .A1(evfCount[9]), .Z(remStepPO[9]));
Q_MX02 U4559 ( .S(oneStepPIi), .A0(ixcSimTime[8]), .A1(evfCount[8]), .Z(remStepPO[8]));
Q_MX02 U4560 ( .S(oneStepPIi), .A0(ixcSimTime[7]), .A1(evfCount[7]), .Z(remStepPO[7]));
Q_MX02 U4561 ( .S(oneStepPIi), .A0(ixcSimTime[6]), .A1(evfCount[6]), .Z(remStepPO[6]));
Q_MX02 U4562 ( .S(oneStepPIi), .A0(ixcSimTime[5]), .A1(evfCount[5]), .Z(remStepPO[5]));
Q_MX02 U4563 ( .S(oneStepPIi), .A0(ixcSimTime[4]), .A1(evfCount[4]), .Z(remStepPO[4]));
Q_MX02 U4564 ( .S(oneStepPIi), .A0(ixcSimTime[3]), .A1(evfCount[3]), .Z(remStepPO[3]));
Q_MX02 U4565 ( .S(oneStepPIi), .A0(ixcSimTime[2]), .A1(evfCount[2]), .Z(remStepPO[2]));
Q_MX02 U4566 ( .S(oneStepPIi), .A0(ixcSimTime[1]), .A1(evfCount[1]), .Z(remStepPO[1]));
Q_MX02 U4567 ( .S(oneStepPIi), .A0(ixcSimTime[0]), .A1(evfCount[0]), .Z(remStepPO[0]));
Q_MX02 U4568 ( .S(n3832), .A0(n3833), .A1(stopTLd), .Z(stopTL));
Q_MX02 U4569 ( .S(n3834), .A0(stop4POd), .A1(stop4R), .Z(stop4PO));
Q_MX02 U4570 ( .S(n3835), .A0(stop2POd), .A1(stop2R), .Z(stop2PO));
Q_MX02 U4571 ( .S(n3836), .A0(stop1POd), .A1(stop1R), .Z(stop1PO));
Q_OR02 U4572 ( .A0(callEmuPre), .A1(stop4R), .Z(n3834));
Q_OR02 U4573 ( .A0(callEmuPre), .A1(stop2R), .Z(n3835));
Q_OR02 U4574 ( .A0(callEmuPre), .A1(stop1R), .Z(n3836));
Q_AO21 U4575 ( .A0(n3555), .A1(tbcPOReg), .B0(GFLock1), .Z(GFLock2R));
Q_OA21 U4576 ( .A0(GFLock2R), .A1(xcReplayOn), .B0(n3045), .Z(GFLock2));
Q_OR02 U4577 ( .A0(GFLBfull), .A1(GFGBfullBw), .Z(n3837));
Q_BUFZP U4578 ( .OE(n3837), .A(n3552), .Z(GFBw));
Q_OR02 U4579 ( .A0(callEmuWait), .A1(callEmuEv), .Z(n3839));
Q_AN02 U4580 ( .A0(callEmuWaitC), .A1(n3839), .Z(callEmuWaitN));
Q_INV U4581 ( .A(callEmuWaitC), .Z(n3838));
Q_AN02 U4582 ( .A0(n3839), .A1(n3838), .Z(callEmu));
Q_OR02 U4583 ( .A0(oneStepPIi), .A1(n2955), .Z(n3843));
Q_MX02 U4584 ( .S(callEmuEv), .A0(simTimeOn), .A1(n3843), .Z(n3844));
Q_OR03 U4585 ( .A0(hwClkDbgTime), .A1(lockTraceOn), .A2(n3844), .Z(n3840));
Q_OR03 U4586 ( .A0(lockTraceOn), .A1(callEmuEv), .A2(hwClkDbgTime), .Z(n3845));
Q_OR02 U4587 ( .A0(n3555), .A1(oneStepPIi), .Z(n3848));
Q_INV U4588 ( .A(lockTraceOn), .Z(n3846));
Q_AO21 U4589 ( .A0(n3846), .A1(n3848), .B0(hwClkDbgTime), .Z(n3847));
Q_INV U4590 ( .A(n3847), .Z(n3841));
Q_NR02 U4591 ( .A0(lockTraceOn), .A1(n3848), .Z(n3849));
Q_OR02 U4592 ( .A0(hwClkDbgTime), .A1(n3849), .Z(n3842));
Q_LDP0 \simTime_REG[0] ( .G(n3840), .D(n3976), .Q(simTime[0]), .QN( ));
Q_LDP0 \simTime_REG[1] ( .G(n3840), .D(n3974), .Q(simTime[1]), .QN( ));
Q_LDP0 \simTime_REG[2] ( .G(n3840), .D(n3972), .Q(simTime[2]), .QN(n3277));
Q_LDP0 \simTime_REG[3] ( .G(n3840), .D(n3970), .Q(simTime[3]), .QN( ));
Q_LDP0 \simTime_REG[4] ( .G(n3840), .D(n3968), .Q(simTime[4]), .QN( ));
Q_LDP0 \simTime_REG[5] ( .G(n3840), .D(n3966), .Q(simTime[5]), .QN( ));
Q_LDP0 \simTime_REG[6] ( .G(n3840), .D(n3964), .Q(simTime[6]), .QN( ));
Q_LDP0 \simTime_REG[7] ( .G(n3840), .D(n3962), .Q(simTime[7]), .QN( ));
Q_LDP0 \simTime_REG[8] ( .G(n3840), .D(n3960), .Q(simTime[8]), .QN( ));
Q_LDP0 \simTime_REG[9] ( .G(n3840), .D(n3958), .Q(simTime[9]), .QN( ));
Q_LDP0 \simTime_REG[10] ( .G(n3840), .D(n3956), .Q(simTime[10]), .QN( ));
Q_LDP0 \simTime_REG[11] ( .G(n3840), .D(n3954), .Q(simTime[11]), .QN( ));
Q_LDP0 \simTime_REG[12] ( .G(n3840), .D(n3952), .Q(simTime[12]), .QN( ));
Q_LDP0 \simTime_REG[13] ( .G(n3840), .D(n3950), .Q(simTime[13]), .QN( ));
Q_LDP0 \simTime_REG[14] ( .G(n3840), .D(n3948), .Q(simTime[14]), .QN( ));
Q_LDP0 \simTime_REG[15] ( .G(n3840), .D(n3946), .Q(simTime[15]), .QN( ));
Q_LDP0 \simTime_REG[16] ( .G(n3840), .D(n3944), .Q(simTime[16]), .QN( ));
Q_LDP0 \simTime_REG[17] ( .G(n3840), .D(n3942), .Q(simTime[17]), .QN( ));
Q_LDP0 \simTime_REG[18] ( .G(n3840), .D(n3940), .Q(simTime[18]), .QN( ));
Q_LDP0 \simTime_REG[19] ( .G(n3840), .D(n3938), .Q(simTime[19]), .QN( ));
Q_LDP0 \simTime_REG[20] ( .G(n3840), .D(n3936), .Q(simTime[20]), .QN( ));
Q_LDP0 \simTime_REG[21] ( .G(n3840), .D(n3934), .Q(simTime[21]), .QN( ));
Q_LDP0 \simTime_REG[22] ( .G(n3840), .D(n3932), .Q(simTime[22]), .QN( ));
Q_LDP0 \simTime_REG[23] ( .G(n3840), .D(n3930), .Q(simTime[23]), .QN( ));
Q_LDP0 \simTime_REG[24] ( .G(n3840), .D(n3928), .Q(simTime[24]), .QN( ));
Q_LDP0 \simTime_REG[25] ( .G(n3840), .D(n3926), .Q(simTime[25]), .QN( ));
Q_LDP0 \simTime_REG[26] ( .G(n3840), .D(n3924), .Q(simTime[26]), .QN( ));
Q_LDP0 \simTime_REG[27] ( .G(n3840), .D(n3922), .Q(simTime[27]), .QN( ));
Q_LDP0 \simTime_REG[28] ( .G(n3840), .D(n3920), .Q(simTime[28]), .QN( ));
Q_LDP0 \simTime_REG[29] ( .G(n3840), .D(n3918), .Q(simTime[29]), .QN( ));
Q_LDP0 \simTime_REG[30] ( .G(n3840), .D(n3916), .Q(simTime[30]), .QN( ));
Q_LDP0 \simTime_REG[31] ( .G(n3840), .D(n3914), .Q(simTime[31]), .QN( ));
Q_LDP0 \simTime_REG[32] ( .G(n3840), .D(n3912), .Q(simTime[32]), .QN( ));
Q_LDP0 \simTime_REG[33] ( .G(n3840), .D(n3910), .Q(simTime[33]), .QN( ));
Q_LDP0 \simTime_REG[34] ( .G(n3840), .D(n3908), .Q(simTime[34]), .QN( ));
Q_LDP0 \simTime_REG[35] ( .G(n3840), .D(n3906), .Q(simTime[35]), .QN( ));
Q_LDP0 \simTime_REG[36] ( .G(n3840), .D(n3904), .Q(simTime[36]), .QN( ));
Q_LDP0 \simTime_REG[37] ( .G(n3840), .D(n3902), .Q(simTime[37]), .QN( ));
Q_LDP0 \simTime_REG[38] ( .G(n3840), .D(n3900), .Q(simTime[38]), .QN( ));
Q_LDP0 \simTime_REG[39] ( .G(n3840), .D(n3898), .Q(simTime[39]), .QN( ));
Q_LDP0 \simTime_REG[40] ( .G(n3840), .D(n3896), .Q(simTime[40]), .QN( ));
Q_LDP0 \simTime_REG[41] ( .G(n3840), .D(n3894), .Q(simTime[41]), .QN( ));
Q_LDP0 \simTime_REG[42] ( .G(n3840), .D(n3892), .Q(simTime[42]), .QN( ));
Q_LDP0 \simTime_REG[43] ( .G(n3840), .D(n3890), .Q(simTime[43]), .QN( ));
Q_LDP0 \simTime_REG[44] ( .G(n3840), .D(n3888), .Q(simTime[44]), .QN( ));
Q_LDP0 \simTime_REG[45] ( .G(n3840), .D(n3886), .Q(simTime[45]), .QN( ));
Q_LDP0 \simTime_REG[46] ( .G(n3840), .D(n3884), .Q(simTime[46]), .QN( ));
Q_LDP0 \simTime_REG[47] ( .G(n3840), .D(n3882), .Q(simTime[47]), .QN( ));
Q_LDP0 \simTime_REG[48] ( .G(n3840), .D(n3880), .Q(simTime[48]), .QN( ));
Q_LDP0 \simTime_REG[49] ( .G(n3840), .D(n3878), .Q(simTime[49]), .QN( ));
Q_LDP0 \simTime_REG[50] ( .G(n3840), .D(n3876), .Q(simTime[50]), .QN( ));
Q_LDP0 \simTime_REG[51] ( .G(n3840), .D(n3874), .Q(simTime[51]), .QN( ));
Q_LDP0 \simTime_REG[52] ( .G(n3840), .D(n3872), .Q(simTime[52]), .QN( ));
Q_LDP0 \simTime_REG[53] ( .G(n3840), .D(n3870), .Q(simTime[53]), .QN( ));
Q_LDP0 \simTime_REG[54] ( .G(n3840), .D(n3868), .Q(simTime[54]), .QN( ));
Q_LDP0 \simTime_REG[55] ( .G(n3840), .D(n3866), .Q(simTime[55]), .QN( ));
Q_LDP0 \simTime_REG[56] ( .G(n3840), .D(n3864), .Q(simTime[56]), .QN( ));
Q_LDP0 \simTime_REG[57] ( .G(n3840), .D(n3862), .Q(simTime[57]), .QN( ));
Q_LDP0 \simTime_REG[58] ( .G(n3840), .D(n3860), .Q(simTime[58]), .QN( ));
Q_LDP0 \simTime_REG[59] ( .G(n3840), .D(n3858), .Q(simTime[59]), .QN( ));
Q_LDP0 \simTime_REG[60] ( .G(n3840), .D(n3856), .Q(simTime[60]), .QN( ));
Q_LDP0 \simTime_REG[61] ( .G(n3840), .D(n3854), .Q(simTime[61]), .QN( ));
Q_LDP0 \simTime_REG[62] ( .G(n3840), .D(n3852), .Q(simTime[62]), .QN( ));
Q_LDP0 \simTime_REG[63] ( .G(n3840), .D(n3850), .Q(simTime[63]), .QN( ));
Q_MX02 U4657 ( .S(n3845), .A0(ixcSimTime[63]), .A1(n3851), .Z(n3850));
Q_MX04 U4658 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[63]), .A1(hwSimTime[63]), .A2(lockTraceTime[63]), .A3(nextDutTimeS[63]), .Z(n3851));
Q_MX02 U4659 ( .S(n3845), .A0(ixcSimTime[62]), .A1(n3853), .Z(n3852));
Q_MX04 U4660 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[62]), .A1(hwSimTime[62]), .A2(lockTraceTime[62]), .A3(nextDutTimeS[62]), .Z(n3853));
Q_MX02 U4661 ( .S(n3845), .A0(ixcSimTime[61]), .A1(n3855), .Z(n3854));
Q_MX04 U4662 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[61]), .A1(hwSimTime[61]), .A2(lockTraceTime[61]), .A3(nextDutTimeS[61]), .Z(n3855));
Q_MX02 U4663 ( .S(n3845), .A0(ixcSimTime[60]), .A1(n3857), .Z(n3856));
Q_MX04 U4664 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[60]), .A1(hwSimTime[60]), .A2(lockTraceTime[60]), .A3(nextDutTimeS[60]), .Z(n3857));
Q_MX02 U4665 ( .S(n3845), .A0(ixcSimTime[59]), .A1(n3859), .Z(n3858));
Q_MX04 U4666 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[59]), .A1(hwSimTime[59]), .A2(lockTraceTime[59]), .A3(nextDutTimeS[59]), .Z(n3859));
Q_MX02 U4667 ( .S(n3845), .A0(ixcSimTime[58]), .A1(n3861), .Z(n3860));
Q_MX04 U4668 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[58]), .A1(hwSimTime[58]), .A2(lockTraceTime[58]), .A3(nextDutTimeS[58]), .Z(n3861));
Q_MX02 U4669 ( .S(n3845), .A0(ixcSimTime[57]), .A1(n3863), .Z(n3862));
Q_MX04 U4670 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[57]), .A1(hwSimTime[57]), .A2(lockTraceTime[57]), .A3(nextDutTimeS[57]), .Z(n3863));
Q_MX02 U4671 ( .S(n3845), .A0(ixcSimTime[56]), .A1(n3865), .Z(n3864));
Q_MX04 U4672 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[56]), .A1(hwSimTime[56]), .A2(lockTraceTime[56]), .A3(nextDutTimeS[56]), .Z(n3865));
Q_MX02 U4673 ( .S(n3845), .A0(ixcSimTime[55]), .A1(n3867), .Z(n3866));
Q_MX04 U4674 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[55]), .A1(hwSimTime[55]), .A2(lockTraceTime[55]), .A3(nextDutTimeS[55]), .Z(n3867));
Q_MX02 U4675 ( .S(n3845), .A0(ixcSimTime[54]), .A1(n3869), .Z(n3868));
Q_MX04 U4676 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[54]), .A1(hwSimTime[54]), .A2(lockTraceTime[54]), .A3(nextDutTimeS[54]), .Z(n3869));
Q_MX02 U4677 ( .S(n3845), .A0(ixcSimTime[53]), .A1(n3871), .Z(n3870));
Q_MX04 U4678 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[53]), .A1(hwSimTime[53]), .A2(lockTraceTime[53]), .A3(nextDutTimeS[53]), .Z(n3871));
Q_MX02 U4679 ( .S(n3845), .A0(ixcSimTime[52]), .A1(n3873), .Z(n3872));
Q_MX04 U4680 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[52]), .A1(hwSimTime[52]), .A2(lockTraceTime[52]), .A3(nextDutTimeS[52]), .Z(n3873));
Q_MX02 U4681 ( .S(n3845), .A0(ixcSimTime[51]), .A1(n3875), .Z(n3874));
Q_MX04 U4682 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[51]), .A1(hwSimTime[51]), .A2(lockTraceTime[51]), .A3(nextDutTimeS[51]), .Z(n3875));
Q_MX02 U4683 ( .S(n3845), .A0(ixcSimTime[50]), .A1(n3877), .Z(n3876));
Q_MX04 U4684 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[50]), .A1(hwSimTime[50]), .A2(lockTraceTime[50]), .A3(nextDutTimeS[50]), .Z(n3877));
Q_MX02 U4685 ( .S(n3845), .A0(ixcSimTime[49]), .A1(n3879), .Z(n3878));
Q_MX04 U4686 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[49]), .A1(hwSimTime[49]), .A2(lockTraceTime[49]), .A3(nextDutTimeS[49]), .Z(n3879));
Q_MX02 U4687 ( .S(n3845), .A0(ixcSimTime[48]), .A1(n3881), .Z(n3880));
Q_MX04 U4688 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[48]), .A1(hwSimTime[48]), .A2(lockTraceTime[48]), .A3(nextDutTimeS[48]), .Z(n3881));
Q_MX02 U4689 ( .S(n3845), .A0(ixcSimTime[47]), .A1(n3883), .Z(n3882));
Q_MX04 U4690 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[47]), .A1(hwSimTime[47]), .A2(lockTraceTime[47]), .A3(nextDutTimeS[47]), .Z(n3883));
Q_MX02 U4691 ( .S(n3845), .A0(ixcSimTime[46]), .A1(n3885), .Z(n3884));
Q_MX04 U4692 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[46]), .A1(hwSimTime[46]), .A2(lockTraceTime[46]), .A3(nextDutTimeS[46]), .Z(n3885));
Q_MX02 U4693 ( .S(n3845), .A0(ixcSimTime[45]), .A1(n3887), .Z(n3886));
Q_MX04 U4694 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[45]), .A1(hwSimTime[45]), .A2(lockTraceTime[45]), .A3(nextDutTimeS[45]), .Z(n3887));
Q_MX02 U4695 ( .S(n3845), .A0(ixcSimTime[44]), .A1(n3889), .Z(n3888));
Q_MX04 U4696 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[44]), .A1(hwSimTime[44]), .A2(lockTraceTime[44]), .A3(nextDutTimeS[44]), .Z(n3889));
Q_MX02 U4697 ( .S(n3845), .A0(ixcSimTime[43]), .A1(n3891), .Z(n3890));
Q_MX04 U4698 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[43]), .A1(hwSimTime[43]), .A2(lockTraceTime[43]), .A3(nextDutTimeS[43]), .Z(n3891));
Q_MX02 U4699 ( .S(n3845), .A0(ixcSimTime[42]), .A1(n3893), .Z(n3892));
Q_MX04 U4700 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[42]), .A1(hwSimTime[42]), .A2(lockTraceTime[42]), .A3(nextDutTimeS[42]), .Z(n3893));
Q_MX02 U4701 ( .S(n3845), .A0(ixcSimTime[41]), .A1(n3895), .Z(n3894));
Q_MX04 U4702 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[41]), .A1(hwSimTime[41]), .A2(lockTraceTime[41]), .A3(nextDutTimeS[41]), .Z(n3895));
Q_MX02 U4703 ( .S(n3845), .A0(ixcSimTime[40]), .A1(n3897), .Z(n3896));
Q_MX04 U4704 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[40]), .A1(hwSimTime[40]), .A2(lockTraceTime[40]), .A3(nextDutTimeS[40]), .Z(n3897));
Q_MX02 U4705 ( .S(n3845), .A0(ixcSimTime[39]), .A1(n3899), .Z(n3898));
Q_MX04 U4706 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[39]), .A1(hwSimTime[39]), .A2(lockTraceTime[39]), .A3(nextDutTimeS[39]), .Z(n3899));
Q_MX02 U4707 ( .S(n3845), .A0(ixcSimTime[38]), .A1(n3901), .Z(n3900));
Q_MX04 U4708 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[38]), .A1(hwSimTime[38]), .A2(lockTraceTime[38]), .A3(nextDutTimeS[38]), .Z(n3901));
Q_MX02 U4709 ( .S(n3845), .A0(ixcSimTime[37]), .A1(n3903), .Z(n3902));
Q_MX04 U4710 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[37]), .A1(hwSimTime[37]), .A2(lockTraceTime[37]), .A3(nextDutTimeS[37]), .Z(n3903));
Q_MX02 U4711 ( .S(n3845), .A0(ixcSimTime[36]), .A1(n3905), .Z(n3904));
Q_MX04 U4712 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[36]), .A1(hwSimTime[36]), .A2(lockTraceTime[36]), .A3(nextDutTimeS[36]), .Z(n3905));
Q_MX02 U4713 ( .S(n3845), .A0(ixcSimTime[35]), .A1(n3907), .Z(n3906));
Q_MX04 U4714 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[35]), .A1(hwSimTime[35]), .A2(lockTraceTime[35]), .A3(nextDutTimeS[35]), .Z(n3907));
Q_MX02 U4715 ( .S(n3845), .A0(ixcSimTime[34]), .A1(n3909), .Z(n3908));
Q_MX04 U4716 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[34]), .A1(hwSimTime[34]), .A2(lockTraceTime[34]), .A3(nextDutTimeS[34]), .Z(n3909));
Q_MX02 U4717 ( .S(n3845), .A0(ixcSimTime[33]), .A1(n3911), .Z(n3910));
Q_MX04 U4718 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[33]), .A1(hwSimTime[33]), .A2(lockTraceTime[33]), .A3(nextDutTimeS[33]), .Z(n3911));
Q_MX02 U4719 ( .S(n3845), .A0(ixcSimTime[32]), .A1(n3913), .Z(n3912));
Q_MX04 U4720 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[32]), .A1(hwSimTime[32]), .A2(lockTraceTime[32]), .A3(nextDutTimeS[32]), .Z(n3913));
Q_MX02 U4721 ( .S(n3845), .A0(ixcSimTime[31]), .A1(n3915), .Z(n3914));
Q_MX04 U4722 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[31]), .A1(hwSimTime[31]), .A2(lockTraceTime[31]), .A3(nextDutTimeS[31]), .Z(n3915));
Q_MX02 U4723 ( .S(n3845), .A0(ixcSimTime[30]), .A1(n3917), .Z(n3916));
Q_MX04 U4724 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[30]), .A1(hwSimTime[30]), .A2(lockTraceTime[30]), .A3(nextDutTimeS[30]), .Z(n3917));
Q_MX02 U4725 ( .S(n3845), .A0(ixcSimTime[29]), .A1(n3919), .Z(n3918));
Q_MX04 U4726 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[29]), .A1(hwSimTime[29]), .A2(lockTraceTime[29]), .A3(nextDutTimeS[29]), .Z(n3919));
Q_MX02 U4727 ( .S(n3845), .A0(ixcSimTime[28]), .A1(n3921), .Z(n3920));
Q_MX04 U4728 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[28]), .A1(hwSimTime[28]), .A2(lockTraceTime[28]), .A3(nextDutTimeS[28]), .Z(n3921));
Q_MX02 U4729 ( .S(n3845), .A0(ixcSimTime[27]), .A1(n3923), .Z(n3922));
Q_MX04 U4730 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[27]), .A1(hwSimTime[27]), .A2(lockTraceTime[27]), .A3(nextDutTimeS[27]), .Z(n3923));
Q_MX02 U4731 ( .S(n3845), .A0(ixcSimTime[26]), .A1(n3925), .Z(n3924));
Q_MX04 U4732 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[26]), .A1(hwSimTime[26]), .A2(lockTraceTime[26]), .A3(nextDutTimeS[26]), .Z(n3925));
Q_MX02 U4733 ( .S(n3845), .A0(ixcSimTime[25]), .A1(n3927), .Z(n3926));
Q_MX04 U4734 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[25]), .A1(hwSimTime[25]), .A2(lockTraceTime[25]), .A3(nextDutTimeS[25]), .Z(n3927));
Q_MX02 U4735 ( .S(n3845), .A0(ixcSimTime[24]), .A1(n3929), .Z(n3928));
Q_MX04 U4736 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[24]), .A1(hwSimTime[24]), .A2(lockTraceTime[24]), .A3(nextDutTimeS[24]), .Z(n3929));
Q_MX02 U4737 ( .S(n3845), .A0(ixcSimTime[23]), .A1(n3931), .Z(n3930));
Q_MX04 U4738 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[23]), .A1(hwSimTime[23]), .A2(lockTraceTime[23]), .A3(nextDutTimeS[23]), .Z(n3931));
Q_MX02 U4739 ( .S(n3845), .A0(ixcSimTime[22]), .A1(n3933), .Z(n3932));
Q_MX04 U4740 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[22]), .A1(hwSimTime[22]), .A2(lockTraceTime[22]), .A3(nextDutTimeS[22]), .Z(n3933));
Q_MX02 U4741 ( .S(n3845), .A0(ixcSimTime[21]), .A1(n3935), .Z(n3934));
Q_MX04 U4742 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[21]), .A1(hwSimTime[21]), .A2(lockTraceTime[21]), .A3(nextDutTimeS[21]), .Z(n3935));
Q_MX02 U4743 ( .S(n3845), .A0(ixcSimTime[20]), .A1(n3937), .Z(n3936));
Q_MX04 U4744 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[20]), .A1(hwSimTime[20]), .A2(lockTraceTime[20]), .A3(nextDutTimeS[20]), .Z(n3937));
Q_MX02 U4745 ( .S(n3845), .A0(ixcSimTime[19]), .A1(n3939), .Z(n3938));
Q_MX04 U4746 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[19]), .A1(hwSimTime[19]), .A2(lockTraceTime[19]), .A3(nextDutTimeS[19]), .Z(n3939));
Q_MX02 U4747 ( .S(n3845), .A0(ixcSimTime[18]), .A1(n3941), .Z(n3940));
Q_MX04 U4748 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[18]), .A1(hwSimTime[18]), .A2(lockTraceTime[18]), .A3(nextDutTimeS[18]), .Z(n3941));
Q_MX02 U4749 ( .S(n3845), .A0(ixcSimTime[17]), .A1(n3943), .Z(n3942));
Q_MX04 U4750 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[17]), .A1(hwSimTime[17]), .A2(lockTraceTime[17]), .A3(nextDutTimeS[17]), .Z(n3943));
Q_MX02 U4751 ( .S(n3845), .A0(ixcSimTime[16]), .A1(n3945), .Z(n3944));
Q_MX04 U4752 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[16]), .A1(hwSimTime[16]), .A2(lockTraceTime[16]), .A3(nextDutTimeS[16]), .Z(n3945));
Q_MX02 U4753 ( .S(n3845), .A0(ixcSimTime[15]), .A1(n3947), .Z(n3946));
Q_MX04 U4754 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[15]), .A1(hwSimTime[15]), .A2(lockTraceTime[15]), .A3(nextDutTimeS[15]), .Z(n3947));
Q_MX02 U4755 ( .S(n3845), .A0(ixcSimTime[14]), .A1(n3949), .Z(n3948));
Q_MX04 U4756 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[14]), .A1(hwSimTime[14]), .A2(lockTraceTime[14]), .A3(nextDutTimeS[14]), .Z(n3949));
Q_MX02 U4757 ( .S(n3845), .A0(ixcSimTime[13]), .A1(n3951), .Z(n3950));
Q_MX04 U4758 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[13]), .A1(hwSimTime[13]), .A2(lockTraceTime[13]), .A3(nextDutTimeS[13]), .Z(n3951));
Q_MX02 U4759 ( .S(n3845), .A0(ixcSimTime[12]), .A1(n3953), .Z(n3952));
Q_MX04 U4760 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[12]), .A1(hwSimTime[12]), .A2(lockTraceTime[12]), .A3(nextDutTimeS[12]), .Z(n3953));
Q_MX02 U4761 ( .S(n3845), .A0(ixcSimTime[11]), .A1(n3955), .Z(n3954));
Q_MX04 U4762 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[11]), .A1(hwSimTime[11]), .A2(lockTraceTime[11]), .A3(nextDutTimeS[11]), .Z(n3955));
Q_MX02 U4763 ( .S(n3845), .A0(ixcSimTime[10]), .A1(n3957), .Z(n3956));
Q_MX04 U4764 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[10]), .A1(hwSimTime[10]), .A2(lockTraceTime[10]), .A3(nextDutTimeS[10]), .Z(n3957));
Q_MX02 U4765 ( .S(n3845), .A0(ixcSimTime[9]), .A1(n3959), .Z(n3958));
Q_MX04 U4766 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[9]), .A1(hwSimTime[9]), .A2(lockTraceTime[9]), .A3(nextDutTimeS[9]), .Z(n3959));
Q_MX02 U4767 ( .S(n3845), .A0(ixcSimTime[8]), .A1(n3961), .Z(n3960));
Q_MX04 U4768 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[8]), .A1(hwSimTime[8]), .A2(lockTraceTime[8]), .A3(nextDutTimeS[8]), .Z(n3961));
Q_MX02 U4769 ( .S(n3845), .A0(ixcSimTime[7]), .A1(n3963), .Z(n3962));
Q_MX04 U4770 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[7]), .A1(hwSimTime[7]), .A2(lockTraceTime[7]), .A3(nextDutTimeS[7]), .Z(n3963));
Q_MX02 U4771 ( .S(n3845), .A0(ixcSimTime[6]), .A1(n3965), .Z(n3964));
Q_MX04 U4772 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[6]), .A1(hwSimTime[6]), .A2(lockTraceTime[6]), .A3(nextDutTimeS[6]), .Z(n3965));
Q_MX02 U4773 ( .S(n3845), .A0(ixcSimTime[5]), .A1(n3967), .Z(n3966));
Q_MX04 U4774 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[5]), .A1(hwSimTime[5]), .A2(lockTraceTime[5]), .A3(nextDutTimeS[5]), .Z(n3967));
Q_MX02 U4775 ( .S(n3845), .A0(ixcSimTime[4]), .A1(n3969), .Z(n3968));
Q_MX04 U4776 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[4]), .A1(hwSimTime[4]), .A2(lockTraceTime[4]), .A3(nextDutTimeS[4]), .Z(n3969));
Q_MX02 U4777 ( .S(n3845), .A0(ixcSimTime[3]), .A1(n3971), .Z(n3970));
Q_MX04 U4778 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[3]), .A1(hwSimTime[3]), .A2(lockTraceTime[3]), .A3(nextDutTimeS[3]), .Z(n3971));
Q_MX02 U4779 ( .S(n3845), .A0(ixcSimTime[2]), .A1(n3973), .Z(n3972));
Q_MX04 U4780 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[2]), .A1(hwSimTime[2]), .A2(lockTraceTime[2]), .A3(nextDutTimeS[2]), .Z(n3973));
Q_MX02 U4781 ( .S(n3845), .A0(ixcSimTime[1]), .A1(n3975), .Z(n3974));
Q_MX04 U4782 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[1]), .A1(hwSimTime[1]), .A2(lockTraceTime[1]), .A3(nextDutTimeS[1]), .Z(n3975));
Q_MX02 U4783 ( .S(n3845), .A0(ixcSimTime[0]), .A1(n3977), .Z(n3976));
Q_MX04 U4784 ( .S0(n3842), .S1(n3841), .A0(ixc_time.nextTbTime[0]), .A1(hwSimTime[0]), .A2(lockTraceTime[0]), .A3(nextDutTimeS[0]), .Z(n3977));
Q_MX02 U4785 ( .S(oneStepPIi), .A0(ixc_time.simTime[63]), .A1(ixc_time.nextTbTime[63]), .Z(ixcSimTime[63]));
Q_MX02 U4786 ( .S(oneStepPIi), .A0(ixc_time.simTime[62]), .A1(ixc_time.nextTbTime[62]), .Z(ixcSimTime[62]));
Q_MX02 U4787 ( .S(oneStepPIi), .A0(ixc_time.simTime[61]), .A1(ixc_time.nextTbTime[61]), .Z(ixcSimTime[61]));
Q_MX02 U4788 ( .S(oneStepPIi), .A0(ixc_time.simTime[60]), .A1(ixc_time.nextTbTime[60]), .Z(ixcSimTime[60]));
Q_MX02 U4789 ( .S(oneStepPIi), .A0(ixc_time.simTime[59]), .A1(ixc_time.nextTbTime[59]), .Z(ixcSimTime[59]));
Q_MX02 U4790 ( .S(oneStepPIi), .A0(ixc_time.simTime[58]), .A1(ixc_time.nextTbTime[58]), .Z(ixcSimTime[58]));
Q_MX02 U4791 ( .S(oneStepPIi), .A0(ixc_time.simTime[57]), .A1(ixc_time.nextTbTime[57]), .Z(ixcSimTime[57]));
Q_MX02 U4792 ( .S(oneStepPIi), .A0(ixc_time.simTime[56]), .A1(ixc_time.nextTbTime[56]), .Z(ixcSimTime[56]));
Q_MX02 U4793 ( .S(oneStepPIi), .A0(ixc_time.simTime[55]), .A1(ixc_time.nextTbTime[55]), .Z(ixcSimTime[55]));
Q_MX02 U4794 ( .S(oneStepPIi), .A0(ixc_time.simTime[54]), .A1(ixc_time.nextTbTime[54]), .Z(ixcSimTime[54]));
Q_MX02 U4795 ( .S(oneStepPIi), .A0(ixc_time.simTime[53]), .A1(ixc_time.nextTbTime[53]), .Z(ixcSimTime[53]));
Q_MX02 U4796 ( .S(oneStepPIi), .A0(ixc_time.simTime[52]), .A1(ixc_time.nextTbTime[52]), .Z(ixcSimTime[52]));
Q_MX02 U4797 ( .S(oneStepPIi), .A0(ixc_time.simTime[51]), .A1(ixc_time.nextTbTime[51]), .Z(ixcSimTime[51]));
Q_MX02 U4798 ( .S(oneStepPIi), .A0(ixc_time.simTime[50]), .A1(ixc_time.nextTbTime[50]), .Z(ixcSimTime[50]));
Q_MX02 U4799 ( .S(oneStepPIi), .A0(ixc_time.simTime[49]), .A1(ixc_time.nextTbTime[49]), .Z(ixcSimTime[49]));
Q_MX02 U4800 ( .S(oneStepPIi), .A0(ixc_time.simTime[48]), .A1(ixc_time.nextTbTime[48]), .Z(ixcSimTime[48]));
Q_MX02 U4801 ( .S(oneStepPIi), .A0(ixc_time.simTime[47]), .A1(ixc_time.nextTbTime[47]), .Z(ixcSimTime[47]));
Q_MX02 U4802 ( .S(oneStepPIi), .A0(ixc_time.simTime[46]), .A1(ixc_time.nextTbTime[46]), .Z(ixcSimTime[46]));
Q_MX02 U4803 ( .S(oneStepPIi), .A0(ixc_time.simTime[45]), .A1(ixc_time.nextTbTime[45]), .Z(ixcSimTime[45]));
Q_MX02 U4804 ( .S(oneStepPIi), .A0(ixc_time.simTime[44]), .A1(ixc_time.nextTbTime[44]), .Z(ixcSimTime[44]));
Q_MX02 U4805 ( .S(oneStepPIi), .A0(ixc_time.simTime[43]), .A1(ixc_time.nextTbTime[43]), .Z(ixcSimTime[43]));
Q_MX02 U4806 ( .S(oneStepPIi), .A0(ixc_time.simTime[42]), .A1(ixc_time.nextTbTime[42]), .Z(ixcSimTime[42]));
Q_MX02 U4807 ( .S(oneStepPIi), .A0(ixc_time.simTime[41]), .A1(ixc_time.nextTbTime[41]), .Z(ixcSimTime[41]));
Q_MX02 U4808 ( .S(oneStepPIi), .A0(ixc_time.simTime[40]), .A1(ixc_time.nextTbTime[40]), .Z(ixcSimTime[40]));
Q_MX02 U4809 ( .S(oneStepPIi), .A0(ixc_time.simTime[39]), .A1(ixc_time.nextTbTime[39]), .Z(ixcSimTime[39]));
Q_MX02 U4810 ( .S(oneStepPIi), .A0(ixc_time.simTime[38]), .A1(ixc_time.nextTbTime[38]), .Z(ixcSimTime[38]));
Q_MX02 U4811 ( .S(oneStepPIi), .A0(ixc_time.simTime[37]), .A1(ixc_time.nextTbTime[37]), .Z(ixcSimTime[37]));
Q_MX02 U4812 ( .S(oneStepPIi), .A0(ixc_time.simTime[36]), .A1(ixc_time.nextTbTime[36]), .Z(ixcSimTime[36]));
Q_MX02 U4813 ( .S(oneStepPIi), .A0(ixc_time.simTime[35]), .A1(ixc_time.nextTbTime[35]), .Z(ixcSimTime[35]));
Q_MX02 U4814 ( .S(oneStepPIi), .A0(ixc_time.simTime[34]), .A1(ixc_time.nextTbTime[34]), .Z(ixcSimTime[34]));
Q_MX02 U4815 ( .S(oneStepPIi), .A0(ixc_time.simTime[33]), .A1(ixc_time.nextTbTime[33]), .Z(ixcSimTime[33]));
Q_MX02 U4816 ( .S(oneStepPIi), .A0(ixc_time.simTime[32]), .A1(ixc_time.nextTbTime[32]), .Z(ixcSimTime[32]));
Q_MX02 U4817 ( .S(oneStepPIi), .A0(ixc_time.simTime[31]), .A1(ixc_time.nextTbTime[31]), .Z(ixcSimTime[31]));
Q_MX02 U4818 ( .S(oneStepPIi), .A0(ixc_time.simTime[30]), .A1(ixc_time.nextTbTime[30]), .Z(ixcSimTime[30]));
Q_MX02 U4819 ( .S(oneStepPIi), .A0(ixc_time.simTime[29]), .A1(ixc_time.nextTbTime[29]), .Z(ixcSimTime[29]));
Q_MX02 U4820 ( .S(oneStepPIi), .A0(ixc_time.simTime[28]), .A1(ixc_time.nextTbTime[28]), .Z(ixcSimTime[28]));
Q_MX02 U4821 ( .S(oneStepPIi), .A0(ixc_time.simTime[27]), .A1(ixc_time.nextTbTime[27]), .Z(ixcSimTime[27]));
Q_MX02 U4822 ( .S(oneStepPIi), .A0(ixc_time.simTime[26]), .A1(ixc_time.nextTbTime[26]), .Z(ixcSimTime[26]));
Q_MX02 U4823 ( .S(oneStepPIi), .A0(ixc_time.simTime[25]), .A1(ixc_time.nextTbTime[25]), .Z(ixcSimTime[25]));
Q_MX02 U4824 ( .S(oneStepPIi), .A0(ixc_time.simTime[24]), .A1(ixc_time.nextTbTime[24]), .Z(ixcSimTime[24]));
Q_MX02 U4825 ( .S(oneStepPIi), .A0(ixc_time.simTime[23]), .A1(ixc_time.nextTbTime[23]), .Z(ixcSimTime[23]));
Q_MX02 U4826 ( .S(oneStepPIi), .A0(ixc_time.simTime[22]), .A1(ixc_time.nextTbTime[22]), .Z(ixcSimTime[22]));
Q_MX02 U4827 ( .S(oneStepPIi), .A0(ixc_time.simTime[21]), .A1(ixc_time.nextTbTime[21]), .Z(ixcSimTime[21]));
Q_MX02 U4828 ( .S(oneStepPIi), .A0(ixc_time.simTime[20]), .A1(ixc_time.nextTbTime[20]), .Z(ixcSimTime[20]));
Q_MX02 U4829 ( .S(oneStepPIi), .A0(ixc_time.simTime[19]), .A1(ixc_time.nextTbTime[19]), .Z(ixcSimTime[19]));
Q_MX02 U4830 ( .S(oneStepPIi), .A0(ixc_time.simTime[18]), .A1(ixc_time.nextTbTime[18]), .Z(ixcSimTime[18]));
Q_MX02 U4831 ( .S(oneStepPIi), .A0(ixc_time.simTime[17]), .A1(ixc_time.nextTbTime[17]), .Z(ixcSimTime[17]));
Q_MX02 U4832 ( .S(oneStepPIi), .A0(ixc_time.simTime[16]), .A1(ixc_time.nextTbTime[16]), .Z(ixcSimTime[16]));
Q_MX02 U4833 ( .S(oneStepPIi), .A0(ixc_time.simTime[15]), .A1(ixc_time.nextTbTime[15]), .Z(ixcSimTime[15]));
Q_MX02 U4834 ( .S(oneStepPIi), .A0(ixc_time.simTime[14]), .A1(ixc_time.nextTbTime[14]), .Z(ixcSimTime[14]));
Q_MX02 U4835 ( .S(oneStepPIi), .A0(ixc_time.simTime[13]), .A1(ixc_time.nextTbTime[13]), .Z(ixcSimTime[13]));
Q_MX02 U4836 ( .S(oneStepPIi), .A0(ixc_time.simTime[12]), .A1(ixc_time.nextTbTime[12]), .Z(ixcSimTime[12]));
Q_MX02 U4837 ( .S(oneStepPIi), .A0(ixc_time.simTime[11]), .A1(ixc_time.nextTbTime[11]), .Z(ixcSimTime[11]));
Q_MX02 U4838 ( .S(oneStepPIi), .A0(ixc_time.simTime[10]), .A1(ixc_time.nextTbTime[10]), .Z(ixcSimTime[10]));
Q_MX02 U4839 ( .S(oneStepPIi), .A0(ixc_time.simTime[9]), .A1(ixc_time.nextTbTime[9]), .Z(ixcSimTime[9]));
Q_MX02 U4840 ( .S(oneStepPIi), .A0(ixc_time.simTime[8]), .A1(ixc_time.nextTbTime[8]), .Z(ixcSimTime[8]));
Q_MX02 U4841 ( .S(oneStepPIi), .A0(ixc_time.simTime[7]), .A1(ixc_time.nextTbTime[7]), .Z(ixcSimTime[7]));
Q_MX02 U4842 ( .S(oneStepPIi), .A0(ixc_time.simTime[6]), .A1(ixc_time.nextTbTime[6]), .Z(ixcSimTime[6]));
Q_MX02 U4843 ( .S(oneStepPIi), .A0(ixc_time.simTime[5]), .A1(ixc_time.nextTbTime[5]), .Z(ixcSimTime[5]));
Q_MX02 U4844 ( .S(oneStepPIi), .A0(ixc_time.simTime[4]), .A1(ixc_time.nextTbTime[4]), .Z(ixcSimTime[4]));
Q_MX02 U4845 ( .S(oneStepPIi), .A0(ixc_time.simTime[3]), .A1(ixc_time.nextTbTime[3]), .Z(ixcSimTime[3]));
Q_MX02 U4846 ( .S(oneStepPIi), .A0(ixc_time.simTime[2]), .A1(ixc_time.nextTbTime[2]), .Z(ixcSimTime[2]));
Q_MX02 U4847 ( .S(oneStepPIi), .A0(ixc_time.simTime[1]), .A1(ixc_time.nextTbTime[1]), .Z(ixcSimTime[1]));
Q_MX02 U4848 ( .S(oneStepPIi), .A0(ixc_time.simTime[0]), .A1(ixc_time.nextTbTime[0]), .Z(ixcSimTime[0]));
Q_LDP0 oneStepPImio_REG  ( .G(n3978), .D(mioPIW_1[4]), .Q(oneStepPImio), .QN( ));
Q_LDP0 ckgHoldPImio_REG  ( .G(n3978), .D(mioPIW_1[2]), .Q(ckgHoldPImio), .QN( ));
Q_LDP0 callEmuPImio_REG  ( .G(n3978), .D(mioPIW_1[1]), .Q(callEmuPImio), .QN( ));
Q_LDP0 \evalStepPImio_REG[0] ( .G(n3978), .D(mioPIW_0[0]), .Q(evalStepPImio[0]), .QN( ));
Q_LDP0 \evalStepPImio_REG[1] ( .G(n3978), .D(mioPIW_0[1]), .Q(evalStepPImio[1]), .QN( ));
Q_LDP0 \evalStepPImio_REG[2] ( .G(n3978), .D(mioPIW_0[2]), .Q(evalStepPImio[2]), .QN( ));
Q_LDP0 \evalStepPImio_REG[3] ( .G(n3978), .D(mioPIW_0[3]), .Q(evalStepPImio[3]), .QN( ));
Q_LDP0 \evalStepPImio_REG[4] ( .G(n3978), .D(mioPIW_0[4]), .Q(evalStepPImio[4]), .QN( ));
Q_LDP0 \evalStepPImio_REG[5] ( .G(n3978), .D(mioPIW_0[5]), .Q(evalStepPImio[5]), .QN( ));
Q_LDP0 \evalStepPImio_REG[6] ( .G(n3978), .D(mioPIW_0[6]), .Q(evalStepPImio[6]), .QN( ));
Q_LDP0 \evalStepPImio_REG[7] ( .G(n3978), .D(mioPIW_0[7]), .Q(evalStepPImio[7]), .QN( ));
Q_LDP0 \evalStepPImio_REG[8] ( .G(n3978), .D(mioPIW_0[8]), .Q(evalStepPImio[8]), .QN( ));
Q_LDP0 \evalStepPImio_REG[9] ( .G(n3978), .D(mioPIW_0[9]), .Q(evalStepPImio[9]), .QN( ));
Q_LDP0 \evalStepPImio_REG[10] ( .G(n3978), .D(mioPIW_0[10]), .Q(evalStepPImio[10]), .QN( ));
Q_LDP0 \evalStepPImio_REG[11] ( .G(n3978), .D(mioPIW_0[11]), .Q(evalStepPImio[11]), .QN( ));
Q_LDP0 \evalStepPImio_REG[12] ( .G(n3978), .D(mioPIW_0[12]), .Q(evalStepPImio[12]), .QN( ));
Q_LDP0 \evalStepPImio_REG[13] ( .G(n3978), .D(mioPIW_0[13]), .Q(evalStepPImio[13]), .QN( ));
Q_LDP0 \evalStepPImio_REG[14] ( .G(n3978), .D(mioPIW_0[14]), .Q(evalStepPImio[14]), .QN( ));
Q_LDP0 \evalStepPImio_REG[15] ( .G(n3978), .D(mioPIW_0[15]), .Q(evalStepPImio[15]), .QN( ));
Q_LDP0 \evalStepPImio_REG[16] ( .G(n3978), .D(mioPIW_0[16]), .Q(evalStepPImio[16]), .QN( ));
Q_LDP0 \evalStepPImio_REG[17] ( .G(n3978), .D(mioPIW_0[17]), .Q(evalStepPImio[17]), .QN( ));
Q_LDP0 \evalStepPImio_REG[18] ( .G(n3978), .D(mioPIW_0[18]), .Q(evalStepPImio[18]), .QN( ));
Q_LDP0 \evalStepPImio_REG[19] ( .G(n3978), .D(mioPIW_0[19]), .Q(evalStepPImio[19]), .QN( ));
Q_LDP0 \evalStepPImio_REG[20] ( .G(n3978), .D(mioPIW_0[20]), .Q(evalStepPImio[20]), .QN( ));
Q_LDP0 \evalStepPImio_REG[21] ( .G(n3978), .D(mioPIW_0[21]), .Q(evalStepPImio[21]), .QN( ));
Q_LDP0 \evalStepPImio_REG[22] ( .G(n3978), .D(mioPIW_0[22]), .Q(evalStepPImio[22]), .QN( ));
Q_LDP0 \evalStepPImio_REG[23] ( .G(n3978), .D(mioPIW_0[23]), .Q(evalStepPImio[23]), .QN( ));
Q_LDP0 \evalStepPImio_REG[24] ( .G(n3978), .D(mioPIW_0[24]), .Q(evalStepPImio[24]), .QN( ));
Q_LDP0 \evalStepPImio_REG[25] ( .G(n3978), .D(mioPIW_0[25]), .Q(evalStepPImio[25]), .QN( ));
Q_LDP0 \evalStepPImio_REG[26] ( .G(n3978), .D(mioPIW_0[26]), .Q(evalStepPImio[26]), .QN( ));
Q_LDP0 \evalStepPImio_REG[27] ( .G(n3978), .D(mioPIW_0[27]), .Q(evalStepPImio[27]), .QN( ));
Q_LDP0 \evalStepPImio_REG[28] ( .G(n3978), .D(mioPIW_0[28]), .Q(evalStepPImio[28]), .QN( ));
Q_LDP0 \evalStepPImio_REG[29] ( .G(n3978), .D(mioPIW_0[29]), .Q(evalStepPImio[29]), .QN( ));
Q_LDP0 \evalStepPImio_REG[30] ( .G(n3978), .D(mioPIW_0[30]), .Q(evalStepPImio[30]), .QN( ));
Q_LDP0 \evalStepPImio_REG[31] ( .G(n3978), .D(mioPIW_0[31]), .Q(evalStepPImio[31]), .QN( ));
Q_LDP0 \evalStepPImio_REG[32] ( .G(n3978), .D(mioPIW_0[32]), .Q(evalStepPImio[32]), .QN( ));
Q_LDP0 \evalStepPImio_REG[33] ( .G(n3978), .D(mioPIW_0[33]), .Q(evalStepPImio[33]), .QN( ));
Q_LDP0 \evalStepPImio_REG[34] ( .G(n3978), .D(mioPIW_0[34]), .Q(evalStepPImio[34]), .QN( ));
Q_LDP0 \evalStepPImio_REG[35] ( .G(n3978), .D(mioPIW_0[35]), .Q(evalStepPImio[35]), .QN( ));
Q_LDP0 \evalStepPImio_REG[36] ( .G(n3978), .D(mioPIW_0[36]), .Q(evalStepPImio[36]), .QN( ));
Q_LDP0 \evalStepPImio_REG[37] ( .G(n3978), .D(mioPIW_0[37]), .Q(evalStepPImio[37]), .QN( ));
Q_LDP0 \evalStepPImio_REG[38] ( .G(n3978), .D(mioPIW_0[38]), .Q(evalStepPImio[38]), .QN( ));
Q_LDP0 \evalStepPImio_REG[39] ( .G(n3978), .D(mioPIW_0[39]), .Q(evalStepPImio[39]), .QN( ));
Q_LDP0 \evalStepPImio_REG[40] ( .G(n3978), .D(mioPIW_0[40]), .Q(evalStepPImio[40]), .QN( ));
Q_LDP0 \evalStepPImio_REG[41] ( .G(n3978), .D(mioPIW_0[41]), .Q(evalStepPImio[41]), .QN( ));
Q_LDP0 \evalStepPImio_REG[42] ( .G(n3978), .D(mioPIW_0[42]), .Q(evalStepPImio[42]), .QN( ));
Q_LDP0 \evalStepPImio_REG[43] ( .G(n3978), .D(mioPIW_0[43]), .Q(evalStepPImio[43]), .QN( ));
Q_LDP0 \evalStepPImio_REG[44] ( .G(n3978), .D(mioPIW_0[44]), .Q(evalStepPImio[44]), .QN( ));
Q_LDP0 \evalStepPImio_REG[45] ( .G(n3978), .D(mioPIW_0[45]), .Q(evalStepPImio[45]), .QN( ));
Q_LDP0 \evalStepPImio_REG[46] ( .G(n3978), .D(mioPIW_0[46]), .Q(evalStepPImio[46]), .QN( ));
Q_LDP0 \evalStepPImio_REG[47] ( .G(n3978), .D(mioPIW_0[47]), .Q(evalStepPImio[47]), .QN( ));
Q_LDP0 \evalStepPImio_REG[48] ( .G(n3978), .D(mioPIW_0[48]), .Q(evalStepPImio[48]), .QN( ));
Q_LDP0 \evalStepPImio_REG[49] ( .G(n3978), .D(mioPIW_0[49]), .Q(evalStepPImio[49]), .QN( ));
Q_LDP0 \evalStepPImio_REG[50] ( .G(n3978), .D(mioPIW_0[50]), .Q(evalStepPImio[50]), .QN( ));
Q_LDP0 \evalStepPImio_REG[51] ( .G(n3978), .D(mioPIW_0[51]), .Q(evalStepPImio[51]), .QN( ));
Q_LDP0 \evalStepPImio_REG[52] ( .G(n3978), .D(mioPIW_0[52]), .Q(evalStepPImio[52]), .QN( ));
Q_LDP0 \evalStepPImio_REG[53] ( .G(n3978), .D(mioPIW_0[53]), .Q(evalStepPImio[53]), .QN( ));
Q_LDP0 \evalStepPImio_REG[54] ( .G(n3978), .D(mioPIW_0[54]), .Q(evalStepPImio[54]), .QN( ));
Q_LDP0 \evalStepPImio_REG[55] ( .G(n3978), .D(mioPIW_0[55]), .Q(evalStepPImio[55]), .QN( ));
Q_LDP0 \evalStepPImio_REG[56] ( .G(n3978), .D(mioPIW_0[56]), .Q(evalStepPImio[56]), .QN( ));
Q_LDP0 \evalStepPImio_REG[57] ( .G(n3978), .D(mioPIW_0[57]), .Q(evalStepPImio[57]), .QN( ));
Q_LDP0 \evalStepPImio_REG[58] ( .G(n3978), .D(mioPIW_0[58]), .Q(evalStepPImio[58]), .QN( ));
Q_LDP0 \evalStepPImio_REG[59] ( .G(n3978), .D(mioPIW_0[59]), .Q(evalStepPImio[59]), .QN( ));
Q_LDP0 \evalStepPImio_REG[60] ( .G(n3978), .D(mioPIW_0[60]), .Q(evalStepPImio[60]), .QN( ));
Q_LDP0 \evalStepPImio_REG[61] ( .G(n3978), .D(mioPIW_0[61]), .Q(evalStepPImio[61]), .QN( ));
Q_LDP0 \evalStepPImio_REG[62] ( .G(n3978), .D(mioPIW_0[62]), .Q(evalStepPImio[62]), .QN( ));
Q_LDP0 \evalStepPImio_REG[63] ( .G(n3978), .D(mioPIW_0[63]), .Q(evalStepPImio[63]), .QN( ));
Q_XOR2 U4916 ( .A0(mioPICnt), .A1(mioPICntd), .Z(n3978));
Q_MX02 U4917 ( .S(xc_mioOn), .A0(oneStepPI), .A1(oneStepPImio), .Z(oneStepPIi));
Q_MX02 U4918 ( .S(xc_mioOn), .A0(stopEmuPI), .A1(mioPIW_1[3]), .Z(stopEmuPIi));
Q_MX02 U4919 ( .S(xc_mioOn), .A0(ckgHoldPI), .A1(ckgHoldPImio), .Z(ckgHoldPIi));
Q_MX02 U4920 ( .S(xc_mioOn), .A0(callEmuPI), .A1(callEmuPImio), .Z(callEmuPIi));
Q_MX02 U4921 ( .S(xc_mioOn), .A0(evalStepPI[63]), .A1(evalStepPImio[63]), .Z(evalStepPIi[63]));
Q_MX02 U4922 ( .S(xc_mioOn), .A0(evalStepPI[62]), .A1(evalStepPImio[62]), .Z(evalStepPIi[62]));
Q_MX02 U4923 ( .S(xc_mioOn), .A0(evalStepPI[61]), .A1(evalStepPImio[61]), .Z(evalStepPIi[61]));
Q_MX02 U4924 ( .S(xc_mioOn), .A0(evalStepPI[60]), .A1(evalStepPImio[60]), .Z(evalStepPIi[60]));
Q_MX02 U4925 ( .S(xc_mioOn), .A0(evalStepPI[59]), .A1(evalStepPImio[59]), .Z(evalStepPIi[59]));
Q_MX02 U4926 ( .S(xc_mioOn), .A0(evalStepPI[58]), .A1(evalStepPImio[58]), .Z(evalStepPIi[58]));
Q_MX02 U4927 ( .S(xc_mioOn), .A0(evalStepPI[57]), .A1(evalStepPImio[57]), .Z(evalStepPIi[57]));
Q_MX02 U4928 ( .S(xc_mioOn), .A0(evalStepPI[56]), .A1(evalStepPImio[56]), .Z(evalStepPIi[56]));
Q_MX02 U4929 ( .S(xc_mioOn), .A0(evalStepPI[55]), .A1(evalStepPImio[55]), .Z(evalStepPIi[55]));
Q_MX02 U4930 ( .S(xc_mioOn), .A0(evalStepPI[54]), .A1(evalStepPImio[54]), .Z(evalStepPIi[54]));
Q_MX02 U4931 ( .S(xc_mioOn), .A0(evalStepPI[53]), .A1(evalStepPImio[53]), .Z(evalStepPIi[53]));
Q_MX02 U4932 ( .S(xc_mioOn), .A0(evalStepPI[52]), .A1(evalStepPImio[52]), .Z(evalStepPIi[52]));
Q_MX02 U4933 ( .S(xc_mioOn), .A0(evalStepPI[51]), .A1(evalStepPImio[51]), .Z(evalStepPIi[51]));
Q_MX02 U4934 ( .S(xc_mioOn), .A0(evalStepPI[50]), .A1(evalStepPImio[50]), .Z(evalStepPIi[50]));
Q_MX02 U4935 ( .S(xc_mioOn), .A0(evalStepPI[49]), .A1(evalStepPImio[49]), .Z(evalStepPIi[49]));
Q_MX02 U4936 ( .S(xc_mioOn), .A0(evalStepPI[48]), .A1(evalStepPImio[48]), .Z(evalStepPIi[48]));
Q_MX02 U4937 ( .S(xc_mioOn), .A0(evalStepPI[47]), .A1(evalStepPImio[47]), .Z(evalStepPIi[47]));
Q_MX02 U4938 ( .S(xc_mioOn), .A0(evalStepPI[46]), .A1(evalStepPImio[46]), .Z(evalStepPIi[46]));
Q_MX02 U4939 ( .S(xc_mioOn), .A0(evalStepPI[45]), .A1(evalStepPImio[45]), .Z(evalStepPIi[45]));
Q_MX02 U4940 ( .S(xc_mioOn), .A0(evalStepPI[44]), .A1(evalStepPImio[44]), .Z(evalStepPIi[44]));
Q_MX02 U4941 ( .S(xc_mioOn), .A0(evalStepPI[43]), .A1(evalStepPImio[43]), .Z(evalStepPIi[43]));
Q_MX02 U4942 ( .S(xc_mioOn), .A0(evalStepPI[42]), .A1(evalStepPImio[42]), .Z(evalStepPIi[42]));
Q_MX02 U4943 ( .S(xc_mioOn), .A0(evalStepPI[41]), .A1(evalStepPImio[41]), .Z(evalStepPIi[41]));
Q_MX02 U4944 ( .S(xc_mioOn), .A0(evalStepPI[40]), .A1(evalStepPImio[40]), .Z(evalStepPIi[40]));
Q_MX02 U4945 ( .S(xc_mioOn), .A0(evalStepPI[39]), .A1(evalStepPImio[39]), .Z(evalStepPIi[39]));
Q_MX02 U4946 ( .S(xc_mioOn), .A0(evalStepPI[38]), .A1(evalStepPImio[38]), .Z(evalStepPIi[38]));
Q_MX02 U4947 ( .S(xc_mioOn), .A0(evalStepPI[37]), .A1(evalStepPImio[37]), .Z(evalStepPIi[37]));
Q_MX02 U4948 ( .S(xc_mioOn), .A0(evalStepPI[36]), .A1(evalStepPImio[36]), .Z(evalStepPIi[36]));
Q_MX02 U4949 ( .S(xc_mioOn), .A0(evalStepPI[35]), .A1(evalStepPImio[35]), .Z(evalStepPIi[35]));
Q_MX02 U4950 ( .S(xc_mioOn), .A0(evalStepPI[34]), .A1(evalStepPImio[34]), .Z(evalStepPIi[34]));
Q_MX02 U4951 ( .S(xc_mioOn), .A0(evalStepPI[33]), .A1(evalStepPImio[33]), .Z(evalStepPIi[33]));
Q_MX02 U4952 ( .S(xc_mioOn), .A0(evalStepPI[32]), .A1(evalStepPImio[32]), .Z(evalStepPIi[32]));
Q_MX02 U4953 ( .S(xc_mioOn), .A0(evalStepPI[31]), .A1(evalStepPImio[31]), .Z(evalStepPIi[31]));
Q_MX02 U4954 ( .S(xc_mioOn), .A0(evalStepPI[30]), .A1(evalStepPImio[30]), .Z(evalStepPIi[30]));
Q_MX02 U4955 ( .S(xc_mioOn), .A0(evalStepPI[29]), .A1(evalStepPImio[29]), .Z(evalStepPIi[29]));
Q_MX02 U4956 ( .S(xc_mioOn), .A0(evalStepPI[28]), .A1(evalStepPImio[28]), .Z(evalStepPIi[28]));
Q_MX02 U4957 ( .S(xc_mioOn), .A0(evalStepPI[27]), .A1(evalStepPImio[27]), .Z(evalStepPIi[27]));
Q_MX02 U4958 ( .S(xc_mioOn), .A0(evalStepPI[26]), .A1(evalStepPImio[26]), .Z(evalStepPIi[26]));
Q_MX02 U4959 ( .S(xc_mioOn), .A0(evalStepPI[25]), .A1(evalStepPImio[25]), .Z(evalStepPIi[25]));
Q_MX02 U4960 ( .S(xc_mioOn), .A0(evalStepPI[24]), .A1(evalStepPImio[24]), .Z(evalStepPIi[24]));
Q_MX02 U4961 ( .S(xc_mioOn), .A0(evalStepPI[23]), .A1(evalStepPImio[23]), .Z(evalStepPIi[23]));
Q_MX02 U4962 ( .S(xc_mioOn), .A0(evalStepPI[22]), .A1(evalStepPImio[22]), .Z(evalStepPIi[22]));
Q_MX02 U4963 ( .S(xc_mioOn), .A0(evalStepPI[21]), .A1(evalStepPImio[21]), .Z(evalStepPIi[21]));
Q_MX02 U4964 ( .S(xc_mioOn), .A0(evalStepPI[20]), .A1(evalStepPImio[20]), .Z(evalStepPIi[20]));
Q_MX02 U4965 ( .S(xc_mioOn), .A0(evalStepPI[19]), .A1(evalStepPImio[19]), .Z(evalStepPIi[19]));
Q_MX02 U4966 ( .S(xc_mioOn), .A0(evalStepPI[18]), .A1(evalStepPImio[18]), .Z(evalStepPIi[18]));
Q_MX02 U4967 ( .S(xc_mioOn), .A0(evalStepPI[17]), .A1(evalStepPImio[17]), .Z(evalStepPIi[17]));
Q_MX02 U4968 ( .S(xc_mioOn), .A0(evalStepPI[16]), .A1(evalStepPImio[16]), .Z(evalStepPIi[16]));
Q_MX02 U4969 ( .S(xc_mioOn), .A0(evalStepPI[15]), .A1(evalStepPImio[15]), .Z(evalStepPIi[15]));
Q_MX02 U4970 ( .S(xc_mioOn), .A0(evalStepPI[14]), .A1(evalStepPImio[14]), .Z(evalStepPIi[14]));
Q_MX02 U4971 ( .S(xc_mioOn), .A0(evalStepPI[13]), .A1(evalStepPImio[13]), .Z(evalStepPIi[13]));
Q_MX02 U4972 ( .S(xc_mioOn), .A0(evalStepPI[12]), .A1(evalStepPImio[12]), .Z(evalStepPIi[12]));
Q_MX02 U4973 ( .S(xc_mioOn), .A0(evalStepPI[11]), .A1(evalStepPImio[11]), .Z(evalStepPIi[11]));
Q_MX02 U4974 ( .S(xc_mioOn), .A0(evalStepPI[10]), .A1(evalStepPImio[10]), .Z(evalStepPIi[10]));
Q_MX02 U4975 ( .S(xc_mioOn), .A0(evalStepPI[9]), .A1(evalStepPImio[9]), .Z(evalStepPIi[9]));
Q_MX02 U4976 ( .S(xc_mioOn), .A0(evalStepPI[8]), .A1(evalStepPImio[8]), .Z(evalStepPIi[8]));
Q_MX02 U4977 ( .S(xc_mioOn), .A0(evalStepPI[7]), .A1(evalStepPImio[7]), .Z(evalStepPIi[7]));
Q_MX02 U4978 ( .S(xc_mioOn), .A0(evalStepPI[6]), .A1(evalStepPImio[6]), .Z(evalStepPIi[6]));
Q_MX02 U4979 ( .S(xc_mioOn), .A0(evalStepPI[5]), .A1(evalStepPImio[5]), .Z(evalStepPIi[5]));
Q_MX02 U4980 ( .S(xc_mioOn), .A0(evalStepPI[4]), .A1(evalStepPImio[4]), .Z(evalStepPIi[4]));
Q_MX02 U4981 ( .S(xc_mioOn), .A0(evalStepPI[3]), .A1(evalStepPImio[3]), .Z(evalStepPIi[3]));
Q_MX02 U4982 ( .S(xc_mioOn), .A0(evalStepPI[2]), .A1(evalStepPImio[2]), .Z(evalStepPIi[2]));
Q_MX02 U4983 ( .S(xc_mioOn), .A0(evalStepPI[1]), .A1(evalStepPImio[1]), .Z(evalStepPIi[1]));
Q_MX02 U4984 ( .S(xc_mioOn), .A0(evalStepPI[0]), .A1(evalStepPImio[0]), .Z(evalStepPIi[0]));
Q_OR02 U4985 ( .A0(hssReset), .A1(hotSwapOnPI), .Z(GFReset));
Q_RDN U4986 ( .Z(ixcHoldClk));
Q_RDN U4987 ( .Z(ptxBusy));
Q_INV U4988 ( .A(maxBpCycle[15]), .Z(n4178));
Q_AN02 U4989 ( .A0(bHaltCnt[15]), .A1(n4178), .Z(n4177));
Q_OR02 U4990 ( .A0(bHaltCnt[15]), .A1(n4178), .Z(n4176));
Q_INV U4991 ( .A(maxBpCycle[14]), .Z(n4175));
Q_AN03 U4992 ( .A0(bHaltCnt[14]), .A1(n4175), .A2(n4176), .Z(n4167));
Q_OA21 U4993 ( .A0(bHaltCnt[14]), .A1(n4175), .B0(n4176), .Z(n4171));
Q_INV U4994 ( .A(maxBpCycle[13]), .Z(n4174));
Q_AN02 U4995 ( .A0(bHaltCnt[13]), .A1(n4174), .Z(n4173));
Q_OA21 U4996 ( .A0(bHaltCnt[13]), .A1(n4174), .B0(n4171), .Z(n4170));
Q_INV U4997 ( .A(maxBpCycle[12]), .Z(n4172));
Q_AN03 U4998 ( .A0(bHaltCnt[12]), .A1(n4172), .A2(n4170), .Z(n4169));
Q_OA21 U4999 ( .A0(bHaltCnt[12]), .A1(n4172), .B0(n4170), .Z(n4165));
Q_AO21 U5000 ( .A0(n4171), .A1(n4173), .B0(n4169), .Z(n4168));
Q_OR03 U5001 ( .A0(n4177), .A1(n4167), .A2(n4168), .Z(n4166));
Q_INV U5002 ( .A(maxBpCycle[11]), .Z(n4164));
Q_AN02 U5003 ( .A0(bHaltCnt[11]), .A1(n4164), .Z(n4163));
Q_OR02 U5004 ( .A0(bHaltCnt[11]), .A1(n4164), .Z(n4162));
Q_INV U5005 ( .A(maxBpCycle[10]), .Z(n4161));
Q_AN02 U5006 ( .A0(bHaltCnt[10]), .A1(n4161), .Z(n4160));
Q_OA21 U5007 ( .A0(bHaltCnt[10]), .A1(n4161), .B0(n4162), .Z(n4155));
Q_INV U5008 ( .A(maxBpCycle[9]), .Z(n4159));
Q_AN02 U5009 ( .A0(bHaltCnt[9]), .A1(n4159), .Z(n4158));
Q_OA21 U5010 ( .A0(bHaltCnt[9]), .A1(n4159), .B0(n4155), .Z(n4154));
Q_INV U5011 ( .A(maxBpCycle[8]), .Z(n4157));
Q_AN03 U5012 ( .A0(bHaltCnt[8]), .A1(n4157), .A2(n4154), .Z(n4153));
Q_OR02 U5013 ( .A0(bHaltCnt[8]), .A1(n4157), .Z(n4156));
Q_AO21 U5014 ( .A0(n4155), .A1(n4158), .B0(n4153), .Z(n4152));
Q_AO21 U5015 ( .A0(n4162), .A1(n4160), .B0(n4163), .Z(n4151));
Q_OA21 U5016 ( .A0(n4151), .A1(n4152), .B0(n4165), .Z(n4119));
Q_AN03 U5017 ( .A0(n4154), .A1(n4156), .A2(n4165), .Z(n4122));
Q_INV U5018 ( .A(maxBpCycle[7]), .Z(n4150));
Q_AN02 U5019 ( .A0(bHaltCnt[7]), .A1(n4150), .Z(n4149));
Q_OR02 U5020 ( .A0(bHaltCnt[7]), .A1(n4150), .Z(n4148));
Q_INV U5021 ( .A(maxBpCycle[6]), .Z(n4147));
Q_AN03 U5022 ( .A0(bHaltCnt[6]), .A1(n4147), .A2(n4148), .Z(n4139));
Q_OA21 U5023 ( .A0(bHaltCnt[6]), .A1(n4147), .B0(n4148), .Z(n4143));
Q_INV U5024 ( .A(maxBpCycle[5]), .Z(n4146));
Q_AN02 U5025 ( .A0(bHaltCnt[5]), .A1(n4146), .Z(n4145));
Q_OA21 U5026 ( .A0(bHaltCnt[5]), .A1(n4146), .B0(n4143), .Z(n4142));
Q_INV U5027 ( .A(maxBpCycle[4]), .Z(n4144));
Q_AN03 U5028 ( .A0(bHaltCnt[4]), .A1(n4144), .A2(n4142), .Z(n4141));
Q_OA21 U5029 ( .A0(bHaltCnt[4]), .A1(n4144), .B0(n4142), .Z(n4137));
Q_AO21 U5030 ( .A0(n4143), .A1(n4145), .B0(n4141), .Z(n4140));
Q_OR03 U5031 ( .A0(n4149), .A1(n4139), .A2(n4140), .Z(n4138));
Q_INV U5032 ( .A(maxBpCycle[3]), .Z(n4136));
Q_AN02 U5033 ( .A0(bHaltCnt[3]), .A1(n4136), .Z(n4135));
Q_OR02 U5034 ( .A0(bHaltCnt[3]), .A1(n4136), .Z(n4134));
Q_INV U5035 ( .A(maxBpCycle[2]), .Z(n4133));
Q_AN03 U5036 ( .A0(bHaltCnt[2]), .A1(n4133), .A2(n4134), .Z(n4124));
Q_OA21 U5037 ( .A0(bHaltCnt[2]), .A1(n4133), .B0(n4134), .Z(n4127));
Q_INV U5038 ( .A(maxBpCycle[1]), .Z(n4132));
Q_AN02 U5039 ( .A0(bHaltCnt[1]), .A1(n4132), .Z(n4131));
Q_OR02 U5040 ( .A0(bHaltCnt[1]), .A1(n4132), .Z(n4130));
Q_INV U5041 ( .A(maxBpCycle[0]), .Z(n4129));
Q_AN02 U5042 ( .A0(bHaltCnt[0]), .A1(n4129), .Z(n4128));
Q_AN03 U5043 ( .A0(n4127), .A1(n4130), .A2(n4128), .Z(n4126));
Q_AO21 U5044 ( .A0(n4127), .A1(n4131), .B0(n4126), .Z(n4125));
Q_OR03 U5045 ( .A0(n4135), .A1(n4124), .A2(n4125), .Z(n4123));
Q_AN03 U5046 ( .A0(n4122), .A1(n4137), .A2(n4123), .Z(n4121));
Q_AO21 U5047 ( .A0(n4122), .A1(n4138), .B0(n4121), .Z(n4120));
Q_OR03 U5048 ( .A0(n4166), .A1(n4119), .A2(n4120), .Z(n4118));
Q_OR03 U5049 ( .A0(maxBpCycle[15]), .A1(maxBpCycle[14]), .A2(maxBpCycle[13]), .Z(n4117));
Q_OR03 U5050 ( .A0(maxBpCycle[12]), .A1(maxBpCycle[11]), .A2(maxBpCycle[10]), .Z(n4116));
Q_OR03 U5051 ( .A0(maxBpCycle[9]), .A1(maxBpCycle[8]), .A2(maxBpCycle[7]), .Z(n4115));
Q_OR03 U5052 ( .A0(maxBpCycle[6]), .A1(maxBpCycle[5]), .A2(maxBpCycle[4]), .Z(n4114));
Q_OR03 U5053 ( .A0(maxBpCycle[3]), .A1(maxBpCycle[2]), .A2(maxBpCycle[1]), .Z(n4113));
Q_OR03 U5054 ( .A0(maxBpCycle[0]), .A1(n4117), .A2(n4116), .Z(n4112));
Q_OR03 U5055 ( .A0(n4115), .A1(n4114), .A2(n4113), .Z(n4111));
Q_OA21 U5056 ( .A0(n4112), .A1(n4111), .B0(n4118), .Z(bpHalt));
Q_INV U5057 ( .A(maxAcCycle[15]), .Z(n4110));
Q_AN02 U5058 ( .A0(aHaltCnt[15]), .A1(n4110), .Z(n4109));
Q_OR02 U5059 ( .A0(aHaltCnt[15]), .A1(n4110), .Z(n4108));
Q_INV U5060 ( .A(maxAcCycle[14]), .Z(n4107));
Q_AN03 U5061 ( .A0(aHaltCnt[14]), .A1(n4107), .A2(n4108), .Z(n4099));
Q_OA21 U5062 ( .A0(aHaltCnt[14]), .A1(n4107), .B0(n4108), .Z(n4103));
Q_INV U5063 ( .A(maxAcCycle[13]), .Z(n4106));
Q_AN02 U5064 ( .A0(aHaltCnt[13]), .A1(n4106), .Z(n4105));
Q_OA21 U5065 ( .A0(aHaltCnt[13]), .A1(n4106), .B0(n4103), .Z(n4102));
Q_INV U5066 ( .A(maxAcCycle[12]), .Z(n4104));
Q_AN03 U5067 ( .A0(aHaltCnt[12]), .A1(n4104), .A2(n4102), .Z(n4101));
Q_OA21 U5068 ( .A0(aHaltCnt[12]), .A1(n4104), .B0(n4102), .Z(n4097));
Q_AO21 U5069 ( .A0(n4103), .A1(n4105), .B0(n4101), .Z(n4100));
Q_OR03 U5070 ( .A0(n4109), .A1(n4099), .A2(n4100), .Z(n4098));
Q_INV U5071 ( .A(maxAcCycle[11]), .Z(n4096));
Q_AN02 U5072 ( .A0(aHaltCnt[11]), .A1(n4096), .Z(n4095));
Q_OR02 U5073 ( .A0(aHaltCnt[11]), .A1(n4096), .Z(n4094));
Q_INV U5074 ( .A(maxAcCycle[10]), .Z(n4093));
Q_AN02 U5075 ( .A0(aHaltCnt[10]), .A1(n4093), .Z(n4092));
Q_OA21 U5076 ( .A0(aHaltCnt[10]), .A1(n4093), .B0(n4094), .Z(n4087));
Q_INV U5077 ( .A(maxAcCycle[9]), .Z(n4091));
Q_AN02 U5078 ( .A0(aHaltCnt[9]), .A1(n4091), .Z(n4090));
Q_OA21 U5079 ( .A0(aHaltCnt[9]), .A1(n4091), .B0(n4087), .Z(n4086));
Q_INV U5080 ( .A(maxAcCycle[8]), .Z(n4089));
Q_AN03 U5081 ( .A0(aHaltCnt[8]), .A1(n4089), .A2(n4086), .Z(n4085));
Q_OR02 U5082 ( .A0(aHaltCnt[8]), .A1(n4089), .Z(n4088));
Q_AO21 U5083 ( .A0(n4087), .A1(n4090), .B0(n4085), .Z(n4084));
Q_AO21 U5084 ( .A0(n4094), .A1(n4092), .B0(n4095), .Z(n4083));
Q_OA21 U5085 ( .A0(n4083), .A1(n4084), .B0(n4097), .Z(n4051));
Q_AN03 U5086 ( .A0(n4086), .A1(n4088), .A2(n4097), .Z(n4054));
Q_INV U5087 ( .A(maxAcCycle[7]), .Z(n4082));
Q_AN02 U5088 ( .A0(aHaltCnt[7]), .A1(n4082), .Z(n4081));
Q_OR02 U5089 ( .A0(aHaltCnt[7]), .A1(n4082), .Z(n4080));
Q_INV U5090 ( .A(maxAcCycle[6]), .Z(n4079));
Q_AN03 U5091 ( .A0(aHaltCnt[6]), .A1(n4079), .A2(n4080), .Z(n4071));
Q_OA21 U5092 ( .A0(aHaltCnt[6]), .A1(n4079), .B0(n4080), .Z(n4075));
Q_INV U5093 ( .A(maxAcCycle[5]), .Z(n4078));
Q_AN02 U5094 ( .A0(aHaltCnt[5]), .A1(n4078), .Z(n4077));
Q_OA21 U5095 ( .A0(aHaltCnt[5]), .A1(n4078), .B0(n4075), .Z(n4074));
Q_INV U5096 ( .A(maxAcCycle[4]), .Z(n4076));
Q_AN03 U5097 ( .A0(aHaltCnt[4]), .A1(n4076), .A2(n4074), .Z(n4073));
Q_OA21 U5098 ( .A0(aHaltCnt[4]), .A1(n4076), .B0(n4074), .Z(n4069));
Q_AO21 U5099 ( .A0(n4075), .A1(n4077), .B0(n4073), .Z(n4072));
Q_OR03 U5100 ( .A0(n4081), .A1(n4071), .A2(n4072), .Z(n4070));
Q_INV U5101 ( .A(maxAcCycle[3]), .Z(n4068));
Q_AN02 U5102 ( .A0(aHaltCnt[3]), .A1(n4068), .Z(n4067));
Q_OR02 U5103 ( .A0(aHaltCnt[3]), .A1(n4068), .Z(n4066));
Q_INV U5104 ( .A(maxAcCycle[2]), .Z(n4065));
Q_AN03 U5105 ( .A0(aHaltCnt[2]), .A1(n4065), .A2(n4066), .Z(n4056));
Q_OA21 U5106 ( .A0(aHaltCnt[2]), .A1(n4065), .B0(n4066), .Z(n4059));
Q_INV U5107 ( .A(maxAcCycle[1]), .Z(n4064));
Q_AN02 U5108 ( .A0(aHaltCnt[1]), .A1(n4064), .Z(n4063));
Q_OR02 U5109 ( .A0(aHaltCnt[1]), .A1(n4064), .Z(n4062));
Q_INV U5110 ( .A(maxAcCycle[0]), .Z(n4061));
Q_AN02 U5111 ( .A0(aHaltCnt[0]), .A1(n4061), .Z(n4060));
Q_AN03 U5112 ( .A0(n4059), .A1(n4062), .A2(n4060), .Z(n4058));
Q_AO21 U5113 ( .A0(n4059), .A1(n4063), .B0(n4058), .Z(n4057));
Q_OR03 U5114 ( .A0(n4067), .A1(n4056), .A2(n4057), .Z(n4055));
Q_AN03 U5115 ( .A0(n4054), .A1(n4069), .A2(n4055), .Z(n4053));
Q_AO21 U5116 ( .A0(n4054), .A1(n4070), .B0(n4053), .Z(n4052));
Q_OR03 U5117 ( .A0(n4098), .A1(n4051), .A2(n4052), .Z(n4050));
Q_OR03 U5118 ( .A0(maxAcCycle[15]), .A1(maxAcCycle[14]), .A2(maxAcCycle[13]), .Z(n4049));
Q_OR03 U5119 ( .A0(maxAcCycle[12]), .A1(maxAcCycle[11]), .A2(maxAcCycle[10]), .Z(n4048));
Q_OR03 U5120 ( .A0(maxAcCycle[9]), .A1(maxAcCycle[8]), .A2(maxAcCycle[7]), .Z(n4047));
Q_OR03 U5121 ( .A0(maxAcCycle[6]), .A1(maxAcCycle[5]), .A2(maxAcCycle[4]), .Z(n4046));
Q_OR03 U5122 ( .A0(maxAcCycle[3]), .A1(maxAcCycle[2]), .A2(maxAcCycle[1]), .Z(n4045));
Q_OR03 U5123 ( .A0(maxAcCycle[0]), .A1(n4049), .A2(n4048), .Z(n4044));
Q_OR03 U5124 ( .A0(n4047), .A1(n4046), .A2(n4045), .Z(n4043));
Q_OA21 U5125 ( .A0(n4044), .A1(n4043), .B0(n4050), .Z(acHalt));
Q_XOR2 U5126 ( .A0(callEmuPIi), .A1(callEmuR), .Z(callEmuEv));
Q_OR02 U5127 ( .A0(lbrOn), .A1(hotSwapOnPI), .Z(lbrOnAll));
Q_INV U5128 ( .A(gfifoAsyncOff), .Z(n4042));
Q_AN02 U5129 ( .A0(GFGBfull), .A1(n4042), .Z(GFGBfullBw));
Q_RDN U5130 ( .Z(GFAck));
Q_OR02 U5131 ( .A0(bClkR), .A1(bpHalt), .Z(bClkRH));
Q_OR03 U5132 ( .A0(n628), .A1(n642), .A2(n641), .Z(n4041));
Q_OR02 U5133 ( .A0(n4041), .A1(n636), .Z(n4040));
Q_OR03 U5134 ( .A0(n598), .A1(n635), .A2(n634), .Z(n4039));
Q_OR02 U5135 ( .A0(n4039), .A1(n629), .Z(n4038));
Q_ND02 U5136 ( .A0(n4040), .A1(n4038), .Z(syncEn));
Q_RDN U5137 ( .Z(svGFbusy));
Q_RDN U5138 ( .Z(otbGFbusy));
Q_RDN U5139 ( .Z(svAsyncCall));
Q_RDN U5140 ( .Z(otbAsyncCall));
Q_RDN U5141 ( .Z(ecmHoldBusy));
Q_EV_WOR qstp1 ( .A(stop1));
Q_EV_WOR qstp2 ( .A(stop2));
Q_EV_WOR qstp4 ( .A(stop4));
Q_RDN U5145 ( .Z(stop1));
Q_RDN U5146 ( .Z(stop2));
Q_RDN U5147 ( .Z(stop4));
Q_AO21 U5148 ( .A0(otbGFbusy), .A1(hasGFIFO1), .B0(svGFbusy), .Z(GFbusy));
Q_AO21 U5149 ( .A0(otbAsyncCall), .A1(syncOtbChannels), .B0(svAsyncCall), .Z(asyncCall));
Q_RDN U5150 ( .Z(isfWait));
Q_RDN U5151 ( .Z(osfWait));
Q_OR03 U5152 ( .A0(fclkPerEval[7]), .A1(fclkPerEval[6]), .A2(fclkPerEval[5]), .Z(n4037));
Q_OR03 U5153 ( .A0(fclkPerEval[4]), .A1(fclkPerEval[3]), .A2(fclkPerEval[2]), .Z(n4036));
Q_OR03 U5154 ( .A0(fclkPerEval[1]), .A1(fclkPerEval[0]), .A2(n4037), .Z(n4035));
Q_NR02 U5155 ( .A0(n4036), .A1(n4035), .Z(oneFclkEval));
Q_AN02 U5156 ( .A0(ixc_time.runClk), .A1(simTimeEnable), .Z(cakeCcEnable));
Q_PULSE U5157 ( .A(eClkR), .Z(eClk));
Q_BUF U5158 ( .A(_ET3_COMPILER_RESERVED_NAME_DBI_APPLY_), .Z(APPLY_PI));
Q_BUF U5159 ( .A(lbrOnAll), .Z(_ET3_COMPILER_RESERVED_NAME_LBRKER_ON_));
Q_RDN U5160 ( .Z(GFLBfull));
Q_RDN U5161 ( .Z(GFGBfull));
Q_RDN U5162 ( .Z(GFBw));
Q_EV_WOR_START gbf ( .A(GFGBfullBw));
Q_OA21 U5164 ( .A0(gfifoOff), .A1(hotSwapOnPI), .B0(n3045), .Z(GFLock1));
Q_OR03 U5165 ( .A0(GFbusy), .A1(GFbusyD), .A2(GFbusyD2), .Z(gfifoWait));
Q_RDN U5166 ( .Z(bpWait));
Q_RDN U5167 ( .Z(bWait));
Q_RDN U5168 ( .Z(eClkHold));
Q_RDN U5169 ( .Z(sampleXpChg));
Q_EV_WOR qbwi ( .A(bpWait));
Q_EV_WOR qxci ( .A(sampleXpChg));
Q_PULSE U5172 ( .A(bClkRH), .Z(bClk));
Q_OR03 U5173 ( .A0(bWait), .A1(bWaitExtend), .A2(holdEcmC), .Z(n4034));
Q_OR03 U5174 ( .A0(bClkHoldD), .A1(ixcHoldClk), .A2(GFBw), .Z(n4033));
Q_OR02 U5175 ( .A0(n4034), .A1(n4033), .Z(xpHold));
Q_EV_WOR_START bkh ( .A(bClkHoldD));
Q_EV_WOR_START hec ( .A(holdEcmC));
Q_BUF intrBuf ( .A(intr), .Z(_ET3_COMPILER_RESERVED_NAME_ORION_INTERRUPT_));
Q_OA21 U5179 ( .A0(it_capture), .A1(it_replay), .B0(it_endBuf), .Z(it_newBuf));
Q_RBUFZN  dum1 ( dummyW, n4032, n4031);
Q_RBUFZP  dum2 ( dummyW, n4030, n1);
Q_OR03 U5182 ( .A0(mioPOW_2[4]), .A1(stopTL), .A2(mioPOW_2[5]), .Z(n4028));
Q_OR03 U5183 ( .A0(mioPOW_2[3]), .A1(mioPOW_2[2]), .A2(n4028), .Z(anyStop));
Q_EV_WOR_START qsynci ( .A(syncEn));
Q_OR02 U5185 ( .A0(callEmuPre), .A1(simTimeEnable), .Z(ecmOn));
Q_OR03 U5186 ( .A0(svAsyncCall), .A1(otbAsyncCall), .A2(ptxBusy), .Z(ecmNotSync));
Q_RDN U5187 ( .Z(holdEcmTb));
Q_RDN U5188 ( .Z(ptxHoldEcm));
Q_OR03 U5189 ( .A0(holdEcmTb), .A1(holdEcmPtxOn), .A2(holdEcmSync), .Z(holdEcm));
Q_PULSE U5190 ( .A(clockMC), .Z(mcp));
Q_XNR2 U5191 ( .A0(ixc_time.nextDutTime[0]), .A1(n4027), .Z(mcDelta[0]));
Q_OR02 U5192 ( .A0(ixc_time.nextDutTime[0]), .A1(n4027), .Z(n3996));
Q_AD02 U5193 ( .CI(n3996), .A0(ixc_time.nextDutTime[1]), .A1(ixc_time.nextDutTime[2]), .B0(n4026), .B1(n4025), .S0(mcDelta[1]), .S1(mcDelta[2]), .CO(n3995));
Q_AD02 U5194 ( .CI(n3995), .A0(ixc_time.nextDutTime[3]), .A1(ixc_time.nextDutTime[4]), .B0(n4024), .B1(n4023), .S0(mcDelta[3]), .S1(mcDelta[4]), .CO(n3994));
Q_AD02 U5195 ( .CI(n3994), .A0(ixc_time.nextDutTime[5]), .A1(ixc_time.nextDutTime[6]), .B0(n4022), .B1(n4021), .S0(mcDelta[5]), .S1(mcDelta[6]), .CO(n3993));
Q_AD02 U5196 ( .CI(n3993), .A0(ixc_time.nextDutTime[7]), .A1(ixc_time.nextDutTime[8]), .B0(n4020), .B1(n4019), .S0(mcDelta[7]), .S1(mcDelta[8]), .CO(n3992));
Q_AD02 U5197 ( .CI(n3992), .A0(ixc_time.nextDutTime[9]), .A1(ixc_time.nextDutTime[10]), .B0(n4018), .B1(n4017), .S0(mcDelta[9]), .S1(mcDelta[10]), .CO(n3991));
Q_AD02 U5198 ( .CI(n3991), .A0(ixc_time.nextDutTime[11]), .A1(ixc_time.nextDutTime[12]), .B0(n4016), .B1(n4015), .S0(mcDelta[11]), .S1(mcDelta[12]), .CO(n3990));
Q_AD02 U5199 ( .CI(n3990), .A0(ixc_time.nextDutTime[13]), .A1(ixc_time.nextDutTime[14]), .B0(n4014), .B1(n4013), .S0(mcDelta[13]), .S1(mcDelta[14]), .CO(n3989));
Q_AD02 U5200 ( .CI(n3989), .A0(ixc_time.nextDutTime[15]), .A1(ixc_time.nextDutTime[16]), .B0(n4012), .B1(n4011), .S0(mcDelta[15]), .S1(mcDelta[16]), .CO(n3988));
Q_AD02 U5201 ( .CI(n3988), .A0(ixc_time.nextDutTime[17]), .A1(ixc_time.nextDutTime[18]), .B0(n4010), .B1(n4009), .S0(mcDelta[17]), .S1(mcDelta[18]), .CO(n3987));
Q_AD02 U5202 ( .CI(n3987), .A0(ixc_time.nextDutTime[19]), .A1(ixc_time.nextDutTime[20]), .B0(n4008), .B1(n4007), .S0(mcDelta[19]), .S1(mcDelta[20]), .CO(n3986));
Q_AD02 U5203 ( .CI(n3986), .A0(ixc_time.nextDutTime[21]), .A1(ixc_time.nextDutTime[22]), .B0(n4006), .B1(n4005), .S0(mcDelta[21]), .S1(mcDelta[22]), .CO(n3985));
Q_AD02 U5204 ( .CI(n3985), .A0(ixc_time.nextDutTime[23]), .A1(ixc_time.nextDutTime[24]), .B0(n4004), .B1(n4003), .S0(mcDelta[23]), .S1(mcDelta[24]), .CO(n3984));
Q_AD02 U5205 ( .CI(n3984), .A0(ixc_time.nextDutTime[25]), .A1(ixc_time.nextDutTime[26]), .B0(n4002), .B1(n4001), .S0(mcDelta[25]), .S1(mcDelta[26]), .CO(n3983));
Q_AD02 U5206 ( .CI(n3983), .A0(ixc_time.nextDutTime[27]), .A1(ixc_time.nextDutTime[28]), .B0(n4000), .B1(n3999), .S0(mcDelta[27]), .S1(mcDelta[28]), .CO(n3982));
Q_AD02 U5207 ( .CI(n3982), .A0(ixc_time.nextDutTime[29]), .A1(ixc_time.nextDutTime[30]), .B0(n3998), .B1(n3997), .S0(mcDelta[29]), .S1(mcDelta[30]), .CO(n3981));
Q_PULSE U5208 ( .A(uClkT), .Z(uClk));
Q_NOT_TOUCH _zzqnthw ( .sig());
Q_INV U5210 ( .A(xpHold), .Z(n3980));
Q_AN02 U5211 ( .A0(lastDelta), .A1(n3980), .Z(mpEnable));
Q_EV_WOR qxhi ( .A(xpHold));
Q_OR02 U5213 ( .A0(ecmNotSync), .A1(ecmNotSyncD), .Z(n3979));
Q_INV U5214 ( .A(n3979), .Z(ecmSync));
Q_INV U5215 ( .A(n2917), .Z(sampleXpV));
Q_INV U5216 ( .A(eCount[63]), .Z(n5489));
Q_FDP4EP \eCount_REG[63] ( .CK(eClk), .CE(n3809), .R(n4029), .D(n5489), .Q(eCount[63]));
Q_INV U5218 ( .A(bpCount[63]), .Z(n5490));
Q_FDP4EP \bpCount_REG[63] ( .CK(bClk), .CE(n3684), .R(n4029), .D(n5490), .Q(bpCount[63]));
Q_INV U5220 ( .A(uClkCntr[0]), .Z(n5491));
Q_FDP4EP \uClkCntr_REG[0] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n5491), .Q(uClkCntr[0]));
Q_FDP4EP \uClkCntr_REG[1] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3428), .Q(uClkCntr[1]));
Q_FDP4EP \uClkCntr_REG[2] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3430), .Q(uClkCntr[2]));
Q_FDP4EP \uClkCntr_REG[3] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3432), .Q(uClkCntr[3]));
Q_FDP4EP \uClkCntr_REG[4] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3434), .Q(uClkCntr[4]));
Q_FDP4EP \uClkCntr_REG[5] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3436), .Q(uClkCntr[5]));
Q_FDP4EP \uClkCntr_REG[6] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3438), .Q(uClkCntr[6]));
Q_FDP4EP \uClkCntr_REG[7] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3440), .Q(uClkCntr[7]));
Q_FDP4EP \uClkCntr_REG[8] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3442), .Q(uClkCntr[8]));
Q_FDP4EP \uClkCntr_REG[9] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3444), .Q(uClkCntr[9]));
Q_FDP4EP \uClkCntr_REG[10] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3446), .Q(uClkCntr[10]));
Q_FDP4EP \uClkCntr_REG[11] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3448), .Q(uClkCntr[11]));
Q_FDP4EP \uClkCntr_REG[12] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3450), .Q(uClkCntr[12]));
Q_FDP4EP \uClkCntr_REG[13] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3452), .Q(uClkCntr[13]));
Q_FDP4EP \uClkCntr_REG[14] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3454), .Q(uClkCntr[14]));
Q_FDP4EP \uClkCntr_REG[15] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3456), .Q(uClkCntr[15]));
Q_FDP4EP \uClkCntr_REG[16] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3458), .Q(uClkCntr[16]));
Q_FDP4EP \uClkCntr_REG[17] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3460), .Q(uClkCntr[17]));
Q_FDP4EP \uClkCntr_REG[18] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3462), .Q(uClkCntr[18]));
Q_FDP4EP \uClkCntr_REG[19] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3464), .Q(uClkCntr[19]));
Q_FDP4EP \uClkCntr_REG[20] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3466), .Q(uClkCntr[20]));
Q_FDP4EP \uClkCntr_REG[21] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3468), .Q(uClkCntr[21]));
Q_FDP4EP \uClkCntr_REG[22] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3470), .Q(uClkCntr[22]));
Q_FDP4EP \uClkCntr_REG[23] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3472), .Q(uClkCntr[23]));
Q_FDP4EP \uClkCntr_REG[24] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3474), .Q(uClkCntr[24]));
Q_FDP4EP \uClkCntr_REG[25] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3476), .Q(uClkCntr[25]));
Q_FDP4EP \uClkCntr_REG[26] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3478), .Q(uClkCntr[26]));
Q_FDP4EP \uClkCntr_REG[27] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3480), .Q(uClkCntr[27]));
Q_FDP4EP \uClkCntr_REG[28] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3482), .Q(uClkCntr[28]));
Q_FDP4EP \uClkCntr_REG[29] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3484), .Q(uClkCntr[29]));
Q_FDP4EP \uClkCntr_REG[30] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3486), .Q(uClkCntr[30]));
Q_FDP4EP \uClkCntr_REG[31] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3488), .Q(uClkCntr[31]));
Q_FDP4EP \uClkCntr_REG[32] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3490), .Q(uClkCntr[32]));
Q_FDP4EP \uClkCntr_REG[33] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3492), .Q(uClkCntr[33]));
Q_FDP4EP \uClkCntr_REG[34] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3494), .Q(uClkCntr[34]));
Q_FDP4EP \uClkCntr_REG[35] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3496), .Q(uClkCntr[35]));
Q_FDP4EP \uClkCntr_REG[36] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3498), .Q(uClkCntr[36]));
Q_FDP4EP \uClkCntr_REG[37] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3500), .Q(uClkCntr[37]));
Q_FDP4EP \uClkCntr_REG[38] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3502), .Q(uClkCntr[38]));
Q_FDP4EP \uClkCntr_REG[39] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3504), .Q(uClkCntr[39]));
Q_FDP4EP \uClkCntr_REG[40] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3506), .Q(uClkCntr[40]));
Q_FDP4EP \uClkCntr_REG[41] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3508), .Q(uClkCntr[41]));
Q_FDP4EP \uClkCntr_REG[42] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3510), .Q(uClkCntr[42]));
Q_FDP4EP \uClkCntr_REG[43] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3512), .Q(uClkCntr[43]));
Q_FDP4EP \uClkCntr_REG[44] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3514), .Q(uClkCntr[44]));
Q_FDP4EP \uClkCntr_REG[45] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3516), .Q(uClkCntr[45]));
Q_FDP4EP \uClkCntr_REG[46] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3518), .Q(uClkCntr[46]));
Q_FDP4EP \uClkCntr_REG[47] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3520), .Q(uClkCntr[47]));
Q_FDP4EP \uClkCntr_REG[48] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3522), .Q(uClkCntr[48]));
Q_FDP4EP \uClkCntr_REG[49] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3524), .Q(uClkCntr[49]));
Q_FDP4EP \uClkCntr_REG[50] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3526), .Q(uClkCntr[50]));
Q_FDP4EP \uClkCntr_REG[51] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3528), .Q(uClkCntr[51]));
Q_FDP4EP \uClkCntr_REG[52] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3530), .Q(uClkCntr[52]));
Q_FDP4EP \uClkCntr_REG[53] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3532), .Q(uClkCntr[53]));
Q_FDP4EP \uClkCntr_REG[54] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3534), .Q(uClkCntr[54]));
Q_FDP4EP \uClkCntr_REG[55] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3536), .Q(uClkCntr[55]));
Q_FDP4EP \uClkCntr_REG[56] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3538), .Q(uClkCntr[56]));
Q_FDP4EP \uClkCntr_REG[57] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3540), .Q(uClkCntr[57]));
Q_FDP4EP \uClkCntr_REG[58] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3542), .Q(uClkCntr[58]));
Q_FDP4EP \uClkCntr_REG[59] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3544), .Q(uClkCntr[59]));
Q_FDP4EP \uClkCntr_REG[60] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3546), .Q(uClkCntr[60]));
Q_FDP4EP \uClkCntr_REG[61] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3548), .Q(uClkCntr[61]));
Q_FDP4EP \uClkCntr_REG[62] ( .CK(uClk), .CE(initClock), .R(n4029), .D(n3550), .Q(uClkCntr[62]));
Q_INV U5284 ( .A(uClkCntr[63]), .Z(n5492));
Q_FDP4EP \uClkCntr_REG[63] ( .CK(uClk), .CE(n2), .R(n4029), .D(n5492), .Q(uClkCntr[63]));
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE "xc_top"
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE_LIB "IXCOM_TEMP_LIBRARY"
// pragma CVASTRPROP MODULE HDLICE PROP_IXCOM_MOD TRUE
// pragma CVASTRPROP MODULE HDLICE PROP_RANOFF TRUE
endmodule
