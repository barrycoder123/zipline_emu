
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
(* celldefine = 1 *) 
module nx_rbus_apb ( rbus_addr_o, rbus_wr_strb_o, rbus_wr_data_o, 
	rbus_rd_strb_o, apb_prdata, apb_pready, apb_pslverr, clk, rst_n, 
	rbus_rd_data_i, rbus_ack_i, rbus_err_ack_i, rbus_wr_strb_i, 
	rbus_rd_strb_i, apb_paddr, apb_psel, apb_penable, apb_pwrite, 
	apb_pwdata);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output [15:0] rbus_addr_o;
output rbus_wr_strb_o;
output [31:0] rbus_wr_data_o;
output rbus_rd_strb_o;
output [31:0] apb_prdata;
output apb_pready;
output apb_pslverr;
input clk;
input rst_n;
input [31:0] rbus_rd_data_i;
input rbus_ack_i;
input rbus_err_ack_i;
input rbus_wr_strb_i;
input rbus_rd_strb_i;
input [15:0] apb_paddr;
input apb_psel;
input apb_penable;
input apb_pwrite;
input [31:0] apb_pwdata;
wire [0:15] _zy_simnet_rbus_addr_o_0_w$;
wire _zy_simnet_rbus_wr_strb_o_1_w$;
wire [0:31] _zy_simnet_rbus_wr_data_o_2_w$;
wire _zy_simnet_rbus_rd_strb_o_3_w$;
wire [0:31] _zy_simnet_apb_prdata_4_w$;
wire _zy_simnet_apb_pready_5_w$;
wire _zy_simnet_apb_pslverr_6_w$;
wire [15:0] apb_paddr_reg;
wire apb_penable_reg;
wire apb_psel_reg;
wire [31:0] apb_pwdata_reg;
wire apb_pwrite_reg;
wire apb_active;
wire apb_active_reg;
ixc_assign _zz_strnp_6 ( _zy_simnet_apb_pslverr_6_w$, apb_pslverr);
ixc_assign _zz_strnp_5 ( _zy_simnet_apb_pready_5_w$, apb_pready);
ixc_assign_32 _zz_strnp_4 ( _zy_simnet_apb_prdata_4_w$[0:31], 
	apb_prdata[31:0]);
ixc_assign _zz_strnp_3 ( _zy_simnet_rbus_rd_strb_o_3_w$, rbus_rd_strb_o);
ixc_assign_32 _zz_strnp_2 ( _zy_simnet_rbus_wr_data_o_2_w$[0:31], 
	rbus_wr_data_o[31:0]);
ixc_assign _zz_strnp_1 ( _zy_simnet_rbus_wr_strb_o_1_w$, rbus_wr_strb_o);
ixc_assign_16 _zz_strnp_0 ( _zy_simnet_rbus_addr_o_0_w$[0:15], 
	rbus_addr_o[15:0]);
Q_FDP1 \apb_paddr_reg_REG[15] ( .CK(clk), .R(rst_n), .D(apb_paddr[15]), .Q(apb_paddr_reg[15]), .QN( ));
Q_FDP1 \apb_paddr_reg_REG[14] ( .CK(clk), .R(rst_n), .D(apb_paddr[14]), .Q(apb_paddr_reg[14]), .QN( ));
Q_FDP1 \apb_paddr_reg_REG[13] ( .CK(clk), .R(rst_n), .D(apb_paddr[13]), .Q(apb_paddr_reg[13]), .QN( ));
Q_FDP1 \apb_paddr_reg_REG[12] ( .CK(clk), .R(rst_n), .D(apb_paddr[12]), .Q(apb_paddr_reg[12]), .QN( ));
Q_FDP1 \apb_paddr_reg_REG[11] ( .CK(clk), .R(rst_n), .D(apb_paddr[11]), .Q(apb_paddr_reg[11]), .QN( ));
Q_FDP1 \apb_paddr_reg_REG[10] ( .CK(clk), .R(rst_n), .D(apb_paddr[10]), .Q(apb_paddr_reg[10]), .QN( ));
Q_FDP1 \apb_paddr_reg_REG[9] ( .CK(clk), .R(rst_n), .D(apb_paddr[9]), .Q(apb_paddr_reg[9]), .QN( ));
Q_FDP1 \apb_paddr_reg_REG[8] ( .CK(clk), .R(rst_n), .D(apb_paddr[8]), .Q(apb_paddr_reg[8]), .QN( ));
Q_FDP1 \apb_paddr_reg_REG[7] ( .CK(clk), .R(rst_n), .D(apb_paddr[7]), .Q(apb_paddr_reg[7]), .QN( ));
Q_FDP1 \apb_paddr_reg_REG[6] ( .CK(clk), .R(rst_n), .D(apb_paddr[6]), .Q(apb_paddr_reg[6]), .QN( ));
Q_FDP1 \apb_paddr_reg_REG[5] ( .CK(clk), .R(rst_n), .D(apb_paddr[5]), .Q(apb_paddr_reg[5]), .QN( ));
Q_FDP1 \apb_paddr_reg_REG[4] ( .CK(clk), .R(rst_n), .D(apb_paddr[4]), .Q(apb_paddr_reg[4]), .QN( ));
Q_FDP1 \apb_paddr_reg_REG[3] ( .CK(clk), .R(rst_n), .D(apb_paddr[3]), .Q(apb_paddr_reg[3]), .QN( ));
Q_FDP1 \apb_paddr_reg_REG[2] ( .CK(clk), .R(rst_n), .D(apb_paddr[2]), .Q(apb_paddr_reg[2]), .QN( ));
Q_FDP1 \apb_paddr_reg_REG[1] ( .CK(clk), .R(rst_n), .D(apb_paddr[1]), .Q(apb_paddr_reg[1]), .QN( ));
Q_FDP1 \apb_paddr_reg_REG[0] ( .CK(clk), .R(rst_n), .D(apb_paddr[0]), .Q(apb_paddr_reg[0]), .QN( ));
Q_FDP1 apb_penable_reg_REG  ( .CK(clk), .R(rst_n), .D(apb_penable), .Q(apb_penable_reg), .QN( ));
Q_FDP1 apb_psel_reg_REG  ( .CK(clk), .R(rst_n), .D(apb_psel), .Q(apb_psel_reg), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[31] ( .CK(clk), .R(rst_n), .D(apb_pwdata[31]), .Q(apb_pwdata_reg[31]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[30] ( .CK(clk), .R(rst_n), .D(apb_pwdata[30]), .Q(apb_pwdata_reg[30]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[29] ( .CK(clk), .R(rst_n), .D(apb_pwdata[29]), .Q(apb_pwdata_reg[29]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[28] ( .CK(clk), .R(rst_n), .D(apb_pwdata[28]), .Q(apb_pwdata_reg[28]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[27] ( .CK(clk), .R(rst_n), .D(apb_pwdata[27]), .Q(apb_pwdata_reg[27]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[26] ( .CK(clk), .R(rst_n), .D(apb_pwdata[26]), .Q(apb_pwdata_reg[26]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[25] ( .CK(clk), .R(rst_n), .D(apb_pwdata[25]), .Q(apb_pwdata_reg[25]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[24] ( .CK(clk), .R(rst_n), .D(apb_pwdata[24]), .Q(apb_pwdata_reg[24]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[23] ( .CK(clk), .R(rst_n), .D(apb_pwdata[23]), .Q(apb_pwdata_reg[23]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[22] ( .CK(clk), .R(rst_n), .D(apb_pwdata[22]), .Q(apb_pwdata_reg[22]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[21] ( .CK(clk), .R(rst_n), .D(apb_pwdata[21]), .Q(apb_pwdata_reg[21]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[20] ( .CK(clk), .R(rst_n), .D(apb_pwdata[20]), .Q(apb_pwdata_reg[20]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[19] ( .CK(clk), .R(rst_n), .D(apb_pwdata[19]), .Q(apb_pwdata_reg[19]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[18] ( .CK(clk), .R(rst_n), .D(apb_pwdata[18]), .Q(apb_pwdata_reg[18]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[17] ( .CK(clk), .R(rst_n), .D(apb_pwdata[17]), .Q(apb_pwdata_reg[17]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[16] ( .CK(clk), .R(rst_n), .D(apb_pwdata[16]), .Q(apb_pwdata_reg[16]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[15] ( .CK(clk), .R(rst_n), .D(apb_pwdata[15]), .Q(apb_pwdata_reg[15]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[14] ( .CK(clk), .R(rst_n), .D(apb_pwdata[14]), .Q(apb_pwdata_reg[14]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[13] ( .CK(clk), .R(rst_n), .D(apb_pwdata[13]), .Q(apb_pwdata_reg[13]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[12] ( .CK(clk), .R(rst_n), .D(apb_pwdata[12]), .Q(apb_pwdata_reg[12]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[11] ( .CK(clk), .R(rst_n), .D(apb_pwdata[11]), .Q(apb_pwdata_reg[11]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[10] ( .CK(clk), .R(rst_n), .D(apb_pwdata[10]), .Q(apb_pwdata_reg[10]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[9] ( .CK(clk), .R(rst_n), .D(apb_pwdata[9]), .Q(apb_pwdata_reg[9]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[8] ( .CK(clk), .R(rst_n), .D(apb_pwdata[8]), .Q(apb_pwdata_reg[8]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[7] ( .CK(clk), .R(rst_n), .D(apb_pwdata[7]), .Q(apb_pwdata_reg[7]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[6] ( .CK(clk), .R(rst_n), .D(apb_pwdata[6]), .Q(apb_pwdata_reg[6]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[5] ( .CK(clk), .R(rst_n), .D(apb_pwdata[5]), .Q(apb_pwdata_reg[5]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[4] ( .CK(clk), .R(rst_n), .D(apb_pwdata[4]), .Q(apb_pwdata_reg[4]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[3] ( .CK(clk), .R(rst_n), .D(apb_pwdata[3]), .Q(apb_pwdata_reg[3]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[2] ( .CK(clk), .R(rst_n), .D(apb_pwdata[2]), .Q(apb_pwdata_reg[2]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[1] ( .CK(clk), .R(rst_n), .D(apb_pwdata[1]), .Q(apb_pwdata_reg[1]), .QN( ));
Q_FDP1 \apb_pwdata_reg_REG[0] ( .CK(clk), .R(rst_n), .D(apb_pwdata[0]), .Q(apb_pwdata_reg[0]), .QN( ));
Q_FDP1 apb_pwrite_reg_REG  ( .CK(clk), .R(rst_n), .D(apb_pwrite), .Q(apb_pwrite_reg), .QN(n1));
Q_FDP1 apb_active_reg_REG  ( .CK(clk), .R(rst_n), .D(apb_active), .Q(apb_active_reg), .QN(n3));
Q_AN03 U59 ( .A0(n3), .A1(n2), .A2(apb_penable_reg), .Z(n4));
Q_AN02 U60 ( .A0(apb_psel_reg), .A1(n4), .Z(n13));
Q_OR03 U61 ( .A0(rbus_rd_strb_i), .A1(rbus_wr_strb_i), .A2(rbus_err_ack_i), .Z(n5));
Q_OR02 U62 ( .A0(rbus_ack_i), .A1(n5), .Z(n11));
Q_AN02 U63 ( .A0(n11), .A1(n5), .Z(n6));
Q_AN02 U64 ( .A0(n12), .A1(n1), .Z(n7));
Q_AN02 U65 ( .A0(n12), .A1(apb_pwrite_reg), .Z(n8));
Q_FDP1 rbus_wr_strb_o_REG  ( .CK(clk), .R(rst_n), .D(n8), .Q(rbus_wr_strb_o), .QN( ));
Q_FDP1 rbus_rd_strb_o_REG  ( .CK(clk), .R(rst_n), .D(n7), .Q(rbus_rd_strb_o), .QN( ));
Q_FDP1 apb_pslverr_REG  ( .CK(clk), .R(rst_n), .D(n6), .Q(apb_pslverr), .QN( ));
Q_FDP1 apb_pready_REG  ( .CK(clk), .R(rst_n), .D(n11), .Q(apb_pready), .QN(n9));
Q_AN02 U70 ( .A0(n13), .A1(n9), .Z(n12));
Q_OR02 U71 ( .A0(n13), .A1(apb_pready), .Z(n10));
Q_FDP4EP apb_active_REG_inst  ( .CK(clk), .CE(n10), .R(n14), .D(n9), .Q(apb_active));
Q_INV U73 ( .A(rst_n), .Z(n14));
Q_INV U74 ( .A(apb_active), .Z(n2));
Q_FDP4EP \apb_prdata_REG[0] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[0]), .Q(apb_prdata[0]));
Q_FDP4EP \apb_prdata_REG[1] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[1]), .Q(apb_prdata[1]));
Q_FDP4EP \apb_prdata_REG[2] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[2]), .Q(apb_prdata[2]));
Q_FDP4EP \apb_prdata_REG[3] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[3]), .Q(apb_prdata[3]));
Q_FDP4EP \apb_prdata_REG[4] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[4]), .Q(apb_prdata[4]));
Q_FDP4EP \apb_prdata_REG[5] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[5]), .Q(apb_prdata[5]));
Q_FDP4EP \apb_prdata_REG[6] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[6]), .Q(apb_prdata[6]));
Q_FDP4EP \apb_prdata_REG[7] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[7]), .Q(apb_prdata[7]));
Q_FDP4EP \apb_prdata_REG[8] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[8]), .Q(apb_prdata[8]));
Q_FDP4EP \apb_prdata_REG[9] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[9]), .Q(apb_prdata[9]));
Q_FDP4EP \apb_prdata_REG[10] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[10]), .Q(apb_prdata[10]));
Q_FDP4EP \apb_prdata_REG[11] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[11]), .Q(apb_prdata[11]));
Q_FDP4EP \apb_prdata_REG[12] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[12]), .Q(apb_prdata[12]));
Q_FDP4EP \apb_prdata_REG[13] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[13]), .Q(apb_prdata[13]));
Q_FDP4EP \apb_prdata_REG[14] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[14]), .Q(apb_prdata[14]));
Q_FDP4EP \apb_prdata_REG[15] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[15]), .Q(apb_prdata[15]));
Q_FDP4EP \apb_prdata_REG[16] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[16]), .Q(apb_prdata[16]));
Q_FDP4EP \apb_prdata_REG[17] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[17]), .Q(apb_prdata[17]));
Q_FDP4EP \apb_prdata_REG[18] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[18]), .Q(apb_prdata[18]));
Q_FDP4EP \apb_prdata_REG[19] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[19]), .Q(apb_prdata[19]));
Q_FDP4EP \apb_prdata_REG[20] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[20]), .Q(apb_prdata[20]));
Q_FDP4EP \apb_prdata_REG[21] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[21]), .Q(apb_prdata[21]));
Q_FDP4EP \apb_prdata_REG[22] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[22]), .Q(apb_prdata[22]));
Q_FDP4EP \apb_prdata_REG[23] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[23]), .Q(apb_prdata[23]));
Q_FDP4EP \apb_prdata_REG[24] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[24]), .Q(apb_prdata[24]));
Q_FDP4EP \apb_prdata_REG[25] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[25]), .Q(apb_prdata[25]));
Q_FDP4EP \apb_prdata_REG[26] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[26]), .Q(apb_prdata[26]));
Q_FDP4EP \apb_prdata_REG[27] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[27]), .Q(apb_prdata[27]));
Q_FDP4EP \apb_prdata_REG[28] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[28]), .Q(apb_prdata[28]));
Q_FDP4EP \apb_prdata_REG[29] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[29]), .Q(apb_prdata[29]));
Q_FDP4EP \apb_prdata_REG[30] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[30]), .Q(apb_prdata[30]));
Q_FDP4EP \apb_prdata_REG[31] ( .CK(clk), .CE(n11), .R(n14), .D(rbus_rd_data_i[31]), .Q(apb_prdata[31]));
Q_FDP4EP \rbus_wr_data_o_REG[0] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[0]), .Q(rbus_wr_data_o[0]));
Q_FDP4EP \rbus_wr_data_o_REG[1] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[1]), .Q(rbus_wr_data_o[1]));
Q_FDP4EP \rbus_wr_data_o_REG[2] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[2]), .Q(rbus_wr_data_o[2]));
Q_FDP4EP \rbus_wr_data_o_REG[3] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[3]), .Q(rbus_wr_data_o[3]));
Q_FDP4EP \rbus_wr_data_o_REG[4] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[4]), .Q(rbus_wr_data_o[4]));
Q_FDP4EP \rbus_wr_data_o_REG[5] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[5]), .Q(rbus_wr_data_o[5]));
Q_FDP4EP \rbus_wr_data_o_REG[6] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[6]), .Q(rbus_wr_data_o[6]));
Q_FDP4EP \rbus_wr_data_o_REG[7] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[7]), .Q(rbus_wr_data_o[7]));
Q_FDP4EP \rbus_wr_data_o_REG[8] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[8]), .Q(rbus_wr_data_o[8]));
Q_FDP4EP \rbus_wr_data_o_REG[9] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[9]), .Q(rbus_wr_data_o[9]));
Q_FDP4EP \rbus_wr_data_o_REG[10] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[10]), .Q(rbus_wr_data_o[10]));
Q_FDP4EP \rbus_wr_data_o_REG[11] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[11]), .Q(rbus_wr_data_o[11]));
Q_FDP4EP \rbus_wr_data_o_REG[12] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[12]), .Q(rbus_wr_data_o[12]));
Q_FDP4EP \rbus_wr_data_o_REG[13] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[13]), .Q(rbus_wr_data_o[13]));
Q_FDP4EP \rbus_wr_data_o_REG[14] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[14]), .Q(rbus_wr_data_o[14]));
Q_FDP4EP \rbus_wr_data_o_REG[15] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[15]), .Q(rbus_wr_data_o[15]));
Q_FDP4EP \rbus_wr_data_o_REG[16] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[16]), .Q(rbus_wr_data_o[16]));
Q_FDP4EP \rbus_wr_data_o_REG[17] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[17]), .Q(rbus_wr_data_o[17]));
Q_FDP4EP \rbus_wr_data_o_REG[18] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[18]), .Q(rbus_wr_data_o[18]));
Q_FDP4EP \rbus_wr_data_o_REG[19] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[19]), .Q(rbus_wr_data_o[19]));
Q_FDP4EP \rbus_wr_data_o_REG[20] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[20]), .Q(rbus_wr_data_o[20]));
Q_FDP4EP \rbus_wr_data_o_REG[21] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[21]), .Q(rbus_wr_data_o[21]));
Q_FDP4EP \rbus_wr_data_o_REG[22] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[22]), .Q(rbus_wr_data_o[22]));
Q_FDP4EP \rbus_wr_data_o_REG[23] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[23]), .Q(rbus_wr_data_o[23]));
Q_FDP4EP \rbus_wr_data_o_REG[24] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[24]), .Q(rbus_wr_data_o[24]));
Q_FDP4EP \rbus_wr_data_o_REG[25] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[25]), .Q(rbus_wr_data_o[25]));
Q_FDP4EP \rbus_wr_data_o_REG[26] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[26]), .Q(rbus_wr_data_o[26]));
Q_FDP4EP \rbus_wr_data_o_REG[27] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[27]), .Q(rbus_wr_data_o[27]));
Q_FDP4EP \rbus_wr_data_o_REG[28] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[28]), .Q(rbus_wr_data_o[28]));
Q_FDP4EP \rbus_wr_data_o_REG[29] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[29]), .Q(rbus_wr_data_o[29]));
Q_FDP4EP \rbus_wr_data_o_REG[30] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[30]), .Q(rbus_wr_data_o[30]));
Q_FDP4EP \rbus_wr_data_o_REG[31] ( .CK(clk), .CE(n12), .R(n14), .D(apb_pwdata_reg[31]), .Q(rbus_wr_data_o[31]));
Q_FDP4EP \rbus_addr_o_REG[0] ( .CK(clk), .CE(n12), .R(n14), .D(apb_paddr_reg[0]), .Q(rbus_addr_o[0]));
Q_FDP4EP \rbus_addr_o_REG[1] ( .CK(clk), .CE(n12), .R(n14), .D(apb_paddr_reg[1]), .Q(rbus_addr_o[1]));
Q_FDP4EP \rbus_addr_o_REG[2] ( .CK(clk), .CE(n12), .R(n14), .D(apb_paddr_reg[2]), .Q(rbus_addr_o[2]));
Q_FDP4EP \rbus_addr_o_REG[3] ( .CK(clk), .CE(n12), .R(n14), .D(apb_paddr_reg[3]), .Q(rbus_addr_o[3]));
Q_FDP4EP \rbus_addr_o_REG[4] ( .CK(clk), .CE(n12), .R(n14), .D(apb_paddr_reg[4]), .Q(rbus_addr_o[4]));
Q_FDP4EP \rbus_addr_o_REG[5] ( .CK(clk), .CE(n12), .R(n14), .D(apb_paddr_reg[5]), .Q(rbus_addr_o[5]));
Q_FDP4EP \rbus_addr_o_REG[6] ( .CK(clk), .CE(n12), .R(n14), .D(apb_paddr_reg[6]), .Q(rbus_addr_o[6]));
Q_FDP4EP \rbus_addr_o_REG[7] ( .CK(clk), .CE(n12), .R(n14), .D(apb_paddr_reg[7]), .Q(rbus_addr_o[7]));
Q_FDP4EP \rbus_addr_o_REG[8] ( .CK(clk), .CE(n12), .R(n14), .D(apb_paddr_reg[8]), .Q(rbus_addr_o[8]));
Q_FDP4EP \rbus_addr_o_REG[9] ( .CK(clk), .CE(n12), .R(n14), .D(apb_paddr_reg[9]), .Q(rbus_addr_o[9]));
Q_FDP4EP \rbus_addr_o_REG[10] ( .CK(clk), .CE(n12), .R(n14), .D(apb_paddr_reg[10]), .Q(rbus_addr_o[10]));
Q_FDP4EP \rbus_addr_o_REG[11] ( .CK(clk), .CE(n12), .R(n14), .D(apb_paddr_reg[11]), .Q(rbus_addr_o[11]));
Q_FDP4EP \rbus_addr_o_REG[12] ( .CK(clk), .CE(n12), .R(n14), .D(apb_paddr_reg[12]), .Q(rbus_addr_o[12]));
Q_FDP4EP \rbus_addr_o_REG[13] ( .CK(clk), .CE(n12), .R(n14), .D(apb_paddr_reg[13]), .Q(rbus_addr_o[13]));
Q_FDP4EP \rbus_addr_o_REG[14] ( .CK(clk), .CE(n12), .R(n14), .D(apb_paddr_reg[14]), .Q(rbus_addr_o[14]));
Q_FDP4EP \rbus_addr_o_REG[15] ( .CK(clk), .CE(n12), .R(n14), .D(apb_paddr_reg[15]), .Q(rbus_addr_o[15]));
endmodule
