
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module cr_kme_drng ( drng_health_fail, drng_seed_expired, drng_256_out, 
	drng_valid, seed0_invalidate, seed1_invalidate, stat_drbg_reseed, 
	drng_idle, clk, rst_n, drng_ack, seed0_valid, 
	seed0_internal_state_key, seed0_internal_state_value, 
	seed0_reseed_interval, seed1_valid, seed1_internal_state_key, 
	seed1_internal_state_value, seed1_reseed_interval);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output drng_health_fail;
output drng_seed_expired;
output [127:0] drng_256_out;
output drng_valid;
output seed0_invalidate;
output seed1_invalidate;
output stat_drbg_reseed;
output drng_idle;
input clk;
input rst_n;
input drng_ack;
input seed0_valid;
input [255:0] seed0_internal_state_key;
input [127:0] seed0_internal_state_value;
input [47:0] seed0_reseed_interval;
input seed1_valid;
input [255:0] seed1_internal_state_key;
input [127:0] seed1_internal_state_value;
input [47:0] seed1_reseed_interval;
wire seed_expired;
wire drng_health_test;
wire [127:0] drng_256_out_pre;
wire _zy_simnet_drng_health_fail_0_w$;
wire _zy_simnet_dio_1;
wire _zy_simnet_dio_2;
wire _zy_simnet_seed_valid_3_w$;
wire [0:383] _zy_simnet_seed_4_w$;
wire [0:47] _zy_simnet_seed_life_5_w$;
wire [127:0] drng_256_last;
wire drng_first;
wire [0:0] seed_entry;
supply1 n1;
Q_MX02 U0 ( .S(seed_entry[0]), .A0(\seed_valid[0][0] ), .A1(\seed_valid[1][0] ), .Z(n435));
Q_MX02 U1 ( .S(seed_entry[0]), .A0(\seed_life[0][47] ), .A1(\seed_life[1][47] ), .Z(n2));
Q_MX02 U2 ( .S(seed_entry[0]), .A0(\seed_life[0][46] ), .A1(\seed_life[1][46] ), .Z(n3));
Q_MX02 U3 ( .S(seed_entry[0]), .A0(\seed_life[0][45] ), .A1(\seed_life[1][45] ), .Z(n4));
Q_MX02 U4 ( .S(seed_entry[0]), .A0(\seed_life[0][44] ), .A1(\seed_life[1][44] ), .Z(n5));
Q_MX02 U5 ( .S(seed_entry[0]), .A0(\seed_life[0][43] ), .A1(\seed_life[1][43] ), .Z(n6));
Q_MX02 U6 ( .S(seed_entry[0]), .A0(\seed_life[0][42] ), .A1(\seed_life[1][42] ), .Z(n7));
Q_MX02 U7 ( .S(seed_entry[0]), .A0(\seed_life[0][41] ), .A1(\seed_life[1][41] ), .Z(n8));
Q_MX02 U8 ( .S(seed_entry[0]), .A0(\seed_life[0][40] ), .A1(\seed_life[1][40] ), .Z(n9));
Q_MX02 U9 ( .S(seed_entry[0]), .A0(\seed_life[0][39] ), .A1(\seed_life[1][39] ), .Z(n10));
Q_MX02 U10 ( .S(seed_entry[0]), .A0(\seed_life[0][38] ), .A1(\seed_life[1][38] ), .Z(n11));
Q_MX02 U11 ( .S(seed_entry[0]), .A0(\seed_life[0][37] ), .A1(\seed_life[1][37] ), .Z(n12));
Q_MX02 U12 ( .S(seed_entry[0]), .A0(\seed_life[0][36] ), .A1(\seed_life[1][36] ), .Z(n13));
Q_MX02 U13 ( .S(seed_entry[0]), .A0(\seed_life[0][35] ), .A1(\seed_life[1][35] ), .Z(n14));
Q_MX02 U14 ( .S(seed_entry[0]), .A0(\seed_life[0][34] ), .A1(\seed_life[1][34] ), .Z(n15));
Q_MX02 U15 ( .S(seed_entry[0]), .A0(\seed_life[0][33] ), .A1(\seed_life[1][33] ), .Z(n16));
Q_MX02 U16 ( .S(seed_entry[0]), .A0(\seed_life[0][32] ), .A1(\seed_life[1][32] ), .Z(n17));
Q_MX02 U17 ( .S(seed_entry[0]), .A0(\seed_life[0][31] ), .A1(\seed_life[1][31] ), .Z(n18));
Q_MX02 U18 ( .S(seed_entry[0]), .A0(\seed_life[0][30] ), .A1(\seed_life[1][30] ), .Z(n19));
Q_MX02 U19 ( .S(seed_entry[0]), .A0(\seed_life[0][29] ), .A1(\seed_life[1][29] ), .Z(n20));
Q_MX02 U20 ( .S(seed_entry[0]), .A0(\seed_life[0][28] ), .A1(\seed_life[1][28] ), .Z(n21));
Q_MX02 U21 ( .S(seed_entry[0]), .A0(\seed_life[0][27] ), .A1(\seed_life[1][27] ), .Z(n22));
Q_MX02 U22 ( .S(seed_entry[0]), .A0(\seed_life[0][26] ), .A1(\seed_life[1][26] ), .Z(n23));
Q_MX02 U23 ( .S(seed_entry[0]), .A0(\seed_life[0][25] ), .A1(\seed_life[1][25] ), .Z(n24));
Q_MX02 U24 ( .S(seed_entry[0]), .A0(\seed_life[0][24] ), .A1(\seed_life[1][24] ), .Z(n25));
Q_MX02 U25 ( .S(seed_entry[0]), .A0(\seed_life[0][23] ), .A1(\seed_life[1][23] ), .Z(n26));
Q_MX02 U26 ( .S(seed_entry[0]), .A0(\seed_life[0][22] ), .A1(\seed_life[1][22] ), .Z(n27));
Q_MX02 U27 ( .S(seed_entry[0]), .A0(\seed_life[0][21] ), .A1(\seed_life[1][21] ), .Z(n28));
Q_MX02 U28 ( .S(seed_entry[0]), .A0(\seed_life[0][20] ), .A1(\seed_life[1][20] ), .Z(n29));
Q_MX02 U29 ( .S(seed_entry[0]), .A0(\seed_life[0][19] ), .A1(\seed_life[1][19] ), .Z(n30));
Q_MX02 U30 ( .S(seed_entry[0]), .A0(\seed_life[0][18] ), .A1(\seed_life[1][18] ), .Z(n31));
Q_MX02 U31 ( .S(seed_entry[0]), .A0(\seed_life[0][17] ), .A1(\seed_life[1][17] ), .Z(n32));
Q_MX02 U32 ( .S(seed_entry[0]), .A0(\seed_life[0][16] ), .A1(\seed_life[1][16] ), .Z(n33));
Q_MX02 U33 ( .S(seed_entry[0]), .A0(\seed_life[0][15] ), .A1(\seed_life[1][15] ), .Z(n34));
Q_MX02 U34 ( .S(seed_entry[0]), .A0(\seed_life[0][14] ), .A1(\seed_life[1][14] ), .Z(n35));
Q_MX02 U35 ( .S(seed_entry[0]), .A0(\seed_life[0][13] ), .A1(\seed_life[1][13] ), .Z(n36));
Q_MX02 U36 ( .S(seed_entry[0]), .A0(\seed_life[0][12] ), .A1(\seed_life[1][12] ), .Z(n37));
Q_MX02 U37 ( .S(seed_entry[0]), .A0(\seed_life[0][11] ), .A1(\seed_life[1][11] ), .Z(n38));
Q_MX02 U38 ( .S(seed_entry[0]), .A0(\seed_life[0][10] ), .A1(\seed_life[1][10] ), .Z(n39));
Q_MX02 U39 ( .S(seed_entry[0]), .A0(\seed_life[0][9] ), .A1(\seed_life[1][9] ), .Z(n40));
Q_MX02 U40 ( .S(seed_entry[0]), .A0(\seed_life[0][8] ), .A1(\seed_life[1][8] ), .Z(n41));
Q_MX02 U41 ( .S(seed_entry[0]), .A0(\seed_life[0][7] ), .A1(\seed_life[1][7] ), .Z(n42));
Q_MX02 U42 ( .S(seed_entry[0]), .A0(\seed_life[0][6] ), .A1(\seed_life[1][6] ), .Z(n43));
Q_MX02 U43 ( .S(seed_entry[0]), .A0(\seed_life[0][5] ), .A1(\seed_life[1][5] ), .Z(n44));
Q_MX02 U44 ( .S(seed_entry[0]), .A0(\seed_life[0][4] ), .A1(\seed_life[1][4] ), .Z(n45));
Q_MX02 U45 ( .S(seed_entry[0]), .A0(\seed_life[0][3] ), .A1(\seed_life[1][3] ), .Z(n46));
Q_MX02 U46 ( .S(seed_entry[0]), .A0(\seed_life[0][2] ), .A1(\seed_life[1][2] ), .Z(n47));
Q_MX02 U47 ( .S(seed_entry[0]), .A0(\seed_life[0][1] ), .A1(\seed_life[1][1] ), .Z(n48));
Q_MX02 U48 ( .S(seed_entry[0]), .A0(\seed_life[0][0] ), .A1(\seed_life[1][0] ), .Z(n49));
Q_MX02 U49 ( .S(seed_entry[0]), .A0(\seed[0][383] ), .A1(\seed[1][383] ), .Z(n50));
Q_MX02 U50 ( .S(seed_entry[0]), .A0(\seed[0][382] ), .A1(\seed[1][382] ), .Z(n51));
Q_MX02 U51 ( .S(seed_entry[0]), .A0(\seed[0][381] ), .A1(\seed[1][381] ), .Z(n52));
Q_MX02 U52 ( .S(seed_entry[0]), .A0(\seed[0][380] ), .A1(\seed[1][380] ), .Z(n53));
Q_MX02 U53 ( .S(seed_entry[0]), .A0(\seed[0][379] ), .A1(\seed[1][379] ), .Z(n54));
Q_MX02 U54 ( .S(seed_entry[0]), .A0(\seed[0][378] ), .A1(\seed[1][378] ), .Z(n55));
Q_MX02 U55 ( .S(seed_entry[0]), .A0(\seed[0][377] ), .A1(\seed[1][377] ), .Z(n56));
Q_MX02 U56 ( .S(seed_entry[0]), .A0(\seed[0][376] ), .A1(\seed[1][376] ), .Z(n57));
Q_MX02 U57 ( .S(seed_entry[0]), .A0(\seed[0][375] ), .A1(\seed[1][375] ), .Z(n58));
Q_MX02 U58 ( .S(seed_entry[0]), .A0(\seed[0][374] ), .A1(\seed[1][374] ), .Z(n59));
Q_MX02 U59 ( .S(seed_entry[0]), .A0(\seed[0][373] ), .A1(\seed[1][373] ), .Z(n60));
Q_MX02 U60 ( .S(seed_entry[0]), .A0(\seed[0][372] ), .A1(\seed[1][372] ), .Z(n61));
Q_MX02 U61 ( .S(seed_entry[0]), .A0(\seed[0][371] ), .A1(\seed[1][371] ), .Z(n62));
Q_MX02 U62 ( .S(seed_entry[0]), .A0(\seed[0][370] ), .A1(\seed[1][370] ), .Z(n63));
Q_MX02 U63 ( .S(seed_entry[0]), .A0(\seed[0][369] ), .A1(\seed[1][369] ), .Z(n64));
Q_MX02 U64 ( .S(seed_entry[0]), .A0(\seed[0][368] ), .A1(\seed[1][368] ), .Z(n65));
Q_MX02 U65 ( .S(seed_entry[0]), .A0(\seed[0][367] ), .A1(\seed[1][367] ), .Z(n66));
Q_MX02 U66 ( .S(seed_entry[0]), .A0(\seed[0][366] ), .A1(\seed[1][366] ), .Z(n67));
Q_MX02 U67 ( .S(seed_entry[0]), .A0(\seed[0][365] ), .A1(\seed[1][365] ), .Z(n68));
Q_MX02 U68 ( .S(seed_entry[0]), .A0(\seed[0][364] ), .A1(\seed[1][364] ), .Z(n69));
Q_MX02 U69 ( .S(seed_entry[0]), .A0(\seed[0][363] ), .A1(\seed[1][363] ), .Z(n70));
Q_MX02 U70 ( .S(seed_entry[0]), .A0(\seed[0][362] ), .A1(\seed[1][362] ), .Z(n71));
Q_MX02 U71 ( .S(seed_entry[0]), .A0(\seed[0][361] ), .A1(\seed[1][361] ), .Z(n72));
Q_MX02 U72 ( .S(seed_entry[0]), .A0(\seed[0][360] ), .A1(\seed[1][360] ), .Z(n73));
Q_MX02 U73 ( .S(seed_entry[0]), .A0(\seed[0][359] ), .A1(\seed[1][359] ), .Z(n74));
Q_MX02 U74 ( .S(seed_entry[0]), .A0(\seed[0][358] ), .A1(\seed[1][358] ), .Z(n75));
Q_MX02 U75 ( .S(seed_entry[0]), .A0(\seed[0][357] ), .A1(\seed[1][357] ), .Z(n76));
Q_MX02 U76 ( .S(seed_entry[0]), .A0(\seed[0][356] ), .A1(\seed[1][356] ), .Z(n77));
Q_MX02 U77 ( .S(seed_entry[0]), .A0(\seed[0][355] ), .A1(\seed[1][355] ), .Z(n78));
Q_MX02 U78 ( .S(seed_entry[0]), .A0(\seed[0][354] ), .A1(\seed[1][354] ), .Z(n79));
Q_MX02 U79 ( .S(seed_entry[0]), .A0(\seed[0][353] ), .A1(\seed[1][353] ), .Z(n80));
Q_MX02 U80 ( .S(seed_entry[0]), .A0(\seed[0][352] ), .A1(\seed[1][352] ), .Z(n81));
Q_MX02 U81 ( .S(seed_entry[0]), .A0(\seed[0][351] ), .A1(\seed[1][351] ), .Z(n82));
Q_MX02 U82 ( .S(seed_entry[0]), .A0(\seed[0][350] ), .A1(\seed[1][350] ), .Z(n83));
Q_MX02 U83 ( .S(seed_entry[0]), .A0(\seed[0][349] ), .A1(\seed[1][349] ), .Z(n84));
Q_MX02 U84 ( .S(seed_entry[0]), .A0(\seed[0][348] ), .A1(\seed[1][348] ), .Z(n85));
Q_MX02 U85 ( .S(seed_entry[0]), .A0(\seed[0][347] ), .A1(\seed[1][347] ), .Z(n86));
Q_MX02 U86 ( .S(seed_entry[0]), .A0(\seed[0][346] ), .A1(\seed[1][346] ), .Z(n87));
Q_MX02 U87 ( .S(seed_entry[0]), .A0(\seed[0][345] ), .A1(\seed[1][345] ), .Z(n88));
Q_MX02 U88 ( .S(seed_entry[0]), .A0(\seed[0][344] ), .A1(\seed[1][344] ), .Z(n89));
Q_MX02 U89 ( .S(seed_entry[0]), .A0(\seed[0][343] ), .A1(\seed[1][343] ), .Z(n90));
Q_MX02 U90 ( .S(seed_entry[0]), .A0(\seed[0][342] ), .A1(\seed[1][342] ), .Z(n91));
Q_MX02 U91 ( .S(seed_entry[0]), .A0(\seed[0][341] ), .A1(\seed[1][341] ), .Z(n92));
Q_MX02 U92 ( .S(seed_entry[0]), .A0(\seed[0][340] ), .A1(\seed[1][340] ), .Z(n93));
Q_MX02 U93 ( .S(seed_entry[0]), .A0(\seed[0][339] ), .A1(\seed[1][339] ), .Z(n94));
Q_MX02 U94 ( .S(seed_entry[0]), .A0(\seed[0][338] ), .A1(\seed[1][338] ), .Z(n95));
Q_MX02 U95 ( .S(seed_entry[0]), .A0(\seed[0][337] ), .A1(\seed[1][337] ), .Z(n96));
Q_MX02 U96 ( .S(seed_entry[0]), .A0(\seed[0][336] ), .A1(\seed[1][336] ), .Z(n97));
Q_MX02 U97 ( .S(seed_entry[0]), .A0(\seed[0][335] ), .A1(\seed[1][335] ), .Z(n98));
Q_MX02 U98 ( .S(seed_entry[0]), .A0(\seed[0][334] ), .A1(\seed[1][334] ), .Z(n99));
Q_MX02 U99 ( .S(seed_entry[0]), .A0(\seed[0][333] ), .A1(\seed[1][333] ), .Z(n100));
Q_MX02 U100 ( .S(seed_entry[0]), .A0(\seed[0][332] ), .A1(\seed[1][332] ), .Z(n101));
Q_MX02 U101 ( .S(seed_entry[0]), .A0(\seed[0][331] ), .A1(\seed[1][331] ), .Z(n102));
Q_MX02 U102 ( .S(seed_entry[0]), .A0(\seed[0][330] ), .A1(\seed[1][330] ), .Z(n103));
Q_MX02 U103 ( .S(seed_entry[0]), .A0(\seed[0][329] ), .A1(\seed[1][329] ), .Z(n104));
Q_MX02 U104 ( .S(seed_entry[0]), .A0(\seed[0][328] ), .A1(\seed[1][328] ), .Z(n105));
Q_MX02 U105 ( .S(seed_entry[0]), .A0(\seed[0][327] ), .A1(\seed[1][327] ), .Z(n106));
Q_MX02 U106 ( .S(seed_entry[0]), .A0(\seed[0][326] ), .A1(\seed[1][326] ), .Z(n107));
Q_MX02 U107 ( .S(seed_entry[0]), .A0(\seed[0][325] ), .A1(\seed[1][325] ), .Z(n108));
Q_MX02 U108 ( .S(seed_entry[0]), .A0(\seed[0][324] ), .A1(\seed[1][324] ), .Z(n109));
Q_MX02 U109 ( .S(seed_entry[0]), .A0(\seed[0][323] ), .A1(\seed[1][323] ), .Z(n110));
Q_MX02 U110 ( .S(seed_entry[0]), .A0(\seed[0][322] ), .A1(\seed[1][322] ), .Z(n111));
Q_MX02 U111 ( .S(seed_entry[0]), .A0(\seed[0][321] ), .A1(\seed[1][321] ), .Z(n112));
Q_MX02 U112 ( .S(seed_entry[0]), .A0(\seed[0][320] ), .A1(\seed[1][320] ), .Z(n113));
Q_MX02 U113 ( .S(seed_entry[0]), .A0(\seed[0][319] ), .A1(\seed[1][319] ), .Z(n114));
Q_MX02 U114 ( .S(seed_entry[0]), .A0(\seed[0][318] ), .A1(\seed[1][318] ), .Z(n115));
Q_MX02 U115 ( .S(seed_entry[0]), .A0(\seed[0][317] ), .A1(\seed[1][317] ), .Z(n116));
Q_MX02 U116 ( .S(seed_entry[0]), .A0(\seed[0][316] ), .A1(\seed[1][316] ), .Z(n117));
Q_MX02 U117 ( .S(seed_entry[0]), .A0(\seed[0][315] ), .A1(\seed[1][315] ), .Z(n118));
Q_MX02 U118 ( .S(seed_entry[0]), .A0(\seed[0][314] ), .A1(\seed[1][314] ), .Z(n119));
Q_MX02 U119 ( .S(seed_entry[0]), .A0(\seed[0][313] ), .A1(\seed[1][313] ), .Z(n120));
Q_MX02 U120 ( .S(seed_entry[0]), .A0(\seed[0][312] ), .A1(\seed[1][312] ), .Z(n121));
Q_MX02 U121 ( .S(seed_entry[0]), .A0(\seed[0][311] ), .A1(\seed[1][311] ), .Z(n122));
Q_MX02 U122 ( .S(seed_entry[0]), .A0(\seed[0][310] ), .A1(\seed[1][310] ), .Z(n123));
Q_MX02 U123 ( .S(seed_entry[0]), .A0(\seed[0][309] ), .A1(\seed[1][309] ), .Z(n124));
Q_MX02 U124 ( .S(seed_entry[0]), .A0(\seed[0][308] ), .A1(\seed[1][308] ), .Z(n125));
Q_MX02 U125 ( .S(seed_entry[0]), .A0(\seed[0][307] ), .A1(\seed[1][307] ), .Z(n126));
Q_MX02 U126 ( .S(seed_entry[0]), .A0(\seed[0][306] ), .A1(\seed[1][306] ), .Z(n127));
Q_MX02 U127 ( .S(seed_entry[0]), .A0(\seed[0][305] ), .A1(\seed[1][305] ), .Z(n128));
Q_MX02 U128 ( .S(seed_entry[0]), .A0(\seed[0][304] ), .A1(\seed[1][304] ), .Z(n129));
Q_MX02 U129 ( .S(seed_entry[0]), .A0(\seed[0][303] ), .A1(\seed[1][303] ), .Z(n130));
Q_MX02 U130 ( .S(seed_entry[0]), .A0(\seed[0][302] ), .A1(\seed[1][302] ), .Z(n131));
Q_MX02 U131 ( .S(seed_entry[0]), .A0(\seed[0][301] ), .A1(\seed[1][301] ), .Z(n132));
Q_MX02 U132 ( .S(seed_entry[0]), .A0(\seed[0][300] ), .A1(\seed[1][300] ), .Z(n133));
Q_MX02 U133 ( .S(seed_entry[0]), .A0(\seed[0][299] ), .A1(\seed[1][299] ), .Z(n134));
Q_MX02 U134 ( .S(seed_entry[0]), .A0(\seed[0][298] ), .A1(\seed[1][298] ), .Z(n135));
Q_MX02 U135 ( .S(seed_entry[0]), .A0(\seed[0][297] ), .A1(\seed[1][297] ), .Z(n136));
Q_MX02 U136 ( .S(seed_entry[0]), .A0(\seed[0][296] ), .A1(\seed[1][296] ), .Z(n137));
Q_MX02 U137 ( .S(seed_entry[0]), .A0(\seed[0][295] ), .A1(\seed[1][295] ), .Z(n138));
Q_MX02 U138 ( .S(seed_entry[0]), .A0(\seed[0][294] ), .A1(\seed[1][294] ), .Z(n139));
Q_MX02 U139 ( .S(seed_entry[0]), .A0(\seed[0][293] ), .A1(\seed[1][293] ), .Z(n140));
Q_MX02 U140 ( .S(seed_entry[0]), .A0(\seed[0][292] ), .A1(\seed[1][292] ), .Z(n141));
Q_MX02 U141 ( .S(seed_entry[0]), .A0(\seed[0][291] ), .A1(\seed[1][291] ), .Z(n142));
Q_MX02 U142 ( .S(seed_entry[0]), .A0(\seed[0][290] ), .A1(\seed[1][290] ), .Z(n143));
Q_MX02 U143 ( .S(seed_entry[0]), .A0(\seed[0][289] ), .A1(\seed[1][289] ), .Z(n144));
Q_MX02 U144 ( .S(seed_entry[0]), .A0(\seed[0][288] ), .A1(\seed[1][288] ), .Z(n145));
Q_MX02 U145 ( .S(seed_entry[0]), .A0(\seed[0][287] ), .A1(\seed[1][287] ), .Z(n146));
Q_MX02 U146 ( .S(seed_entry[0]), .A0(\seed[0][286] ), .A1(\seed[1][286] ), .Z(n147));
Q_MX02 U147 ( .S(seed_entry[0]), .A0(\seed[0][285] ), .A1(\seed[1][285] ), .Z(n148));
Q_MX02 U148 ( .S(seed_entry[0]), .A0(\seed[0][284] ), .A1(\seed[1][284] ), .Z(n149));
Q_MX02 U149 ( .S(seed_entry[0]), .A0(\seed[0][283] ), .A1(\seed[1][283] ), .Z(n150));
Q_MX02 U150 ( .S(seed_entry[0]), .A0(\seed[0][282] ), .A1(\seed[1][282] ), .Z(n151));
Q_MX02 U151 ( .S(seed_entry[0]), .A0(\seed[0][281] ), .A1(\seed[1][281] ), .Z(n152));
Q_MX02 U152 ( .S(seed_entry[0]), .A0(\seed[0][280] ), .A1(\seed[1][280] ), .Z(n153));
Q_MX02 U153 ( .S(seed_entry[0]), .A0(\seed[0][279] ), .A1(\seed[1][279] ), .Z(n154));
Q_MX02 U154 ( .S(seed_entry[0]), .A0(\seed[0][278] ), .A1(\seed[1][278] ), .Z(n155));
Q_MX02 U155 ( .S(seed_entry[0]), .A0(\seed[0][277] ), .A1(\seed[1][277] ), .Z(n156));
Q_MX02 U156 ( .S(seed_entry[0]), .A0(\seed[0][276] ), .A1(\seed[1][276] ), .Z(n157));
Q_MX02 U157 ( .S(seed_entry[0]), .A0(\seed[0][275] ), .A1(\seed[1][275] ), .Z(n158));
Q_MX02 U158 ( .S(seed_entry[0]), .A0(\seed[0][274] ), .A1(\seed[1][274] ), .Z(n159));
Q_MX02 U159 ( .S(seed_entry[0]), .A0(\seed[0][273] ), .A1(\seed[1][273] ), .Z(n160));
Q_MX02 U160 ( .S(seed_entry[0]), .A0(\seed[0][272] ), .A1(\seed[1][272] ), .Z(n161));
Q_MX02 U161 ( .S(seed_entry[0]), .A0(\seed[0][271] ), .A1(\seed[1][271] ), .Z(n162));
Q_MX02 U162 ( .S(seed_entry[0]), .A0(\seed[0][270] ), .A1(\seed[1][270] ), .Z(n163));
Q_MX02 U163 ( .S(seed_entry[0]), .A0(\seed[0][269] ), .A1(\seed[1][269] ), .Z(n164));
Q_MX02 U164 ( .S(seed_entry[0]), .A0(\seed[0][268] ), .A1(\seed[1][268] ), .Z(n165));
Q_MX02 U165 ( .S(seed_entry[0]), .A0(\seed[0][267] ), .A1(\seed[1][267] ), .Z(n166));
Q_MX02 U166 ( .S(seed_entry[0]), .A0(\seed[0][266] ), .A1(\seed[1][266] ), .Z(n167));
Q_MX02 U167 ( .S(seed_entry[0]), .A0(\seed[0][265] ), .A1(\seed[1][265] ), .Z(n168));
Q_MX02 U168 ( .S(seed_entry[0]), .A0(\seed[0][264] ), .A1(\seed[1][264] ), .Z(n169));
Q_MX02 U169 ( .S(seed_entry[0]), .A0(\seed[0][263] ), .A1(\seed[1][263] ), .Z(n170));
Q_MX02 U170 ( .S(seed_entry[0]), .A0(\seed[0][262] ), .A1(\seed[1][262] ), .Z(n171));
Q_MX02 U171 ( .S(seed_entry[0]), .A0(\seed[0][261] ), .A1(\seed[1][261] ), .Z(n172));
Q_MX02 U172 ( .S(seed_entry[0]), .A0(\seed[0][260] ), .A1(\seed[1][260] ), .Z(n173));
Q_MX02 U173 ( .S(seed_entry[0]), .A0(\seed[0][259] ), .A1(\seed[1][259] ), .Z(n174));
Q_MX02 U174 ( .S(seed_entry[0]), .A0(\seed[0][258] ), .A1(\seed[1][258] ), .Z(n175));
Q_MX02 U175 ( .S(seed_entry[0]), .A0(\seed[0][257] ), .A1(\seed[1][257] ), .Z(n176));
Q_MX02 U176 ( .S(seed_entry[0]), .A0(\seed[0][256] ), .A1(\seed[1][256] ), .Z(n177));
Q_MX02 U177 ( .S(seed_entry[0]), .A0(\seed[0][255] ), .A1(\seed[1][255] ), .Z(n178));
Q_MX02 U178 ( .S(seed_entry[0]), .A0(\seed[0][254] ), .A1(\seed[1][254] ), .Z(n179));
Q_MX02 U179 ( .S(seed_entry[0]), .A0(\seed[0][253] ), .A1(\seed[1][253] ), .Z(n180));
Q_MX02 U180 ( .S(seed_entry[0]), .A0(\seed[0][252] ), .A1(\seed[1][252] ), .Z(n181));
Q_MX02 U181 ( .S(seed_entry[0]), .A0(\seed[0][251] ), .A1(\seed[1][251] ), .Z(n182));
Q_MX02 U182 ( .S(seed_entry[0]), .A0(\seed[0][250] ), .A1(\seed[1][250] ), .Z(n183));
Q_MX02 U183 ( .S(seed_entry[0]), .A0(\seed[0][249] ), .A1(\seed[1][249] ), .Z(n184));
Q_MX02 U184 ( .S(seed_entry[0]), .A0(\seed[0][248] ), .A1(\seed[1][248] ), .Z(n185));
Q_MX02 U185 ( .S(seed_entry[0]), .A0(\seed[0][247] ), .A1(\seed[1][247] ), .Z(n186));
Q_MX02 U186 ( .S(seed_entry[0]), .A0(\seed[0][246] ), .A1(\seed[1][246] ), .Z(n187));
Q_MX02 U187 ( .S(seed_entry[0]), .A0(\seed[0][245] ), .A1(\seed[1][245] ), .Z(n188));
Q_MX02 U188 ( .S(seed_entry[0]), .A0(\seed[0][244] ), .A1(\seed[1][244] ), .Z(n189));
Q_MX02 U189 ( .S(seed_entry[0]), .A0(\seed[0][243] ), .A1(\seed[1][243] ), .Z(n190));
Q_MX02 U190 ( .S(seed_entry[0]), .A0(\seed[0][242] ), .A1(\seed[1][242] ), .Z(n191));
Q_MX02 U191 ( .S(seed_entry[0]), .A0(\seed[0][241] ), .A1(\seed[1][241] ), .Z(n192));
Q_MX02 U192 ( .S(seed_entry[0]), .A0(\seed[0][240] ), .A1(\seed[1][240] ), .Z(n193));
Q_MX02 U193 ( .S(seed_entry[0]), .A0(\seed[0][239] ), .A1(\seed[1][239] ), .Z(n194));
Q_MX02 U194 ( .S(seed_entry[0]), .A0(\seed[0][238] ), .A1(\seed[1][238] ), .Z(n195));
Q_MX02 U195 ( .S(seed_entry[0]), .A0(\seed[0][237] ), .A1(\seed[1][237] ), .Z(n196));
Q_MX02 U196 ( .S(seed_entry[0]), .A0(\seed[0][236] ), .A1(\seed[1][236] ), .Z(n197));
Q_MX02 U197 ( .S(seed_entry[0]), .A0(\seed[0][235] ), .A1(\seed[1][235] ), .Z(n198));
Q_MX02 U198 ( .S(seed_entry[0]), .A0(\seed[0][234] ), .A1(\seed[1][234] ), .Z(n199));
Q_MX02 U199 ( .S(seed_entry[0]), .A0(\seed[0][233] ), .A1(\seed[1][233] ), .Z(n200));
Q_MX02 U200 ( .S(seed_entry[0]), .A0(\seed[0][232] ), .A1(\seed[1][232] ), .Z(n201));
Q_MX02 U201 ( .S(seed_entry[0]), .A0(\seed[0][231] ), .A1(\seed[1][231] ), .Z(n202));
Q_MX02 U202 ( .S(seed_entry[0]), .A0(\seed[0][230] ), .A1(\seed[1][230] ), .Z(n203));
Q_MX02 U203 ( .S(seed_entry[0]), .A0(\seed[0][229] ), .A1(\seed[1][229] ), .Z(n204));
Q_MX02 U204 ( .S(seed_entry[0]), .A0(\seed[0][228] ), .A1(\seed[1][228] ), .Z(n205));
Q_MX02 U205 ( .S(seed_entry[0]), .A0(\seed[0][227] ), .A1(\seed[1][227] ), .Z(n206));
Q_MX02 U206 ( .S(seed_entry[0]), .A0(\seed[0][226] ), .A1(\seed[1][226] ), .Z(n207));
Q_MX02 U207 ( .S(seed_entry[0]), .A0(\seed[0][225] ), .A1(\seed[1][225] ), .Z(n208));
Q_MX02 U208 ( .S(seed_entry[0]), .A0(\seed[0][224] ), .A1(\seed[1][224] ), .Z(n209));
Q_MX02 U209 ( .S(seed_entry[0]), .A0(\seed[0][223] ), .A1(\seed[1][223] ), .Z(n210));
Q_MX02 U210 ( .S(seed_entry[0]), .A0(\seed[0][222] ), .A1(\seed[1][222] ), .Z(n211));
Q_MX02 U211 ( .S(seed_entry[0]), .A0(\seed[0][221] ), .A1(\seed[1][221] ), .Z(n212));
Q_MX02 U212 ( .S(seed_entry[0]), .A0(\seed[0][220] ), .A1(\seed[1][220] ), .Z(n213));
Q_MX02 U213 ( .S(seed_entry[0]), .A0(\seed[0][219] ), .A1(\seed[1][219] ), .Z(n214));
Q_MX02 U214 ( .S(seed_entry[0]), .A0(\seed[0][218] ), .A1(\seed[1][218] ), .Z(n215));
Q_MX02 U215 ( .S(seed_entry[0]), .A0(\seed[0][217] ), .A1(\seed[1][217] ), .Z(n216));
Q_MX02 U216 ( .S(seed_entry[0]), .A0(\seed[0][216] ), .A1(\seed[1][216] ), .Z(n217));
Q_MX02 U217 ( .S(seed_entry[0]), .A0(\seed[0][215] ), .A1(\seed[1][215] ), .Z(n218));
Q_MX02 U218 ( .S(seed_entry[0]), .A0(\seed[0][214] ), .A1(\seed[1][214] ), .Z(n219));
Q_MX02 U219 ( .S(seed_entry[0]), .A0(\seed[0][213] ), .A1(\seed[1][213] ), .Z(n220));
Q_MX02 U220 ( .S(seed_entry[0]), .A0(\seed[0][212] ), .A1(\seed[1][212] ), .Z(n221));
Q_MX02 U221 ( .S(seed_entry[0]), .A0(\seed[0][211] ), .A1(\seed[1][211] ), .Z(n222));
Q_MX02 U222 ( .S(seed_entry[0]), .A0(\seed[0][210] ), .A1(\seed[1][210] ), .Z(n223));
Q_MX02 U223 ( .S(seed_entry[0]), .A0(\seed[0][209] ), .A1(\seed[1][209] ), .Z(n224));
Q_MX02 U224 ( .S(seed_entry[0]), .A0(\seed[0][208] ), .A1(\seed[1][208] ), .Z(n225));
Q_MX02 U225 ( .S(seed_entry[0]), .A0(\seed[0][207] ), .A1(\seed[1][207] ), .Z(n226));
Q_MX02 U226 ( .S(seed_entry[0]), .A0(\seed[0][206] ), .A1(\seed[1][206] ), .Z(n227));
Q_MX02 U227 ( .S(seed_entry[0]), .A0(\seed[0][205] ), .A1(\seed[1][205] ), .Z(n228));
Q_MX02 U228 ( .S(seed_entry[0]), .A0(\seed[0][204] ), .A1(\seed[1][204] ), .Z(n229));
Q_MX02 U229 ( .S(seed_entry[0]), .A0(\seed[0][203] ), .A1(\seed[1][203] ), .Z(n230));
Q_MX02 U230 ( .S(seed_entry[0]), .A0(\seed[0][202] ), .A1(\seed[1][202] ), .Z(n231));
Q_MX02 U231 ( .S(seed_entry[0]), .A0(\seed[0][201] ), .A1(\seed[1][201] ), .Z(n232));
Q_MX02 U232 ( .S(seed_entry[0]), .A0(\seed[0][200] ), .A1(\seed[1][200] ), .Z(n233));
Q_MX02 U233 ( .S(seed_entry[0]), .A0(\seed[0][199] ), .A1(\seed[1][199] ), .Z(n234));
Q_MX02 U234 ( .S(seed_entry[0]), .A0(\seed[0][198] ), .A1(\seed[1][198] ), .Z(n235));
Q_MX02 U235 ( .S(seed_entry[0]), .A0(\seed[0][197] ), .A1(\seed[1][197] ), .Z(n236));
Q_MX02 U236 ( .S(seed_entry[0]), .A0(\seed[0][196] ), .A1(\seed[1][196] ), .Z(n237));
Q_MX02 U237 ( .S(seed_entry[0]), .A0(\seed[0][195] ), .A1(\seed[1][195] ), .Z(n238));
Q_MX02 U238 ( .S(seed_entry[0]), .A0(\seed[0][194] ), .A1(\seed[1][194] ), .Z(n239));
Q_MX02 U239 ( .S(seed_entry[0]), .A0(\seed[0][193] ), .A1(\seed[1][193] ), .Z(n240));
Q_MX02 U240 ( .S(seed_entry[0]), .A0(\seed[0][192] ), .A1(\seed[1][192] ), .Z(n241));
Q_MX02 U241 ( .S(seed_entry[0]), .A0(\seed[0][191] ), .A1(\seed[1][191] ), .Z(n242));
Q_MX02 U242 ( .S(seed_entry[0]), .A0(\seed[0][190] ), .A1(\seed[1][190] ), .Z(n243));
Q_MX02 U243 ( .S(seed_entry[0]), .A0(\seed[0][189] ), .A1(\seed[1][189] ), .Z(n244));
Q_MX02 U244 ( .S(seed_entry[0]), .A0(\seed[0][188] ), .A1(\seed[1][188] ), .Z(n245));
Q_MX02 U245 ( .S(seed_entry[0]), .A0(\seed[0][187] ), .A1(\seed[1][187] ), .Z(n246));
Q_MX02 U246 ( .S(seed_entry[0]), .A0(\seed[0][186] ), .A1(\seed[1][186] ), .Z(n247));
Q_MX02 U247 ( .S(seed_entry[0]), .A0(\seed[0][185] ), .A1(\seed[1][185] ), .Z(n248));
Q_MX02 U248 ( .S(seed_entry[0]), .A0(\seed[0][184] ), .A1(\seed[1][184] ), .Z(n249));
Q_MX02 U249 ( .S(seed_entry[0]), .A0(\seed[0][183] ), .A1(\seed[1][183] ), .Z(n250));
Q_MX02 U250 ( .S(seed_entry[0]), .A0(\seed[0][182] ), .A1(\seed[1][182] ), .Z(n251));
Q_MX02 U251 ( .S(seed_entry[0]), .A0(\seed[0][181] ), .A1(\seed[1][181] ), .Z(n252));
Q_MX02 U252 ( .S(seed_entry[0]), .A0(\seed[0][180] ), .A1(\seed[1][180] ), .Z(n253));
Q_MX02 U253 ( .S(seed_entry[0]), .A0(\seed[0][179] ), .A1(\seed[1][179] ), .Z(n254));
Q_MX02 U254 ( .S(seed_entry[0]), .A0(\seed[0][178] ), .A1(\seed[1][178] ), .Z(n255));
Q_MX02 U255 ( .S(seed_entry[0]), .A0(\seed[0][177] ), .A1(\seed[1][177] ), .Z(n256));
Q_MX02 U256 ( .S(seed_entry[0]), .A0(\seed[0][176] ), .A1(\seed[1][176] ), .Z(n257));
Q_MX02 U257 ( .S(seed_entry[0]), .A0(\seed[0][175] ), .A1(\seed[1][175] ), .Z(n258));
Q_MX02 U258 ( .S(seed_entry[0]), .A0(\seed[0][174] ), .A1(\seed[1][174] ), .Z(n259));
Q_MX02 U259 ( .S(seed_entry[0]), .A0(\seed[0][173] ), .A1(\seed[1][173] ), .Z(n260));
Q_MX02 U260 ( .S(seed_entry[0]), .A0(\seed[0][172] ), .A1(\seed[1][172] ), .Z(n261));
Q_MX02 U261 ( .S(seed_entry[0]), .A0(\seed[0][171] ), .A1(\seed[1][171] ), .Z(n262));
Q_MX02 U262 ( .S(seed_entry[0]), .A0(\seed[0][170] ), .A1(\seed[1][170] ), .Z(n263));
Q_MX02 U263 ( .S(seed_entry[0]), .A0(\seed[0][169] ), .A1(\seed[1][169] ), .Z(n264));
Q_MX02 U264 ( .S(seed_entry[0]), .A0(\seed[0][168] ), .A1(\seed[1][168] ), .Z(n265));
Q_MX02 U265 ( .S(seed_entry[0]), .A0(\seed[0][167] ), .A1(\seed[1][167] ), .Z(n266));
Q_MX02 U266 ( .S(seed_entry[0]), .A0(\seed[0][166] ), .A1(\seed[1][166] ), .Z(n267));
Q_MX02 U267 ( .S(seed_entry[0]), .A0(\seed[0][165] ), .A1(\seed[1][165] ), .Z(n268));
Q_MX02 U268 ( .S(seed_entry[0]), .A0(\seed[0][164] ), .A1(\seed[1][164] ), .Z(n269));
Q_MX02 U269 ( .S(seed_entry[0]), .A0(\seed[0][163] ), .A1(\seed[1][163] ), .Z(n270));
Q_MX02 U270 ( .S(seed_entry[0]), .A0(\seed[0][162] ), .A1(\seed[1][162] ), .Z(n271));
Q_MX02 U271 ( .S(seed_entry[0]), .A0(\seed[0][161] ), .A1(\seed[1][161] ), .Z(n272));
Q_MX02 U272 ( .S(seed_entry[0]), .A0(\seed[0][160] ), .A1(\seed[1][160] ), .Z(n273));
Q_MX02 U273 ( .S(seed_entry[0]), .A0(\seed[0][159] ), .A1(\seed[1][159] ), .Z(n274));
Q_MX02 U274 ( .S(seed_entry[0]), .A0(\seed[0][158] ), .A1(\seed[1][158] ), .Z(n275));
Q_MX02 U275 ( .S(seed_entry[0]), .A0(\seed[0][157] ), .A1(\seed[1][157] ), .Z(n276));
Q_MX02 U276 ( .S(seed_entry[0]), .A0(\seed[0][156] ), .A1(\seed[1][156] ), .Z(n277));
Q_MX02 U277 ( .S(seed_entry[0]), .A0(\seed[0][155] ), .A1(\seed[1][155] ), .Z(n278));
Q_MX02 U278 ( .S(seed_entry[0]), .A0(\seed[0][154] ), .A1(\seed[1][154] ), .Z(n279));
Q_MX02 U279 ( .S(seed_entry[0]), .A0(\seed[0][153] ), .A1(\seed[1][153] ), .Z(n280));
Q_MX02 U280 ( .S(seed_entry[0]), .A0(\seed[0][152] ), .A1(\seed[1][152] ), .Z(n281));
Q_MX02 U281 ( .S(seed_entry[0]), .A0(\seed[0][151] ), .A1(\seed[1][151] ), .Z(n282));
Q_MX02 U282 ( .S(seed_entry[0]), .A0(\seed[0][150] ), .A1(\seed[1][150] ), .Z(n283));
Q_MX02 U283 ( .S(seed_entry[0]), .A0(\seed[0][149] ), .A1(\seed[1][149] ), .Z(n284));
Q_MX02 U284 ( .S(seed_entry[0]), .A0(\seed[0][148] ), .A1(\seed[1][148] ), .Z(n285));
Q_MX02 U285 ( .S(seed_entry[0]), .A0(\seed[0][147] ), .A1(\seed[1][147] ), .Z(n286));
Q_MX02 U286 ( .S(seed_entry[0]), .A0(\seed[0][146] ), .A1(\seed[1][146] ), .Z(n287));
Q_MX02 U287 ( .S(seed_entry[0]), .A0(\seed[0][145] ), .A1(\seed[1][145] ), .Z(n288));
Q_MX02 U288 ( .S(seed_entry[0]), .A0(\seed[0][144] ), .A1(\seed[1][144] ), .Z(n289));
Q_MX02 U289 ( .S(seed_entry[0]), .A0(\seed[0][143] ), .A1(\seed[1][143] ), .Z(n290));
Q_MX02 U290 ( .S(seed_entry[0]), .A0(\seed[0][142] ), .A1(\seed[1][142] ), .Z(n291));
Q_MX02 U291 ( .S(seed_entry[0]), .A0(\seed[0][141] ), .A1(\seed[1][141] ), .Z(n292));
Q_MX02 U292 ( .S(seed_entry[0]), .A0(\seed[0][140] ), .A1(\seed[1][140] ), .Z(n293));
Q_MX02 U293 ( .S(seed_entry[0]), .A0(\seed[0][139] ), .A1(\seed[1][139] ), .Z(n294));
Q_MX02 U294 ( .S(seed_entry[0]), .A0(\seed[0][138] ), .A1(\seed[1][138] ), .Z(n295));
Q_MX02 U295 ( .S(seed_entry[0]), .A0(\seed[0][137] ), .A1(\seed[1][137] ), .Z(n296));
Q_MX02 U296 ( .S(seed_entry[0]), .A0(\seed[0][136] ), .A1(\seed[1][136] ), .Z(n297));
Q_MX02 U297 ( .S(seed_entry[0]), .A0(\seed[0][135] ), .A1(\seed[1][135] ), .Z(n298));
Q_MX02 U298 ( .S(seed_entry[0]), .A0(\seed[0][134] ), .A1(\seed[1][134] ), .Z(n299));
Q_MX02 U299 ( .S(seed_entry[0]), .A0(\seed[0][133] ), .A1(\seed[1][133] ), .Z(n300));
Q_MX02 U300 ( .S(seed_entry[0]), .A0(\seed[0][132] ), .A1(\seed[1][132] ), .Z(n301));
Q_MX02 U301 ( .S(seed_entry[0]), .A0(\seed[0][131] ), .A1(\seed[1][131] ), .Z(n302));
Q_MX02 U302 ( .S(seed_entry[0]), .A0(\seed[0][130] ), .A1(\seed[1][130] ), .Z(n303));
Q_MX02 U303 ( .S(seed_entry[0]), .A0(\seed[0][129] ), .A1(\seed[1][129] ), .Z(n304));
Q_MX02 U304 ( .S(seed_entry[0]), .A0(\seed[0][128] ), .A1(\seed[1][128] ), .Z(n305));
Q_MX02 U305 ( .S(seed_entry[0]), .A0(\seed[0][127] ), .A1(\seed[1][127] ), .Z(n306));
Q_MX02 U306 ( .S(seed_entry[0]), .A0(\seed[0][126] ), .A1(\seed[1][126] ), .Z(n307));
Q_MX02 U307 ( .S(seed_entry[0]), .A0(\seed[0][125] ), .A1(\seed[1][125] ), .Z(n308));
Q_MX02 U308 ( .S(seed_entry[0]), .A0(\seed[0][124] ), .A1(\seed[1][124] ), .Z(n309));
Q_MX02 U309 ( .S(seed_entry[0]), .A0(\seed[0][123] ), .A1(\seed[1][123] ), .Z(n310));
Q_MX02 U310 ( .S(seed_entry[0]), .A0(\seed[0][122] ), .A1(\seed[1][122] ), .Z(n311));
Q_MX02 U311 ( .S(seed_entry[0]), .A0(\seed[0][121] ), .A1(\seed[1][121] ), .Z(n312));
Q_MX02 U312 ( .S(seed_entry[0]), .A0(\seed[0][120] ), .A1(\seed[1][120] ), .Z(n313));
Q_MX02 U313 ( .S(seed_entry[0]), .A0(\seed[0][119] ), .A1(\seed[1][119] ), .Z(n314));
Q_MX02 U314 ( .S(seed_entry[0]), .A0(\seed[0][118] ), .A1(\seed[1][118] ), .Z(n315));
Q_MX02 U315 ( .S(seed_entry[0]), .A0(\seed[0][117] ), .A1(\seed[1][117] ), .Z(n316));
Q_MX02 U316 ( .S(seed_entry[0]), .A0(\seed[0][116] ), .A1(\seed[1][116] ), .Z(n317));
Q_MX02 U317 ( .S(seed_entry[0]), .A0(\seed[0][115] ), .A1(\seed[1][115] ), .Z(n318));
Q_MX02 U318 ( .S(seed_entry[0]), .A0(\seed[0][114] ), .A1(\seed[1][114] ), .Z(n319));
Q_MX02 U319 ( .S(seed_entry[0]), .A0(\seed[0][113] ), .A1(\seed[1][113] ), .Z(n320));
Q_MX02 U320 ( .S(seed_entry[0]), .A0(\seed[0][112] ), .A1(\seed[1][112] ), .Z(n321));
Q_MX02 U321 ( .S(seed_entry[0]), .A0(\seed[0][111] ), .A1(\seed[1][111] ), .Z(n322));
Q_MX02 U322 ( .S(seed_entry[0]), .A0(\seed[0][110] ), .A1(\seed[1][110] ), .Z(n323));
Q_MX02 U323 ( .S(seed_entry[0]), .A0(\seed[0][109] ), .A1(\seed[1][109] ), .Z(n324));
Q_MX02 U324 ( .S(seed_entry[0]), .A0(\seed[0][108] ), .A1(\seed[1][108] ), .Z(n325));
Q_MX02 U325 ( .S(seed_entry[0]), .A0(\seed[0][107] ), .A1(\seed[1][107] ), .Z(n326));
Q_MX02 U326 ( .S(seed_entry[0]), .A0(\seed[0][106] ), .A1(\seed[1][106] ), .Z(n327));
Q_MX02 U327 ( .S(seed_entry[0]), .A0(\seed[0][105] ), .A1(\seed[1][105] ), .Z(n328));
Q_MX02 U328 ( .S(seed_entry[0]), .A0(\seed[0][104] ), .A1(\seed[1][104] ), .Z(n329));
Q_MX02 U329 ( .S(seed_entry[0]), .A0(\seed[0][103] ), .A1(\seed[1][103] ), .Z(n330));
Q_MX02 U330 ( .S(seed_entry[0]), .A0(\seed[0][102] ), .A1(\seed[1][102] ), .Z(n331));
Q_MX02 U331 ( .S(seed_entry[0]), .A0(\seed[0][101] ), .A1(\seed[1][101] ), .Z(n332));
Q_MX02 U332 ( .S(seed_entry[0]), .A0(\seed[0][100] ), .A1(\seed[1][100] ), .Z(n333));
Q_MX02 U333 ( .S(seed_entry[0]), .A0(\seed[0][99] ), .A1(\seed[1][99] ), .Z(n334));
Q_MX02 U334 ( .S(seed_entry[0]), .A0(\seed[0][98] ), .A1(\seed[1][98] ), .Z(n335));
Q_MX02 U335 ( .S(seed_entry[0]), .A0(\seed[0][97] ), .A1(\seed[1][97] ), .Z(n336));
Q_MX02 U336 ( .S(seed_entry[0]), .A0(\seed[0][96] ), .A1(\seed[1][96] ), .Z(n337));
Q_MX02 U337 ( .S(seed_entry[0]), .A0(\seed[0][95] ), .A1(\seed[1][95] ), .Z(n338));
Q_MX02 U338 ( .S(seed_entry[0]), .A0(\seed[0][94] ), .A1(\seed[1][94] ), .Z(n339));
Q_MX02 U339 ( .S(seed_entry[0]), .A0(\seed[0][93] ), .A1(\seed[1][93] ), .Z(n340));
Q_MX02 U340 ( .S(seed_entry[0]), .A0(\seed[0][92] ), .A1(\seed[1][92] ), .Z(n341));
Q_MX02 U341 ( .S(seed_entry[0]), .A0(\seed[0][91] ), .A1(\seed[1][91] ), .Z(n342));
Q_MX02 U342 ( .S(seed_entry[0]), .A0(\seed[0][90] ), .A1(\seed[1][90] ), .Z(n343));
Q_MX02 U343 ( .S(seed_entry[0]), .A0(\seed[0][89] ), .A1(\seed[1][89] ), .Z(n344));
Q_MX02 U344 ( .S(seed_entry[0]), .A0(\seed[0][88] ), .A1(\seed[1][88] ), .Z(n345));
Q_MX02 U345 ( .S(seed_entry[0]), .A0(\seed[0][87] ), .A1(\seed[1][87] ), .Z(n346));
Q_MX02 U346 ( .S(seed_entry[0]), .A0(\seed[0][86] ), .A1(\seed[1][86] ), .Z(n347));
Q_MX02 U347 ( .S(seed_entry[0]), .A0(\seed[0][85] ), .A1(\seed[1][85] ), .Z(n348));
Q_MX02 U348 ( .S(seed_entry[0]), .A0(\seed[0][84] ), .A1(\seed[1][84] ), .Z(n349));
Q_MX02 U349 ( .S(seed_entry[0]), .A0(\seed[0][83] ), .A1(\seed[1][83] ), .Z(n350));
Q_MX02 U350 ( .S(seed_entry[0]), .A0(\seed[0][82] ), .A1(\seed[1][82] ), .Z(n351));
Q_MX02 U351 ( .S(seed_entry[0]), .A0(\seed[0][81] ), .A1(\seed[1][81] ), .Z(n352));
Q_MX02 U352 ( .S(seed_entry[0]), .A0(\seed[0][80] ), .A1(\seed[1][80] ), .Z(n353));
Q_MX02 U353 ( .S(seed_entry[0]), .A0(\seed[0][79] ), .A1(\seed[1][79] ), .Z(n354));
Q_MX02 U354 ( .S(seed_entry[0]), .A0(\seed[0][78] ), .A1(\seed[1][78] ), .Z(n355));
Q_MX02 U355 ( .S(seed_entry[0]), .A0(\seed[0][77] ), .A1(\seed[1][77] ), .Z(n356));
Q_MX02 U356 ( .S(seed_entry[0]), .A0(\seed[0][76] ), .A1(\seed[1][76] ), .Z(n357));
Q_MX02 U357 ( .S(seed_entry[0]), .A0(\seed[0][75] ), .A1(\seed[1][75] ), .Z(n358));
Q_MX02 U358 ( .S(seed_entry[0]), .A0(\seed[0][74] ), .A1(\seed[1][74] ), .Z(n359));
Q_MX02 U359 ( .S(seed_entry[0]), .A0(\seed[0][73] ), .A1(\seed[1][73] ), .Z(n360));
Q_MX02 U360 ( .S(seed_entry[0]), .A0(\seed[0][72] ), .A1(\seed[1][72] ), .Z(n361));
Q_MX02 U361 ( .S(seed_entry[0]), .A0(\seed[0][71] ), .A1(\seed[1][71] ), .Z(n362));
Q_MX02 U362 ( .S(seed_entry[0]), .A0(\seed[0][70] ), .A1(\seed[1][70] ), .Z(n363));
Q_MX02 U363 ( .S(seed_entry[0]), .A0(\seed[0][69] ), .A1(\seed[1][69] ), .Z(n364));
Q_MX02 U364 ( .S(seed_entry[0]), .A0(\seed[0][68] ), .A1(\seed[1][68] ), .Z(n365));
Q_MX02 U365 ( .S(seed_entry[0]), .A0(\seed[0][67] ), .A1(\seed[1][67] ), .Z(n366));
Q_MX02 U366 ( .S(seed_entry[0]), .A0(\seed[0][66] ), .A1(\seed[1][66] ), .Z(n367));
Q_MX02 U367 ( .S(seed_entry[0]), .A0(\seed[0][65] ), .A1(\seed[1][65] ), .Z(n368));
Q_MX02 U368 ( .S(seed_entry[0]), .A0(\seed[0][64] ), .A1(\seed[1][64] ), .Z(n369));
Q_MX02 U369 ( .S(seed_entry[0]), .A0(\seed[0][63] ), .A1(\seed[1][63] ), .Z(n370));
Q_MX02 U370 ( .S(seed_entry[0]), .A0(\seed[0][62] ), .A1(\seed[1][62] ), .Z(n371));
Q_MX02 U371 ( .S(seed_entry[0]), .A0(\seed[0][61] ), .A1(\seed[1][61] ), .Z(n372));
Q_MX02 U372 ( .S(seed_entry[0]), .A0(\seed[0][60] ), .A1(\seed[1][60] ), .Z(n373));
Q_MX02 U373 ( .S(seed_entry[0]), .A0(\seed[0][59] ), .A1(\seed[1][59] ), .Z(n374));
Q_MX02 U374 ( .S(seed_entry[0]), .A0(\seed[0][58] ), .A1(\seed[1][58] ), .Z(n375));
Q_MX02 U375 ( .S(seed_entry[0]), .A0(\seed[0][57] ), .A1(\seed[1][57] ), .Z(n376));
Q_MX02 U376 ( .S(seed_entry[0]), .A0(\seed[0][56] ), .A1(\seed[1][56] ), .Z(n377));
Q_MX02 U377 ( .S(seed_entry[0]), .A0(\seed[0][55] ), .A1(\seed[1][55] ), .Z(n378));
Q_MX02 U378 ( .S(seed_entry[0]), .A0(\seed[0][54] ), .A1(\seed[1][54] ), .Z(n379));
Q_MX02 U379 ( .S(seed_entry[0]), .A0(\seed[0][53] ), .A1(\seed[1][53] ), .Z(n380));
Q_MX02 U380 ( .S(seed_entry[0]), .A0(\seed[0][52] ), .A1(\seed[1][52] ), .Z(n381));
Q_MX02 U381 ( .S(seed_entry[0]), .A0(\seed[0][51] ), .A1(\seed[1][51] ), .Z(n382));
Q_MX02 U382 ( .S(seed_entry[0]), .A0(\seed[0][50] ), .A1(\seed[1][50] ), .Z(n383));
Q_MX02 U383 ( .S(seed_entry[0]), .A0(\seed[0][49] ), .A1(\seed[1][49] ), .Z(n384));
Q_MX02 U384 ( .S(seed_entry[0]), .A0(\seed[0][48] ), .A1(\seed[1][48] ), .Z(n385));
Q_MX02 U385 ( .S(seed_entry[0]), .A0(\seed[0][47] ), .A1(\seed[1][47] ), .Z(n386));
Q_MX02 U386 ( .S(seed_entry[0]), .A0(\seed[0][46] ), .A1(\seed[1][46] ), .Z(n387));
Q_MX02 U387 ( .S(seed_entry[0]), .A0(\seed[0][45] ), .A1(\seed[1][45] ), .Z(n388));
Q_MX02 U388 ( .S(seed_entry[0]), .A0(\seed[0][44] ), .A1(\seed[1][44] ), .Z(n389));
Q_MX02 U389 ( .S(seed_entry[0]), .A0(\seed[0][43] ), .A1(\seed[1][43] ), .Z(n390));
Q_MX02 U390 ( .S(seed_entry[0]), .A0(\seed[0][42] ), .A1(\seed[1][42] ), .Z(n391));
Q_MX02 U391 ( .S(seed_entry[0]), .A0(\seed[0][41] ), .A1(\seed[1][41] ), .Z(n392));
Q_MX02 U392 ( .S(seed_entry[0]), .A0(\seed[0][40] ), .A1(\seed[1][40] ), .Z(n393));
Q_MX02 U393 ( .S(seed_entry[0]), .A0(\seed[0][39] ), .A1(\seed[1][39] ), .Z(n394));
Q_MX02 U394 ( .S(seed_entry[0]), .A0(\seed[0][38] ), .A1(\seed[1][38] ), .Z(n395));
Q_MX02 U395 ( .S(seed_entry[0]), .A0(\seed[0][37] ), .A1(\seed[1][37] ), .Z(n396));
Q_MX02 U396 ( .S(seed_entry[0]), .A0(\seed[0][36] ), .A1(\seed[1][36] ), .Z(n397));
Q_MX02 U397 ( .S(seed_entry[0]), .A0(\seed[0][35] ), .A1(\seed[1][35] ), .Z(n398));
Q_MX02 U398 ( .S(seed_entry[0]), .A0(\seed[0][34] ), .A1(\seed[1][34] ), .Z(n399));
Q_MX02 U399 ( .S(seed_entry[0]), .A0(\seed[0][33] ), .A1(\seed[1][33] ), .Z(n400));
Q_MX02 U400 ( .S(seed_entry[0]), .A0(\seed[0][32] ), .A1(\seed[1][32] ), .Z(n401));
Q_MX02 U401 ( .S(seed_entry[0]), .A0(\seed[0][31] ), .A1(\seed[1][31] ), .Z(n402));
Q_MX02 U402 ( .S(seed_entry[0]), .A0(\seed[0][30] ), .A1(\seed[1][30] ), .Z(n403));
Q_MX02 U403 ( .S(seed_entry[0]), .A0(\seed[0][29] ), .A1(\seed[1][29] ), .Z(n404));
Q_MX02 U404 ( .S(seed_entry[0]), .A0(\seed[0][28] ), .A1(\seed[1][28] ), .Z(n405));
Q_MX02 U405 ( .S(seed_entry[0]), .A0(\seed[0][27] ), .A1(\seed[1][27] ), .Z(n406));
Q_MX02 U406 ( .S(seed_entry[0]), .A0(\seed[0][26] ), .A1(\seed[1][26] ), .Z(n407));
Q_MX02 U407 ( .S(seed_entry[0]), .A0(\seed[0][25] ), .A1(\seed[1][25] ), .Z(n408));
Q_MX02 U408 ( .S(seed_entry[0]), .A0(\seed[0][24] ), .A1(\seed[1][24] ), .Z(n409));
Q_MX02 U409 ( .S(seed_entry[0]), .A0(\seed[0][23] ), .A1(\seed[1][23] ), .Z(n410));
Q_MX02 U410 ( .S(seed_entry[0]), .A0(\seed[0][22] ), .A1(\seed[1][22] ), .Z(n411));
Q_MX02 U411 ( .S(seed_entry[0]), .A0(\seed[0][21] ), .A1(\seed[1][21] ), .Z(n412));
Q_MX02 U412 ( .S(seed_entry[0]), .A0(\seed[0][20] ), .A1(\seed[1][20] ), .Z(n413));
Q_MX02 U413 ( .S(seed_entry[0]), .A0(\seed[0][19] ), .A1(\seed[1][19] ), .Z(n414));
Q_MX02 U414 ( .S(seed_entry[0]), .A0(\seed[0][18] ), .A1(\seed[1][18] ), .Z(n415));
Q_MX02 U415 ( .S(seed_entry[0]), .A0(\seed[0][17] ), .A1(\seed[1][17] ), .Z(n416));
Q_MX02 U416 ( .S(seed_entry[0]), .A0(\seed[0][16] ), .A1(\seed[1][16] ), .Z(n417));
Q_MX02 U417 ( .S(seed_entry[0]), .A0(\seed[0][15] ), .A1(\seed[1][15] ), .Z(n418));
Q_MX02 U418 ( .S(seed_entry[0]), .A0(\seed[0][14] ), .A1(\seed[1][14] ), .Z(n419));
Q_MX02 U419 ( .S(seed_entry[0]), .A0(\seed[0][13] ), .A1(\seed[1][13] ), .Z(n420));
Q_MX02 U420 ( .S(seed_entry[0]), .A0(\seed[0][12] ), .A1(\seed[1][12] ), .Z(n421));
Q_MX02 U421 ( .S(seed_entry[0]), .A0(\seed[0][11] ), .A1(\seed[1][11] ), .Z(n422));
Q_MX02 U422 ( .S(seed_entry[0]), .A0(\seed[0][10] ), .A1(\seed[1][10] ), .Z(n423));
Q_MX02 U423 ( .S(seed_entry[0]), .A0(\seed[0][9] ), .A1(\seed[1][9] ), .Z(n424));
Q_MX02 U424 ( .S(seed_entry[0]), .A0(\seed[0][8] ), .A1(\seed[1][8] ), .Z(n425));
Q_MX02 U425 ( .S(seed_entry[0]), .A0(\seed[0][7] ), .A1(\seed[1][7] ), .Z(n426));
Q_MX02 U426 ( .S(seed_entry[0]), .A0(\seed[0][6] ), .A1(\seed[1][6] ), .Z(n427));
Q_MX02 U427 ( .S(seed_entry[0]), .A0(\seed[0][5] ), .A1(\seed[1][5] ), .Z(n428));
Q_MX02 U428 ( .S(seed_entry[0]), .A0(\seed[0][4] ), .A1(\seed[1][4] ), .Z(n429));
Q_MX02 U429 ( .S(seed_entry[0]), .A0(\seed[0][3] ), .A1(\seed[1][3] ), .Z(n430));
Q_MX02 U430 ( .S(seed_entry[0]), .A0(\seed[0][2] ), .A1(\seed[1][2] ), .Z(n431));
Q_MX02 U431 ( .S(seed_entry[0]), .A0(\seed[0][1] ), .A1(\seed[1][1] ), .Z(n432));
Q_MX02 U432 ( .S(seed_entry[0]), .A0(\seed[0][0] ), .A1(\seed[1][0] ), .Z(n433));
Q_INV U433 ( .A(drng_health_test), .Z(n434));
Q_AN02 U434 ( .A0(n434), .A1(drng_256_out_pre[127]), .Z(drng_256_out[127]));
Q_AN02 U435 ( .A0(n434), .A1(drng_256_out_pre[126]), .Z(drng_256_out[126]));
Q_AN02 U436 ( .A0(n434), .A1(drng_256_out_pre[125]), .Z(drng_256_out[125]));
Q_AN02 U437 ( .A0(n434), .A1(drng_256_out_pre[124]), .Z(drng_256_out[124]));
Q_AN02 U438 ( .A0(n434), .A1(drng_256_out_pre[123]), .Z(drng_256_out[123]));
Q_AN02 U439 ( .A0(n434), .A1(drng_256_out_pre[122]), .Z(drng_256_out[122]));
Q_AN02 U440 ( .A0(n434), .A1(drng_256_out_pre[121]), .Z(drng_256_out[121]));
Q_AN02 U441 ( .A0(n434), .A1(drng_256_out_pre[120]), .Z(drng_256_out[120]));
Q_AN02 U442 ( .A0(n434), .A1(drng_256_out_pre[119]), .Z(drng_256_out[119]));
Q_AN02 U443 ( .A0(n434), .A1(drng_256_out_pre[118]), .Z(drng_256_out[118]));
Q_AN02 U444 ( .A0(n434), .A1(drng_256_out_pre[117]), .Z(drng_256_out[117]));
Q_AN02 U445 ( .A0(n434), .A1(drng_256_out_pre[116]), .Z(drng_256_out[116]));
Q_AN02 U446 ( .A0(n434), .A1(drng_256_out_pre[115]), .Z(drng_256_out[115]));
Q_AN02 U447 ( .A0(n434), .A1(drng_256_out_pre[114]), .Z(drng_256_out[114]));
Q_AN02 U448 ( .A0(n434), .A1(drng_256_out_pre[113]), .Z(drng_256_out[113]));
Q_AN02 U449 ( .A0(n434), .A1(drng_256_out_pre[112]), .Z(drng_256_out[112]));
Q_AN02 U450 ( .A0(n434), .A1(drng_256_out_pre[111]), .Z(drng_256_out[111]));
Q_AN02 U451 ( .A0(n434), .A1(drng_256_out_pre[110]), .Z(drng_256_out[110]));
Q_AN02 U452 ( .A0(n434), .A1(drng_256_out_pre[109]), .Z(drng_256_out[109]));
Q_AN02 U453 ( .A0(n434), .A1(drng_256_out_pre[108]), .Z(drng_256_out[108]));
Q_AN02 U454 ( .A0(n434), .A1(drng_256_out_pre[107]), .Z(drng_256_out[107]));
Q_AN02 U455 ( .A0(n434), .A1(drng_256_out_pre[106]), .Z(drng_256_out[106]));
Q_AN02 U456 ( .A0(n434), .A1(drng_256_out_pre[105]), .Z(drng_256_out[105]));
Q_AN02 U457 ( .A0(n434), .A1(drng_256_out_pre[104]), .Z(drng_256_out[104]));
Q_AN02 U458 ( .A0(n434), .A1(drng_256_out_pre[103]), .Z(drng_256_out[103]));
Q_AN02 U459 ( .A0(n434), .A1(drng_256_out_pre[102]), .Z(drng_256_out[102]));
Q_AN02 U460 ( .A0(n434), .A1(drng_256_out_pre[101]), .Z(drng_256_out[101]));
Q_AN02 U461 ( .A0(n434), .A1(drng_256_out_pre[100]), .Z(drng_256_out[100]));
Q_AN02 U462 ( .A0(n434), .A1(drng_256_out_pre[99]), .Z(drng_256_out[99]));
Q_AN02 U463 ( .A0(n434), .A1(drng_256_out_pre[98]), .Z(drng_256_out[98]));
Q_AN02 U464 ( .A0(n434), .A1(drng_256_out_pre[97]), .Z(drng_256_out[97]));
Q_AN02 U465 ( .A0(n434), .A1(drng_256_out_pre[96]), .Z(drng_256_out[96]));
Q_AN02 U466 ( .A0(n434), .A1(drng_256_out_pre[95]), .Z(drng_256_out[95]));
Q_AN02 U467 ( .A0(n434), .A1(drng_256_out_pre[94]), .Z(drng_256_out[94]));
Q_AN02 U468 ( .A0(n434), .A1(drng_256_out_pre[93]), .Z(drng_256_out[93]));
Q_AN02 U469 ( .A0(n434), .A1(drng_256_out_pre[92]), .Z(drng_256_out[92]));
Q_AN02 U470 ( .A0(n434), .A1(drng_256_out_pre[91]), .Z(drng_256_out[91]));
Q_AN02 U471 ( .A0(n434), .A1(drng_256_out_pre[90]), .Z(drng_256_out[90]));
Q_AN02 U472 ( .A0(n434), .A1(drng_256_out_pre[89]), .Z(drng_256_out[89]));
Q_AN02 U473 ( .A0(n434), .A1(drng_256_out_pre[88]), .Z(drng_256_out[88]));
Q_AN02 U474 ( .A0(n434), .A1(drng_256_out_pre[87]), .Z(drng_256_out[87]));
Q_AN02 U475 ( .A0(n434), .A1(drng_256_out_pre[86]), .Z(drng_256_out[86]));
Q_AN02 U476 ( .A0(n434), .A1(drng_256_out_pre[85]), .Z(drng_256_out[85]));
Q_AN02 U477 ( .A0(n434), .A1(drng_256_out_pre[84]), .Z(drng_256_out[84]));
Q_AN02 U478 ( .A0(n434), .A1(drng_256_out_pre[83]), .Z(drng_256_out[83]));
Q_AN02 U479 ( .A0(n434), .A1(drng_256_out_pre[82]), .Z(drng_256_out[82]));
Q_AN02 U480 ( .A0(n434), .A1(drng_256_out_pre[81]), .Z(drng_256_out[81]));
Q_AN02 U481 ( .A0(n434), .A1(drng_256_out_pre[80]), .Z(drng_256_out[80]));
Q_AN02 U482 ( .A0(n434), .A1(drng_256_out_pre[79]), .Z(drng_256_out[79]));
Q_AN02 U483 ( .A0(n434), .A1(drng_256_out_pre[78]), .Z(drng_256_out[78]));
Q_AN02 U484 ( .A0(n434), .A1(drng_256_out_pre[77]), .Z(drng_256_out[77]));
Q_AN02 U485 ( .A0(n434), .A1(drng_256_out_pre[76]), .Z(drng_256_out[76]));
Q_AN02 U486 ( .A0(n434), .A1(drng_256_out_pre[75]), .Z(drng_256_out[75]));
Q_AN02 U487 ( .A0(n434), .A1(drng_256_out_pre[74]), .Z(drng_256_out[74]));
Q_AN02 U488 ( .A0(n434), .A1(drng_256_out_pre[73]), .Z(drng_256_out[73]));
Q_AN02 U489 ( .A0(n434), .A1(drng_256_out_pre[72]), .Z(drng_256_out[72]));
Q_AN02 U490 ( .A0(n434), .A1(drng_256_out_pre[71]), .Z(drng_256_out[71]));
Q_AN02 U491 ( .A0(n434), .A1(drng_256_out_pre[70]), .Z(drng_256_out[70]));
Q_AN02 U492 ( .A0(n434), .A1(drng_256_out_pre[69]), .Z(drng_256_out[69]));
Q_AN02 U493 ( .A0(n434), .A1(drng_256_out_pre[68]), .Z(drng_256_out[68]));
Q_AN02 U494 ( .A0(n434), .A1(drng_256_out_pre[67]), .Z(drng_256_out[67]));
Q_AN02 U495 ( .A0(n434), .A1(drng_256_out_pre[66]), .Z(drng_256_out[66]));
Q_AN02 U496 ( .A0(n434), .A1(drng_256_out_pre[65]), .Z(drng_256_out[65]));
Q_AN02 U497 ( .A0(n434), .A1(drng_256_out_pre[64]), .Z(drng_256_out[64]));
Q_AN02 U498 ( .A0(n434), .A1(drng_256_out_pre[63]), .Z(drng_256_out[63]));
Q_AN02 U499 ( .A0(n434), .A1(drng_256_out_pre[62]), .Z(drng_256_out[62]));
Q_AN02 U500 ( .A0(n434), .A1(drng_256_out_pre[61]), .Z(drng_256_out[61]));
Q_AN02 U501 ( .A0(n434), .A1(drng_256_out_pre[60]), .Z(drng_256_out[60]));
Q_AN02 U502 ( .A0(n434), .A1(drng_256_out_pre[59]), .Z(drng_256_out[59]));
Q_AN02 U503 ( .A0(n434), .A1(drng_256_out_pre[58]), .Z(drng_256_out[58]));
Q_AN02 U504 ( .A0(n434), .A1(drng_256_out_pre[57]), .Z(drng_256_out[57]));
Q_AN02 U505 ( .A0(n434), .A1(drng_256_out_pre[56]), .Z(drng_256_out[56]));
Q_AN02 U506 ( .A0(n434), .A1(drng_256_out_pre[55]), .Z(drng_256_out[55]));
Q_AN02 U507 ( .A0(n434), .A1(drng_256_out_pre[54]), .Z(drng_256_out[54]));
Q_AN02 U508 ( .A0(n434), .A1(drng_256_out_pre[53]), .Z(drng_256_out[53]));
Q_AN02 U509 ( .A0(n434), .A1(drng_256_out_pre[52]), .Z(drng_256_out[52]));
Q_AN02 U510 ( .A0(n434), .A1(drng_256_out_pre[51]), .Z(drng_256_out[51]));
Q_AN02 U511 ( .A0(n434), .A1(drng_256_out_pre[50]), .Z(drng_256_out[50]));
Q_AN02 U512 ( .A0(n434), .A1(drng_256_out_pre[49]), .Z(drng_256_out[49]));
Q_AN02 U513 ( .A0(n434), .A1(drng_256_out_pre[48]), .Z(drng_256_out[48]));
Q_AN02 U514 ( .A0(n434), .A1(drng_256_out_pre[47]), .Z(drng_256_out[47]));
Q_AN02 U515 ( .A0(n434), .A1(drng_256_out_pre[46]), .Z(drng_256_out[46]));
Q_AN02 U516 ( .A0(n434), .A1(drng_256_out_pre[45]), .Z(drng_256_out[45]));
Q_AN02 U517 ( .A0(n434), .A1(drng_256_out_pre[44]), .Z(drng_256_out[44]));
Q_AN02 U518 ( .A0(n434), .A1(drng_256_out_pre[43]), .Z(drng_256_out[43]));
Q_AN02 U519 ( .A0(n434), .A1(drng_256_out_pre[42]), .Z(drng_256_out[42]));
Q_AN02 U520 ( .A0(n434), .A1(drng_256_out_pre[41]), .Z(drng_256_out[41]));
Q_AN02 U521 ( .A0(n434), .A1(drng_256_out_pre[40]), .Z(drng_256_out[40]));
Q_AN02 U522 ( .A0(n434), .A1(drng_256_out_pre[39]), .Z(drng_256_out[39]));
Q_AN02 U523 ( .A0(n434), .A1(drng_256_out_pre[38]), .Z(drng_256_out[38]));
Q_AN02 U524 ( .A0(n434), .A1(drng_256_out_pre[37]), .Z(drng_256_out[37]));
Q_AN02 U525 ( .A0(n434), .A1(drng_256_out_pre[36]), .Z(drng_256_out[36]));
Q_AN02 U526 ( .A0(n434), .A1(drng_256_out_pre[35]), .Z(drng_256_out[35]));
Q_AN02 U527 ( .A0(n434), .A1(drng_256_out_pre[34]), .Z(drng_256_out[34]));
Q_AN02 U528 ( .A0(n434), .A1(drng_256_out_pre[33]), .Z(drng_256_out[33]));
Q_AN02 U529 ( .A0(n434), .A1(drng_256_out_pre[32]), .Z(drng_256_out[32]));
Q_AN02 U530 ( .A0(n434), .A1(drng_256_out_pre[31]), .Z(drng_256_out[31]));
Q_AN02 U531 ( .A0(n434), .A1(drng_256_out_pre[30]), .Z(drng_256_out[30]));
Q_AN02 U532 ( .A0(n434), .A1(drng_256_out_pre[29]), .Z(drng_256_out[29]));
Q_AN02 U533 ( .A0(n434), .A1(drng_256_out_pre[28]), .Z(drng_256_out[28]));
Q_AN02 U534 ( .A0(n434), .A1(drng_256_out_pre[27]), .Z(drng_256_out[27]));
Q_AN02 U535 ( .A0(n434), .A1(drng_256_out_pre[26]), .Z(drng_256_out[26]));
Q_AN02 U536 ( .A0(n434), .A1(drng_256_out_pre[25]), .Z(drng_256_out[25]));
Q_AN02 U537 ( .A0(n434), .A1(drng_256_out_pre[24]), .Z(drng_256_out[24]));
Q_AN02 U538 ( .A0(n434), .A1(drng_256_out_pre[23]), .Z(drng_256_out[23]));
Q_AN02 U539 ( .A0(n434), .A1(drng_256_out_pre[22]), .Z(drng_256_out[22]));
Q_AN02 U540 ( .A0(n434), .A1(drng_256_out_pre[21]), .Z(drng_256_out[21]));
Q_AN02 U541 ( .A0(n434), .A1(drng_256_out_pre[20]), .Z(drng_256_out[20]));
Q_AN02 U542 ( .A0(n434), .A1(drng_256_out_pre[19]), .Z(drng_256_out[19]));
Q_AN02 U543 ( .A0(n434), .A1(drng_256_out_pre[18]), .Z(drng_256_out[18]));
Q_AN02 U544 ( .A0(n434), .A1(drng_256_out_pre[17]), .Z(drng_256_out[17]));
Q_AN02 U545 ( .A0(n434), .A1(drng_256_out_pre[16]), .Z(drng_256_out[16]));
Q_AN02 U546 ( .A0(n434), .A1(drng_256_out_pre[15]), .Z(drng_256_out[15]));
Q_AN02 U547 ( .A0(n434), .A1(drng_256_out_pre[14]), .Z(drng_256_out[14]));
Q_AN02 U548 ( .A0(n434), .A1(drng_256_out_pre[13]), .Z(drng_256_out[13]));
Q_AN02 U549 ( .A0(n434), .A1(drng_256_out_pre[12]), .Z(drng_256_out[12]));
Q_AN02 U550 ( .A0(n434), .A1(drng_256_out_pre[11]), .Z(drng_256_out[11]));
Q_AN02 U551 ( .A0(n434), .A1(drng_256_out_pre[10]), .Z(drng_256_out[10]));
Q_AN02 U552 ( .A0(n434), .A1(drng_256_out_pre[9]), .Z(drng_256_out[9]));
Q_AN02 U553 ( .A0(n434), .A1(drng_256_out_pre[8]), .Z(drng_256_out[8]));
Q_AN02 U554 ( .A0(n434), .A1(drng_256_out_pre[7]), .Z(drng_256_out[7]));
Q_AN02 U555 ( .A0(n434), .A1(drng_256_out_pre[6]), .Z(drng_256_out[6]));
Q_AN02 U556 ( .A0(n434), .A1(drng_256_out_pre[5]), .Z(drng_256_out[5]));
Q_AN02 U557 ( .A0(n434), .A1(drng_256_out_pre[4]), .Z(drng_256_out[4]));
Q_AN02 U558 ( .A0(n434), .A1(drng_256_out_pre[3]), .Z(drng_256_out[3]));
Q_AN02 U559 ( .A0(n434), .A1(drng_256_out_pre[2]), .Z(drng_256_out[2]));
Q_AN02 U560 ( .A0(n434), .A1(drng_256_out_pre[1]), .Z(drng_256_out[1]));
Q_AN02 U561 ( .A0(n434), .A1(drng_256_out_pre[0]), .Z(drng_256_out[0]));
Q_INV U562 ( .A(n437), .Z(n438));
Q_MX02 U563 ( .S(seed_entry[0]), .A0(seed0_invalidate), .A1(seed1_invalidate), .Z(n437));
Q_MX02 U564 ( .S(n435), .A0(drng_seed_expired), .A1(n438), .Z(n439));
Q_FDP1 \seed_entry_REG[0] ( .CK(clk), .R(rst_n), .D(n440), .Q(seed_entry[0]), .QN(n655));
Q_AN03 U566 ( .A0(n442), .A1(n441), .A2(drng_first), .Z(n436));
Q_AN03 U567 ( .A0(n445), .A1(n444), .A2(n443), .Z(n441));
Q_AN03 U568 ( .A0(n448), .A1(n447), .A2(n446), .Z(n442));
Q_AN03 U569 ( .A0(n451), .A1(n450), .A2(n449), .Z(n443));
Q_AN03 U570 ( .A0(n454), .A1(n453), .A2(n452), .Z(n444));
Q_AN03 U571 ( .A0(n457), .A1(n456), .A2(n455), .Z(n445));
Q_AN03 U572 ( .A0(n460), .A1(n459), .A2(n458), .Z(n446));
Q_AN03 U573 ( .A0(n463), .A1(n462), .A2(n461), .Z(n447));
Q_AN03 U574 ( .A0(n466), .A1(n465), .A2(n464), .Z(n448));
Q_AN03 U575 ( .A0(n469), .A1(n468), .A2(n467), .Z(n449));
Q_AN03 U576 ( .A0(n472), .A1(n471), .A2(n470), .Z(n450));
Q_AN03 U577 ( .A0(n475), .A1(n474), .A2(n473), .Z(n451));
Q_AN03 U578 ( .A0(n478), .A1(n477), .A2(n476), .Z(n452));
Q_AN03 U579 ( .A0(n481), .A1(n480), .A2(n479), .Z(n453));
Q_AN03 U580 ( .A0(n484), .A1(n483), .A2(n482), .Z(n454));
Q_AN03 U581 ( .A0(n487), .A1(n486), .A2(n485), .Z(n455));
Q_AN03 U582 ( .A0(n490), .A1(n489), .A2(n488), .Z(n456));
Q_AN03 U583 ( .A0(n493), .A1(n492), .A2(n491), .Z(n457));
Q_AN03 U584 ( .A0(n496), .A1(n495), .A2(n494), .Z(n458));
Q_AN03 U585 ( .A0(n499), .A1(n498), .A2(n497), .Z(n459));
Q_AN03 U586 ( .A0(n502), .A1(n501), .A2(n500), .Z(n460));
Q_AN03 U587 ( .A0(n630), .A1(n631), .A2(n503), .Z(n461));
Q_AN03 U588 ( .A0(n627), .A1(n628), .A2(n629), .Z(n462));
Q_AN03 U589 ( .A0(n624), .A1(n625), .A2(n626), .Z(n463));
Q_AN03 U590 ( .A0(n621), .A1(n622), .A2(n623), .Z(n464));
Q_AN03 U591 ( .A0(n618), .A1(n619), .A2(n620), .Z(n465));
Q_AN03 U592 ( .A0(n615), .A1(n616), .A2(n617), .Z(n466));
Q_AN03 U593 ( .A0(n612), .A1(n613), .A2(n614), .Z(n467));
Q_AN03 U594 ( .A0(n609), .A1(n610), .A2(n611), .Z(n468));
Q_AN03 U595 ( .A0(n606), .A1(n607), .A2(n608), .Z(n469));
Q_AN03 U596 ( .A0(n603), .A1(n604), .A2(n605), .Z(n470));
Q_AN03 U597 ( .A0(n600), .A1(n601), .A2(n602), .Z(n471));
Q_AN03 U598 ( .A0(n597), .A1(n598), .A2(n599), .Z(n472));
Q_AN03 U599 ( .A0(n594), .A1(n595), .A2(n596), .Z(n473));
Q_AN03 U600 ( .A0(n591), .A1(n592), .A2(n593), .Z(n474));
Q_AN03 U601 ( .A0(n588), .A1(n589), .A2(n590), .Z(n475));
Q_AN03 U602 ( .A0(n585), .A1(n586), .A2(n587), .Z(n476));
Q_AN03 U603 ( .A0(n582), .A1(n583), .A2(n584), .Z(n477));
Q_AN03 U604 ( .A0(n579), .A1(n580), .A2(n581), .Z(n478));
Q_AN03 U605 ( .A0(n576), .A1(n577), .A2(n578), .Z(n479));
Q_AN03 U606 ( .A0(n573), .A1(n574), .A2(n575), .Z(n480));
Q_AN03 U607 ( .A0(n570), .A1(n571), .A2(n572), .Z(n481));
Q_AN03 U608 ( .A0(n567), .A1(n568), .A2(n569), .Z(n482));
Q_AN03 U609 ( .A0(n564), .A1(n565), .A2(n566), .Z(n483));
Q_AN03 U610 ( .A0(n561), .A1(n562), .A2(n563), .Z(n484));
Q_AN03 U611 ( .A0(n558), .A1(n559), .A2(n560), .Z(n485));
Q_AN03 U612 ( .A0(n555), .A1(n556), .A2(n557), .Z(n486));
Q_AN03 U613 ( .A0(n552), .A1(n553), .A2(n554), .Z(n487));
Q_AN03 U614 ( .A0(n549), .A1(n550), .A2(n551), .Z(n488));
Q_AN03 U615 ( .A0(n546), .A1(n547), .A2(n548), .Z(n489));
Q_AN03 U616 ( .A0(n543), .A1(n544), .A2(n545), .Z(n490));
Q_AN03 U617 ( .A0(n540), .A1(n541), .A2(n542), .Z(n491));
Q_AN03 U618 ( .A0(n537), .A1(n538), .A2(n539), .Z(n492));
Q_AN03 U619 ( .A0(n534), .A1(n535), .A2(n536), .Z(n493));
Q_AN03 U620 ( .A0(n531), .A1(n532), .A2(n533), .Z(n494));
Q_AN03 U621 ( .A0(n528), .A1(n529), .A2(n530), .Z(n495));
Q_AN03 U622 ( .A0(n525), .A1(n526), .A2(n527), .Z(n496));
Q_AN03 U623 ( .A0(n522), .A1(n523), .A2(n524), .Z(n497));
Q_AN03 U624 ( .A0(n519), .A1(n520), .A2(n521), .Z(n498));
Q_AN03 U625 ( .A0(n516), .A1(n517), .A2(n518), .Z(n499));
Q_AN03 U626 ( .A0(n513), .A1(n514), .A2(n515), .Z(n500));
Q_AN03 U627 ( .A0(n510), .A1(n511), .A2(n512), .Z(n501));
Q_AN03 U628 ( .A0(n507), .A1(n508), .A2(n509), .Z(n502));
Q_AN03 U629 ( .A0(n504), .A1(n505), .A2(n506), .Z(n503));
Q_XNR2 U630 ( .A0(drng_256_last[127]), .A1(drng_256_out[127]), .Z(n504));
Q_XNR2 U631 ( .A0(drng_256_last[126]), .A1(drng_256_out[126]), .Z(n505));
Q_XNR2 U632 ( .A0(drng_256_last[125]), .A1(drng_256_out[125]), .Z(n506));
Q_XNR2 U633 ( .A0(drng_256_last[124]), .A1(drng_256_out[124]), .Z(n507));
Q_XNR2 U634 ( .A0(drng_256_last[123]), .A1(drng_256_out[123]), .Z(n508));
Q_XNR2 U635 ( .A0(drng_256_last[122]), .A1(drng_256_out[122]), .Z(n509));
Q_XNR2 U636 ( .A0(drng_256_last[121]), .A1(drng_256_out[121]), .Z(n510));
Q_XNR2 U637 ( .A0(drng_256_last[120]), .A1(drng_256_out[120]), .Z(n511));
Q_XNR2 U638 ( .A0(drng_256_last[119]), .A1(drng_256_out[119]), .Z(n512));
Q_XNR2 U639 ( .A0(drng_256_last[118]), .A1(drng_256_out[118]), .Z(n513));
Q_XNR2 U640 ( .A0(drng_256_last[117]), .A1(drng_256_out[117]), .Z(n514));
Q_XNR2 U641 ( .A0(drng_256_last[116]), .A1(drng_256_out[116]), .Z(n515));
Q_XNR2 U642 ( .A0(drng_256_last[115]), .A1(drng_256_out[115]), .Z(n516));
Q_XNR2 U643 ( .A0(drng_256_last[114]), .A1(drng_256_out[114]), .Z(n517));
Q_XNR2 U644 ( .A0(drng_256_last[113]), .A1(drng_256_out[113]), .Z(n518));
Q_XNR2 U645 ( .A0(drng_256_last[112]), .A1(drng_256_out[112]), .Z(n519));
Q_XNR2 U646 ( .A0(drng_256_last[111]), .A1(drng_256_out[111]), .Z(n520));
Q_XNR2 U647 ( .A0(drng_256_last[110]), .A1(drng_256_out[110]), .Z(n521));
Q_XNR2 U648 ( .A0(drng_256_last[109]), .A1(drng_256_out[109]), .Z(n522));
Q_XNR2 U649 ( .A0(drng_256_last[108]), .A1(drng_256_out[108]), .Z(n523));
Q_XNR2 U650 ( .A0(drng_256_last[107]), .A1(drng_256_out[107]), .Z(n524));
Q_XNR2 U651 ( .A0(drng_256_last[106]), .A1(drng_256_out[106]), .Z(n525));
Q_XNR2 U652 ( .A0(drng_256_last[105]), .A1(drng_256_out[105]), .Z(n526));
Q_XNR2 U653 ( .A0(drng_256_last[104]), .A1(drng_256_out[104]), .Z(n527));
Q_XNR2 U654 ( .A0(drng_256_last[103]), .A1(drng_256_out[103]), .Z(n528));
Q_XNR2 U655 ( .A0(drng_256_last[102]), .A1(drng_256_out[102]), .Z(n529));
Q_XNR2 U656 ( .A0(drng_256_last[101]), .A1(drng_256_out[101]), .Z(n530));
Q_XNR2 U657 ( .A0(drng_256_last[100]), .A1(drng_256_out[100]), .Z(n531));
Q_XNR2 U658 ( .A0(drng_256_last[99]), .A1(drng_256_out[99]), .Z(n532));
Q_XNR2 U659 ( .A0(drng_256_last[98]), .A1(drng_256_out[98]), .Z(n533));
Q_XNR2 U660 ( .A0(drng_256_last[97]), .A1(drng_256_out[97]), .Z(n534));
Q_XNR2 U661 ( .A0(drng_256_last[96]), .A1(drng_256_out[96]), .Z(n535));
Q_XNR2 U662 ( .A0(drng_256_last[95]), .A1(drng_256_out[95]), .Z(n536));
Q_XNR2 U663 ( .A0(drng_256_last[94]), .A1(drng_256_out[94]), .Z(n537));
Q_XNR2 U664 ( .A0(drng_256_last[93]), .A1(drng_256_out[93]), .Z(n538));
Q_XNR2 U665 ( .A0(drng_256_last[92]), .A1(drng_256_out[92]), .Z(n539));
Q_XNR2 U666 ( .A0(drng_256_last[91]), .A1(drng_256_out[91]), .Z(n540));
Q_XNR2 U667 ( .A0(drng_256_last[90]), .A1(drng_256_out[90]), .Z(n541));
Q_XNR2 U668 ( .A0(drng_256_last[89]), .A1(drng_256_out[89]), .Z(n542));
Q_XNR2 U669 ( .A0(drng_256_last[88]), .A1(drng_256_out[88]), .Z(n543));
Q_XNR2 U670 ( .A0(drng_256_last[87]), .A1(drng_256_out[87]), .Z(n544));
Q_XNR2 U671 ( .A0(drng_256_last[86]), .A1(drng_256_out[86]), .Z(n545));
Q_XNR2 U672 ( .A0(drng_256_last[85]), .A1(drng_256_out[85]), .Z(n546));
Q_XNR2 U673 ( .A0(drng_256_last[84]), .A1(drng_256_out[84]), .Z(n547));
Q_XNR2 U674 ( .A0(drng_256_last[83]), .A1(drng_256_out[83]), .Z(n548));
Q_XNR2 U675 ( .A0(drng_256_last[82]), .A1(drng_256_out[82]), .Z(n549));
Q_XNR2 U676 ( .A0(drng_256_last[81]), .A1(drng_256_out[81]), .Z(n550));
Q_XNR2 U677 ( .A0(drng_256_last[80]), .A1(drng_256_out[80]), .Z(n551));
Q_XNR2 U678 ( .A0(drng_256_last[79]), .A1(drng_256_out[79]), .Z(n552));
Q_XNR2 U679 ( .A0(drng_256_last[78]), .A1(drng_256_out[78]), .Z(n553));
Q_XNR2 U680 ( .A0(drng_256_last[77]), .A1(drng_256_out[77]), .Z(n554));
Q_XNR2 U681 ( .A0(drng_256_last[76]), .A1(drng_256_out[76]), .Z(n555));
Q_XNR2 U682 ( .A0(drng_256_last[75]), .A1(drng_256_out[75]), .Z(n556));
Q_XNR2 U683 ( .A0(drng_256_last[74]), .A1(drng_256_out[74]), .Z(n557));
Q_XNR2 U684 ( .A0(drng_256_last[73]), .A1(drng_256_out[73]), .Z(n558));
Q_XNR2 U685 ( .A0(drng_256_last[72]), .A1(drng_256_out[72]), .Z(n559));
Q_XNR2 U686 ( .A0(drng_256_last[71]), .A1(drng_256_out[71]), .Z(n560));
Q_XNR2 U687 ( .A0(drng_256_last[70]), .A1(drng_256_out[70]), .Z(n561));
Q_XNR2 U688 ( .A0(drng_256_last[69]), .A1(drng_256_out[69]), .Z(n562));
Q_XNR2 U689 ( .A0(drng_256_last[68]), .A1(drng_256_out[68]), .Z(n563));
Q_XNR2 U690 ( .A0(drng_256_last[67]), .A1(drng_256_out[67]), .Z(n564));
Q_XNR2 U691 ( .A0(drng_256_last[66]), .A1(drng_256_out[66]), .Z(n565));
Q_XNR2 U692 ( .A0(drng_256_last[65]), .A1(drng_256_out[65]), .Z(n566));
Q_XNR2 U693 ( .A0(drng_256_last[64]), .A1(drng_256_out[64]), .Z(n567));
Q_XNR2 U694 ( .A0(drng_256_last[63]), .A1(drng_256_out[63]), .Z(n568));
Q_XNR2 U695 ( .A0(drng_256_last[62]), .A1(drng_256_out[62]), .Z(n569));
Q_XNR2 U696 ( .A0(drng_256_last[61]), .A1(drng_256_out[61]), .Z(n570));
Q_XNR2 U697 ( .A0(drng_256_last[60]), .A1(drng_256_out[60]), .Z(n571));
Q_XNR2 U698 ( .A0(drng_256_last[59]), .A1(drng_256_out[59]), .Z(n572));
Q_XNR2 U699 ( .A0(drng_256_last[58]), .A1(drng_256_out[58]), .Z(n573));
Q_XNR2 U700 ( .A0(drng_256_last[57]), .A1(drng_256_out[57]), .Z(n574));
Q_XNR2 U701 ( .A0(drng_256_last[56]), .A1(drng_256_out[56]), .Z(n575));
Q_XNR2 U702 ( .A0(drng_256_last[55]), .A1(drng_256_out[55]), .Z(n576));
Q_XNR2 U703 ( .A0(drng_256_last[54]), .A1(drng_256_out[54]), .Z(n577));
Q_XNR2 U704 ( .A0(drng_256_last[53]), .A1(drng_256_out[53]), .Z(n578));
Q_XNR2 U705 ( .A0(drng_256_last[52]), .A1(drng_256_out[52]), .Z(n579));
Q_XNR2 U706 ( .A0(drng_256_last[51]), .A1(drng_256_out[51]), .Z(n580));
Q_XNR2 U707 ( .A0(drng_256_last[50]), .A1(drng_256_out[50]), .Z(n581));
Q_XNR2 U708 ( .A0(drng_256_last[49]), .A1(drng_256_out[49]), .Z(n582));
Q_XNR2 U709 ( .A0(drng_256_last[48]), .A1(drng_256_out[48]), .Z(n583));
Q_XNR2 U710 ( .A0(drng_256_last[47]), .A1(drng_256_out[47]), .Z(n584));
Q_XNR2 U711 ( .A0(drng_256_last[46]), .A1(drng_256_out[46]), .Z(n585));
Q_XNR2 U712 ( .A0(drng_256_last[45]), .A1(drng_256_out[45]), .Z(n586));
Q_XNR2 U713 ( .A0(drng_256_last[44]), .A1(drng_256_out[44]), .Z(n587));
Q_XNR2 U714 ( .A0(drng_256_last[43]), .A1(drng_256_out[43]), .Z(n588));
Q_XNR2 U715 ( .A0(drng_256_last[42]), .A1(drng_256_out[42]), .Z(n589));
Q_XNR2 U716 ( .A0(drng_256_last[41]), .A1(drng_256_out[41]), .Z(n590));
Q_XNR2 U717 ( .A0(drng_256_last[40]), .A1(drng_256_out[40]), .Z(n591));
Q_XNR2 U718 ( .A0(drng_256_last[39]), .A1(drng_256_out[39]), .Z(n592));
Q_XNR2 U719 ( .A0(drng_256_last[38]), .A1(drng_256_out[38]), .Z(n593));
Q_XNR2 U720 ( .A0(drng_256_last[37]), .A1(drng_256_out[37]), .Z(n594));
Q_XNR2 U721 ( .A0(drng_256_last[36]), .A1(drng_256_out[36]), .Z(n595));
Q_XNR2 U722 ( .A0(drng_256_last[35]), .A1(drng_256_out[35]), .Z(n596));
Q_XNR2 U723 ( .A0(drng_256_last[34]), .A1(drng_256_out[34]), .Z(n597));
Q_XNR2 U724 ( .A0(drng_256_last[33]), .A1(drng_256_out[33]), .Z(n598));
Q_XNR2 U725 ( .A0(drng_256_last[32]), .A1(drng_256_out[32]), .Z(n599));
Q_XNR2 U726 ( .A0(drng_256_last[31]), .A1(drng_256_out[31]), .Z(n600));
Q_XNR2 U727 ( .A0(drng_256_last[30]), .A1(drng_256_out[30]), .Z(n601));
Q_XNR2 U728 ( .A0(drng_256_last[29]), .A1(drng_256_out[29]), .Z(n602));
Q_XNR2 U729 ( .A0(drng_256_last[28]), .A1(drng_256_out[28]), .Z(n603));
Q_XNR2 U730 ( .A0(drng_256_last[27]), .A1(drng_256_out[27]), .Z(n604));
Q_XNR2 U731 ( .A0(drng_256_last[26]), .A1(drng_256_out[26]), .Z(n605));
Q_XNR2 U732 ( .A0(drng_256_last[25]), .A1(drng_256_out[25]), .Z(n606));
Q_XNR2 U733 ( .A0(drng_256_last[24]), .A1(drng_256_out[24]), .Z(n607));
Q_XNR2 U734 ( .A0(drng_256_last[23]), .A1(drng_256_out[23]), .Z(n608));
Q_XNR2 U735 ( .A0(drng_256_last[22]), .A1(drng_256_out[22]), .Z(n609));
Q_XNR2 U736 ( .A0(drng_256_last[21]), .A1(drng_256_out[21]), .Z(n610));
Q_XNR2 U737 ( .A0(drng_256_last[20]), .A1(drng_256_out[20]), .Z(n611));
Q_XNR2 U738 ( .A0(drng_256_last[19]), .A1(drng_256_out[19]), .Z(n612));
Q_XNR2 U739 ( .A0(drng_256_last[18]), .A1(drng_256_out[18]), .Z(n613));
Q_XNR2 U740 ( .A0(drng_256_last[17]), .A1(drng_256_out[17]), .Z(n614));
Q_XNR2 U741 ( .A0(drng_256_last[16]), .A1(drng_256_out[16]), .Z(n615));
Q_XNR2 U742 ( .A0(drng_256_last[15]), .A1(drng_256_out[15]), .Z(n616));
Q_XNR2 U743 ( .A0(drng_256_last[14]), .A1(drng_256_out[14]), .Z(n617));
Q_XNR2 U744 ( .A0(drng_256_last[13]), .A1(drng_256_out[13]), .Z(n618));
Q_XNR2 U745 ( .A0(drng_256_last[12]), .A1(drng_256_out[12]), .Z(n619));
Q_XNR2 U746 ( .A0(drng_256_last[11]), .A1(drng_256_out[11]), .Z(n620));
Q_XNR2 U747 ( .A0(drng_256_last[10]), .A1(drng_256_out[10]), .Z(n621));
Q_XNR2 U748 ( .A0(drng_256_last[9]), .A1(drng_256_out[9]), .Z(n622));
Q_XNR2 U749 ( .A0(drng_256_last[8]), .A1(drng_256_out[8]), .Z(n623));
Q_XNR2 U750 ( .A0(drng_256_last[7]), .A1(drng_256_out[7]), .Z(n624));
Q_XNR2 U751 ( .A0(drng_256_last[6]), .A1(drng_256_out[6]), .Z(n625));
Q_XNR2 U752 ( .A0(drng_256_last[5]), .A1(drng_256_out[5]), .Z(n626));
Q_XNR2 U753 ( .A0(drng_256_last[4]), .A1(drng_256_out[4]), .Z(n627));
Q_XNR2 U754 ( .A0(drng_256_last[3]), .A1(drng_256_out[3]), .Z(n628));
Q_XNR2 U755 ( .A0(drng_256_last[2]), .A1(drng_256_out[2]), .Z(n629));
Q_XNR2 U756 ( .A0(drng_256_last[1]), .A1(drng_256_out[1]), .Z(n630));
Q_XNR2 U757 ( .A0(drng_256_last[0]), .A1(drng_256_out[0]), .Z(n631));
ixc_assign_384 _zz_strnp_0 ( { \seed[0][383] , \seed[0][382] , \seed[0][381] , 
	\seed[0][380] , \seed[0][379] , \seed[0][378] , \seed[0][377] , 
	\seed[0][376] , \seed[0][375] , \seed[0][374] , \seed[0][373] , 
	\seed[0][372] , \seed[0][371] , \seed[0][370] , \seed[0][369] , 
	\seed[0][368] , \seed[0][367] , \seed[0][366] , \seed[0][365] , 
	\seed[0][364] , \seed[0][363] , \seed[0][362] , \seed[0][361] , 
	\seed[0][360] , \seed[0][359] , \seed[0][358] , \seed[0][357] , 
	\seed[0][356] , \seed[0][355] , \seed[0][354] , \seed[0][353] , 
	\seed[0][352] , \seed[0][351] , \seed[0][350] , \seed[0][349] , 
	\seed[0][348] , \seed[0][347] , \seed[0][346] , \seed[0][345] , 
	\seed[0][344] , \seed[0][343] , \seed[0][342] , \seed[0][341] , 
	\seed[0][340] , \seed[0][339] , \seed[0][338] , \seed[0][337] , 
	\seed[0][336] , \seed[0][335] , \seed[0][334] , \seed[0][333] , 
	\seed[0][332] , \seed[0][331] , \seed[0][330] , \seed[0][329] , 
	\seed[0][328] , \seed[0][327] , \seed[0][326] , \seed[0][325] , 
	\seed[0][324] , \seed[0][323] , \seed[0][322] , \seed[0][321] , 
	\seed[0][320] , \seed[0][319] , \seed[0][318] , \seed[0][317] , 
	\seed[0][316] , \seed[0][315] , \seed[0][314] , \seed[0][313] , 
	\seed[0][312] , \seed[0][311] , \seed[0][310] , \seed[0][309] , 
	\seed[0][308] , \seed[0][307] , \seed[0][306] , \seed[0][305] , 
	\seed[0][304] , \seed[0][303] , \seed[0][302] , \seed[0][301] , 
	\seed[0][300] , \seed[0][299] , \seed[0][298] , \seed[0][297] , 
	\seed[0][296] , \seed[0][295] , \seed[0][294] , \seed[0][293] , 
	\seed[0][292] , \seed[0][291] , \seed[0][290] , \seed[0][289] , 
	\seed[0][288] , \seed[0][287] , \seed[0][286] , \seed[0][285] , 
	\seed[0][284] , \seed[0][283] , \seed[0][282] , \seed[0][281] , 
	\seed[0][280] , \seed[0][279] , \seed[0][278] , \seed[0][277] , 
	\seed[0][276] , \seed[0][275] , \seed[0][274] , \seed[0][273] , 
	\seed[0][272] , \seed[0][271] , \seed[0][270] , \seed[0][269] , 
	\seed[0][268] , \seed[0][267] , \seed[0][266] , \seed[0][265] , 
	\seed[0][264] , \seed[0][263] , \seed[0][262] , \seed[0][261] , 
	\seed[0][260] , \seed[0][259] , \seed[0][258] , \seed[0][257] , 
	\seed[0][256] , \seed[0][255] , \seed[0][254] , \seed[0][253] , 
	\seed[0][252] , \seed[0][251] , \seed[0][250] , \seed[0][249] , 
	\seed[0][248] , \seed[0][247] , \seed[0][246] , \seed[0][245] , 
	\seed[0][244] , \seed[0][243] , \seed[0][242] , \seed[0][241] , 
	\seed[0][240] , \seed[0][239] , \seed[0][238] , \seed[0][237] , 
	\seed[0][236] , \seed[0][235] , \seed[0][234] , \seed[0][233] , 
	\seed[0][232] , \seed[0][231] , \seed[0][230] , \seed[0][229] , 
	\seed[0][228] , \seed[0][227] , \seed[0][226] , \seed[0][225] , 
	\seed[0][224] , \seed[0][223] , \seed[0][222] , \seed[0][221] , 
	\seed[0][220] , \seed[0][219] , \seed[0][218] , \seed[0][217] , 
	\seed[0][216] , \seed[0][215] , \seed[0][214] , \seed[0][213] , 
	\seed[0][212] , \seed[0][211] , \seed[0][210] , \seed[0][209] , 
	\seed[0][208] , \seed[0][207] , \seed[0][206] , \seed[0][205] , 
	\seed[0][204] , \seed[0][203] , \seed[0][202] , \seed[0][201] , 
	\seed[0][200] , \seed[0][199] , \seed[0][198] , \seed[0][197] , 
	\seed[0][196] , \seed[0][195] , \seed[0][194] , \seed[0][193] , 
	\seed[0][192] , \seed[0][191] , \seed[0][190] , \seed[0][189] , 
	\seed[0][188] , \seed[0][187] , \seed[0][186] , \seed[0][185] , 
	\seed[0][184] , \seed[0][183] , \seed[0][182] , \seed[0][181] , 
	\seed[0][180] , \seed[0][179] , \seed[0][178] , \seed[0][177] , 
	\seed[0][176] , \seed[0][175] , \seed[0][174] , \seed[0][173] , 
	\seed[0][172] , \seed[0][171] , \seed[0][170] , \seed[0][169] , 
	\seed[0][168] , \seed[0][167] , \seed[0][166] , \seed[0][165] , 
	\seed[0][164] , \seed[0][163] , \seed[0][162] , \seed[0][161] , 
	\seed[0][160] , \seed[0][159] , \seed[0][158] , \seed[0][157] , 
	\seed[0][156] , \seed[0][155] , \seed[0][154] , \seed[0][153] , 
	\seed[0][152] , \seed[0][151] , \seed[0][150] , \seed[0][149] , 
	\seed[0][148] , \seed[0][147] , \seed[0][146] , \seed[0][145] , 
	\seed[0][144] , \seed[0][143] , \seed[0][142] , \seed[0][141] , 
	\seed[0][140] , \seed[0][139] , \seed[0][138] , \seed[0][137] , 
	\seed[0][136] , \seed[0][135] , \seed[0][134] , \seed[0][133] , 
	\seed[0][132] , \seed[0][131] , \seed[0][130] , \seed[0][129] , 
	\seed[0][128] , \seed[0][127] , \seed[0][126] , \seed[0][125] , 
	\seed[0][124] , \seed[0][123] , \seed[0][122] , \seed[0][121] , 
	\seed[0][120] , \seed[0][119] , \seed[0][118] , \seed[0][117] , 
	\seed[0][116] , \seed[0][115] , \seed[0][114] , \seed[0][113] , 
	\seed[0][112] , \seed[0][111] , \seed[0][110] , \seed[0][109] , 
	\seed[0][108] , \seed[0][107] , \seed[0][106] , \seed[0][105] , 
	\seed[0][104] , \seed[0][103] , \seed[0][102] , \seed[0][101] , 
	\seed[0][100] , \seed[0][99] , \seed[0][98] , \seed[0][97] , 
	\seed[0][96] , \seed[0][95] , \seed[0][94] , \seed[0][93] , 
	\seed[0][92] , \seed[0][91] , \seed[0][90] , \seed[0][89] , 
	\seed[0][88] , \seed[0][87] , \seed[0][86] , \seed[0][85] , 
	\seed[0][84] , \seed[0][83] , \seed[0][82] , \seed[0][81] , 
	\seed[0][80] , \seed[0][79] , \seed[0][78] , \seed[0][77] , 
	\seed[0][76] , \seed[0][75] , \seed[0][74] , \seed[0][73] , 
	\seed[0][72] , \seed[0][71] , \seed[0][70] , \seed[0][69] , 
	\seed[0][68] , \seed[0][67] , \seed[0][66] , \seed[0][65] , 
	\seed[0][64] , \seed[0][63] , \seed[0][62] , \seed[0][61] , 
	\seed[0][60] , \seed[0][59] , \seed[0][58] , \seed[0][57] , 
	\seed[0][56] , \seed[0][55] , \seed[0][54] , \seed[0][53] , 
	\seed[0][52] , \seed[0][51] , \seed[0][50] , \seed[0][49] , 
	\seed[0][48] , \seed[0][47] , \seed[0][46] , \seed[0][45] , 
	\seed[0][44] , \seed[0][43] , \seed[0][42] , \seed[0][41] , 
	\seed[0][40] , \seed[0][39] , \seed[0][38] , \seed[0][37] , 
	\seed[0][36] , \seed[0][35] , \seed[0][34] , \seed[0][33] , 
	\seed[0][32] , \seed[0][31] , \seed[0][30] , \seed[0][29] , 
	\seed[0][28] , \seed[0][27] , \seed[0][26] , \seed[0][25] , 
	\seed[0][24] , \seed[0][23] , \seed[0][22] , \seed[0][21] , 
	\seed[0][20] , \seed[0][19] , \seed[0][18] , \seed[0][17] , 
	\seed[0][16] , \seed[0][15] , \seed[0][14] , \seed[0][13] , 
	\seed[0][12] , \seed[0][11] , \seed[0][10] , \seed[0][9] , 
	\seed[0][8] , \seed[0][7] , \seed[0][6] , \seed[0][5] , \seed[0][4] , 
	\seed[0][3] , \seed[0][2] , \seed[0][1] , \seed[0][0] }, { 
	seed0_internal_state_key[255], seed0_internal_state_key[254], 
	seed0_internal_state_key[253], seed0_internal_state_key[252], 
	seed0_internal_state_key[251], seed0_internal_state_key[250], 
	seed0_internal_state_key[249], seed0_internal_state_key[248], 
	seed0_internal_state_key[247], seed0_internal_state_key[246], 
	seed0_internal_state_key[245], seed0_internal_state_key[244], 
	seed0_internal_state_key[243], seed0_internal_state_key[242], 
	seed0_internal_state_key[241], seed0_internal_state_key[240], 
	seed0_internal_state_key[239], seed0_internal_state_key[238], 
	seed0_internal_state_key[237], seed0_internal_state_key[236], 
	seed0_internal_state_key[235], seed0_internal_state_key[234], 
	seed0_internal_state_key[233], seed0_internal_state_key[232], 
	seed0_internal_state_key[231], seed0_internal_state_key[230], 
	seed0_internal_state_key[229], seed0_internal_state_key[228], 
	seed0_internal_state_key[227], seed0_internal_state_key[226], 
	seed0_internal_state_key[225], seed0_internal_state_key[224], 
	seed0_internal_state_key[223], seed0_internal_state_key[222], 
	seed0_internal_state_key[221], seed0_internal_state_key[220], 
	seed0_internal_state_key[219], seed0_internal_state_key[218], 
	seed0_internal_state_key[217], seed0_internal_state_key[216], 
	seed0_internal_state_key[215], seed0_internal_state_key[214], 
	seed0_internal_state_key[213], seed0_internal_state_key[212], 
	seed0_internal_state_key[211], seed0_internal_state_key[210], 
	seed0_internal_state_key[209], seed0_internal_state_key[208], 
	seed0_internal_state_key[207], seed0_internal_state_key[206], 
	seed0_internal_state_key[205], seed0_internal_state_key[204], 
	seed0_internal_state_key[203], seed0_internal_state_key[202], 
	seed0_internal_state_key[201], seed0_internal_state_key[200], 
	seed0_internal_state_key[199], seed0_internal_state_key[198], 
	seed0_internal_state_key[197], seed0_internal_state_key[196], 
	seed0_internal_state_key[195], seed0_internal_state_key[194], 
	seed0_internal_state_key[193], seed0_internal_state_key[192], 
	seed0_internal_state_key[191], seed0_internal_state_key[190], 
	seed0_internal_state_key[189], seed0_internal_state_key[188], 
	seed0_internal_state_key[187], seed0_internal_state_key[186], 
	seed0_internal_state_key[185], seed0_internal_state_key[184], 
	seed0_internal_state_key[183], seed0_internal_state_key[182], 
	seed0_internal_state_key[181], seed0_internal_state_key[180], 
	seed0_internal_state_key[179], seed0_internal_state_key[178], 
	seed0_internal_state_key[177], seed0_internal_state_key[176], 
	seed0_internal_state_key[175], seed0_internal_state_key[174], 
	seed0_internal_state_key[173], seed0_internal_state_key[172], 
	seed0_internal_state_key[171], seed0_internal_state_key[170], 
	seed0_internal_state_key[169], seed0_internal_state_key[168], 
	seed0_internal_state_key[167], seed0_internal_state_key[166], 
	seed0_internal_state_key[165], seed0_internal_state_key[164], 
	seed0_internal_state_key[163], seed0_internal_state_key[162], 
	seed0_internal_state_key[161], seed0_internal_state_key[160], 
	seed0_internal_state_key[159], seed0_internal_state_key[158], 
	seed0_internal_state_key[157], seed0_internal_state_key[156], 
	seed0_internal_state_key[155], seed0_internal_state_key[154], 
	seed0_internal_state_key[153], seed0_internal_state_key[152], 
	seed0_internal_state_key[151], seed0_internal_state_key[150], 
	seed0_internal_state_key[149], seed0_internal_state_key[148], 
	seed0_internal_state_key[147], seed0_internal_state_key[146], 
	seed0_internal_state_key[145], seed0_internal_state_key[144], 
	seed0_internal_state_key[143], seed0_internal_state_key[142], 
	seed0_internal_state_key[141], seed0_internal_state_key[140], 
	seed0_internal_state_key[139], seed0_internal_state_key[138], 
	seed0_internal_state_key[137], seed0_internal_state_key[136], 
	seed0_internal_state_key[135], seed0_internal_state_key[134], 
	seed0_internal_state_key[133], seed0_internal_state_key[132], 
	seed0_internal_state_key[131], seed0_internal_state_key[130], 
	seed0_internal_state_key[129], seed0_internal_state_key[128], 
	seed0_internal_state_key[127], seed0_internal_state_key[126], 
	seed0_internal_state_key[125], seed0_internal_state_key[124], 
	seed0_internal_state_key[123], seed0_internal_state_key[122], 
	seed0_internal_state_key[121], seed0_internal_state_key[120], 
	seed0_internal_state_key[119], seed0_internal_state_key[118], 
	seed0_internal_state_key[117], seed0_internal_state_key[116], 
	seed0_internal_state_key[115], seed0_internal_state_key[114], 
	seed0_internal_state_key[113], seed0_internal_state_key[112], 
	seed0_internal_state_key[111], seed0_internal_state_key[110], 
	seed0_internal_state_key[109], seed0_internal_state_key[108], 
	seed0_internal_state_key[107], seed0_internal_state_key[106], 
	seed0_internal_state_key[105], seed0_internal_state_key[104], 
	seed0_internal_state_key[103], seed0_internal_state_key[102], 
	seed0_internal_state_key[101], seed0_internal_state_key[100], 
	seed0_internal_state_key[99], seed0_internal_state_key[98], 
	seed0_internal_state_key[97], seed0_internal_state_key[96], 
	seed0_internal_state_key[95], seed0_internal_state_key[94], 
	seed0_internal_state_key[93], seed0_internal_state_key[92], 
	seed0_internal_state_key[91], seed0_internal_state_key[90], 
	seed0_internal_state_key[89], seed0_internal_state_key[88], 
	seed0_internal_state_key[87], seed0_internal_state_key[86], 
	seed0_internal_state_key[85], seed0_internal_state_key[84], 
	seed0_internal_state_key[83], seed0_internal_state_key[82], 
	seed0_internal_state_key[81], seed0_internal_state_key[80], 
	seed0_internal_state_key[79], seed0_internal_state_key[78], 
	seed0_internal_state_key[77], seed0_internal_state_key[76], 
	seed0_internal_state_key[75], seed0_internal_state_key[74], 
	seed0_internal_state_key[73], seed0_internal_state_key[72], 
	seed0_internal_state_key[71], seed0_internal_state_key[70], 
	seed0_internal_state_key[69], seed0_internal_state_key[68], 
	seed0_internal_state_key[67], seed0_internal_state_key[66], 
	seed0_internal_state_key[65], seed0_internal_state_key[64], 
	seed0_internal_state_key[63], seed0_internal_state_key[62], 
	seed0_internal_state_key[61], seed0_internal_state_key[60], 
	seed0_internal_state_key[59], seed0_internal_state_key[58], 
	seed0_internal_state_key[57], seed0_internal_state_key[56], 
	seed0_internal_state_key[55], seed0_internal_state_key[54], 
	seed0_internal_state_key[53], seed0_internal_state_key[52], 
	seed0_internal_state_key[51], seed0_internal_state_key[50], 
	seed0_internal_state_key[49], seed0_internal_state_key[48], 
	seed0_internal_state_key[47], seed0_internal_state_key[46], 
	seed0_internal_state_key[45], seed0_internal_state_key[44], 
	seed0_internal_state_key[43], seed0_internal_state_key[42], 
	seed0_internal_state_key[41], seed0_internal_state_key[40], 
	seed0_internal_state_key[39], seed0_internal_state_key[38], 
	seed0_internal_state_key[37], seed0_internal_state_key[36], 
	seed0_internal_state_key[35], seed0_internal_state_key[34], 
	seed0_internal_state_key[33], seed0_internal_state_key[32], 
	seed0_internal_state_key[31], seed0_internal_state_key[30], 
	seed0_internal_state_key[29], seed0_internal_state_key[28], 
	seed0_internal_state_key[27], seed0_internal_state_key[26], 
	seed0_internal_state_key[25], seed0_internal_state_key[24], 
	seed0_internal_state_key[23], seed0_internal_state_key[22], 
	seed0_internal_state_key[21], seed0_internal_state_key[20], 
	seed0_internal_state_key[19], seed0_internal_state_key[18], 
	seed0_internal_state_key[17], seed0_internal_state_key[16], 
	seed0_internal_state_key[15], seed0_internal_state_key[14], 
	seed0_internal_state_key[13], seed0_internal_state_key[12], 
	seed0_internal_state_key[11], seed0_internal_state_key[10], 
	seed0_internal_state_key[9], seed0_internal_state_key[8], 
	seed0_internal_state_key[7], seed0_internal_state_key[6], 
	seed0_internal_state_key[5], seed0_internal_state_key[4], 
	seed0_internal_state_key[3], seed0_internal_state_key[2], 
	seed0_internal_state_key[1], seed0_internal_state_key[0], 
	seed0_internal_state_value[127], seed0_internal_state_value[126], 
	seed0_internal_state_value[125], seed0_internal_state_value[124], 
	seed0_internal_state_value[123], seed0_internal_state_value[122], 
	seed0_internal_state_value[121], seed0_internal_state_value[120], 
	seed0_internal_state_value[119], seed0_internal_state_value[118], 
	seed0_internal_state_value[117], seed0_internal_state_value[116], 
	seed0_internal_state_value[115], seed0_internal_state_value[114], 
	seed0_internal_state_value[113], seed0_internal_state_value[112], 
	seed0_internal_state_value[111], seed0_internal_state_value[110], 
	seed0_internal_state_value[109], seed0_internal_state_value[108], 
	seed0_internal_state_value[107], seed0_internal_state_value[106], 
	seed0_internal_state_value[105], seed0_internal_state_value[104], 
	seed0_internal_state_value[103], seed0_internal_state_value[102], 
	seed0_internal_state_value[101], seed0_internal_state_value[100], 
	seed0_internal_state_value[99], seed0_internal_state_value[98], 
	seed0_internal_state_value[97], seed0_internal_state_value[96], 
	seed0_internal_state_value[95], seed0_internal_state_value[94], 
	seed0_internal_state_value[93], seed0_internal_state_value[92], 
	seed0_internal_state_value[91], seed0_internal_state_value[90], 
	seed0_internal_state_value[89], seed0_internal_state_value[88], 
	seed0_internal_state_value[87], seed0_internal_state_value[86], 
	seed0_internal_state_value[85], seed0_internal_state_value[84], 
	seed0_internal_state_value[83], seed0_internal_state_value[82], 
	seed0_internal_state_value[81], seed0_internal_state_value[80], 
	seed0_internal_state_value[79], seed0_internal_state_value[78], 
	seed0_internal_state_value[77], seed0_internal_state_value[76], 
	seed0_internal_state_value[75], seed0_internal_state_value[74], 
	seed0_internal_state_value[73], seed0_internal_state_value[72], 
	seed0_internal_state_value[71], seed0_internal_state_value[70], 
	seed0_internal_state_value[69], seed0_internal_state_value[68], 
	seed0_internal_state_value[67], seed0_internal_state_value[66], 
	seed0_internal_state_value[65], seed0_internal_state_value[64], 
	seed0_internal_state_value[63], seed0_internal_state_value[62], 
	seed0_internal_state_value[61], seed0_internal_state_value[60], 
	seed0_internal_state_value[59], seed0_internal_state_value[58], 
	seed0_internal_state_value[57], seed0_internal_state_value[56], 
	seed0_internal_state_value[55], seed0_internal_state_value[54], 
	seed0_internal_state_value[53], seed0_internal_state_value[52], 
	seed0_internal_state_value[51], seed0_internal_state_value[50], 
	seed0_internal_state_value[49], seed0_internal_state_value[48], 
	seed0_internal_state_value[47], seed0_internal_state_value[46], 
	seed0_internal_state_value[45], seed0_internal_state_value[44], 
	seed0_internal_state_value[43], seed0_internal_state_value[42], 
	seed0_internal_state_value[41], seed0_internal_state_value[40], 
	seed0_internal_state_value[39], seed0_internal_state_value[38], 
	seed0_internal_state_value[37], seed0_internal_state_value[36], 
	seed0_internal_state_value[35], seed0_internal_state_value[34], 
	seed0_internal_state_value[33], seed0_internal_state_value[32], 
	seed0_internal_state_value[31], seed0_internal_state_value[30], 
	seed0_internal_state_value[29], seed0_internal_state_value[28], 
	seed0_internal_state_value[27], seed0_internal_state_value[26], 
	seed0_internal_state_value[25], seed0_internal_state_value[24], 
	seed0_internal_state_value[23], seed0_internal_state_value[22], 
	seed0_internal_state_value[21], seed0_internal_state_value[20], 
	seed0_internal_state_value[19], seed0_internal_state_value[18], 
	seed0_internal_state_value[17], seed0_internal_state_value[16], 
	seed0_internal_state_value[15], seed0_internal_state_value[14], 
	seed0_internal_state_value[13], seed0_internal_state_value[12], 
	seed0_internal_state_value[11], seed0_internal_state_value[10], 
	seed0_internal_state_value[9], seed0_internal_state_value[8], 
	seed0_internal_state_value[7], seed0_internal_state_value[6], 
	seed0_internal_state_value[5], seed0_internal_state_value[4], 
	seed0_internal_state_value[3], seed0_internal_state_value[2], 
	seed0_internal_state_value[1], seed0_internal_state_value[0]});
ixc_assign_384 _zz_strnp_1 ( { \seed[1][383] , \seed[1][382] , \seed[1][381] , 
	\seed[1][380] , \seed[1][379] , \seed[1][378] , \seed[1][377] , 
	\seed[1][376] , \seed[1][375] , \seed[1][374] , \seed[1][373] , 
	\seed[1][372] , \seed[1][371] , \seed[1][370] , \seed[1][369] , 
	\seed[1][368] , \seed[1][367] , \seed[1][366] , \seed[1][365] , 
	\seed[1][364] , \seed[1][363] , \seed[1][362] , \seed[1][361] , 
	\seed[1][360] , \seed[1][359] , \seed[1][358] , \seed[1][357] , 
	\seed[1][356] , \seed[1][355] , \seed[1][354] , \seed[1][353] , 
	\seed[1][352] , \seed[1][351] , \seed[1][350] , \seed[1][349] , 
	\seed[1][348] , \seed[1][347] , \seed[1][346] , \seed[1][345] , 
	\seed[1][344] , \seed[1][343] , \seed[1][342] , \seed[1][341] , 
	\seed[1][340] , \seed[1][339] , \seed[1][338] , \seed[1][337] , 
	\seed[1][336] , \seed[1][335] , \seed[1][334] , \seed[1][333] , 
	\seed[1][332] , \seed[1][331] , \seed[1][330] , \seed[1][329] , 
	\seed[1][328] , \seed[1][327] , \seed[1][326] , \seed[1][325] , 
	\seed[1][324] , \seed[1][323] , \seed[1][322] , \seed[1][321] , 
	\seed[1][320] , \seed[1][319] , \seed[1][318] , \seed[1][317] , 
	\seed[1][316] , \seed[1][315] , \seed[1][314] , \seed[1][313] , 
	\seed[1][312] , \seed[1][311] , \seed[1][310] , \seed[1][309] , 
	\seed[1][308] , \seed[1][307] , \seed[1][306] , \seed[1][305] , 
	\seed[1][304] , \seed[1][303] , \seed[1][302] , \seed[1][301] , 
	\seed[1][300] , \seed[1][299] , \seed[1][298] , \seed[1][297] , 
	\seed[1][296] , \seed[1][295] , \seed[1][294] , \seed[1][293] , 
	\seed[1][292] , \seed[1][291] , \seed[1][290] , \seed[1][289] , 
	\seed[1][288] , \seed[1][287] , \seed[1][286] , \seed[1][285] , 
	\seed[1][284] , \seed[1][283] , \seed[1][282] , \seed[1][281] , 
	\seed[1][280] , \seed[1][279] , \seed[1][278] , \seed[1][277] , 
	\seed[1][276] , \seed[1][275] , \seed[1][274] , \seed[1][273] , 
	\seed[1][272] , \seed[1][271] , \seed[1][270] , \seed[1][269] , 
	\seed[1][268] , \seed[1][267] , \seed[1][266] , \seed[1][265] , 
	\seed[1][264] , \seed[1][263] , \seed[1][262] , \seed[1][261] , 
	\seed[1][260] , \seed[1][259] , \seed[1][258] , \seed[1][257] , 
	\seed[1][256] , \seed[1][255] , \seed[1][254] , \seed[1][253] , 
	\seed[1][252] , \seed[1][251] , \seed[1][250] , \seed[1][249] , 
	\seed[1][248] , \seed[1][247] , \seed[1][246] , \seed[1][245] , 
	\seed[1][244] , \seed[1][243] , \seed[1][242] , \seed[1][241] , 
	\seed[1][240] , \seed[1][239] , \seed[1][238] , \seed[1][237] , 
	\seed[1][236] , \seed[1][235] , \seed[1][234] , \seed[1][233] , 
	\seed[1][232] , \seed[1][231] , \seed[1][230] , \seed[1][229] , 
	\seed[1][228] , \seed[1][227] , \seed[1][226] , \seed[1][225] , 
	\seed[1][224] , \seed[1][223] , \seed[1][222] , \seed[1][221] , 
	\seed[1][220] , \seed[1][219] , \seed[1][218] , \seed[1][217] , 
	\seed[1][216] , \seed[1][215] , \seed[1][214] , \seed[1][213] , 
	\seed[1][212] , \seed[1][211] , \seed[1][210] , \seed[1][209] , 
	\seed[1][208] , \seed[1][207] , \seed[1][206] , \seed[1][205] , 
	\seed[1][204] , \seed[1][203] , \seed[1][202] , \seed[1][201] , 
	\seed[1][200] , \seed[1][199] , \seed[1][198] , \seed[1][197] , 
	\seed[1][196] , \seed[1][195] , \seed[1][194] , \seed[1][193] , 
	\seed[1][192] , \seed[1][191] , \seed[1][190] , \seed[1][189] , 
	\seed[1][188] , \seed[1][187] , \seed[1][186] , \seed[1][185] , 
	\seed[1][184] , \seed[1][183] , \seed[1][182] , \seed[1][181] , 
	\seed[1][180] , \seed[1][179] , \seed[1][178] , \seed[1][177] , 
	\seed[1][176] , \seed[1][175] , \seed[1][174] , \seed[1][173] , 
	\seed[1][172] , \seed[1][171] , \seed[1][170] , \seed[1][169] , 
	\seed[1][168] , \seed[1][167] , \seed[1][166] , \seed[1][165] , 
	\seed[1][164] , \seed[1][163] , \seed[1][162] , \seed[1][161] , 
	\seed[1][160] , \seed[1][159] , \seed[1][158] , \seed[1][157] , 
	\seed[1][156] , \seed[1][155] , \seed[1][154] , \seed[1][153] , 
	\seed[1][152] , \seed[1][151] , \seed[1][150] , \seed[1][149] , 
	\seed[1][148] , \seed[1][147] , \seed[1][146] , \seed[1][145] , 
	\seed[1][144] , \seed[1][143] , \seed[1][142] , \seed[1][141] , 
	\seed[1][140] , \seed[1][139] , \seed[1][138] , \seed[1][137] , 
	\seed[1][136] , \seed[1][135] , \seed[1][134] , \seed[1][133] , 
	\seed[1][132] , \seed[1][131] , \seed[1][130] , \seed[1][129] , 
	\seed[1][128] , \seed[1][127] , \seed[1][126] , \seed[1][125] , 
	\seed[1][124] , \seed[1][123] , \seed[1][122] , \seed[1][121] , 
	\seed[1][120] , \seed[1][119] , \seed[1][118] , \seed[1][117] , 
	\seed[1][116] , \seed[1][115] , \seed[1][114] , \seed[1][113] , 
	\seed[1][112] , \seed[1][111] , \seed[1][110] , \seed[1][109] , 
	\seed[1][108] , \seed[1][107] , \seed[1][106] , \seed[1][105] , 
	\seed[1][104] , \seed[1][103] , \seed[1][102] , \seed[1][101] , 
	\seed[1][100] , \seed[1][99] , \seed[1][98] , \seed[1][97] , 
	\seed[1][96] , \seed[1][95] , \seed[1][94] , \seed[1][93] , 
	\seed[1][92] , \seed[1][91] , \seed[1][90] , \seed[1][89] , 
	\seed[1][88] , \seed[1][87] , \seed[1][86] , \seed[1][85] , 
	\seed[1][84] , \seed[1][83] , \seed[1][82] , \seed[1][81] , 
	\seed[1][80] , \seed[1][79] , \seed[1][78] , \seed[1][77] , 
	\seed[1][76] , \seed[1][75] , \seed[1][74] , \seed[1][73] , 
	\seed[1][72] , \seed[1][71] , \seed[1][70] , \seed[1][69] , 
	\seed[1][68] , \seed[1][67] , \seed[1][66] , \seed[1][65] , 
	\seed[1][64] , \seed[1][63] , \seed[1][62] , \seed[1][61] , 
	\seed[1][60] , \seed[1][59] , \seed[1][58] , \seed[1][57] , 
	\seed[1][56] , \seed[1][55] , \seed[1][54] , \seed[1][53] , 
	\seed[1][52] , \seed[1][51] , \seed[1][50] , \seed[1][49] , 
	\seed[1][48] , \seed[1][47] , \seed[1][46] , \seed[1][45] , 
	\seed[1][44] , \seed[1][43] , \seed[1][42] , \seed[1][41] , 
	\seed[1][40] , \seed[1][39] , \seed[1][38] , \seed[1][37] , 
	\seed[1][36] , \seed[1][35] , \seed[1][34] , \seed[1][33] , 
	\seed[1][32] , \seed[1][31] , \seed[1][30] , \seed[1][29] , 
	\seed[1][28] , \seed[1][27] , \seed[1][26] , \seed[1][25] , 
	\seed[1][24] , \seed[1][23] , \seed[1][22] , \seed[1][21] , 
	\seed[1][20] , \seed[1][19] , \seed[1][18] , \seed[1][17] , 
	\seed[1][16] , \seed[1][15] , \seed[1][14] , \seed[1][13] , 
	\seed[1][12] , \seed[1][11] , \seed[1][10] , \seed[1][9] , 
	\seed[1][8] , \seed[1][7] , \seed[1][6] , \seed[1][5] , \seed[1][4] , 
	\seed[1][3] , \seed[1][2] , \seed[1][1] , \seed[1][0] }, { 
	seed1_internal_state_key[255], seed1_internal_state_key[254], 
	seed1_internal_state_key[253], seed1_internal_state_key[252], 
	seed1_internal_state_key[251], seed1_internal_state_key[250], 
	seed1_internal_state_key[249], seed1_internal_state_key[248], 
	seed1_internal_state_key[247], seed1_internal_state_key[246], 
	seed1_internal_state_key[245], seed1_internal_state_key[244], 
	seed1_internal_state_key[243], seed1_internal_state_key[242], 
	seed1_internal_state_key[241], seed1_internal_state_key[240], 
	seed1_internal_state_key[239], seed1_internal_state_key[238], 
	seed1_internal_state_key[237], seed1_internal_state_key[236], 
	seed1_internal_state_key[235], seed1_internal_state_key[234], 
	seed1_internal_state_key[233], seed1_internal_state_key[232], 
	seed1_internal_state_key[231], seed1_internal_state_key[230], 
	seed1_internal_state_key[229], seed1_internal_state_key[228], 
	seed1_internal_state_key[227], seed1_internal_state_key[226], 
	seed1_internal_state_key[225], seed1_internal_state_key[224], 
	seed1_internal_state_key[223], seed1_internal_state_key[222], 
	seed1_internal_state_key[221], seed1_internal_state_key[220], 
	seed1_internal_state_key[219], seed1_internal_state_key[218], 
	seed1_internal_state_key[217], seed1_internal_state_key[216], 
	seed1_internal_state_key[215], seed1_internal_state_key[214], 
	seed1_internal_state_key[213], seed1_internal_state_key[212], 
	seed1_internal_state_key[211], seed1_internal_state_key[210], 
	seed1_internal_state_key[209], seed1_internal_state_key[208], 
	seed1_internal_state_key[207], seed1_internal_state_key[206], 
	seed1_internal_state_key[205], seed1_internal_state_key[204], 
	seed1_internal_state_key[203], seed1_internal_state_key[202], 
	seed1_internal_state_key[201], seed1_internal_state_key[200], 
	seed1_internal_state_key[199], seed1_internal_state_key[198], 
	seed1_internal_state_key[197], seed1_internal_state_key[196], 
	seed1_internal_state_key[195], seed1_internal_state_key[194], 
	seed1_internal_state_key[193], seed1_internal_state_key[192], 
	seed1_internal_state_key[191], seed1_internal_state_key[190], 
	seed1_internal_state_key[189], seed1_internal_state_key[188], 
	seed1_internal_state_key[187], seed1_internal_state_key[186], 
	seed1_internal_state_key[185], seed1_internal_state_key[184], 
	seed1_internal_state_key[183], seed1_internal_state_key[182], 
	seed1_internal_state_key[181], seed1_internal_state_key[180], 
	seed1_internal_state_key[179], seed1_internal_state_key[178], 
	seed1_internal_state_key[177], seed1_internal_state_key[176], 
	seed1_internal_state_key[175], seed1_internal_state_key[174], 
	seed1_internal_state_key[173], seed1_internal_state_key[172], 
	seed1_internal_state_key[171], seed1_internal_state_key[170], 
	seed1_internal_state_key[169], seed1_internal_state_key[168], 
	seed1_internal_state_key[167], seed1_internal_state_key[166], 
	seed1_internal_state_key[165], seed1_internal_state_key[164], 
	seed1_internal_state_key[163], seed1_internal_state_key[162], 
	seed1_internal_state_key[161], seed1_internal_state_key[160], 
	seed1_internal_state_key[159], seed1_internal_state_key[158], 
	seed1_internal_state_key[157], seed1_internal_state_key[156], 
	seed1_internal_state_key[155], seed1_internal_state_key[154], 
	seed1_internal_state_key[153], seed1_internal_state_key[152], 
	seed1_internal_state_key[151], seed1_internal_state_key[150], 
	seed1_internal_state_key[149], seed1_internal_state_key[148], 
	seed1_internal_state_key[147], seed1_internal_state_key[146], 
	seed1_internal_state_key[145], seed1_internal_state_key[144], 
	seed1_internal_state_key[143], seed1_internal_state_key[142], 
	seed1_internal_state_key[141], seed1_internal_state_key[140], 
	seed1_internal_state_key[139], seed1_internal_state_key[138], 
	seed1_internal_state_key[137], seed1_internal_state_key[136], 
	seed1_internal_state_key[135], seed1_internal_state_key[134], 
	seed1_internal_state_key[133], seed1_internal_state_key[132], 
	seed1_internal_state_key[131], seed1_internal_state_key[130], 
	seed1_internal_state_key[129], seed1_internal_state_key[128], 
	seed1_internal_state_key[127], seed1_internal_state_key[126], 
	seed1_internal_state_key[125], seed1_internal_state_key[124], 
	seed1_internal_state_key[123], seed1_internal_state_key[122], 
	seed1_internal_state_key[121], seed1_internal_state_key[120], 
	seed1_internal_state_key[119], seed1_internal_state_key[118], 
	seed1_internal_state_key[117], seed1_internal_state_key[116], 
	seed1_internal_state_key[115], seed1_internal_state_key[114], 
	seed1_internal_state_key[113], seed1_internal_state_key[112], 
	seed1_internal_state_key[111], seed1_internal_state_key[110], 
	seed1_internal_state_key[109], seed1_internal_state_key[108], 
	seed1_internal_state_key[107], seed1_internal_state_key[106], 
	seed1_internal_state_key[105], seed1_internal_state_key[104], 
	seed1_internal_state_key[103], seed1_internal_state_key[102], 
	seed1_internal_state_key[101], seed1_internal_state_key[100], 
	seed1_internal_state_key[99], seed1_internal_state_key[98], 
	seed1_internal_state_key[97], seed1_internal_state_key[96], 
	seed1_internal_state_key[95], seed1_internal_state_key[94], 
	seed1_internal_state_key[93], seed1_internal_state_key[92], 
	seed1_internal_state_key[91], seed1_internal_state_key[90], 
	seed1_internal_state_key[89], seed1_internal_state_key[88], 
	seed1_internal_state_key[87], seed1_internal_state_key[86], 
	seed1_internal_state_key[85], seed1_internal_state_key[84], 
	seed1_internal_state_key[83], seed1_internal_state_key[82], 
	seed1_internal_state_key[81], seed1_internal_state_key[80], 
	seed1_internal_state_key[79], seed1_internal_state_key[78], 
	seed1_internal_state_key[77], seed1_internal_state_key[76], 
	seed1_internal_state_key[75], seed1_internal_state_key[74], 
	seed1_internal_state_key[73], seed1_internal_state_key[72], 
	seed1_internal_state_key[71], seed1_internal_state_key[70], 
	seed1_internal_state_key[69], seed1_internal_state_key[68], 
	seed1_internal_state_key[67], seed1_internal_state_key[66], 
	seed1_internal_state_key[65], seed1_internal_state_key[64], 
	seed1_internal_state_key[63], seed1_internal_state_key[62], 
	seed1_internal_state_key[61], seed1_internal_state_key[60], 
	seed1_internal_state_key[59], seed1_internal_state_key[58], 
	seed1_internal_state_key[57], seed1_internal_state_key[56], 
	seed1_internal_state_key[55], seed1_internal_state_key[54], 
	seed1_internal_state_key[53], seed1_internal_state_key[52], 
	seed1_internal_state_key[51], seed1_internal_state_key[50], 
	seed1_internal_state_key[49], seed1_internal_state_key[48], 
	seed1_internal_state_key[47], seed1_internal_state_key[46], 
	seed1_internal_state_key[45], seed1_internal_state_key[44], 
	seed1_internal_state_key[43], seed1_internal_state_key[42], 
	seed1_internal_state_key[41], seed1_internal_state_key[40], 
	seed1_internal_state_key[39], seed1_internal_state_key[38], 
	seed1_internal_state_key[37], seed1_internal_state_key[36], 
	seed1_internal_state_key[35], seed1_internal_state_key[34], 
	seed1_internal_state_key[33], seed1_internal_state_key[32], 
	seed1_internal_state_key[31], seed1_internal_state_key[30], 
	seed1_internal_state_key[29], seed1_internal_state_key[28], 
	seed1_internal_state_key[27], seed1_internal_state_key[26], 
	seed1_internal_state_key[25], seed1_internal_state_key[24], 
	seed1_internal_state_key[23], seed1_internal_state_key[22], 
	seed1_internal_state_key[21], seed1_internal_state_key[20], 
	seed1_internal_state_key[19], seed1_internal_state_key[18], 
	seed1_internal_state_key[17], seed1_internal_state_key[16], 
	seed1_internal_state_key[15], seed1_internal_state_key[14], 
	seed1_internal_state_key[13], seed1_internal_state_key[12], 
	seed1_internal_state_key[11], seed1_internal_state_key[10], 
	seed1_internal_state_key[9], seed1_internal_state_key[8], 
	seed1_internal_state_key[7], seed1_internal_state_key[6], 
	seed1_internal_state_key[5], seed1_internal_state_key[4], 
	seed1_internal_state_key[3], seed1_internal_state_key[2], 
	seed1_internal_state_key[1], seed1_internal_state_key[0], 
	seed1_internal_state_value[127], seed1_internal_state_value[126], 
	seed1_internal_state_value[125], seed1_internal_state_value[124], 
	seed1_internal_state_value[123], seed1_internal_state_value[122], 
	seed1_internal_state_value[121], seed1_internal_state_value[120], 
	seed1_internal_state_value[119], seed1_internal_state_value[118], 
	seed1_internal_state_value[117], seed1_internal_state_value[116], 
	seed1_internal_state_value[115], seed1_internal_state_value[114], 
	seed1_internal_state_value[113], seed1_internal_state_value[112], 
	seed1_internal_state_value[111], seed1_internal_state_value[110], 
	seed1_internal_state_value[109], seed1_internal_state_value[108], 
	seed1_internal_state_value[107], seed1_internal_state_value[106], 
	seed1_internal_state_value[105], seed1_internal_state_value[104], 
	seed1_internal_state_value[103], seed1_internal_state_value[102], 
	seed1_internal_state_value[101], seed1_internal_state_value[100], 
	seed1_internal_state_value[99], seed1_internal_state_value[98], 
	seed1_internal_state_value[97], seed1_internal_state_value[96], 
	seed1_internal_state_value[95], seed1_internal_state_value[94], 
	seed1_internal_state_value[93], seed1_internal_state_value[92], 
	seed1_internal_state_value[91], seed1_internal_state_value[90], 
	seed1_internal_state_value[89], seed1_internal_state_value[88], 
	seed1_internal_state_value[87], seed1_internal_state_value[86], 
	seed1_internal_state_value[85], seed1_internal_state_value[84], 
	seed1_internal_state_value[83], seed1_internal_state_value[82], 
	seed1_internal_state_value[81], seed1_internal_state_value[80], 
	seed1_internal_state_value[79], seed1_internal_state_value[78], 
	seed1_internal_state_value[77], seed1_internal_state_value[76], 
	seed1_internal_state_value[75], seed1_internal_state_value[74], 
	seed1_internal_state_value[73], seed1_internal_state_value[72], 
	seed1_internal_state_value[71], seed1_internal_state_value[70], 
	seed1_internal_state_value[69], seed1_internal_state_value[68], 
	seed1_internal_state_value[67], seed1_internal_state_value[66], 
	seed1_internal_state_value[65], seed1_internal_state_value[64], 
	seed1_internal_state_value[63], seed1_internal_state_value[62], 
	seed1_internal_state_value[61], seed1_internal_state_value[60], 
	seed1_internal_state_value[59], seed1_internal_state_value[58], 
	seed1_internal_state_value[57], seed1_internal_state_value[56], 
	seed1_internal_state_value[55], seed1_internal_state_value[54], 
	seed1_internal_state_value[53], seed1_internal_state_value[52], 
	seed1_internal_state_value[51], seed1_internal_state_value[50], 
	seed1_internal_state_value[49], seed1_internal_state_value[48], 
	seed1_internal_state_value[47], seed1_internal_state_value[46], 
	seed1_internal_state_value[45], seed1_internal_state_value[44], 
	seed1_internal_state_value[43], seed1_internal_state_value[42], 
	seed1_internal_state_value[41], seed1_internal_state_value[40], 
	seed1_internal_state_value[39], seed1_internal_state_value[38], 
	seed1_internal_state_value[37], seed1_internal_state_value[36], 
	seed1_internal_state_value[35], seed1_internal_state_value[34], 
	seed1_internal_state_value[33], seed1_internal_state_value[32], 
	seed1_internal_state_value[31], seed1_internal_state_value[30], 
	seed1_internal_state_value[29], seed1_internal_state_value[28], 
	seed1_internal_state_value[27], seed1_internal_state_value[26], 
	seed1_internal_state_value[25], seed1_internal_state_value[24], 
	seed1_internal_state_value[23], seed1_internal_state_value[22], 
	seed1_internal_state_value[21], seed1_internal_state_value[20], 
	seed1_internal_state_value[19], seed1_internal_state_value[18], 
	seed1_internal_state_value[17], seed1_internal_state_value[16], 
	seed1_internal_state_value[15], seed1_internal_state_value[14], 
	seed1_internal_state_value[13], seed1_internal_state_value[12], 
	seed1_internal_state_value[11], seed1_internal_state_value[10], 
	seed1_internal_state_value[9], seed1_internal_state_value[8], 
	seed1_internal_state_value[7], seed1_internal_state_value[6], 
	seed1_internal_state_value[5], seed1_internal_state_value[4], 
	seed1_internal_state_value[3], seed1_internal_state_value[2], 
	seed1_internal_state_value[1], seed1_internal_state_value[0]});
ixc_assign_48 _zz_strnp_2 ( { \seed_life[0][47] , \seed_life[0][46] , 
	\seed_life[0][45] , \seed_life[0][44] , \seed_life[0][43] , 
	\seed_life[0][42] , \seed_life[0][41] , \seed_life[0][40] , 
	\seed_life[0][39] , \seed_life[0][38] , \seed_life[0][37] , 
	\seed_life[0][36] , \seed_life[0][35] , \seed_life[0][34] , 
	\seed_life[0][33] , \seed_life[0][32] , \seed_life[0][31] , 
	\seed_life[0][30] , \seed_life[0][29] , \seed_life[0][28] , 
	\seed_life[0][27] , \seed_life[0][26] , \seed_life[0][25] , 
	\seed_life[0][24] , \seed_life[0][23] , \seed_life[0][22] , 
	\seed_life[0][21] , \seed_life[0][20] , \seed_life[0][19] , 
	\seed_life[0][18] , \seed_life[0][17] , \seed_life[0][16] , 
	\seed_life[0][15] , \seed_life[0][14] , \seed_life[0][13] , 
	\seed_life[0][12] , \seed_life[0][11] , \seed_life[0][10] , 
	\seed_life[0][9] , \seed_life[0][8] , \seed_life[0][7] , 
	\seed_life[0][6] , \seed_life[0][5] , \seed_life[0][4] , 
	\seed_life[0][3] , \seed_life[0][2] , \seed_life[0][1] , 
	\seed_life[0][0] }, seed0_reseed_interval[47:0]);
ixc_assign_48 _zz_strnp_3 ( { \seed_life[1][47] , \seed_life[1][46] , 
	\seed_life[1][45] , \seed_life[1][44] , \seed_life[1][43] , 
	\seed_life[1][42] , \seed_life[1][41] , \seed_life[1][40] , 
	\seed_life[1][39] , \seed_life[1][38] , \seed_life[1][37] , 
	\seed_life[1][36] , \seed_life[1][35] , \seed_life[1][34] , 
	\seed_life[1][33] , \seed_life[1][32] , \seed_life[1][31] , 
	\seed_life[1][30] , \seed_life[1][29] , \seed_life[1][28] , 
	\seed_life[1][27] , \seed_life[1][26] , \seed_life[1][25] , 
	\seed_life[1][24] , \seed_life[1][23] , \seed_life[1][22] , 
	\seed_life[1][21] , \seed_life[1][20] , \seed_life[1][19] , 
	\seed_life[1][18] , \seed_life[1][17] , \seed_life[1][16] , 
	\seed_life[1][15] , \seed_life[1][14] , \seed_life[1][13] , 
	\seed_life[1][12] , \seed_life[1][11] , \seed_life[1][10] , 
	\seed_life[1][9] , \seed_life[1][8] , \seed_life[1][7] , 
	\seed_life[1][6] , \seed_life[1][5] , \seed_life[1][4] , 
	\seed_life[1][3] , \seed_life[1][2] , \seed_life[1][1] , 
	\seed_life[1][0] }, seed1_reseed_interval[47:0]);
ixc_assign _zz_strnp_4 ( \seed_valid[0][0] , seed0_valid);
ixc_assign _zz_strnp_5 ( \seed_valid[1][0] , seed1_valid);
Q_AN03 U764 ( .A0(seed0_valid), .A1(seed_expired), .A2(n655), .Z(seed0_invalidate));
Q_AN03 U765 ( .A0(seed1_valid), .A1(seed_expired), .A2(seed_entry[0]), .Z(seed1_invalidate));
Q_NR02 U766 ( .A0(seed0_valid), .A1(seed1_valid), .Z(drng_seed_expired));
Q_OR02 U767 ( .A0(seed0_invalidate), .A1(seed1_invalidate), .Z(stat_drbg_reseed));
Q_AN03 U768 ( .A0(n2), .A1(n3), .A2(n4), .Z(n654));
Q_AN03 U769 ( .A0(n5), .A1(n6), .A2(n7), .Z(n653));
Q_AN03 U770 ( .A0(n8), .A1(n9), .A2(n10), .Z(n652));
Q_AN03 U771 ( .A0(n11), .A1(n12), .A2(n13), .Z(n651));
Q_AN03 U772 ( .A0(n14), .A1(n15), .A2(n16), .Z(n650));
Q_AN03 U773 ( .A0(n17), .A1(n18), .A2(n19), .Z(n649));
Q_AN03 U774 ( .A0(n20), .A1(n21), .A2(n22), .Z(n648));
Q_AN03 U775 ( .A0(n23), .A1(n24), .A2(n25), .Z(n647));
Q_AN03 U776 ( .A0(n26), .A1(n27), .A2(n28), .Z(n646));
Q_AN03 U777 ( .A0(n29), .A1(n30), .A2(n31), .Z(n645));
Q_AN03 U778 ( .A0(n32), .A1(n33), .A2(n34), .Z(n644));
Q_AN03 U779 ( .A0(n35), .A1(n36), .A2(n37), .Z(n643));
Q_AN03 U780 ( .A0(n38), .A1(n39), .A2(n40), .Z(n642));
Q_AN03 U781 ( .A0(n41), .A1(n42), .A2(n43), .Z(n641));
Q_AN03 U782 ( .A0(n44), .A1(n45), .A2(n46), .Z(n640));
Q_AN03 U783 ( .A0(n47), .A1(n48), .A2(n49), .Z(n639));
Q_AN03 U784 ( .A0(n654), .A1(n653), .A2(n652), .Z(n638));
Q_AN03 U785 ( .A0(n651), .A1(n650), .A2(n649), .Z(n637));
Q_AN03 U786 ( .A0(n648), .A1(n647), .A2(n646), .Z(n636));
Q_AN03 U787 ( .A0(n645), .A1(n644), .A2(n643), .Z(n635));
Q_AN03 U788 ( .A0(n642), .A1(n641), .A2(n640), .Z(n634));
Q_AN03 U789 ( .A0(n639), .A1(n638), .A2(n637), .Z(n633));
Q_AN03 U790 ( .A0(n636), .A1(n635), .A2(n634), .Z(n632));
Q_AN02 U791 ( .A0(n633), .A1(n632), .Z(drng_health_test));
ixc_assign _zz_strnp_6 ( _zy_simnet_drng_health_fail_0_w$, drng_health_fail);
ixc_assign _zz_strnp_7 ( _zy_simnet_seed_valid_3_w$, n435);
ixc_assign_384 _zz_strnp_8 ( _zy_simnet_seed_4_w$[0:383], { n50, n51, n52, n53, 
	n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, 
	n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
	n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
	n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
	n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, 
	n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, 
	n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, 
	n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
	n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
	n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
	n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, 
	n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
	n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
	n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, 
	n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, 
	n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, 
	n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, 
	n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, 
	n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, 
	n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
	n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
	n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, 
	n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, 
	n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, 
	n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, 
	n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, 
	n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, 
	n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, 
	n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, 
	n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, 
	n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, 
	n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, 
	n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
	n427, n428, n429, n430, n431, n432, n433});
ixc_assign_48 _zz_strnp_9 ( _zy_simnet_seed_life_5_w$[0:47], { n2, n3, n4, n5, 
	n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, 
	n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, 
	n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
	n48, n49});
cr_kme_aes_256_drng drng ( .seed_expired( seed_expired), .drng_valid( 
	drng_valid), .drng_256_out( drng_256_out_pre[127:0]), 
	.drng_fifo_overflow( _zy_simnet_dio_1), .drng_fifo_underflow( 
	_zy_simnet_dio_2), .drng_idle( drng_idle), .start( 
	_zy_simnet_seed_valid_3_w$), .seed( _zy_simnet_seed_4_w$[0:383]), 
	.seed_life( _zy_simnet_seed_life_5_w$[0:47]), .drng_ack( drng_ack), 
	.clk( clk), .rst_n( rst_n));
Q_XOR2 U797 ( .A0(n439), .A1(n655), .Z(n440));
Q_FDP4EP \drng_256_last_REG[127] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[127]), .Q(drng_256_last[127]));
Q_INV U799 ( .A(rst_n), .Z(n656));
Q_FDP4EP \drng_256_last_REG[126] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[126]), .Q(drng_256_last[126]));
Q_FDP4EP \drng_256_last_REG[125] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[125]), .Q(drng_256_last[125]));
Q_FDP4EP \drng_256_last_REG[124] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[124]), .Q(drng_256_last[124]));
Q_FDP4EP \drng_256_last_REG[123] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[123]), .Q(drng_256_last[123]));
Q_FDP4EP \drng_256_last_REG[122] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[122]), .Q(drng_256_last[122]));
Q_FDP4EP \drng_256_last_REG[121] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[121]), .Q(drng_256_last[121]));
Q_FDP4EP \drng_256_last_REG[120] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[120]), .Q(drng_256_last[120]));
Q_FDP4EP \drng_256_last_REG[119] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[119]), .Q(drng_256_last[119]));
Q_FDP4EP \drng_256_last_REG[118] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[118]), .Q(drng_256_last[118]));
Q_FDP4EP \drng_256_last_REG[117] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[117]), .Q(drng_256_last[117]));
Q_FDP4EP \drng_256_last_REG[116] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[116]), .Q(drng_256_last[116]));
Q_FDP4EP \drng_256_last_REG[115] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[115]), .Q(drng_256_last[115]));
Q_FDP4EP \drng_256_last_REG[114] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[114]), .Q(drng_256_last[114]));
Q_FDP4EP \drng_256_last_REG[113] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[113]), .Q(drng_256_last[113]));
Q_FDP4EP \drng_256_last_REG[112] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[112]), .Q(drng_256_last[112]));
Q_FDP4EP \drng_256_last_REG[111] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[111]), .Q(drng_256_last[111]));
Q_FDP4EP \drng_256_last_REG[110] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[110]), .Q(drng_256_last[110]));
Q_FDP4EP \drng_256_last_REG[109] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[109]), .Q(drng_256_last[109]));
Q_FDP4EP \drng_256_last_REG[108] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[108]), .Q(drng_256_last[108]));
Q_FDP4EP \drng_256_last_REG[107] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[107]), .Q(drng_256_last[107]));
Q_FDP4EP \drng_256_last_REG[106] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[106]), .Q(drng_256_last[106]));
Q_FDP4EP \drng_256_last_REG[105] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[105]), .Q(drng_256_last[105]));
Q_FDP4EP \drng_256_last_REG[104] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[104]), .Q(drng_256_last[104]));
Q_FDP4EP \drng_256_last_REG[103] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[103]), .Q(drng_256_last[103]));
Q_FDP4EP \drng_256_last_REG[102] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[102]), .Q(drng_256_last[102]));
Q_FDP4EP \drng_256_last_REG[101] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[101]), .Q(drng_256_last[101]));
Q_FDP4EP \drng_256_last_REG[100] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[100]), .Q(drng_256_last[100]));
Q_FDP4EP \drng_256_last_REG[99] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[99]), .Q(drng_256_last[99]));
Q_FDP4EP \drng_256_last_REG[98] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[98]), .Q(drng_256_last[98]));
Q_FDP4EP \drng_256_last_REG[97] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[97]), .Q(drng_256_last[97]));
Q_FDP4EP \drng_256_last_REG[96] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[96]), .Q(drng_256_last[96]));
Q_FDP4EP \drng_256_last_REG[95] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[95]), .Q(drng_256_last[95]));
Q_FDP4EP \drng_256_last_REG[94] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[94]), .Q(drng_256_last[94]));
Q_FDP4EP \drng_256_last_REG[93] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[93]), .Q(drng_256_last[93]));
Q_FDP4EP \drng_256_last_REG[92] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[92]), .Q(drng_256_last[92]));
Q_FDP4EP \drng_256_last_REG[91] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[91]), .Q(drng_256_last[91]));
Q_FDP4EP \drng_256_last_REG[90] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[90]), .Q(drng_256_last[90]));
Q_FDP4EP \drng_256_last_REG[89] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[89]), .Q(drng_256_last[89]));
Q_FDP4EP \drng_256_last_REG[88] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[88]), .Q(drng_256_last[88]));
Q_FDP4EP \drng_256_last_REG[87] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[87]), .Q(drng_256_last[87]));
Q_FDP4EP \drng_256_last_REG[86] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[86]), .Q(drng_256_last[86]));
Q_FDP4EP \drng_256_last_REG[85] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[85]), .Q(drng_256_last[85]));
Q_FDP4EP \drng_256_last_REG[84] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[84]), .Q(drng_256_last[84]));
Q_FDP4EP \drng_256_last_REG[83] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[83]), .Q(drng_256_last[83]));
Q_FDP4EP \drng_256_last_REG[82] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[82]), .Q(drng_256_last[82]));
Q_FDP4EP \drng_256_last_REG[81] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[81]), .Q(drng_256_last[81]));
Q_FDP4EP \drng_256_last_REG[80] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[80]), .Q(drng_256_last[80]));
Q_FDP4EP \drng_256_last_REG[79] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[79]), .Q(drng_256_last[79]));
Q_FDP4EP \drng_256_last_REG[78] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[78]), .Q(drng_256_last[78]));
Q_FDP4EP \drng_256_last_REG[77] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[77]), .Q(drng_256_last[77]));
Q_FDP4EP \drng_256_last_REG[76] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[76]), .Q(drng_256_last[76]));
Q_FDP4EP \drng_256_last_REG[75] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[75]), .Q(drng_256_last[75]));
Q_FDP4EP \drng_256_last_REG[74] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[74]), .Q(drng_256_last[74]));
Q_FDP4EP \drng_256_last_REG[73] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[73]), .Q(drng_256_last[73]));
Q_FDP4EP \drng_256_last_REG[72] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[72]), .Q(drng_256_last[72]));
Q_FDP4EP \drng_256_last_REG[71] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[71]), .Q(drng_256_last[71]));
Q_FDP4EP \drng_256_last_REG[70] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[70]), .Q(drng_256_last[70]));
Q_FDP4EP \drng_256_last_REG[69] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[69]), .Q(drng_256_last[69]));
Q_FDP4EP \drng_256_last_REG[68] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[68]), .Q(drng_256_last[68]));
Q_FDP4EP \drng_256_last_REG[67] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[67]), .Q(drng_256_last[67]));
Q_FDP4EP \drng_256_last_REG[66] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[66]), .Q(drng_256_last[66]));
Q_FDP4EP \drng_256_last_REG[65] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[65]), .Q(drng_256_last[65]));
Q_FDP4EP \drng_256_last_REG[64] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[64]), .Q(drng_256_last[64]));
Q_FDP4EP \drng_256_last_REG[63] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[63]), .Q(drng_256_last[63]));
Q_FDP4EP \drng_256_last_REG[62] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[62]), .Q(drng_256_last[62]));
Q_FDP4EP \drng_256_last_REG[61] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[61]), .Q(drng_256_last[61]));
Q_FDP4EP \drng_256_last_REG[60] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[60]), .Q(drng_256_last[60]));
Q_FDP4EP \drng_256_last_REG[59] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[59]), .Q(drng_256_last[59]));
Q_FDP4EP \drng_256_last_REG[58] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[58]), .Q(drng_256_last[58]));
Q_FDP4EP \drng_256_last_REG[57] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[57]), .Q(drng_256_last[57]));
Q_FDP4EP \drng_256_last_REG[56] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[56]), .Q(drng_256_last[56]));
Q_FDP4EP \drng_256_last_REG[55] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[55]), .Q(drng_256_last[55]));
Q_FDP4EP \drng_256_last_REG[54] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[54]), .Q(drng_256_last[54]));
Q_FDP4EP \drng_256_last_REG[53] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[53]), .Q(drng_256_last[53]));
Q_FDP4EP \drng_256_last_REG[52] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[52]), .Q(drng_256_last[52]));
Q_FDP4EP \drng_256_last_REG[51] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[51]), .Q(drng_256_last[51]));
Q_FDP4EP \drng_256_last_REG[50] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[50]), .Q(drng_256_last[50]));
Q_FDP4EP \drng_256_last_REG[49] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[49]), .Q(drng_256_last[49]));
Q_FDP4EP \drng_256_last_REG[48] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[48]), .Q(drng_256_last[48]));
Q_FDP4EP \drng_256_last_REG[47] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[47]), .Q(drng_256_last[47]));
Q_FDP4EP \drng_256_last_REG[46] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[46]), .Q(drng_256_last[46]));
Q_FDP4EP \drng_256_last_REG[45] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[45]), .Q(drng_256_last[45]));
Q_FDP4EP \drng_256_last_REG[44] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[44]), .Q(drng_256_last[44]));
Q_FDP4EP \drng_256_last_REG[43] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[43]), .Q(drng_256_last[43]));
Q_FDP4EP \drng_256_last_REG[42] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[42]), .Q(drng_256_last[42]));
Q_FDP4EP \drng_256_last_REG[41] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[41]), .Q(drng_256_last[41]));
Q_FDP4EP \drng_256_last_REG[40] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[40]), .Q(drng_256_last[40]));
Q_FDP4EP \drng_256_last_REG[39] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[39]), .Q(drng_256_last[39]));
Q_FDP4EP \drng_256_last_REG[38] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[38]), .Q(drng_256_last[38]));
Q_FDP4EP \drng_256_last_REG[37] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[37]), .Q(drng_256_last[37]));
Q_FDP4EP \drng_256_last_REG[36] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[36]), .Q(drng_256_last[36]));
Q_FDP4EP \drng_256_last_REG[35] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[35]), .Q(drng_256_last[35]));
Q_FDP4EP \drng_256_last_REG[34] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[34]), .Q(drng_256_last[34]));
Q_FDP4EP \drng_256_last_REG[33] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[33]), .Q(drng_256_last[33]));
Q_FDP4EP \drng_256_last_REG[32] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[32]), .Q(drng_256_last[32]));
Q_FDP4EP \drng_256_last_REG[31] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[31]), .Q(drng_256_last[31]));
Q_FDP4EP \drng_256_last_REG[30] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[30]), .Q(drng_256_last[30]));
Q_FDP4EP \drng_256_last_REG[29] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[29]), .Q(drng_256_last[29]));
Q_FDP4EP \drng_256_last_REG[28] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[28]), .Q(drng_256_last[28]));
Q_FDP4EP \drng_256_last_REG[27] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[27]), .Q(drng_256_last[27]));
Q_FDP4EP \drng_256_last_REG[26] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[26]), .Q(drng_256_last[26]));
Q_FDP4EP \drng_256_last_REG[25] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[25]), .Q(drng_256_last[25]));
Q_FDP4EP \drng_256_last_REG[24] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[24]), .Q(drng_256_last[24]));
Q_FDP4EP \drng_256_last_REG[23] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[23]), .Q(drng_256_last[23]));
Q_FDP4EP \drng_256_last_REG[22] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[22]), .Q(drng_256_last[22]));
Q_FDP4EP \drng_256_last_REG[21] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[21]), .Q(drng_256_last[21]));
Q_FDP4EP \drng_256_last_REG[20] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[20]), .Q(drng_256_last[20]));
Q_FDP4EP \drng_256_last_REG[19] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[19]), .Q(drng_256_last[19]));
Q_FDP4EP \drng_256_last_REG[18] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[18]), .Q(drng_256_last[18]));
Q_FDP4EP \drng_256_last_REG[17] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[17]), .Q(drng_256_last[17]));
Q_FDP4EP \drng_256_last_REG[16] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[16]), .Q(drng_256_last[16]));
Q_FDP4EP \drng_256_last_REG[15] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[15]), .Q(drng_256_last[15]));
Q_FDP4EP \drng_256_last_REG[14] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[14]), .Q(drng_256_last[14]));
Q_FDP4EP \drng_256_last_REG[13] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[13]), .Q(drng_256_last[13]));
Q_FDP4EP \drng_256_last_REG[12] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[12]), .Q(drng_256_last[12]));
Q_FDP4EP \drng_256_last_REG[11] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[11]), .Q(drng_256_last[11]));
Q_FDP4EP \drng_256_last_REG[10] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[10]), .Q(drng_256_last[10]));
Q_FDP4EP \drng_256_last_REG[9] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[9]), .Q(drng_256_last[9]));
Q_FDP4EP \drng_256_last_REG[8] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[8]), .Q(drng_256_last[8]));
Q_FDP4EP \drng_256_last_REG[7] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[7]), .Q(drng_256_last[7]));
Q_FDP4EP \drng_256_last_REG[6] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[6]), .Q(drng_256_last[6]));
Q_FDP4EP \drng_256_last_REG[5] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[5]), .Q(drng_256_last[5]));
Q_FDP4EP \drng_256_last_REG[4] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[4]), .Q(drng_256_last[4]));
Q_FDP4EP \drng_256_last_REG[3] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[3]), .Q(drng_256_last[3]));
Q_FDP4EP \drng_256_last_REG[2] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[2]), .Q(drng_256_last[2]));
Q_FDP4EP \drng_256_last_REG[1] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[1]), .Q(drng_256_last[1]));
Q_FDP4EP \drng_256_last_REG[0] ( .CK(clk), .CE(drng_ack), .R(n656), .D(drng_256_out[0]), .Q(drng_256_last[0]));
Q_FDP4EP drng_first_REG  ( .CK(clk), .CE(drng_ack), .R(n656), .D(n1), .Q(drng_first));
Q_FDP4EP drng_health_fail_REG  ( .CK(clk), .CE(drng_ack), .R(n656), .D(n436), .Q(drng_health_fail));
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m1 "seed 1 383 0 1 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m2 "seed_life 1 47 0 1 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m3 "seed_valid 1 0 0 1 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_NON_CMM "3"
endmodule
