module ifsyn_conns();
wire i_0_0_0, ip_0_0_0;
// quickturn name_map i_0_0_0  kme_tb.apb_xactor._zyixc_port_0_0_isf
// quickturn name_map ip_0_0_0 xcva_top.IXC_GFIFO.ISF.pvec[0]
  wire o_0_0_0, op_0_0_0;
// quickturn name_map op_0_0_0 xcva_top.IXC_GFIFO.OSF.pvecEv[0]
// quickturn name_map o_0_0_0  kme_tb.apb_xactor._zyixc_port_0_0_osf
wire i_0_1_1, ip_0_1_1;
// quickturn name_map i_0_1_1  kme_tb.apb_xactor._zyixc_port_0_1_isf
// quickturn name_map ip_0_1_1 xcva_top.IXC_GFIFO.ISF.pvec[1]
  wire o_0_1_1, op_0_1_1;
// quickturn name_map op_0_1_1 xcva_top.IXC_GFIFO.OSF.pvecEv[1]
// quickturn name_map o_0_1_1  kme_tb.apb_xactor._zyixc_port_0_1_osf
  wire o_1_0_0, op_1_0_0;
// quickturn name_map op_1_0_0 xcva_top.IXC_GFIFO.OSF1.pvecEv[0]
// quickturn name_map o_1_0_0  kme_tb.kme_dut.u_cr_kme_core.\kme_is_core.txc_axi_intf .u_cr_fifo_wrap2.\ram_fifo.u_nx_fifo_ram_1r1w .fifo_ctrl._zyixc_port_1_0_osf
  wire o_1_1_0, op_1_1_0;
// quickturn name_map op_1_1_0 xcva_top.IXC_GFIFO.OSF1.pvecEv[1]
// quickturn name_map o_1_1_0  kme_tb.kme_dut.u_cr_kme_core.\kme_is_core.cceip_encrypt_kop_fifo .ram_fifo.\ram_fifo.u_nx_fifo_ram_1r1w .fifo_ctrl._zyixc_port_1_0_osf
  wire o_1_2_0, op_1_2_0;
// quickturn name_map op_1_2_0 xcva_top.IXC_GFIFO.OSF1.pvecEv[2]
// quickturn name_map o_1_2_0  kme_tb.kme_dut.u_cr_kme_core.\kme_is_core.cceip_validate_kop_fifo .ram_fifo.\ram_fifo.u_nx_fifo_ram_1r1w .fifo_ctrl._zyixc_port_1_0_osf
  wire o_1_3_0, op_1_3_0;
// quickturn name_map op_1_3_0 xcva_top.IXC_GFIFO.OSF1.pvecEv[3]
// quickturn name_map o_1_3_0  kme_tb.kme_dut.u_cr_kme_core.\kme_is_core.cceip0_key_tlv_rsm .u_cr_tlvp2_rsm.u_cr_fifo_wrap2_tob.\ram_fifo.u_nx_fifo_ram_1r1w .fifo_ctrl._zyixc_port_1_0_osf
  wire o_1_4_0, op_1_4_0;
// quickturn name_map op_1_4_0 xcva_top.IXC_GFIFO.OSF1.pvecEv[4]
// quickturn name_map o_1_4_0  kme_tb.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cceip0.u_nx_credit_manager._zyixc_port_1_0_osf
  wire o_1_5_1, op_1_5_1;
// quickturn name_map op_1_5_1 xcva_top.IXC_GFIFO.OSF1.pvecEv[5]
// quickturn name_map o_1_5_1  kme_tb.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cceip0.u_nx_credit_manager._zyixc_port_1_1_osf
  wire o_1_6_0, op_1_6_0;
// quickturn name_map op_1_6_0 xcva_top.IXC_GFIFO.OSF1.pvecEv[6]
// quickturn name_map o_1_6_0  kme_tb.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cceip1.u_nx_credit_manager._zyixc_port_1_0_osf
  wire o_1_7_1, op_1_7_1;
// quickturn name_map op_1_7_1 xcva_top.IXC_GFIFO.OSF1.pvecEv[7]
// quickturn name_map o_1_7_1  kme_tb.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cceip1.u_nx_credit_manager._zyixc_port_1_1_osf
  wire o_1_8_0, op_1_8_0;
// quickturn name_map op_1_8_0 xcva_top.IXC_GFIFO.OSF1.pvecEv[8]
// quickturn name_map o_1_8_0  kme_tb.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cceip2.u_nx_credit_manager._zyixc_port_1_0_osf
  wire o_1_9_1, op_1_9_1;
// quickturn name_map op_1_9_1 xcva_top.IXC_GFIFO.OSF1.pvecEv[9]
// quickturn name_map o_1_9_1  kme_tb.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cceip2.u_nx_credit_manager._zyixc_port_1_1_osf
  wire o_1_10_0, op_1_10_0;
// quickturn name_map op_1_10_0 xcva_top.IXC_GFIFO.OSF1.pvecEv[10]
// quickturn name_map o_1_10_0  kme_tb.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cceip3.u_nx_credit_manager._zyixc_port_1_0_osf
  wire o_1_11_1, op_1_11_1;
// quickturn name_map op_1_11_1 xcva_top.IXC_GFIFO.OSF1.pvecEv[11]
// quickturn name_map o_1_11_1  kme_tb.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cceip3.u_nx_credit_manager._zyixc_port_1_1_osf
  wire o_1_12_0, op_1_12_0;
// quickturn name_map op_1_12_0 xcva_top.IXC_GFIFO.OSF1.pvecEv[12]
// quickturn name_map o_1_12_0  kme_tb.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cddip0.u_nx_credit_manager._zyixc_port_1_0_osf
  wire o_1_13_1, op_1_13_1;
// quickturn name_map op_1_13_1 xcva_top.IXC_GFIFO.OSF1.pvecEv[13]
// quickturn name_map o_1_13_1  kme_tb.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cddip0.u_nx_credit_manager._zyixc_port_1_1_osf
  wire o_1_14_0, op_1_14_0;
// quickturn name_map op_1_14_0 xcva_top.IXC_GFIFO.OSF1.pvecEv[14]
// quickturn name_map o_1_14_0  kme_tb.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cddip1.u_nx_credit_manager._zyixc_port_1_0_osf
  wire o_1_15_1, op_1_15_1;
// quickturn name_map op_1_15_1 xcva_top.IXC_GFIFO.OSF1.pvecEv[15]
// quickturn name_map o_1_15_1  kme_tb.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cddip1.u_nx_credit_manager._zyixc_port_1_1_osf
  wire o_1_16_0, op_1_16_0;
// quickturn name_map op_1_16_0 xcva_top.IXC_GFIFO.OSF1.pvecEv[16]
// quickturn name_map o_1_16_0  kme_tb.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cddip2.u_nx_credit_manager._zyixc_port_1_0_osf
  wire o_1_17_1, op_1_17_1;
// quickturn name_map op_1_17_1 xcva_top.IXC_GFIFO.OSF1.pvecEv[17]
// quickturn name_map o_1_17_1  kme_tb.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cddip2.u_nx_credit_manager._zyixc_port_1_1_osf
  wire o_1_18_0, op_1_18_0;
// quickturn name_map op_1_18_0 xcva_top.IXC_GFIFO.OSF1.pvecEv[18]
// quickturn name_map o_1_18_0  kme_tb.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cddip3.u_nx_credit_manager._zyixc_port_1_0_osf
  wire o_1_19_1, op_1_19_1;
// quickturn name_map op_1_19_1 xcva_top.IXC_GFIFO.OSF1.pvecEv[19]
// quickturn name_map o_1_19_1  kme_tb.kme_dut.u_cr_kme_regfile.u_nx_interface_monitor_cddip3.u_nx_credit_manager._zyixc_port_1_1_osf
  ixc_assign isfasgn_0_0_0(i_0_0_0, ip_0_0_0);
  ixc_assign osfasgn_0_0_0(op_0_0_0, o_0_0_0);
  ixc_assign isfasgn_0_1_1(i_0_1_1, ip_0_1_1);
  ixc_assign osfasgn_0_1_1(op_0_1_1, o_0_1_1);
  ixc_assign osfasgn_1_0_0(op_1_0_0, o_1_0_0);
  ixc_assign osfasgn_1_1_0(op_1_1_0, o_1_1_0);
  ixc_assign osfasgn_1_2_0(op_1_2_0, o_1_2_0);
  ixc_assign osfasgn_1_3_0(op_1_3_0, o_1_3_0);
  ixc_assign osfasgn_1_4_0(op_1_4_0, o_1_4_0);
  ixc_assign osfasgn_1_5_1(op_1_5_1, o_1_5_1);
  ixc_assign osfasgn_1_6_0(op_1_6_0, o_1_6_0);
  ixc_assign osfasgn_1_7_1(op_1_7_1, o_1_7_1);
  ixc_assign osfasgn_1_8_0(op_1_8_0, o_1_8_0);
  ixc_assign osfasgn_1_9_1(op_1_9_1, o_1_9_1);
  ixc_assign osfasgn_1_10_0(op_1_10_0, o_1_10_0);
  ixc_assign osfasgn_1_11_1(op_1_11_1, o_1_11_1);
  ixc_assign osfasgn_1_12_0(op_1_12_0, o_1_12_0);
  ixc_assign osfasgn_1_13_1(op_1_13_1, o_1_13_1);
  ixc_assign osfasgn_1_14_0(op_1_14_0, o_1_14_0);
  ixc_assign osfasgn_1_15_1(op_1_15_1, o_1_15_1);
  ixc_assign osfasgn_1_16_0(op_1_16_0, o_1_16_0);
  ixc_assign osfasgn_1_17_1(op_1_17_1, o_1_17_1);
  ixc_assign osfasgn_1_18_0(op_1_18_0, o_1_18_0);
  ixc_assign osfasgn_1_19_1(op_1_19_1, o_1_19_1);
endmodule