// xc_work/v/140.sv
// /lan/cva_rel/ixcom23h1/23.03.131.s001/tools.lnx86/etc/ixcom/IXCSF.sv:556
// NOTE: This file corresponds to a module in the Hardware/DUT partition.
`timescale 1ps/1ps
 (* upf_always_on = 1, _2_state_ = 1 *) module IXC_PTXTOP;
tri0  xptRtn;
bit callEvOn;
wire  callEv;
wire  uClk;
wire  hasPTX;
bit [1:0] dly ;
// pragma CVASTRPROP MODULE IXC_PTXTOP PROP_IXCOM_MOD TRUE
endmodule

