architecture module of ixc_sfifo_bind_4_2 is

begin
end module;
