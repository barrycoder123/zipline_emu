
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
`_2_ (* upf_always_on = 1 *) 
module ixc_sfifo_port_32_0 ( call, iarg, oarg, tid, fen, CiData, CtId, CoData, 
	CoDataEn, CoDataLen);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output call;
`_2_ output [31:0] iarg;
input [0:0] oarg;
input [21:0] tid;
`_2_ output fen;
input [511:0] CiData;
input [21:0] CtId;
output [511:0] CoData;
output CoDataEn;
output [3:0] CoDataLen;
wire fclk;
`_2_ wire fenN;
`_2_ wire callr;
`_2_ wire callrN;
`_2_ wire [15:0] argl;
`_2_ wire [15:0] arglN;
`_2_ wire [0:0] lden;
`_2_ wire [0:0] ldenN;
wire [31:0] i;
`_2_ wire [511:0] oargB;
`_2_ wire oen;
`_2_ wire [15:0] opktl;
`_2_ wire [0:0] sten;
`_2_ wire [3:0] wlen;
`_2_ wire oState;
Q_FDP0UA U0 ( .D(callrN), .QTFCLK( ), .Q(callr));
Q_FDP0UA U1 ( .D(arglN[15]), .QTFCLK( ), .Q(argl[15]));
Q_FDP0UA U2 ( .D(arglN[14]), .QTFCLK( ), .Q(argl[14]));
Q_FDP0UA U3 ( .D(arglN[13]), .QTFCLK( ), .Q(argl[13]));
Q_FDP0UA U4 ( .D(arglN[12]), .QTFCLK( ), .Q(argl[12]));
Q_FDP0UA U5 ( .D(arglN[11]), .QTFCLK( ), .Q(argl[11]));
Q_FDP0UA U6 ( .D(arglN[10]), .QTFCLK( ), .Q(argl[10]));
Q_FDP0UA U7 ( .D(arglN[9]), .QTFCLK( ), .Q(argl[9]));
Q_FDP0UA U8 ( .D(arglN[8]), .QTFCLK( ), .Q(argl[8]));
Q_FDP0UA U9 ( .D(arglN[7]), .QTFCLK( ), .Q(argl[7]));
Q_FDP0UA U10 ( .D(arglN[6]), .QTFCLK( ), .Q(argl[6]));
Q_FDP0UA U11 ( .D(arglN[5]), .QTFCLK( ), .Q(argl[5]));
Q_FDP0UA U12 ( .D(arglN[4]), .QTFCLK( ), .Q(argl[4]));
Q_FDP0UA U13 ( .D(arglN[3]), .QTFCLK( ), .Q(argl[3]));
Q_FDP0UA U14 ( .D(arglN[2]), .QTFCLK( ), .Q(argl[2]));
Q_FDP0UA U15 ( .D(arglN[1]), .QTFCLK( ), .Q(argl[1]));
Q_FDP0UA U16 ( .D(arglN[0]), .QTFCLK( ), .Q(argl[0]));
Q_FDP0UA U17 ( .D(ldenN[0]), .QTFCLK( ), .Q(lden[0]));
Q_FDP0UA U18 ( .D(fenN), .QTFCLK( ), .Q(fen));
Q_NR02 U19 ( .A0(n2), .A1(n3), .Z(n6));
Q_OR02 U20 ( .A0(n6), .A1(n5), .Z(n4));
Q_INV U21 ( .A(n4), .Z(fenN));
Q_XNR2 U22 ( .A0(n4), .A1(callr), .Z(callrN));
Q_AN02 U23 ( .A0(n5), .A1(n7), .Z(arglN[15]));
Q_AN02 U24 ( .A0(n5), .A1(n9), .Z(arglN[14]));
Q_AN02 U25 ( .A0(n5), .A1(n11), .Z(arglN[13]));
Q_AN02 U26 ( .A0(n5), .A1(n13), .Z(arglN[12]));
Q_AN02 U27 ( .A0(n5), .A1(n15), .Z(arglN[11]));
Q_AN02 U28 ( .A0(n5), .A1(n17), .Z(arglN[10]));
Q_AN02 U29 ( .A0(n5), .A1(n19), .Z(arglN[9]));
Q_AN02 U30 ( .A0(n5), .A1(n21), .Z(arglN[8]));
Q_AN02 U31 ( .A0(n5), .A1(n23), .Z(arglN[7]));
Q_AN02 U32 ( .A0(n5), .A1(n25), .Z(arglN[6]));
Q_AN02 U33 ( .A0(n5), .A1(n27), .Z(arglN[5]));
Q_AN02 U34 ( .A0(n5), .A1(n29), .Z(arglN[4]));
Q_AN02 U35 ( .A0(n5), .A1(n31), .Z(arglN[3]));
Q_AN02 U36 ( .A0(n5), .A1(n33), .Z(arglN[2]));
Q_AN02 U37 ( .A0(n5), .A1(n35), .Z(arglN[1]));
Q_AN02 U38 ( .A0(n5), .A1(n36), .Z(arglN[0]));
Q_INV U39 ( .A(n5), .Z(ldenN[0]));
Q_XNR2 U40 ( .A0(argl[15]), .A1(n8), .Z(n7));
Q_OR02 U41 ( .A0(argl[14]), .A1(n10), .Z(n8));
Q_XNR2 U42 ( .A0(argl[14]), .A1(n10), .Z(n9));
Q_OR02 U43 ( .A0(argl[13]), .A1(n12), .Z(n10));
Q_XNR2 U44 ( .A0(argl[13]), .A1(n12), .Z(n11));
Q_OR02 U45 ( .A0(argl[12]), .A1(n14), .Z(n12));
Q_XNR2 U46 ( .A0(argl[12]), .A1(n14), .Z(n13));
Q_OR02 U47 ( .A0(argl[11]), .A1(n16), .Z(n14));
Q_XNR2 U48 ( .A0(argl[11]), .A1(n16), .Z(n15));
Q_OR02 U49 ( .A0(argl[10]), .A1(n18), .Z(n16));
Q_XNR2 U50 ( .A0(argl[10]), .A1(n18), .Z(n17));
Q_OR02 U51 ( .A0(argl[9]), .A1(n20), .Z(n18));
Q_XNR2 U52 ( .A0(argl[9]), .A1(n20), .Z(n19));
Q_OR02 U53 ( .A0(argl[8]), .A1(n22), .Z(n20));
Q_XNR2 U54 ( .A0(argl[8]), .A1(n22), .Z(n21));
Q_OR02 U55 ( .A0(argl[7]), .A1(n24), .Z(n22));
Q_XNR2 U56 ( .A0(argl[7]), .A1(n24), .Z(n23));
Q_OR02 U57 ( .A0(argl[6]), .A1(n26), .Z(n24));
Q_XNR2 U58 ( .A0(argl[6]), .A1(n26), .Z(n25));
Q_OR02 U59 ( .A0(argl[5]), .A1(n28), .Z(n26));
Q_XNR2 U60 ( .A0(argl[5]), .A1(n28), .Z(n27));
Q_OR02 U61 ( .A0(argl[4]), .A1(n30), .Z(n28));
Q_XNR2 U62 ( .A0(argl[4]), .A1(n30), .Z(n29));
Q_OR02 U63 ( .A0(argl[3]), .A1(n32), .Z(n30));
Q_XNR2 U64 ( .A0(argl[3]), .A1(n32), .Z(n31));
Q_OR02 U65 ( .A0(argl[2]), .A1(n34), .Z(n32));
Q_XNR2 U66 ( .A0(argl[2]), .A1(n34), .Z(n33));
Q_OR02 U67 ( .A0(argl[1]), .A1(argl[0]), .Z(n34));
Q_XNR2 U68 ( .A0(argl[1]), .A1(argl[0]), .Z(n35));
Q_INV U69 ( .A(argl[0]), .Z(n36));
Q_OA21 U70 ( .A0(n37), .A1(n38), .B0(n2), .Z(n5));
Q_OR03 U71 ( .A0(n39), .A1(argl[1]), .A2(n40), .Z(n38));
Q_OR02 U72 ( .A0(argl[3]), .A1(argl[2]), .Z(n39));
Q_OR03 U73 ( .A0(argl[7]), .A1(argl[6]), .A2(n41), .Z(n40));
Q_OR02 U74 ( .A0(argl[5]), .A1(argl[4]), .Z(n41));
Q_OR03 U75 ( .A0(n42), .A1(n43), .A2(n44), .Z(n37));
Q_OR02 U76 ( .A0(argl[11]), .A1(argl[10]), .Z(n42));
Q_OR02 U77 ( .A0(argl[9]), .A1(argl[8]), .Z(n43));
Q_OR03 U78 ( .A0(argl[15]), .A1(argl[14]), .A2(n45), .Z(n44));
Q_OR02 U79 ( .A0(argl[13]), .A1(argl[12]), .Z(n45));
Q_OR02 U80 ( .A0(n47), .A1(n46), .Z(n2));
Q_OR03 U81 ( .A0(n50), .A1(n49), .A2(n48), .Z(n46));
Q_OR03 U82 ( .A0(argl[0]), .A1(n52), .A2(n51), .Z(n47));
Q_OR03 U83 ( .A0(argl[3]), .A1(argl[2]), .A2(argl[1]), .Z(n48));
Q_OR03 U84 ( .A0(argl[6]), .A1(argl[5]), .A2(argl[4]), .Z(n49));
Q_OR03 U85 ( .A0(argl[9]), .A1(argl[8]), .A2(argl[7]), .Z(n50));
Q_OR03 U86 ( .A0(argl[12]), .A1(argl[11]), .A2(argl[10]), .Z(n51));
Q_OR03 U87 ( .A0(argl[15]), .A1(argl[14]), .A2(argl[13]), .Z(n52));
Q_INV U88 ( .A(xc_top.GFReset), .Z(n53));
Q_AN03 U89 ( .A0(n55), .A1(n54), .A2(n53), .Z(n3));
Q_AN03 U90 ( .A0(n58), .A1(n57), .A2(n56), .Z(n54));
Q_AN03 U91 ( .A0(n61), .A1(n60), .A2(n59), .Z(n55));
Q_AN03 U92 ( .A0(n85), .A1(n63), .A2(n62), .Z(n56));
Q_AN03 U93 ( .A0(n82), .A1(n83), .A2(n84), .Z(n57));
Q_AN03 U94 ( .A0(n79), .A1(n80), .A2(n81), .Z(n58));
Q_AN03 U95 ( .A0(n76), .A1(n77), .A2(n78), .Z(n59));
Q_AN03 U96 ( .A0(n73), .A1(n74), .A2(n75), .Z(n60));
Q_AN03 U97 ( .A0(n70), .A1(n71), .A2(n72), .Z(n61));
Q_AN03 U98 ( .A0(n67), .A1(n68), .A2(n69), .Z(n62));
Q_AN03 U99 ( .A0(n64), .A1(n65), .A2(n66), .Z(n63));
Q_XNR2 U100 ( .A0(CtId[21]), .A1(tid[21]), .Z(n64));
Q_XNR2 U101 ( .A0(CtId[20]), .A1(tid[20]), .Z(n65));
Q_XNR2 U102 ( .A0(CtId[19]), .A1(tid[19]), .Z(n66));
Q_XNR2 U103 ( .A0(CtId[18]), .A1(tid[18]), .Z(n67));
Q_XNR2 U104 ( .A0(CtId[17]), .A1(tid[17]), .Z(n68));
Q_XNR2 U105 ( .A0(CtId[16]), .A1(tid[16]), .Z(n69));
Q_XNR2 U106 ( .A0(CtId[15]), .A1(tid[15]), .Z(n70));
Q_XNR2 U107 ( .A0(CtId[14]), .A1(tid[14]), .Z(n71));
Q_XNR2 U108 ( .A0(CtId[13]), .A1(tid[13]), .Z(n72));
Q_XNR2 U109 ( .A0(CtId[12]), .A1(tid[12]), .Z(n73));
Q_XNR2 U110 ( .A0(CtId[11]), .A1(tid[11]), .Z(n74));
Q_XNR2 U111 ( .A0(CtId[10]), .A1(tid[10]), .Z(n75));
Q_XNR2 U112 ( .A0(CtId[9]), .A1(tid[9]), .Z(n76));
Q_XNR2 U113 ( .A0(CtId[8]), .A1(tid[8]), .Z(n77));
Q_XNR2 U114 ( .A0(CtId[7]), .A1(tid[7]), .Z(n78));
Q_XNR2 U115 ( .A0(CtId[6]), .A1(tid[6]), .Z(n79));
Q_XNR2 U116 ( .A0(CtId[5]), .A1(tid[5]), .Z(n80));
Q_XNR2 U117 ( .A0(CtId[4]), .A1(tid[4]), .Z(n81));
Q_XNR2 U118 ( .A0(CtId[3]), .A1(tid[3]), .Z(n82));
Q_XNR2 U119 ( .A0(CtId[2]), .A1(tid[2]), .Z(n83));
Q_XNR2 U120 ( .A0(CtId[1]), .A1(tid[1]), .Z(n84));
Q_XNR2 U121 ( .A0(CtId[0]), .A1(tid[0]), .Z(n85));
Q_LDP0 \iarg_REG[0] ( .G(lden[0]), .D(CiData[0]), .Q(iarg[0]), .QN( ));
Q_LDP0 \iarg_REG[1] ( .G(lden[0]), .D(CiData[1]), .Q(iarg[1]), .QN( ));
Q_LDP0 \iarg_REG[2] ( .G(lden[0]), .D(CiData[2]), .Q(iarg[2]), .QN( ));
Q_LDP0 \iarg_REG[3] ( .G(lden[0]), .D(CiData[3]), .Q(iarg[3]), .QN( ));
Q_LDP0 \iarg_REG[4] ( .G(lden[0]), .D(CiData[4]), .Q(iarg[4]), .QN( ));
Q_LDP0 \iarg_REG[5] ( .G(lden[0]), .D(CiData[5]), .Q(iarg[5]), .QN( ));
Q_LDP0 \iarg_REG[6] ( .G(lden[0]), .D(CiData[6]), .Q(iarg[6]), .QN( ));
Q_LDP0 \iarg_REG[7] ( .G(lden[0]), .D(CiData[7]), .Q(iarg[7]), .QN( ));
Q_LDP0 \iarg_REG[8] ( .G(lden[0]), .D(CiData[8]), .Q(iarg[8]), .QN( ));
Q_LDP0 \iarg_REG[9] ( .G(lden[0]), .D(CiData[9]), .Q(iarg[9]), .QN( ));
Q_LDP0 \iarg_REG[10] ( .G(lden[0]), .D(CiData[10]), .Q(iarg[10]), .QN( ));
Q_LDP0 \iarg_REG[11] ( .G(lden[0]), .D(CiData[11]), .Q(iarg[11]), .QN( ));
Q_LDP0 \iarg_REG[12] ( .G(lden[0]), .D(CiData[12]), .Q(iarg[12]), .QN( ));
Q_LDP0 \iarg_REG[13] ( .G(lden[0]), .D(CiData[13]), .Q(iarg[13]), .QN( ));
Q_LDP0 \iarg_REG[14] ( .G(lden[0]), .D(CiData[14]), .Q(iarg[14]), .QN( ));
Q_LDP0 \iarg_REG[15] ( .G(lden[0]), .D(CiData[15]), .Q(iarg[15]), .QN( ));
Q_LDP0 \iarg_REG[16] ( .G(lden[0]), .D(CiData[16]), .Q(iarg[16]), .QN( ));
Q_LDP0 \iarg_REG[17] ( .G(lden[0]), .D(CiData[17]), .Q(iarg[17]), .QN( ));
Q_LDP0 \iarg_REG[18] ( .G(lden[0]), .D(CiData[18]), .Q(iarg[18]), .QN( ));
Q_LDP0 \iarg_REG[19] ( .G(lden[0]), .D(CiData[19]), .Q(iarg[19]), .QN( ));
Q_LDP0 \iarg_REG[20] ( .G(lden[0]), .D(CiData[20]), .Q(iarg[20]), .QN( ));
Q_LDP0 \iarg_REG[21] ( .G(lden[0]), .D(CiData[21]), .Q(iarg[21]), .QN( ));
Q_LDP0 \iarg_REG[22] ( .G(lden[0]), .D(CiData[22]), .Q(iarg[22]), .QN( ));
Q_LDP0 \iarg_REG[23] ( .G(lden[0]), .D(CiData[23]), .Q(iarg[23]), .QN( ));
Q_LDP0 \iarg_REG[24] ( .G(lden[0]), .D(CiData[24]), .Q(iarg[24]), .QN( ));
Q_LDP0 \iarg_REG[25] ( .G(lden[0]), .D(CiData[25]), .Q(iarg[25]), .QN( ));
Q_LDP0 \iarg_REG[26] ( .G(lden[0]), .D(CiData[26]), .Q(iarg[26]), .QN( ));
Q_LDP0 \iarg_REG[27] ( .G(lden[0]), .D(CiData[27]), .Q(iarg[27]), .QN( ));
Q_LDP0 \iarg_REG[28] ( .G(lden[0]), .D(CiData[28]), .Q(iarg[28]), .QN( ));
Q_LDP0 \iarg_REG[29] ( .G(lden[0]), .D(CiData[29]), .Q(iarg[29]), .QN( ));
Q_LDP0 \iarg_REG[30] ( .G(lden[0]), .D(CiData[30]), .Q(iarg[30]), .QN( ));
Q_LDP0 \iarg_REG[31] ( .G(lden[0]), .D(CiData[31]), .Q(iarg[31]), .QN( ));
Q_PULSE U154 ( .A(callr), .Z(call));
Q_NOT_TOUCH _zzqnthw ( .sig());
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE "ixc_sfifo_port"
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE_LIB "IXCOM_TEMP_LIBRARY"
// pragma CVASTRPROP MODULE HDLICE PROP_IXCOM_MOD TRUE
endmodule
