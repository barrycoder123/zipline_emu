
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
`_2_ (* upf_always_on = 1 *) 
module ixc_context_read_2048 ( rdata);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
input [2047:0] rdata;
supply1 n1;
supply0 n2;
Q_NOT_TOUCH _zzqnthw ( .sig());
`ifdef CBV

reg [511:0] _zymem [0:3];
always @(n2 or rdata[511] or rdata[510] or rdata[509] or rdata[508]
 or rdata[507] or rdata[506] or rdata[505] or rdata[504] or rdata[503] or rdata[502] or rdata[501] or rdata[500]
 or rdata[499] or rdata[498] or rdata[497] or rdata[496] or rdata[495] or rdata[494] or rdata[493] or rdata[492]
 or rdata[491] or rdata[490] or rdata[489] or rdata[488] or rdata[487] or rdata[486] or rdata[485] or rdata[484]
 or rdata[483] or rdata[482] or rdata[481] or rdata[480] or rdata[479] or rdata[478] or rdata[477] or rdata[476]
 or rdata[475] or rdata[474] or rdata[473] or rdata[472] or rdata[471] or rdata[470] or rdata[469] or rdata[468]
 or rdata[467] or rdata[466] or rdata[465] or rdata[464] or rdata[463] or rdata[462] or rdata[461] or rdata[460]
 or rdata[459] or rdata[458] or rdata[457] or rdata[456] or rdata[455] or rdata[454] or rdata[453] or rdata[452]
 or rdata[451] or rdata[450] or rdata[449] or rdata[448] or rdata[447] or rdata[446] or rdata[445] or rdata[444]
 or rdata[443] or rdata[442] or rdata[441] or rdata[440] or rdata[439] or rdata[438] or rdata[437] or rdata[436]
 or rdata[435] or rdata[434] or rdata[433] or rdata[432] or rdata[431] or rdata[430] or rdata[429] or rdata[428]
 or rdata[427] or rdata[426] or rdata[425] or rdata[424] or rdata[423] or rdata[422] or rdata[421] or rdata[420]
 or rdata[419] or rdata[418] or rdata[417] or rdata[416] or rdata[415] or rdata[414] or rdata[413] or rdata[412]
 or rdata[411] or rdata[410] or rdata[409] or rdata[408] or rdata[407] or rdata[406] or rdata[405] or rdata[404]
 or rdata[403] or rdata[402] or rdata[401] or rdata[400] or rdata[399] or rdata[398] or rdata[397] or rdata[396]
 or rdata[395] or rdata[394] or rdata[393] or rdata[392] or rdata[391] or rdata[390] or rdata[389] or rdata[388]
 or rdata[387] or rdata[386] or rdata[385] or rdata[384] or rdata[383] or rdata[382] or rdata[381] or rdata[380]
 or rdata[379] or rdata[378] or rdata[377] or rdata[376] or rdata[375] or rdata[374] or rdata[373] or rdata[372]
 or rdata[371] or rdata[370] or rdata[369] or rdata[368] or rdata[367] or rdata[366] or rdata[365] or rdata[364]
 or rdata[363] or rdata[362] or rdata[361] or rdata[360] or rdata[359] or rdata[358] or rdata[357] or rdata[356]
 or rdata[355] or rdata[354] or rdata[353] or rdata[352] or rdata[351] or rdata[350] or rdata[349] or rdata[348]
 or rdata[347] or rdata[346] or rdata[345] or rdata[344] or rdata[343] or rdata[342] or rdata[341] or rdata[340]
 or rdata[339] or rdata[338] or rdata[337] or rdata[336] or rdata[335] or rdata[334] or rdata[333] or rdata[332]
 or rdata[331] or rdata[330] or rdata[329] or rdata[328] or rdata[327] or rdata[326] or rdata[325] or rdata[324]
 or rdata[323] or rdata[322] or rdata[321] or rdata[320] or rdata[319] or rdata[318] or rdata[317] or rdata[316]
 or rdata[315] or rdata[314] or rdata[313] or rdata[312] or rdata[311] or rdata[310] or rdata[309] or rdata[308]
 or rdata[307] or rdata[306] or rdata[305] or rdata[304] or rdata[303] or rdata[302] or rdata[301] or rdata[300]
 or rdata[299] or rdata[298] or rdata[297] or rdata[296] or rdata[295] or rdata[294] or rdata[293] or rdata[292]
 or rdata[291] or rdata[290] or rdata[289] or rdata[288] or rdata[287] or rdata[286] or rdata[285] or rdata[284]
 or rdata[283] or rdata[282] or rdata[281] or rdata[280] or rdata[279] or rdata[278] or rdata[277] or rdata[276]
 or rdata[275] or rdata[274] or rdata[273] or rdata[272] or rdata[271] or rdata[270] or rdata[269] or rdata[268]
 or rdata[267] or rdata[266] or rdata[265] or rdata[264] or rdata[263] or rdata[262] or rdata[261] or rdata[260]
 or rdata[259] or rdata[258] or rdata[257] or rdata[256] or rdata[255] or rdata[254] or rdata[253] or rdata[252]
 or rdata[251] or rdata[250] or rdata[249] or rdata[248] or rdata[247] or rdata[246] or rdata[245] or rdata[244]
 or rdata[243] or rdata[242] or rdata[241] or rdata[240] or rdata[239] or rdata[238] or rdata[237] or rdata[236]
 or rdata[235] or rdata[234] or rdata[233] or rdata[232] or rdata[231] or rdata[230] or rdata[229] or rdata[228]
 or rdata[227] or rdata[226] or rdata[225] or rdata[224] or rdata[223] or rdata[222] or rdata[221] or rdata[220]
 or rdata[219] or rdata[218] or rdata[217] or rdata[216] or rdata[215] or rdata[214] or rdata[213] or rdata[212]
 or rdata[211] or rdata[210] or rdata[209] or rdata[208] or rdata[207] or rdata[206] or rdata[205] or rdata[204]
 or rdata[203] or rdata[202] or rdata[201] or rdata[200] or rdata[199] or rdata[198] or rdata[197] or rdata[196]
 or rdata[195] or rdata[194] or rdata[193] or rdata[192] or rdata[191] or rdata[190] or rdata[189] or rdata[188]
 or rdata[187] or rdata[186] or rdata[185] or rdata[184] or rdata[183] or rdata[182] or rdata[181] or rdata[180]
 or rdata[179] or rdata[178] or rdata[177] or rdata[176] or rdata[175] or rdata[174] or rdata[173] or rdata[172]
 or rdata[171] or rdata[170] or rdata[169] or rdata[168] or rdata[167] or rdata[166] or rdata[165] or rdata[164]
 or rdata[163] or rdata[162] or rdata[161] or rdata[160] or rdata[159] or rdata[158] or rdata[157] or rdata[156]
 or rdata[155] or rdata[154] or rdata[153] or rdata[152] or rdata[151] or rdata[150] or rdata[149] or rdata[148]
 or rdata[147] or rdata[146] or rdata[145] or rdata[144] or rdata[143] or rdata[142] or rdata[141] or rdata[140]
 or rdata[139] or rdata[138] or rdata[137] or rdata[136] or rdata[135] or rdata[134] or rdata[133] or rdata[132]
 or rdata[131] or rdata[130] or rdata[129] or rdata[128] or rdata[127] or rdata[126] or rdata[125] or rdata[124]
 or rdata[123] or rdata[122] or rdata[121] or rdata[120] or rdata[119] or rdata[118] or rdata[117] or rdata[116]
 or rdata[115] or rdata[114] or rdata[113] or rdata[112] or rdata[111] or rdata[110] or rdata[109] or rdata[108]
 or rdata[107] or rdata[106] or rdata[105] or rdata[104] or rdata[103] or rdata[102] or rdata[101] or rdata[100]
 or rdata[99] or rdata[98] or rdata[97] or rdata[96] or rdata[95] or rdata[94] or rdata[93] or rdata[92]
 or rdata[91] or rdata[90] or rdata[89] or rdata[88] or rdata[87] or rdata[86] or rdata[85] or rdata[84]
 or rdata[83] or rdata[82] or rdata[81] or rdata[80] or rdata[79] or rdata[78] or rdata[77] or rdata[76]
 or rdata[75] or rdata[74] or rdata[73] or rdata[72] or rdata[71] or rdata[70] or rdata[69] or rdata[68]
 or rdata[67] or rdata[66] or rdata[65] or rdata[64] or rdata[63] or rdata[62] or rdata[61] or rdata[60]
 or rdata[59] or rdata[58] or rdata[57] or rdata[56] or rdata[55] or rdata[54] or rdata[53] or rdata[52]
 or rdata[51] or rdata[50] or rdata[49] or rdata[48] or rdata[47] or rdata[46] or rdata[45] or rdata[44]
 or rdata[43] or rdata[42] or rdata[41] or rdata[40] or rdata[39] or rdata[38] or rdata[37] or rdata[36]
 or rdata[35] or rdata[34] or rdata[33] or rdata[32] or rdata[31] or rdata[30] or rdata[29] or rdata[28]
 or rdata[27] or rdata[26] or rdata[25] or rdata[24] or rdata[23] or rdata[22] or rdata[21] or rdata[20]
 or rdata[19] or rdata[18] or rdata[17] or rdata[16] or rdata[15] or rdata[14] or rdata[13] or rdata[12]
 or rdata[11] or rdata[10] or rdata[9] or rdata[8] or rdata[7] or rdata[6] or rdata[5] or rdata[4]
 or rdata[3] or rdata[2] or rdata[1] or rdata[0] or n1 or rdata[1023] or rdata[1022] or rdata[1021]
 or rdata[1020] or rdata[1019] or rdata[1018] or rdata[1017] or rdata[1016] or rdata[1015] or rdata[1014] or rdata[1013]
 or rdata[1012] or rdata[1011] or rdata[1010] or rdata[1009] or rdata[1008] or rdata[1007] or rdata[1006] or rdata[1005]
 or rdata[1004] or rdata[1003] or rdata[1002] or rdata[1001] or rdata[1000] or rdata[999] or rdata[998] or rdata[997]
 or rdata[996] or rdata[995] or rdata[994] or rdata[993] or rdata[992] or rdata[991] or rdata[990] or rdata[989]
 or rdata[988] or rdata[987] or rdata[986] or rdata[985] or rdata[984] or rdata[983] or rdata[982] or rdata[981]
 or rdata[980] or rdata[979] or rdata[978] or rdata[977] or rdata[976] or rdata[975] or rdata[974] or rdata[973]
 or rdata[972] or rdata[971] or rdata[970] or rdata[969] or rdata[968] or rdata[967] or rdata[966] or rdata[965]
 or rdata[964] or rdata[963] or rdata[962] or rdata[961] or rdata[960] or rdata[959] or rdata[958] or rdata[957]
 or rdata[956] or rdata[955] or rdata[954] or rdata[953] or rdata[952] or rdata[951] or rdata[950] or rdata[949]
 or rdata[948] or rdata[947] or rdata[946] or rdata[945] or rdata[944] or rdata[943] or rdata[942] or rdata[941]
 or rdata[940] or rdata[939] or rdata[938] or rdata[937] or rdata[936] or rdata[935] or rdata[934] or rdata[933]
 or rdata[932] or rdata[931] or rdata[930] or rdata[929] or rdata[928] or rdata[927] or rdata[926] or rdata[925]
 or rdata[924] or rdata[923] or rdata[922] or rdata[921] or rdata[920] or rdata[919] or rdata[918] or rdata[917]
 or rdata[916] or rdata[915] or rdata[914] or rdata[913] or rdata[912] or rdata[911] or rdata[910] or rdata[909]
 or rdata[908] or rdata[907] or rdata[906] or rdata[905] or rdata[904] or rdata[903] or rdata[902] or rdata[901]
 or rdata[900] or rdata[899] or rdata[898] or rdata[897] or rdata[896] or rdata[895] or rdata[894] or rdata[893]
 or rdata[892] or rdata[891] or rdata[890] or rdata[889] or rdata[888] or rdata[887] or rdata[886] or rdata[885]
 or rdata[884] or rdata[883] or rdata[882] or rdata[881] or rdata[880] or rdata[879] or rdata[878] or rdata[877]
 or rdata[876] or rdata[875] or rdata[874] or rdata[873] or rdata[872] or rdata[871] or rdata[870] or rdata[869]
 or rdata[868] or rdata[867] or rdata[866] or rdata[865] or rdata[864] or rdata[863] or rdata[862] or rdata[861]
 or rdata[860] or rdata[859] or rdata[858] or rdata[857] or rdata[856] or rdata[855] or rdata[854] or rdata[853]
 or rdata[852] or rdata[851] or rdata[850] or rdata[849] or rdata[848] or rdata[847] or rdata[846] or rdata[845]
 or rdata[844] or rdata[843] or rdata[842] or rdata[841] or rdata[840] or rdata[839] or rdata[838] or rdata[837]
 or rdata[836] or rdata[835] or rdata[834] or rdata[833] or rdata[832] or rdata[831] or rdata[830] or rdata[829]
 or rdata[828] or rdata[827] or rdata[826] or rdata[825] or rdata[824] or rdata[823] or rdata[822] or rdata[821]
 or rdata[820] or rdata[819] or rdata[818] or rdata[817] or rdata[816] or rdata[815] or rdata[814] or rdata[813]
 or rdata[812] or rdata[811] or rdata[810] or rdata[809] or rdata[808] or rdata[807] or rdata[806] or rdata[805]
 or rdata[804] or rdata[803] or rdata[802] or rdata[801] or rdata[800] or rdata[799] or rdata[798] or rdata[797]
 or rdata[796] or rdata[795] or rdata[794] or rdata[793] or rdata[792] or rdata[791] or rdata[790] or rdata[789]
 or rdata[788] or rdata[787] or rdata[786] or rdata[785] or rdata[784] or rdata[783] or rdata[782] or rdata[781]
 or rdata[780] or rdata[779] or rdata[778] or rdata[777] or rdata[776] or rdata[775] or rdata[774] or rdata[773]
 or rdata[772] or rdata[771] or rdata[770] or rdata[769] or rdata[768] or rdata[767] or rdata[766] or rdata[765]
 or rdata[764] or rdata[763] or rdata[762] or rdata[761] or rdata[760] or rdata[759] or rdata[758] or rdata[757]
 or rdata[756] or rdata[755] or rdata[754] or rdata[753] or rdata[752] or rdata[751] or rdata[750] or rdata[749]
 or rdata[748] or rdata[747] or rdata[746] or rdata[745] or rdata[744] or rdata[743] or rdata[742] or rdata[741]
 or rdata[740] or rdata[739] or rdata[738] or rdata[737] or rdata[736] or rdata[735] or rdata[734] or rdata[733]
 or rdata[732] or rdata[731] or rdata[730] or rdata[729] or rdata[728] or rdata[727] or rdata[726] or rdata[725]
 or rdata[724] or rdata[723] or rdata[722] or rdata[721] or rdata[720] or rdata[719] or rdata[718] or rdata[717]
 or rdata[716] or rdata[715] or rdata[714] or rdata[713] or rdata[712] or rdata[711] or rdata[710] or rdata[709]
 or rdata[708] or rdata[707] or rdata[706] or rdata[705] or rdata[704] or rdata[703] or rdata[702] or rdata[701]
 or rdata[700] or rdata[699] or rdata[698] or rdata[697] or rdata[696] or rdata[695] or rdata[694] or rdata[693]
 or rdata[692] or rdata[691] or rdata[690] or rdata[689] or rdata[688] or rdata[687] or rdata[686] or rdata[685]
 or rdata[684] or rdata[683] or rdata[682] or rdata[681] or rdata[680] or rdata[679] or rdata[678] or rdata[677]
 or rdata[676] or rdata[675] or rdata[674] or rdata[673] or rdata[672] or rdata[671] or rdata[670] or rdata[669]
 or rdata[668] or rdata[667] or rdata[666] or rdata[665] or rdata[664] or rdata[663] or rdata[662] or rdata[661]
 or rdata[660] or rdata[659] or rdata[658] or rdata[657] or rdata[656] or rdata[655] or rdata[654] or rdata[653]
 or rdata[652] or rdata[651] or rdata[650] or rdata[649] or rdata[648] or rdata[647] or rdata[646] or rdata[645]
 or rdata[644] or rdata[643] or rdata[642] or rdata[641] or rdata[640] or rdata[639] or rdata[638] or rdata[637]
 or rdata[636] or rdata[635] or rdata[634] or rdata[633] or rdata[632] or rdata[631] or rdata[630] or rdata[629]
 or rdata[628] or rdata[627] or rdata[626] or rdata[625] or rdata[624] or rdata[623] or rdata[622] or rdata[621]
 or rdata[620] or rdata[619] or rdata[618] or rdata[617] or rdata[616] or rdata[615] or rdata[614] or rdata[613]
 or rdata[612] or rdata[611] or rdata[610] or rdata[609] or rdata[608] or rdata[607] or rdata[606] or rdata[605]
 or rdata[604] or rdata[603] or rdata[602] or rdata[601] or rdata[600] or rdata[599] or rdata[598] or rdata[597]
 or rdata[596] or rdata[595] or rdata[594] or rdata[593] or rdata[592] or rdata[591] or rdata[590] or rdata[589]
 or rdata[588] or rdata[587] or rdata[586] or rdata[585] or rdata[584] or rdata[583] or rdata[582] or rdata[581]
 or rdata[580] or rdata[579] or rdata[578] or rdata[577] or rdata[576] or rdata[575] or rdata[574] or rdata[573]
 or rdata[572] or rdata[571] or rdata[570] or rdata[569] or rdata[568] or rdata[567] or rdata[566] or rdata[565]
 or rdata[564] or rdata[563] or rdata[562] or rdata[561] or rdata[560] or rdata[559] or rdata[558] or rdata[557]
 or rdata[556] or rdata[555] or rdata[554] or rdata[553] or rdata[552] or rdata[551] or rdata[550] or rdata[549]
 or rdata[548] or rdata[547] or rdata[546] or rdata[545] or rdata[544] or rdata[543] or rdata[542] or rdata[541]
 or rdata[540] or rdata[539] or rdata[538] or rdata[537] or rdata[536] or rdata[535] or rdata[534] or rdata[533]
 or rdata[532] or rdata[531] or rdata[530] or rdata[529] or rdata[528] or rdata[527] or rdata[526] or rdata[525]
 or rdata[524] or rdata[523] or rdata[522] or rdata[521] or rdata[520] or rdata[519] or rdata[518] or rdata[517]
 or rdata[516] or rdata[515] or rdata[514] or rdata[513] or rdata[512] or rdata[1535] or rdata[1534] or rdata[1533]
 or rdata[1532] or rdata[1531] or rdata[1530] or rdata[1529] or rdata[1528] or rdata[1527] or rdata[1526] or rdata[1525]
 or rdata[1524] or rdata[1523] or rdata[1522] or rdata[1521] or rdata[1520] or rdata[1519] or rdata[1518] or rdata[1517]
 or rdata[1516] or rdata[1515] or rdata[1514] or rdata[1513] or rdata[1512] or rdata[1511] or rdata[1510] or rdata[1509]
 or rdata[1508] or rdata[1507] or rdata[1506] or rdata[1505] or rdata[1504] or rdata[1503] or rdata[1502] or rdata[1501]
 or rdata[1500] or rdata[1499] or rdata[1498] or rdata[1497] or rdata[1496] or rdata[1495] or rdata[1494] or rdata[1493]
 or rdata[1492] or rdata[1491] or rdata[1490] or rdata[1489] or rdata[1488] or rdata[1487] or rdata[1486] or rdata[1485]
 or rdata[1484] or rdata[1483] or rdata[1482] or rdata[1481] or rdata[1480] or rdata[1479] or rdata[1478] or rdata[1477]
 or rdata[1476] or rdata[1475] or rdata[1474] or rdata[1473] or rdata[1472] or rdata[1471] or rdata[1470] or rdata[1469]
 or rdata[1468] or rdata[1467] or rdata[1466] or rdata[1465] or rdata[1464] or rdata[1463] or rdata[1462] or rdata[1461]
 or rdata[1460] or rdata[1459] or rdata[1458] or rdata[1457] or rdata[1456] or rdata[1455] or rdata[1454] or rdata[1453]
 or rdata[1452] or rdata[1451] or rdata[1450] or rdata[1449] or rdata[1448] or rdata[1447] or rdata[1446] or rdata[1445]
 or rdata[1444] or rdata[1443] or rdata[1442] or rdata[1441] or rdata[1440] or rdata[1439] or rdata[1438] or rdata[1437]
 or rdata[1436] or rdata[1435] or rdata[1434] or rdata[1433] or rdata[1432] or rdata[1431] or rdata[1430] or rdata[1429]
 or rdata[1428] or rdata[1427] or rdata[1426] or rdata[1425] or rdata[1424] or rdata[1423] or rdata[1422] or rdata[1421]
 or rdata[1420] or rdata[1419] or rdata[1418] or rdata[1417] or rdata[1416] or rdata[1415] or rdata[1414] or rdata[1413]
 or rdata[1412] or rdata[1411] or rdata[1410] or rdata[1409] or rdata[1408] or rdata[1407] or rdata[1406] or rdata[1405]
 or rdata[1404] or rdata[1403] or rdata[1402] or rdata[1401] or rdata[1400] or rdata[1399] or rdata[1398] or rdata[1397]
 or rdata[1396] or rdata[1395] or rdata[1394] or rdata[1393] or rdata[1392] or rdata[1391] or rdata[1390] or rdata[1389]
 or rdata[1388] or rdata[1387] or rdata[1386] or rdata[1385] or rdata[1384] or rdata[1383] or rdata[1382] or rdata[1381]
 or rdata[1380] or rdata[1379] or rdata[1378] or rdata[1377] or rdata[1376] or rdata[1375] or rdata[1374] or rdata[1373]
 or rdata[1372] or rdata[1371] or rdata[1370] or rdata[1369] or rdata[1368] or rdata[1367] or rdata[1366] or rdata[1365]
 or rdata[1364] or rdata[1363] or rdata[1362] or rdata[1361] or rdata[1360] or rdata[1359] or rdata[1358] or rdata[1357]
 or rdata[1356] or rdata[1355] or rdata[1354] or rdata[1353] or rdata[1352] or rdata[1351] or rdata[1350] or rdata[1349]
 or rdata[1348] or rdata[1347] or rdata[1346] or rdata[1345] or rdata[1344] or rdata[1343] or rdata[1342] or rdata[1341]
 or rdata[1340] or rdata[1339] or rdata[1338] or rdata[1337] or rdata[1336] or rdata[1335] or rdata[1334] or rdata[1333]
 or rdata[1332] or rdata[1331] or rdata[1330] or rdata[1329] or rdata[1328] or rdata[1327] or rdata[1326] or rdata[1325]
 or rdata[1324] or rdata[1323] or rdata[1322] or rdata[1321] or rdata[1320] or rdata[1319] or rdata[1318] or rdata[1317]
 or rdata[1316] or rdata[1315] or rdata[1314] or rdata[1313] or rdata[1312] or rdata[1311] or rdata[1310] or rdata[1309]
 or rdata[1308] or rdata[1307] or rdata[1306] or rdata[1305] or rdata[1304] or rdata[1303] or rdata[1302] or rdata[1301]
 or rdata[1300] or rdata[1299] or rdata[1298] or rdata[1297] or rdata[1296] or rdata[1295] or rdata[1294] or rdata[1293]
 or rdata[1292] or rdata[1291] or rdata[1290] or rdata[1289] or rdata[1288] or rdata[1287] or rdata[1286] or rdata[1285]
 or rdata[1284] or rdata[1283] or rdata[1282] or rdata[1281] or rdata[1280] or rdata[1279] or rdata[1278] or rdata[1277]
 or rdata[1276] or rdata[1275] or rdata[1274] or rdata[1273] or rdata[1272] or rdata[1271] or rdata[1270] or rdata[1269]
 or rdata[1268] or rdata[1267] or rdata[1266] or rdata[1265] or rdata[1264] or rdata[1263] or rdata[1262] or rdata[1261]
 or rdata[1260] or rdata[1259] or rdata[1258] or rdata[1257] or rdata[1256] or rdata[1255] or rdata[1254] or rdata[1253]
 or rdata[1252] or rdata[1251] or rdata[1250] or rdata[1249] or rdata[1248] or rdata[1247] or rdata[1246] or rdata[1245]
 or rdata[1244] or rdata[1243] or rdata[1242] or rdata[1241] or rdata[1240] or rdata[1239] or rdata[1238] or rdata[1237]
 or rdata[1236] or rdata[1235] or rdata[1234] or rdata[1233] or rdata[1232] or rdata[1231] or rdata[1230] or rdata[1229]
 or rdata[1228] or rdata[1227] or rdata[1226] or rdata[1225] or rdata[1224] or rdata[1223] or rdata[1222] or rdata[1221]
 or rdata[1220] or rdata[1219] or rdata[1218] or rdata[1217] or rdata[1216] or rdata[1215] or rdata[1214] or rdata[1213]
 or rdata[1212] or rdata[1211] or rdata[1210] or rdata[1209] or rdata[1208] or rdata[1207] or rdata[1206] or rdata[1205]
 or rdata[1204] or rdata[1203] or rdata[1202] or rdata[1201] or rdata[1200] or rdata[1199] or rdata[1198] or rdata[1197]
 or rdata[1196] or rdata[1195] or rdata[1194] or rdata[1193] or rdata[1192] or rdata[1191] or rdata[1190] or rdata[1189]
 or rdata[1188] or rdata[1187] or rdata[1186] or rdata[1185] or rdata[1184] or rdata[1183] or rdata[1182] or rdata[1181]
 or rdata[1180] or rdata[1179] or rdata[1178] or rdata[1177] or rdata[1176] or rdata[1175] or rdata[1174] or rdata[1173]
 or rdata[1172] or rdata[1171] or rdata[1170] or rdata[1169] or rdata[1168] or rdata[1167] or rdata[1166] or rdata[1165]
 or rdata[1164] or rdata[1163] or rdata[1162] or rdata[1161] or rdata[1160] or rdata[1159] or rdata[1158] or rdata[1157]
 or rdata[1156] or rdata[1155] or rdata[1154] or rdata[1153] or rdata[1152] or rdata[1151] or rdata[1150] or rdata[1149]
 or rdata[1148] or rdata[1147] or rdata[1146] or rdata[1145] or rdata[1144] or rdata[1143] or rdata[1142] or rdata[1141]
 or rdata[1140] or rdata[1139] or rdata[1138] or rdata[1137] or rdata[1136] or rdata[1135] or rdata[1134] or rdata[1133]
 or rdata[1132] or rdata[1131] or rdata[1130] or rdata[1129] or rdata[1128] or rdata[1127] or rdata[1126] or rdata[1125]
 or rdata[1124] or rdata[1123] or rdata[1122] or rdata[1121] or rdata[1120] or rdata[1119] or rdata[1118] or rdata[1117]
 or rdata[1116] or rdata[1115] or rdata[1114] or rdata[1113] or rdata[1112] or rdata[1111] or rdata[1110] or rdata[1109]
 or rdata[1108] or rdata[1107] or rdata[1106] or rdata[1105] or rdata[1104] or rdata[1103] or rdata[1102] or rdata[1101]
 or rdata[1100] or rdata[1099] or rdata[1098] or rdata[1097] or rdata[1096] or rdata[1095] or rdata[1094] or rdata[1093]
 or rdata[1092] or rdata[1091] or rdata[1090] or rdata[1089] or rdata[1088] or rdata[1087] or rdata[1086] or rdata[1085]
 or rdata[1084] or rdata[1083] or rdata[1082] or rdata[1081] or rdata[1080] or rdata[1079] or rdata[1078] or rdata[1077]
 or rdata[1076] or rdata[1075] or rdata[1074] or rdata[1073] or rdata[1072] or rdata[1071] or rdata[1070] or rdata[1069]
 or rdata[1068] or rdata[1067] or rdata[1066] or rdata[1065] or rdata[1064] or rdata[1063] or rdata[1062] or rdata[1061]
 or rdata[1060] or rdata[1059] or rdata[1058] or rdata[1057] or rdata[1056] or rdata[1055] or rdata[1054] or rdata[1053]
 or rdata[1052] or rdata[1051] or rdata[1050] or rdata[1049] or rdata[1048] or rdata[1047] or rdata[1046] or rdata[1045]
 or rdata[1044] or rdata[1043] or rdata[1042] or rdata[1041] or rdata[1040] or rdata[1039] or rdata[1038] or rdata[1037]
 or rdata[1036] or rdata[1035] or rdata[1034] or rdata[1033] or rdata[1032] or rdata[1031] or rdata[1030] or rdata[1029]
 or rdata[1028] or rdata[1027] or rdata[1026] or rdata[1025] or rdata[1024] or rdata[2047] or rdata[2046] or rdata[2045]
 or rdata[2044] or rdata[2043] or rdata[2042] or rdata[2041] or rdata[2040] or rdata[2039] or rdata[2038] or rdata[2037]
 or rdata[2036] or rdata[2035] or rdata[2034] or rdata[2033] or rdata[2032] or rdata[2031] or rdata[2030] or rdata[2029]
 or rdata[2028] or rdata[2027] or rdata[2026] or rdata[2025] or rdata[2024] or rdata[2023] or rdata[2022] or rdata[2021]
 or rdata[2020] or rdata[2019] or rdata[2018] or rdata[2017] or rdata[2016] or rdata[2015] or rdata[2014] or rdata[2013]
 or rdata[2012] or rdata[2011] or rdata[2010] or rdata[2009] or rdata[2008] or rdata[2007] or rdata[2006] or rdata[2005]
 or rdata[2004] or rdata[2003] or rdata[2002] or rdata[2001] or rdata[2000] or rdata[1999] or rdata[1998] or rdata[1997]
 or rdata[1996] or rdata[1995] or rdata[1994] or rdata[1993] or rdata[1992] or rdata[1991] or rdata[1990] or rdata[1989]
 or rdata[1988] or rdata[1987] or rdata[1986] or rdata[1985] or rdata[1984] or rdata[1983] or rdata[1982] or rdata[1981]
 or rdata[1980] or rdata[1979] or rdata[1978] or rdata[1977] or rdata[1976] or rdata[1975] or rdata[1974] or rdata[1973]
 or rdata[1972] or rdata[1971] or rdata[1970] or rdata[1969] or rdata[1968] or rdata[1967] or rdata[1966] or rdata[1965]
 or rdata[1964] or rdata[1963] or rdata[1962] or rdata[1961] or rdata[1960] or rdata[1959] or rdata[1958] or rdata[1957]
 or rdata[1956] or rdata[1955] or rdata[1954] or rdata[1953] or rdata[1952] or rdata[1951] or rdata[1950] or rdata[1949]
 or rdata[1948] or rdata[1947] or rdata[1946] or rdata[1945] or rdata[1944] or rdata[1943] or rdata[1942] or rdata[1941]
 or rdata[1940] or rdata[1939] or rdata[1938] or rdata[1937] or rdata[1936] or rdata[1935] or rdata[1934] or rdata[1933]
 or rdata[1932] or rdata[1931] or rdata[1930] or rdata[1929] or rdata[1928] or rdata[1927] or rdata[1926] or rdata[1925]
 or rdata[1924] or rdata[1923] or rdata[1922] or rdata[1921] or rdata[1920] or rdata[1919] or rdata[1918] or rdata[1917]
 or rdata[1916] or rdata[1915] or rdata[1914] or rdata[1913] or rdata[1912] or rdata[1911] or rdata[1910] or rdata[1909]
 or rdata[1908] or rdata[1907] or rdata[1906] or rdata[1905] or rdata[1904] or rdata[1903] or rdata[1902] or rdata[1901]
 or rdata[1900] or rdata[1899] or rdata[1898] or rdata[1897] or rdata[1896] or rdata[1895] or rdata[1894] or rdata[1893]
 or rdata[1892] or rdata[1891] or rdata[1890] or rdata[1889] or rdata[1888] or rdata[1887] or rdata[1886] or rdata[1885]
 or rdata[1884] or rdata[1883] or rdata[1882] or rdata[1881] or rdata[1880] or rdata[1879] or rdata[1878] or rdata[1877]
 or rdata[1876] or rdata[1875] or rdata[1874] or rdata[1873] or rdata[1872] or rdata[1871] or rdata[1870] or rdata[1869]
 or rdata[1868] or rdata[1867] or rdata[1866] or rdata[1865] or rdata[1864] or rdata[1863] or rdata[1862] or rdata[1861]
 or rdata[1860] or rdata[1859] or rdata[1858] or rdata[1857] or rdata[1856] or rdata[1855] or rdata[1854] or rdata[1853]
 or rdata[1852] or rdata[1851] or rdata[1850] or rdata[1849] or rdata[1848] or rdata[1847] or rdata[1846] or rdata[1845]
 or rdata[1844] or rdata[1843] or rdata[1842] or rdata[1841] or rdata[1840] or rdata[1839] or rdata[1838] or rdata[1837]
 or rdata[1836] or rdata[1835] or rdata[1834] or rdata[1833] or rdata[1832] or rdata[1831] or rdata[1830] or rdata[1829]
 or rdata[1828] or rdata[1827] or rdata[1826] or rdata[1825] or rdata[1824] or rdata[1823] or rdata[1822] or rdata[1821]
 or rdata[1820] or rdata[1819] or rdata[1818] or rdata[1817] or rdata[1816] or rdata[1815] or rdata[1814] or rdata[1813]
 or rdata[1812] or rdata[1811] or rdata[1810] or rdata[1809] or rdata[1808] or rdata[1807] or rdata[1806] or rdata[1805]
 or rdata[1804] or rdata[1803] or rdata[1802] or rdata[1801] or rdata[1800] or rdata[1799] or rdata[1798] or rdata[1797]
 or rdata[1796] or rdata[1795] or rdata[1794] or rdata[1793] or rdata[1792] or rdata[1791] or rdata[1790] or rdata[1789]
 or rdata[1788] or rdata[1787] or rdata[1786] or rdata[1785] or rdata[1784] or rdata[1783] or rdata[1782] or rdata[1781]
 or rdata[1780] or rdata[1779] or rdata[1778] or rdata[1777] or rdata[1776] or rdata[1775] or rdata[1774] or rdata[1773]
 or rdata[1772] or rdata[1771] or rdata[1770] or rdata[1769] or rdata[1768] or rdata[1767] or rdata[1766] or rdata[1765]
 or rdata[1764] or rdata[1763] or rdata[1762] or rdata[1761] or rdata[1760] or rdata[1759] or rdata[1758] or rdata[1757]
 or rdata[1756] or rdata[1755] or rdata[1754] or rdata[1753] or rdata[1752] or rdata[1751] or rdata[1750] or rdata[1749]
 or rdata[1748] or rdata[1747] or rdata[1746] or rdata[1745] or rdata[1744] or rdata[1743] or rdata[1742] or rdata[1741]
 or rdata[1740] or rdata[1739] or rdata[1738] or rdata[1737] or rdata[1736] or rdata[1735] or rdata[1734] or rdata[1733]
 or rdata[1732] or rdata[1731] or rdata[1730] or rdata[1729] or rdata[1728] or rdata[1727] or rdata[1726] or rdata[1725]
 or rdata[1724] or rdata[1723] or rdata[1722] or rdata[1721] or rdata[1720] or rdata[1719] or rdata[1718] or rdata[1717]
 or rdata[1716] or rdata[1715] or rdata[1714] or rdata[1713] or rdata[1712] or rdata[1711] or rdata[1710] or rdata[1709]
 or rdata[1708] or rdata[1707] or rdata[1706] or rdata[1705] or rdata[1704] or rdata[1703] or rdata[1702] or rdata[1701]
 or rdata[1700] or rdata[1699] or rdata[1698] or rdata[1697] or rdata[1696] or rdata[1695] or rdata[1694] or rdata[1693]
 or rdata[1692] or rdata[1691] or rdata[1690] or rdata[1689] or rdata[1688] or rdata[1687] or rdata[1686] or rdata[1685]
 or rdata[1684] or rdata[1683] or rdata[1682] or rdata[1681] or rdata[1680] or rdata[1679] or rdata[1678] or rdata[1677]
 or rdata[1676] or rdata[1675] or rdata[1674] or rdata[1673] or rdata[1672] or rdata[1671] or rdata[1670] or rdata[1669]
 or rdata[1668] or rdata[1667] or rdata[1666] or rdata[1665] or rdata[1664] or rdata[1663] or rdata[1662] or rdata[1661]
 or rdata[1660] or rdata[1659] or rdata[1658] or rdata[1657] or rdata[1656] or rdata[1655] or rdata[1654] or rdata[1653]
 or rdata[1652] or rdata[1651] or rdata[1650] or rdata[1649] or rdata[1648] or rdata[1647] or rdata[1646] or rdata[1645]
 or rdata[1644] or rdata[1643] or rdata[1642] or rdata[1641] or rdata[1640] or rdata[1639] or rdata[1638] or rdata[1637]
 or rdata[1636] or rdata[1635] or rdata[1634] or rdata[1633] or rdata[1632] or rdata[1631] or rdata[1630] or rdata[1629]
 or rdata[1628] or rdata[1627] or rdata[1626] or rdata[1625] or rdata[1624] or rdata[1623] or rdata[1622] or rdata[1621]
 or rdata[1620] or rdata[1619] or rdata[1618] or rdata[1617] or rdata[1616] or rdata[1615] or rdata[1614] or rdata[1613]
 or rdata[1612] or rdata[1611] or rdata[1610] or rdata[1609] or rdata[1608] or rdata[1607] or rdata[1606] or rdata[1605]
 or rdata[1604] or rdata[1603] or rdata[1602] or rdata[1601] or rdata[1600] or rdata[1599] or rdata[1598] or rdata[1597]
 or rdata[1596] or rdata[1595] or rdata[1594] or rdata[1593] or rdata[1592] or rdata[1591] or rdata[1590] or rdata[1589]
 or rdata[1588] or rdata[1587] or rdata[1586] or rdata[1585] or rdata[1584] or rdata[1583] or rdata[1582] or rdata[1581]
 or rdata[1580] or rdata[1579] or rdata[1578] or rdata[1577] or rdata[1576] or rdata[1575] or rdata[1574] or rdata[1573]
 or rdata[1572] or rdata[1571] or rdata[1570] or rdata[1569] or rdata[1568] or rdata[1567] or rdata[1566] or rdata[1565]
 or rdata[1564] or rdata[1563] or rdata[1562] or rdata[1561] or rdata[1560] or rdata[1559] or rdata[1558] or rdata[1557]
 or rdata[1556] or rdata[1555] or rdata[1554] or rdata[1553] or rdata[1552] or rdata[1551] or rdata[1550] or rdata[1549]
 or rdata[1548] or rdata[1547] or rdata[1546] or rdata[1545] or rdata[1544] or rdata[1543] or rdata[1542] or rdata[1541]
 or rdata[1540] or rdata[1539] or rdata[1538] or rdata[1537] or rdata[1536])
#0 begin
if (n1)
_zymem[{n2, n2}] =
{rdata[511], rdata[510], rdata[509], rdata[508], rdata[507],
 rdata[506], rdata[505], rdata[504], rdata[503], rdata[502], rdata[501], rdata[500], rdata[499],
 rdata[498], rdata[497], rdata[496], rdata[495], rdata[494], rdata[493], rdata[492], rdata[491],
 rdata[490], rdata[489], rdata[488], rdata[487], rdata[486], rdata[485], rdata[484], rdata[483],
 rdata[482], rdata[481], rdata[480], rdata[479], rdata[478], rdata[477], rdata[476], rdata[475],
 rdata[474], rdata[473], rdata[472], rdata[471], rdata[470], rdata[469], rdata[468], rdata[467],
 rdata[466], rdata[465], rdata[464], rdata[463], rdata[462], rdata[461], rdata[460], rdata[459],
 rdata[458], rdata[457], rdata[456], rdata[455], rdata[454], rdata[453], rdata[452], rdata[451],
 rdata[450], rdata[449], rdata[448], rdata[447], rdata[446], rdata[445], rdata[444], rdata[443],
 rdata[442], rdata[441], rdata[440], rdata[439], rdata[438], rdata[437], rdata[436], rdata[435],
 rdata[434], rdata[433], rdata[432], rdata[431], rdata[430], rdata[429], rdata[428], rdata[427],
 rdata[426], rdata[425], rdata[424], rdata[423], rdata[422], rdata[421], rdata[420], rdata[419],
 rdata[418], rdata[417], rdata[416], rdata[415], rdata[414], rdata[413], rdata[412], rdata[411],
 rdata[410], rdata[409], rdata[408], rdata[407], rdata[406], rdata[405], rdata[404], rdata[403],
 rdata[402], rdata[401], rdata[400], rdata[399], rdata[398], rdata[397], rdata[396], rdata[395],
 rdata[394], rdata[393], rdata[392], rdata[391], rdata[390], rdata[389], rdata[388], rdata[387],
 rdata[386], rdata[385], rdata[384], rdata[383], rdata[382], rdata[381], rdata[380], rdata[379],
 rdata[378], rdata[377], rdata[376], rdata[375], rdata[374], rdata[373], rdata[372], rdata[371],
 rdata[370], rdata[369], rdata[368], rdata[367], rdata[366], rdata[365], rdata[364], rdata[363],
 rdata[362], rdata[361], rdata[360], rdata[359], rdata[358], rdata[357], rdata[356], rdata[355],
 rdata[354], rdata[353], rdata[352], rdata[351], rdata[350], rdata[349], rdata[348], rdata[347],
 rdata[346], rdata[345], rdata[344], rdata[343], rdata[342], rdata[341], rdata[340], rdata[339],
 rdata[338], rdata[337], rdata[336], rdata[335], rdata[334], rdata[333], rdata[332], rdata[331],
 rdata[330], rdata[329], rdata[328], rdata[327], rdata[326], rdata[325], rdata[324], rdata[323],
 rdata[322], rdata[321], rdata[320], rdata[319], rdata[318], rdata[317], rdata[316], rdata[315],
 rdata[314], rdata[313], rdata[312], rdata[311], rdata[310], rdata[309], rdata[308], rdata[307],
 rdata[306], rdata[305], rdata[304], rdata[303], rdata[302], rdata[301], rdata[300], rdata[299],
 rdata[298], rdata[297], rdata[296], rdata[295], rdata[294], rdata[293], rdata[292], rdata[291],
 rdata[290], rdata[289], rdata[288], rdata[287], rdata[286], rdata[285], rdata[284], rdata[283],
 rdata[282], rdata[281], rdata[280], rdata[279], rdata[278], rdata[277], rdata[276], rdata[275],
 rdata[274], rdata[273], rdata[272], rdata[271], rdata[270], rdata[269], rdata[268], rdata[267],
 rdata[266], rdata[265], rdata[264], rdata[263], rdata[262], rdata[261], rdata[260], rdata[259],
 rdata[258], rdata[257], rdata[256], rdata[255], rdata[254], rdata[253], rdata[252], rdata[251],
 rdata[250], rdata[249], rdata[248], rdata[247], rdata[246], rdata[245], rdata[244], rdata[243],
 rdata[242], rdata[241], rdata[240], rdata[239], rdata[238], rdata[237], rdata[236], rdata[235],
 rdata[234], rdata[233], rdata[232], rdata[231], rdata[230], rdata[229], rdata[228], rdata[227],
 rdata[226], rdata[225], rdata[224], rdata[223], rdata[222], rdata[221], rdata[220], rdata[219],
 rdata[218], rdata[217], rdata[216], rdata[215], rdata[214], rdata[213], rdata[212], rdata[211],
 rdata[210], rdata[209], rdata[208], rdata[207], rdata[206], rdata[205], rdata[204], rdata[203],
 rdata[202], rdata[201], rdata[200], rdata[199], rdata[198], rdata[197], rdata[196], rdata[195],
 rdata[194], rdata[193], rdata[192], rdata[191], rdata[190], rdata[189], rdata[188], rdata[187],
 rdata[186], rdata[185], rdata[184], rdata[183], rdata[182], rdata[181], rdata[180], rdata[179],
 rdata[178], rdata[177], rdata[176], rdata[175], rdata[174], rdata[173], rdata[172], rdata[171],
 rdata[170], rdata[169], rdata[168], rdata[167], rdata[166], rdata[165], rdata[164], rdata[163],
 rdata[162], rdata[161], rdata[160], rdata[159], rdata[158], rdata[157], rdata[156], rdata[155],
 rdata[154], rdata[153], rdata[152], rdata[151], rdata[150], rdata[149], rdata[148], rdata[147],
 rdata[146], rdata[145], rdata[144], rdata[143], rdata[142], rdata[141], rdata[140], rdata[139],
 rdata[138], rdata[137], rdata[136], rdata[135], rdata[134], rdata[133], rdata[132], rdata[131],
 rdata[130], rdata[129], rdata[128], rdata[127], rdata[126], rdata[125], rdata[124], rdata[123],
 rdata[122], rdata[121], rdata[120], rdata[119], rdata[118], rdata[117], rdata[116], rdata[115],
 rdata[114], rdata[113], rdata[112], rdata[111], rdata[110], rdata[109], rdata[108], rdata[107],
 rdata[106], rdata[105], rdata[104], rdata[103], rdata[102], rdata[101], rdata[100], rdata[99],
 rdata[98], rdata[97], rdata[96], rdata[95], rdata[94], rdata[93], rdata[92], rdata[91],
 rdata[90], rdata[89], rdata[88], rdata[87], rdata[86], rdata[85], rdata[84], rdata[83],
 rdata[82], rdata[81], rdata[80], rdata[79], rdata[78], rdata[77], rdata[76], rdata[75],
 rdata[74], rdata[73], rdata[72], rdata[71], rdata[70], rdata[69], rdata[68], rdata[67],
 rdata[66], rdata[65], rdata[64], rdata[63], rdata[62], rdata[61], rdata[60], rdata[59],
 rdata[58], rdata[57], rdata[56], rdata[55], rdata[54], rdata[53], rdata[52], rdata[51],
 rdata[50], rdata[49], rdata[48], rdata[47], rdata[46], rdata[45], rdata[44], rdata[43],
 rdata[42], rdata[41], rdata[40], rdata[39], rdata[38], rdata[37], rdata[36], rdata[35],
 rdata[34], rdata[33], rdata[32], rdata[31], rdata[30], rdata[29], rdata[28], rdata[27],
 rdata[26], rdata[25], rdata[24], rdata[23], rdata[22], rdata[21], rdata[20], rdata[19],
 rdata[18], rdata[17], rdata[16], rdata[15], rdata[14], rdata[13], rdata[12], rdata[11],
 rdata[10], rdata[9], rdata[8], rdata[7], rdata[6], rdata[5], rdata[4], rdata[3],
 rdata[2], rdata[1], rdata[0]};
if (n1)
_zymem[{n2, n1}] =
{rdata[1023], rdata[1022], rdata[1021], rdata[1020], rdata[1019],
 rdata[1018], rdata[1017], rdata[1016], rdata[1015], rdata[1014], rdata[1013], rdata[1012], rdata[1011],
 rdata[1010], rdata[1009], rdata[1008], rdata[1007], rdata[1006], rdata[1005], rdata[1004], rdata[1003],
 rdata[1002], rdata[1001], rdata[1000], rdata[999], rdata[998], rdata[997], rdata[996], rdata[995],
 rdata[994], rdata[993], rdata[992], rdata[991], rdata[990], rdata[989], rdata[988], rdata[987],
 rdata[986], rdata[985], rdata[984], rdata[983], rdata[982], rdata[981], rdata[980], rdata[979],
 rdata[978], rdata[977], rdata[976], rdata[975], rdata[974], rdata[973], rdata[972], rdata[971],
 rdata[970], rdata[969], rdata[968], rdata[967], rdata[966], rdata[965], rdata[964], rdata[963],
 rdata[962], rdata[961], rdata[960], rdata[959], rdata[958], rdata[957], rdata[956], rdata[955],
 rdata[954], rdata[953], rdata[952], rdata[951], rdata[950], rdata[949], rdata[948], rdata[947],
 rdata[946], rdata[945], rdata[944], rdata[943], rdata[942], rdata[941], rdata[940], rdata[939],
 rdata[938], rdata[937], rdata[936], rdata[935], rdata[934], rdata[933], rdata[932], rdata[931],
 rdata[930], rdata[929], rdata[928], rdata[927], rdata[926], rdata[925], rdata[924], rdata[923],
 rdata[922], rdata[921], rdata[920], rdata[919], rdata[918], rdata[917], rdata[916], rdata[915],
 rdata[914], rdata[913], rdata[912], rdata[911], rdata[910], rdata[909], rdata[908], rdata[907],
 rdata[906], rdata[905], rdata[904], rdata[903], rdata[902], rdata[901], rdata[900], rdata[899],
 rdata[898], rdata[897], rdata[896], rdata[895], rdata[894], rdata[893], rdata[892], rdata[891],
 rdata[890], rdata[889], rdata[888], rdata[887], rdata[886], rdata[885], rdata[884], rdata[883],
 rdata[882], rdata[881], rdata[880], rdata[879], rdata[878], rdata[877], rdata[876], rdata[875],
 rdata[874], rdata[873], rdata[872], rdata[871], rdata[870], rdata[869], rdata[868], rdata[867],
 rdata[866], rdata[865], rdata[864], rdata[863], rdata[862], rdata[861], rdata[860], rdata[859],
 rdata[858], rdata[857], rdata[856], rdata[855], rdata[854], rdata[853], rdata[852], rdata[851],
 rdata[850], rdata[849], rdata[848], rdata[847], rdata[846], rdata[845], rdata[844], rdata[843],
 rdata[842], rdata[841], rdata[840], rdata[839], rdata[838], rdata[837], rdata[836], rdata[835],
 rdata[834], rdata[833], rdata[832], rdata[831], rdata[830], rdata[829], rdata[828], rdata[827],
 rdata[826], rdata[825], rdata[824], rdata[823], rdata[822], rdata[821], rdata[820], rdata[819],
 rdata[818], rdata[817], rdata[816], rdata[815], rdata[814], rdata[813], rdata[812], rdata[811],
 rdata[810], rdata[809], rdata[808], rdata[807], rdata[806], rdata[805], rdata[804], rdata[803],
 rdata[802], rdata[801], rdata[800], rdata[799], rdata[798], rdata[797], rdata[796], rdata[795],
 rdata[794], rdata[793], rdata[792], rdata[791], rdata[790], rdata[789], rdata[788], rdata[787],
 rdata[786], rdata[785], rdata[784], rdata[783], rdata[782], rdata[781], rdata[780], rdata[779],
 rdata[778], rdata[777], rdata[776], rdata[775], rdata[774], rdata[773], rdata[772], rdata[771],
 rdata[770], rdata[769], rdata[768], rdata[767], rdata[766], rdata[765], rdata[764], rdata[763],
 rdata[762], rdata[761], rdata[760], rdata[759], rdata[758], rdata[757], rdata[756], rdata[755],
 rdata[754], rdata[753], rdata[752], rdata[751], rdata[750], rdata[749], rdata[748], rdata[747],
 rdata[746], rdata[745], rdata[744], rdata[743], rdata[742], rdata[741], rdata[740], rdata[739],
 rdata[738], rdata[737], rdata[736], rdata[735], rdata[734], rdata[733], rdata[732], rdata[731],
 rdata[730], rdata[729], rdata[728], rdata[727], rdata[726], rdata[725], rdata[724], rdata[723],
 rdata[722], rdata[721], rdata[720], rdata[719], rdata[718], rdata[717], rdata[716], rdata[715],
 rdata[714], rdata[713], rdata[712], rdata[711], rdata[710], rdata[709], rdata[708], rdata[707],
 rdata[706], rdata[705], rdata[704], rdata[703], rdata[702], rdata[701], rdata[700], rdata[699],
 rdata[698], rdata[697], rdata[696], rdata[695], rdata[694], rdata[693], rdata[692], rdata[691],
 rdata[690], rdata[689], rdata[688], rdata[687], rdata[686], rdata[685], rdata[684], rdata[683],
 rdata[682], rdata[681], rdata[680], rdata[679], rdata[678], rdata[677], rdata[676], rdata[675],
 rdata[674], rdata[673], rdata[672], rdata[671], rdata[670], rdata[669], rdata[668], rdata[667],
 rdata[666], rdata[665], rdata[664], rdata[663], rdata[662], rdata[661], rdata[660], rdata[659],
 rdata[658], rdata[657], rdata[656], rdata[655], rdata[654], rdata[653], rdata[652], rdata[651],
 rdata[650], rdata[649], rdata[648], rdata[647], rdata[646], rdata[645], rdata[644], rdata[643],
 rdata[642], rdata[641], rdata[640], rdata[639], rdata[638], rdata[637], rdata[636], rdata[635],
 rdata[634], rdata[633], rdata[632], rdata[631], rdata[630], rdata[629], rdata[628], rdata[627],
 rdata[626], rdata[625], rdata[624], rdata[623], rdata[622], rdata[621], rdata[620], rdata[619],
 rdata[618], rdata[617], rdata[616], rdata[615], rdata[614], rdata[613], rdata[612], rdata[611],
 rdata[610], rdata[609], rdata[608], rdata[607], rdata[606], rdata[605], rdata[604], rdata[603],
 rdata[602], rdata[601], rdata[600], rdata[599], rdata[598], rdata[597], rdata[596], rdata[595],
 rdata[594], rdata[593], rdata[592], rdata[591], rdata[590], rdata[589], rdata[588], rdata[587],
 rdata[586], rdata[585], rdata[584], rdata[583], rdata[582], rdata[581], rdata[580], rdata[579],
 rdata[578], rdata[577], rdata[576], rdata[575], rdata[574], rdata[573], rdata[572], rdata[571],
 rdata[570], rdata[569], rdata[568], rdata[567], rdata[566], rdata[565], rdata[564], rdata[563],
 rdata[562], rdata[561], rdata[560], rdata[559], rdata[558], rdata[557], rdata[556], rdata[555],
 rdata[554], rdata[553], rdata[552], rdata[551], rdata[550], rdata[549], rdata[548], rdata[547],
 rdata[546], rdata[545], rdata[544], rdata[543], rdata[542], rdata[541], rdata[540], rdata[539],
 rdata[538], rdata[537], rdata[536], rdata[535], rdata[534], rdata[533], rdata[532], rdata[531],
 rdata[530], rdata[529], rdata[528], rdata[527], rdata[526], rdata[525], rdata[524], rdata[523],
 rdata[522], rdata[521], rdata[520], rdata[519], rdata[518], rdata[517], rdata[516], rdata[515],
 rdata[514], rdata[513], rdata[512]};
if (n1)
_zymem[{n1, n2}] =
{rdata[1535], rdata[1534], rdata[1533], rdata[1532], rdata[1531],
 rdata[1530], rdata[1529], rdata[1528], rdata[1527], rdata[1526], rdata[1525], rdata[1524], rdata[1523],
 rdata[1522], rdata[1521], rdata[1520], rdata[1519], rdata[1518], rdata[1517], rdata[1516], rdata[1515],
 rdata[1514], rdata[1513], rdata[1512], rdata[1511], rdata[1510], rdata[1509], rdata[1508], rdata[1507],
 rdata[1506], rdata[1505], rdata[1504], rdata[1503], rdata[1502], rdata[1501], rdata[1500], rdata[1499],
 rdata[1498], rdata[1497], rdata[1496], rdata[1495], rdata[1494], rdata[1493], rdata[1492], rdata[1491],
 rdata[1490], rdata[1489], rdata[1488], rdata[1487], rdata[1486], rdata[1485], rdata[1484], rdata[1483],
 rdata[1482], rdata[1481], rdata[1480], rdata[1479], rdata[1478], rdata[1477], rdata[1476], rdata[1475],
 rdata[1474], rdata[1473], rdata[1472], rdata[1471], rdata[1470], rdata[1469], rdata[1468], rdata[1467],
 rdata[1466], rdata[1465], rdata[1464], rdata[1463], rdata[1462], rdata[1461], rdata[1460], rdata[1459],
 rdata[1458], rdata[1457], rdata[1456], rdata[1455], rdata[1454], rdata[1453], rdata[1452], rdata[1451],
 rdata[1450], rdata[1449], rdata[1448], rdata[1447], rdata[1446], rdata[1445], rdata[1444], rdata[1443],
 rdata[1442], rdata[1441], rdata[1440], rdata[1439], rdata[1438], rdata[1437], rdata[1436], rdata[1435],
 rdata[1434], rdata[1433], rdata[1432], rdata[1431], rdata[1430], rdata[1429], rdata[1428], rdata[1427],
 rdata[1426], rdata[1425], rdata[1424], rdata[1423], rdata[1422], rdata[1421], rdata[1420], rdata[1419],
 rdata[1418], rdata[1417], rdata[1416], rdata[1415], rdata[1414], rdata[1413], rdata[1412], rdata[1411],
 rdata[1410], rdata[1409], rdata[1408], rdata[1407], rdata[1406], rdata[1405], rdata[1404], rdata[1403],
 rdata[1402], rdata[1401], rdata[1400], rdata[1399], rdata[1398], rdata[1397], rdata[1396], rdata[1395],
 rdata[1394], rdata[1393], rdata[1392], rdata[1391], rdata[1390], rdata[1389], rdata[1388], rdata[1387],
 rdata[1386], rdata[1385], rdata[1384], rdata[1383], rdata[1382], rdata[1381], rdata[1380], rdata[1379],
 rdata[1378], rdata[1377], rdata[1376], rdata[1375], rdata[1374], rdata[1373], rdata[1372], rdata[1371],
 rdata[1370], rdata[1369], rdata[1368], rdata[1367], rdata[1366], rdata[1365], rdata[1364], rdata[1363],
 rdata[1362], rdata[1361], rdata[1360], rdata[1359], rdata[1358], rdata[1357], rdata[1356], rdata[1355],
 rdata[1354], rdata[1353], rdata[1352], rdata[1351], rdata[1350], rdata[1349], rdata[1348], rdata[1347],
 rdata[1346], rdata[1345], rdata[1344], rdata[1343], rdata[1342], rdata[1341], rdata[1340], rdata[1339],
 rdata[1338], rdata[1337], rdata[1336], rdata[1335], rdata[1334], rdata[1333], rdata[1332], rdata[1331],
 rdata[1330], rdata[1329], rdata[1328], rdata[1327], rdata[1326], rdata[1325], rdata[1324], rdata[1323],
 rdata[1322], rdata[1321], rdata[1320], rdata[1319], rdata[1318], rdata[1317], rdata[1316], rdata[1315],
 rdata[1314], rdata[1313], rdata[1312], rdata[1311], rdata[1310], rdata[1309], rdata[1308], rdata[1307],
 rdata[1306], rdata[1305], rdata[1304], rdata[1303], rdata[1302], rdata[1301], rdata[1300], rdata[1299],
 rdata[1298], rdata[1297], rdata[1296], rdata[1295], rdata[1294], rdata[1293], rdata[1292], rdata[1291],
 rdata[1290], rdata[1289], rdata[1288], rdata[1287], rdata[1286], rdata[1285], rdata[1284], rdata[1283],
 rdata[1282], rdata[1281], rdata[1280], rdata[1279], rdata[1278], rdata[1277], rdata[1276], rdata[1275],
 rdata[1274], rdata[1273], rdata[1272], rdata[1271], rdata[1270], rdata[1269], rdata[1268], rdata[1267],
 rdata[1266], rdata[1265], rdata[1264], rdata[1263], rdata[1262], rdata[1261], rdata[1260], rdata[1259],
 rdata[1258], rdata[1257], rdata[1256], rdata[1255], rdata[1254], rdata[1253], rdata[1252], rdata[1251],
 rdata[1250], rdata[1249], rdata[1248], rdata[1247], rdata[1246], rdata[1245], rdata[1244], rdata[1243],
 rdata[1242], rdata[1241], rdata[1240], rdata[1239], rdata[1238], rdata[1237], rdata[1236], rdata[1235],
 rdata[1234], rdata[1233], rdata[1232], rdata[1231], rdata[1230], rdata[1229], rdata[1228], rdata[1227],
 rdata[1226], rdata[1225], rdata[1224], rdata[1223], rdata[1222], rdata[1221], rdata[1220], rdata[1219],
 rdata[1218], rdata[1217], rdata[1216], rdata[1215], rdata[1214], rdata[1213], rdata[1212], rdata[1211],
 rdata[1210], rdata[1209], rdata[1208], rdata[1207], rdata[1206], rdata[1205], rdata[1204], rdata[1203],
 rdata[1202], rdata[1201], rdata[1200], rdata[1199], rdata[1198], rdata[1197], rdata[1196], rdata[1195],
 rdata[1194], rdata[1193], rdata[1192], rdata[1191], rdata[1190], rdata[1189], rdata[1188], rdata[1187],
 rdata[1186], rdata[1185], rdata[1184], rdata[1183], rdata[1182], rdata[1181], rdata[1180], rdata[1179],
 rdata[1178], rdata[1177], rdata[1176], rdata[1175], rdata[1174], rdata[1173], rdata[1172], rdata[1171],
 rdata[1170], rdata[1169], rdata[1168], rdata[1167], rdata[1166], rdata[1165], rdata[1164], rdata[1163],
 rdata[1162], rdata[1161], rdata[1160], rdata[1159], rdata[1158], rdata[1157], rdata[1156], rdata[1155],
 rdata[1154], rdata[1153], rdata[1152], rdata[1151], rdata[1150], rdata[1149], rdata[1148], rdata[1147],
 rdata[1146], rdata[1145], rdata[1144], rdata[1143], rdata[1142], rdata[1141], rdata[1140], rdata[1139],
 rdata[1138], rdata[1137], rdata[1136], rdata[1135], rdata[1134], rdata[1133], rdata[1132], rdata[1131],
 rdata[1130], rdata[1129], rdata[1128], rdata[1127], rdata[1126], rdata[1125], rdata[1124], rdata[1123],
 rdata[1122], rdata[1121], rdata[1120], rdata[1119], rdata[1118], rdata[1117], rdata[1116], rdata[1115],
 rdata[1114], rdata[1113], rdata[1112], rdata[1111], rdata[1110], rdata[1109], rdata[1108], rdata[1107],
 rdata[1106], rdata[1105], rdata[1104], rdata[1103], rdata[1102], rdata[1101], rdata[1100], rdata[1099],
 rdata[1098], rdata[1097], rdata[1096], rdata[1095], rdata[1094], rdata[1093], rdata[1092], rdata[1091],
 rdata[1090], rdata[1089], rdata[1088], rdata[1087], rdata[1086], rdata[1085], rdata[1084], rdata[1083],
 rdata[1082], rdata[1081], rdata[1080], rdata[1079], rdata[1078], rdata[1077], rdata[1076], rdata[1075],
 rdata[1074], rdata[1073], rdata[1072], rdata[1071], rdata[1070], rdata[1069], rdata[1068], rdata[1067],
 rdata[1066], rdata[1065], rdata[1064], rdata[1063], rdata[1062], rdata[1061], rdata[1060], rdata[1059],
 rdata[1058], rdata[1057], rdata[1056], rdata[1055], rdata[1054], rdata[1053], rdata[1052], rdata[1051],
 rdata[1050], rdata[1049], rdata[1048], rdata[1047], rdata[1046], rdata[1045], rdata[1044], rdata[1043],
 rdata[1042], rdata[1041], rdata[1040], rdata[1039], rdata[1038], rdata[1037], rdata[1036], rdata[1035],
 rdata[1034], rdata[1033], rdata[1032], rdata[1031], rdata[1030], rdata[1029], rdata[1028], rdata[1027],
 rdata[1026], rdata[1025], rdata[1024]};
if (n1)
_zymem[{n1, n1}] =
{rdata[2047], rdata[2046], rdata[2045], rdata[2044], rdata[2043],
 rdata[2042], rdata[2041], rdata[2040], rdata[2039], rdata[2038], rdata[2037], rdata[2036], rdata[2035],
 rdata[2034], rdata[2033], rdata[2032], rdata[2031], rdata[2030], rdata[2029], rdata[2028], rdata[2027],
 rdata[2026], rdata[2025], rdata[2024], rdata[2023], rdata[2022], rdata[2021], rdata[2020], rdata[2019],
 rdata[2018], rdata[2017], rdata[2016], rdata[2015], rdata[2014], rdata[2013], rdata[2012], rdata[2011],
 rdata[2010], rdata[2009], rdata[2008], rdata[2007], rdata[2006], rdata[2005], rdata[2004], rdata[2003],
 rdata[2002], rdata[2001], rdata[2000], rdata[1999], rdata[1998], rdata[1997], rdata[1996], rdata[1995],
 rdata[1994], rdata[1993], rdata[1992], rdata[1991], rdata[1990], rdata[1989], rdata[1988], rdata[1987],
 rdata[1986], rdata[1985], rdata[1984], rdata[1983], rdata[1982], rdata[1981], rdata[1980], rdata[1979],
 rdata[1978], rdata[1977], rdata[1976], rdata[1975], rdata[1974], rdata[1973], rdata[1972], rdata[1971],
 rdata[1970], rdata[1969], rdata[1968], rdata[1967], rdata[1966], rdata[1965], rdata[1964], rdata[1963],
 rdata[1962], rdata[1961], rdata[1960], rdata[1959], rdata[1958], rdata[1957], rdata[1956], rdata[1955],
 rdata[1954], rdata[1953], rdata[1952], rdata[1951], rdata[1950], rdata[1949], rdata[1948], rdata[1947],
 rdata[1946], rdata[1945], rdata[1944], rdata[1943], rdata[1942], rdata[1941], rdata[1940], rdata[1939],
 rdata[1938], rdata[1937], rdata[1936], rdata[1935], rdata[1934], rdata[1933], rdata[1932], rdata[1931],
 rdata[1930], rdata[1929], rdata[1928], rdata[1927], rdata[1926], rdata[1925], rdata[1924], rdata[1923],
 rdata[1922], rdata[1921], rdata[1920], rdata[1919], rdata[1918], rdata[1917], rdata[1916], rdata[1915],
 rdata[1914], rdata[1913], rdata[1912], rdata[1911], rdata[1910], rdata[1909], rdata[1908], rdata[1907],
 rdata[1906], rdata[1905], rdata[1904], rdata[1903], rdata[1902], rdata[1901], rdata[1900], rdata[1899],
 rdata[1898], rdata[1897], rdata[1896], rdata[1895], rdata[1894], rdata[1893], rdata[1892], rdata[1891],
 rdata[1890], rdata[1889], rdata[1888], rdata[1887], rdata[1886], rdata[1885], rdata[1884], rdata[1883],
 rdata[1882], rdata[1881], rdata[1880], rdata[1879], rdata[1878], rdata[1877], rdata[1876], rdata[1875],
 rdata[1874], rdata[1873], rdata[1872], rdata[1871], rdata[1870], rdata[1869], rdata[1868], rdata[1867],
 rdata[1866], rdata[1865], rdata[1864], rdata[1863], rdata[1862], rdata[1861], rdata[1860], rdata[1859],
 rdata[1858], rdata[1857], rdata[1856], rdata[1855], rdata[1854], rdata[1853], rdata[1852], rdata[1851],
 rdata[1850], rdata[1849], rdata[1848], rdata[1847], rdata[1846], rdata[1845], rdata[1844], rdata[1843],
 rdata[1842], rdata[1841], rdata[1840], rdata[1839], rdata[1838], rdata[1837], rdata[1836], rdata[1835],
 rdata[1834], rdata[1833], rdata[1832], rdata[1831], rdata[1830], rdata[1829], rdata[1828], rdata[1827],
 rdata[1826], rdata[1825], rdata[1824], rdata[1823], rdata[1822], rdata[1821], rdata[1820], rdata[1819],
 rdata[1818], rdata[1817], rdata[1816], rdata[1815], rdata[1814], rdata[1813], rdata[1812], rdata[1811],
 rdata[1810], rdata[1809], rdata[1808], rdata[1807], rdata[1806], rdata[1805], rdata[1804], rdata[1803],
 rdata[1802], rdata[1801], rdata[1800], rdata[1799], rdata[1798], rdata[1797], rdata[1796], rdata[1795],
 rdata[1794], rdata[1793], rdata[1792], rdata[1791], rdata[1790], rdata[1789], rdata[1788], rdata[1787],
 rdata[1786], rdata[1785], rdata[1784], rdata[1783], rdata[1782], rdata[1781], rdata[1780], rdata[1779],
 rdata[1778], rdata[1777], rdata[1776], rdata[1775], rdata[1774], rdata[1773], rdata[1772], rdata[1771],
 rdata[1770], rdata[1769], rdata[1768], rdata[1767], rdata[1766], rdata[1765], rdata[1764], rdata[1763],
 rdata[1762], rdata[1761], rdata[1760], rdata[1759], rdata[1758], rdata[1757], rdata[1756], rdata[1755],
 rdata[1754], rdata[1753], rdata[1752], rdata[1751], rdata[1750], rdata[1749], rdata[1748], rdata[1747],
 rdata[1746], rdata[1745], rdata[1744], rdata[1743], rdata[1742], rdata[1741], rdata[1740], rdata[1739],
 rdata[1738], rdata[1737], rdata[1736], rdata[1735], rdata[1734], rdata[1733], rdata[1732], rdata[1731],
 rdata[1730], rdata[1729], rdata[1728], rdata[1727], rdata[1726], rdata[1725], rdata[1724], rdata[1723],
 rdata[1722], rdata[1721], rdata[1720], rdata[1719], rdata[1718], rdata[1717], rdata[1716], rdata[1715],
 rdata[1714], rdata[1713], rdata[1712], rdata[1711], rdata[1710], rdata[1709], rdata[1708], rdata[1707],
 rdata[1706], rdata[1705], rdata[1704], rdata[1703], rdata[1702], rdata[1701], rdata[1700], rdata[1699],
 rdata[1698], rdata[1697], rdata[1696], rdata[1695], rdata[1694], rdata[1693], rdata[1692], rdata[1691],
 rdata[1690], rdata[1689], rdata[1688], rdata[1687], rdata[1686], rdata[1685], rdata[1684], rdata[1683],
 rdata[1682], rdata[1681], rdata[1680], rdata[1679], rdata[1678], rdata[1677], rdata[1676], rdata[1675],
 rdata[1674], rdata[1673], rdata[1672], rdata[1671], rdata[1670], rdata[1669], rdata[1668], rdata[1667],
 rdata[1666], rdata[1665], rdata[1664], rdata[1663], rdata[1662], rdata[1661], rdata[1660], rdata[1659],
 rdata[1658], rdata[1657], rdata[1656], rdata[1655], rdata[1654], rdata[1653], rdata[1652], rdata[1651],
 rdata[1650], rdata[1649], rdata[1648], rdata[1647], rdata[1646], rdata[1645], rdata[1644], rdata[1643],
 rdata[1642], rdata[1641], rdata[1640], rdata[1639], rdata[1638], rdata[1637], rdata[1636], rdata[1635],
 rdata[1634], rdata[1633], rdata[1632], rdata[1631], rdata[1630], rdata[1629], rdata[1628], rdata[1627],
 rdata[1626], rdata[1625], rdata[1624], rdata[1623], rdata[1622], rdata[1621], rdata[1620], rdata[1619],
 rdata[1618], rdata[1617], rdata[1616], rdata[1615], rdata[1614], rdata[1613], rdata[1612], rdata[1611],
 rdata[1610], rdata[1609], rdata[1608], rdata[1607], rdata[1606], rdata[1605], rdata[1604], rdata[1603],
 rdata[1602], rdata[1601], rdata[1600], rdata[1599], rdata[1598], rdata[1597], rdata[1596], rdata[1595],
 rdata[1594], rdata[1593], rdata[1592], rdata[1591], rdata[1590], rdata[1589], rdata[1588], rdata[1587],
 rdata[1586], rdata[1585], rdata[1584], rdata[1583], rdata[1582], rdata[1581], rdata[1580], rdata[1579],
 rdata[1578], rdata[1577], rdata[1576], rdata[1575], rdata[1574], rdata[1573], rdata[1572], rdata[1571],
 rdata[1570], rdata[1569], rdata[1568], rdata[1567], rdata[1566], rdata[1565], rdata[1564], rdata[1563],
 rdata[1562], rdata[1561], rdata[1560], rdata[1559], rdata[1558], rdata[1557], rdata[1556], rdata[1555],
 rdata[1554], rdata[1553], rdata[1552], rdata[1551], rdata[1550], rdata[1549], rdata[1548], rdata[1547],
 rdata[1546], rdata[1545], rdata[1544], rdata[1543], rdata[1542], rdata[1541], rdata[1540], rdata[1539],
 rdata[1538], rdata[1537], rdata[1536]};
end
`else

MPW4X512 _zymem ( .A1(n2), .A0(n2), .DI511(rdata[511]), .DI510(rdata[510]), .DI509(rdata[509]), .DI508(rdata[508]),
 .DI507(rdata[507]), .DI506(rdata[506]), .DI505(rdata[505]), .DI504(rdata[504]), .DI503(rdata[503]), .DI502(rdata[502]), .DI501(rdata[501]), .DI500(rdata[500]),
 .DI499(rdata[499]), .DI498(rdata[498]), .DI497(rdata[497]), .DI496(rdata[496]), .DI495(rdata[495]), .DI494(rdata[494]), .DI493(rdata[493]), .DI492(rdata[492]),
 .DI491(rdata[491]), .DI490(rdata[490]), .DI489(rdata[489]), .DI488(rdata[488]), .DI487(rdata[487]), .DI486(rdata[486]), .DI485(rdata[485]), .DI484(rdata[484]),
 .DI483(rdata[483]), .DI482(rdata[482]), .DI481(rdata[481]), .DI480(rdata[480]), .DI479(rdata[479]), .DI478(rdata[478]), .DI477(rdata[477]), .DI476(rdata[476]),
 .DI475(rdata[475]), .DI474(rdata[474]), .DI473(rdata[473]), .DI472(rdata[472]), .DI471(rdata[471]), .DI470(rdata[470]), .DI469(rdata[469]), .DI468(rdata[468]),
 .DI467(rdata[467]), .DI466(rdata[466]), .DI465(rdata[465]), .DI464(rdata[464]), .DI463(rdata[463]), .DI462(rdata[462]), .DI461(rdata[461]), .DI460(rdata[460]),
 .DI459(rdata[459]), .DI458(rdata[458]), .DI457(rdata[457]), .DI456(rdata[456]), .DI455(rdata[455]), .DI454(rdata[454]), .DI453(rdata[453]), .DI452(rdata[452]),
 .DI451(rdata[451]), .DI450(rdata[450]), .DI449(rdata[449]), .DI448(rdata[448]), .DI447(rdata[447]), .DI446(rdata[446]), .DI445(rdata[445]), .DI444(rdata[444]),
 .DI443(rdata[443]), .DI442(rdata[442]), .DI441(rdata[441]), .DI440(rdata[440]), .DI439(rdata[439]), .DI438(rdata[438]), .DI437(rdata[437]), .DI436(rdata[436]),
 .DI435(rdata[435]), .DI434(rdata[434]), .DI433(rdata[433]), .DI432(rdata[432]), .DI431(rdata[431]), .DI430(rdata[430]), .DI429(rdata[429]), .DI428(rdata[428]),
 .DI427(rdata[427]), .DI426(rdata[426]), .DI425(rdata[425]), .DI424(rdata[424]), .DI423(rdata[423]), .DI422(rdata[422]), .DI421(rdata[421]), .DI420(rdata[420]),
 .DI419(rdata[419]), .DI418(rdata[418]), .DI417(rdata[417]), .DI416(rdata[416]), .DI415(rdata[415]), .DI414(rdata[414]), .DI413(rdata[413]), .DI412(rdata[412]),
 .DI411(rdata[411]), .DI410(rdata[410]), .DI409(rdata[409]), .DI408(rdata[408]), .DI407(rdata[407]), .DI406(rdata[406]), .DI405(rdata[405]), .DI404(rdata[404]),
 .DI403(rdata[403]), .DI402(rdata[402]), .DI401(rdata[401]), .DI400(rdata[400]), .DI399(rdata[399]), .DI398(rdata[398]), .DI397(rdata[397]), .DI396(rdata[396]),
 .DI395(rdata[395]), .DI394(rdata[394]), .DI393(rdata[393]), .DI392(rdata[392]), .DI391(rdata[391]), .DI390(rdata[390]), .DI389(rdata[389]), .DI388(rdata[388]),
 .DI387(rdata[387]), .DI386(rdata[386]), .DI385(rdata[385]), .DI384(rdata[384]), .DI383(rdata[383]), .DI382(rdata[382]), .DI381(rdata[381]), .DI380(rdata[380]),
 .DI379(rdata[379]), .DI378(rdata[378]), .DI377(rdata[377]), .DI376(rdata[376]), .DI375(rdata[375]), .DI374(rdata[374]), .DI373(rdata[373]), .DI372(rdata[372]),
 .DI371(rdata[371]), .DI370(rdata[370]), .DI369(rdata[369]), .DI368(rdata[368]), .DI367(rdata[367]), .DI366(rdata[366]), .DI365(rdata[365]), .DI364(rdata[364]),
 .DI363(rdata[363]), .DI362(rdata[362]), .DI361(rdata[361]), .DI360(rdata[360]), .DI359(rdata[359]), .DI358(rdata[358]), .DI357(rdata[357]), .DI356(rdata[356]),
 .DI355(rdata[355]), .DI354(rdata[354]), .DI353(rdata[353]), .DI352(rdata[352]), .DI351(rdata[351]), .DI350(rdata[350]), .DI349(rdata[349]), .DI348(rdata[348]),
 .DI347(rdata[347]), .DI346(rdata[346]), .DI345(rdata[345]), .DI344(rdata[344]), .DI343(rdata[343]), .DI342(rdata[342]), .DI341(rdata[341]), .DI340(rdata[340]),
 .DI339(rdata[339]), .DI338(rdata[338]), .DI337(rdata[337]), .DI336(rdata[336]), .DI335(rdata[335]), .DI334(rdata[334]), .DI333(rdata[333]), .DI332(rdata[332]),
 .DI331(rdata[331]), .DI330(rdata[330]), .DI329(rdata[329]), .DI328(rdata[328]), .DI327(rdata[327]), .DI326(rdata[326]), .DI325(rdata[325]), .DI324(rdata[324]),
 .DI323(rdata[323]), .DI322(rdata[322]), .DI321(rdata[321]), .DI320(rdata[320]), .DI319(rdata[319]), .DI318(rdata[318]), .DI317(rdata[317]), .DI316(rdata[316]),
 .DI315(rdata[315]), .DI314(rdata[314]), .DI313(rdata[313]), .DI312(rdata[312]), .DI311(rdata[311]), .DI310(rdata[310]), .DI309(rdata[309]), .DI308(rdata[308]),
 .DI307(rdata[307]), .DI306(rdata[306]), .DI305(rdata[305]), .DI304(rdata[304]), .DI303(rdata[303]), .DI302(rdata[302]), .DI301(rdata[301]), .DI300(rdata[300]),
 .DI299(rdata[299]), .DI298(rdata[298]), .DI297(rdata[297]), .DI296(rdata[296]), .DI295(rdata[295]), .DI294(rdata[294]), .DI293(rdata[293]), .DI292(rdata[292]),
 .DI291(rdata[291]), .DI290(rdata[290]), .DI289(rdata[289]), .DI288(rdata[288]), .DI287(rdata[287]), .DI286(rdata[286]), .DI285(rdata[285]), .DI284(rdata[284]),
 .DI283(rdata[283]), .DI282(rdata[282]), .DI281(rdata[281]), .DI280(rdata[280]), .DI279(rdata[279]), .DI278(rdata[278]), .DI277(rdata[277]), .DI276(rdata[276]),
 .DI275(rdata[275]), .DI274(rdata[274]), .DI273(rdata[273]), .DI272(rdata[272]), .DI271(rdata[271]), .DI270(rdata[270]), .DI269(rdata[269]), .DI268(rdata[268]),
 .DI267(rdata[267]), .DI266(rdata[266]), .DI265(rdata[265]), .DI264(rdata[264]), .DI263(rdata[263]), .DI262(rdata[262]), .DI261(rdata[261]), .DI260(rdata[260]),
 .DI259(rdata[259]), .DI258(rdata[258]), .DI257(rdata[257]), .DI256(rdata[256]), .DI255(rdata[255]), .DI254(rdata[254]), .DI253(rdata[253]), .DI252(rdata[252]),
 .DI251(rdata[251]), .DI250(rdata[250]), .DI249(rdata[249]), .DI248(rdata[248]), .DI247(rdata[247]), .DI246(rdata[246]), .DI245(rdata[245]), .DI244(rdata[244]),
 .DI243(rdata[243]), .DI242(rdata[242]), .DI241(rdata[241]), .DI240(rdata[240]), .DI239(rdata[239]), .DI238(rdata[238]), .DI237(rdata[237]), .DI236(rdata[236]),
 .DI235(rdata[235]), .DI234(rdata[234]), .DI233(rdata[233]), .DI232(rdata[232]), .DI231(rdata[231]), .DI230(rdata[230]), .DI229(rdata[229]), .DI228(rdata[228]),
 .DI227(rdata[227]), .DI226(rdata[226]), .DI225(rdata[225]), .DI224(rdata[224]), .DI223(rdata[223]), .DI222(rdata[222]), .DI221(rdata[221]), .DI220(rdata[220]),
 .DI219(rdata[219]), .DI218(rdata[218]), .DI217(rdata[217]), .DI216(rdata[216]), .DI215(rdata[215]), .DI214(rdata[214]), .DI213(rdata[213]), .DI212(rdata[212]),
 .DI211(rdata[211]), .DI210(rdata[210]), .DI209(rdata[209]), .DI208(rdata[208]), .DI207(rdata[207]), .DI206(rdata[206]), .DI205(rdata[205]), .DI204(rdata[204]),
 .DI203(rdata[203]), .DI202(rdata[202]), .DI201(rdata[201]), .DI200(rdata[200]), .DI199(rdata[199]), .DI198(rdata[198]), .DI197(rdata[197]), .DI196(rdata[196]),
 .DI195(rdata[195]), .DI194(rdata[194]), .DI193(rdata[193]), .DI192(rdata[192]), .DI191(rdata[191]), .DI190(rdata[190]), .DI189(rdata[189]), .DI188(rdata[188]),
 .DI187(rdata[187]), .DI186(rdata[186]), .DI185(rdata[185]), .DI184(rdata[184]), .DI183(rdata[183]), .DI182(rdata[182]), .DI181(rdata[181]), .DI180(rdata[180]),
 .DI179(rdata[179]), .DI178(rdata[178]), .DI177(rdata[177]), .DI176(rdata[176]), .DI175(rdata[175]), .DI174(rdata[174]), .DI173(rdata[173]), .DI172(rdata[172]),
 .DI171(rdata[171]), .DI170(rdata[170]), .DI169(rdata[169]), .DI168(rdata[168]), .DI167(rdata[167]), .DI166(rdata[166]), .DI165(rdata[165]), .DI164(rdata[164]),
 .DI163(rdata[163]), .DI162(rdata[162]), .DI161(rdata[161]), .DI160(rdata[160]), .DI159(rdata[159]), .DI158(rdata[158]), .DI157(rdata[157]), .DI156(rdata[156]),
 .DI155(rdata[155]), .DI154(rdata[154]), .DI153(rdata[153]), .DI152(rdata[152]), .DI151(rdata[151]), .DI150(rdata[150]), .DI149(rdata[149]), .DI148(rdata[148]),
 .DI147(rdata[147]), .DI146(rdata[146]), .DI145(rdata[145]), .DI144(rdata[144]), .DI143(rdata[143]), .DI142(rdata[142]), .DI141(rdata[141]), .DI140(rdata[140]),
 .DI139(rdata[139]), .DI138(rdata[138]), .DI137(rdata[137]), .DI136(rdata[136]), .DI135(rdata[135]), .DI134(rdata[134]), .DI133(rdata[133]), .DI132(rdata[132]),
 .DI131(rdata[131]), .DI130(rdata[130]), .DI129(rdata[129]), .DI128(rdata[128]), .DI127(rdata[127]), .DI126(rdata[126]), .DI125(rdata[125]), .DI124(rdata[124]),
 .DI123(rdata[123]), .DI122(rdata[122]), .DI121(rdata[121]), .DI120(rdata[120]), .DI119(rdata[119]), .DI118(rdata[118]), .DI117(rdata[117]), .DI116(rdata[116]),
 .DI115(rdata[115]), .DI114(rdata[114]), .DI113(rdata[113]), .DI112(rdata[112]), .DI111(rdata[111]), .DI110(rdata[110]), .DI109(rdata[109]), .DI108(rdata[108]),
 .DI107(rdata[107]), .DI106(rdata[106]), .DI105(rdata[105]), .DI104(rdata[104]), .DI103(rdata[103]), .DI102(rdata[102]), .DI101(rdata[101]), .DI100(rdata[100]),
 .DI99(rdata[99]), .DI98(rdata[98]), .DI97(rdata[97]), .DI96(rdata[96]), .DI95(rdata[95]), .DI94(rdata[94]), .DI93(rdata[93]), .DI92(rdata[92]),
 .DI91(rdata[91]), .DI90(rdata[90]), .DI89(rdata[89]), .DI88(rdata[88]), .DI87(rdata[87]), .DI86(rdata[86]), .DI85(rdata[85]), .DI84(rdata[84]),
 .DI83(rdata[83]), .DI82(rdata[82]), .DI81(rdata[81]), .DI80(rdata[80]), .DI79(rdata[79]), .DI78(rdata[78]), .DI77(rdata[77]), .DI76(rdata[76]),
 .DI75(rdata[75]), .DI74(rdata[74]), .DI73(rdata[73]), .DI72(rdata[72]), .DI71(rdata[71]), .DI70(rdata[70]), .DI69(rdata[69]), .DI68(rdata[68]),
 .DI67(rdata[67]), .DI66(rdata[66]), .DI65(rdata[65]), .DI64(rdata[64]), .DI63(rdata[63]), .DI62(rdata[62]), .DI61(rdata[61]), .DI60(rdata[60]),
 .DI59(rdata[59]), .DI58(rdata[58]), .DI57(rdata[57]), .DI56(rdata[56]), .DI55(rdata[55]), .DI54(rdata[54]), .DI53(rdata[53]), .DI52(rdata[52]),
 .DI51(rdata[51]), .DI50(rdata[50]), .DI49(rdata[49]), .DI48(rdata[48]), .DI47(rdata[47]), .DI46(rdata[46]), .DI45(rdata[45]), .DI44(rdata[44]),
 .DI43(rdata[43]), .DI42(rdata[42]), .DI41(rdata[41]), .DI40(rdata[40]), .DI39(rdata[39]), .DI38(rdata[38]), .DI37(rdata[37]), .DI36(rdata[36]),
 .DI35(rdata[35]), .DI34(rdata[34]), .DI33(rdata[33]), .DI32(rdata[32]), .DI31(rdata[31]), .DI30(rdata[30]), .DI29(rdata[29]), .DI28(rdata[28]),
 .DI27(rdata[27]), .DI26(rdata[26]), .DI25(rdata[25]), .DI24(rdata[24]), .DI23(rdata[23]), .DI22(rdata[22]), .DI21(rdata[21]), .DI20(rdata[20]),
 .DI19(rdata[19]), .DI18(rdata[18]), .DI17(rdata[17]), .DI16(rdata[16]), .DI15(rdata[15]), .DI14(rdata[14]), .DI13(rdata[13]), .DI12(rdata[12]),
 .DI11(rdata[11]), .DI10(rdata[10]), .DI9(rdata[9]), .DI8(rdata[8]), .DI7(rdata[7]), .DI6(rdata[6]), .DI5(rdata[5]), .DI4(rdata[4]),
 .DI3(rdata[3]), .DI2(rdata[2]), .DI1(rdata[1]), .DI0(rdata[0]), .WE(n1), .SYNC_IN(n2), .SYNC_OUT(n4));
// pragma CVASTRPROP INSTANCE "_zymem" HDL_MEMORY_DECL "1 511 0 0 3"
MPW4X512 U2 ( .A1(n2), .A0(n1), .DI511(rdata[1023]), .DI510(rdata[1022]), .DI509(rdata[1021]), .DI508(rdata[1020]),
 .DI507(rdata[1019]), .DI506(rdata[1018]), .DI505(rdata[1017]), .DI504(rdata[1016]), .DI503(rdata[1015]), .DI502(rdata[1014]), .DI501(rdata[1013]), .DI500(rdata[1012]),
 .DI499(rdata[1011]), .DI498(rdata[1010]), .DI497(rdata[1009]), .DI496(rdata[1008]), .DI495(rdata[1007]), .DI494(rdata[1006]), .DI493(rdata[1005]), .DI492(rdata[1004]),
 .DI491(rdata[1003]), .DI490(rdata[1002]), .DI489(rdata[1001]), .DI488(rdata[1000]), .DI487(rdata[999]), .DI486(rdata[998]), .DI485(rdata[997]), .DI484(rdata[996]),
 .DI483(rdata[995]), .DI482(rdata[994]), .DI481(rdata[993]), .DI480(rdata[992]), .DI479(rdata[991]), .DI478(rdata[990]), .DI477(rdata[989]), .DI476(rdata[988]),
 .DI475(rdata[987]), .DI474(rdata[986]), .DI473(rdata[985]), .DI472(rdata[984]), .DI471(rdata[983]), .DI470(rdata[982]), .DI469(rdata[981]), .DI468(rdata[980]),
 .DI467(rdata[979]), .DI466(rdata[978]), .DI465(rdata[977]), .DI464(rdata[976]), .DI463(rdata[975]), .DI462(rdata[974]), .DI461(rdata[973]), .DI460(rdata[972]),
 .DI459(rdata[971]), .DI458(rdata[970]), .DI457(rdata[969]), .DI456(rdata[968]), .DI455(rdata[967]), .DI454(rdata[966]), .DI453(rdata[965]), .DI452(rdata[964]),
 .DI451(rdata[963]), .DI450(rdata[962]), .DI449(rdata[961]), .DI448(rdata[960]), .DI447(rdata[959]), .DI446(rdata[958]), .DI445(rdata[957]), .DI444(rdata[956]),
 .DI443(rdata[955]), .DI442(rdata[954]), .DI441(rdata[953]), .DI440(rdata[952]), .DI439(rdata[951]), .DI438(rdata[950]), .DI437(rdata[949]), .DI436(rdata[948]),
 .DI435(rdata[947]), .DI434(rdata[946]), .DI433(rdata[945]), .DI432(rdata[944]), .DI431(rdata[943]), .DI430(rdata[942]), .DI429(rdata[941]), .DI428(rdata[940]),
 .DI427(rdata[939]), .DI426(rdata[938]), .DI425(rdata[937]), .DI424(rdata[936]), .DI423(rdata[935]), .DI422(rdata[934]), .DI421(rdata[933]), .DI420(rdata[932]),
 .DI419(rdata[931]), .DI418(rdata[930]), .DI417(rdata[929]), .DI416(rdata[928]), .DI415(rdata[927]), .DI414(rdata[926]), .DI413(rdata[925]), .DI412(rdata[924]),
 .DI411(rdata[923]), .DI410(rdata[922]), .DI409(rdata[921]), .DI408(rdata[920]), .DI407(rdata[919]), .DI406(rdata[918]), .DI405(rdata[917]), .DI404(rdata[916]),
 .DI403(rdata[915]), .DI402(rdata[914]), .DI401(rdata[913]), .DI400(rdata[912]), .DI399(rdata[911]), .DI398(rdata[910]), .DI397(rdata[909]), .DI396(rdata[908]),
 .DI395(rdata[907]), .DI394(rdata[906]), .DI393(rdata[905]), .DI392(rdata[904]), .DI391(rdata[903]), .DI390(rdata[902]), .DI389(rdata[901]), .DI388(rdata[900]),
 .DI387(rdata[899]), .DI386(rdata[898]), .DI385(rdata[897]), .DI384(rdata[896]), .DI383(rdata[895]), .DI382(rdata[894]), .DI381(rdata[893]), .DI380(rdata[892]),
 .DI379(rdata[891]), .DI378(rdata[890]), .DI377(rdata[889]), .DI376(rdata[888]), .DI375(rdata[887]), .DI374(rdata[886]), .DI373(rdata[885]), .DI372(rdata[884]),
 .DI371(rdata[883]), .DI370(rdata[882]), .DI369(rdata[881]), .DI368(rdata[880]), .DI367(rdata[879]), .DI366(rdata[878]), .DI365(rdata[877]), .DI364(rdata[876]),
 .DI363(rdata[875]), .DI362(rdata[874]), .DI361(rdata[873]), .DI360(rdata[872]), .DI359(rdata[871]), .DI358(rdata[870]), .DI357(rdata[869]), .DI356(rdata[868]),
 .DI355(rdata[867]), .DI354(rdata[866]), .DI353(rdata[865]), .DI352(rdata[864]), .DI351(rdata[863]), .DI350(rdata[862]), .DI349(rdata[861]), .DI348(rdata[860]),
 .DI347(rdata[859]), .DI346(rdata[858]), .DI345(rdata[857]), .DI344(rdata[856]), .DI343(rdata[855]), .DI342(rdata[854]), .DI341(rdata[853]), .DI340(rdata[852]),
 .DI339(rdata[851]), .DI338(rdata[850]), .DI337(rdata[849]), .DI336(rdata[848]), .DI335(rdata[847]), .DI334(rdata[846]), .DI333(rdata[845]), .DI332(rdata[844]),
 .DI331(rdata[843]), .DI330(rdata[842]), .DI329(rdata[841]), .DI328(rdata[840]), .DI327(rdata[839]), .DI326(rdata[838]), .DI325(rdata[837]), .DI324(rdata[836]),
 .DI323(rdata[835]), .DI322(rdata[834]), .DI321(rdata[833]), .DI320(rdata[832]), .DI319(rdata[831]), .DI318(rdata[830]), .DI317(rdata[829]), .DI316(rdata[828]),
 .DI315(rdata[827]), .DI314(rdata[826]), .DI313(rdata[825]), .DI312(rdata[824]), .DI311(rdata[823]), .DI310(rdata[822]), .DI309(rdata[821]), .DI308(rdata[820]),
 .DI307(rdata[819]), .DI306(rdata[818]), .DI305(rdata[817]), .DI304(rdata[816]), .DI303(rdata[815]), .DI302(rdata[814]), .DI301(rdata[813]), .DI300(rdata[812]),
 .DI299(rdata[811]), .DI298(rdata[810]), .DI297(rdata[809]), .DI296(rdata[808]), .DI295(rdata[807]), .DI294(rdata[806]), .DI293(rdata[805]), .DI292(rdata[804]),
 .DI291(rdata[803]), .DI290(rdata[802]), .DI289(rdata[801]), .DI288(rdata[800]), .DI287(rdata[799]), .DI286(rdata[798]), .DI285(rdata[797]), .DI284(rdata[796]),
 .DI283(rdata[795]), .DI282(rdata[794]), .DI281(rdata[793]), .DI280(rdata[792]), .DI279(rdata[791]), .DI278(rdata[790]), .DI277(rdata[789]), .DI276(rdata[788]),
 .DI275(rdata[787]), .DI274(rdata[786]), .DI273(rdata[785]), .DI272(rdata[784]), .DI271(rdata[783]), .DI270(rdata[782]), .DI269(rdata[781]), .DI268(rdata[780]),
 .DI267(rdata[779]), .DI266(rdata[778]), .DI265(rdata[777]), .DI264(rdata[776]), .DI263(rdata[775]), .DI262(rdata[774]), .DI261(rdata[773]), .DI260(rdata[772]),
 .DI259(rdata[771]), .DI258(rdata[770]), .DI257(rdata[769]), .DI256(rdata[768]), .DI255(rdata[767]), .DI254(rdata[766]), .DI253(rdata[765]), .DI252(rdata[764]),
 .DI251(rdata[763]), .DI250(rdata[762]), .DI249(rdata[761]), .DI248(rdata[760]), .DI247(rdata[759]), .DI246(rdata[758]), .DI245(rdata[757]), .DI244(rdata[756]),
 .DI243(rdata[755]), .DI242(rdata[754]), .DI241(rdata[753]), .DI240(rdata[752]), .DI239(rdata[751]), .DI238(rdata[750]), .DI237(rdata[749]), .DI236(rdata[748]),
 .DI235(rdata[747]), .DI234(rdata[746]), .DI233(rdata[745]), .DI232(rdata[744]), .DI231(rdata[743]), .DI230(rdata[742]), .DI229(rdata[741]), .DI228(rdata[740]),
 .DI227(rdata[739]), .DI226(rdata[738]), .DI225(rdata[737]), .DI224(rdata[736]), .DI223(rdata[735]), .DI222(rdata[734]), .DI221(rdata[733]), .DI220(rdata[732]),
 .DI219(rdata[731]), .DI218(rdata[730]), .DI217(rdata[729]), .DI216(rdata[728]), .DI215(rdata[727]), .DI214(rdata[726]), .DI213(rdata[725]), .DI212(rdata[724]),
 .DI211(rdata[723]), .DI210(rdata[722]), .DI209(rdata[721]), .DI208(rdata[720]), .DI207(rdata[719]), .DI206(rdata[718]), .DI205(rdata[717]), .DI204(rdata[716]),
 .DI203(rdata[715]), .DI202(rdata[714]), .DI201(rdata[713]), .DI200(rdata[712]), .DI199(rdata[711]), .DI198(rdata[710]), .DI197(rdata[709]), .DI196(rdata[708]),
 .DI195(rdata[707]), .DI194(rdata[706]), .DI193(rdata[705]), .DI192(rdata[704]), .DI191(rdata[703]), .DI190(rdata[702]), .DI189(rdata[701]), .DI188(rdata[700]),
 .DI187(rdata[699]), .DI186(rdata[698]), .DI185(rdata[697]), .DI184(rdata[696]), .DI183(rdata[695]), .DI182(rdata[694]), .DI181(rdata[693]), .DI180(rdata[692]),
 .DI179(rdata[691]), .DI178(rdata[690]), .DI177(rdata[689]), .DI176(rdata[688]), .DI175(rdata[687]), .DI174(rdata[686]), .DI173(rdata[685]), .DI172(rdata[684]),
 .DI171(rdata[683]), .DI170(rdata[682]), .DI169(rdata[681]), .DI168(rdata[680]), .DI167(rdata[679]), .DI166(rdata[678]), .DI165(rdata[677]), .DI164(rdata[676]),
 .DI163(rdata[675]), .DI162(rdata[674]), .DI161(rdata[673]), .DI160(rdata[672]), .DI159(rdata[671]), .DI158(rdata[670]), .DI157(rdata[669]), .DI156(rdata[668]),
 .DI155(rdata[667]), .DI154(rdata[666]), .DI153(rdata[665]), .DI152(rdata[664]), .DI151(rdata[663]), .DI150(rdata[662]), .DI149(rdata[661]), .DI148(rdata[660]),
 .DI147(rdata[659]), .DI146(rdata[658]), .DI145(rdata[657]), .DI144(rdata[656]), .DI143(rdata[655]), .DI142(rdata[654]), .DI141(rdata[653]), .DI140(rdata[652]),
 .DI139(rdata[651]), .DI138(rdata[650]), .DI137(rdata[649]), .DI136(rdata[648]), .DI135(rdata[647]), .DI134(rdata[646]), .DI133(rdata[645]), .DI132(rdata[644]),
 .DI131(rdata[643]), .DI130(rdata[642]), .DI129(rdata[641]), .DI128(rdata[640]), .DI127(rdata[639]), .DI126(rdata[638]), .DI125(rdata[637]), .DI124(rdata[636]),
 .DI123(rdata[635]), .DI122(rdata[634]), .DI121(rdata[633]), .DI120(rdata[632]), .DI119(rdata[631]), .DI118(rdata[630]), .DI117(rdata[629]), .DI116(rdata[628]),
 .DI115(rdata[627]), .DI114(rdata[626]), .DI113(rdata[625]), .DI112(rdata[624]), .DI111(rdata[623]), .DI110(rdata[622]), .DI109(rdata[621]), .DI108(rdata[620]),
 .DI107(rdata[619]), .DI106(rdata[618]), .DI105(rdata[617]), .DI104(rdata[616]), .DI103(rdata[615]), .DI102(rdata[614]), .DI101(rdata[613]), .DI100(rdata[612]),
 .DI99(rdata[611]), .DI98(rdata[610]), .DI97(rdata[609]), .DI96(rdata[608]), .DI95(rdata[607]), .DI94(rdata[606]), .DI93(rdata[605]), .DI92(rdata[604]),
 .DI91(rdata[603]), .DI90(rdata[602]), .DI89(rdata[601]), .DI88(rdata[600]), .DI87(rdata[599]), .DI86(rdata[598]), .DI85(rdata[597]), .DI84(rdata[596]),
 .DI83(rdata[595]), .DI82(rdata[594]), .DI81(rdata[593]), .DI80(rdata[592]), .DI79(rdata[591]), .DI78(rdata[590]), .DI77(rdata[589]), .DI76(rdata[588]),
 .DI75(rdata[587]), .DI74(rdata[586]), .DI73(rdata[585]), .DI72(rdata[584]), .DI71(rdata[583]), .DI70(rdata[582]), .DI69(rdata[581]), .DI68(rdata[580]),
 .DI67(rdata[579]), .DI66(rdata[578]), .DI65(rdata[577]), .DI64(rdata[576]), .DI63(rdata[575]), .DI62(rdata[574]), .DI61(rdata[573]), .DI60(rdata[572]),
 .DI59(rdata[571]), .DI58(rdata[570]), .DI57(rdata[569]), .DI56(rdata[568]), .DI55(rdata[567]), .DI54(rdata[566]), .DI53(rdata[565]), .DI52(rdata[564]),
 .DI51(rdata[563]), .DI50(rdata[562]), .DI49(rdata[561]), .DI48(rdata[560]), .DI47(rdata[559]), .DI46(rdata[558]), .DI45(rdata[557]), .DI44(rdata[556]),
 .DI43(rdata[555]), .DI42(rdata[554]), .DI41(rdata[553]), .DI40(rdata[552]), .DI39(rdata[551]), .DI38(rdata[550]), .DI37(rdata[549]), .DI36(rdata[548]),
 .DI35(rdata[547]), .DI34(rdata[546]), .DI33(rdata[545]), .DI32(rdata[544]), .DI31(rdata[543]), .DI30(rdata[542]), .DI29(rdata[541]), .DI28(rdata[540]),
 .DI27(rdata[539]), .DI26(rdata[538]), .DI25(rdata[537]), .DI24(rdata[536]), .DI23(rdata[535]), .DI22(rdata[534]), .DI21(rdata[533]), .DI20(rdata[532]),
 .DI19(rdata[531]), .DI18(rdata[530]), .DI17(rdata[529]), .DI16(rdata[528]), .DI15(rdata[527]), .DI14(rdata[526]), .DI13(rdata[525]), .DI12(rdata[524]),
 .DI11(rdata[523]), .DI10(rdata[522]), .DI9(rdata[521]), .DI8(rdata[520]), .DI7(rdata[519]), .DI6(rdata[518]), .DI5(rdata[517]), .DI4(rdata[516]),
 .DI3(rdata[515]), .DI2(rdata[514]), .DI1(rdata[513]), .DI0(rdata[512]), .WE(n1), .SYNC_IN(n4), .SYNC_OUT(n5));
MPW4X512 U3 ( .A1(n1), .A0(n2), .DI511(rdata[1535]), .DI510(rdata[1534]), .DI509(rdata[1533]), .DI508(rdata[1532]),
 .DI507(rdata[1531]), .DI506(rdata[1530]), .DI505(rdata[1529]), .DI504(rdata[1528]), .DI503(rdata[1527]), .DI502(rdata[1526]), .DI501(rdata[1525]), .DI500(rdata[1524]),
 .DI499(rdata[1523]), .DI498(rdata[1522]), .DI497(rdata[1521]), .DI496(rdata[1520]), .DI495(rdata[1519]), .DI494(rdata[1518]), .DI493(rdata[1517]), .DI492(rdata[1516]),
 .DI491(rdata[1515]), .DI490(rdata[1514]), .DI489(rdata[1513]), .DI488(rdata[1512]), .DI487(rdata[1511]), .DI486(rdata[1510]), .DI485(rdata[1509]), .DI484(rdata[1508]),
 .DI483(rdata[1507]), .DI482(rdata[1506]), .DI481(rdata[1505]), .DI480(rdata[1504]), .DI479(rdata[1503]), .DI478(rdata[1502]), .DI477(rdata[1501]), .DI476(rdata[1500]),
 .DI475(rdata[1499]), .DI474(rdata[1498]), .DI473(rdata[1497]), .DI472(rdata[1496]), .DI471(rdata[1495]), .DI470(rdata[1494]), .DI469(rdata[1493]), .DI468(rdata[1492]),
 .DI467(rdata[1491]), .DI466(rdata[1490]), .DI465(rdata[1489]), .DI464(rdata[1488]), .DI463(rdata[1487]), .DI462(rdata[1486]), .DI461(rdata[1485]), .DI460(rdata[1484]),
 .DI459(rdata[1483]), .DI458(rdata[1482]), .DI457(rdata[1481]), .DI456(rdata[1480]), .DI455(rdata[1479]), .DI454(rdata[1478]), .DI453(rdata[1477]), .DI452(rdata[1476]),
 .DI451(rdata[1475]), .DI450(rdata[1474]), .DI449(rdata[1473]), .DI448(rdata[1472]), .DI447(rdata[1471]), .DI446(rdata[1470]), .DI445(rdata[1469]), .DI444(rdata[1468]),
 .DI443(rdata[1467]), .DI442(rdata[1466]), .DI441(rdata[1465]), .DI440(rdata[1464]), .DI439(rdata[1463]), .DI438(rdata[1462]), .DI437(rdata[1461]), .DI436(rdata[1460]),
 .DI435(rdata[1459]), .DI434(rdata[1458]), .DI433(rdata[1457]), .DI432(rdata[1456]), .DI431(rdata[1455]), .DI430(rdata[1454]), .DI429(rdata[1453]), .DI428(rdata[1452]),
 .DI427(rdata[1451]), .DI426(rdata[1450]), .DI425(rdata[1449]), .DI424(rdata[1448]), .DI423(rdata[1447]), .DI422(rdata[1446]), .DI421(rdata[1445]), .DI420(rdata[1444]),
 .DI419(rdata[1443]), .DI418(rdata[1442]), .DI417(rdata[1441]), .DI416(rdata[1440]), .DI415(rdata[1439]), .DI414(rdata[1438]), .DI413(rdata[1437]), .DI412(rdata[1436]),
 .DI411(rdata[1435]), .DI410(rdata[1434]), .DI409(rdata[1433]), .DI408(rdata[1432]), .DI407(rdata[1431]), .DI406(rdata[1430]), .DI405(rdata[1429]), .DI404(rdata[1428]),
 .DI403(rdata[1427]), .DI402(rdata[1426]), .DI401(rdata[1425]), .DI400(rdata[1424]), .DI399(rdata[1423]), .DI398(rdata[1422]), .DI397(rdata[1421]), .DI396(rdata[1420]),
 .DI395(rdata[1419]), .DI394(rdata[1418]), .DI393(rdata[1417]), .DI392(rdata[1416]), .DI391(rdata[1415]), .DI390(rdata[1414]), .DI389(rdata[1413]), .DI388(rdata[1412]),
 .DI387(rdata[1411]), .DI386(rdata[1410]), .DI385(rdata[1409]), .DI384(rdata[1408]), .DI383(rdata[1407]), .DI382(rdata[1406]), .DI381(rdata[1405]), .DI380(rdata[1404]),
 .DI379(rdata[1403]), .DI378(rdata[1402]), .DI377(rdata[1401]), .DI376(rdata[1400]), .DI375(rdata[1399]), .DI374(rdata[1398]), .DI373(rdata[1397]), .DI372(rdata[1396]),
 .DI371(rdata[1395]), .DI370(rdata[1394]), .DI369(rdata[1393]), .DI368(rdata[1392]), .DI367(rdata[1391]), .DI366(rdata[1390]), .DI365(rdata[1389]), .DI364(rdata[1388]),
 .DI363(rdata[1387]), .DI362(rdata[1386]), .DI361(rdata[1385]), .DI360(rdata[1384]), .DI359(rdata[1383]), .DI358(rdata[1382]), .DI357(rdata[1381]), .DI356(rdata[1380]),
 .DI355(rdata[1379]), .DI354(rdata[1378]), .DI353(rdata[1377]), .DI352(rdata[1376]), .DI351(rdata[1375]), .DI350(rdata[1374]), .DI349(rdata[1373]), .DI348(rdata[1372]),
 .DI347(rdata[1371]), .DI346(rdata[1370]), .DI345(rdata[1369]), .DI344(rdata[1368]), .DI343(rdata[1367]), .DI342(rdata[1366]), .DI341(rdata[1365]), .DI340(rdata[1364]),
 .DI339(rdata[1363]), .DI338(rdata[1362]), .DI337(rdata[1361]), .DI336(rdata[1360]), .DI335(rdata[1359]), .DI334(rdata[1358]), .DI333(rdata[1357]), .DI332(rdata[1356]),
 .DI331(rdata[1355]), .DI330(rdata[1354]), .DI329(rdata[1353]), .DI328(rdata[1352]), .DI327(rdata[1351]), .DI326(rdata[1350]), .DI325(rdata[1349]), .DI324(rdata[1348]),
 .DI323(rdata[1347]), .DI322(rdata[1346]), .DI321(rdata[1345]), .DI320(rdata[1344]), .DI319(rdata[1343]), .DI318(rdata[1342]), .DI317(rdata[1341]), .DI316(rdata[1340]),
 .DI315(rdata[1339]), .DI314(rdata[1338]), .DI313(rdata[1337]), .DI312(rdata[1336]), .DI311(rdata[1335]), .DI310(rdata[1334]), .DI309(rdata[1333]), .DI308(rdata[1332]),
 .DI307(rdata[1331]), .DI306(rdata[1330]), .DI305(rdata[1329]), .DI304(rdata[1328]), .DI303(rdata[1327]), .DI302(rdata[1326]), .DI301(rdata[1325]), .DI300(rdata[1324]),
 .DI299(rdata[1323]), .DI298(rdata[1322]), .DI297(rdata[1321]), .DI296(rdata[1320]), .DI295(rdata[1319]), .DI294(rdata[1318]), .DI293(rdata[1317]), .DI292(rdata[1316]),
 .DI291(rdata[1315]), .DI290(rdata[1314]), .DI289(rdata[1313]), .DI288(rdata[1312]), .DI287(rdata[1311]), .DI286(rdata[1310]), .DI285(rdata[1309]), .DI284(rdata[1308]),
 .DI283(rdata[1307]), .DI282(rdata[1306]), .DI281(rdata[1305]), .DI280(rdata[1304]), .DI279(rdata[1303]), .DI278(rdata[1302]), .DI277(rdata[1301]), .DI276(rdata[1300]),
 .DI275(rdata[1299]), .DI274(rdata[1298]), .DI273(rdata[1297]), .DI272(rdata[1296]), .DI271(rdata[1295]), .DI270(rdata[1294]), .DI269(rdata[1293]), .DI268(rdata[1292]),
 .DI267(rdata[1291]), .DI266(rdata[1290]), .DI265(rdata[1289]), .DI264(rdata[1288]), .DI263(rdata[1287]), .DI262(rdata[1286]), .DI261(rdata[1285]), .DI260(rdata[1284]),
 .DI259(rdata[1283]), .DI258(rdata[1282]), .DI257(rdata[1281]), .DI256(rdata[1280]), .DI255(rdata[1279]), .DI254(rdata[1278]), .DI253(rdata[1277]), .DI252(rdata[1276]),
 .DI251(rdata[1275]), .DI250(rdata[1274]), .DI249(rdata[1273]), .DI248(rdata[1272]), .DI247(rdata[1271]), .DI246(rdata[1270]), .DI245(rdata[1269]), .DI244(rdata[1268]),
 .DI243(rdata[1267]), .DI242(rdata[1266]), .DI241(rdata[1265]), .DI240(rdata[1264]), .DI239(rdata[1263]), .DI238(rdata[1262]), .DI237(rdata[1261]), .DI236(rdata[1260]),
 .DI235(rdata[1259]), .DI234(rdata[1258]), .DI233(rdata[1257]), .DI232(rdata[1256]), .DI231(rdata[1255]), .DI230(rdata[1254]), .DI229(rdata[1253]), .DI228(rdata[1252]),
 .DI227(rdata[1251]), .DI226(rdata[1250]), .DI225(rdata[1249]), .DI224(rdata[1248]), .DI223(rdata[1247]), .DI222(rdata[1246]), .DI221(rdata[1245]), .DI220(rdata[1244]),
 .DI219(rdata[1243]), .DI218(rdata[1242]), .DI217(rdata[1241]), .DI216(rdata[1240]), .DI215(rdata[1239]), .DI214(rdata[1238]), .DI213(rdata[1237]), .DI212(rdata[1236]),
 .DI211(rdata[1235]), .DI210(rdata[1234]), .DI209(rdata[1233]), .DI208(rdata[1232]), .DI207(rdata[1231]), .DI206(rdata[1230]), .DI205(rdata[1229]), .DI204(rdata[1228]),
 .DI203(rdata[1227]), .DI202(rdata[1226]), .DI201(rdata[1225]), .DI200(rdata[1224]), .DI199(rdata[1223]), .DI198(rdata[1222]), .DI197(rdata[1221]), .DI196(rdata[1220]),
 .DI195(rdata[1219]), .DI194(rdata[1218]), .DI193(rdata[1217]), .DI192(rdata[1216]), .DI191(rdata[1215]), .DI190(rdata[1214]), .DI189(rdata[1213]), .DI188(rdata[1212]),
 .DI187(rdata[1211]), .DI186(rdata[1210]), .DI185(rdata[1209]), .DI184(rdata[1208]), .DI183(rdata[1207]), .DI182(rdata[1206]), .DI181(rdata[1205]), .DI180(rdata[1204]),
 .DI179(rdata[1203]), .DI178(rdata[1202]), .DI177(rdata[1201]), .DI176(rdata[1200]), .DI175(rdata[1199]), .DI174(rdata[1198]), .DI173(rdata[1197]), .DI172(rdata[1196]),
 .DI171(rdata[1195]), .DI170(rdata[1194]), .DI169(rdata[1193]), .DI168(rdata[1192]), .DI167(rdata[1191]), .DI166(rdata[1190]), .DI165(rdata[1189]), .DI164(rdata[1188]),
 .DI163(rdata[1187]), .DI162(rdata[1186]), .DI161(rdata[1185]), .DI160(rdata[1184]), .DI159(rdata[1183]), .DI158(rdata[1182]), .DI157(rdata[1181]), .DI156(rdata[1180]),
 .DI155(rdata[1179]), .DI154(rdata[1178]), .DI153(rdata[1177]), .DI152(rdata[1176]), .DI151(rdata[1175]), .DI150(rdata[1174]), .DI149(rdata[1173]), .DI148(rdata[1172]),
 .DI147(rdata[1171]), .DI146(rdata[1170]), .DI145(rdata[1169]), .DI144(rdata[1168]), .DI143(rdata[1167]), .DI142(rdata[1166]), .DI141(rdata[1165]), .DI140(rdata[1164]),
 .DI139(rdata[1163]), .DI138(rdata[1162]), .DI137(rdata[1161]), .DI136(rdata[1160]), .DI135(rdata[1159]), .DI134(rdata[1158]), .DI133(rdata[1157]), .DI132(rdata[1156]),
 .DI131(rdata[1155]), .DI130(rdata[1154]), .DI129(rdata[1153]), .DI128(rdata[1152]), .DI127(rdata[1151]), .DI126(rdata[1150]), .DI125(rdata[1149]), .DI124(rdata[1148]),
 .DI123(rdata[1147]), .DI122(rdata[1146]), .DI121(rdata[1145]), .DI120(rdata[1144]), .DI119(rdata[1143]), .DI118(rdata[1142]), .DI117(rdata[1141]), .DI116(rdata[1140]),
 .DI115(rdata[1139]), .DI114(rdata[1138]), .DI113(rdata[1137]), .DI112(rdata[1136]), .DI111(rdata[1135]), .DI110(rdata[1134]), .DI109(rdata[1133]), .DI108(rdata[1132]),
 .DI107(rdata[1131]), .DI106(rdata[1130]), .DI105(rdata[1129]), .DI104(rdata[1128]), .DI103(rdata[1127]), .DI102(rdata[1126]), .DI101(rdata[1125]), .DI100(rdata[1124]),
 .DI99(rdata[1123]), .DI98(rdata[1122]), .DI97(rdata[1121]), .DI96(rdata[1120]), .DI95(rdata[1119]), .DI94(rdata[1118]), .DI93(rdata[1117]), .DI92(rdata[1116]),
 .DI91(rdata[1115]), .DI90(rdata[1114]), .DI89(rdata[1113]), .DI88(rdata[1112]), .DI87(rdata[1111]), .DI86(rdata[1110]), .DI85(rdata[1109]), .DI84(rdata[1108]),
 .DI83(rdata[1107]), .DI82(rdata[1106]), .DI81(rdata[1105]), .DI80(rdata[1104]), .DI79(rdata[1103]), .DI78(rdata[1102]), .DI77(rdata[1101]), .DI76(rdata[1100]),
 .DI75(rdata[1099]), .DI74(rdata[1098]), .DI73(rdata[1097]), .DI72(rdata[1096]), .DI71(rdata[1095]), .DI70(rdata[1094]), .DI69(rdata[1093]), .DI68(rdata[1092]),
 .DI67(rdata[1091]), .DI66(rdata[1090]), .DI65(rdata[1089]), .DI64(rdata[1088]), .DI63(rdata[1087]), .DI62(rdata[1086]), .DI61(rdata[1085]), .DI60(rdata[1084]),
 .DI59(rdata[1083]), .DI58(rdata[1082]), .DI57(rdata[1081]), .DI56(rdata[1080]), .DI55(rdata[1079]), .DI54(rdata[1078]), .DI53(rdata[1077]), .DI52(rdata[1076]),
 .DI51(rdata[1075]), .DI50(rdata[1074]), .DI49(rdata[1073]), .DI48(rdata[1072]), .DI47(rdata[1071]), .DI46(rdata[1070]), .DI45(rdata[1069]), .DI44(rdata[1068]),
 .DI43(rdata[1067]), .DI42(rdata[1066]), .DI41(rdata[1065]), .DI40(rdata[1064]), .DI39(rdata[1063]), .DI38(rdata[1062]), .DI37(rdata[1061]), .DI36(rdata[1060]),
 .DI35(rdata[1059]), .DI34(rdata[1058]), .DI33(rdata[1057]), .DI32(rdata[1056]), .DI31(rdata[1055]), .DI30(rdata[1054]), .DI29(rdata[1053]), .DI28(rdata[1052]),
 .DI27(rdata[1051]), .DI26(rdata[1050]), .DI25(rdata[1049]), .DI24(rdata[1048]), .DI23(rdata[1047]), .DI22(rdata[1046]), .DI21(rdata[1045]), .DI20(rdata[1044]),
 .DI19(rdata[1043]), .DI18(rdata[1042]), .DI17(rdata[1041]), .DI16(rdata[1040]), .DI15(rdata[1039]), .DI14(rdata[1038]), .DI13(rdata[1037]), .DI12(rdata[1036]),
 .DI11(rdata[1035]), .DI10(rdata[1034]), .DI9(rdata[1033]), .DI8(rdata[1032]), .DI7(rdata[1031]), .DI6(rdata[1030]), .DI5(rdata[1029]), .DI4(rdata[1028]),
 .DI3(rdata[1027]), .DI2(rdata[1026]), .DI1(rdata[1025]), .DI0(rdata[1024]), .WE(n1), .SYNC_IN(n5), .SYNC_OUT(n6));
MPW4X512 U4 ( .A1(n1), .A0(n1), .DI511(rdata[2047]), .DI510(rdata[2046]), .DI509(rdata[2045]), .DI508(rdata[2044]),
 .DI507(rdata[2043]), .DI506(rdata[2042]), .DI505(rdata[2041]), .DI504(rdata[2040]), .DI503(rdata[2039]), .DI502(rdata[2038]), .DI501(rdata[2037]), .DI500(rdata[2036]),
 .DI499(rdata[2035]), .DI498(rdata[2034]), .DI497(rdata[2033]), .DI496(rdata[2032]), .DI495(rdata[2031]), .DI494(rdata[2030]), .DI493(rdata[2029]), .DI492(rdata[2028]),
 .DI491(rdata[2027]), .DI490(rdata[2026]), .DI489(rdata[2025]), .DI488(rdata[2024]), .DI487(rdata[2023]), .DI486(rdata[2022]), .DI485(rdata[2021]), .DI484(rdata[2020]),
 .DI483(rdata[2019]), .DI482(rdata[2018]), .DI481(rdata[2017]), .DI480(rdata[2016]), .DI479(rdata[2015]), .DI478(rdata[2014]), .DI477(rdata[2013]), .DI476(rdata[2012]),
 .DI475(rdata[2011]), .DI474(rdata[2010]), .DI473(rdata[2009]), .DI472(rdata[2008]), .DI471(rdata[2007]), .DI470(rdata[2006]), .DI469(rdata[2005]), .DI468(rdata[2004]),
 .DI467(rdata[2003]), .DI466(rdata[2002]), .DI465(rdata[2001]), .DI464(rdata[2000]), .DI463(rdata[1999]), .DI462(rdata[1998]), .DI461(rdata[1997]), .DI460(rdata[1996]),
 .DI459(rdata[1995]), .DI458(rdata[1994]), .DI457(rdata[1993]), .DI456(rdata[1992]), .DI455(rdata[1991]), .DI454(rdata[1990]), .DI453(rdata[1989]), .DI452(rdata[1988]),
 .DI451(rdata[1987]), .DI450(rdata[1986]), .DI449(rdata[1985]), .DI448(rdata[1984]), .DI447(rdata[1983]), .DI446(rdata[1982]), .DI445(rdata[1981]), .DI444(rdata[1980]),
 .DI443(rdata[1979]), .DI442(rdata[1978]), .DI441(rdata[1977]), .DI440(rdata[1976]), .DI439(rdata[1975]), .DI438(rdata[1974]), .DI437(rdata[1973]), .DI436(rdata[1972]),
 .DI435(rdata[1971]), .DI434(rdata[1970]), .DI433(rdata[1969]), .DI432(rdata[1968]), .DI431(rdata[1967]), .DI430(rdata[1966]), .DI429(rdata[1965]), .DI428(rdata[1964]),
 .DI427(rdata[1963]), .DI426(rdata[1962]), .DI425(rdata[1961]), .DI424(rdata[1960]), .DI423(rdata[1959]), .DI422(rdata[1958]), .DI421(rdata[1957]), .DI420(rdata[1956]),
 .DI419(rdata[1955]), .DI418(rdata[1954]), .DI417(rdata[1953]), .DI416(rdata[1952]), .DI415(rdata[1951]), .DI414(rdata[1950]), .DI413(rdata[1949]), .DI412(rdata[1948]),
 .DI411(rdata[1947]), .DI410(rdata[1946]), .DI409(rdata[1945]), .DI408(rdata[1944]), .DI407(rdata[1943]), .DI406(rdata[1942]), .DI405(rdata[1941]), .DI404(rdata[1940]),
 .DI403(rdata[1939]), .DI402(rdata[1938]), .DI401(rdata[1937]), .DI400(rdata[1936]), .DI399(rdata[1935]), .DI398(rdata[1934]), .DI397(rdata[1933]), .DI396(rdata[1932]),
 .DI395(rdata[1931]), .DI394(rdata[1930]), .DI393(rdata[1929]), .DI392(rdata[1928]), .DI391(rdata[1927]), .DI390(rdata[1926]), .DI389(rdata[1925]), .DI388(rdata[1924]),
 .DI387(rdata[1923]), .DI386(rdata[1922]), .DI385(rdata[1921]), .DI384(rdata[1920]), .DI383(rdata[1919]), .DI382(rdata[1918]), .DI381(rdata[1917]), .DI380(rdata[1916]),
 .DI379(rdata[1915]), .DI378(rdata[1914]), .DI377(rdata[1913]), .DI376(rdata[1912]), .DI375(rdata[1911]), .DI374(rdata[1910]), .DI373(rdata[1909]), .DI372(rdata[1908]),
 .DI371(rdata[1907]), .DI370(rdata[1906]), .DI369(rdata[1905]), .DI368(rdata[1904]), .DI367(rdata[1903]), .DI366(rdata[1902]), .DI365(rdata[1901]), .DI364(rdata[1900]),
 .DI363(rdata[1899]), .DI362(rdata[1898]), .DI361(rdata[1897]), .DI360(rdata[1896]), .DI359(rdata[1895]), .DI358(rdata[1894]), .DI357(rdata[1893]), .DI356(rdata[1892]),
 .DI355(rdata[1891]), .DI354(rdata[1890]), .DI353(rdata[1889]), .DI352(rdata[1888]), .DI351(rdata[1887]), .DI350(rdata[1886]), .DI349(rdata[1885]), .DI348(rdata[1884]),
 .DI347(rdata[1883]), .DI346(rdata[1882]), .DI345(rdata[1881]), .DI344(rdata[1880]), .DI343(rdata[1879]), .DI342(rdata[1878]), .DI341(rdata[1877]), .DI340(rdata[1876]),
 .DI339(rdata[1875]), .DI338(rdata[1874]), .DI337(rdata[1873]), .DI336(rdata[1872]), .DI335(rdata[1871]), .DI334(rdata[1870]), .DI333(rdata[1869]), .DI332(rdata[1868]),
 .DI331(rdata[1867]), .DI330(rdata[1866]), .DI329(rdata[1865]), .DI328(rdata[1864]), .DI327(rdata[1863]), .DI326(rdata[1862]), .DI325(rdata[1861]), .DI324(rdata[1860]),
 .DI323(rdata[1859]), .DI322(rdata[1858]), .DI321(rdata[1857]), .DI320(rdata[1856]), .DI319(rdata[1855]), .DI318(rdata[1854]), .DI317(rdata[1853]), .DI316(rdata[1852]),
 .DI315(rdata[1851]), .DI314(rdata[1850]), .DI313(rdata[1849]), .DI312(rdata[1848]), .DI311(rdata[1847]), .DI310(rdata[1846]), .DI309(rdata[1845]), .DI308(rdata[1844]),
 .DI307(rdata[1843]), .DI306(rdata[1842]), .DI305(rdata[1841]), .DI304(rdata[1840]), .DI303(rdata[1839]), .DI302(rdata[1838]), .DI301(rdata[1837]), .DI300(rdata[1836]),
 .DI299(rdata[1835]), .DI298(rdata[1834]), .DI297(rdata[1833]), .DI296(rdata[1832]), .DI295(rdata[1831]), .DI294(rdata[1830]), .DI293(rdata[1829]), .DI292(rdata[1828]),
 .DI291(rdata[1827]), .DI290(rdata[1826]), .DI289(rdata[1825]), .DI288(rdata[1824]), .DI287(rdata[1823]), .DI286(rdata[1822]), .DI285(rdata[1821]), .DI284(rdata[1820]),
 .DI283(rdata[1819]), .DI282(rdata[1818]), .DI281(rdata[1817]), .DI280(rdata[1816]), .DI279(rdata[1815]), .DI278(rdata[1814]), .DI277(rdata[1813]), .DI276(rdata[1812]),
 .DI275(rdata[1811]), .DI274(rdata[1810]), .DI273(rdata[1809]), .DI272(rdata[1808]), .DI271(rdata[1807]), .DI270(rdata[1806]), .DI269(rdata[1805]), .DI268(rdata[1804]),
 .DI267(rdata[1803]), .DI266(rdata[1802]), .DI265(rdata[1801]), .DI264(rdata[1800]), .DI263(rdata[1799]), .DI262(rdata[1798]), .DI261(rdata[1797]), .DI260(rdata[1796]),
 .DI259(rdata[1795]), .DI258(rdata[1794]), .DI257(rdata[1793]), .DI256(rdata[1792]), .DI255(rdata[1791]), .DI254(rdata[1790]), .DI253(rdata[1789]), .DI252(rdata[1788]),
 .DI251(rdata[1787]), .DI250(rdata[1786]), .DI249(rdata[1785]), .DI248(rdata[1784]), .DI247(rdata[1783]), .DI246(rdata[1782]), .DI245(rdata[1781]), .DI244(rdata[1780]),
 .DI243(rdata[1779]), .DI242(rdata[1778]), .DI241(rdata[1777]), .DI240(rdata[1776]), .DI239(rdata[1775]), .DI238(rdata[1774]), .DI237(rdata[1773]), .DI236(rdata[1772]),
 .DI235(rdata[1771]), .DI234(rdata[1770]), .DI233(rdata[1769]), .DI232(rdata[1768]), .DI231(rdata[1767]), .DI230(rdata[1766]), .DI229(rdata[1765]), .DI228(rdata[1764]),
 .DI227(rdata[1763]), .DI226(rdata[1762]), .DI225(rdata[1761]), .DI224(rdata[1760]), .DI223(rdata[1759]), .DI222(rdata[1758]), .DI221(rdata[1757]), .DI220(rdata[1756]),
 .DI219(rdata[1755]), .DI218(rdata[1754]), .DI217(rdata[1753]), .DI216(rdata[1752]), .DI215(rdata[1751]), .DI214(rdata[1750]), .DI213(rdata[1749]), .DI212(rdata[1748]),
 .DI211(rdata[1747]), .DI210(rdata[1746]), .DI209(rdata[1745]), .DI208(rdata[1744]), .DI207(rdata[1743]), .DI206(rdata[1742]), .DI205(rdata[1741]), .DI204(rdata[1740]),
 .DI203(rdata[1739]), .DI202(rdata[1738]), .DI201(rdata[1737]), .DI200(rdata[1736]), .DI199(rdata[1735]), .DI198(rdata[1734]), .DI197(rdata[1733]), .DI196(rdata[1732]),
 .DI195(rdata[1731]), .DI194(rdata[1730]), .DI193(rdata[1729]), .DI192(rdata[1728]), .DI191(rdata[1727]), .DI190(rdata[1726]), .DI189(rdata[1725]), .DI188(rdata[1724]),
 .DI187(rdata[1723]), .DI186(rdata[1722]), .DI185(rdata[1721]), .DI184(rdata[1720]), .DI183(rdata[1719]), .DI182(rdata[1718]), .DI181(rdata[1717]), .DI180(rdata[1716]),
 .DI179(rdata[1715]), .DI178(rdata[1714]), .DI177(rdata[1713]), .DI176(rdata[1712]), .DI175(rdata[1711]), .DI174(rdata[1710]), .DI173(rdata[1709]), .DI172(rdata[1708]),
 .DI171(rdata[1707]), .DI170(rdata[1706]), .DI169(rdata[1705]), .DI168(rdata[1704]), .DI167(rdata[1703]), .DI166(rdata[1702]), .DI165(rdata[1701]), .DI164(rdata[1700]),
 .DI163(rdata[1699]), .DI162(rdata[1698]), .DI161(rdata[1697]), .DI160(rdata[1696]), .DI159(rdata[1695]), .DI158(rdata[1694]), .DI157(rdata[1693]), .DI156(rdata[1692]),
 .DI155(rdata[1691]), .DI154(rdata[1690]), .DI153(rdata[1689]), .DI152(rdata[1688]), .DI151(rdata[1687]), .DI150(rdata[1686]), .DI149(rdata[1685]), .DI148(rdata[1684]),
 .DI147(rdata[1683]), .DI146(rdata[1682]), .DI145(rdata[1681]), .DI144(rdata[1680]), .DI143(rdata[1679]), .DI142(rdata[1678]), .DI141(rdata[1677]), .DI140(rdata[1676]),
 .DI139(rdata[1675]), .DI138(rdata[1674]), .DI137(rdata[1673]), .DI136(rdata[1672]), .DI135(rdata[1671]), .DI134(rdata[1670]), .DI133(rdata[1669]), .DI132(rdata[1668]),
 .DI131(rdata[1667]), .DI130(rdata[1666]), .DI129(rdata[1665]), .DI128(rdata[1664]), .DI127(rdata[1663]), .DI126(rdata[1662]), .DI125(rdata[1661]), .DI124(rdata[1660]),
 .DI123(rdata[1659]), .DI122(rdata[1658]), .DI121(rdata[1657]), .DI120(rdata[1656]), .DI119(rdata[1655]), .DI118(rdata[1654]), .DI117(rdata[1653]), .DI116(rdata[1652]),
 .DI115(rdata[1651]), .DI114(rdata[1650]), .DI113(rdata[1649]), .DI112(rdata[1648]), .DI111(rdata[1647]), .DI110(rdata[1646]), .DI109(rdata[1645]), .DI108(rdata[1644]),
 .DI107(rdata[1643]), .DI106(rdata[1642]), .DI105(rdata[1641]), .DI104(rdata[1640]), .DI103(rdata[1639]), .DI102(rdata[1638]), .DI101(rdata[1637]), .DI100(rdata[1636]),
 .DI99(rdata[1635]), .DI98(rdata[1634]), .DI97(rdata[1633]), .DI96(rdata[1632]), .DI95(rdata[1631]), .DI94(rdata[1630]), .DI93(rdata[1629]), .DI92(rdata[1628]),
 .DI91(rdata[1627]), .DI90(rdata[1626]), .DI89(rdata[1625]), .DI88(rdata[1624]), .DI87(rdata[1623]), .DI86(rdata[1622]), .DI85(rdata[1621]), .DI84(rdata[1620]),
 .DI83(rdata[1619]), .DI82(rdata[1618]), .DI81(rdata[1617]), .DI80(rdata[1616]), .DI79(rdata[1615]), .DI78(rdata[1614]), .DI77(rdata[1613]), .DI76(rdata[1612]),
 .DI75(rdata[1611]), .DI74(rdata[1610]), .DI73(rdata[1609]), .DI72(rdata[1608]), .DI71(rdata[1607]), .DI70(rdata[1606]), .DI69(rdata[1605]), .DI68(rdata[1604]),
 .DI67(rdata[1603]), .DI66(rdata[1602]), .DI65(rdata[1601]), .DI64(rdata[1600]), .DI63(rdata[1599]), .DI62(rdata[1598]), .DI61(rdata[1597]), .DI60(rdata[1596]),
 .DI59(rdata[1595]), .DI58(rdata[1594]), .DI57(rdata[1593]), .DI56(rdata[1592]), .DI55(rdata[1591]), .DI54(rdata[1590]), .DI53(rdata[1589]), .DI52(rdata[1588]),
 .DI51(rdata[1587]), .DI50(rdata[1586]), .DI49(rdata[1585]), .DI48(rdata[1584]), .DI47(rdata[1583]), .DI46(rdata[1582]), .DI45(rdata[1581]), .DI44(rdata[1580]),
 .DI43(rdata[1579]), .DI42(rdata[1578]), .DI41(rdata[1577]), .DI40(rdata[1576]), .DI39(rdata[1575]), .DI38(rdata[1574]), .DI37(rdata[1573]), .DI36(rdata[1572]),
 .DI35(rdata[1571]), .DI34(rdata[1570]), .DI33(rdata[1569]), .DI32(rdata[1568]), .DI31(rdata[1567]), .DI30(rdata[1566]), .DI29(rdata[1565]), .DI28(rdata[1564]),
 .DI27(rdata[1563]), .DI26(rdata[1562]), .DI25(rdata[1561]), .DI24(rdata[1560]), .DI23(rdata[1559]), .DI22(rdata[1558]), .DI21(rdata[1557]), .DI20(rdata[1556]),
 .DI19(rdata[1555]), .DI18(rdata[1554]), .DI17(rdata[1553]), .DI16(rdata[1552]), .DI15(rdata[1551]), .DI14(rdata[1550]), .DI13(rdata[1549]), .DI12(rdata[1548]),
 .DI11(rdata[1547]), .DI10(rdata[1546]), .DI9(rdata[1545]), .DI8(rdata[1544]), .DI7(rdata[1543]), .DI6(rdata[1542]), .DI5(rdata[1541]), .DI4(rdata[1540]),
 .DI3(rdata[1539]), .DI2(rdata[1538]), .DI1(rdata[1537]), .DI0(rdata[1536]), .WE(n1), .SYNC_IN(n6), .SYNC_OUT( ));
`endif
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "_zymem 1 511 0 0 3"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "1"
// pragma CVASTRPROP MODULE HDLICE CVAIUSNAMES_FORGEN_LABEL "genblk1"
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE "ixc_context_read"
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE_LIB "IXCOM_TEMP_LIBRARY"
// pragma CVASTRPROP MODULE HDLICE PROP_IXCOM_MOD TRUE
endmodule
`ifdef CBV
`else
`ifdef MPW4X512_MPR4X512
`else
module MPW4X512( A1, A0, DI511, DI510, DI509, DI508, DI507,
 DI506, DI505, DI504, DI503, DI502, DI501, DI500, DI499,
 DI498, DI497, DI496, DI495, DI494, DI493, DI492, DI491,
 DI490, DI489, DI488, DI487, DI486, DI485, DI484, DI483,
 DI482, DI481, DI480, DI479, DI478, DI477, DI476, DI475,
 DI474, DI473, DI472, DI471, DI470, DI469, DI468, DI467,
 DI466, DI465, DI464, DI463, DI462, DI461, DI460, DI459,
 DI458, DI457, DI456, DI455, DI454, DI453, DI452, DI451,
 DI450, DI449, DI448, DI447, DI446, DI445, DI444, DI443,
 DI442, DI441, DI440, DI439, DI438, DI437, DI436, DI435,
 DI434, DI433, DI432, DI431, DI430, DI429, DI428, DI427,
 DI426, DI425, DI424, DI423, DI422, DI421, DI420, DI419,
 DI418, DI417, DI416, DI415, DI414, DI413, DI412, DI411,
 DI410, DI409, DI408, DI407, DI406, DI405, DI404, DI403,
 DI402, DI401, DI400, DI399, DI398, DI397, DI396, DI395,
 DI394, DI393, DI392, DI391, DI390, DI389, DI388, DI387,
 DI386, DI385, DI384, DI383, DI382, DI381, DI380, DI379,
 DI378, DI377, DI376, DI375, DI374, DI373, DI372, DI371,
 DI370, DI369, DI368, DI367, DI366, DI365, DI364, DI363,
 DI362, DI361, DI360, DI359, DI358, DI357, DI356, DI355,
 DI354, DI353, DI352, DI351, DI350, DI349, DI348, DI347,
 DI346, DI345, DI344, DI343, DI342, DI341, DI340, DI339,
 DI338, DI337, DI336, DI335, DI334, DI333, DI332, DI331,
 DI330, DI329, DI328, DI327, DI326, DI325, DI324, DI323,
 DI322, DI321, DI320, DI319, DI318, DI317, DI316, DI315,
 DI314, DI313, DI312, DI311, DI310, DI309, DI308, DI307,
 DI306, DI305, DI304, DI303, DI302, DI301, DI300, DI299,
 DI298, DI297, DI296, DI295, DI294, DI293, DI292, DI291,
 DI290, DI289, DI288, DI287, DI286, DI285, DI284, DI283,
 DI282, DI281, DI280, DI279, DI278, DI277, DI276, DI275,
 DI274, DI273, DI272, DI271, DI270, DI269, DI268, DI267,
 DI266, DI265, DI264, DI263, DI262, DI261, DI260, DI259,
 DI258, DI257, DI256, DI255, DI254, DI253, DI252, DI251,
 DI250, DI249, DI248, DI247, DI246, DI245, DI244, DI243,
 DI242, DI241, DI240, DI239, DI238, DI237, DI236, DI235,
 DI234, DI233, DI232, DI231, DI230, DI229, DI228, DI227,
 DI226, DI225, DI224, DI223, DI222, DI221, DI220, DI219,
 DI218, DI217, DI216, DI215, DI214, DI213, DI212, DI211,
 DI210, DI209, DI208, DI207, DI206, DI205, DI204, DI203,
 DI202, DI201, DI200, DI199, DI198, DI197, DI196, DI195,
 DI194, DI193, DI192, DI191, DI190, DI189, DI188, DI187,
 DI186, DI185, DI184, DI183, DI182, DI181, DI180, DI179,
 DI178, DI177, DI176, DI175, DI174, DI173, DI172, DI171,
 DI170, DI169, DI168, DI167, DI166, DI165, DI164, DI163,
 DI162, DI161, DI160, DI159, DI158, DI157, DI156, DI155,
 DI154, DI153, DI152, DI151, DI150, DI149, DI148, DI147,
 DI146, DI145, DI144, DI143, DI142, DI141, DI140, DI139,
 DI138, DI137, DI136, DI135, DI134, DI133, DI132, DI131,
 DI130, DI129, DI128, DI127, DI126, DI125, DI124, DI123,
 DI122, DI121, DI120, DI119, DI118, DI117, DI116, DI115,
 DI114, DI113, DI112, DI111, DI110, DI109, DI108, DI107,
 DI106, DI105, DI104, DI103, DI102, DI101, DI100, DI99,
 DI98, DI97, DI96, DI95, DI94, DI93, DI92, DI91,
 DI90, DI89, DI88, DI87, DI86, DI85, DI84, DI83,
 DI82, DI81, DI80, DI79, DI78, DI77, DI76, DI75,
 DI74, DI73, DI72, DI71, DI70, DI69, DI68, DI67,
 DI66, DI65, DI64, DI63, DI62, DI61, DI60, DI59,
 DI58, DI57, DI56, DI55, DI54, DI53, DI52, DI51,
 DI50, DI49, DI48, DI47, DI46, DI45, DI44, DI43,
 DI42, DI41, DI40, DI39, DI38, DI37, DI36, DI35,
 DI34, DI33, DI32, DI31, DI30, DI29, DI28, DI27,
 DI26, DI25, DI24, DI23, DI22, DI21, DI20, DI19,
 DI18, DI17, DI16, DI15, DI14, DI13, DI12, DI11,
 DI10, DI9, DI8, DI7, DI6, DI5, DI4, DI3,
 DI2, DI1, DI0, WE, SYNC_IN, SYNC_OUT);
input  A1, A0, DI511, DI510, DI509, DI508, DI507, DI506,
 DI505, DI504, DI503, DI502, DI501, DI500, DI499, DI498, DI497, DI496,
 DI495, DI494, DI493, DI492, DI491, DI490, DI489, DI488, DI487, DI486,
 DI485, DI484, DI483, DI482, DI481, DI480, DI479, DI478, DI477, DI476,
 DI475, DI474, DI473, DI472, DI471, DI470, DI469, DI468, DI467, DI466,
 DI465, DI464, DI463, DI462, DI461, DI460, DI459, DI458, DI457, DI456,
 DI455, DI454, DI453, DI452, DI451, DI450, DI449, DI448, DI447, DI446,
 DI445, DI444, DI443, DI442, DI441, DI440, DI439, DI438, DI437, DI436,
 DI435, DI434, DI433, DI432, DI431, DI430, DI429, DI428, DI427, DI426,
 DI425, DI424, DI423, DI422, DI421, DI420, DI419, DI418, DI417, DI416,
 DI415, DI414, DI413, DI412, DI411, DI410, DI409, DI408, DI407, DI406,
 DI405, DI404, DI403, DI402, DI401, DI400, DI399, DI398, DI397, DI396,
 DI395, DI394, DI393, DI392, DI391, DI390, DI389, DI388, DI387, DI386,
 DI385, DI384, DI383, DI382, DI381, DI380, DI379, DI378, DI377, DI376,
 DI375, DI374, DI373, DI372, DI371, DI370, DI369, DI368, DI367, DI366,
 DI365, DI364, DI363, DI362, DI361, DI360, DI359, DI358, DI357, DI356,
 DI355, DI354, DI353, DI352, DI351, DI350, DI349, DI348, DI347, DI346,
 DI345, DI344, DI343, DI342, DI341, DI340, DI339, DI338, DI337, DI336,
 DI335, DI334, DI333, DI332, DI331, DI330, DI329, DI328, DI327, DI326,
 DI325, DI324, DI323, DI322, DI321, DI320, DI319, DI318, DI317, DI316,
 DI315, DI314, DI313, DI312, DI311, DI310, DI309, DI308, DI307, DI306,
 DI305, DI304, DI303, DI302, DI301, DI300, DI299, DI298, DI297, DI296,
 DI295, DI294, DI293, DI292, DI291, DI290, DI289, DI288, DI287, DI286,
 DI285, DI284, DI283, DI282, DI281, DI280, DI279, DI278, DI277, DI276,
 DI275, DI274, DI273, DI272, DI271, DI270, DI269, DI268, DI267, DI266,
 DI265, DI264, DI263, DI262, DI261, DI260, DI259, DI258, DI257, DI256,
 DI255, DI254, DI253, DI252, DI251, DI250, DI249, DI248, DI247, DI246,
 DI245, DI244, DI243, DI242, DI241, DI240, DI239, DI238, DI237, DI236,
 DI235, DI234, DI233, DI232, DI231, DI230, DI229, DI228, DI227, DI226,
 DI225, DI224, DI223, DI222, DI221, DI220, DI219, DI218, DI217, DI216,
 DI215, DI214, DI213, DI212, DI211, DI210, DI209, DI208, DI207, DI206,
 DI205, DI204, DI203, DI202, DI201, DI200, DI199, DI198, DI197, DI196,
 DI195, DI194, DI193, DI192, DI191, DI190, DI189, DI188, DI187, DI186,
 DI185, DI184, DI183, DI182, DI181, DI180, DI179, DI178, DI177, DI176,
 DI175, DI174, DI173, DI172, DI171, DI170, DI169, DI168, DI167, DI166,
 DI165, DI164, DI163, DI162, DI161, DI160, DI159, DI158, DI157, DI156,
 DI155, DI154, DI153, DI152, DI151, DI150, DI149, DI148, DI147, DI146,
 DI145, DI144, DI143, DI142, DI141, DI140, DI139, DI138, DI137, DI136,
 DI135, DI134, DI133, DI132, DI131, DI130, DI129, DI128, DI127, DI126,
 DI125, DI124, DI123, DI122, DI121, DI120, DI119, DI118, DI117, DI116,
 DI115, DI114, DI113, DI112, DI111, DI110, DI109, DI108, DI107, DI106,
 DI105, DI104, DI103, DI102, DI101, DI100, DI99, DI98, DI97, DI96,
 DI95, DI94, DI93, DI92, DI91, DI90, DI89, DI88, DI87, DI86,
 DI85, DI84, DI83, DI82, DI81, DI80, DI79, DI78, DI77, DI76,
 DI75, DI74, DI73, DI72, DI71, DI70, DI69, DI68, DI67, DI66,
 DI65, DI64, DI63, DI62, DI61, DI60, DI59, DI58, DI57, DI56,
 DI55, DI54, DI53, DI52, DI51, DI50, DI49, DI48, DI47, DI46,
 DI45, DI44, DI43, DI42, DI41, DI40, DI39, DI38, DI37, DI36,
 DI35, DI34, DI33, DI32, DI31, DI30, DI29, DI28, DI27, DI26,
 DI25, DI24, DI23, DI22, DI21, DI20, DI19, DI18, DI17, DI16,
 DI15, DI14, DI13, DI12, DI11, DI10, DI9, DI8, DI7, DI6,
 DI5, DI4, DI3, DI2, DI1, DI0, WE, SYNC_IN;
output  SYNC_OUT;
endmodule
`ifdef _MPR4X512_
`else
module MPR4X512( A1, A0, SYNC_IN, DO511, DO510, DO509, DO508,
 DO507, DO506, DO505, DO504, DO503, DO502, DO501, DO500,
 DO499, DO498, DO497, DO496, DO495, DO494, DO493, DO492,
 DO491, DO490, DO489, DO488, DO487, DO486, DO485, DO484,
 DO483, DO482, DO481, DO480, DO479, DO478, DO477, DO476,
 DO475, DO474, DO473, DO472, DO471, DO470, DO469, DO468,
 DO467, DO466, DO465, DO464, DO463, DO462, DO461, DO460,
 DO459, DO458, DO457, DO456, DO455, DO454, DO453, DO452,
 DO451, DO450, DO449, DO448, DO447, DO446, DO445, DO444,
 DO443, DO442, DO441, DO440, DO439, DO438, DO437, DO436,
 DO435, DO434, DO433, DO432, DO431, DO430, DO429, DO428,
 DO427, DO426, DO425, DO424, DO423, DO422, DO421, DO420,
 DO419, DO418, DO417, DO416, DO415, DO414, DO413, DO412,
 DO411, DO410, DO409, DO408, DO407, DO406, DO405, DO404,
 DO403, DO402, DO401, DO400, DO399, DO398, DO397, DO396,
 DO395, DO394, DO393, DO392, DO391, DO390, DO389, DO388,
 DO387, DO386, DO385, DO384, DO383, DO382, DO381, DO380,
 DO379, DO378, DO377, DO376, DO375, DO374, DO373, DO372,
 DO371, DO370, DO369, DO368, DO367, DO366, DO365, DO364,
 DO363, DO362, DO361, DO360, DO359, DO358, DO357, DO356,
 DO355, DO354, DO353, DO352, DO351, DO350, DO349, DO348,
 DO347, DO346, DO345, DO344, DO343, DO342, DO341, DO340,
 DO339, DO338, DO337, DO336, DO335, DO334, DO333, DO332,
 DO331, DO330, DO329, DO328, DO327, DO326, DO325, DO324,
 DO323, DO322, DO321, DO320, DO319, DO318, DO317, DO316,
 DO315, DO314, DO313, DO312, DO311, DO310, DO309, DO308,
 DO307, DO306, DO305, DO304, DO303, DO302, DO301, DO300,
 DO299, DO298, DO297, DO296, DO295, DO294, DO293, DO292,
 DO291, DO290, DO289, DO288, DO287, DO286, DO285, DO284,
 DO283, DO282, DO281, DO280, DO279, DO278, DO277, DO276,
 DO275, DO274, DO273, DO272, DO271, DO270, DO269, DO268,
 DO267, DO266, DO265, DO264, DO263, DO262, DO261, DO260,
 DO259, DO258, DO257, DO256, DO255, DO254, DO253, DO252,
 DO251, DO250, DO249, DO248, DO247, DO246, DO245, DO244,
 DO243, DO242, DO241, DO240, DO239, DO238, DO237, DO236,
 DO235, DO234, DO233, DO232, DO231, DO230, DO229, DO228,
 DO227, DO226, DO225, DO224, DO223, DO222, DO221, DO220,
 DO219, DO218, DO217, DO216, DO215, DO214, DO213, DO212,
 DO211, DO210, DO209, DO208, DO207, DO206, DO205, DO204,
 DO203, DO202, DO201, DO200, DO199, DO198, DO197, DO196,
 DO195, DO194, DO193, DO192, DO191, DO190, DO189, DO188,
 DO187, DO186, DO185, DO184, DO183, DO182, DO181, DO180,
 DO179, DO178, DO177, DO176, DO175, DO174, DO173, DO172,
 DO171, DO170, DO169, DO168, DO167, DO166, DO165, DO164,
 DO163, DO162, DO161, DO160, DO159, DO158, DO157, DO156,
 DO155, DO154, DO153, DO152, DO151, DO150, DO149, DO148,
 DO147, DO146, DO145, DO144, DO143, DO142, DO141, DO140,
 DO139, DO138, DO137, DO136, DO135, DO134, DO133, DO132,
 DO131, DO130, DO129, DO128, DO127, DO126, DO125, DO124,
 DO123, DO122, DO121, DO120, DO119, DO118, DO117, DO116,
 DO115, DO114, DO113, DO112, DO111, DO110, DO109, DO108,
 DO107, DO106, DO105, DO104, DO103, DO102, DO101, DO100,
 DO99, DO98, DO97, DO96, DO95, DO94, DO93, DO92,
 DO91, DO90, DO89, DO88, DO87, DO86, DO85, DO84,
 DO83, DO82, DO81, DO80, DO79, DO78, DO77, DO76,
 DO75, DO74, DO73, DO72, DO71, DO70, DO69, DO68,
 DO67, DO66, DO65, DO64, DO63, DO62, DO61, DO60,
 DO59, DO58, DO57, DO56, DO55, DO54, DO53, DO52,
 DO51, DO50, DO49, DO48, DO47, DO46, DO45, DO44,
 DO43, DO42, DO41, DO40, DO39, DO38, DO37, DO36,
 DO35, DO34, DO33, DO32, DO31, DO30, DO29, DO28,
 DO27, DO26, DO25, DO24, DO23, DO22, DO21, DO20,
 DO19, DO18, DO17, DO16, DO15, DO14, DO13, DO12,
 DO11, DO10, DO9, DO8, DO7, DO6, DO5, DO4,
 DO3, DO2, DO1, DO0, SYNC_OUT);
input  A1, A0, SYNC_IN;
output  DO511, DO510, DO509, DO508, DO507, DO506, DO505, DO504,
 DO503, DO502, DO501, DO500, DO499, DO498, DO497, DO496, DO495, DO494,
 DO493, DO492, DO491, DO490, DO489, DO488, DO487, DO486, DO485, DO484,
 DO483, DO482, DO481, DO480, DO479, DO478, DO477, DO476, DO475, DO474,
 DO473, DO472, DO471, DO470, DO469, DO468, DO467, DO466, DO465, DO464,
 DO463, DO462, DO461, DO460, DO459, DO458, DO457, DO456, DO455, DO454,
 DO453, DO452, DO451, DO450, DO449, DO448, DO447, DO446, DO445, DO444,
 DO443, DO442, DO441, DO440, DO439, DO438, DO437, DO436, DO435, DO434,
 DO433, DO432, DO431, DO430, DO429, DO428, DO427, DO426, DO425, DO424,
 DO423, DO422, DO421, DO420, DO419, DO418, DO417, DO416, DO415, DO414,
 DO413, DO412, DO411, DO410, DO409, DO408, DO407, DO406, DO405, DO404,
 DO403, DO402, DO401, DO400, DO399, DO398, DO397, DO396, DO395, DO394,
 DO393, DO392, DO391, DO390, DO389, DO388, DO387, DO386, DO385, DO384,
 DO383, DO382, DO381, DO380, DO379, DO378, DO377, DO376, DO375, DO374,
 DO373, DO372, DO371, DO370, DO369, DO368, DO367, DO366, DO365, DO364,
 DO363, DO362, DO361, DO360, DO359, DO358, DO357, DO356, DO355, DO354,
 DO353, DO352, DO351, DO350, DO349, DO348, DO347, DO346, DO345, DO344,
 DO343, DO342, DO341, DO340, DO339, DO338, DO337, DO336, DO335, DO334,
 DO333, DO332, DO331, DO330, DO329, DO328, DO327, DO326, DO325, DO324,
 DO323, DO322, DO321, DO320, DO319, DO318, DO317, DO316, DO315, DO314,
 DO313, DO312, DO311, DO310, DO309, DO308, DO307, DO306, DO305, DO304,
 DO303, DO302, DO301, DO300, DO299, DO298, DO297, DO296, DO295, DO294,
 DO293, DO292, DO291, DO290, DO289, DO288, DO287, DO286, DO285, DO284,
 DO283, DO282, DO281, DO280, DO279, DO278, DO277, DO276, DO275, DO274,
 DO273, DO272, DO271, DO270, DO269, DO268, DO267, DO266, DO265, DO264,
 DO263, DO262, DO261, DO260, DO259, DO258, DO257, DO256, DO255, DO254,
 DO253, DO252, DO251, DO250, DO249, DO248, DO247, DO246, DO245, DO244,
 DO243, DO242, DO241, DO240, DO239, DO238, DO237, DO236, DO235, DO234,
 DO233, DO232, DO231, DO230, DO229, DO228, DO227, DO226, DO225, DO224,
 DO223, DO222, DO221, DO220, DO219, DO218, DO217, DO216, DO215, DO214,
 DO213, DO212, DO211, DO210, DO209, DO208, DO207, DO206, DO205, DO204,
 DO203, DO202, DO201, DO200, DO199, DO198, DO197, DO196, DO195, DO194,
 DO193, DO192, DO191, DO190, DO189, DO188, DO187, DO186, DO185, DO184,
 DO183, DO182, DO181, DO180, DO179, DO178, DO177, DO176, DO175, DO174,
 DO173, DO172, DO171, DO170, DO169, DO168, DO167, DO166, DO165, DO164,
 DO163, DO162, DO161, DO160, DO159, DO158, DO157, DO156, DO155, DO154,
 DO153, DO152, DO151, DO150, DO149, DO148, DO147, DO146, DO145, DO144,
 DO143, DO142, DO141, DO140, DO139, DO138, DO137, DO136, DO135, DO134,
 DO133, DO132, DO131, DO130, DO129, DO128, DO127, DO126, DO125, DO124,
 DO123, DO122, DO121, DO120, DO119, DO118, DO117, DO116, DO115, DO114,
 DO113, DO112, DO111, DO110, DO109, DO108, DO107, DO106, DO105, DO104,
 DO103, DO102, DO101, DO100, DO99, DO98, DO97, DO96, DO95, DO94,
 DO93, DO92, DO91, DO90, DO89, DO88, DO87, DO86, DO85, DO84,
 DO83, DO82, DO81, DO80, DO79, DO78, DO77, DO76, DO75, DO74,
 DO73, DO72, DO71, DO70, DO69, DO68, DO67, DO66, DO65, DO64,
 DO63, DO62, DO61, DO60, DO59, DO58, DO57, DO56, DO55, DO54,
 DO53, DO52, DO51, DO50, DO49, DO48, DO47, DO46, DO45, DO44,
 DO43, DO42, DO41, DO40, DO39, DO38, DO37, DO36, DO35, DO34,
 DO33, DO32, DO31, DO30, DO29, DO28, DO27, DO26, DO25, DO24,
 DO23, DO22, DO21, DO20, DO19, DO18, DO17, DO16, DO15, DO14,
 DO13, DO12, DO11, DO10, DO9, DO8, DO7, DO6, DO5, DO4,
 DO3, DO2, DO1, DO0, SYNC_OUT;
endmodule
`define _MPR4X512_
`endif
`define MPW4X512_MPR4X512
`endif
`endif
