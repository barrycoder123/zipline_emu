
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
`_2_ (* upf_always_on = 1 *) 
module ixc_gfifo_port_96_3 ( tkout, tkin, ireq, cbid, len, idata, CGFtsReq, 
	CGFcbid, CGFlen, CGFidata, CGFfull, CLBreq, CLBrd, CLBwr, CLBfull, 
	Rtkin);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output tkout;
input tkin;
input ireq;
input [19:0] cbid;
input [11:0] len;
input [95:0] idata;
output CGFtsReq;
output [19:0] CGFcbid;
output [11:0] CGFlen;
output [511:0] CGFidata;
input CGFfull;
output CLBreq;
input [3:0] CLBrd;
input [3:0] CLBwr;
input CLBfull;
input Rtkin;
wire fclk;
wire enq;
wire CLBreqWhileFull;
`_2_ wire en;
`_2_ wire ack;
`_2_ wire [95:0] odata;
`_2_ wire oreq;
`_2_ wire [19:0] ocbid;
`_2_ wire [19:0] xcbid;
`_2_ wire [11:0] olen;
`_2_ wire [11:0] xlen;
`_2_ wire [0:0] sel;
`_2_ wire [95:0] xdata;
wire [31:0] i;
`_2_ wire ireqR;
supply1 n5;
Q_BUF U0 ( .A(olen[0]), .Z(xlen[0]));
Q_BUF U1 ( .A(olen[1]), .Z(xlen[1]));
Q_BUF U2 ( .A(olen[2]), .Z(xlen[2]));
Q_BUF U3 ( .A(olen[3]), .Z(xlen[3]));
Q_BUF U4 ( .A(olen[4]), .Z(xlen[4]));
Q_BUF U5 ( .A(olen[5]), .Z(xlen[5]));
Q_BUF U6 ( .A(olen[6]), .Z(xlen[6]));
Q_BUF U7 ( .A(olen[7]), .Z(xlen[7]));
Q_BUF U8 ( .A(olen[8]), .Z(xlen[8]));
Q_BUF U9 ( .A(olen[9]), .Z(xlen[9]));
Q_BUF U10 ( .A(olen[10]), .Z(xlen[10]));
Q_BUF U11 ( .A(olen[11]), .Z(xlen[11]));
Q_BUF U12 ( .A(ocbid[0]), .Z(xcbid[0]));
Q_BUF U13 ( .A(ocbid[1]), .Z(xcbid[1]));
Q_BUF U14 ( .A(ocbid[2]), .Z(xcbid[2]));
Q_BUF U15 ( .A(ocbid[3]), .Z(xcbid[3]));
Q_BUF U16 ( .A(ocbid[4]), .Z(xcbid[4]));
Q_BUF U17 ( .A(ocbid[5]), .Z(xcbid[5]));
Q_BUF U18 ( .A(ocbid[6]), .Z(xcbid[6]));
Q_BUF U19 ( .A(ocbid[7]), .Z(xcbid[7]));
Q_BUF U20 ( .A(ocbid[8]), .Z(xcbid[8]));
Q_BUF U21 ( .A(ocbid[9]), .Z(xcbid[9]));
Q_BUF U22 ( .A(ocbid[10]), .Z(xcbid[10]));
Q_BUF U23 ( .A(ocbid[11]), .Z(xcbid[11]));
Q_BUF U24 ( .A(ocbid[12]), .Z(xcbid[12]));
Q_BUF U25 ( .A(ocbid[13]), .Z(xcbid[13]));
Q_BUF U26 ( .A(ocbid[14]), .Z(xcbid[14]));
Q_BUF U27 ( .A(ocbid[15]), .Z(xcbid[15]));
Q_BUF U28 ( .A(ocbid[16]), .Z(xcbid[16]));
Q_BUF U29 ( .A(ocbid[17]), .Z(xcbid[17]));
Q_BUF U30 ( .A(ocbid[18]), .Z(xcbid[18]));
Q_BUF U31 ( .A(ocbid[19]), .Z(xcbid[19]));
Q_BUF U32 ( .A(odata[0]), .Z(xdata[0]));
Q_BUF U33 ( .A(odata[1]), .Z(xdata[1]));
Q_BUF U34 ( .A(odata[2]), .Z(xdata[2]));
Q_BUF U35 ( .A(odata[3]), .Z(xdata[3]));
Q_BUF U36 ( .A(odata[4]), .Z(xdata[4]));
Q_BUF U37 ( .A(odata[5]), .Z(xdata[5]));
Q_BUF U38 ( .A(odata[6]), .Z(xdata[6]));
Q_BUF U39 ( .A(odata[7]), .Z(xdata[7]));
Q_BUF U40 ( .A(odata[8]), .Z(xdata[8]));
Q_BUF U41 ( .A(odata[9]), .Z(xdata[9]));
Q_BUF U42 ( .A(odata[10]), .Z(xdata[10]));
Q_BUF U43 ( .A(odata[11]), .Z(xdata[11]));
Q_BUF U44 ( .A(odata[12]), .Z(xdata[12]));
Q_BUF U45 ( .A(odata[13]), .Z(xdata[13]));
Q_BUF U46 ( .A(odata[14]), .Z(xdata[14]));
Q_BUF U47 ( .A(odata[15]), .Z(xdata[15]));
Q_BUF U48 ( .A(odata[16]), .Z(xdata[16]));
Q_BUF U49 ( .A(odata[17]), .Z(xdata[17]));
Q_BUF U50 ( .A(odata[18]), .Z(xdata[18]));
Q_BUF U51 ( .A(odata[19]), .Z(xdata[19]));
Q_BUF U52 ( .A(odata[20]), .Z(xdata[20]));
Q_BUF U53 ( .A(odata[21]), .Z(xdata[21]));
Q_BUF U54 ( .A(odata[22]), .Z(xdata[22]));
Q_BUF U55 ( .A(odata[23]), .Z(xdata[23]));
Q_BUF U56 ( .A(odata[24]), .Z(xdata[24]));
Q_BUF U57 ( .A(odata[25]), .Z(xdata[25]));
Q_BUF U58 ( .A(odata[26]), .Z(xdata[26]));
Q_BUF U59 ( .A(odata[27]), .Z(xdata[27]));
Q_BUF U60 ( .A(odata[28]), .Z(xdata[28]));
Q_BUF U61 ( .A(odata[29]), .Z(xdata[29]));
Q_BUF U62 ( .A(odata[30]), .Z(xdata[30]));
Q_BUF U63 ( .A(odata[31]), .Z(xdata[31]));
Q_BUF U64 ( .A(odata[32]), .Z(xdata[32]));
Q_BUF U65 ( .A(odata[33]), .Z(xdata[33]));
Q_BUF U66 ( .A(odata[34]), .Z(xdata[34]));
Q_BUF U67 ( .A(odata[35]), .Z(xdata[35]));
Q_BUF U68 ( .A(odata[36]), .Z(xdata[36]));
Q_BUF U69 ( .A(odata[37]), .Z(xdata[37]));
Q_BUF U70 ( .A(odata[38]), .Z(xdata[38]));
Q_BUF U71 ( .A(odata[39]), .Z(xdata[39]));
Q_BUF U72 ( .A(odata[40]), .Z(xdata[40]));
Q_BUF U73 ( .A(odata[41]), .Z(xdata[41]));
Q_BUF U74 ( .A(odata[42]), .Z(xdata[42]));
Q_BUF U75 ( .A(odata[43]), .Z(xdata[43]));
Q_BUF U76 ( .A(odata[44]), .Z(xdata[44]));
Q_BUF U77 ( .A(odata[45]), .Z(xdata[45]));
Q_BUF U78 ( .A(odata[46]), .Z(xdata[46]));
Q_BUF U79 ( .A(odata[47]), .Z(xdata[47]));
Q_BUF U80 ( .A(odata[48]), .Z(xdata[48]));
Q_BUF U81 ( .A(odata[49]), .Z(xdata[49]));
Q_BUF U82 ( .A(odata[50]), .Z(xdata[50]));
Q_BUF U83 ( .A(odata[51]), .Z(xdata[51]));
Q_BUF U84 ( .A(odata[52]), .Z(xdata[52]));
Q_BUF U85 ( .A(odata[53]), .Z(xdata[53]));
Q_BUF U86 ( .A(odata[54]), .Z(xdata[54]));
Q_BUF U87 ( .A(odata[55]), .Z(xdata[55]));
Q_BUF U88 ( .A(odata[56]), .Z(xdata[56]));
Q_BUF U89 ( .A(odata[57]), .Z(xdata[57]));
Q_BUF U90 ( .A(odata[58]), .Z(xdata[58]));
Q_BUF U91 ( .A(odata[59]), .Z(xdata[59]));
Q_BUF U92 ( .A(odata[60]), .Z(xdata[60]));
Q_BUF U93 ( .A(odata[61]), .Z(xdata[61]));
Q_BUF U94 ( .A(odata[62]), .Z(xdata[62]));
Q_BUF U95 ( .A(odata[63]), .Z(xdata[63]));
Q_BUF U96 ( .A(odata[64]), .Z(xdata[64]));
Q_BUF U97 ( .A(odata[65]), .Z(xdata[65]));
Q_BUF U98 ( .A(odata[66]), .Z(xdata[66]));
Q_BUF U99 ( .A(odata[67]), .Z(xdata[67]));
Q_BUF U100 ( .A(odata[68]), .Z(xdata[68]));
Q_BUF U101 ( .A(odata[69]), .Z(xdata[69]));
Q_BUF U102 ( .A(odata[70]), .Z(xdata[70]));
Q_BUF U103 ( .A(odata[71]), .Z(xdata[71]));
Q_BUF U104 ( .A(odata[72]), .Z(xdata[72]));
Q_BUF U105 ( .A(odata[73]), .Z(xdata[73]));
Q_BUF U106 ( .A(odata[74]), .Z(xdata[74]));
Q_BUF U107 ( .A(odata[75]), .Z(xdata[75]));
Q_BUF U108 ( .A(odata[76]), .Z(xdata[76]));
Q_BUF U109 ( .A(odata[77]), .Z(xdata[77]));
Q_BUF U110 ( .A(odata[78]), .Z(xdata[78]));
Q_BUF U111 ( .A(odata[79]), .Z(xdata[79]));
Q_BUF U112 ( .A(odata[80]), .Z(xdata[80]));
Q_BUF U113 ( .A(odata[81]), .Z(xdata[81]));
Q_BUF U114 ( .A(odata[82]), .Z(xdata[82]));
Q_BUF U115 ( .A(odata[83]), .Z(xdata[83]));
Q_BUF U116 ( .A(odata[84]), .Z(xdata[84]));
Q_BUF U117 ( .A(odata[85]), .Z(xdata[85]));
Q_BUF U118 ( .A(odata[86]), .Z(xdata[86]));
Q_BUF U119 ( .A(odata[87]), .Z(xdata[87]));
Q_BUF U120 ( .A(odata[88]), .Z(xdata[88]));
Q_BUF U121 ( .A(odata[89]), .Z(xdata[89]));
Q_BUF U122 ( .A(odata[90]), .Z(xdata[90]));
Q_BUF U123 ( .A(odata[91]), .Z(xdata[91]));
Q_BUF U124 ( .A(odata[92]), .Z(xdata[92]));
Q_BUF U125 ( .A(odata[93]), .Z(xdata[93]));
Q_BUF U126 ( .A(odata[94]), .Z(xdata[94]));
Q_BUF U127 ( .A(odata[95]), .Z(xdata[95]));
Q_NOT_TOUCH _zzqnthw ( .sig());
Q_EV_WOR_START qi ( .A(CLBreqWhileFull));
Q_INV U130 ( .A(n4), .Z(tkout));
Q_XNR2 U131 ( .A0(oreq), .A1(ack), .Z(n4));
Q_CCLKCHK cchk ( .sig(ireq));
Q_AN02 U133 ( .A0(enq), .A1(CLBfull), .Z(CLBreqWhileFull));
Q_AN02 U134 ( .A0(n2), .A1(n3), .Z(enq));
Q_INV U135 ( .A(xc_top.GFLock2), .Z(n3));
Q_XOR2 U136 ( .A0(ireq), .A1(ireqR), .Z(n2));
Q_BUFZP U137 ( .OE(CLBreqWhileFull), .A(n5), .Z(xc_top.GFLBfull));
Q_BUFZP U138 ( .OE(en), .A(xcbid[0]), .Z(CGFcbid[0]));
Q_BUFZP U139 ( .OE(en), .A(xcbid[1]), .Z(CGFcbid[1]));
Q_BUFZP U140 ( .OE(en), .A(xcbid[2]), .Z(CGFcbid[2]));
Q_BUFZP U141 ( .OE(en), .A(xcbid[3]), .Z(CGFcbid[3]));
Q_BUFZP U142 ( .OE(en), .A(xcbid[4]), .Z(CGFcbid[4]));
Q_BUFZP U143 ( .OE(en), .A(xcbid[5]), .Z(CGFcbid[5]));
Q_BUFZP U144 ( .OE(en), .A(xcbid[6]), .Z(CGFcbid[6]));
Q_BUFZP U145 ( .OE(en), .A(xcbid[7]), .Z(CGFcbid[7]));
Q_BUFZP U146 ( .OE(en), .A(xcbid[8]), .Z(CGFcbid[8]));
Q_BUFZP U147 ( .OE(en), .A(xcbid[9]), .Z(CGFcbid[9]));
Q_BUFZP U148 ( .OE(en), .A(xcbid[10]), .Z(CGFcbid[10]));
Q_BUFZP U149 ( .OE(en), .A(xcbid[11]), .Z(CGFcbid[11]));
Q_BUFZP U150 ( .OE(en), .A(xcbid[12]), .Z(CGFcbid[12]));
Q_BUFZP U151 ( .OE(en), .A(xcbid[13]), .Z(CGFcbid[13]));
Q_BUFZP U152 ( .OE(en), .A(xcbid[14]), .Z(CGFcbid[14]));
Q_BUFZP U153 ( .OE(en), .A(xcbid[15]), .Z(CGFcbid[15]));
Q_BUFZP U154 ( .OE(en), .A(xcbid[16]), .Z(CGFcbid[16]));
Q_BUFZP U155 ( .OE(en), .A(xcbid[17]), .Z(CGFcbid[17]));
Q_BUFZP U156 ( .OE(en), .A(xcbid[18]), .Z(CGFcbid[18]));
Q_BUFZP U157 ( .OE(en), .A(xcbid[19]), .Z(CGFcbid[19]));
Q_BUFZP U158 ( .OE(en), .A(xlen[0]), .Z(CGFlen[0]));
Q_BUFZP U159 ( .OE(en), .A(xlen[1]), .Z(CGFlen[1]));
Q_BUFZP U160 ( .OE(en), .A(xlen[2]), .Z(CGFlen[2]));
Q_BUFZP U161 ( .OE(en), .A(xlen[3]), .Z(CGFlen[3]));
Q_BUFZP U162 ( .OE(en), .A(xlen[4]), .Z(CGFlen[4]));
Q_BUFZP U163 ( .OE(en), .A(xlen[5]), .Z(CGFlen[5]));
Q_BUFZP U164 ( .OE(en), .A(xlen[6]), .Z(CGFlen[6]));
Q_BUFZP U165 ( .OE(en), .A(xlen[7]), .Z(CGFlen[7]));
Q_BUFZP U166 ( .OE(en), .A(xlen[8]), .Z(CGFlen[8]));
Q_BUFZP U167 ( .OE(en), .A(xlen[9]), .Z(CGFlen[9]));
Q_BUFZP U168 ( .OE(en), .A(xlen[10]), .Z(CGFlen[10]));
Q_BUFZP U169 ( .OE(en), .A(xlen[11]), .Z(CGFlen[11]));
Q_BUFZP U170 ( .OE(en), .A(xdata[0]), .Z(CGFidata[0]));
Q_BUFZP U171 ( .OE(en), .A(xdata[1]), .Z(CGFidata[1]));
Q_BUFZP U172 ( .OE(en), .A(xdata[2]), .Z(CGFidata[2]));
Q_BUFZP U173 ( .OE(en), .A(xdata[3]), .Z(CGFidata[3]));
Q_BUFZP U174 ( .OE(en), .A(xdata[4]), .Z(CGFidata[4]));
Q_BUFZP U175 ( .OE(en), .A(xdata[5]), .Z(CGFidata[5]));
Q_BUFZP U176 ( .OE(en), .A(xdata[6]), .Z(CGFidata[6]));
Q_BUFZP U177 ( .OE(en), .A(xdata[7]), .Z(CGFidata[7]));
Q_BUFZP U178 ( .OE(en), .A(xdata[8]), .Z(CGFidata[8]));
Q_BUFZP U179 ( .OE(en), .A(xdata[9]), .Z(CGFidata[9]));
Q_BUFZP U180 ( .OE(en), .A(xdata[10]), .Z(CGFidata[10]));
Q_BUFZP U181 ( .OE(en), .A(xdata[11]), .Z(CGFidata[11]));
Q_BUFZP U182 ( .OE(en), .A(xdata[12]), .Z(CGFidata[12]));
Q_BUFZP U183 ( .OE(en), .A(xdata[13]), .Z(CGFidata[13]));
Q_BUFZP U184 ( .OE(en), .A(xdata[14]), .Z(CGFidata[14]));
Q_BUFZP U185 ( .OE(en), .A(xdata[15]), .Z(CGFidata[15]));
Q_BUFZP U186 ( .OE(en), .A(xdata[16]), .Z(CGFidata[16]));
Q_BUFZP U187 ( .OE(en), .A(xdata[17]), .Z(CGFidata[17]));
Q_BUFZP U188 ( .OE(en), .A(xdata[18]), .Z(CGFidata[18]));
Q_BUFZP U189 ( .OE(en), .A(xdata[19]), .Z(CGFidata[19]));
Q_BUFZP U190 ( .OE(en), .A(xdata[20]), .Z(CGFidata[20]));
Q_BUFZP U191 ( .OE(en), .A(xdata[21]), .Z(CGFidata[21]));
Q_BUFZP U192 ( .OE(en), .A(xdata[22]), .Z(CGFidata[22]));
Q_BUFZP U193 ( .OE(en), .A(xdata[23]), .Z(CGFidata[23]));
Q_BUFZP U194 ( .OE(en), .A(xdata[24]), .Z(CGFidata[24]));
Q_BUFZP U195 ( .OE(en), .A(xdata[25]), .Z(CGFidata[25]));
Q_BUFZP U196 ( .OE(en), .A(xdata[26]), .Z(CGFidata[26]));
Q_BUFZP U197 ( .OE(en), .A(xdata[27]), .Z(CGFidata[27]));
Q_BUFZP U198 ( .OE(en), .A(xdata[28]), .Z(CGFidata[28]));
Q_BUFZP U199 ( .OE(en), .A(xdata[29]), .Z(CGFidata[29]));
Q_BUFZP U200 ( .OE(en), .A(xdata[30]), .Z(CGFidata[30]));
Q_BUFZP U201 ( .OE(en), .A(xdata[31]), .Z(CGFidata[31]));
Q_BUFZP U202 ( .OE(en), .A(xdata[32]), .Z(CGFidata[32]));
Q_BUFZP U203 ( .OE(en), .A(xdata[33]), .Z(CGFidata[33]));
Q_BUFZP U204 ( .OE(en), .A(xdata[34]), .Z(CGFidata[34]));
Q_BUFZP U205 ( .OE(en), .A(xdata[35]), .Z(CGFidata[35]));
Q_BUFZP U206 ( .OE(en), .A(xdata[36]), .Z(CGFidata[36]));
Q_BUFZP U207 ( .OE(en), .A(xdata[37]), .Z(CGFidata[37]));
Q_BUFZP U208 ( .OE(en), .A(xdata[38]), .Z(CGFidata[38]));
Q_BUFZP U209 ( .OE(en), .A(xdata[39]), .Z(CGFidata[39]));
Q_BUFZP U210 ( .OE(en), .A(xdata[40]), .Z(CGFidata[40]));
Q_BUFZP U211 ( .OE(en), .A(xdata[41]), .Z(CGFidata[41]));
Q_BUFZP U212 ( .OE(en), .A(xdata[42]), .Z(CGFidata[42]));
Q_BUFZP U213 ( .OE(en), .A(xdata[43]), .Z(CGFidata[43]));
Q_BUFZP U214 ( .OE(en), .A(xdata[44]), .Z(CGFidata[44]));
Q_BUFZP U215 ( .OE(en), .A(xdata[45]), .Z(CGFidata[45]));
Q_BUFZP U216 ( .OE(en), .A(xdata[46]), .Z(CGFidata[46]));
Q_BUFZP U217 ( .OE(en), .A(xdata[47]), .Z(CGFidata[47]));
Q_BUFZP U218 ( .OE(en), .A(xdata[48]), .Z(CGFidata[48]));
Q_BUFZP U219 ( .OE(en), .A(xdata[49]), .Z(CGFidata[49]));
Q_BUFZP U220 ( .OE(en), .A(xdata[50]), .Z(CGFidata[50]));
Q_BUFZP U221 ( .OE(en), .A(xdata[51]), .Z(CGFidata[51]));
Q_BUFZP U222 ( .OE(en), .A(xdata[52]), .Z(CGFidata[52]));
Q_BUFZP U223 ( .OE(en), .A(xdata[53]), .Z(CGFidata[53]));
Q_BUFZP U224 ( .OE(en), .A(xdata[54]), .Z(CGFidata[54]));
Q_BUFZP U225 ( .OE(en), .A(xdata[55]), .Z(CGFidata[55]));
Q_BUFZP U226 ( .OE(en), .A(xdata[56]), .Z(CGFidata[56]));
Q_BUFZP U227 ( .OE(en), .A(xdata[57]), .Z(CGFidata[57]));
Q_BUFZP U228 ( .OE(en), .A(xdata[58]), .Z(CGFidata[58]));
Q_BUFZP U229 ( .OE(en), .A(xdata[59]), .Z(CGFidata[59]));
Q_BUFZP U230 ( .OE(en), .A(xdata[60]), .Z(CGFidata[60]));
Q_BUFZP U231 ( .OE(en), .A(xdata[61]), .Z(CGFidata[61]));
Q_BUFZP U232 ( .OE(en), .A(xdata[62]), .Z(CGFidata[62]));
Q_BUFZP U233 ( .OE(en), .A(xdata[63]), .Z(CGFidata[63]));
Q_BUFZP U234 ( .OE(en), .A(xdata[64]), .Z(CGFidata[64]));
Q_BUFZP U235 ( .OE(en), .A(xdata[65]), .Z(CGFidata[65]));
Q_BUFZP U236 ( .OE(en), .A(xdata[66]), .Z(CGFidata[66]));
Q_BUFZP U237 ( .OE(en), .A(xdata[67]), .Z(CGFidata[67]));
Q_BUFZP U238 ( .OE(en), .A(xdata[68]), .Z(CGFidata[68]));
Q_BUFZP U239 ( .OE(en), .A(xdata[69]), .Z(CGFidata[69]));
Q_BUFZP U240 ( .OE(en), .A(xdata[70]), .Z(CGFidata[70]));
Q_BUFZP U241 ( .OE(en), .A(xdata[71]), .Z(CGFidata[71]));
Q_BUFZP U242 ( .OE(en), .A(xdata[72]), .Z(CGFidata[72]));
Q_BUFZP U243 ( .OE(en), .A(xdata[73]), .Z(CGFidata[73]));
Q_BUFZP U244 ( .OE(en), .A(xdata[74]), .Z(CGFidata[74]));
Q_BUFZP U245 ( .OE(en), .A(xdata[75]), .Z(CGFidata[75]));
Q_BUFZP U246 ( .OE(en), .A(xdata[76]), .Z(CGFidata[76]));
Q_BUFZP U247 ( .OE(en), .A(xdata[77]), .Z(CGFidata[77]));
Q_BUFZP U248 ( .OE(en), .A(xdata[78]), .Z(CGFidata[78]));
Q_BUFZP U249 ( .OE(en), .A(xdata[79]), .Z(CGFidata[79]));
Q_BUFZP U250 ( .OE(en), .A(xdata[80]), .Z(CGFidata[80]));
Q_BUFZP U251 ( .OE(en), .A(xdata[81]), .Z(CGFidata[81]));
Q_BUFZP U252 ( .OE(en), .A(xdata[82]), .Z(CGFidata[82]));
Q_BUFZP U253 ( .OE(en), .A(xdata[83]), .Z(CGFidata[83]));
Q_BUFZP U254 ( .OE(en), .A(xdata[84]), .Z(CGFidata[84]));
Q_BUFZP U255 ( .OE(en), .A(xdata[85]), .Z(CGFidata[85]));
Q_BUFZP U256 ( .OE(en), .A(xdata[86]), .Z(CGFidata[86]));
Q_BUFZP U257 ( .OE(en), .A(xdata[87]), .Z(CGFidata[87]));
Q_BUFZP U258 ( .OE(en), .A(xdata[88]), .Z(CGFidata[88]));
Q_BUFZP U259 ( .OE(en), .A(xdata[89]), .Z(CGFidata[89]));
Q_BUFZP U260 ( .OE(en), .A(xdata[90]), .Z(CGFidata[90]));
Q_BUFZP U261 ( .OE(en), .A(xdata[91]), .Z(CGFidata[91]));
Q_BUFZP U262 ( .OE(en), .A(xdata[92]), .Z(CGFidata[92]));
Q_BUFZP U263 ( .OE(en), .A(xdata[93]), .Z(CGFidata[93]));
Q_BUFZP U264 ( .OE(en), .A(xdata[94]), .Z(CGFidata[94]));
Q_BUFZP U265 ( .OE(en), .A(xdata[95]), .Z(CGFidata[95]));
Q_BUFZP U266 ( .OE(enq), .A(n5), .Z(CLBreq));
Q_BUFZP U267 ( .OE(enq), .A(n5), .Z(CGFtsReq));
Q_INV U268 ( .A(CLBwr[2]), .Z(n6));
ixc_bind \genblk3.b5 ( CLBfull, IXC_GFIFO.O.O.LBfull);
ixc_bind_4 \genblk3.b4 ( CLBwr[3:0], IXC_GFIFO.O.O.LBwr[3:0]);
ixc_bind_4 \genblk3.b3 ( CLBrd[3:0], IXC_GFIFO.O.O.LBrd[3:0]);
ixc_bind \genblk3.b2 ( CLBreq, IXC_GFIFO.O.O.LBreq);
ixc_bind \genblk3.b1 ( CGFfull, IXC_GFIFO.O.O.GFfull);
ixc_bind \genblk3.b0 ( CGFtsReq, IXC_GFIFO.O.O.GFtsReq);
Q_MX02 U275 ( .S(xc_top.GFLock2), .A0(oreq), .A1(ireq), .Z(n8));
Q_FDP0UA U276 ( .D(n9), .QTFCLK( ), .Q(ack));
Q_MX02 U277 ( .S(n14), .A0(ack), .A1(n8), .Z(n9));
Q_FDP0UA U278 ( .D(n10), .QTFCLK( ), .Q(en));
Q_NR02 U279 ( .A0(xc_top.GFLock2), .A1(n11), .Z(n10));
Q_OR02 U280 ( .A0(xc_top.GFLock2), .A1(n12), .Z(n14));
Q_INV U281 ( .A(n11), .Z(n12));
Q_OR03 U282 ( .A0(n4), .A1(tkin), .A2(n13), .Z(n11));
Q_OR02 U283 ( .A0(Rtkin), .A1(CGFfull), .Z(n13));
Q_MX02 U284 ( .S(CLBfull), .A0(ireq), .A1(ireqR), .Z(n15));
Q_FDP0UA U285 ( .D(n15), .QTFCLK( ), .Q(ireqR));
Q_AN02 U286 ( .A0(CLBwr[0]), .A1(n6), .Z(n16));
Q_AN02 U287 ( .A0(CLBwr[1]), .A1(n6), .Z(n17));
Q_INV U288 ( .A(n16), .Z(n18));
Q_INV U289 ( .A(n17), .Z(n19));
Q_NR02 U290 ( .A0(n17), .A1(n16), .Z(n20));
Q_AN02 U291 ( .A0(n19), .A1(n16), .Z(n21));
Q_AN02 U292 ( .A0(n17), .A1(n18), .Z(n22));
Q_AN02 U293 ( .A0(n17), .A1(n16), .Z(n23));
Q_AN02 U294 ( .A0(n20), .A1(n6), .Z(n24));
Q_LDP0 \_zzLB_REG[0][0] ( .G(n24), .D(len[0]), .Q(\_zzLB[0][0] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][1] ( .G(n24), .D(len[1]), .Q(\_zzLB[0][1] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][2] ( .G(n24), .D(len[2]), .Q(\_zzLB[0][2] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][3] ( .G(n24), .D(len[3]), .Q(\_zzLB[0][3] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][4] ( .G(n24), .D(len[4]), .Q(\_zzLB[0][4] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][5] ( .G(n24), .D(len[5]), .Q(\_zzLB[0][5] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][6] ( .G(n24), .D(len[6]), .Q(\_zzLB[0][6] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][7] ( .G(n24), .D(len[7]), .Q(\_zzLB[0][7] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][8] ( .G(n24), .D(len[8]), .Q(\_zzLB[0][8] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][9] ( .G(n24), .D(len[9]), .Q(\_zzLB[0][9] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][10] ( .G(n24), .D(len[10]), .Q(\_zzLB[0][10] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][11] ( .G(n24), .D(len[11]), .Q(\_zzLB[0][11] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][12] ( .G(n24), .D(cbid[0]), .Q(\_zzLB[0][12] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][13] ( .G(n24), .D(cbid[1]), .Q(\_zzLB[0][13] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][14] ( .G(n24), .D(cbid[2]), .Q(\_zzLB[0][14] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][15] ( .G(n24), .D(cbid[3]), .Q(\_zzLB[0][15] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][16] ( .G(n24), .D(cbid[4]), .Q(\_zzLB[0][16] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][17] ( .G(n24), .D(cbid[5]), .Q(\_zzLB[0][17] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][18] ( .G(n24), .D(cbid[6]), .Q(\_zzLB[0][18] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][19] ( .G(n24), .D(cbid[7]), .Q(\_zzLB[0][19] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][20] ( .G(n24), .D(cbid[8]), .Q(\_zzLB[0][20] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][21] ( .G(n24), .D(cbid[9]), .Q(\_zzLB[0][21] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][22] ( .G(n24), .D(cbid[10]), .Q(\_zzLB[0][22] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][23] ( .G(n24), .D(cbid[11]), .Q(\_zzLB[0][23] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][24] ( .G(n24), .D(cbid[12]), .Q(\_zzLB[0][24] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][25] ( .G(n24), .D(cbid[13]), .Q(\_zzLB[0][25] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][26] ( .G(n24), .D(cbid[14]), .Q(\_zzLB[0][26] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][27] ( .G(n24), .D(cbid[15]), .Q(\_zzLB[0][27] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][28] ( .G(n24), .D(cbid[16]), .Q(\_zzLB[0][28] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][29] ( .G(n24), .D(cbid[17]), .Q(\_zzLB[0][29] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][30] ( .G(n24), .D(cbid[18]), .Q(\_zzLB[0][30] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][31] ( .G(n24), .D(cbid[19]), .Q(\_zzLB[0][31] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][32] ( .G(n24), .D(idata[0]), .Q(\_zzLB[0][32] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][33] ( .G(n24), .D(idata[1]), .Q(\_zzLB[0][33] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][34] ( .G(n24), .D(idata[2]), .Q(\_zzLB[0][34] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][35] ( .G(n24), .D(idata[3]), .Q(\_zzLB[0][35] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][36] ( .G(n24), .D(idata[4]), .Q(\_zzLB[0][36] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][37] ( .G(n24), .D(idata[5]), .Q(\_zzLB[0][37] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][38] ( .G(n24), .D(idata[6]), .Q(\_zzLB[0][38] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][39] ( .G(n24), .D(idata[7]), .Q(\_zzLB[0][39] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][40] ( .G(n24), .D(idata[8]), .Q(\_zzLB[0][40] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][41] ( .G(n24), .D(idata[9]), .Q(\_zzLB[0][41] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][42] ( .G(n24), .D(idata[10]), .Q(\_zzLB[0][42] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][43] ( .G(n24), .D(idata[11]), .Q(\_zzLB[0][43] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][44] ( .G(n24), .D(idata[12]), .Q(\_zzLB[0][44] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][45] ( .G(n24), .D(idata[13]), .Q(\_zzLB[0][45] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][46] ( .G(n24), .D(idata[14]), .Q(\_zzLB[0][46] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][47] ( .G(n24), .D(idata[15]), .Q(\_zzLB[0][47] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][48] ( .G(n24), .D(idata[16]), .Q(\_zzLB[0][48] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][49] ( .G(n24), .D(idata[17]), .Q(\_zzLB[0][49] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][50] ( .G(n24), .D(idata[18]), .Q(\_zzLB[0][50] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][51] ( .G(n24), .D(idata[19]), .Q(\_zzLB[0][51] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][52] ( .G(n24), .D(idata[20]), .Q(\_zzLB[0][52] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][53] ( .G(n24), .D(idata[21]), .Q(\_zzLB[0][53] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][54] ( .G(n24), .D(idata[22]), .Q(\_zzLB[0][54] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][55] ( .G(n24), .D(idata[23]), .Q(\_zzLB[0][55] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][56] ( .G(n24), .D(idata[24]), .Q(\_zzLB[0][56] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][57] ( .G(n24), .D(idata[25]), .Q(\_zzLB[0][57] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][58] ( .G(n24), .D(idata[26]), .Q(\_zzLB[0][58] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][59] ( .G(n24), .D(idata[27]), .Q(\_zzLB[0][59] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][60] ( .G(n24), .D(idata[28]), .Q(\_zzLB[0][60] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][61] ( .G(n24), .D(idata[29]), .Q(\_zzLB[0][61] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][62] ( .G(n24), .D(idata[30]), .Q(\_zzLB[0][62] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][63] ( .G(n24), .D(idata[31]), .Q(\_zzLB[0][63] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][64] ( .G(n24), .D(idata[32]), .Q(\_zzLB[0][64] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][65] ( .G(n24), .D(idata[33]), .Q(\_zzLB[0][65] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][66] ( .G(n24), .D(idata[34]), .Q(\_zzLB[0][66] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][67] ( .G(n24), .D(idata[35]), .Q(\_zzLB[0][67] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][68] ( .G(n24), .D(idata[36]), .Q(\_zzLB[0][68] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][69] ( .G(n24), .D(idata[37]), .Q(\_zzLB[0][69] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][70] ( .G(n24), .D(idata[38]), .Q(\_zzLB[0][70] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][71] ( .G(n24), .D(idata[39]), .Q(\_zzLB[0][71] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][72] ( .G(n24), .D(idata[40]), .Q(\_zzLB[0][72] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][73] ( .G(n24), .D(idata[41]), .Q(\_zzLB[0][73] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][74] ( .G(n24), .D(idata[42]), .Q(\_zzLB[0][74] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][75] ( .G(n24), .D(idata[43]), .Q(\_zzLB[0][75] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][76] ( .G(n24), .D(idata[44]), .Q(\_zzLB[0][76] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][77] ( .G(n24), .D(idata[45]), .Q(\_zzLB[0][77] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][78] ( .G(n24), .D(idata[46]), .Q(\_zzLB[0][78] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][79] ( .G(n24), .D(idata[47]), .Q(\_zzLB[0][79] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][80] ( .G(n24), .D(idata[48]), .Q(\_zzLB[0][80] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][81] ( .G(n24), .D(idata[49]), .Q(\_zzLB[0][81] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][82] ( .G(n24), .D(idata[50]), .Q(\_zzLB[0][82] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][83] ( .G(n24), .D(idata[51]), .Q(\_zzLB[0][83] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][84] ( .G(n24), .D(idata[52]), .Q(\_zzLB[0][84] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][85] ( .G(n24), .D(idata[53]), .Q(\_zzLB[0][85] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][86] ( .G(n24), .D(idata[54]), .Q(\_zzLB[0][86] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][87] ( .G(n24), .D(idata[55]), .Q(\_zzLB[0][87] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][88] ( .G(n24), .D(idata[56]), .Q(\_zzLB[0][88] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][89] ( .G(n24), .D(idata[57]), .Q(\_zzLB[0][89] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][90] ( .G(n24), .D(idata[58]), .Q(\_zzLB[0][90] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][91] ( .G(n24), .D(idata[59]), .Q(\_zzLB[0][91] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][92] ( .G(n24), .D(idata[60]), .Q(\_zzLB[0][92] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][93] ( .G(n24), .D(idata[61]), .Q(\_zzLB[0][93] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][94] ( .G(n24), .D(idata[62]), .Q(\_zzLB[0][94] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][95] ( .G(n24), .D(idata[63]), .Q(\_zzLB[0][95] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][96] ( .G(n24), .D(idata[64]), .Q(\_zzLB[0][96] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][97] ( .G(n24), .D(idata[65]), .Q(\_zzLB[0][97] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][98] ( .G(n24), .D(idata[66]), .Q(\_zzLB[0][98] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][99] ( .G(n24), .D(idata[67]), .Q(\_zzLB[0][99] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][100] ( .G(n24), .D(idata[68]), .Q(\_zzLB[0][100] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][101] ( .G(n24), .D(idata[69]), .Q(\_zzLB[0][101] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][102] ( .G(n24), .D(idata[70]), .Q(\_zzLB[0][102] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][103] ( .G(n24), .D(idata[71]), .Q(\_zzLB[0][103] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][104] ( .G(n24), .D(idata[72]), .Q(\_zzLB[0][104] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][105] ( .G(n24), .D(idata[73]), .Q(\_zzLB[0][105] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][106] ( .G(n24), .D(idata[74]), .Q(\_zzLB[0][106] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][107] ( .G(n24), .D(idata[75]), .Q(\_zzLB[0][107] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][108] ( .G(n24), .D(idata[76]), .Q(\_zzLB[0][108] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][109] ( .G(n24), .D(idata[77]), .Q(\_zzLB[0][109] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][110] ( .G(n24), .D(idata[78]), .Q(\_zzLB[0][110] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][111] ( .G(n24), .D(idata[79]), .Q(\_zzLB[0][111] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][112] ( .G(n24), .D(idata[80]), .Q(\_zzLB[0][112] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][113] ( .G(n24), .D(idata[81]), .Q(\_zzLB[0][113] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][114] ( .G(n24), .D(idata[82]), .Q(\_zzLB[0][114] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][115] ( .G(n24), .D(idata[83]), .Q(\_zzLB[0][115] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][116] ( .G(n24), .D(idata[84]), .Q(\_zzLB[0][116] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][117] ( .G(n24), .D(idata[85]), .Q(\_zzLB[0][117] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][118] ( .G(n24), .D(idata[86]), .Q(\_zzLB[0][118] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][119] ( .G(n24), .D(idata[87]), .Q(\_zzLB[0][119] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][120] ( .G(n24), .D(idata[88]), .Q(\_zzLB[0][120] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][121] ( .G(n24), .D(idata[89]), .Q(\_zzLB[0][121] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][122] ( .G(n24), .D(idata[90]), .Q(\_zzLB[0][122] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][123] ( .G(n24), .D(idata[91]), .Q(\_zzLB[0][123] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][124] ( .G(n24), .D(idata[92]), .Q(\_zzLB[0][124] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][125] ( .G(n24), .D(idata[93]), .Q(\_zzLB[0][125] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][126] ( .G(n24), .D(idata[94]), .Q(\_zzLB[0][126] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][127] ( .G(n24), .D(idata[95]), .Q(\_zzLB[0][127] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][128] ( .G(n24), .D(ireq), .Q(\_zzLB[0][128] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][0] ( .G(n21), .D(len[0]), .Q(\_zzLB[1][0] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][1] ( .G(n21), .D(len[1]), .Q(\_zzLB[1][1] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][2] ( .G(n21), .D(len[2]), .Q(\_zzLB[1][2] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][3] ( .G(n21), .D(len[3]), .Q(\_zzLB[1][3] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][4] ( .G(n21), .D(len[4]), .Q(\_zzLB[1][4] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][5] ( .G(n21), .D(len[5]), .Q(\_zzLB[1][5] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][6] ( .G(n21), .D(len[6]), .Q(\_zzLB[1][6] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][7] ( .G(n21), .D(len[7]), .Q(\_zzLB[1][7] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][8] ( .G(n21), .D(len[8]), .Q(\_zzLB[1][8] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][9] ( .G(n21), .D(len[9]), .Q(\_zzLB[1][9] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][10] ( .G(n21), .D(len[10]), .Q(\_zzLB[1][10] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][11] ( .G(n21), .D(len[11]), .Q(\_zzLB[1][11] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][12] ( .G(n21), .D(cbid[0]), .Q(\_zzLB[1][12] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][13] ( .G(n21), .D(cbid[1]), .Q(\_zzLB[1][13] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][14] ( .G(n21), .D(cbid[2]), .Q(\_zzLB[1][14] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][15] ( .G(n21), .D(cbid[3]), .Q(\_zzLB[1][15] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][16] ( .G(n21), .D(cbid[4]), .Q(\_zzLB[1][16] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][17] ( .G(n21), .D(cbid[5]), .Q(\_zzLB[1][17] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][18] ( .G(n21), .D(cbid[6]), .Q(\_zzLB[1][18] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][19] ( .G(n21), .D(cbid[7]), .Q(\_zzLB[1][19] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][20] ( .G(n21), .D(cbid[8]), .Q(\_zzLB[1][20] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][21] ( .G(n21), .D(cbid[9]), .Q(\_zzLB[1][21] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][22] ( .G(n21), .D(cbid[10]), .Q(\_zzLB[1][22] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][23] ( .G(n21), .D(cbid[11]), .Q(\_zzLB[1][23] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][24] ( .G(n21), .D(cbid[12]), .Q(\_zzLB[1][24] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][25] ( .G(n21), .D(cbid[13]), .Q(\_zzLB[1][25] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][26] ( .G(n21), .D(cbid[14]), .Q(\_zzLB[1][26] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][27] ( .G(n21), .D(cbid[15]), .Q(\_zzLB[1][27] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][28] ( .G(n21), .D(cbid[16]), .Q(\_zzLB[1][28] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][29] ( .G(n21), .D(cbid[17]), .Q(\_zzLB[1][29] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][30] ( .G(n21), .D(cbid[18]), .Q(\_zzLB[1][30] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][31] ( .G(n21), .D(cbid[19]), .Q(\_zzLB[1][31] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][32] ( .G(n21), .D(idata[0]), .Q(\_zzLB[1][32] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][33] ( .G(n21), .D(idata[1]), .Q(\_zzLB[1][33] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][34] ( .G(n21), .D(idata[2]), .Q(\_zzLB[1][34] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][35] ( .G(n21), .D(idata[3]), .Q(\_zzLB[1][35] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][36] ( .G(n21), .D(idata[4]), .Q(\_zzLB[1][36] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][37] ( .G(n21), .D(idata[5]), .Q(\_zzLB[1][37] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][38] ( .G(n21), .D(idata[6]), .Q(\_zzLB[1][38] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][39] ( .G(n21), .D(idata[7]), .Q(\_zzLB[1][39] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][40] ( .G(n21), .D(idata[8]), .Q(\_zzLB[1][40] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][41] ( .G(n21), .D(idata[9]), .Q(\_zzLB[1][41] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][42] ( .G(n21), .D(idata[10]), .Q(\_zzLB[1][42] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][43] ( .G(n21), .D(idata[11]), .Q(\_zzLB[1][43] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][44] ( .G(n21), .D(idata[12]), .Q(\_zzLB[1][44] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][45] ( .G(n21), .D(idata[13]), .Q(\_zzLB[1][45] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][46] ( .G(n21), .D(idata[14]), .Q(\_zzLB[1][46] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][47] ( .G(n21), .D(idata[15]), .Q(\_zzLB[1][47] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][48] ( .G(n21), .D(idata[16]), .Q(\_zzLB[1][48] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][49] ( .G(n21), .D(idata[17]), .Q(\_zzLB[1][49] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][50] ( .G(n21), .D(idata[18]), .Q(\_zzLB[1][50] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][51] ( .G(n21), .D(idata[19]), .Q(\_zzLB[1][51] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][52] ( .G(n21), .D(idata[20]), .Q(\_zzLB[1][52] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][53] ( .G(n21), .D(idata[21]), .Q(\_zzLB[1][53] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][54] ( .G(n21), .D(idata[22]), .Q(\_zzLB[1][54] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][55] ( .G(n21), .D(idata[23]), .Q(\_zzLB[1][55] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][56] ( .G(n21), .D(idata[24]), .Q(\_zzLB[1][56] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][57] ( .G(n21), .D(idata[25]), .Q(\_zzLB[1][57] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][58] ( .G(n21), .D(idata[26]), .Q(\_zzLB[1][58] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][59] ( .G(n21), .D(idata[27]), .Q(\_zzLB[1][59] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][60] ( .G(n21), .D(idata[28]), .Q(\_zzLB[1][60] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][61] ( .G(n21), .D(idata[29]), .Q(\_zzLB[1][61] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][62] ( .G(n21), .D(idata[30]), .Q(\_zzLB[1][62] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][63] ( .G(n21), .D(idata[31]), .Q(\_zzLB[1][63] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][64] ( .G(n21), .D(idata[32]), .Q(\_zzLB[1][64] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][65] ( .G(n21), .D(idata[33]), .Q(\_zzLB[1][65] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][66] ( .G(n21), .D(idata[34]), .Q(\_zzLB[1][66] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][67] ( .G(n21), .D(idata[35]), .Q(\_zzLB[1][67] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][68] ( .G(n21), .D(idata[36]), .Q(\_zzLB[1][68] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][69] ( .G(n21), .D(idata[37]), .Q(\_zzLB[1][69] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][70] ( .G(n21), .D(idata[38]), .Q(\_zzLB[1][70] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][71] ( .G(n21), .D(idata[39]), .Q(\_zzLB[1][71] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][72] ( .G(n21), .D(idata[40]), .Q(\_zzLB[1][72] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][73] ( .G(n21), .D(idata[41]), .Q(\_zzLB[1][73] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][74] ( .G(n21), .D(idata[42]), .Q(\_zzLB[1][74] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][75] ( .G(n21), .D(idata[43]), .Q(\_zzLB[1][75] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][76] ( .G(n21), .D(idata[44]), .Q(\_zzLB[1][76] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][77] ( .G(n21), .D(idata[45]), .Q(\_zzLB[1][77] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][78] ( .G(n21), .D(idata[46]), .Q(\_zzLB[1][78] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][79] ( .G(n21), .D(idata[47]), .Q(\_zzLB[1][79] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][80] ( .G(n21), .D(idata[48]), .Q(\_zzLB[1][80] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][81] ( .G(n21), .D(idata[49]), .Q(\_zzLB[1][81] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][82] ( .G(n21), .D(idata[50]), .Q(\_zzLB[1][82] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][83] ( .G(n21), .D(idata[51]), .Q(\_zzLB[1][83] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][84] ( .G(n21), .D(idata[52]), .Q(\_zzLB[1][84] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][85] ( .G(n21), .D(idata[53]), .Q(\_zzLB[1][85] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][86] ( .G(n21), .D(idata[54]), .Q(\_zzLB[1][86] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][87] ( .G(n21), .D(idata[55]), .Q(\_zzLB[1][87] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][88] ( .G(n21), .D(idata[56]), .Q(\_zzLB[1][88] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][89] ( .G(n21), .D(idata[57]), .Q(\_zzLB[1][89] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][90] ( .G(n21), .D(idata[58]), .Q(\_zzLB[1][90] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][91] ( .G(n21), .D(idata[59]), .Q(\_zzLB[1][91] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][92] ( .G(n21), .D(idata[60]), .Q(\_zzLB[1][92] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][93] ( .G(n21), .D(idata[61]), .Q(\_zzLB[1][93] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][94] ( .G(n21), .D(idata[62]), .Q(\_zzLB[1][94] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][95] ( .G(n21), .D(idata[63]), .Q(\_zzLB[1][95] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][96] ( .G(n21), .D(idata[64]), .Q(\_zzLB[1][96] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][97] ( .G(n21), .D(idata[65]), .Q(\_zzLB[1][97] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][98] ( .G(n21), .D(idata[66]), .Q(\_zzLB[1][98] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][99] ( .G(n21), .D(idata[67]), .Q(\_zzLB[1][99] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][100] ( .G(n21), .D(idata[68]), .Q(\_zzLB[1][100] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][101] ( .G(n21), .D(idata[69]), .Q(\_zzLB[1][101] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][102] ( .G(n21), .D(idata[70]), .Q(\_zzLB[1][102] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][103] ( .G(n21), .D(idata[71]), .Q(\_zzLB[1][103] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][104] ( .G(n21), .D(idata[72]), .Q(\_zzLB[1][104] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][105] ( .G(n21), .D(idata[73]), .Q(\_zzLB[1][105] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][106] ( .G(n21), .D(idata[74]), .Q(\_zzLB[1][106] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][107] ( .G(n21), .D(idata[75]), .Q(\_zzLB[1][107] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][108] ( .G(n21), .D(idata[76]), .Q(\_zzLB[1][108] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][109] ( .G(n21), .D(idata[77]), .Q(\_zzLB[1][109] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][110] ( .G(n21), .D(idata[78]), .Q(\_zzLB[1][110] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][111] ( .G(n21), .D(idata[79]), .Q(\_zzLB[1][111] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][112] ( .G(n21), .D(idata[80]), .Q(\_zzLB[1][112] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][113] ( .G(n21), .D(idata[81]), .Q(\_zzLB[1][113] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][114] ( .G(n21), .D(idata[82]), .Q(\_zzLB[1][114] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][115] ( .G(n21), .D(idata[83]), .Q(\_zzLB[1][115] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][116] ( .G(n21), .D(idata[84]), .Q(\_zzLB[1][116] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][117] ( .G(n21), .D(idata[85]), .Q(\_zzLB[1][117] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][118] ( .G(n21), .D(idata[86]), .Q(\_zzLB[1][118] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][119] ( .G(n21), .D(idata[87]), .Q(\_zzLB[1][119] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][120] ( .G(n21), .D(idata[88]), .Q(\_zzLB[1][120] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][121] ( .G(n21), .D(idata[89]), .Q(\_zzLB[1][121] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][122] ( .G(n21), .D(idata[90]), .Q(\_zzLB[1][122] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][123] ( .G(n21), .D(idata[91]), .Q(\_zzLB[1][123] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][124] ( .G(n21), .D(idata[92]), .Q(\_zzLB[1][124] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][125] ( .G(n21), .D(idata[93]), .Q(\_zzLB[1][125] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][126] ( .G(n21), .D(idata[94]), .Q(\_zzLB[1][126] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][127] ( .G(n21), .D(idata[95]), .Q(\_zzLB[1][127] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][128] ( .G(n21), .D(ireq), .Q(\_zzLB[1][128] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][0] ( .G(n22), .D(len[0]), .Q(\_zzLB[2][0] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][1] ( .G(n22), .D(len[1]), .Q(\_zzLB[2][1] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][2] ( .G(n22), .D(len[2]), .Q(\_zzLB[2][2] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][3] ( .G(n22), .D(len[3]), .Q(\_zzLB[2][3] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][4] ( .G(n22), .D(len[4]), .Q(\_zzLB[2][4] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][5] ( .G(n22), .D(len[5]), .Q(\_zzLB[2][5] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][6] ( .G(n22), .D(len[6]), .Q(\_zzLB[2][6] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][7] ( .G(n22), .D(len[7]), .Q(\_zzLB[2][7] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][8] ( .G(n22), .D(len[8]), .Q(\_zzLB[2][8] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][9] ( .G(n22), .D(len[9]), .Q(\_zzLB[2][9] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][10] ( .G(n22), .D(len[10]), .Q(\_zzLB[2][10] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][11] ( .G(n22), .D(len[11]), .Q(\_zzLB[2][11] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][12] ( .G(n22), .D(cbid[0]), .Q(\_zzLB[2][12] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][13] ( .G(n22), .D(cbid[1]), .Q(\_zzLB[2][13] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][14] ( .G(n22), .D(cbid[2]), .Q(\_zzLB[2][14] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][15] ( .G(n22), .D(cbid[3]), .Q(\_zzLB[2][15] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][16] ( .G(n22), .D(cbid[4]), .Q(\_zzLB[2][16] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][17] ( .G(n22), .D(cbid[5]), .Q(\_zzLB[2][17] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][18] ( .G(n22), .D(cbid[6]), .Q(\_zzLB[2][18] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][19] ( .G(n22), .D(cbid[7]), .Q(\_zzLB[2][19] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][20] ( .G(n22), .D(cbid[8]), .Q(\_zzLB[2][20] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][21] ( .G(n22), .D(cbid[9]), .Q(\_zzLB[2][21] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][22] ( .G(n22), .D(cbid[10]), .Q(\_zzLB[2][22] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][23] ( .G(n22), .D(cbid[11]), .Q(\_zzLB[2][23] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][24] ( .G(n22), .D(cbid[12]), .Q(\_zzLB[2][24] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][25] ( .G(n22), .D(cbid[13]), .Q(\_zzLB[2][25] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][26] ( .G(n22), .D(cbid[14]), .Q(\_zzLB[2][26] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][27] ( .G(n22), .D(cbid[15]), .Q(\_zzLB[2][27] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][28] ( .G(n22), .D(cbid[16]), .Q(\_zzLB[2][28] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][29] ( .G(n22), .D(cbid[17]), .Q(\_zzLB[2][29] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][30] ( .G(n22), .D(cbid[18]), .Q(\_zzLB[2][30] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][31] ( .G(n22), .D(cbid[19]), .Q(\_zzLB[2][31] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][32] ( .G(n22), .D(idata[0]), .Q(\_zzLB[2][32] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][33] ( .G(n22), .D(idata[1]), .Q(\_zzLB[2][33] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][34] ( .G(n22), .D(idata[2]), .Q(\_zzLB[2][34] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][35] ( .G(n22), .D(idata[3]), .Q(\_zzLB[2][35] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][36] ( .G(n22), .D(idata[4]), .Q(\_zzLB[2][36] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][37] ( .G(n22), .D(idata[5]), .Q(\_zzLB[2][37] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][38] ( .G(n22), .D(idata[6]), .Q(\_zzLB[2][38] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][39] ( .G(n22), .D(idata[7]), .Q(\_zzLB[2][39] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][40] ( .G(n22), .D(idata[8]), .Q(\_zzLB[2][40] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][41] ( .G(n22), .D(idata[9]), .Q(\_zzLB[2][41] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][42] ( .G(n22), .D(idata[10]), .Q(\_zzLB[2][42] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][43] ( .G(n22), .D(idata[11]), .Q(\_zzLB[2][43] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][44] ( .G(n22), .D(idata[12]), .Q(\_zzLB[2][44] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][45] ( .G(n22), .D(idata[13]), .Q(\_zzLB[2][45] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][46] ( .G(n22), .D(idata[14]), .Q(\_zzLB[2][46] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][47] ( .G(n22), .D(idata[15]), .Q(\_zzLB[2][47] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][48] ( .G(n22), .D(idata[16]), .Q(\_zzLB[2][48] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][49] ( .G(n22), .D(idata[17]), .Q(\_zzLB[2][49] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][50] ( .G(n22), .D(idata[18]), .Q(\_zzLB[2][50] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][51] ( .G(n22), .D(idata[19]), .Q(\_zzLB[2][51] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][52] ( .G(n22), .D(idata[20]), .Q(\_zzLB[2][52] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][53] ( .G(n22), .D(idata[21]), .Q(\_zzLB[2][53] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][54] ( .G(n22), .D(idata[22]), .Q(\_zzLB[2][54] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][55] ( .G(n22), .D(idata[23]), .Q(\_zzLB[2][55] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][56] ( .G(n22), .D(idata[24]), .Q(\_zzLB[2][56] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][57] ( .G(n22), .D(idata[25]), .Q(\_zzLB[2][57] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][58] ( .G(n22), .D(idata[26]), .Q(\_zzLB[2][58] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][59] ( .G(n22), .D(idata[27]), .Q(\_zzLB[2][59] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][60] ( .G(n22), .D(idata[28]), .Q(\_zzLB[2][60] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][61] ( .G(n22), .D(idata[29]), .Q(\_zzLB[2][61] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][62] ( .G(n22), .D(idata[30]), .Q(\_zzLB[2][62] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][63] ( .G(n22), .D(idata[31]), .Q(\_zzLB[2][63] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][64] ( .G(n22), .D(idata[32]), .Q(\_zzLB[2][64] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][65] ( .G(n22), .D(idata[33]), .Q(\_zzLB[2][65] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][66] ( .G(n22), .D(idata[34]), .Q(\_zzLB[2][66] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][67] ( .G(n22), .D(idata[35]), .Q(\_zzLB[2][67] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][68] ( .G(n22), .D(idata[36]), .Q(\_zzLB[2][68] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][69] ( .G(n22), .D(idata[37]), .Q(\_zzLB[2][69] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][70] ( .G(n22), .D(idata[38]), .Q(\_zzLB[2][70] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][71] ( .G(n22), .D(idata[39]), .Q(\_zzLB[2][71] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][72] ( .G(n22), .D(idata[40]), .Q(\_zzLB[2][72] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][73] ( .G(n22), .D(idata[41]), .Q(\_zzLB[2][73] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][74] ( .G(n22), .D(idata[42]), .Q(\_zzLB[2][74] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][75] ( .G(n22), .D(idata[43]), .Q(\_zzLB[2][75] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][76] ( .G(n22), .D(idata[44]), .Q(\_zzLB[2][76] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][77] ( .G(n22), .D(idata[45]), .Q(\_zzLB[2][77] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][78] ( .G(n22), .D(idata[46]), .Q(\_zzLB[2][78] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][79] ( .G(n22), .D(idata[47]), .Q(\_zzLB[2][79] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][80] ( .G(n22), .D(idata[48]), .Q(\_zzLB[2][80] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][81] ( .G(n22), .D(idata[49]), .Q(\_zzLB[2][81] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][82] ( .G(n22), .D(idata[50]), .Q(\_zzLB[2][82] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][83] ( .G(n22), .D(idata[51]), .Q(\_zzLB[2][83] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][84] ( .G(n22), .D(idata[52]), .Q(\_zzLB[2][84] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][85] ( .G(n22), .D(idata[53]), .Q(\_zzLB[2][85] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][86] ( .G(n22), .D(idata[54]), .Q(\_zzLB[2][86] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][87] ( .G(n22), .D(idata[55]), .Q(\_zzLB[2][87] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][88] ( .G(n22), .D(idata[56]), .Q(\_zzLB[2][88] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][89] ( .G(n22), .D(idata[57]), .Q(\_zzLB[2][89] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][90] ( .G(n22), .D(idata[58]), .Q(\_zzLB[2][90] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][91] ( .G(n22), .D(idata[59]), .Q(\_zzLB[2][91] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][92] ( .G(n22), .D(idata[60]), .Q(\_zzLB[2][92] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][93] ( .G(n22), .D(idata[61]), .Q(\_zzLB[2][93] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][94] ( .G(n22), .D(idata[62]), .Q(\_zzLB[2][94] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][95] ( .G(n22), .D(idata[63]), .Q(\_zzLB[2][95] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][96] ( .G(n22), .D(idata[64]), .Q(\_zzLB[2][96] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][97] ( .G(n22), .D(idata[65]), .Q(\_zzLB[2][97] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][98] ( .G(n22), .D(idata[66]), .Q(\_zzLB[2][98] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][99] ( .G(n22), .D(idata[67]), .Q(\_zzLB[2][99] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][100] ( .G(n22), .D(idata[68]), .Q(\_zzLB[2][100] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][101] ( .G(n22), .D(idata[69]), .Q(\_zzLB[2][101] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][102] ( .G(n22), .D(idata[70]), .Q(\_zzLB[2][102] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][103] ( .G(n22), .D(idata[71]), .Q(\_zzLB[2][103] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][104] ( .G(n22), .D(idata[72]), .Q(\_zzLB[2][104] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][105] ( .G(n22), .D(idata[73]), .Q(\_zzLB[2][105] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][106] ( .G(n22), .D(idata[74]), .Q(\_zzLB[2][106] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][107] ( .G(n22), .D(idata[75]), .Q(\_zzLB[2][107] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][108] ( .G(n22), .D(idata[76]), .Q(\_zzLB[2][108] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][109] ( .G(n22), .D(idata[77]), .Q(\_zzLB[2][109] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][110] ( .G(n22), .D(idata[78]), .Q(\_zzLB[2][110] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][111] ( .G(n22), .D(idata[79]), .Q(\_zzLB[2][111] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][112] ( .G(n22), .D(idata[80]), .Q(\_zzLB[2][112] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][113] ( .G(n22), .D(idata[81]), .Q(\_zzLB[2][113] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][114] ( .G(n22), .D(idata[82]), .Q(\_zzLB[2][114] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][115] ( .G(n22), .D(idata[83]), .Q(\_zzLB[2][115] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][116] ( .G(n22), .D(idata[84]), .Q(\_zzLB[2][116] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][117] ( .G(n22), .D(idata[85]), .Q(\_zzLB[2][117] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][118] ( .G(n22), .D(idata[86]), .Q(\_zzLB[2][118] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][119] ( .G(n22), .D(idata[87]), .Q(\_zzLB[2][119] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][120] ( .G(n22), .D(idata[88]), .Q(\_zzLB[2][120] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][121] ( .G(n22), .D(idata[89]), .Q(\_zzLB[2][121] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][122] ( .G(n22), .D(idata[90]), .Q(\_zzLB[2][122] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][123] ( .G(n22), .D(idata[91]), .Q(\_zzLB[2][123] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][124] ( .G(n22), .D(idata[92]), .Q(\_zzLB[2][124] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][125] ( .G(n22), .D(idata[93]), .Q(\_zzLB[2][125] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][126] ( .G(n22), .D(idata[94]), .Q(\_zzLB[2][126] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][127] ( .G(n22), .D(idata[95]), .Q(\_zzLB[2][127] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][128] ( .G(n22), .D(ireq), .Q(\_zzLB[2][128] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][0] ( .G(n23), .D(len[0]), .Q(\_zzLB[3][0] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][1] ( .G(n23), .D(len[1]), .Q(\_zzLB[3][1] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][2] ( .G(n23), .D(len[2]), .Q(\_zzLB[3][2] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][3] ( .G(n23), .D(len[3]), .Q(\_zzLB[3][3] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][4] ( .G(n23), .D(len[4]), .Q(\_zzLB[3][4] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][5] ( .G(n23), .D(len[5]), .Q(\_zzLB[3][5] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][6] ( .G(n23), .D(len[6]), .Q(\_zzLB[3][6] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][7] ( .G(n23), .D(len[7]), .Q(\_zzLB[3][7] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][8] ( .G(n23), .D(len[8]), .Q(\_zzLB[3][8] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][9] ( .G(n23), .D(len[9]), .Q(\_zzLB[3][9] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][10] ( .G(n23), .D(len[10]), .Q(\_zzLB[3][10] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][11] ( .G(n23), .D(len[11]), .Q(\_zzLB[3][11] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][12] ( .G(n23), .D(cbid[0]), .Q(\_zzLB[3][12] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][13] ( .G(n23), .D(cbid[1]), .Q(\_zzLB[3][13] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][14] ( .G(n23), .D(cbid[2]), .Q(\_zzLB[3][14] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][15] ( .G(n23), .D(cbid[3]), .Q(\_zzLB[3][15] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][16] ( .G(n23), .D(cbid[4]), .Q(\_zzLB[3][16] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][17] ( .G(n23), .D(cbid[5]), .Q(\_zzLB[3][17] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][18] ( .G(n23), .D(cbid[6]), .Q(\_zzLB[3][18] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][19] ( .G(n23), .D(cbid[7]), .Q(\_zzLB[3][19] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][20] ( .G(n23), .D(cbid[8]), .Q(\_zzLB[3][20] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][21] ( .G(n23), .D(cbid[9]), .Q(\_zzLB[3][21] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][22] ( .G(n23), .D(cbid[10]), .Q(\_zzLB[3][22] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][23] ( .G(n23), .D(cbid[11]), .Q(\_zzLB[3][23] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][24] ( .G(n23), .D(cbid[12]), .Q(\_zzLB[3][24] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][25] ( .G(n23), .D(cbid[13]), .Q(\_zzLB[3][25] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][26] ( .G(n23), .D(cbid[14]), .Q(\_zzLB[3][26] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][27] ( .G(n23), .D(cbid[15]), .Q(\_zzLB[3][27] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][28] ( .G(n23), .D(cbid[16]), .Q(\_zzLB[3][28] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][29] ( .G(n23), .D(cbid[17]), .Q(\_zzLB[3][29] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][30] ( .G(n23), .D(cbid[18]), .Q(\_zzLB[3][30] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][31] ( .G(n23), .D(cbid[19]), .Q(\_zzLB[3][31] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][32] ( .G(n23), .D(idata[0]), .Q(\_zzLB[3][32] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][33] ( .G(n23), .D(idata[1]), .Q(\_zzLB[3][33] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][34] ( .G(n23), .D(idata[2]), .Q(\_zzLB[3][34] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][35] ( .G(n23), .D(idata[3]), .Q(\_zzLB[3][35] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][36] ( .G(n23), .D(idata[4]), .Q(\_zzLB[3][36] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][37] ( .G(n23), .D(idata[5]), .Q(\_zzLB[3][37] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][38] ( .G(n23), .D(idata[6]), .Q(\_zzLB[3][38] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][39] ( .G(n23), .D(idata[7]), .Q(\_zzLB[3][39] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][40] ( .G(n23), .D(idata[8]), .Q(\_zzLB[3][40] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][41] ( .G(n23), .D(idata[9]), .Q(\_zzLB[3][41] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][42] ( .G(n23), .D(idata[10]), .Q(\_zzLB[3][42] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][43] ( .G(n23), .D(idata[11]), .Q(\_zzLB[3][43] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][44] ( .G(n23), .D(idata[12]), .Q(\_zzLB[3][44] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][45] ( .G(n23), .D(idata[13]), .Q(\_zzLB[3][45] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][46] ( .G(n23), .D(idata[14]), .Q(\_zzLB[3][46] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][47] ( .G(n23), .D(idata[15]), .Q(\_zzLB[3][47] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][48] ( .G(n23), .D(idata[16]), .Q(\_zzLB[3][48] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][49] ( .G(n23), .D(idata[17]), .Q(\_zzLB[3][49] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][50] ( .G(n23), .D(idata[18]), .Q(\_zzLB[3][50] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][51] ( .G(n23), .D(idata[19]), .Q(\_zzLB[3][51] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][52] ( .G(n23), .D(idata[20]), .Q(\_zzLB[3][52] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][53] ( .G(n23), .D(idata[21]), .Q(\_zzLB[3][53] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][54] ( .G(n23), .D(idata[22]), .Q(\_zzLB[3][54] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][55] ( .G(n23), .D(idata[23]), .Q(\_zzLB[3][55] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][56] ( .G(n23), .D(idata[24]), .Q(\_zzLB[3][56] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][57] ( .G(n23), .D(idata[25]), .Q(\_zzLB[3][57] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][58] ( .G(n23), .D(idata[26]), .Q(\_zzLB[3][58] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][59] ( .G(n23), .D(idata[27]), .Q(\_zzLB[3][59] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][60] ( .G(n23), .D(idata[28]), .Q(\_zzLB[3][60] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][61] ( .G(n23), .D(idata[29]), .Q(\_zzLB[3][61] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][62] ( .G(n23), .D(idata[30]), .Q(\_zzLB[3][62] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][63] ( .G(n23), .D(idata[31]), .Q(\_zzLB[3][63] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][64] ( .G(n23), .D(idata[32]), .Q(\_zzLB[3][64] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][65] ( .G(n23), .D(idata[33]), .Q(\_zzLB[3][65] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][66] ( .G(n23), .D(idata[34]), .Q(\_zzLB[3][66] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][67] ( .G(n23), .D(idata[35]), .Q(\_zzLB[3][67] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][68] ( .G(n23), .D(idata[36]), .Q(\_zzLB[3][68] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][69] ( .G(n23), .D(idata[37]), .Q(\_zzLB[3][69] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][70] ( .G(n23), .D(idata[38]), .Q(\_zzLB[3][70] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][71] ( .G(n23), .D(idata[39]), .Q(\_zzLB[3][71] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][72] ( .G(n23), .D(idata[40]), .Q(\_zzLB[3][72] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][73] ( .G(n23), .D(idata[41]), .Q(\_zzLB[3][73] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][74] ( .G(n23), .D(idata[42]), .Q(\_zzLB[3][74] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][75] ( .G(n23), .D(idata[43]), .Q(\_zzLB[3][75] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][76] ( .G(n23), .D(idata[44]), .Q(\_zzLB[3][76] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][77] ( .G(n23), .D(idata[45]), .Q(\_zzLB[3][77] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][78] ( .G(n23), .D(idata[46]), .Q(\_zzLB[3][78] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][79] ( .G(n23), .D(idata[47]), .Q(\_zzLB[3][79] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][80] ( .G(n23), .D(idata[48]), .Q(\_zzLB[3][80] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][81] ( .G(n23), .D(idata[49]), .Q(\_zzLB[3][81] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][82] ( .G(n23), .D(idata[50]), .Q(\_zzLB[3][82] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][83] ( .G(n23), .D(idata[51]), .Q(\_zzLB[3][83] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][84] ( .G(n23), .D(idata[52]), .Q(\_zzLB[3][84] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][85] ( .G(n23), .D(idata[53]), .Q(\_zzLB[3][85] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][86] ( .G(n23), .D(idata[54]), .Q(\_zzLB[3][86] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][87] ( .G(n23), .D(idata[55]), .Q(\_zzLB[3][87] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][88] ( .G(n23), .D(idata[56]), .Q(\_zzLB[3][88] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][89] ( .G(n23), .D(idata[57]), .Q(\_zzLB[3][89] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][90] ( .G(n23), .D(idata[58]), .Q(\_zzLB[3][90] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][91] ( .G(n23), .D(idata[59]), .Q(\_zzLB[3][91] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][92] ( .G(n23), .D(idata[60]), .Q(\_zzLB[3][92] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][93] ( .G(n23), .D(idata[61]), .Q(\_zzLB[3][93] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][94] ( .G(n23), .D(idata[62]), .Q(\_zzLB[3][94] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][95] ( .G(n23), .D(idata[63]), .Q(\_zzLB[3][95] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][96] ( .G(n23), .D(idata[64]), .Q(\_zzLB[3][96] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][97] ( .G(n23), .D(idata[65]), .Q(\_zzLB[3][97] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][98] ( .G(n23), .D(idata[66]), .Q(\_zzLB[3][98] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][99] ( .G(n23), .D(idata[67]), .Q(\_zzLB[3][99] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][100] ( .G(n23), .D(idata[68]), .Q(\_zzLB[3][100] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][101] ( .G(n23), .D(idata[69]), .Q(\_zzLB[3][101] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][102] ( .G(n23), .D(idata[70]), .Q(\_zzLB[3][102] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][103] ( .G(n23), .D(idata[71]), .Q(\_zzLB[3][103] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][104] ( .G(n23), .D(idata[72]), .Q(\_zzLB[3][104] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][105] ( .G(n23), .D(idata[73]), .Q(\_zzLB[3][105] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][106] ( .G(n23), .D(idata[74]), .Q(\_zzLB[3][106] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][107] ( .G(n23), .D(idata[75]), .Q(\_zzLB[3][107] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][108] ( .G(n23), .D(idata[76]), .Q(\_zzLB[3][108] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][109] ( .G(n23), .D(idata[77]), .Q(\_zzLB[3][109] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][110] ( .G(n23), .D(idata[78]), .Q(\_zzLB[3][110] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][111] ( .G(n23), .D(idata[79]), .Q(\_zzLB[3][111] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][112] ( .G(n23), .D(idata[80]), .Q(\_zzLB[3][112] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][113] ( .G(n23), .D(idata[81]), .Q(\_zzLB[3][113] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][114] ( .G(n23), .D(idata[82]), .Q(\_zzLB[3][114] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][115] ( .G(n23), .D(idata[83]), .Q(\_zzLB[3][115] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][116] ( .G(n23), .D(idata[84]), .Q(\_zzLB[3][116] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][117] ( .G(n23), .D(idata[85]), .Q(\_zzLB[3][117] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][118] ( .G(n23), .D(idata[86]), .Q(\_zzLB[3][118] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][119] ( .G(n23), .D(idata[87]), .Q(\_zzLB[3][119] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][120] ( .G(n23), .D(idata[88]), .Q(\_zzLB[3][120] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][121] ( .G(n23), .D(idata[89]), .Q(\_zzLB[3][121] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][122] ( .G(n23), .D(idata[90]), .Q(\_zzLB[3][122] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][123] ( .G(n23), .D(idata[91]), .Q(\_zzLB[3][123] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][124] ( .G(n23), .D(idata[92]), .Q(\_zzLB[3][124] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][125] ( .G(n23), .D(idata[93]), .Q(\_zzLB[3][125] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][126] ( .G(n23), .D(idata[94]), .Q(\_zzLB[3][126] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][127] ( .G(n23), .D(idata[95]), .Q(\_zzLB[3][127] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][128] ( .G(n23), .D(ireq), .Q(\_zzLB[3][128] ), .QN( ));
Q_MX04 U811 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][0] ), .A1(\_zzLB[1][0] ), .A2(\_zzLB[2][0] ), .A3(\_zzLB[3][0] ), .Z(olen[0]));
Q_MX04 U812 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][1] ), .A1(\_zzLB[1][1] ), .A2(\_zzLB[2][1] ), .A3(\_zzLB[3][1] ), .Z(olen[1]));
Q_MX04 U813 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][2] ), .A1(\_zzLB[1][2] ), .A2(\_zzLB[2][2] ), .A3(\_zzLB[3][2] ), .Z(olen[2]));
Q_MX04 U814 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][3] ), .A1(\_zzLB[1][3] ), .A2(\_zzLB[2][3] ), .A3(\_zzLB[3][3] ), .Z(olen[3]));
Q_MX04 U815 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][4] ), .A1(\_zzLB[1][4] ), .A2(\_zzLB[2][4] ), .A3(\_zzLB[3][4] ), .Z(olen[4]));
Q_MX04 U816 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][5] ), .A1(\_zzLB[1][5] ), .A2(\_zzLB[2][5] ), .A3(\_zzLB[3][5] ), .Z(olen[5]));
Q_MX04 U817 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][6] ), .A1(\_zzLB[1][6] ), .A2(\_zzLB[2][6] ), .A3(\_zzLB[3][6] ), .Z(olen[6]));
Q_MX04 U818 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][7] ), .A1(\_zzLB[1][7] ), .A2(\_zzLB[2][7] ), .A3(\_zzLB[3][7] ), .Z(olen[7]));
Q_MX04 U819 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][8] ), .A1(\_zzLB[1][8] ), .A2(\_zzLB[2][8] ), .A3(\_zzLB[3][8] ), .Z(olen[8]));
Q_MX04 U820 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][9] ), .A1(\_zzLB[1][9] ), .A2(\_zzLB[2][9] ), .A3(\_zzLB[3][9] ), .Z(olen[9]));
Q_MX04 U821 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][10] ), .A1(\_zzLB[1][10] ), .A2(\_zzLB[2][10] ), .A3(\_zzLB[3][10] ), .Z(olen[10]));
Q_MX04 U822 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][11] ), .A1(\_zzLB[1][11] ), .A2(\_zzLB[2][11] ), .A3(\_zzLB[3][11] ), .Z(olen[11]));
Q_MX04 U823 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][12] ), .A1(\_zzLB[1][12] ), .A2(\_zzLB[2][12] ), .A3(\_zzLB[3][12] ), .Z(ocbid[0]));
Q_MX04 U824 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][13] ), .A1(\_zzLB[1][13] ), .A2(\_zzLB[2][13] ), .A3(\_zzLB[3][13] ), .Z(ocbid[1]));
Q_MX04 U825 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][14] ), .A1(\_zzLB[1][14] ), .A2(\_zzLB[2][14] ), .A3(\_zzLB[3][14] ), .Z(ocbid[2]));
Q_MX04 U826 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][15] ), .A1(\_zzLB[1][15] ), .A2(\_zzLB[2][15] ), .A3(\_zzLB[3][15] ), .Z(ocbid[3]));
Q_MX04 U827 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][16] ), .A1(\_zzLB[1][16] ), .A2(\_zzLB[2][16] ), .A3(\_zzLB[3][16] ), .Z(ocbid[4]));
Q_MX04 U828 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][17] ), .A1(\_zzLB[1][17] ), .A2(\_zzLB[2][17] ), .A3(\_zzLB[3][17] ), .Z(ocbid[5]));
Q_MX04 U829 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][18] ), .A1(\_zzLB[1][18] ), .A2(\_zzLB[2][18] ), .A3(\_zzLB[3][18] ), .Z(ocbid[6]));
Q_MX04 U830 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][19] ), .A1(\_zzLB[1][19] ), .A2(\_zzLB[2][19] ), .A3(\_zzLB[3][19] ), .Z(ocbid[7]));
Q_MX04 U831 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][20] ), .A1(\_zzLB[1][20] ), .A2(\_zzLB[2][20] ), .A3(\_zzLB[3][20] ), .Z(ocbid[8]));
Q_MX04 U832 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][21] ), .A1(\_zzLB[1][21] ), .A2(\_zzLB[2][21] ), .A3(\_zzLB[3][21] ), .Z(ocbid[9]));
Q_MX04 U833 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][22] ), .A1(\_zzLB[1][22] ), .A2(\_zzLB[2][22] ), .A3(\_zzLB[3][22] ), .Z(ocbid[10]));
Q_MX04 U834 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][23] ), .A1(\_zzLB[1][23] ), .A2(\_zzLB[2][23] ), .A3(\_zzLB[3][23] ), .Z(ocbid[11]));
Q_MX04 U835 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][24] ), .A1(\_zzLB[1][24] ), .A2(\_zzLB[2][24] ), .A3(\_zzLB[3][24] ), .Z(ocbid[12]));
Q_MX04 U836 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][25] ), .A1(\_zzLB[1][25] ), .A2(\_zzLB[2][25] ), .A3(\_zzLB[3][25] ), .Z(ocbid[13]));
Q_MX04 U837 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][26] ), .A1(\_zzLB[1][26] ), .A2(\_zzLB[2][26] ), .A3(\_zzLB[3][26] ), .Z(ocbid[14]));
Q_MX04 U838 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][27] ), .A1(\_zzLB[1][27] ), .A2(\_zzLB[2][27] ), .A3(\_zzLB[3][27] ), .Z(ocbid[15]));
Q_MX04 U839 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][28] ), .A1(\_zzLB[1][28] ), .A2(\_zzLB[2][28] ), .A3(\_zzLB[3][28] ), .Z(ocbid[16]));
Q_MX04 U840 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][29] ), .A1(\_zzLB[1][29] ), .A2(\_zzLB[2][29] ), .A3(\_zzLB[3][29] ), .Z(ocbid[17]));
Q_MX04 U841 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][30] ), .A1(\_zzLB[1][30] ), .A2(\_zzLB[2][30] ), .A3(\_zzLB[3][30] ), .Z(ocbid[18]));
Q_MX04 U842 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][31] ), .A1(\_zzLB[1][31] ), .A2(\_zzLB[2][31] ), .A3(\_zzLB[3][31] ), .Z(ocbid[19]));
Q_MX04 U843 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][32] ), .A1(\_zzLB[1][32] ), .A2(\_zzLB[2][32] ), .A3(\_zzLB[3][32] ), .Z(odata[0]));
Q_MX04 U844 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][33] ), .A1(\_zzLB[1][33] ), .A2(\_zzLB[2][33] ), .A3(\_zzLB[3][33] ), .Z(odata[1]));
Q_MX04 U845 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][34] ), .A1(\_zzLB[1][34] ), .A2(\_zzLB[2][34] ), .A3(\_zzLB[3][34] ), .Z(odata[2]));
Q_MX04 U846 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][35] ), .A1(\_zzLB[1][35] ), .A2(\_zzLB[2][35] ), .A3(\_zzLB[3][35] ), .Z(odata[3]));
Q_MX04 U847 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][36] ), .A1(\_zzLB[1][36] ), .A2(\_zzLB[2][36] ), .A3(\_zzLB[3][36] ), .Z(odata[4]));
Q_MX04 U848 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][37] ), .A1(\_zzLB[1][37] ), .A2(\_zzLB[2][37] ), .A3(\_zzLB[3][37] ), .Z(odata[5]));
Q_MX04 U849 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][38] ), .A1(\_zzLB[1][38] ), .A2(\_zzLB[2][38] ), .A3(\_zzLB[3][38] ), .Z(odata[6]));
Q_MX04 U850 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][39] ), .A1(\_zzLB[1][39] ), .A2(\_zzLB[2][39] ), .A3(\_zzLB[3][39] ), .Z(odata[7]));
Q_MX04 U851 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][40] ), .A1(\_zzLB[1][40] ), .A2(\_zzLB[2][40] ), .A3(\_zzLB[3][40] ), .Z(odata[8]));
Q_MX04 U852 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][41] ), .A1(\_zzLB[1][41] ), .A2(\_zzLB[2][41] ), .A3(\_zzLB[3][41] ), .Z(odata[9]));
Q_MX04 U853 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][42] ), .A1(\_zzLB[1][42] ), .A2(\_zzLB[2][42] ), .A3(\_zzLB[3][42] ), .Z(odata[10]));
Q_MX04 U854 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][43] ), .A1(\_zzLB[1][43] ), .A2(\_zzLB[2][43] ), .A3(\_zzLB[3][43] ), .Z(odata[11]));
Q_MX04 U855 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][44] ), .A1(\_zzLB[1][44] ), .A2(\_zzLB[2][44] ), .A3(\_zzLB[3][44] ), .Z(odata[12]));
Q_MX04 U856 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][45] ), .A1(\_zzLB[1][45] ), .A2(\_zzLB[2][45] ), .A3(\_zzLB[3][45] ), .Z(odata[13]));
Q_MX04 U857 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][46] ), .A1(\_zzLB[1][46] ), .A2(\_zzLB[2][46] ), .A3(\_zzLB[3][46] ), .Z(odata[14]));
Q_MX04 U858 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][47] ), .A1(\_zzLB[1][47] ), .A2(\_zzLB[2][47] ), .A3(\_zzLB[3][47] ), .Z(odata[15]));
Q_MX04 U859 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][48] ), .A1(\_zzLB[1][48] ), .A2(\_zzLB[2][48] ), .A3(\_zzLB[3][48] ), .Z(odata[16]));
Q_MX04 U860 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][49] ), .A1(\_zzLB[1][49] ), .A2(\_zzLB[2][49] ), .A3(\_zzLB[3][49] ), .Z(odata[17]));
Q_MX04 U861 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][50] ), .A1(\_zzLB[1][50] ), .A2(\_zzLB[2][50] ), .A3(\_zzLB[3][50] ), .Z(odata[18]));
Q_MX04 U862 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][51] ), .A1(\_zzLB[1][51] ), .A2(\_zzLB[2][51] ), .A3(\_zzLB[3][51] ), .Z(odata[19]));
Q_MX04 U863 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][52] ), .A1(\_zzLB[1][52] ), .A2(\_zzLB[2][52] ), .A3(\_zzLB[3][52] ), .Z(odata[20]));
Q_MX04 U864 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][53] ), .A1(\_zzLB[1][53] ), .A2(\_zzLB[2][53] ), .A3(\_zzLB[3][53] ), .Z(odata[21]));
Q_MX04 U865 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][54] ), .A1(\_zzLB[1][54] ), .A2(\_zzLB[2][54] ), .A3(\_zzLB[3][54] ), .Z(odata[22]));
Q_MX04 U866 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][55] ), .A1(\_zzLB[1][55] ), .A2(\_zzLB[2][55] ), .A3(\_zzLB[3][55] ), .Z(odata[23]));
Q_MX04 U867 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][56] ), .A1(\_zzLB[1][56] ), .A2(\_zzLB[2][56] ), .A3(\_zzLB[3][56] ), .Z(odata[24]));
Q_MX04 U868 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][57] ), .A1(\_zzLB[1][57] ), .A2(\_zzLB[2][57] ), .A3(\_zzLB[3][57] ), .Z(odata[25]));
Q_MX04 U869 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][58] ), .A1(\_zzLB[1][58] ), .A2(\_zzLB[2][58] ), .A3(\_zzLB[3][58] ), .Z(odata[26]));
Q_MX04 U870 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][59] ), .A1(\_zzLB[1][59] ), .A2(\_zzLB[2][59] ), .A3(\_zzLB[3][59] ), .Z(odata[27]));
Q_MX04 U871 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][60] ), .A1(\_zzLB[1][60] ), .A2(\_zzLB[2][60] ), .A3(\_zzLB[3][60] ), .Z(odata[28]));
Q_MX04 U872 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][61] ), .A1(\_zzLB[1][61] ), .A2(\_zzLB[2][61] ), .A3(\_zzLB[3][61] ), .Z(odata[29]));
Q_MX04 U873 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][62] ), .A1(\_zzLB[1][62] ), .A2(\_zzLB[2][62] ), .A3(\_zzLB[3][62] ), .Z(odata[30]));
Q_MX04 U874 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][63] ), .A1(\_zzLB[1][63] ), .A2(\_zzLB[2][63] ), .A3(\_zzLB[3][63] ), .Z(odata[31]));
Q_MX04 U875 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][64] ), .A1(\_zzLB[1][64] ), .A2(\_zzLB[2][64] ), .A3(\_zzLB[3][64] ), .Z(odata[32]));
Q_MX04 U876 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][65] ), .A1(\_zzLB[1][65] ), .A2(\_zzLB[2][65] ), .A3(\_zzLB[3][65] ), .Z(odata[33]));
Q_MX04 U877 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][66] ), .A1(\_zzLB[1][66] ), .A2(\_zzLB[2][66] ), .A3(\_zzLB[3][66] ), .Z(odata[34]));
Q_MX04 U878 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][67] ), .A1(\_zzLB[1][67] ), .A2(\_zzLB[2][67] ), .A3(\_zzLB[3][67] ), .Z(odata[35]));
Q_MX04 U879 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][68] ), .A1(\_zzLB[1][68] ), .A2(\_zzLB[2][68] ), .A3(\_zzLB[3][68] ), .Z(odata[36]));
Q_MX04 U880 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][69] ), .A1(\_zzLB[1][69] ), .A2(\_zzLB[2][69] ), .A3(\_zzLB[3][69] ), .Z(odata[37]));
Q_MX04 U881 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][70] ), .A1(\_zzLB[1][70] ), .A2(\_zzLB[2][70] ), .A3(\_zzLB[3][70] ), .Z(odata[38]));
Q_MX04 U882 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][71] ), .A1(\_zzLB[1][71] ), .A2(\_zzLB[2][71] ), .A3(\_zzLB[3][71] ), .Z(odata[39]));
Q_MX04 U883 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][72] ), .A1(\_zzLB[1][72] ), .A2(\_zzLB[2][72] ), .A3(\_zzLB[3][72] ), .Z(odata[40]));
Q_MX04 U884 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][73] ), .A1(\_zzLB[1][73] ), .A2(\_zzLB[2][73] ), .A3(\_zzLB[3][73] ), .Z(odata[41]));
Q_MX04 U885 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][74] ), .A1(\_zzLB[1][74] ), .A2(\_zzLB[2][74] ), .A3(\_zzLB[3][74] ), .Z(odata[42]));
Q_MX04 U886 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][75] ), .A1(\_zzLB[1][75] ), .A2(\_zzLB[2][75] ), .A3(\_zzLB[3][75] ), .Z(odata[43]));
Q_MX04 U887 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][76] ), .A1(\_zzLB[1][76] ), .A2(\_zzLB[2][76] ), .A3(\_zzLB[3][76] ), .Z(odata[44]));
Q_MX04 U888 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][77] ), .A1(\_zzLB[1][77] ), .A2(\_zzLB[2][77] ), .A3(\_zzLB[3][77] ), .Z(odata[45]));
Q_MX04 U889 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][78] ), .A1(\_zzLB[1][78] ), .A2(\_zzLB[2][78] ), .A3(\_zzLB[3][78] ), .Z(odata[46]));
Q_MX04 U890 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][79] ), .A1(\_zzLB[1][79] ), .A2(\_zzLB[2][79] ), .A3(\_zzLB[3][79] ), .Z(odata[47]));
Q_MX04 U891 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][80] ), .A1(\_zzLB[1][80] ), .A2(\_zzLB[2][80] ), .A3(\_zzLB[3][80] ), .Z(odata[48]));
Q_MX04 U892 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][81] ), .A1(\_zzLB[1][81] ), .A2(\_zzLB[2][81] ), .A3(\_zzLB[3][81] ), .Z(odata[49]));
Q_MX04 U893 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][82] ), .A1(\_zzLB[1][82] ), .A2(\_zzLB[2][82] ), .A3(\_zzLB[3][82] ), .Z(odata[50]));
Q_MX04 U894 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][83] ), .A1(\_zzLB[1][83] ), .A2(\_zzLB[2][83] ), .A3(\_zzLB[3][83] ), .Z(odata[51]));
Q_MX04 U895 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][84] ), .A1(\_zzLB[1][84] ), .A2(\_zzLB[2][84] ), .A3(\_zzLB[3][84] ), .Z(odata[52]));
Q_MX04 U896 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][85] ), .A1(\_zzLB[1][85] ), .A2(\_zzLB[2][85] ), .A3(\_zzLB[3][85] ), .Z(odata[53]));
Q_MX04 U897 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][86] ), .A1(\_zzLB[1][86] ), .A2(\_zzLB[2][86] ), .A3(\_zzLB[3][86] ), .Z(odata[54]));
Q_MX04 U898 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][87] ), .A1(\_zzLB[1][87] ), .A2(\_zzLB[2][87] ), .A3(\_zzLB[3][87] ), .Z(odata[55]));
Q_MX04 U899 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][88] ), .A1(\_zzLB[1][88] ), .A2(\_zzLB[2][88] ), .A3(\_zzLB[3][88] ), .Z(odata[56]));
Q_MX04 U900 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][89] ), .A1(\_zzLB[1][89] ), .A2(\_zzLB[2][89] ), .A3(\_zzLB[3][89] ), .Z(odata[57]));
Q_MX04 U901 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][90] ), .A1(\_zzLB[1][90] ), .A2(\_zzLB[2][90] ), .A3(\_zzLB[3][90] ), .Z(odata[58]));
Q_MX04 U902 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][91] ), .A1(\_zzLB[1][91] ), .A2(\_zzLB[2][91] ), .A3(\_zzLB[3][91] ), .Z(odata[59]));
Q_MX04 U903 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][92] ), .A1(\_zzLB[1][92] ), .A2(\_zzLB[2][92] ), .A3(\_zzLB[3][92] ), .Z(odata[60]));
Q_MX04 U904 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][93] ), .A1(\_zzLB[1][93] ), .A2(\_zzLB[2][93] ), .A3(\_zzLB[3][93] ), .Z(odata[61]));
Q_MX04 U905 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][94] ), .A1(\_zzLB[1][94] ), .A2(\_zzLB[2][94] ), .A3(\_zzLB[3][94] ), .Z(odata[62]));
Q_MX04 U906 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][95] ), .A1(\_zzLB[1][95] ), .A2(\_zzLB[2][95] ), .A3(\_zzLB[3][95] ), .Z(odata[63]));
Q_MX04 U907 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][96] ), .A1(\_zzLB[1][96] ), .A2(\_zzLB[2][96] ), .A3(\_zzLB[3][96] ), .Z(odata[64]));
Q_MX04 U908 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][97] ), .A1(\_zzLB[1][97] ), .A2(\_zzLB[2][97] ), .A3(\_zzLB[3][97] ), .Z(odata[65]));
Q_MX04 U909 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][98] ), .A1(\_zzLB[1][98] ), .A2(\_zzLB[2][98] ), .A3(\_zzLB[3][98] ), .Z(odata[66]));
Q_MX04 U910 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][99] ), .A1(\_zzLB[1][99] ), .A2(\_zzLB[2][99] ), .A3(\_zzLB[3][99] ), .Z(odata[67]));
Q_MX04 U911 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][100] ), .A1(\_zzLB[1][100] ), .A2(\_zzLB[2][100] ), .A3(\_zzLB[3][100] ), .Z(odata[68]));
Q_MX04 U912 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][101] ), .A1(\_zzLB[1][101] ), .A2(\_zzLB[2][101] ), .A3(\_zzLB[3][101] ), .Z(odata[69]));
Q_MX04 U913 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][102] ), .A1(\_zzLB[1][102] ), .A2(\_zzLB[2][102] ), .A3(\_zzLB[3][102] ), .Z(odata[70]));
Q_MX04 U914 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][103] ), .A1(\_zzLB[1][103] ), .A2(\_zzLB[2][103] ), .A3(\_zzLB[3][103] ), .Z(odata[71]));
Q_MX04 U915 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][104] ), .A1(\_zzLB[1][104] ), .A2(\_zzLB[2][104] ), .A3(\_zzLB[3][104] ), .Z(odata[72]));
Q_MX04 U916 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][105] ), .A1(\_zzLB[1][105] ), .A2(\_zzLB[2][105] ), .A3(\_zzLB[3][105] ), .Z(odata[73]));
Q_MX04 U917 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][106] ), .A1(\_zzLB[1][106] ), .A2(\_zzLB[2][106] ), .A3(\_zzLB[3][106] ), .Z(odata[74]));
Q_MX04 U918 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][107] ), .A1(\_zzLB[1][107] ), .A2(\_zzLB[2][107] ), .A3(\_zzLB[3][107] ), .Z(odata[75]));
Q_MX04 U919 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][108] ), .A1(\_zzLB[1][108] ), .A2(\_zzLB[2][108] ), .A3(\_zzLB[3][108] ), .Z(odata[76]));
Q_MX04 U920 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][109] ), .A1(\_zzLB[1][109] ), .A2(\_zzLB[2][109] ), .A3(\_zzLB[3][109] ), .Z(odata[77]));
Q_MX04 U921 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][110] ), .A1(\_zzLB[1][110] ), .A2(\_zzLB[2][110] ), .A3(\_zzLB[3][110] ), .Z(odata[78]));
Q_MX04 U922 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][111] ), .A1(\_zzLB[1][111] ), .A2(\_zzLB[2][111] ), .A3(\_zzLB[3][111] ), .Z(odata[79]));
Q_MX04 U923 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][112] ), .A1(\_zzLB[1][112] ), .A2(\_zzLB[2][112] ), .A3(\_zzLB[3][112] ), .Z(odata[80]));
Q_MX04 U924 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][113] ), .A1(\_zzLB[1][113] ), .A2(\_zzLB[2][113] ), .A3(\_zzLB[3][113] ), .Z(odata[81]));
Q_MX04 U925 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][114] ), .A1(\_zzLB[1][114] ), .A2(\_zzLB[2][114] ), .A3(\_zzLB[3][114] ), .Z(odata[82]));
Q_MX04 U926 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][115] ), .A1(\_zzLB[1][115] ), .A2(\_zzLB[2][115] ), .A3(\_zzLB[3][115] ), .Z(odata[83]));
Q_MX04 U927 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][116] ), .A1(\_zzLB[1][116] ), .A2(\_zzLB[2][116] ), .A3(\_zzLB[3][116] ), .Z(odata[84]));
Q_MX04 U928 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][117] ), .A1(\_zzLB[1][117] ), .A2(\_zzLB[2][117] ), .A3(\_zzLB[3][117] ), .Z(odata[85]));
Q_MX04 U929 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][118] ), .A1(\_zzLB[1][118] ), .A2(\_zzLB[2][118] ), .A3(\_zzLB[3][118] ), .Z(odata[86]));
Q_MX04 U930 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][119] ), .A1(\_zzLB[1][119] ), .A2(\_zzLB[2][119] ), .A3(\_zzLB[3][119] ), .Z(odata[87]));
Q_MX04 U931 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][120] ), .A1(\_zzLB[1][120] ), .A2(\_zzLB[2][120] ), .A3(\_zzLB[3][120] ), .Z(odata[88]));
Q_MX04 U932 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][121] ), .A1(\_zzLB[1][121] ), .A2(\_zzLB[2][121] ), .A3(\_zzLB[3][121] ), .Z(odata[89]));
Q_MX04 U933 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][122] ), .A1(\_zzLB[1][122] ), .A2(\_zzLB[2][122] ), .A3(\_zzLB[3][122] ), .Z(odata[90]));
Q_MX04 U934 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][123] ), .A1(\_zzLB[1][123] ), .A2(\_zzLB[2][123] ), .A3(\_zzLB[3][123] ), .Z(odata[91]));
Q_MX04 U935 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][124] ), .A1(\_zzLB[1][124] ), .A2(\_zzLB[2][124] ), .A3(\_zzLB[3][124] ), .Z(odata[92]));
Q_MX04 U936 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][125] ), .A1(\_zzLB[1][125] ), .A2(\_zzLB[2][125] ), .A3(\_zzLB[3][125] ), .Z(odata[93]));
Q_MX04 U937 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][126] ), .A1(\_zzLB[1][126] ), .A2(\_zzLB[2][126] ), .A3(\_zzLB[3][126] ), .Z(odata[94]));
Q_MX04 U938 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][127] ), .A1(\_zzLB[1][127] ), .A2(\_zzLB[2][127] ), .A3(\_zzLB[3][127] ), .Z(odata[95]));
Q_MX04 U939 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][128] ), .A1(\_zzLB[1][128] ), .A2(\_zzLB[2][128] ), .A3(\_zzLB[3][128] ), .Z(oreq));
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m1 "_zzLB 1 128 0 0 3"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_NON_CMM "1"
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE "ixc_gfifo_port"
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE_LIB "IXCOM_TEMP_LIBRARY"
// pragma CVASTRPROP MODULE HDLICE PROP_IXCOM_MOD TRUE
endmodule
