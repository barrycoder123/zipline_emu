
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
`_2_ (* upf_always_on = 1 *) 
module ixcEcmHold ;
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
wire fclk;
wire uclk;
`_2_ wire holdEcm;
`_2_ wire hc;
`_2_ wire hs;
`_2_ wire [63:0] ecmTs;
`_2_ wire [63:0] ecmTsP;
`_2_ wire [255:0] ctrlR;
`_2_ wire [255:0] ctrlW;
`_2_ wire [1:0] ctrlEv;
`_2_ wire [1:0] ctrlEvP;
`_2_ wire newCtrl;
`_2_ wire [7:0] cmdC;
`_2_ wire [7:0] cmdR;
`_2_ wire [7:0] cmdCnt;
`_2_ wire [7:0] cmdCntP;
`_2_ wire [63:0] argTc;
`_2_ wire [63:0] argTs;
`_2_ wire [63:0] cRet;
`_2_ wire newCmd;
`_2_ wire busyOn;
`_2_ wire [7:0] busyCnt;
`_2_ wire [7:0] syncId;
`_2_ wire [7:0] syncIdP;
`_2_ wire newSync;
`_2_ wire [3:0] holdEcmD;
`_2_ wire holdEcmBusy;
`_2_ wire sdlStopRply;
`_2_ wire [63:0] simTime;
wire [0:0] _zyL692_meState0;
wire [0:0] _zyL739_meState1;
supply1 n337;
supply0 n594;
Q_BUF U0 ( .A(cRet[0]), .Z(ctrlW[0]));
Q_BUF U1 ( .A(cRet[1]), .Z(ctrlW[1]));
Q_BUF U2 ( .A(cRet[2]), .Z(ctrlW[2]));
Q_BUF U3 ( .A(cRet[3]), .Z(ctrlW[3]));
Q_ASSIGN U4 ( .B(cRet[4]), .A(ctrlW[4]));
Q_ASSIGN U5 ( .B(cRet[5]), .A(ctrlW[5]));
Q_ASSIGN U6 ( .B(cRet[6]), .A(ctrlW[6]));
Q_ASSIGN U7 ( .B(cRet[7]), .A(ctrlW[7]));
Q_BUF U8 ( .A(cRet[8]), .Z(ctrlW[8]));
Q_BUF U9 ( .A(cRet[9]), .Z(ctrlW[9]));
Q_BUF U10 ( .A(cRet[10]), .Z(ctrlW[10]));
Q_BUF U11 ( .A(cRet[11]), .Z(ctrlW[11]));
Q_BUF U12 ( .A(cRet[12]), .Z(ctrlW[12]));
Q_BUF U13 ( .A(cRet[13]), .Z(ctrlW[13]));
Q_BUF U14 ( .A(cRet[14]), .Z(ctrlW[14]));
Q_BUF U15 ( .A(cRet[15]), .Z(ctrlW[15]));
Q_ASSIGN U16 ( .B(cRet[16]), .A(ctrlW[16]));
Q_ASSIGN U17 ( .B(cRet[17]), .A(ctrlW[17]));
Q_ASSIGN U18 ( .B(cRet[18]), .A(ctrlW[18]));
Q_ASSIGN U19 ( .B(cRet[19]), .A(ctrlW[19]));
Q_ASSIGN U20 ( .B(cRet[20]), .A(ctrlW[20]));
Q_ASSIGN U21 ( .B(cRet[21]), .A(ctrlW[21]));
Q_ASSIGN U22 ( .B(cRet[22]), .A(ctrlW[22]));
Q_ASSIGN U23 ( .B(cRet[23]), .A(ctrlW[23]));
Q_ASSIGN U24 ( .B(cRet[24]), .A(ctrlW[24]));
Q_ASSIGN U25 ( .B(cRet[25]), .A(ctrlW[25]));
Q_ASSIGN U26 ( .B(cRet[26]), .A(ctrlW[26]));
Q_ASSIGN U27 ( .B(cRet[27]), .A(ctrlW[27]));
Q_ASSIGN U28 ( .B(cRet[28]), .A(ctrlW[28]));
Q_ASSIGN U29 ( .B(cRet[29]), .A(ctrlW[29]));
Q_ASSIGN U30 ( .B(cRet[30]), .A(ctrlW[30]));
Q_ASSIGN U31 ( .B(cRet[31]), .A(ctrlW[31]));
Q_ASSIGN U32 ( .B(cRet[32]), .A(ctrlW[32]));
Q_ASSIGN U33 ( .B(cRet[33]), .A(ctrlW[33]));
Q_ASSIGN U34 ( .B(cRet[34]), .A(ctrlW[34]));
Q_ASSIGN U35 ( .B(cRet[35]), .A(ctrlW[35]));
Q_ASSIGN U36 ( .B(cRet[36]), .A(ctrlW[36]));
Q_ASSIGN U37 ( .B(cRet[37]), .A(ctrlW[37]));
Q_ASSIGN U38 ( .B(cRet[38]), .A(ctrlW[38]));
Q_ASSIGN U39 ( .B(cRet[39]), .A(ctrlW[39]));
Q_ASSIGN U40 ( .B(cRet[40]), .A(ctrlW[40]));
Q_ASSIGN U41 ( .B(cRet[41]), .A(ctrlW[41]));
Q_ASSIGN U42 ( .B(cRet[42]), .A(ctrlW[42]));
Q_ASSIGN U43 ( .B(cRet[43]), .A(ctrlW[43]));
Q_ASSIGN U44 ( .B(cRet[44]), .A(ctrlW[44]));
Q_ASSIGN U45 ( .B(cRet[45]), .A(ctrlW[45]));
Q_ASSIGN U46 ( .B(cRet[46]), .A(ctrlW[46]));
Q_ASSIGN U47 ( .B(cRet[47]), .A(ctrlW[47]));
Q_ASSIGN U48 ( .B(cRet[48]), .A(ctrlW[48]));
Q_ASSIGN U49 ( .B(cRet[49]), .A(ctrlW[49]));
Q_ASSIGN U50 ( .B(cRet[50]), .A(ctrlW[50]));
Q_ASSIGN U51 ( .B(cRet[51]), .A(ctrlW[51]));
Q_ASSIGN U52 ( .B(cRet[52]), .A(ctrlW[52]));
Q_ASSIGN U53 ( .B(cRet[53]), .A(ctrlW[53]));
Q_ASSIGN U54 ( .B(cRet[54]), .A(ctrlW[54]));
Q_ASSIGN U55 ( .B(cRet[55]), .A(ctrlW[55]));
Q_ASSIGN U56 ( .B(cRet[56]), .A(ctrlW[56]));
Q_ASSIGN U57 ( .B(cRet[57]), .A(ctrlW[57]));
Q_ASSIGN U58 ( .B(cRet[58]), .A(ctrlW[58]));
Q_ASSIGN U59 ( .B(cRet[59]), .A(ctrlW[59]));
Q_ASSIGN U60 ( .B(cRet[60]), .A(ctrlW[60]));
Q_ASSIGN U61 ( .B(cRet[61]), .A(ctrlW[61]));
Q_ASSIGN U62 ( .B(cRet[62]), .A(ctrlW[62]));
Q_ASSIGN U63 ( .B(cRet[63]), .A(ctrlW[63]));
Q_ASSIGN U64 ( .B(xcva_top.xc_top.simTime[0]), .A(ctrlW[128]));
Q_ASSIGN U65 ( .B(xcva_top.xc_top.simTime[0]), .A(simTime[0]));
Q_ASSIGN U66 ( .B(xcva_top.xc_top.simTime[1]), .A(ctrlW[129]));
Q_ASSIGN U67 ( .B(xcva_top.xc_top.simTime[1]), .A(simTime[1]));
Q_ASSIGN U68 ( .B(xcva_top.xc_top.simTime[2]), .A(ctrlW[130]));
Q_ASSIGN U69 ( .B(xcva_top.xc_top.simTime[2]), .A(simTime[2]));
Q_ASSIGN U70 ( .B(xcva_top.xc_top.simTime[3]), .A(ctrlW[131]));
Q_ASSIGN U71 ( .B(xcva_top.xc_top.simTime[3]), .A(simTime[3]));
Q_ASSIGN U72 ( .B(xcva_top.xc_top.simTime[4]), .A(ctrlW[132]));
Q_ASSIGN U73 ( .B(xcva_top.xc_top.simTime[4]), .A(simTime[4]));
Q_ASSIGN U74 ( .B(xcva_top.xc_top.simTime[5]), .A(ctrlW[133]));
Q_ASSIGN U75 ( .B(xcva_top.xc_top.simTime[5]), .A(simTime[5]));
Q_ASSIGN U76 ( .B(xcva_top.xc_top.simTime[6]), .A(ctrlW[134]));
Q_ASSIGN U77 ( .B(xcva_top.xc_top.simTime[6]), .A(simTime[6]));
Q_ASSIGN U78 ( .B(xcva_top.xc_top.simTime[7]), .A(ctrlW[135]));
Q_ASSIGN U79 ( .B(xcva_top.xc_top.simTime[7]), .A(simTime[7]));
Q_ASSIGN U80 ( .B(xcva_top.xc_top.simTime[8]), .A(ctrlW[136]));
Q_ASSIGN U81 ( .B(xcva_top.xc_top.simTime[8]), .A(simTime[8]));
Q_ASSIGN U82 ( .B(xcva_top.xc_top.simTime[9]), .A(ctrlW[137]));
Q_ASSIGN U83 ( .B(xcva_top.xc_top.simTime[9]), .A(simTime[9]));
Q_ASSIGN U84 ( .B(xcva_top.xc_top.simTime[10]), .A(ctrlW[138]));
Q_ASSIGN U85 ( .B(xcva_top.xc_top.simTime[10]), .A(simTime[10]));
Q_ASSIGN U86 ( .B(xcva_top.xc_top.simTime[11]), .A(ctrlW[139]));
Q_ASSIGN U87 ( .B(xcva_top.xc_top.simTime[11]), .A(simTime[11]));
Q_ASSIGN U88 ( .B(xcva_top.xc_top.simTime[12]), .A(ctrlW[140]));
Q_ASSIGN U89 ( .B(xcva_top.xc_top.simTime[12]), .A(simTime[12]));
Q_ASSIGN U90 ( .B(xcva_top.xc_top.simTime[13]), .A(ctrlW[141]));
Q_ASSIGN U91 ( .B(xcva_top.xc_top.simTime[13]), .A(simTime[13]));
Q_ASSIGN U92 ( .B(xcva_top.xc_top.simTime[14]), .A(ctrlW[142]));
Q_ASSIGN U93 ( .B(xcva_top.xc_top.simTime[14]), .A(simTime[14]));
Q_ASSIGN U94 ( .B(xcva_top.xc_top.simTime[15]), .A(ctrlW[143]));
Q_ASSIGN U95 ( .B(xcva_top.xc_top.simTime[15]), .A(simTime[15]));
Q_ASSIGN U96 ( .B(xcva_top.xc_top.simTime[16]), .A(ctrlW[144]));
Q_ASSIGN U97 ( .B(xcva_top.xc_top.simTime[16]), .A(simTime[16]));
Q_ASSIGN U98 ( .B(xcva_top.xc_top.simTime[17]), .A(ctrlW[145]));
Q_ASSIGN U99 ( .B(xcva_top.xc_top.simTime[17]), .A(simTime[17]));
Q_ASSIGN U100 ( .B(xcva_top.xc_top.simTime[18]), .A(ctrlW[146]));
Q_ASSIGN U101 ( .B(xcva_top.xc_top.simTime[18]), .A(simTime[18]));
Q_ASSIGN U102 ( .B(xcva_top.xc_top.simTime[19]), .A(ctrlW[147]));
Q_ASSIGN U103 ( .B(xcva_top.xc_top.simTime[19]), .A(simTime[19]));
Q_ASSIGN U104 ( .B(xcva_top.xc_top.simTime[20]), .A(ctrlW[148]));
Q_ASSIGN U105 ( .B(xcva_top.xc_top.simTime[20]), .A(simTime[20]));
Q_ASSIGN U106 ( .B(xcva_top.xc_top.simTime[21]), .A(ctrlW[149]));
Q_ASSIGN U107 ( .B(xcva_top.xc_top.simTime[21]), .A(simTime[21]));
Q_ASSIGN U108 ( .B(xcva_top.xc_top.simTime[22]), .A(ctrlW[150]));
Q_ASSIGN U109 ( .B(xcva_top.xc_top.simTime[22]), .A(simTime[22]));
Q_ASSIGN U110 ( .B(xcva_top.xc_top.simTime[23]), .A(ctrlW[151]));
Q_ASSIGN U111 ( .B(xcva_top.xc_top.simTime[23]), .A(simTime[23]));
Q_ASSIGN U112 ( .B(xcva_top.xc_top.simTime[24]), .A(ctrlW[152]));
Q_ASSIGN U113 ( .B(xcva_top.xc_top.simTime[24]), .A(simTime[24]));
Q_ASSIGN U114 ( .B(xcva_top.xc_top.simTime[25]), .A(ctrlW[153]));
Q_ASSIGN U115 ( .B(xcva_top.xc_top.simTime[25]), .A(simTime[25]));
Q_ASSIGN U116 ( .B(xcva_top.xc_top.simTime[26]), .A(ctrlW[154]));
Q_ASSIGN U117 ( .B(xcva_top.xc_top.simTime[26]), .A(simTime[26]));
Q_ASSIGN U118 ( .B(xcva_top.xc_top.simTime[27]), .A(ctrlW[155]));
Q_ASSIGN U119 ( .B(xcva_top.xc_top.simTime[27]), .A(simTime[27]));
Q_ASSIGN U120 ( .B(xcva_top.xc_top.simTime[28]), .A(ctrlW[156]));
Q_ASSIGN U121 ( .B(xcva_top.xc_top.simTime[28]), .A(simTime[28]));
Q_ASSIGN U122 ( .B(xcva_top.xc_top.simTime[29]), .A(ctrlW[157]));
Q_ASSIGN U123 ( .B(xcva_top.xc_top.simTime[29]), .A(simTime[29]));
Q_ASSIGN U124 ( .B(xcva_top.xc_top.simTime[30]), .A(ctrlW[158]));
Q_ASSIGN U125 ( .B(xcva_top.xc_top.simTime[30]), .A(simTime[30]));
Q_ASSIGN U126 ( .B(xcva_top.xc_top.simTime[31]), .A(ctrlW[159]));
Q_ASSIGN U127 ( .B(xcva_top.xc_top.simTime[31]), .A(simTime[31]));
Q_ASSIGN U128 ( .B(xcva_top.xc_top.simTime[32]), .A(ctrlW[160]));
Q_ASSIGN U129 ( .B(xcva_top.xc_top.simTime[32]), .A(simTime[32]));
Q_ASSIGN U130 ( .B(xcva_top.xc_top.simTime[33]), .A(ctrlW[161]));
Q_ASSIGN U131 ( .B(xcva_top.xc_top.simTime[33]), .A(simTime[33]));
Q_ASSIGN U132 ( .B(xcva_top.xc_top.simTime[34]), .A(ctrlW[162]));
Q_ASSIGN U133 ( .B(xcva_top.xc_top.simTime[34]), .A(simTime[34]));
Q_ASSIGN U134 ( .B(xcva_top.xc_top.simTime[35]), .A(ctrlW[163]));
Q_ASSIGN U135 ( .B(xcva_top.xc_top.simTime[35]), .A(simTime[35]));
Q_ASSIGN U136 ( .B(xcva_top.xc_top.simTime[36]), .A(ctrlW[164]));
Q_ASSIGN U137 ( .B(xcva_top.xc_top.simTime[36]), .A(simTime[36]));
Q_ASSIGN U138 ( .B(xcva_top.xc_top.simTime[37]), .A(ctrlW[165]));
Q_ASSIGN U139 ( .B(xcva_top.xc_top.simTime[37]), .A(simTime[37]));
Q_ASSIGN U140 ( .B(xcva_top.xc_top.simTime[38]), .A(ctrlW[166]));
Q_ASSIGN U141 ( .B(xcva_top.xc_top.simTime[38]), .A(simTime[38]));
Q_ASSIGN U142 ( .B(xcva_top.xc_top.simTime[39]), .A(ctrlW[167]));
Q_ASSIGN U143 ( .B(xcva_top.xc_top.simTime[39]), .A(simTime[39]));
Q_ASSIGN U144 ( .B(xcva_top.xc_top.simTime[40]), .A(ctrlW[168]));
Q_ASSIGN U145 ( .B(xcva_top.xc_top.simTime[40]), .A(simTime[40]));
Q_ASSIGN U146 ( .B(xcva_top.xc_top.simTime[41]), .A(ctrlW[169]));
Q_ASSIGN U147 ( .B(xcva_top.xc_top.simTime[41]), .A(simTime[41]));
Q_ASSIGN U148 ( .B(xcva_top.xc_top.simTime[42]), .A(ctrlW[170]));
Q_ASSIGN U149 ( .B(xcva_top.xc_top.simTime[42]), .A(simTime[42]));
Q_ASSIGN U150 ( .B(xcva_top.xc_top.simTime[43]), .A(ctrlW[171]));
Q_ASSIGN U151 ( .B(xcva_top.xc_top.simTime[43]), .A(simTime[43]));
Q_ASSIGN U152 ( .B(xcva_top.xc_top.simTime[44]), .A(ctrlW[172]));
Q_ASSIGN U153 ( .B(xcva_top.xc_top.simTime[44]), .A(simTime[44]));
Q_ASSIGN U154 ( .B(xcva_top.xc_top.simTime[45]), .A(ctrlW[173]));
Q_ASSIGN U155 ( .B(xcva_top.xc_top.simTime[45]), .A(simTime[45]));
Q_ASSIGN U156 ( .B(xcva_top.xc_top.simTime[46]), .A(ctrlW[174]));
Q_ASSIGN U157 ( .B(xcva_top.xc_top.simTime[46]), .A(simTime[46]));
Q_ASSIGN U158 ( .B(xcva_top.xc_top.simTime[47]), .A(ctrlW[175]));
Q_ASSIGN U159 ( .B(xcva_top.xc_top.simTime[47]), .A(simTime[47]));
Q_ASSIGN U160 ( .B(xcva_top.xc_top.simTime[48]), .A(ctrlW[176]));
Q_ASSIGN U161 ( .B(xcva_top.xc_top.simTime[48]), .A(simTime[48]));
Q_ASSIGN U162 ( .B(xcva_top.xc_top.simTime[49]), .A(ctrlW[177]));
Q_ASSIGN U163 ( .B(xcva_top.xc_top.simTime[49]), .A(simTime[49]));
Q_ASSIGN U164 ( .B(xcva_top.xc_top.simTime[50]), .A(ctrlW[178]));
Q_ASSIGN U165 ( .B(xcva_top.xc_top.simTime[50]), .A(simTime[50]));
Q_ASSIGN U166 ( .B(xcva_top.xc_top.simTime[51]), .A(ctrlW[179]));
Q_ASSIGN U167 ( .B(xcva_top.xc_top.simTime[51]), .A(simTime[51]));
Q_ASSIGN U168 ( .B(xcva_top.xc_top.simTime[52]), .A(ctrlW[180]));
Q_ASSIGN U169 ( .B(xcva_top.xc_top.simTime[52]), .A(simTime[52]));
Q_ASSIGN U170 ( .B(xcva_top.xc_top.simTime[53]), .A(ctrlW[181]));
Q_ASSIGN U171 ( .B(xcva_top.xc_top.simTime[53]), .A(simTime[53]));
Q_ASSIGN U172 ( .B(xcva_top.xc_top.simTime[54]), .A(ctrlW[182]));
Q_ASSIGN U173 ( .B(xcva_top.xc_top.simTime[54]), .A(simTime[54]));
Q_ASSIGN U174 ( .B(xcva_top.xc_top.simTime[55]), .A(ctrlW[183]));
Q_ASSIGN U175 ( .B(xcva_top.xc_top.simTime[55]), .A(simTime[55]));
Q_ASSIGN U176 ( .B(xcva_top.xc_top.simTime[56]), .A(ctrlW[184]));
Q_ASSIGN U177 ( .B(xcva_top.xc_top.simTime[56]), .A(simTime[56]));
Q_ASSIGN U178 ( .B(xcva_top.xc_top.simTime[57]), .A(ctrlW[185]));
Q_ASSIGN U179 ( .B(xcva_top.xc_top.simTime[57]), .A(simTime[57]));
Q_ASSIGN U180 ( .B(xcva_top.xc_top.simTime[58]), .A(ctrlW[186]));
Q_ASSIGN U181 ( .B(xcva_top.xc_top.simTime[58]), .A(simTime[58]));
Q_ASSIGN U182 ( .B(xcva_top.xc_top.simTime[59]), .A(ctrlW[187]));
Q_ASSIGN U183 ( .B(xcva_top.xc_top.simTime[59]), .A(simTime[59]));
Q_ASSIGN U184 ( .B(xcva_top.xc_top.simTime[60]), .A(ctrlW[188]));
Q_ASSIGN U185 ( .B(xcva_top.xc_top.simTime[60]), .A(simTime[60]));
Q_ASSIGN U186 ( .B(xcva_top.xc_top.simTime[61]), .A(ctrlW[189]));
Q_ASSIGN U187 ( .B(xcva_top.xc_top.simTime[61]), .A(simTime[61]));
Q_ASSIGN U188 ( .B(xcva_top.xc_top.simTime[62]), .A(ctrlW[190]));
Q_ASSIGN U189 ( .B(xcva_top.xc_top.simTime[62]), .A(simTime[62]));
Q_ASSIGN U190 ( .B(xcva_top.xc_top.simTime[63]), .A(ctrlW[191]));
Q_ASSIGN U191 ( .B(xcva_top.xc_top.simTime[63]), .A(simTime[63]));
Q_BUF U192 ( .A(ecmTs[0]), .Z(ctrlW[64]));
Q_BUF U193 ( .A(ecmTs[1]), .Z(ctrlW[65]));
Q_BUF U194 ( .A(ecmTs[2]), .Z(ctrlW[66]));
Q_BUF U195 ( .A(ecmTs[3]), .Z(ctrlW[67]));
Q_BUF U196 ( .A(ecmTs[4]), .Z(ctrlW[68]));
Q_BUF U197 ( .A(ecmTs[5]), .Z(ctrlW[69]));
Q_BUF U198 ( .A(ecmTs[6]), .Z(ctrlW[70]));
Q_BUF U199 ( .A(ecmTs[7]), .Z(ctrlW[71]));
Q_BUF U200 ( .A(ecmTs[8]), .Z(ctrlW[72]));
Q_BUF U201 ( .A(ecmTs[9]), .Z(ctrlW[73]));
Q_BUF U202 ( .A(ecmTs[10]), .Z(ctrlW[74]));
Q_BUF U203 ( .A(ecmTs[11]), .Z(ctrlW[75]));
Q_BUF U204 ( .A(ecmTs[12]), .Z(ctrlW[76]));
Q_BUF U205 ( .A(ecmTs[13]), .Z(ctrlW[77]));
Q_BUF U206 ( .A(ecmTs[14]), .Z(ctrlW[78]));
Q_BUF U207 ( .A(ecmTs[15]), .Z(ctrlW[79]));
Q_BUF U208 ( .A(ecmTs[16]), .Z(ctrlW[80]));
Q_BUF U209 ( .A(ecmTs[17]), .Z(ctrlW[81]));
Q_BUF U210 ( .A(ecmTs[18]), .Z(ctrlW[82]));
Q_BUF U211 ( .A(ecmTs[19]), .Z(ctrlW[83]));
Q_BUF U212 ( .A(ecmTs[20]), .Z(ctrlW[84]));
Q_BUF U213 ( .A(ecmTs[21]), .Z(ctrlW[85]));
Q_BUF U214 ( .A(ecmTs[22]), .Z(ctrlW[86]));
Q_BUF U215 ( .A(ecmTs[23]), .Z(ctrlW[87]));
Q_BUF U216 ( .A(ecmTs[24]), .Z(ctrlW[88]));
Q_BUF U217 ( .A(ecmTs[25]), .Z(ctrlW[89]));
Q_BUF U218 ( .A(ecmTs[26]), .Z(ctrlW[90]));
Q_BUF U219 ( .A(ecmTs[27]), .Z(ctrlW[91]));
Q_BUF U220 ( .A(ecmTs[28]), .Z(ctrlW[92]));
Q_BUF U221 ( .A(ecmTs[29]), .Z(ctrlW[93]));
Q_BUF U222 ( .A(ecmTs[30]), .Z(ctrlW[94]));
Q_BUF U223 ( .A(ecmTs[31]), .Z(ctrlW[95]));
Q_BUF U224 ( .A(ecmTs[32]), .Z(ctrlW[96]));
Q_BUF U225 ( .A(ecmTs[33]), .Z(ctrlW[97]));
Q_BUF U226 ( .A(ecmTs[34]), .Z(ctrlW[98]));
Q_BUF U227 ( .A(ecmTs[35]), .Z(ctrlW[99]));
Q_BUF U228 ( .A(ecmTs[36]), .Z(ctrlW[100]));
Q_BUF U229 ( .A(ecmTs[37]), .Z(ctrlW[101]));
Q_BUF U230 ( .A(ecmTs[38]), .Z(ctrlW[102]));
Q_BUF U231 ( .A(ecmTs[39]), .Z(ctrlW[103]));
Q_BUF U232 ( .A(ecmTs[40]), .Z(ctrlW[104]));
Q_BUF U233 ( .A(ecmTs[41]), .Z(ctrlW[105]));
Q_BUF U234 ( .A(ecmTs[42]), .Z(ctrlW[106]));
Q_BUF U235 ( .A(ecmTs[43]), .Z(ctrlW[107]));
Q_BUF U236 ( .A(ecmTs[44]), .Z(ctrlW[108]));
Q_BUF U237 ( .A(ecmTs[45]), .Z(ctrlW[109]));
Q_BUF U238 ( .A(ecmTs[46]), .Z(ctrlW[110]));
Q_BUF U239 ( .A(ecmTs[47]), .Z(ctrlW[111]));
Q_BUF U240 ( .A(ecmTs[48]), .Z(ctrlW[112]));
Q_BUF U241 ( .A(ecmTs[49]), .Z(ctrlW[113]));
Q_BUF U242 ( .A(ecmTs[50]), .Z(ctrlW[114]));
Q_BUF U243 ( .A(ecmTs[51]), .Z(ctrlW[115]));
Q_BUF U244 ( .A(ecmTs[52]), .Z(ctrlW[116]));
Q_BUF U245 ( .A(ecmTs[53]), .Z(ctrlW[117]));
Q_BUF U246 ( .A(ecmTs[54]), .Z(ctrlW[118]));
Q_BUF U247 ( .A(ecmTs[55]), .Z(ctrlW[119]));
Q_BUF U248 ( .A(ecmTs[56]), .Z(ctrlW[120]));
Q_BUF U249 ( .A(ecmTs[57]), .Z(ctrlW[121]));
Q_BUF U250 ( .A(ecmTs[58]), .Z(ctrlW[122]));
Q_BUF U251 ( .A(ecmTs[59]), .Z(ctrlW[123]));
Q_BUF U252 ( .A(ecmTs[60]), .Z(ctrlW[124]));
Q_BUF U253 ( .A(ecmTs[61]), .Z(ctrlW[125]));
Q_BUF U254 ( .A(ecmTs[62]), .Z(ctrlW[126]));
Q_BUF U255 ( .A(ecmTs[63]), .Z(ctrlW[127]));
Q_BUF U256 ( .A(ctrlR[136]), .Z(ctrlEv[0]));
Q_BUF U257 ( .A(ctrlR[192]), .Z(ctrlEv[1]));
Q_AN02 U258 ( .A0(n1064), .A1(xcva_top.xc_top.ecmOnD), .Z(n1742));
Q_FDP0 U259 ( .CK(uclk), .D(ctrlW[255]), .Q(n1741), .QN( ));
Q_FDP0 U260 ( .CK(uclk), .D(ctrlW[254]), .Q(n1740), .QN( ));
Q_FDP0 U261 ( .CK(uclk), .D(ctrlW[253]), .Q(n1739), .QN( ));
Q_FDP0 U262 ( .CK(uclk), .D(ctrlW[252]), .Q(n1738), .QN( ));
Q_FDP0 U263 ( .CK(uclk), .D(ctrlW[251]), .Q(n1737), .QN( ));
Q_FDP0 U264 ( .CK(uclk), .D(ctrlW[250]), .Q(n1736), .QN( ));
Q_FDP0 U265 ( .CK(uclk), .D(ctrlW[249]), .Q(n1735), .QN( ));
Q_FDP0 U266 ( .CK(uclk), .D(ctrlW[248]), .Q(n1734), .QN( ));
Q_FDP0 U267 ( .CK(uclk), .D(ctrlW[247]), .Q(n1733), .QN( ));
Q_FDP0 U268 ( .CK(uclk), .D(ctrlW[246]), .Q(n1732), .QN( ));
Q_FDP0 U269 ( .CK(uclk), .D(ctrlW[245]), .Q(n1731), .QN( ));
Q_FDP0 U270 ( .CK(uclk), .D(ctrlW[244]), .Q(n1730), .QN( ));
Q_FDP0 U271 ( .CK(uclk), .D(ctrlW[243]), .Q(n1729), .QN( ));
Q_FDP0 U272 ( .CK(uclk), .D(ctrlW[242]), .Q(n1728), .QN( ));
Q_FDP0 U273 ( .CK(uclk), .D(ctrlW[241]), .Q(n1727), .QN( ));
Q_FDP0 U274 ( .CK(uclk), .D(ctrlW[240]), .Q(n1726), .QN( ));
Q_FDP0 U275 ( .CK(uclk), .D(ctrlW[239]), .Q(n1725), .QN( ));
Q_FDP0 U276 ( .CK(uclk), .D(ctrlW[238]), .Q(n1724), .QN( ));
Q_FDP0 U277 ( .CK(uclk), .D(ctrlW[237]), .Q(n1723), .QN( ));
Q_FDP0 U278 ( .CK(uclk), .D(ctrlW[236]), .Q(n1722), .QN( ));
Q_FDP0 U279 ( .CK(uclk), .D(ctrlW[235]), .Q(n1721), .QN( ));
Q_FDP0 U280 ( .CK(uclk), .D(ctrlW[234]), .Q(n1720), .QN( ));
Q_FDP0 U281 ( .CK(uclk), .D(ctrlW[233]), .Q(n1719), .QN( ));
Q_FDP0 U282 ( .CK(uclk), .D(ctrlW[232]), .Q(n1718), .QN( ));
Q_FDP0 U283 ( .CK(uclk), .D(ctrlW[231]), .Q(n1717), .QN( ));
Q_FDP0 U284 ( .CK(uclk), .D(ctrlW[230]), .Q(n1716), .QN( ));
Q_FDP0 U285 ( .CK(uclk), .D(ctrlW[229]), .Q(n1715), .QN( ));
Q_FDP0 U286 ( .CK(uclk), .D(ctrlW[228]), .Q(n1714), .QN( ));
Q_FDP0 U287 ( .CK(uclk), .D(ctrlW[227]), .Q(n1713), .QN( ));
Q_FDP0 U288 ( .CK(uclk), .D(ctrlW[226]), .Q(n1712), .QN( ));
Q_FDP0 U289 ( .CK(uclk), .D(ctrlW[225]), .Q(n1711), .QN( ));
Q_FDP0 U290 ( .CK(uclk), .D(ctrlW[224]), .Q(n1710), .QN( ));
Q_FDP0 U291 ( .CK(uclk), .D(ctrlW[223]), .Q(n1709), .QN( ));
Q_FDP0 U292 ( .CK(uclk), .D(ctrlW[222]), .Q(n1708), .QN( ));
Q_FDP0 U293 ( .CK(uclk), .D(ctrlW[221]), .Q(n1707), .QN( ));
Q_FDP0 U294 ( .CK(uclk), .D(ctrlW[220]), .Q(n1706), .QN( ));
Q_FDP0 U295 ( .CK(uclk), .D(ctrlW[219]), .Q(n1705), .QN( ));
Q_FDP0 U296 ( .CK(uclk), .D(ctrlW[218]), .Q(n1704), .QN( ));
Q_FDP0 U297 ( .CK(uclk), .D(ctrlW[217]), .Q(n1703), .QN( ));
Q_FDP0 U298 ( .CK(uclk), .D(ctrlW[216]), .Q(n1702), .QN( ));
Q_FDP0 U299 ( .CK(uclk), .D(ctrlW[215]), .Q(n1701), .QN( ));
Q_FDP0 U300 ( .CK(uclk), .D(ctrlW[214]), .Q(n1700), .QN( ));
Q_FDP0 U301 ( .CK(uclk), .D(ctrlW[213]), .Q(n1699), .QN( ));
Q_FDP0 U302 ( .CK(uclk), .D(ctrlW[212]), .Q(n1698), .QN( ));
Q_FDP0 U303 ( .CK(uclk), .D(ctrlW[211]), .Q(n1697), .QN( ));
Q_FDP0 U304 ( .CK(uclk), .D(ctrlW[210]), .Q(n1696), .QN( ));
Q_FDP0 U305 ( .CK(uclk), .D(ctrlW[209]), .Q(n1695), .QN( ));
Q_FDP0 U306 ( .CK(uclk), .D(ctrlW[208]), .Q(n1694), .QN( ));
Q_FDP0 U307 ( .CK(uclk), .D(ctrlW[207]), .Q(n1693), .QN( ));
Q_FDP0 U308 ( .CK(uclk), .D(ctrlW[206]), .Q(n1692), .QN( ));
Q_FDP0 U309 ( .CK(uclk), .D(ctrlW[205]), .Q(n1691), .QN( ));
Q_FDP0 U310 ( .CK(uclk), .D(ctrlW[204]), .Q(n1690), .QN( ));
Q_FDP0 U311 ( .CK(uclk), .D(ctrlW[203]), .Q(n1689), .QN( ));
Q_FDP0 U312 ( .CK(uclk), .D(ctrlW[202]), .Q(n1688), .QN( ));
Q_FDP0 U313 ( .CK(uclk), .D(ctrlW[201]), .Q(n1687), .QN( ));
Q_FDP0 U314 ( .CK(uclk), .D(ctrlW[200]), .Q(n1686), .QN( ));
Q_FDP0 U315 ( .CK(uclk), .D(ctrlW[199]), .Q(n1685), .QN( ));
Q_FDP0 U316 ( .CK(uclk), .D(ctrlW[198]), .Q(n1684), .QN( ));
Q_FDP0 U317 ( .CK(uclk), .D(ctrlW[197]), .Q(n1683), .QN( ));
Q_FDP0 U318 ( .CK(uclk), .D(ctrlW[196]), .Q(n1682), .QN( ));
Q_FDP0 U319 ( .CK(uclk), .D(ctrlW[195]), .Q(n1681), .QN( ));
Q_FDP0 U320 ( .CK(uclk), .D(ctrlW[194]), .Q(n1680), .QN( ));
Q_FDP0 U321 ( .CK(uclk), .D(ctrlW[193]), .Q(n1679), .QN( ));
Q_FDP0 U322 ( .CK(uclk), .D(ctrlW[192]), .Q(n1678), .QN( ));
Q_FDP0 U323 ( .CK(uclk), .D(xcva_top.xc_top.simTime[63]), .Q(n1677), .QN( ));
Q_FDP0 U324 ( .CK(uclk), .D(xcva_top.xc_top.simTime[62]), .Q(n1676), .QN( ));
Q_FDP0 U325 ( .CK(uclk), .D(xcva_top.xc_top.simTime[61]), .Q(n1675), .QN( ));
Q_FDP0 U326 ( .CK(uclk), .D(xcva_top.xc_top.simTime[60]), .Q(n1674), .QN( ));
Q_FDP0 U327 ( .CK(uclk), .D(xcva_top.xc_top.simTime[59]), .Q(n1673), .QN( ));
Q_FDP0 U328 ( .CK(uclk), .D(xcva_top.xc_top.simTime[58]), .Q(n1672), .QN( ));
Q_FDP0 U329 ( .CK(uclk), .D(xcva_top.xc_top.simTime[57]), .Q(n1671), .QN( ));
Q_FDP0 U330 ( .CK(uclk), .D(xcva_top.xc_top.simTime[56]), .Q(n1670), .QN( ));
Q_FDP0 U331 ( .CK(uclk), .D(xcva_top.xc_top.simTime[55]), .Q(n1669), .QN( ));
Q_FDP0 U332 ( .CK(uclk), .D(xcva_top.xc_top.simTime[54]), .Q(n1668), .QN( ));
Q_FDP0 U333 ( .CK(uclk), .D(xcva_top.xc_top.simTime[53]), .Q(n1667), .QN( ));
Q_FDP0 U334 ( .CK(uclk), .D(xcva_top.xc_top.simTime[52]), .Q(n1666), .QN( ));
Q_FDP0 U335 ( .CK(uclk), .D(xcva_top.xc_top.simTime[51]), .Q(n1665), .QN( ));
Q_FDP0 U336 ( .CK(uclk), .D(xcva_top.xc_top.simTime[50]), .Q(n1664), .QN( ));
Q_FDP0 U337 ( .CK(uclk), .D(xcva_top.xc_top.simTime[49]), .Q(n1663), .QN( ));
Q_FDP0 U338 ( .CK(uclk), .D(xcva_top.xc_top.simTime[48]), .Q(n1662), .QN( ));
Q_FDP0 U339 ( .CK(uclk), .D(xcva_top.xc_top.simTime[47]), .Q(n1661), .QN( ));
Q_FDP0 U340 ( .CK(uclk), .D(xcva_top.xc_top.simTime[46]), .Q(n1660), .QN( ));
Q_FDP0 U341 ( .CK(uclk), .D(xcva_top.xc_top.simTime[45]), .Q(n1659), .QN( ));
Q_FDP0 U342 ( .CK(uclk), .D(xcva_top.xc_top.simTime[44]), .Q(n1658), .QN( ));
Q_FDP0 U343 ( .CK(uclk), .D(xcva_top.xc_top.simTime[43]), .Q(n1657), .QN( ));
Q_FDP0 U344 ( .CK(uclk), .D(xcva_top.xc_top.simTime[42]), .Q(n1656), .QN( ));
Q_FDP0 U345 ( .CK(uclk), .D(xcva_top.xc_top.simTime[41]), .Q(n1655), .QN( ));
Q_FDP0 U346 ( .CK(uclk), .D(xcva_top.xc_top.simTime[40]), .Q(n1654), .QN( ));
Q_FDP0 U347 ( .CK(uclk), .D(xcva_top.xc_top.simTime[39]), .Q(n1653), .QN( ));
Q_FDP0 U348 ( .CK(uclk), .D(xcva_top.xc_top.simTime[38]), .Q(n1652), .QN( ));
Q_FDP0 U349 ( .CK(uclk), .D(xcva_top.xc_top.simTime[37]), .Q(n1651), .QN( ));
Q_FDP0 U350 ( .CK(uclk), .D(xcva_top.xc_top.simTime[36]), .Q(n1650), .QN( ));
Q_FDP0 U351 ( .CK(uclk), .D(xcva_top.xc_top.simTime[35]), .Q(n1649), .QN( ));
Q_FDP0 U352 ( .CK(uclk), .D(xcva_top.xc_top.simTime[34]), .Q(n1648), .QN( ));
Q_FDP0 U353 ( .CK(uclk), .D(xcva_top.xc_top.simTime[33]), .Q(n1647), .QN( ));
Q_FDP0 U354 ( .CK(uclk), .D(xcva_top.xc_top.simTime[32]), .Q(n1646), .QN( ));
Q_FDP0 U355 ( .CK(uclk), .D(xcva_top.xc_top.simTime[31]), .Q(n1645), .QN( ));
Q_FDP0 U356 ( .CK(uclk), .D(xcva_top.xc_top.simTime[30]), .Q(n1644), .QN( ));
Q_FDP0 U357 ( .CK(uclk), .D(xcva_top.xc_top.simTime[29]), .Q(n1643), .QN( ));
Q_FDP0 U358 ( .CK(uclk), .D(xcva_top.xc_top.simTime[28]), .Q(n1642), .QN( ));
Q_FDP0 U359 ( .CK(uclk), .D(xcva_top.xc_top.simTime[27]), .Q(n1641), .QN( ));
Q_FDP0 U360 ( .CK(uclk), .D(xcva_top.xc_top.simTime[26]), .Q(n1640), .QN( ));
Q_FDP0 U361 ( .CK(uclk), .D(xcva_top.xc_top.simTime[25]), .Q(n1639), .QN( ));
Q_FDP0 U362 ( .CK(uclk), .D(xcva_top.xc_top.simTime[24]), .Q(n1638), .QN( ));
Q_FDP0 U363 ( .CK(uclk), .D(xcva_top.xc_top.simTime[23]), .Q(n1637), .QN( ));
Q_FDP0 U364 ( .CK(uclk), .D(xcva_top.xc_top.simTime[22]), .Q(n1636), .QN( ));
Q_FDP0 U365 ( .CK(uclk), .D(xcva_top.xc_top.simTime[21]), .Q(n1635), .QN( ));
Q_FDP0 U366 ( .CK(uclk), .D(xcva_top.xc_top.simTime[20]), .Q(n1634), .QN( ));
Q_FDP0 U367 ( .CK(uclk), .D(xcva_top.xc_top.simTime[19]), .Q(n1633), .QN( ));
Q_FDP0 U368 ( .CK(uclk), .D(xcva_top.xc_top.simTime[18]), .Q(n1632), .QN( ));
Q_FDP0 U369 ( .CK(uclk), .D(xcva_top.xc_top.simTime[17]), .Q(n1631), .QN( ));
Q_FDP0 U370 ( .CK(uclk), .D(xcva_top.xc_top.simTime[16]), .Q(n1630), .QN( ));
Q_FDP0 U371 ( .CK(uclk), .D(xcva_top.xc_top.simTime[15]), .Q(n1629), .QN( ));
Q_FDP0 U372 ( .CK(uclk), .D(xcva_top.xc_top.simTime[14]), .Q(n1628), .QN( ));
Q_FDP0 U373 ( .CK(uclk), .D(xcva_top.xc_top.simTime[13]), .Q(n1627), .QN( ));
Q_FDP0 U374 ( .CK(uclk), .D(xcva_top.xc_top.simTime[12]), .Q(n1626), .QN( ));
Q_FDP0 U375 ( .CK(uclk), .D(xcva_top.xc_top.simTime[11]), .Q(n1625), .QN( ));
Q_FDP0 U376 ( .CK(uclk), .D(xcva_top.xc_top.simTime[10]), .Q(n1624), .QN( ));
Q_FDP0 U377 ( .CK(uclk), .D(xcva_top.xc_top.simTime[9]), .Q(n1623), .QN( ));
Q_FDP0 U378 ( .CK(uclk), .D(xcva_top.xc_top.simTime[8]), .Q(n1622), .QN( ));
Q_FDP0 U379 ( .CK(uclk), .D(xcva_top.xc_top.simTime[7]), .Q(n1621), .QN( ));
Q_FDP0 U380 ( .CK(uclk), .D(xcva_top.xc_top.simTime[6]), .Q(n1620), .QN( ));
Q_FDP0 U381 ( .CK(uclk), .D(xcva_top.xc_top.simTime[5]), .Q(n1619), .QN( ));
Q_FDP0 U382 ( .CK(uclk), .D(xcva_top.xc_top.simTime[4]), .Q(n1618), .QN( ));
Q_FDP0 U383 ( .CK(uclk), .D(xcva_top.xc_top.simTime[3]), .Q(n1617), .QN( ));
Q_FDP0 U384 ( .CK(uclk), .D(xcva_top.xc_top.simTime[2]), .Q(n1616), .QN( ));
Q_FDP0 U385 ( .CK(uclk), .D(xcva_top.xc_top.simTime[1]), .Q(n1615), .QN( ));
Q_FDP0 U386 ( .CK(uclk), .D(xcva_top.xc_top.simTime[0]), .Q(n1614), .QN( ));
Q_FDP0 U387 ( .CK(uclk), .D(ctrlW[127]), .Q(n1613), .QN( ));
Q_FDP0 U388 ( .CK(uclk), .D(ctrlW[126]), .Q(n1612), .QN( ));
Q_FDP0 U389 ( .CK(uclk), .D(ctrlW[125]), .Q(n1611), .QN( ));
Q_FDP0 U390 ( .CK(uclk), .D(ctrlW[124]), .Q(n1610), .QN( ));
Q_FDP0 U391 ( .CK(uclk), .D(ctrlW[123]), .Q(n1609), .QN( ));
Q_FDP0 U392 ( .CK(uclk), .D(ctrlW[122]), .Q(n1608), .QN( ));
Q_FDP0 U393 ( .CK(uclk), .D(ctrlW[121]), .Q(n1607), .QN( ));
Q_FDP0 U394 ( .CK(uclk), .D(ctrlW[120]), .Q(n1606), .QN( ));
Q_FDP0 U395 ( .CK(uclk), .D(ctrlW[119]), .Q(n1605), .QN( ));
Q_FDP0 U396 ( .CK(uclk), .D(ctrlW[118]), .Q(n1604), .QN( ));
Q_FDP0 U397 ( .CK(uclk), .D(ctrlW[117]), .Q(n1603), .QN( ));
Q_FDP0 U398 ( .CK(uclk), .D(ctrlW[116]), .Q(n1602), .QN( ));
Q_FDP0 U399 ( .CK(uclk), .D(ctrlW[115]), .Q(n1601), .QN( ));
Q_FDP0 U400 ( .CK(uclk), .D(ctrlW[114]), .Q(n1600), .QN( ));
Q_FDP0 U401 ( .CK(uclk), .D(ctrlW[113]), .Q(n1599), .QN( ));
Q_FDP0 U402 ( .CK(uclk), .D(ctrlW[112]), .Q(n1598), .QN( ));
Q_FDP0 U403 ( .CK(uclk), .D(ctrlW[111]), .Q(n1597), .QN( ));
Q_FDP0 U404 ( .CK(uclk), .D(ctrlW[110]), .Q(n1596), .QN( ));
Q_FDP0 U405 ( .CK(uclk), .D(ctrlW[109]), .Q(n1595), .QN( ));
Q_FDP0 U406 ( .CK(uclk), .D(ctrlW[108]), .Q(n1594), .QN( ));
Q_FDP0 U407 ( .CK(uclk), .D(ctrlW[107]), .Q(n1593), .QN( ));
Q_FDP0 U408 ( .CK(uclk), .D(ctrlW[106]), .Q(n1592), .QN( ));
Q_FDP0 U409 ( .CK(uclk), .D(ctrlW[105]), .Q(n1591), .QN( ));
Q_FDP0 U410 ( .CK(uclk), .D(ctrlW[104]), .Q(n1590), .QN( ));
Q_FDP0 U411 ( .CK(uclk), .D(ctrlW[103]), .Q(n1589), .QN( ));
Q_FDP0 U412 ( .CK(uclk), .D(ctrlW[102]), .Q(n1588), .QN( ));
Q_FDP0 U413 ( .CK(uclk), .D(ctrlW[101]), .Q(n1587), .QN( ));
Q_FDP0 U414 ( .CK(uclk), .D(ctrlW[100]), .Q(n1586), .QN( ));
Q_FDP0 U415 ( .CK(uclk), .D(ctrlW[99]), .Q(n1585), .QN( ));
Q_FDP0 U416 ( .CK(uclk), .D(ctrlW[98]), .Q(n1584), .QN( ));
Q_FDP0 U417 ( .CK(uclk), .D(ctrlW[97]), .Q(n1583), .QN( ));
Q_FDP0 U418 ( .CK(uclk), .D(ctrlW[96]), .Q(n1582), .QN( ));
Q_FDP0 U419 ( .CK(uclk), .D(ctrlW[95]), .Q(n1581), .QN( ));
Q_FDP0 U420 ( .CK(uclk), .D(ctrlW[94]), .Q(n1580), .QN( ));
Q_FDP0 U421 ( .CK(uclk), .D(ctrlW[93]), .Q(n1579), .QN( ));
Q_FDP0 U422 ( .CK(uclk), .D(ctrlW[92]), .Q(n1578), .QN( ));
Q_FDP0 U423 ( .CK(uclk), .D(ctrlW[91]), .Q(n1577), .QN( ));
Q_FDP0 U424 ( .CK(uclk), .D(ctrlW[90]), .Q(n1576), .QN( ));
Q_FDP0 U425 ( .CK(uclk), .D(ctrlW[89]), .Q(n1575), .QN( ));
Q_FDP0 U426 ( .CK(uclk), .D(ctrlW[88]), .Q(n1574), .QN( ));
Q_FDP0 U427 ( .CK(uclk), .D(ctrlW[87]), .Q(n1573), .QN( ));
Q_FDP0 U428 ( .CK(uclk), .D(ctrlW[86]), .Q(n1572), .QN( ));
Q_FDP0 U429 ( .CK(uclk), .D(ctrlW[85]), .Q(n1571), .QN( ));
Q_FDP0 U430 ( .CK(uclk), .D(ctrlW[84]), .Q(n1570), .QN( ));
Q_FDP0 U431 ( .CK(uclk), .D(ctrlW[83]), .Q(n1569), .QN( ));
Q_FDP0 U432 ( .CK(uclk), .D(ctrlW[82]), .Q(n1568), .QN( ));
Q_FDP0 U433 ( .CK(uclk), .D(ctrlW[81]), .Q(n1567), .QN( ));
Q_FDP0 U434 ( .CK(uclk), .D(ctrlW[80]), .Q(n1566), .QN( ));
Q_FDP0 U435 ( .CK(uclk), .D(ctrlW[79]), .Q(n1565), .QN( ));
Q_FDP0 U436 ( .CK(uclk), .D(ctrlW[78]), .Q(n1564), .QN( ));
Q_FDP0 U437 ( .CK(uclk), .D(ctrlW[77]), .Q(n1563), .QN( ));
Q_FDP0 U438 ( .CK(uclk), .D(ctrlW[76]), .Q(n1562), .QN( ));
Q_FDP0 U439 ( .CK(uclk), .D(ctrlW[75]), .Q(n1561), .QN( ));
Q_FDP0 U440 ( .CK(uclk), .D(ctrlW[74]), .Q(n1560), .QN( ));
Q_FDP0 U441 ( .CK(uclk), .D(ctrlW[73]), .Q(n1559), .QN( ));
Q_FDP0 U442 ( .CK(uclk), .D(ctrlW[72]), .Q(n1558), .QN( ));
Q_FDP0 U443 ( .CK(uclk), .D(ctrlW[71]), .Q(n1557), .QN( ));
Q_FDP0 U444 ( .CK(uclk), .D(ctrlW[70]), .Q(n1556), .QN( ));
Q_FDP0 U445 ( .CK(uclk), .D(ctrlW[69]), .Q(n1555), .QN( ));
Q_FDP0 U446 ( .CK(uclk), .D(ctrlW[68]), .Q(n1554), .QN( ));
Q_FDP0 U447 ( .CK(uclk), .D(ctrlW[67]), .Q(n1553), .QN( ));
Q_FDP0 U448 ( .CK(uclk), .D(ctrlW[66]), .Q(n1552), .QN( ));
Q_FDP0 U449 ( .CK(uclk), .D(ctrlW[65]), .Q(n1551), .QN( ));
Q_FDP0 U450 ( .CK(uclk), .D(ctrlW[64]), .Q(n1550), .QN( ));
Q_FDP0 U451 ( .CK(uclk), .D(ctrlW[63]), .Q(n1549), .QN( ));
Q_FDP0 U452 ( .CK(uclk), .D(ctrlW[62]), .Q(n1548), .QN( ));
Q_FDP0 U453 ( .CK(uclk), .D(ctrlW[61]), .Q(n1547), .QN( ));
Q_FDP0 U454 ( .CK(uclk), .D(ctrlW[60]), .Q(n1546), .QN( ));
Q_FDP0 U455 ( .CK(uclk), .D(ctrlW[59]), .Q(n1545), .QN( ));
Q_FDP0 U456 ( .CK(uclk), .D(ctrlW[58]), .Q(n1544), .QN( ));
Q_FDP0 U457 ( .CK(uclk), .D(ctrlW[57]), .Q(n1543), .QN( ));
Q_FDP0 U458 ( .CK(uclk), .D(ctrlW[56]), .Q(n1542), .QN( ));
Q_FDP0 U459 ( .CK(uclk), .D(ctrlW[55]), .Q(n1541), .QN( ));
Q_FDP0 U460 ( .CK(uclk), .D(ctrlW[54]), .Q(n1540), .QN( ));
Q_FDP0 U461 ( .CK(uclk), .D(ctrlW[53]), .Q(n1539), .QN( ));
Q_FDP0 U462 ( .CK(uclk), .D(ctrlW[52]), .Q(n1538), .QN( ));
Q_FDP0 U463 ( .CK(uclk), .D(ctrlW[51]), .Q(n1537), .QN( ));
Q_FDP0 U464 ( .CK(uclk), .D(ctrlW[50]), .Q(n1536), .QN( ));
Q_FDP0 U465 ( .CK(uclk), .D(ctrlW[49]), .Q(n1535), .QN( ));
Q_FDP0 U466 ( .CK(uclk), .D(ctrlW[48]), .Q(n1534), .QN( ));
Q_FDP0 U467 ( .CK(uclk), .D(ctrlW[47]), .Q(n1533), .QN( ));
Q_FDP0 U468 ( .CK(uclk), .D(ctrlW[46]), .Q(n1532), .QN( ));
Q_FDP0 U469 ( .CK(uclk), .D(ctrlW[45]), .Q(n1531), .QN( ));
Q_FDP0 U470 ( .CK(uclk), .D(ctrlW[44]), .Q(n1530), .QN( ));
Q_FDP0 U471 ( .CK(uclk), .D(ctrlW[43]), .Q(n1529), .QN( ));
Q_FDP0 U472 ( .CK(uclk), .D(ctrlW[42]), .Q(n1528), .QN( ));
Q_FDP0 U473 ( .CK(uclk), .D(ctrlW[41]), .Q(n1527), .QN( ));
Q_FDP0 U474 ( .CK(uclk), .D(ctrlW[40]), .Q(n1526), .QN( ));
Q_FDP0 U475 ( .CK(uclk), .D(ctrlW[39]), .Q(n1525), .QN( ));
Q_FDP0 U476 ( .CK(uclk), .D(ctrlW[38]), .Q(n1524), .QN( ));
Q_FDP0 U477 ( .CK(uclk), .D(ctrlW[37]), .Q(n1523), .QN( ));
Q_FDP0 U478 ( .CK(uclk), .D(ctrlW[36]), .Q(n1522), .QN( ));
Q_FDP0 U479 ( .CK(uclk), .D(ctrlW[35]), .Q(n1521), .QN( ));
Q_FDP0 U480 ( .CK(uclk), .D(ctrlW[34]), .Q(n1520), .QN( ));
Q_FDP0 U481 ( .CK(uclk), .D(ctrlW[33]), .Q(n1519), .QN( ));
Q_FDP0 U482 ( .CK(uclk), .D(ctrlW[32]), .Q(n1518), .QN( ));
Q_FDP0 U483 ( .CK(uclk), .D(ctrlW[31]), .Q(n1517), .QN( ));
Q_FDP0 U484 ( .CK(uclk), .D(ctrlW[30]), .Q(n1516), .QN( ));
Q_FDP0 U485 ( .CK(uclk), .D(ctrlW[29]), .Q(n1515), .QN( ));
Q_FDP0 U486 ( .CK(uclk), .D(ctrlW[28]), .Q(n1514), .QN( ));
Q_FDP0 U487 ( .CK(uclk), .D(ctrlW[27]), .Q(n1513), .QN( ));
Q_FDP0 U488 ( .CK(uclk), .D(ctrlW[26]), .Q(n1512), .QN( ));
Q_FDP0 U489 ( .CK(uclk), .D(ctrlW[25]), .Q(n1511), .QN( ));
Q_FDP0 U490 ( .CK(uclk), .D(ctrlW[24]), .Q(n1510), .QN( ));
Q_FDP0 U491 ( .CK(uclk), .D(ctrlW[23]), .Q(n1509), .QN( ));
Q_FDP0 U492 ( .CK(uclk), .D(ctrlW[22]), .Q(n1508), .QN( ));
Q_FDP0 U493 ( .CK(uclk), .D(ctrlW[21]), .Q(n1507), .QN( ));
Q_FDP0 U494 ( .CK(uclk), .D(ctrlW[20]), .Q(n1506), .QN( ));
Q_FDP0 U495 ( .CK(uclk), .D(ctrlW[19]), .Q(n1505), .QN( ));
Q_FDP0 U496 ( .CK(uclk), .D(ctrlW[18]), .Q(n1504), .QN( ));
Q_FDP0 U497 ( .CK(uclk), .D(ctrlW[17]), .Q(n1503), .QN( ));
Q_FDP0 U498 ( .CK(uclk), .D(ctrlW[16]), .Q(n1502), .QN( ));
Q_FDP0 U499 ( .CK(uclk), .D(ctrlW[15]), .Q(n1501), .QN( ));
Q_FDP0 U500 ( .CK(uclk), .D(ctrlW[14]), .Q(n1500), .QN( ));
Q_FDP0 U501 ( .CK(uclk), .D(ctrlW[13]), .Q(n1499), .QN( ));
Q_FDP0 U502 ( .CK(uclk), .D(ctrlW[12]), .Q(n1498), .QN( ));
Q_FDP0 U503 ( .CK(uclk), .D(ctrlW[11]), .Q(n1497), .QN( ));
Q_FDP0 U504 ( .CK(uclk), .D(ctrlW[10]), .Q(n1496), .QN( ));
Q_FDP0 U505 ( .CK(uclk), .D(ctrlW[9]), .Q(n1495), .QN( ));
Q_FDP0 U506 ( .CK(uclk), .D(ctrlW[8]), .Q(n1494), .QN( ));
Q_FDP0 U507 ( .CK(uclk), .D(ctrlW[7]), .Q(n1493), .QN( ));
Q_FDP0 U508 ( .CK(uclk), .D(ctrlW[6]), .Q(n1492), .QN( ));
Q_FDP0 U509 ( .CK(uclk), .D(ctrlW[5]), .Q(n1491), .QN( ));
Q_FDP0 U510 ( .CK(uclk), .D(ctrlW[4]), .Q(n1490), .QN( ));
Q_FDP0 U511 ( .CK(uclk), .D(ctrlW[3]), .Q(n1489), .QN( ));
Q_FDP0 U512 ( .CK(uclk), .D(ctrlW[2]), .Q(n1488), .QN( ));
Q_FDP0 U513 ( .CK(uclk), .D(ctrlW[1]), .Q(n1487), .QN( ));
Q_FDP0 U514 ( .CK(uclk), .D(ctrlW[0]), .Q(n1486), .QN( ));
Q_XOR2 U515 ( .A0(n1482), .A1(n1484), .Z(n1485));
// pragma CVAINTPROP NET n1482 _2_state_ 1
// pragma CVAINTPROP INSTANCE U515 NOBREAKS 1
Q_FDP0B U516 ( .D(n1482), .QTFCLK( ), .Q(n1484));
Q_FDP0 U517 ( .CK(uclk), .D(n1483), .Q(n1482), .QN(n1483));
Q_MX02 U518 ( .S(_zyL739_meState1[0]), .A0(n1195), .A1(xcva_top.xc_top.ecmSync), .Z(n1480));
Q_AN02 U519 ( .A0(_zyL739_meState1[0]), .A1(xcva_top.xc_top.ecmSync), .Z(n1481));
Q_FDP0UA U520 ( .D(n1479), .QTFCLK( ), .Q(_zyL739_meState1[0]));
Q_INV U521 ( .A(n1480), .Z(n1479));
Q_MX02 U522 ( .S(n1481), .A0(ctrlW[192]), .A1(syncId[0]), .Z(n1478));
Q_FDP0UA U523 ( .D(n1478), .QTFCLK( ), .Q(ctrlW[192]));
Q_MX02 U524 ( .S(n1481), .A0(ctrlW[193]), .A1(syncId[1]), .Z(n1477));
Q_FDP0UA U525 ( .D(n1477), .QTFCLK( ), .Q(ctrlW[193]));
Q_MX02 U526 ( .S(n1481), .A0(ctrlW[194]), .A1(syncId[2]), .Z(n1476));
Q_FDP0UA U527 ( .D(n1476), .QTFCLK( ), .Q(ctrlW[194]));
Q_MX02 U528 ( .S(n1481), .A0(ctrlW[195]), .A1(syncId[3]), .Z(n1475));
Q_FDP0UA U529 ( .D(n1475), .QTFCLK( ), .Q(ctrlW[195]));
Q_MX02 U530 ( .S(n1481), .A0(ctrlW[196]), .A1(syncId[4]), .Z(n1474));
Q_FDP0UA U531 ( .D(n1474), .QTFCLK( ), .Q(ctrlW[196]));
Q_MX02 U532 ( .S(n1481), .A0(ctrlW[197]), .A1(syncId[5]), .Z(n1473));
Q_FDP0UA U533 ( .D(n1473), .QTFCLK( ), .Q(ctrlW[197]));
Q_MX02 U534 ( .S(n1481), .A0(ctrlW[198]), .A1(syncId[6]), .Z(n1472));
Q_FDP0UA U535 ( .D(n1472), .QTFCLK( ), .Q(ctrlW[198]));
Q_MX02 U536 ( .S(n1481), .A0(ctrlW[199]), .A1(syncId[7]), .Z(n1471));
Q_FDP0UA U537 ( .D(n1471), .QTFCLK( ), .Q(ctrlW[199]));
Q_AN02 U538 ( .A0(n1414), .A1(ctrlW[200]), .Z(n1470));
Q_FDP0UA U539 ( .D(n1470), .QTFCLK( ), .Q(ctrlW[200]));
Q_AN02 U540 ( .A0(n1414), .A1(ctrlW[201]), .Z(n1469));
Q_FDP0UA U541 ( .D(n1469), .QTFCLK( ), .Q(ctrlW[201]));
Q_AN02 U542 ( .A0(n1414), .A1(ctrlW[202]), .Z(n1468));
Q_FDP0UA U543 ( .D(n1468), .QTFCLK( ), .Q(ctrlW[202]));
Q_AN02 U544 ( .A0(n1414), .A1(ctrlW[203]), .Z(n1467));
Q_FDP0UA U545 ( .D(n1467), .QTFCLK( ), .Q(ctrlW[203]));
Q_AN02 U546 ( .A0(n1414), .A1(ctrlW[204]), .Z(n1466));
Q_FDP0UA U547 ( .D(n1466), .QTFCLK( ), .Q(ctrlW[204]));
Q_AN02 U548 ( .A0(n1414), .A1(ctrlW[205]), .Z(n1465));
Q_FDP0UA U549 ( .D(n1465), .QTFCLK( ), .Q(ctrlW[205]));
Q_AN02 U550 ( .A0(n1414), .A1(ctrlW[206]), .Z(n1464));
Q_FDP0UA U551 ( .D(n1464), .QTFCLK( ), .Q(ctrlW[206]));
Q_AN02 U552 ( .A0(n1414), .A1(ctrlW[207]), .Z(n1463));
Q_FDP0UA U553 ( .D(n1463), .QTFCLK( ), .Q(ctrlW[207]));
Q_AN02 U554 ( .A0(n1414), .A1(ctrlW[208]), .Z(n1462));
Q_FDP0UA U555 ( .D(n1462), .QTFCLK( ), .Q(ctrlW[208]));
Q_AN02 U556 ( .A0(n1414), .A1(ctrlW[209]), .Z(n1461));
Q_FDP0UA U557 ( .D(n1461), .QTFCLK( ), .Q(ctrlW[209]));
Q_AN02 U558 ( .A0(n1414), .A1(ctrlW[210]), .Z(n1460));
Q_FDP0UA U559 ( .D(n1460), .QTFCLK( ), .Q(ctrlW[210]));
Q_AN02 U560 ( .A0(n1414), .A1(ctrlW[211]), .Z(n1459));
Q_FDP0UA U561 ( .D(n1459), .QTFCLK( ), .Q(ctrlW[211]));
Q_AN02 U562 ( .A0(n1414), .A1(ctrlW[212]), .Z(n1458));
Q_FDP0UA U563 ( .D(n1458), .QTFCLK( ), .Q(ctrlW[212]));
Q_AN02 U564 ( .A0(n1414), .A1(ctrlW[213]), .Z(n1457));
Q_FDP0UA U565 ( .D(n1457), .QTFCLK( ), .Q(ctrlW[213]));
Q_AN02 U566 ( .A0(n1414), .A1(ctrlW[214]), .Z(n1456));
Q_FDP0UA U567 ( .D(n1456), .QTFCLK( ), .Q(ctrlW[214]));
Q_AN02 U568 ( .A0(n1414), .A1(ctrlW[215]), .Z(n1455));
Q_FDP0UA U569 ( .D(n1455), .QTFCLK( ), .Q(ctrlW[215]));
Q_AN02 U570 ( .A0(n1414), .A1(ctrlW[216]), .Z(n1454));
Q_FDP0UA U571 ( .D(n1454), .QTFCLK( ), .Q(ctrlW[216]));
Q_AN02 U572 ( .A0(n1414), .A1(ctrlW[217]), .Z(n1453));
Q_FDP0UA U573 ( .D(n1453), .QTFCLK( ), .Q(ctrlW[217]));
Q_AN02 U574 ( .A0(n1414), .A1(ctrlW[218]), .Z(n1452));
Q_FDP0UA U575 ( .D(n1452), .QTFCLK( ), .Q(ctrlW[218]));
Q_AN02 U576 ( .A0(n1414), .A1(ctrlW[219]), .Z(n1451));
Q_FDP0UA U577 ( .D(n1451), .QTFCLK( ), .Q(ctrlW[219]));
Q_AN02 U578 ( .A0(n1414), .A1(ctrlW[220]), .Z(n1450));
Q_FDP0UA U579 ( .D(n1450), .QTFCLK( ), .Q(ctrlW[220]));
Q_AN02 U580 ( .A0(n1414), .A1(ctrlW[221]), .Z(n1449));
Q_FDP0UA U581 ( .D(n1449), .QTFCLK( ), .Q(ctrlW[221]));
Q_AN02 U582 ( .A0(n1414), .A1(ctrlW[222]), .Z(n1448));
Q_FDP0UA U583 ( .D(n1448), .QTFCLK( ), .Q(ctrlW[222]));
Q_AN02 U584 ( .A0(n1414), .A1(ctrlW[223]), .Z(n1447));
Q_FDP0UA U585 ( .D(n1447), .QTFCLK( ), .Q(ctrlW[223]));
Q_AN02 U586 ( .A0(n1414), .A1(ctrlW[224]), .Z(n1446));
Q_FDP0UA U587 ( .D(n1446), .QTFCLK( ), .Q(ctrlW[224]));
Q_AN02 U588 ( .A0(n1414), .A1(ctrlW[225]), .Z(n1445));
Q_FDP0UA U589 ( .D(n1445), .QTFCLK( ), .Q(ctrlW[225]));
Q_AN02 U590 ( .A0(n1414), .A1(ctrlW[226]), .Z(n1444));
Q_FDP0UA U591 ( .D(n1444), .QTFCLK( ), .Q(ctrlW[226]));
Q_AN02 U592 ( .A0(n1414), .A1(ctrlW[227]), .Z(n1443));
Q_FDP0UA U593 ( .D(n1443), .QTFCLK( ), .Q(ctrlW[227]));
Q_AN02 U594 ( .A0(n1414), .A1(ctrlW[228]), .Z(n1442));
Q_FDP0UA U595 ( .D(n1442), .QTFCLK( ), .Q(ctrlW[228]));
Q_AN02 U596 ( .A0(n1414), .A1(ctrlW[229]), .Z(n1441));
Q_FDP0UA U597 ( .D(n1441), .QTFCLK( ), .Q(ctrlW[229]));
Q_AN02 U598 ( .A0(n1414), .A1(ctrlW[230]), .Z(n1440));
Q_FDP0UA U599 ( .D(n1440), .QTFCLK( ), .Q(ctrlW[230]));
Q_AN02 U600 ( .A0(n1414), .A1(ctrlW[231]), .Z(n1439));
Q_FDP0UA U601 ( .D(n1439), .QTFCLK( ), .Q(ctrlW[231]));
Q_AN02 U602 ( .A0(n1414), .A1(ctrlW[232]), .Z(n1438));
Q_FDP0UA U603 ( .D(n1438), .QTFCLK( ), .Q(ctrlW[232]));
Q_AN02 U604 ( .A0(n1414), .A1(ctrlW[233]), .Z(n1437));
Q_FDP0UA U605 ( .D(n1437), .QTFCLK( ), .Q(ctrlW[233]));
Q_AN02 U606 ( .A0(n1414), .A1(ctrlW[234]), .Z(n1436));
Q_FDP0UA U607 ( .D(n1436), .QTFCLK( ), .Q(ctrlW[234]));
Q_AN02 U608 ( .A0(n1414), .A1(ctrlW[235]), .Z(n1435));
Q_FDP0UA U609 ( .D(n1435), .QTFCLK( ), .Q(ctrlW[235]));
Q_AN02 U610 ( .A0(n1414), .A1(ctrlW[236]), .Z(n1434));
Q_FDP0UA U611 ( .D(n1434), .QTFCLK( ), .Q(ctrlW[236]));
Q_AN02 U612 ( .A0(n1414), .A1(ctrlW[237]), .Z(n1433));
Q_FDP0UA U613 ( .D(n1433), .QTFCLK( ), .Q(ctrlW[237]));
Q_AN02 U614 ( .A0(n1414), .A1(ctrlW[238]), .Z(n1432));
Q_FDP0UA U615 ( .D(n1432), .QTFCLK( ), .Q(ctrlW[238]));
Q_AN02 U616 ( .A0(n1414), .A1(ctrlW[239]), .Z(n1431));
Q_FDP0UA U617 ( .D(n1431), .QTFCLK( ), .Q(ctrlW[239]));
Q_AN02 U618 ( .A0(n1414), .A1(ctrlW[240]), .Z(n1430));
Q_FDP0UA U619 ( .D(n1430), .QTFCLK( ), .Q(ctrlW[240]));
Q_AN02 U620 ( .A0(n1414), .A1(ctrlW[241]), .Z(n1429));
Q_FDP0UA U621 ( .D(n1429), .QTFCLK( ), .Q(ctrlW[241]));
Q_AN02 U622 ( .A0(n1414), .A1(ctrlW[242]), .Z(n1428));
Q_FDP0UA U623 ( .D(n1428), .QTFCLK( ), .Q(ctrlW[242]));
Q_AN02 U624 ( .A0(n1414), .A1(ctrlW[243]), .Z(n1427));
Q_FDP0UA U625 ( .D(n1427), .QTFCLK( ), .Q(ctrlW[243]));
Q_AN02 U626 ( .A0(n1414), .A1(ctrlW[244]), .Z(n1426));
Q_FDP0UA U627 ( .D(n1426), .QTFCLK( ), .Q(ctrlW[244]));
Q_AN02 U628 ( .A0(n1414), .A1(ctrlW[245]), .Z(n1425));
Q_FDP0UA U629 ( .D(n1425), .QTFCLK( ), .Q(ctrlW[245]));
Q_AN02 U630 ( .A0(n1414), .A1(ctrlW[246]), .Z(n1424));
Q_FDP0UA U631 ( .D(n1424), .QTFCLK( ), .Q(ctrlW[246]));
Q_AN02 U632 ( .A0(n1414), .A1(ctrlW[247]), .Z(n1423));
Q_FDP0UA U633 ( .D(n1423), .QTFCLK( ), .Q(ctrlW[247]));
Q_AN02 U634 ( .A0(n1414), .A1(ctrlW[248]), .Z(n1422));
Q_FDP0UA U635 ( .D(n1422), .QTFCLK( ), .Q(ctrlW[248]));
Q_AN02 U636 ( .A0(n1414), .A1(ctrlW[249]), .Z(n1421));
Q_FDP0UA U637 ( .D(n1421), .QTFCLK( ), .Q(ctrlW[249]));
Q_AN02 U638 ( .A0(n1414), .A1(ctrlW[250]), .Z(n1420));
Q_FDP0UA U639 ( .D(n1420), .QTFCLK( ), .Q(ctrlW[250]));
Q_AN02 U640 ( .A0(n1414), .A1(ctrlW[251]), .Z(n1419));
Q_FDP0UA U641 ( .D(n1419), .QTFCLK( ), .Q(ctrlW[251]));
Q_AN02 U642 ( .A0(n1414), .A1(ctrlW[252]), .Z(n1418));
Q_FDP0UA U643 ( .D(n1418), .QTFCLK( ), .Q(ctrlW[252]));
Q_AN02 U644 ( .A0(n1414), .A1(ctrlW[253]), .Z(n1417));
Q_FDP0UA U645 ( .D(n1417), .QTFCLK( ), .Q(ctrlW[253]));
Q_AN02 U646 ( .A0(n1414), .A1(ctrlW[254]), .Z(n1416));
Q_FDP0UA U647 ( .D(n1416), .QTFCLK( ), .Q(ctrlW[254]));
Q_AN02 U648 ( .A0(n1414), .A1(ctrlW[255]), .Z(n1415));
Q_INV U649 ( .A(n1481), .Z(n1414));
Q_FDP0UA U650 ( .D(n1415), .QTFCLK( ), .Q(ctrlW[255]));
Q_MX02 U651 ( .S(_zyL739_meState1[0]), .A0(syncIdP[0]), .A1(syncId[0]), .Z(n1413));
Q_FDP0UA U652 ( .D(n1413), .QTFCLK( ), .Q(syncIdP[0]));
Q_MX02 U653 ( .S(_zyL739_meState1[0]), .A0(syncIdP[1]), .A1(syncId[1]), .Z(n1412));
Q_FDP0UA U654 ( .D(n1412), .QTFCLK( ), .Q(syncIdP[1]));
Q_MX02 U655 ( .S(_zyL739_meState1[0]), .A0(syncIdP[2]), .A1(syncId[2]), .Z(n1411));
Q_FDP0UA U656 ( .D(n1411), .QTFCLK( ), .Q(syncIdP[2]));
Q_MX02 U657 ( .S(_zyL739_meState1[0]), .A0(syncIdP[3]), .A1(syncId[3]), .Z(n1410));
Q_FDP0UA U658 ( .D(n1410), .QTFCLK( ), .Q(syncIdP[3]));
Q_MX02 U659 ( .S(_zyL739_meState1[0]), .A0(syncIdP[4]), .A1(syncId[4]), .Z(n1409));
Q_FDP0UA U660 ( .D(n1409), .QTFCLK( ), .Q(syncIdP[4]));
Q_MX02 U661 ( .S(_zyL739_meState1[0]), .A0(syncIdP[5]), .A1(syncId[5]), .Z(n1408));
Q_FDP0UA U662 ( .D(n1408), .QTFCLK( ), .Q(syncIdP[5]));
Q_MX02 U663 ( .S(_zyL739_meState1[0]), .A0(syncIdP[6]), .A1(syncId[6]), .Z(n1407));
Q_FDP0UA U664 ( .D(n1407), .QTFCLK( ), .Q(syncIdP[6]));
Q_MX02 U665 ( .S(_zyL739_meState1[0]), .A0(syncIdP[7]), .A1(syncId[7]), .Z(n1406));
Q_FDP0UA U666 ( .D(n1406), .QTFCLK( ), .Q(syncIdP[7]));
Q_MX02 U667 ( .S(n1480), .A0(syncId[0]), .A1(ctrlEv[1]), .Z(n1405));
Q_FDP0UA U668 ( .D(n1405), .QTFCLK( ), .Q(syncId[0]));
Q_MX02 U669 ( .S(n1480), .A0(syncId[1]), .A1(ctrlR[193]), .Z(n1404));
Q_FDP0UA U670 ( .D(n1404), .QTFCLK( ), .Q(syncId[1]));
Q_MX02 U671 ( .S(n1480), .A0(syncId[2]), .A1(ctrlR[194]), .Z(n1403));
Q_FDP0UA U672 ( .D(n1403), .QTFCLK( ), .Q(syncId[2]));
Q_MX02 U673 ( .S(n1480), .A0(syncId[3]), .A1(ctrlR[195]), .Z(n1402));
Q_FDP0UA U674 ( .D(n1402), .QTFCLK( ), .Q(syncId[3]));
Q_MX02 U675 ( .S(n1480), .A0(syncId[4]), .A1(ctrlR[196]), .Z(n1401));
Q_FDP0UA U676 ( .D(n1401), .QTFCLK( ), .Q(syncId[4]));
Q_MX02 U677 ( .S(n1480), .A0(syncId[5]), .A1(ctrlR[197]), .Z(n1400));
Q_FDP0UA U678 ( .D(n1400), .QTFCLK( ), .Q(syncId[5]));
Q_MX02 U679 ( .S(n1480), .A0(syncId[6]), .A1(ctrlR[198]), .Z(n1399));
Q_FDP0UA U680 ( .D(n1399), .QTFCLK( ), .Q(syncId[6]));
Q_MX02 U681 ( .S(n1480), .A0(syncId[7]), .A1(ctrlR[199]), .Z(n1398));
Q_FDP0UA U682 ( .D(n1398), .QTFCLK( ), .Q(syncId[7]));
Q_INV U683 ( .A(xcva_top.xc_top.ptxStop), .Z(n1395));
Q_AN02 U684 ( .A0(n1395), .A1(holdEcm), .Z(n1397));
Q_AN02 U685 ( .A0(n1397), .A1(holdEcmD[3]), .Z(n1394));
Q_INV U686 ( .A(holdEcmD[3]), .Z(n1393));
Q_AN02 U687 ( .A0(n1397), .A1(n1393), .Z(n1396));
Q_FDP0UA U688 ( .D(n1396), .QTFCLK( ), .Q(holdEcmBusy));
Q_MX02 U689 ( .S(n1394), .A0(n1385), .A1(holdEcmD[0]), .Z(n1392));
Q_FDP0UA U690 ( .D(n1392), .QTFCLK( ), .Q(holdEcmD[0]));
Q_MX02 U691 ( .S(n1394), .A0(n1386), .A1(holdEcmD[1]), .Z(n1391));
Q_FDP0UA U692 ( .D(n1391), .QTFCLK( ), .Q(holdEcmD[1]));
Q_MX02 U693 ( .S(n1394), .A0(n1387), .A1(holdEcmD[2]), .Z(n1390));
Q_FDP0UA U694 ( .D(n1390), .QTFCLK( ), .Q(holdEcmD[2]));
Q_MX02 U695 ( .S(n1394), .A0(n1388), .A1(holdEcmD[3]), .Z(n1389));
Q_FDP0UA U696 ( .D(n1389), .QTFCLK( ), .Q(holdEcmD[3]));
Q_AN02 U697 ( .A0(n1397), .A1(n1384), .Z(n1388));
Q_AN02 U698 ( .A0(n1397), .A1(n1382), .Z(n1387));
Q_AN02 U699 ( .A0(n1397), .A1(n1380), .Z(n1386));
Q_AN02 U700 ( .A0(n1397), .A1(n1379), .Z(n1385));
Q_XOR2 U701 ( .A0(holdEcmD[3]), .A1(n1383), .Z(n1384));
Q_AD01HF U702 ( .A0(holdEcmD[2]), .B0(n1381), .S(n1382), .CO(n1383));
Q_AD01HF U703 ( .A0(holdEcmD[1]), .B0(holdEcmD[0]), .S(n1380), .CO(n1381));
Q_INV U704 ( .A(holdEcmD[0]), .Z(n1379));
Q_FDP0UA U705 ( .D(n1378), .QTFCLK( ), .Q(cRet[0]));
Q_FDP0UA U706 ( .D(n1377), .QTFCLK( ), .Q(cRet[2]));
Q_MX02 U707 ( .S(xcva_top.xc_top.ptxStop), .A0(holdEcmD[3]), .A1(n1377), .Z(n1378));
Q_INV U708 ( .A(xcva_top.xc_top.evalOnC), .Z(n1377));
Q_FDP0UA U709 ( .D(xcva_top.xc_top.ecmSync), .QTFCLK( ), .Q(cRet[1]));
Q_FDP0UA U710 ( .D(sdlStopRply), .QTFCLK( ), .Q(cRet[3]));
Q_FDP0UA U711 ( .D(ctrlEv[0]), .QTFCLK( ), .Q(cmdCnt[0]));
Q_FDP0UA U712 ( .D(ctrlR[137]), .QTFCLK( ), .Q(cmdCnt[1]));
Q_FDP0UA U713 ( .D(ctrlR[138]), .QTFCLK( ), .Q(cmdCnt[2]));
Q_FDP0UA U714 ( .D(ctrlR[139]), .QTFCLK( ), .Q(cmdCnt[3]));
Q_FDP0UA U715 ( .D(ctrlR[140]), .QTFCLK( ), .Q(cmdCnt[4]));
Q_FDP0UA U716 ( .D(ctrlR[141]), .QTFCLK( ), .Q(cmdCnt[5]));
Q_FDP0UA U717 ( .D(ctrlR[142]), .QTFCLK( ), .Q(cmdCnt[6]));
Q_FDP0UA U718 ( .D(ctrlR[143]), .QTFCLK( ), .Q(cmdCnt[7]));
Q_FDP0UA U719 ( .D(ctrlR[128]), .QTFCLK( ), .Q(cmdC[0]));
Q_FDP0UA U720 ( .D(ctrlR[129]), .QTFCLK( ), .Q(cmdC[1]));
Q_FDP0UA U721 ( .D(ctrlR[130]), .QTFCLK( ), .Q(cmdC[2]));
Q_FDP0UA U722 ( .D(ctrlR[131]), .QTFCLK( ), .Q(cmdC[3]));
Q_FDP0UA U723 ( .D(ctrlR[132]), .QTFCLK( ), .Q(cmdC[4]));
Q_FDP0UA U724 ( .D(ctrlR[133]), .QTFCLK( ), .Q(cmdC[5]));
Q_FDP0UA U725 ( .D(ctrlR[134]), .QTFCLK( ), .Q(cmdC[6]));
Q_FDP0UA U726 ( .D(ctrlR[135]), .QTFCLK( ), .Q(cmdC[7]));
Q_AN02 U727 ( .A0(_zyL692_meState0[0]), .A1(n1376), .Z(n1375));
Q_INV U728 ( .A(_zyL692_meState0[0]), .Z(n1373));
Q_AN02 U729 ( .A0(n1373), .A1(n1207), .Z(n1372));
Q_NR02 U730 ( .A0(n1372), .A1(n1375), .Z(n1374));
Q_FDP0UA U731 ( .D(n1374), .QTFCLK( ), .Q(_zyL692_meState0[0]));
Q_ND03 U732 ( .A0(cmdC[0]), .A1(xcva_top.xc_top.ptxStop), .A2(xcva_top.xc_top.evalOnC), .Z(n1376));
Q_MX02 U733 ( .S(n1375), .A0(ctrlW[8]), .A1(cmdCnt[0]), .Z(n1371));
Q_FDP0UA U734 ( .D(n1371), .QTFCLK( ), .Q(cRet[8]));
Q_MX02 U735 ( .S(n1375), .A0(ctrlW[9]), .A1(cmdCnt[1]), .Z(n1370));
Q_FDP0UA U736 ( .D(n1370), .QTFCLK( ), .Q(cRet[9]));
Q_MX02 U737 ( .S(n1375), .A0(ctrlW[10]), .A1(cmdCnt[2]), .Z(n1369));
Q_FDP0UA U738 ( .D(n1369), .QTFCLK( ), .Q(cRet[10]));
Q_MX02 U739 ( .S(n1375), .A0(ctrlW[11]), .A1(cmdCnt[3]), .Z(n1368));
Q_FDP0UA U740 ( .D(n1368), .QTFCLK( ), .Q(cRet[11]));
Q_MX02 U741 ( .S(n1375), .A0(ctrlW[12]), .A1(cmdCnt[4]), .Z(n1367));
Q_FDP0UA U742 ( .D(n1367), .QTFCLK( ), .Q(cRet[12]));
Q_MX02 U743 ( .S(n1375), .A0(ctrlW[13]), .A1(cmdCnt[5]), .Z(n1366));
Q_FDP0UA U744 ( .D(n1366), .QTFCLK( ), .Q(cRet[13]));
Q_MX02 U745 ( .S(n1375), .A0(ctrlW[14]), .A1(cmdCnt[6]), .Z(n1365));
Q_FDP0UA U746 ( .D(n1365), .QTFCLK( ), .Q(cRet[14]));
Q_MX02 U747 ( .S(n1375), .A0(ctrlW[15]), .A1(cmdCnt[7]), .Z(n1364));
Q_FDP0UA U748 ( .D(n1364), .QTFCLK( ), .Q(cRet[15]));
Q_MX02 U749 ( .S(n1375), .A0(argTs[0]), .A1(ctrlR[64]), .Z(n1363));
Q_FDP0UA U750 ( .D(n1363), .QTFCLK( ), .Q(argTs[0]));
Q_MX02 U751 ( .S(n1375), .A0(argTs[1]), .A1(ctrlR[65]), .Z(n1362));
Q_FDP0UA U752 ( .D(n1362), .QTFCLK( ), .Q(argTs[1]));
Q_MX02 U753 ( .S(n1375), .A0(argTs[2]), .A1(ctrlR[66]), .Z(n1361));
Q_FDP0UA U754 ( .D(n1361), .QTFCLK( ), .Q(argTs[2]));
Q_MX02 U755 ( .S(n1375), .A0(argTs[3]), .A1(ctrlR[67]), .Z(n1360));
Q_FDP0UA U756 ( .D(n1360), .QTFCLK( ), .Q(argTs[3]));
Q_MX02 U757 ( .S(n1375), .A0(argTs[4]), .A1(ctrlR[68]), .Z(n1359));
Q_FDP0UA U758 ( .D(n1359), .QTFCLK( ), .Q(argTs[4]));
Q_MX02 U759 ( .S(n1375), .A0(argTs[5]), .A1(ctrlR[69]), .Z(n1358));
Q_FDP0UA U760 ( .D(n1358), .QTFCLK( ), .Q(argTs[5]));
Q_MX02 U761 ( .S(n1375), .A0(argTs[6]), .A1(ctrlR[70]), .Z(n1357));
Q_FDP0UA U762 ( .D(n1357), .QTFCLK( ), .Q(argTs[6]));
Q_MX02 U763 ( .S(n1375), .A0(argTs[7]), .A1(ctrlR[71]), .Z(n1356));
Q_FDP0UA U764 ( .D(n1356), .QTFCLK( ), .Q(argTs[7]));
Q_MX02 U765 ( .S(n1375), .A0(argTs[8]), .A1(ctrlR[72]), .Z(n1355));
Q_FDP0UA U766 ( .D(n1355), .QTFCLK( ), .Q(argTs[8]));
Q_MX02 U767 ( .S(n1375), .A0(argTs[9]), .A1(ctrlR[73]), .Z(n1354));
Q_FDP0UA U768 ( .D(n1354), .QTFCLK( ), .Q(argTs[9]));
Q_MX02 U769 ( .S(n1375), .A0(argTs[10]), .A1(ctrlR[74]), .Z(n1353));
Q_FDP0UA U770 ( .D(n1353), .QTFCLK( ), .Q(argTs[10]));
Q_MX02 U771 ( .S(n1375), .A0(argTs[11]), .A1(ctrlR[75]), .Z(n1352));
Q_FDP0UA U772 ( .D(n1352), .QTFCLK( ), .Q(argTs[11]));
Q_MX02 U773 ( .S(n1375), .A0(argTs[12]), .A1(ctrlR[76]), .Z(n1351));
Q_FDP0UA U774 ( .D(n1351), .QTFCLK( ), .Q(argTs[12]));
Q_MX02 U775 ( .S(n1375), .A0(argTs[13]), .A1(ctrlR[77]), .Z(n1350));
Q_FDP0UA U776 ( .D(n1350), .QTFCLK( ), .Q(argTs[13]));
Q_MX02 U777 ( .S(n1375), .A0(argTs[14]), .A1(ctrlR[78]), .Z(n1349));
Q_FDP0UA U778 ( .D(n1349), .QTFCLK( ), .Q(argTs[14]));
Q_MX02 U779 ( .S(n1375), .A0(argTs[15]), .A1(ctrlR[79]), .Z(n1348));
Q_FDP0UA U780 ( .D(n1348), .QTFCLK( ), .Q(argTs[15]));
Q_MX02 U781 ( .S(n1375), .A0(argTs[16]), .A1(ctrlR[80]), .Z(n1347));
Q_FDP0UA U782 ( .D(n1347), .QTFCLK( ), .Q(argTs[16]));
Q_MX02 U783 ( .S(n1375), .A0(argTs[17]), .A1(ctrlR[81]), .Z(n1346));
Q_FDP0UA U784 ( .D(n1346), .QTFCLK( ), .Q(argTs[17]));
Q_MX02 U785 ( .S(n1375), .A0(argTs[18]), .A1(ctrlR[82]), .Z(n1345));
Q_FDP0UA U786 ( .D(n1345), .QTFCLK( ), .Q(argTs[18]));
Q_MX02 U787 ( .S(n1375), .A0(argTs[19]), .A1(ctrlR[83]), .Z(n1344));
Q_FDP0UA U788 ( .D(n1344), .QTFCLK( ), .Q(argTs[19]));
Q_MX02 U789 ( .S(n1375), .A0(argTs[20]), .A1(ctrlR[84]), .Z(n1343));
Q_FDP0UA U790 ( .D(n1343), .QTFCLK( ), .Q(argTs[20]));
Q_MX02 U791 ( .S(n1375), .A0(argTs[21]), .A1(ctrlR[85]), .Z(n1342));
Q_FDP0UA U792 ( .D(n1342), .QTFCLK( ), .Q(argTs[21]));
Q_MX02 U793 ( .S(n1375), .A0(argTs[22]), .A1(ctrlR[86]), .Z(n1341));
Q_FDP0UA U794 ( .D(n1341), .QTFCLK( ), .Q(argTs[22]));
Q_MX02 U795 ( .S(n1375), .A0(argTs[23]), .A1(ctrlR[87]), .Z(n1340));
Q_FDP0UA U796 ( .D(n1340), .QTFCLK( ), .Q(argTs[23]));
Q_MX02 U797 ( .S(n1375), .A0(argTs[24]), .A1(ctrlR[88]), .Z(n1339));
Q_FDP0UA U798 ( .D(n1339), .QTFCLK( ), .Q(argTs[24]));
Q_MX02 U799 ( .S(n1375), .A0(argTs[25]), .A1(ctrlR[89]), .Z(n1338));
Q_FDP0UA U800 ( .D(n1338), .QTFCLK( ), .Q(argTs[25]));
Q_MX02 U801 ( .S(n1375), .A0(argTs[26]), .A1(ctrlR[90]), .Z(n1337));
Q_FDP0UA U802 ( .D(n1337), .QTFCLK( ), .Q(argTs[26]));
Q_MX02 U803 ( .S(n1375), .A0(argTs[27]), .A1(ctrlR[91]), .Z(n1336));
Q_FDP0UA U804 ( .D(n1336), .QTFCLK( ), .Q(argTs[27]));
Q_MX02 U805 ( .S(n1375), .A0(argTs[28]), .A1(ctrlR[92]), .Z(n1335));
Q_FDP0UA U806 ( .D(n1335), .QTFCLK( ), .Q(argTs[28]));
Q_MX02 U807 ( .S(n1375), .A0(argTs[29]), .A1(ctrlR[93]), .Z(n1334));
Q_FDP0UA U808 ( .D(n1334), .QTFCLK( ), .Q(argTs[29]));
Q_MX02 U809 ( .S(n1375), .A0(argTs[30]), .A1(ctrlR[94]), .Z(n1333));
Q_FDP0UA U810 ( .D(n1333), .QTFCLK( ), .Q(argTs[30]));
Q_MX02 U811 ( .S(n1375), .A0(argTs[31]), .A1(ctrlR[95]), .Z(n1332));
Q_FDP0UA U812 ( .D(n1332), .QTFCLK( ), .Q(argTs[31]));
Q_MX02 U813 ( .S(n1375), .A0(argTs[32]), .A1(ctrlR[96]), .Z(n1331));
Q_FDP0UA U814 ( .D(n1331), .QTFCLK( ), .Q(argTs[32]));
Q_MX02 U815 ( .S(n1375), .A0(argTs[33]), .A1(ctrlR[97]), .Z(n1330));
Q_FDP0UA U816 ( .D(n1330), .QTFCLK( ), .Q(argTs[33]));
Q_MX02 U817 ( .S(n1375), .A0(argTs[34]), .A1(ctrlR[98]), .Z(n1329));
Q_FDP0UA U818 ( .D(n1329), .QTFCLK( ), .Q(argTs[34]));
Q_MX02 U819 ( .S(n1375), .A0(argTs[35]), .A1(ctrlR[99]), .Z(n1328));
Q_FDP0UA U820 ( .D(n1328), .QTFCLK( ), .Q(argTs[35]));
Q_MX02 U821 ( .S(n1375), .A0(argTs[36]), .A1(ctrlR[100]), .Z(n1327));
Q_FDP0UA U822 ( .D(n1327), .QTFCLK( ), .Q(argTs[36]));
Q_MX02 U823 ( .S(n1375), .A0(argTs[37]), .A1(ctrlR[101]), .Z(n1326));
Q_FDP0UA U824 ( .D(n1326), .QTFCLK( ), .Q(argTs[37]));
Q_MX02 U825 ( .S(n1375), .A0(argTs[38]), .A1(ctrlR[102]), .Z(n1325));
Q_FDP0UA U826 ( .D(n1325), .QTFCLK( ), .Q(argTs[38]));
Q_MX02 U827 ( .S(n1375), .A0(argTs[39]), .A1(ctrlR[103]), .Z(n1324));
Q_FDP0UA U828 ( .D(n1324), .QTFCLK( ), .Q(argTs[39]));
Q_MX02 U829 ( .S(n1375), .A0(argTs[40]), .A1(ctrlR[104]), .Z(n1323));
Q_FDP0UA U830 ( .D(n1323), .QTFCLK( ), .Q(argTs[40]));
Q_MX02 U831 ( .S(n1375), .A0(argTs[41]), .A1(ctrlR[105]), .Z(n1322));
Q_FDP0UA U832 ( .D(n1322), .QTFCLK( ), .Q(argTs[41]));
Q_MX02 U833 ( .S(n1375), .A0(argTs[42]), .A1(ctrlR[106]), .Z(n1321));
Q_FDP0UA U834 ( .D(n1321), .QTFCLK( ), .Q(argTs[42]));
Q_MX02 U835 ( .S(n1375), .A0(argTs[43]), .A1(ctrlR[107]), .Z(n1320));
Q_FDP0UA U836 ( .D(n1320), .QTFCLK( ), .Q(argTs[43]));
Q_MX02 U837 ( .S(n1375), .A0(argTs[44]), .A1(ctrlR[108]), .Z(n1319));
Q_FDP0UA U838 ( .D(n1319), .QTFCLK( ), .Q(argTs[44]));
Q_MX02 U839 ( .S(n1375), .A0(argTs[45]), .A1(ctrlR[109]), .Z(n1318));
Q_FDP0UA U840 ( .D(n1318), .QTFCLK( ), .Q(argTs[45]));
Q_MX02 U841 ( .S(n1375), .A0(argTs[46]), .A1(ctrlR[110]), .Z(n1317));
Q_FDP0UA U842 ( .D(n1317), .QTFCLK( ), .Q(argTs[46]));
Q_MX02 U843 ( .S(n1375), .A0(argTs[47]), .A1(ctrlR[111]), .Z(n1316));
Q_FDP0UA U844 ( .D(n1316), .QTFCLK( ), .Q(argTs[47]));
Q_MX02 U845 ( .S(n1375), .A0(argTs[48]), .A1(ctrlR[112]), .Z(n1315));
Q_FDP0UA U846 ( .D(n1315), .QTFCLK( ), .Q(argTs[48]));
Q_MX02 U847 ( .S(n1375), .A0(argTs[49]), .A1(ctrlR[113]), .Z(n1314));
Q_FDP0UA U848 ( .D(n1314), .QTFCLK( ), .Q(argTs[49]));
Q_MX02 U849 ( .S(n1375), .A0(argTs[50]), .A1(ctrlR[114]), .Z(n1313));
Q_FDP0UA U850 ( .D(n1313), .QTFCLK( ), .Q(argTs[50]));
Q_MX02 U851 ( .S(n1375), .A0(argTs[51]), .A1(ctrlR[115]), .Z(n1312));
Q_FDP0UA U852 ( .D(n1312), .QTFCLK( ), .Q(argTs[51]));
Q_MX02 U853 ( .S(n1375), .A0(argTs[52]), .A1(ctrlR[116]), .Z(n1311));
Q_FDP0UA U854 ( .D(n1311), .QTFCLK( ), .Q(argTs[52]));
Q_MX02 U855 ( .S(n1375), .A0(argTs[53]), .A1(ctrlR[117]), .Z(n1310));
Q_FDP0UA U856 ( .D(n1310), .QTFCLK( ), .Q(argTs[53]));
Q_MX02 U857 ( .S(n1375), .A0(argTs[54]), .A1(ctrlR[118]), .Z(n1309));
Q_FDP0UA U858 ( .D(n1309), .QTFCLK( ), .Q(argTs[54]));
Q_MX02 U859 ( .S(n1375), .A0(argTs[55]), .A1(ctrlR[119]), .Z(n1308));
Q_FDP0UA U860 ( .D(n1308), .QTFCLK( ), .Q(argTs[55]));
Q_MX02 U861 ( .S(n1375), .A0(argTs[56]), .A1(ctrlR[120]), .Z(n1307));
Q_FDP0UA U862 ( .D(n1307), .QTFCLK( ), .Q(argTs[56]));
Q_MX02 U863 ( .S(n1375), .A0(argTs[57]), .A1(ctrlR[121]), .Z(n1306));
Q_FDP0UA U864 ( .D(n1306), .QTFCLK( ), .Q(argTs[57]));
Q_MX02 U865 ( .S(n1375), .A0(argTs[58]), .A1(ctrlR[122]), .Z(n1305));
Q_FDP0UA U866 ( .D(n1305), .QTFCLK( ), .Q(argTs[58]));
Q_MX02 U867 ( .S(n1375), .A0(argTs[59]), .A1(ctrlR[123]), .Z(n1304));
Q_FDP0UA U868 ( .D(n1304), .QTFCLK( ), .Q(argTs[59]));
Q_MX02 U869 ( .S(n1375), .A0(argTs[60]), .A1(ctrlR[124]), .Z(n1303));
Q_FDP0UA U870 ( .D(n1303), .QTFCLK( ), .Q(argTs[60]));
Q_MX02 U871 ( .S(n1375), .A0(argTs[61]), .A1(ctrlR[125]), .Z(n1302));
Q_FDP0UA U872 ( .D(n1302), .QTFCLK( ), .Q(argTs[61]));
Q_MX02 U873 ( .S(n1375), .A0(argTs[62]), .A1(ctrlR[126]), .Z(n1301));
Q_FDP0UA U874 ( .D(n1301), .QTFCLK( ), .Q(argTs[62]));
Q_MX02 U875 ( .S(n1375), .A0(argTs[63]), .A1(ctrlR[127]), .Z(n1300));
Q_FDP0UA U876 ( .D(n1300), .QTFCLK( ), .Q(argTs[63]));
Q_MX02 U877 ( .S(n1375), .A0(argTc[0]), .A1(ctrlR[0]), .Z(n1299));
Q_FDP0UA U878 ( .D(n1299), .QTFCLK( ), .Q(argTc[0]));
Q_MX02 U879 ( .S(n1375), .A0(argTc[1]), .A1(ctrlR[1]), .Z(n1298));
Q_FDP0UA U880 ( .D(n1298), .QTFCLK( ), .Q(argTc[1]));
Q_MX02 U881 ( .S(n1375), .A0(argTc[2]), .A1(ctrlR[2]), .Z(n1297));
Q_FDP0UA U882 ( .D(n1297), .QTFCLK( ), .Q(argTc[2]));
Q_MX02 U883 ( .S(n1375), .A0(argTc[3]), .A1(ctrlR[3]), .Z(n1296));
Q_FDP0UA U884 ( .D(n1296), .QTFCLK( ), .Q(argTc[3]));
Q_MX02 U885 ( .S(n1375), .A0(argTc[4]), .A1(ctrlR[4]), .Z(n1295));
Q_FDP0UA U886 ( .D(n1295), .QTFCLK( ), .Q(argTc[4]));
Q_MX02 U887 ( .S(n1375), .A0(argTc[5]), .A1(ctrlR[5]), .Z(n1294));
Q_FDP0UA U888 ( .D(n1294), .QTFCLK( ), .Q(argTc[5]));
Q_MX02 U889 ( .S(n1375), .A0(argTc[6]), .A1(ctrlR[6]), .Z(n1293));
Q_FDP0UA U890 ( .D(n1293), .QTFCLK( ), .Q(argTc[6]));
Q_MX02 U891 ( .S(n1375), .A0(argTc[7]), .A1(ctrlR[7]), .Z(n1292));
Q_FDP0UA U892 ( .D(n1292), .QTFCLK( ), .Q(argTc[7]));
Q_MX02 U893 ( .S(n1375), .A0(argTc[8]), .A1(ctrlR[8]), .Z(n1291));
Q_FDP0UA U894 ( .D(n1291), .QTFCLK( ), .Q(argTc[8]));
Q_MX02 U895 ( .S(n1375), .A0(argTc[9]), .A1(ctrlR[9]), .Z(n1290));
Q_FDP0UA U896 ( .D(n1290), .QTFCLK( ), .Q(argTc[9]));
Q_MX02 U897 ( .S(n1375), .A0(argTc[10]), .A1(ctrlR[10]), .Z(n1289));
Q_FDP0UA U898 ( .D(n1289), .QTFCLK( ), .Q(argTc[10]));
Q_MX02 U899 ( .S(n1375), .A0(argTc[11]), .A1(ctrlR[11]), .Z(n1288));
Q_FDP0UA U900 ( .D(n1288), .QTFCLK( ), .Q(argTc[11]));
Q_MX02 U901 ( .S(n1375), .A0(argTc[12]), .A1(ctrlR[12]), .Z(n1287));
Q_FDP0UA U902 ( .D(n1287), .QTFCLK( ), .Q(argTc[12]));
Q_MX02 U903 ( .S(n1375), .A0(argTc[13]), .A1(ctrlR[13]), .Z(n1286));
Q_FDP0UA U904 ( .D(n1286), .QTFCLK( ), .Q(argTc[13]));
Q_MX02 U905 ( .S(n1375), .A0(argTc[14]), .A1(ctrlR[14]), .Z(n1285));
Q_FDP0UA U906 ( .D(n1285), .QTFCLK( ), .Q(argTc[14]));
Q_MX02 U907 ( .S(n1375), .A0(argTc[15]), .A1(ctrlR[15]), .Z(n1284));
Q_FDP0UA U908 ( .D(n1284), .QTFCLK( ), .Q(argTc[15]));
Q_MX02 U909 ( .S(n1375), .A0(argTc[16]), .A1(ctrlR[16]), .Z(n1283));
Q_FDP0UA U910 ( .D(n1283), .QTFCLK( ), .Q(argTc[16]));
Q_MX02 U911 ( .S(n1375), .A0(argTc[17]), .A1(ctrlR[17]), .Z(n1282));
Q_FDP0UA U912 ( .D(n1282), .QTFCLK( ), .Q(argTc[17]));
Q_MX02 U913 ( .S(n1375), .A0(argTc[18]), .A1(ctrlR[18]), .Z(n1281));
Q_FDP0UA U914 ( .D(n1281), .QTFCLK( ), .Q(argTc[18]));
Q_MX02 U915 ( .S(n1375), .A0(argTc[19]), .A1(ctrlR[19]), .Z(n1280));
Q_FDP0UA U916 ( .D(n1280), .QTFCLK( ), .Q(argTc[19]));
Q_MX02 U917 ( .S(n1375), .A0(argTc[20]), .A1(ctrlR[20]), .Z(n1279));
Q_FDP0UA U918 ( .D(n1279), .QTFCLK( ), .Q(argTc[20]));
Q_MX02 U919 ( .S(n1375), .A0(argTc[21]), .A1(ctrlR[21]), .Z(n1278));
Q_FDP0UA U920 ( .D(n1278), .QTFCLK( ), .Q(argTc[21]));
Q_MX02 U921 ( .S(n1375), .A0(argTc[22]), .A1(ctrlR[22]), .Z(n1277));
Q_FDP0UA U922 ( .D(n1277), .QTFCLK( ), .Q(argTc[22]));
Q_MX02 U923 ( .S(n1375), .A0(argTc[23]), .A1(ctrlR[23]), .Z(n1276));
Q_FDP0UA U924 ( .D(n1276), .QTFCLK( ), .Q(argTc[23]));
Q_MX02 U925 ( .S(n1375), .A0(argTc[24]), .A1(ctrlR[24]), .Z(n1275));
Q_FDP0UA U926 ( .D(n1275), .QTFCLK( ), .Q(argTc[24]));
Q_MX02 U927 ( .S(n1375), .A0(argTc[25]), .A1(ctrlR[25]), .Z(n1274));
Q_FDP0UA U928 ( .D(n1274), .QTFCLK( ), .Q(argTc[25]));
Q_MX02 U929 ( .S(n1375), .A0(argTc[26]), .A1(ctrlR[26]), .Z(n1273));
Q_FDP0UA U930 ( .D(n1273), .QTFCLK( ), .Q(argTc[26]));
Q_MX02 U931 ( .S(n1375), .A0(argTc[27]), .A1(ctrlR[27]), .Z(n1272));
Q_FDP0UA U932 ( .D(n1272), .QTFCLK( ), .Q(argTc[27]));
Q_MX02 U933 ( .S(n1375), .A0(argTc[28]), .A1(ctrlR[28]), .Z(n1271));
Q_FDP0UA U934 ( .D(n1271), .QTFCLK( ), .Q(argTc[28]));
Q_MX02 U935 ( .S(n1375), .A0(argTc[29]), .A1(ctrlR[29]), .Z(n1270));
Q_FDP0UA U936 ( .D(n1270), .QTFCLK( ), .Q(argTc[29]));
Q_MX02 U937 ( .S(n1375), .A0(argTc[30]), .A1(ctrlR[30]), .Z(n1269));
Q_FDP0UA U938 ( .D(n1269), .QTFCLK( ), .Q(argTc[30]));
Q_MX02 U939 ( .S(n1375), .A0(argTc[31]), .A1(ctrlR[31]), .Z(n1268));
Q_FDP0UA U940 ( .D(n1268), .QTFCLK( ), .Q(argTc[31]));
Q_MX02 U941 ( .S(n1375), .A0(argTc[32]), .A1(ctrlR[32]), .Z(n1267));
Q_FDP0UA U942 ( .D(n1267), .QTFCLK( ), .Q(argTc[32]));
Q_MX02 U943 ( .S(n1375), .A0(argTc[33]), .A1(ctrlR[33]), .Z(n1266));
Q_FDP0UA U944 ( .D(n1266), .QTFCLK( ), .Q(argTc[33]));
Q_MX02 U945 ( .S(n1375), .A0(argTc[34]), .A1(ctrlR[34]), .Z(n1265));
Q_FDP0UA U946 ( .D(n1265), .QTFCLK( ), .Q(argTc[34]));
Q_MX02 U947 ( .S(n1375), .A0(argTc[35]), .A1(ctrlR[35]), .Z(n1264));
Q_FDP0UA U948 ( .D(n1264), .QTFCLK( ), .Q(argTc[35]));
Q_MX02 U949 ( .S(n1375), .A0(argTc[36]), .A1(ctrlR[36]), .Z(n1263));
Q_FDP0UA U950 ( .D(n1263), .QTFCLK( ), .Q(argTc[36]));
Q_MX02 U951 ( .S(n1375), .A0(argTc[37]), .A1(ctrlR[37]), .Z(n1262));
Q_FDP0UA U952 ( .D(n1262), .QTFCLK( ), .Q(argTc[37]));
Q_MX02 U953 ( .S(n1375), .A0(argTc[38]), .A1(ctrlR[38]), .Z(n1261));
Q_FDP0UA U954 ( .D(n1261), .QTFCLK( ), .Q(argTc[38]));
Q_MX02 U955 ( .S(n1375), .A0(argTc[39]), .A1(ctrlR[39]), .Z(n1260));
Q_FDP0UA U956 ( .D(n1260), .QTFCLK( ), .Q(argTc[39]));
Q_MX02 U957 ( .S(n1375), .A0(argTc[40]), .A1(ctrlR[40]), .Z(n1259));
Q_FDP0UA U958 ( .D(n1259), .QTFCLK( ), .Q(argTc[40]));
Q_MX02 U959 ( .S(n1375), .A0(argTc[41]), .A1(ctrlR[41]), .Z(n1258));
Q_FDP0UA U960 ( .D(n1258), .QTFCLK( ), .Q(argTc[41]));
Q_MX02 U961 ( .S(n1375), .A0(argTc[42]), .A1(ctrlR[42]), .Z(n1257));
Q_FDP0UA U962 ( .D(n1257), .QTFCLK( ), .Q(argTc[42]));
Q_MX02 U963 ( .S(n1375), .A0(argTc[43]), .A1(ctrlR[43]), .Z(n1256));
Q_FDP0UA U964 ( .D(n1256), .QTFCLK( ), .Q(argTc[43]));
Q_MX02 U965 ( .S(n1375), .A0(argTc[44]), .A1(ctrlR[44]), .Z(n1255));
Q_FDP0UA U966 ( .D(n1255), .QTFCLK( ), .Q(argTc[44]));
Q_MX02 U967 ( .S(n1375), .A0(argTc[45]), .A1(ctrlR[45]), .Z(n1254));
Q_FDP0UA U968 ( .D(n1254), .QTFCLK( ), .Q(argTc[45]));
Q_MX02 U969 ( .S(n1375), .A0(argTc[46]), .A1(ctrlR[46]), .Z(n1253));
Q_FDP0UA U970 ( .D(n1253), .QTFCLK( ), .Q(argTc[46]));
Q_MX02 U971 ( .S(n1375), .A0(argTc[47]), .A1(ctrlR[47]), .Z(n1252));
Q_FDP0UA U972 ( .D(n1252), .QTFCLK( ), .Q(argTc[47]));
Q_MX02 U973 ( .S(n1375), .A0(argTc[48]), .A1(ctrlR[48]), .Z(n1251));
Q_FDP0UA U974 ( .D(n1251), .QTFCLK( ), .Q(argTc[48]));
Q_MX02 U975 ( .S(n1375), .A0(argTc[49]), .A1(ctrlR[49]), .Z(n1250));
Q_FDP0UA U976 ( .D(n1250), .QTFCLK( ), .Q(argTc[49]));
Q_MX02 U977 ( .S(n1375), .A0(argTc[50]), .A1(ctrlR[50]), .Z(n1249));
Q_FDP0UA U978 ( .D(n1249), .QTFCLK( ), .Q(argTc[50]));
Q_MX02 U979 ( .S(n1375), .A0(argTc[51]), .A1(ctrlR[51]), .Z(n1248));
Q_FDP0UA U980 ( .D(n1248), .QTFCLK( ), .Q(argTc[51]));
Q_MX02 U981 ( .S(n1375), .A0(argTc[52]), .A1(ctrlR[52]), .Z(n1247));
Q_FDP0UA U982 ( .D(n1247), .QTFCLK( ), .Q(argTc[52]));
Q_MX02 U983 ( .S(n1375), .A0(argTc[53]), .A1(ctrlR[53]), .Z(n1246));
Q_FDP0UA U984 ( .D(n1246), .QTFCLK( ), .Q(argTc[53]));
Q_MX02 U985 ( .S(n1375), .A0(argTc[54]), .A1(ctrlR[54]), .Z(n1245));
Q_FDP0UA U986 ( .D(n1245), .QTFCLK( ), .Q(argTc[54]));
Q_MX02 U987 ( .S(n1375), .A0(argTc[55]), .A1(ctrlR[55]), .Z(n1244));
Q_FDP0UA U988 ( .D(n1244), .QTFCLK( ), .Q(argTc[55]));
Q_MX02 U989 ( .S(n1375), .A0(argTc[56]), .A1(ctrlR[56]), .Z(n1243));
Q_FDP0UA U990 ( .D(n1243), .QTFCLK( ), .Q(argTc[56]));
Q_MX02 U991 ( .S(n1375), .A0(argTc[57]), .A1(ctrlR[57]), .Z(n1242));
Q_FDP0UA U992 ( .D(n1242), .QTFCLK( ), .Q(argTc[57]));
Q_MX02 U993 ( .S(n1375), .A0(argTc[58]), .A1(ctrlR[58]), .Z(n1241));
Q_FDP0UA U994 ( .D(n1241), .QTFCLK( ), .Q(argTc[58]));
Q_MX02 U995 ( .S(n1375), .A0(argTc[59]), .A1(ctrlR[59]), .Z(n1240));
Q_FDP0UA U996 ( .D(n1240), .QTFCLK( ), .Q(argTc[59]));
Q_MX02 U997 ( .S(n1375), .A0(argTc[60]), .A1(ctrlR[60]), .Z(n1239));
Q_FDP0UA U998 ( .D(n1239), .QTFCLK( ), .Q(argTc[60]));
Q_MX02 U999 ( .S(n1375), .A0(argTc[61]), .A1(ctrlR[61]), .Z(n1238));
Q_FDP0UA U1000 ( .D(n1238), .QTFCLK( ), .Q(argTc[61]));
Q_MX02 U1001 ( .S(n1375), .A0(argTc[62]), .A1(ctrlR[62]), .Z(n1237));
Q_FDP0UA U1002 ( .D(n1237), .QTFCLK( ), .Q(argTc[62]));
Q_MX02 U1003 ( .S(n1375), .A0(argTc[63]), .A1(ctrlR[63]), .Z(n1236));
Q_FDP0UA U1004 ( .D(n1236), .QTFCLK( ), .Q(argTc[63]));
Q_MX02 U1005 ( .S(n1375), .A0(cmdCntP[0]), .A1(cmdCnt[0]), .Z(n1235));
Q_FDP0UA U1006 ( .D(n1235), .QTFCLK( ), .Q(cmdCntP[0]));
Q_MX02 U1007 ( .S(n1375), .A0(cmdCntP[1]), .A1(cmdCnt[1]), .Z(n1234));
Q_FDP0UA U1008 ( .D(n1234), .QTFCLK( ), .Q(cmdCntP[1]));
Q_MX02 U1009 ( .S(n1375), .A0(cmdCntP[2]), .A1(cmdCnt[2]), .Z(n1233));
Q_FDP0UA U1010 ( .D(n1233), .QTFCLK( ), .Q(cmdCntP[2]));
Q_MX02 U1011 ( .S(n1375), .A0(cmdCntP[3]), .A1(cmdCnt[3]), .Z(n1232));
Q_FDP0UA U1012 ( .D(n1232), .QTFCLK( ), .Q(cmdCntP[3]));
Q_MX02 U1013 ( .S(n1375), .A0(cmdCntP[4]), .A1(cmdCnt[4]), .Z(n1231));
Q_FDP0UA U1014 ( .D(n1231), .QTFCLK( ), .Q(cmdCntP[4]));
Q_MX02 U1015 ( .S(n1375), .A0(cmdCntP[5]), .A1(cmdCnt[5]), .Z(n1230));
Q_FDP0UA U1016 ( .D(n1230), .QTFCLK( ), .Q(cmdCntP[5]));
Q_MX02 U1017 ( .S(n1375), .A0(cmdCntP[6]), .A1(cmdCnt[6]), .Z(n1229));
Q_FDP0UA U1018 ( .D(n1229), .QTFCLK( ), .Q(cmdCntP[6]));
Q_MX02 U1019 ( .S(n1375), .A0(cmdCntP[7]), .A1(cmdCnt[7]), .Z(n1228));
Q_FDP0UA U1020 ( .D(n1228), .QTFCLK( ), .Q(cmdCntP[7]));
Q_MX02 U1021 ( .S(n1375), .A0(cmdR[0]), .A1(cmdC[0]), .Z(n1227));
Q_FDP0UA U1022 ( .D(n1227), .QTFCLK( ), .Q(cmdR[0]));
Q_MX02 U1023 ( .S(n1375), .A0(cmdR[1]), .A1(cmdC[1]), .Z(n1226));
Q_FDP0UA U1024 ( .D(n1226), .QTFCLK( ), .Q(cmdR[1]));
Q_MX02 U1025 ( .S(n1375), .A0(cmdR[2]), .A1(cmdC[2]), .Z(n1225));
Q_FDP0UA U1026 ( .D(n1225), .QTFCLK( ), .Q(cmdR[2]));
Q_MX02 U1027 ( .S(n1375), .A0(cmdR[3]), .A1(cmdC[3]), .Z(n1224));
Q_FDP0UA U1028 ( .D(n1224), .QTFCLK( ), .Q(cmdR[3]));
Q_MX02 U1029 ( .S(n1375), .A0(cmdR[4]), .A1(cmdC[4]), .Z(n1223));
Q_FDP0UA U1030 ( .D(n1223), .QTFCLK( ), .Q(cmdR[4]));
Q_MX02 U1031 ( .S(n1375), .A0(cmdR[5]), .A1(cmdC[5]), .Z(n1222));
Q_FDP0UA U1032 ( .D(n1222), .QTFCLK( ), .Q(cmdR[5]));
Q_MX02 U1033 ( .S(n1375), .A0(cmdR[6]), .A1(cmdC[6]), .Z(n1221));
Q_FDP0UA U1034 ( .D(n1221), .QTFCLK( ), .Q(cmdR[6]));
Q_MX02 U1035 ( .S(n1375), .A0(cmdR[7]), .A1(cmdC[7]), .Z(n1220));
Q_FDP0UA U1036 ( .D(n1220), .QTFCLK( ), .Q(cmdR[7]));
Q_FDP0UA U1037 ( .D(busyCnt[6]), .QTFCLK( ), .Q(busyCnt[7]));
Q_FDP0UA U1038 ( .D(busyCnt[5]), .QTFCLK( ), .Q(busyCnt[6]));
Q_FDP0UA U1039 ( .D(busyCnt[4]), .QTFCLK( ), .Q(busyCnt[5]));
Q_FDP0UA U1040 ( .D(busyCnt[3]), .QTFCLK( ), .Q(busyCnt[4]));
Q_FDP0UA U1041 ( .D(busyCnt[2]), .QTFCLK( ), .Q(busyCnt[3]));
Q_FDP0UA U1042 ( .D(busyCnt[1]), .QTFCLK( ), .Q(busyCnt[2]));
Q_FDP0UA U1043 ( .D(busyCnt[0]), .QTFCLK( ), .Q(busyCnt[1]));
Q_FDP0UA U1044 ( .D(newCtrl), .QTFCLK( ), .Q(busyCnt[0]));
Q_FDP0UA U1045 ( .D(ctrlW[127]), .QTFCLK( ), .Q(ecmTsP[63]));
Q_FDP0UA U1046 ( .D(ctrlW[126]), .QTFCLK( ), .Q(ecmTsP[62]));
Q_FDP0UA U1047 ( .D(ctrlW[125]), .QTFCLK( ), .Q(ecmTsP[61]));
Q_FDP0UA U1048 ( .D(ctrlW[124]), .QTFCLK( ), .Q(ecmTsP[60]));
Q_FDP0UA U1049 ( .D(ctrlW[123]), .QTFCLK( ), .Q(ecmTsP[59]));
Q_FDP0UA U1050 ( .D(ctrlW[122]), .QTFCLK( ), .Q(ecmTsP[58]));
Q_FDP0UA U1051 ( .D(ctrlW[121]), .QTFCLK( ), .Q(ecmTsP[57]));
Q_FDP0UA U1052 ( .D(ctrlW[120]), .QTFCLK( ), .Q(ecmTsP[56]));
Q_FDP0UA U1053 ( .D(ctrlW[119]), .QTFCLK( ), .Q(ecmTsP[55]));
Q_FDP0UA U1054 ( .D(ctrlW[118]), .QTFCLK( ), .Q(ecmTsP[54]));
Q_FDP0UA U1055 ( .D(ctrlW[117]), .QTFCLK( ), .Q(ecmTsP[53]));
Q_FDP0UA U1056 ( .D(ctrlW[116]), .QTFCLK( ), .Q(ecmTsP[52]));
Q_FDP0UA U1057 ( .D(ctrlW[115]), .QTFCLK( ), .Q(ecmTsP[51]));
Q_FDP0UA U1058 ( .D(ctrlW[114]), .QTFCLK( ), .Q(ecmTsP[50]));
Q_FDP0UA U1059 ( .D(ctrlW[113]), .QTFCLK( ), .Q(ecmTsP[49]));
Q_FDP0UA U1060 ( .D(ctrlW[112]), .QTFCLK( ), .Q(ecmTsP[48]));
Q_FDP0UA U1061 ( .D(ctrlW[111]), .QTFCLK( ), .Q(ecmTsP[47]));
Q_FDP0UA U1062 ( .D(ctrlW[110]), .QTFCLK( ), .Q(ecmTsP[46]));
Q_FDP0UA U1063 ( .D(ctrlW[109]), .QTFCLK( ), .Q(ecmTsP[45]));
Q_FDP0UA U1064 ( .D(ctrlW[108]), .QTFCLK( ), .Q(ecmTsP[44]));
Q_FDP0UA U1065 ( .D(ctrlW[107]), .QTFCLK( ), .Q(ecmTsP[43]));
Q_FDP0UA U1066 ( .D(ctrlW[106]), .QTFCLK( ), .Q(ecmTsP[42]));
Q_FDP0UA U1067 ( .D(ctrlW[105]), .QTFCLK( ), .Q(ecmTsP[41]));
Q_FDP0UA U1068 ( .D(ctrlW[104]), .QTFCLK( ), .Q(ecmTsP[40]));
Q_FDP0UA U1069 ( .D(ctrlW[103]), .QTFCLK( ), .Q(ecmTsP[39]));
Q_FDP0UA U1070 ( .D(ctrlW[102]), .QTFCLK( ), .Q(ecmTsP[38]));
Q_FDP0UA U1071 ( .D(ctrlW[101]), .QTFCLK( ), .Q(ecmTsP[37]));
Q_FDP0UA U1072 ( .D(ctrlW[100]), .QTFCLK( ), .Q(ecmTsP[36]));
Q_FDP0UA U1073 ( .D(ctrlW[99]), .QTFCLK( ), .Q(ecmTsP[35]));
Q_FDP0UA U1074 ( .D(ctrlW[98]), .QTFCLK( ), .Q(ecmTsP[34]));
Q_FDP0UA U1075 ( .D(ctrlW[97]), .QTFCLK( ), .Q(ecmTsP[33]));
Q_FDP0UA U1076 ( .D(ctrlW[96]), .QTFCLK( ), .Q(ecmTsP[32]));
Q_FDP0UA U1077 ( .D(ctrlW[95]), .QTFCLK( ), .Q(ecmTsP[31]));
Q_FDP0UA U1078 ( .D(ctrlW[94]), .QTFCLK( ), .Q(ecmTsP[30]));
Q_FDP0UA U1079 ( .D(ctrlW[93]), .QTFCLK( ), .Q(ecmTsP[29]));
Q_FDP0UA U1080 ( .D(ctrlW[92]), .QTFCLK( ), .Q(ecmTsP[28]));
Q_FDP0UA U1081 ( .D(ctrlW[91]), .QTFCLK( ), .Q(ecmTsP[27]));
Q_FDP0UA U1082 ( .D(ctrlW[90]), .QTFCLK( ), .Q(ecmTsP[26]));
Q_FDP0UA U1083 ( .D(ctrlW[89]), .QTFCLK( ), .Q(ecmTsP[25]));
Q_FDP0UA U1084 ( .D(ctrlW[88]), .QTFCLK( ), .Q(ecmTsP[24]));
Q_FDP0UA U1085 ( .D(ctrlW[87]), .QTFCLK( ), .Q(ecmTsP[23]));
Q_FDP0UA U1086 ( .D(ctrlW[86]), .QTFCLK( ), .Q(ecmTsP[22]));
Q_FDP0UA U1087 ( .D(ctrlW[85]), .QTFCLK( ), .Q(ecmTsP[21]));
Q_FDP0UA U1088 ( .D(ctrlW[84]), .QTFCLK( ), .Q(ecmTsP[20]));
Q_FDP0UA U1089 ( .D(ctrlW[83]), .QTFCLK( ), .Q(ecmTsP[19]));
Q_FDP0UA U1090 ( .D(ctrlW[82]), .QTFCLK( ), .Q(ecmTsP[18]));
Q_FDP0UA U1091 ( .D(ctrlW[81]), .QTFCLK( ), .Q(ecmTsP[17]));
Q_FDP0UA U1092 ( .D(ctrlW[80]), .QTFCLK( ), .Q(ecmTsP[16]));
Q_FDP0UA U1093 ( .D(ctrlW[79]), .QTFCLK( ), .Q(ecmTsP[15]));
Q_FDP0UA U1094 ( .D(ctrlW[78]), .QTFCLK( ), .Q(ecmTsP[14]));
Q_FDP0UA U1095 ( .D(ctrlW[77]), .QTFCLK( ), .Q(ecmTsP[13]));
Q_FDP0UA U1096 ( .D(ctrlW[76]), .QTFCLK( ), .Q(ecmTsP[12]));
Q_FDP0UA U1097 ( .D(ctrlW[75]), .QTFCLK( ), .Q(ecmTsP[11]));
Q_FDP0UA U1098 ( .D(ctrlW[74]), .QTFCLK( ), .Q(ecmTsP[10]));
Q_FDP0UA U1099 ( .D(ctrlW[73]), .QTFCLK( ), .Q(ecmTsP[9]));
Q_FDP0UA U1100 ( .D(ctrlW[72]), .QTFCLK( ), .Q(ecmTsP[8]));
Q_FDP0UA U1101 ( .D(ctrlW[71]), .QTFCLK( ), .Q(ecmTsP[7]));
Q_FDP0UA U1102 ( .D(ctrlW[70]), .QTFCLK( ), .Q(ecmTsP[6]));
Q_FDP0UA U1103 ( .D(ctrlW[69]), .QTFCLK( ), .Q(ecmTsP[5]));
Q_FDP0UA U1104 ( .D(ctrlW[68]), .QTFCLK( ), .Q(ecmTsP[4]));
Q_FDP0UA U1105 ( .D(ctrlW[67]), .QTFCLK( ), .Q(ecmTsP[3]));
Q_FDP0UA U1106 ( .D(ctrlW[66]), .QTFCLK( ), .Q(ecmTsP[2]));
Q_FDP0UA U1107 ( .D(ctrlW[65]), .QTFCLK( ), .Q(ecmTsP[1]));
Q_FDP0UA U1108 ( .D(ctrlW[64]), .QTFCLK( ), .Q(ecmTsP[0]));
Q_FDP0UA U1109 ( .D(ctrlEv[1]), .QTFCLK( ), .Q(ctrlEvP[1]));
Q_FDP0UA U1110 ( .D(ctrlEv[0]), .QTFCLK( ), .Q(ctrlEvP[0]));
Q_FDP0UA U1111 ( .D(xcva_top.xc_top.sdlStopRply), .QTFCLK( ), .Q(sdlStopRply));
Q_XNR2 U1112 ( .A0(cmdCnt[0]), .A1(cmdCntP[0]), .Z(n1218));
Q_XNR2 U1113 ( .A0(cmdCnt[1]), .A1(cmdCntP[1]), .Z(n1217));
Q_XNR2 U1114 ( .A0(cmdCnt[2]), .A1(cmdCntP[2]), .Z(n1216));
Q_XNR2 U1115 ( .A0(cmdCnt[3]), .A1(cmdCntP[3]), .Z(n1215));
Q_XNR2 U1116 ( .A0(cmdCnt[4]), .A1(cmdCntP[4]), .Z(n1214));
Q_XNR2 U1117 ( .A0(cmdCnt[5]), .A1(cmdCntP[5]), .Z(n1213));
Q_XNR2 U1118 ( .A0(cmdCnt[6]), .A1(cmdCntP[6]), .Z(n1212));
Q_XNR2 U1119 ( .A0(cmdCnt[7]), .A1(cmdCntP[7]), .Z(n1211));
Q_AN03 U1120 ( .A0(n1211), .A1(n1212), .A2(n1213), .Z(n1210));
Q_AN03 U1121 ( .A0(n1214), .A1(n1215), .A2(n1216), .Z(n1209));
Q_AN03 U1122 ( .A0(n1217), .A1(n1218), .A2(n1210), .Z(n1208));
Q_AN02 U1123 ( .A0(n1209), .A1(n1208), .Z(n1207));
Q_INV U1124 ( .A(n1207), .Z(newCmd));
Q_XNR2 U1125 ( .A0(syncId[0]), .A1(syncIdP[0]), .Z(n1206));
Q_XNR2 U1126 ( .A0(syncId[1]), .A1(syncIdP[1]), .Z(n1205));
Q_XNR2 U1127 ( .A0(syncId[2]), .A1(syncIdP[2]), .Z(n1204));
Q_XNR2 U1128 ( .A0(syncId[3]), .A1(syncIdP[3]), .Z(n1203));
Q_XNR2 U1129 ( .A0(syncId[4]), .A1(syncIdP[4]), .Z(n1202));
Q_XNR2 U1130 ( .A0(syncId[5]), .A1(syncIdP[5]), .Z(n1201));
Q_XNR2 U1131 ( .A0(syncId[6]), .A1(syncIdP[6]), .Z(n1200));
Q_XNR2 U1132 ( .A0(syncId[7]), .A1(syncIdP[7]), .Z(n1199));
Q_AN03 U1133 ( .A0(n1199), .A1(n1200), .A2(n1201), .Z(n1198));
Q_AN03 U1134 ( .A0(n1202), .A1(n1203), .A2(n1204), .Z(n1197));
Q_AN03 U1135 ( .A0(n1205), .A1(n1206), .A2(n1198), .Z(n1196));
Q_AN02 U1136 ( .A0(n1197), .A1(n1196), .Z(n1195));
Q_INV U1137 ( .A(n1195), .Z(newSync));
Q_XOR2 U1138 ( .A0(ctrlEv[0]), .A1(ctrlEvP[0]), .Z(n1194));
Q_XOR2 U1139 ( .A0(ctrlEv[1]), .A1(ctrlEvP[1]), .Z(n1193));
Q_OR02 U1140 ( .A0(n1194), .A1(n1193), .Z(newCtrl));
Q_OR03 U1141 ( .A0(busyCnt[7]), .A1(busyCnt[6]), .A2(busyCnt[5]), .Z(n1192));
Q_OR03 U1142 ( .A0(busyCnt[4]), .A1(busyCnt[3]), .A2(busyCnt[2]), .Z(n1191));
Q_OR03 U1143 ( .A0(busyCnt[1]), .A1(busyCnt[0]), .A2(n1192), .Z(n1190));
Q_OR02 U1144 ( .A0(n1191), .A1(n1190), .Z(n1189));
Q_AN02 U1145 ( .A0(holdEcmBusy), .A1(n1395), .Z(n1188));
Q_OR03 U1146 ( .A0(newCtrl), .A1(n1189), .A2(n1188), .Z(busyOn));
Q_AD01HF U1147 ( .A0(ecmTsP[1]), .B0(ecmTsP[0]), .S(n1187), .CO(n1186));
Q_AD01HF U1148 ( .A0(ecmTsP[2]), .B0(n1186), .S(n1185), .CO(n1184));
Q_AD01HF U1149 ( .A0(ecmTsP[3]), .B0(n1184), .S(n1183), .CO(n1182));
Q_AD01HF U1150 ( .A0(ecmTsP[4]), .B0(n1182), .S(n1181), .CO(n1180));
Q_AD01HF U1151 ( .A0(ecmTsP[5]), .B0(n1180), .S(n1179), .CO(n1178));
Q_AD01HF U1152 ( .A0(ecmTsP[6]), .B0(n1178), .S(n1177), .CO(n1176));
Q_AD01HF U1153 ( .A0(ecmTsP[7]), .B0(n1176), .S(n1175), .CO(n1174));
Q_AD01HF U1154 ( .A0(ecmTsP[8]), .B0(n1174), .S(n1173), .CO(n1172));
Q_AD01HF U1155 ( .A0(ecmTsP[9]), .B0(n1172), .S(n1171), .CO(n1170));
Q_AD01HF U1156 ( .A0(ecmTsP[10]), .B0(n1170), .S(n1169), .CO(n1168));
Q_AD01HF U1157 ( .A0(ecmTsP[11]), .B0(n1168), .S(n1167), .CO(n1166));
Q_AD01HF U1158 ( .A0(ecmTsP[12]), .B0(n1166), .S(n1165), .CO(n1164));
Q_AD01HF U1159 ( .A0(ecmTsP[13]), .B0(n1164), .S(n1163), .CO(n1162));
Q_AD01HF U1160 ( .A0(ecmTsP[14]), .B0(n1162), .S(n1161), .CO(n1160));
Q_AD01HF U1161 ( .A0(ecmTsP[15]), .B0(n1160), .S(n1159), .CO(n1158));
Q_AD01HF U1162 ( .A0(ecmTsP[16]), .B0(n1158), .S(n1157), .CO(n1156));
Q_AD01HF U1163 ( .A0(ecmTsP[17]), .B0(n1156), .S(n1155), .CO(n1154));
Q_AD01HF U1164 ( .A0(ecmTsP[18]), .B0(n1154), .S(n1153), .CO(n1152));
Q_AD01HF U1165 ( .A0(ecmTsP[19]), .B0(n1152), .S(n1151), .CO(n1150));
Q_AD01HF U1166 ( .A0(ecmTsP[20]), .B0(n1150), .S(n1149), .CO(n1148));
Q_AD01HF U1167 ( .A0(ecmTsP[21]), .B0(n1148), .S(n1147), .CO(n1146));
Q_AD01HF U1168 ( .A0(ecmTsP[22]), .B0(n1146), .S(n1145), .CO(n1144));
Q_AD01HF U1169 ( .A0(ecmTsP[23]), .B0(n1144), .S(n1143), .CO(n1142));
Q_AD01HF U1170 ( .A0(ecmTsP[24]), .B0(n1142), .S(n1141), .CO(n1140));
Q_AD01HF U1171 ( .A0(ecmTsP[25]), .B0(n1140), .S(n1139), .CO(n1138));
Q_AD01HF U1172 ( .A0(ecmTsP[26]), .B0(n1138), .S(n1137), .CO(n1136));
Q_AD01HF U1173 ( .A0(ecmTsP[27]), .B0(n1136), .S(n1135), .CO(n1134));
Q_AD01HF U1174 ( .A0(ecmTsP[28]), .B0(n1134), .S(n1133), .CO(n1132));
Q_AD01HF U1175 ( .A0(ecmTsP[29]), .B0(n1132), .S(n1131), .CO(n1130));
Q_AD01HF U1176 ( .A0(ecmTsP[30]), .B0(n1130), .S(n1129), .CO(n1128));
Q_AD01HF U1177 ( .A0(ecmTsP[31]), .B0(n1128), .S(n1127), .CO(n1126));
Q_AD01HF U1178 ( .A0(ecmTsP[32]), .B0(n1126), .S(n1125), .CO(n1124));
Q_AD01HF U1179 ( .A0(ecmTsP[33]), .B0(n1124), .S(n1123), .CO(n1122));
Q_AD01HF U1180 ( .A0(ecmTsP[34]), .B0(n1122), .S(n1121), .CO(n1120));
Q_AD01HF U1181 ( .A0(ecmTsP[35]), .B0(n1120), .S(n1119), .CO(n1118));
Q_AD01HF U1182 ( .A0(ecmTsP[36]), .B0(n1118), .S(n1117), .CO(n1116));
Q_AD01HF U1183 ( .A0(ecmTsP[37]), .B0(n1116), .S(n1115), .CO(n1114));
Q_AD01HF U1184 ( .A0(ecmTsP[38]), .B0(n1114), .S(n1113), .CO(n1112));
Q_AD01HF U1185 ( .A0(ecmTsP[39]), .B0(n1112), .S(n1111), .CO(n1110));
Q_AD01HF U1186 ( .A0(ecmTsP[40]), .B0(n1110), .S(n1109), .CO(n1108));
Q_AD01HF U1187 ( .A0(ecmTsP[41]), .B0(n1108), .S(n1107), .CO(n1106));
Q_AD01HF U1188 ( .A0(ecmTsP[42]), .B0(n1106), .S(n1105), .CO(n1104));
Q_AD01HF U1189 ( .A0(ecmTsP[43]), .B0(n1104), .S(n1103), .CO(n1102));
Q_AD01HF U1190 ( .A0(ecmTsP[44]), .B0(n1102), .S(n1101), .CO(n1100));
Q_AD01HF U1191 ( .A0(ecmTsP[45]), .B0(n1100), .S(n1099), .CO(n1098));
Q_AD01HF U1192 ( .A0(ecmTsP[46]), .B0(n1098), .S(n1097), .CO(n1096));
Q_AD01HF U1193 ( .A0(ecmTsP[47]), .B0(n1096), .S(n1095), .CO(n1094));
Q_AD01HF U1194 ( .A0(ecmTsP[48]), .B0(n1094), .S(n1093), .CO(n1092));
Q_AD01HF U1195 ( .A0(ecmTsP[49]), .B0(n1092), .S(n1091), .CO(n1090));
Q_AD01HF U1196 ( .A0(ecmTsP[50]), .B0(n1090), .S(n1089), .CO(n1088));
Q_AD01HF U1197 ( .A0(ecmTsP[51]), .B0(n1088), .S(n1087), .CO(n1086));
Q_AD01HF U1198 ( .A0(ecmTsP[52]), .B0(n1086), .S(n1085), .CO(n1084));
Q_AD01HF U1199 ( .A0(ecmTsP[53]), .B0(n1084), .S(n1083), .CO(n1082));
Q_AD01HF U1200 ( .A0(ecmTsP[54]), .B0(n1082), .S(n1081), .CO(n1080));
Q_AD01HF U1201 ( .A0(ecmTsP[55]), .B0(n1080), .S(n1079), .CO(n1078));
Q_AD01HF U1202 ( .A0(ecmTsP[56]), .B0(n1078), .S(n1077), .CO(n1076));
Q_AD01HF U1203 ( .A0(ecmTsP[57]), .B0(n1076), .S(n1075), .CO(n1074));
Q_AD01HF U1204 ( .A0(ecmTsP[58]), .B0(n1074), .S(n1073), .CO(n1072));
Q_AD01HF U1205 ( .A0(ecmTsP[59]), .B0(n1072), .S(n1071), .CO(n1070));
Q_AD01HF U1206 ( .A0(ecmTsP[60]), .B0(n1070), .S(n1069), .CO(n1068));
Q_AD01HF U1207 ( .A0(ecmTsP[61]), .B0(n1068), .S(n1067), .CO(n1066));
Q_AD01HF U1208 ( .A0(ecmTsP[62]), .B0(n1066), .S(n1065), .CO(n1064));
Q_XOR2 U1209 ( .A0(ecmTsP[63]), .A1(n1742), .Z(ecmTs[63]));
Q_XOR2 U1210 ( .A0(xcva_top.xc_top.ecmOnD), .A1(ecmTsP[0]), .Z(ecmTs[0]));
Q_MX02 U1211 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[1]), .A1(n1187), .Z(ecmTs[1]));
Q_MX02 U1212 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[2]), .A1(n1185), .Z(ecmTs[2]));
Q_MX02 U1213 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[3]), .A1(n1183), .Z(ecmTs[3]));
Q_MX02 U1214 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[4]), .A1(n1181), .Z(ecmTs[4]));
Q_MX02 U1215 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[5]), .A1(n1179), .Z(ecmTs[5]));
Q_MX02 U1216 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[6]), .A1(n1177), .Z(ecmTs[6]));
Q_MX02 U1217 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[7]), .A1(n1175), .Z(ecmTs[7]));
Q_MX02 U1218 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[8]), .A1(n1173), .Z(ecmTs[8]));
Q_MX02 U1219 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[9]), .A1(n1171), .Z(ecmTs[9]));
Q_MX02 U1220 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[10]), .A1(n1169), .Z(ecmTs[10]));
Q_MX02 U1221 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[11]), .A1(n1167), .Z(ecmTs[11]));
Q_MX02 U1222 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[12]), .A1(n1165), .Z(ecmTs[12]));
Q_MX02 U1223 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[13]), .A1(n1163), .Z(ecmTs[13]));
Q_MX02 U1224 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[14]), .A1(n1161), .Z(ecmTs[14]));
Q_MX02 U1225 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[15]), .A1(n1159), .Z(ecmTs[15]));
Q_MX02 U1226 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[16]), .A1(n1157), .Z(ecmTs[16]));
Q_MX02 U1227 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[17]), .A1(n1155), .Z(ecmTs[17]));
Q_MX02 U1228 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[18]), .A1(n1153), .Z(ecmTs[18]));
Q_MX02 U1229 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[19]), .A1(n1151), .Z(ecmTs[19]));
Q_MX02 U1230 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[20]), .A1(n1149), .Z(ecmTs[20]));
Q_MX02 U1231 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[21]), .A1(n1147), .Z(ecmTs[21]));
Q_MX02 U1232 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[22]), .A1(n1145), .Z(ecmTs[22]));
Q_MX02 U1233 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[23]), .A1(n1143), .Z(ecmTs[23]));
Q_MX02 U1234 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[24]), .A1(n1141), .Z(ecmTs[24]));
Q_MX02 U1235 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[25]), .A1(n1139), .Z(ecmTs[25]));
Q_MX02 U1236 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[26]), .A1(n1137), .Z(ecmTs[26]));
Q_MX02 U1237 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[27]), .A1(n1135), .Z(ecmTs[27]));
Q_MX02 U1238 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[28]), .A1(n1133), .Z(ecmTs[28]));
Q_MX02 U1239 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[29]), .A1(n1131), .Z(ecmTs[29]));
Q_MX02 U1240 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[30]), .A1(n1129), .Z(ecmTs[30]));
Q_MX02 U1241 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[31]), .A1(n1127), .Z(ecmTs[31]));
Q_MX02 U1242 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[32]), .A1(n1125), .Z(ecmTs[32]));
Q_MX02 U1243 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[33]), .A1(n1123), .Z(ecmTs[33]));
Q_MX02 U1244 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[34]), .A1(n1121), .Z(ecmTs[34]));
Q_MX02 U1245 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[35]), .A1(n1119), .Z(ecmTs[35]));
Q_MX02 U1246 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[36]), .A1(n1117), .Z(ecmTs[36]));
Q_MX02 U1247 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[37]), .A1(n1115), .Z(ecmTs[37]));
Q_MX02 U1248 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[38]), .A1(n1113), .Z(ecmTs[38]));
Q_MX02 U1249 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[39]), .A1(n1111), .Z(ecmTs[39]));
Q_MX02 U1250 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[40]), .A1(n1109), .Z(ecmTs[40]));
Q_MX02 U1251 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[41]), .A1(n1107), .Z(ecmTs[41]));
Q_MX02 U1252 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[42]), .A1(n1105), .Z(ecmTs[42]));
Q_MX02 U1253 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[43]), .A1(n1103), .Z(ecmTs[43]));
Q_MX02 U1254 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[44]), .A1(n1101), .Z(ecmTs[44]));
Q_MX02 U1255 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[45]), .A1(n1099), .Z(ecmTs[45]));
Q_MX02 U1256 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[46]), .A1(n1097), .Z(ecmTs[46]));
Q_MX02 U1257 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[47]), .A1(n1095), .Z(ecmTs[47]));
Q_MX02 U1258 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[48]), .A1(n1093), .Z(ecmTs[48]));
Q_MX02 U1259 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[49]), .A1(n1091), .Z(ecmTs[49]));
Q_MX02 U1260 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[50]), .A1(n1089), .Z(ecmTs[50]));
Q_MX02 U1261 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[51]), .A1(n1087), .Z(ecmTs[51]));
Q_MX02 U1262 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[52]), .A1(n1085), .Z(ecmTs[52]));
Q_MX02 U1263 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[53]), .A1(n1083), .Z(ecmTs[53]));
Q_MX02 U1264 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[54]), .A1(n1081), .Z(ecmTs[54]));
Q_MX02 U1265 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[55]), .A1(n1079), .Z(ecmTs[55]));
Q_MX02 U1266 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[56]), .A1(n1077), .Z(ecmTs[56]));
Q_MX02 U1267 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[57]), .A1(n1075), .Z(ecmTs[57]));
Q_MX02 U1268 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[58]), .A1(n1073), .Z(ecmTs[58]));
Q_MX02 U1269 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[59]), .A1(n1071), .Z(ecmTs[59]));
Q_MX02 U1270 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[60]), .A1(n1069), .Z(ecmTs[60]));
Q_MX02 U1271 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[61]), .A1(n1067), .Z(ecmTs[61]));
Q_MX02 U1272 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[62]), .A1(n1065), .Z(ecmTs[62]));
Q_INV U1273 ( .A(ctrlW[127]), .Z(n1063));
Q_AO21 U1274 ( .A0(argTc[63]), .A1(n1063), .B0(n1054), .Z(n1053));
Q_OR02 U1275 ( .A0(argTc[63]), .A1(n1063), .Z(n1062));
Q_INV U1276 ( .A(ctrlW[126]), .Z(n1061));
Q_AN03 U1277 ( .A0(argTc[62]), .A1(n1061), .A2(n1062), .Z(n1054));
Q_OA21 U1278 ( .A0(argTc[62]), .A1(n1061), .B0(n1062), .Z(n1058));
Q_INV U1279 ( .A(ctrlW[125]), .Z(n1060));
Q_AN03 U1280 ( .A0(argTc[61]), .A1(n1060), .A2(n1058), .Z(n1055));
Q_OA21 U1281 ( .A0(argTc[61]), .A1(n1060), .B0(n1058), .Z(n1057));
Q_INV U1282 ( .A(ctrlW[124]), .Z(n1059));
Q_AN03 U1283 ( .A0(argTc[60]), .A1(n1059), .A2(n1057), .Z(n1056));
Q_OA21 U1284 ( .A0(argTc[60]), .A1(n1059), .B0(n1057), .Z(n1051));
Q_OR03 U1285 ( .A0(n1055), .A1(n1056), .A2(n1053), .Z(n1052));
Q_INV U1286 ( .A(ctrlW[123]), .Z(n1050));
Q_AO21 U1287 ( .A0(argTc[59]), .A1(n1050), .B0(n1041), .Z(n1040));
Q_OR02 U1288 ( .A0(argTc[59]), .A1(n1050), .Z(n1049));
Q_INV U1289 ( .A(ctrlW[122]), .Z(n1048));
Q_AN03 U1290 ( .A0(argTc[58]), .A1(n1048), .A2(n1049), .Z(n1041));
Q_OA21 U1291 ( .A0(argTc[58]), .A1(n1048), .B0(n1049), .Z(n1045));
Q_INV U1292 ( .A(ctrlW[121]), .Z(n1047));
Q_AN03 U1293 ( .A0(argTc[57]), .A1(n1047), .A2(n1045), .Z(n1042));
Q_OA21 U1294 ( .A0(argTc[57]), .A1(n1047), .B0(n1045), .Z(n1044));
Q_INV U1295 ( .A(ctrlW[120]), .Z(n1046));
Q_AN03 U1296 ( .A0(argTc[56]), .A1(n1046), .A2(n1044), .Z(n1043));
Q_OA21 U1297 ( .A0(argTc[56]), .A1(n1046), .B0(n1044), .Z(n1038));
Q_OR03 U1298 ( .A0(n1042), .A1(n1043), .A2(n1040), .Z(n1039));
Q_INV U1299 ( .A(ctrlW[119]), .Z(n1037));
Q_AO21 U1300 ( .A0(argTc[55]), .A1(n1037), .B0(n1028), .Z(n1027));
Q_OR02 U1301 ( .A0(argTc[55]), .A1(n1037), .Z(n1036));
Q_INV U1302 ( .A(ctrlW[118]), .Z(n1035));
Q_AN03 U1303 ( .A0(argTc[54]), .A1(n1035), .A2(n1036), .Z(n1028));
Q_OA21 U1304 ( .A0(argTc[54]), .A1(n1035), .B0(n1036), .Z(n1032));
Q_INV U1305 ( .A(ctrlW[117]), .Z(n1034));
Q_AN03 U1306 ( .A0(argTc[53]), .A1(n1034), .A2(n1032), .Z(n1029));
Q_OA21 U1307 ( .A0(argTc[53]), .A1(n1034), .B0(n1032), .Z(n1031));
Q_INV U1308 ( .A(ctrlW[116]), .Z(n1033));
Q_AN03 U1309 ( .A0(argTc[52]), .A1(n1033), .A2(n1031), .Z(n1030));
Q_OA21 U1310 ( .A0(argTc[52]), .A1(n1033), .B0(n1031), .Z(n1025));
Q_OR03 U1311 ( .A0(n1029), .A1(n1030), .A2(n1027), .Z(n1026));
Q_INV U1312 ( .A(ctrlW[115]), .Z(n1024));
Q_AO21 U1313 ( .A0(argTc[51]), .A1(n1024), .B0(n1015), .Z(n1014));
Q_OR02 U1314 ( .A0(argTc[51]), .A1(n1024), .Z(n1023));
Q_INV U1315 ( .A(ctrlW[114]), .Z(n1022));
Q_AN03 U1316 ( .A0(argTc[50]), .A1(n1022), .A2(n1023), .Z(n1015));
Q_OA21 U1317 ( .A0(argTc[50]), .A1(n1022), .B0(n1023), .Z(n1019));
Q_INV U1318 ( .A(ctrlW[113]), .Z(n1021));
Q_AN03 U1319 ( .A0(argTc[49]), .A1(n1021), .A2(n1019), .Z(n1016));
Q_OA21 U1320 ( .A0(argTc[49]), .A1(n1021), .B0(n1019), .Z(n1018));
Q_INV U1321 ( .A(ctrlW[112]), .Z(n1020));
Q_AN03 U1322 ( .A0(argTc[48]), .A1(n1020), .A2(n1018), .Z(n1017));
Q_OA21 U1323 ( .A0(argTc[48]), .A1(n1020), .B0(n1018), .Z(n1012));
Q_OR03 U1324 ( .A0(n1016), .A1(n1017), .A2(n1014), .Z(n1013));
Q_INV U1325 ( .A(ctrlW[111]), .Z(n1011));
Q_AO21 U1326 ( .A0(argTc[47]), .A1(n1011), .B0(n1002), .Z(n1001));
Q_OR02 U1327 ( .A0(argTc[47]), .A1(n1011), .Z(n1010));
Q_INV U1328 ( .A(ctrlW[110]), .Z(n1009));
Q_AN03 U1329 ( .A0(argTc[46]), .A1(n1009), .A2(n1010), .Z(n1002));
Q_OA21 U1330 ( .A0(argTc[46]), .A1(n1009), .B0(n1010), .Z(n1006));
Q_INV U1331 ( .A(ctrlW[109]), .Z(n1008));
Q_AN03 U1332 ( .A0(argTc[45]), .A1(n1008), .A2(n1006), .Z(n1003));
Q_OA21 U1333 ( .A0(argTc[45]), .A1(n1008), .B0(n1006), .Z(n1005));
Q_INV U1334 ( .A(ctrlW[108]), .Z(n1007));
Q_AN03 U1335 ( .A0(argTc[44]), .A1(n1007), .A2(n1005), .Z(n1004));
Q_OA21 U1336 ( .A0(argTc[44]), .A1(n1007), .B0(n1005), .Z(n999));
Q_OR03 U1337 ( .A0(n1003), .A1(n1004), .A2(n1001), .Z(n1000));
Q_INV U1338 ( .A(ctrlW[107]), .Z(n998));
Q_AO21 U1339 ( .A0(argTc[43]), .A1(n998), .B0(n989), .Z(n988));
Q_OR02 U1340 ( .A0(argTc[43]), .A1(n998), .Z(n997));
Q_INV U1341 ( .A(ctrlW[106]), .Z(n996));
Q_AN03 U1342 ( .A0(argTc[42]), .A1(n996), .A2(n997), .Z(n989));
Q_OA21 U1343 ( .A0(argTc[42]), .A1(n996), .B0(n997), .Z(n993));
Q_INV U1344 ( .A(ctrlW[105]), .Z(n995));
Q_AN03 U1345 ( .A0(argTc[41]), .A1(n995), .A2(n993), .Z(n990));
Q_OA21 U1346 ( .A0(argTc[41]), .A1(n995), .B0(n993), .Z(n992));
Q_INV U1347 ( .A(ctrlW[104]), .Z(n994));
Q_AN03 U1348 ( .A0(argTc[40]), .A1(n994), .A2(n992), .Z(n991));
Q_OA21 U1349 ( .A0(argTc[40]), .A1(n994), .B0(n992), .Z(n986));
Q_OR03 U1350 ( .A0(n990), .A1(n991), .A2(n988), .Z(n987));
Q_INV U1351 ( .A(ctrlW[103]), .Z(n985));
Q_AO21 U1352 ( .A0(argTc[39]), .A1(n985), .B0(n976), .Z(n975));
Q_OR02 U1353 ( .A0(argTc[39]), .A1(n985), .Z(n984));
Q_INV U1354 ( .A(ctrlW[102]), .Z(n983));
Q_AN03 U1355 ( .A0(argTc[38]), .A1(n983), .A2(n984), .Z(n976));
Q_OA21 U1356 ( .A0(argTc[38]), .A1(n983), .B0(n984), .Z(n980));
Q_INV U1357 ( .A(ctrlW[101]), .Z(n982));
Q_AN03 U1358 ( .A0(argTc[37]), .A1(n982), .A2(n980), .Z(n977));
Q_OA21 U1359 ( .A0(argTc[37]), .A1(n982), .B0(n980), .Z(n979));
Q_INV U1360 ( .A(ctrlW[100]), .Z(n981));
Q_AN03 U1361 ( .A0(argTc[36]), .A1(n981), .A2(n979), .Z(n978));
Q_OA21 U1362 ( .A0(argTc[36]), .A1(n981), .B0(n979), .Z(n973));
Q_OR03 U1363 ( .A0(n977), .A1(n978), .A2(n975), .Z(n974));
Q_INV U1364 ( .A(ctrlW[99]), .Z(n972));
Q_AO21 U1365 ( .A0(argTc[35]), .A1(n972), .B0(n963), .Z(n962));
Q_OR02 U1366 ( .A0(argTc[35]), .A1(n972), .Z(n971));
Q_INV U1367 ( .A(ctrlW[98]), .Z(n970));
Q_AN03 U1368 ( .A0(argTc[34]), .A1(n970), .A2(n971), .Z(n963));
Q_OA21 U1369 ( .A0(argTc[34]), .A1(n970), .B0(n971), .Z(n967));
Q_INV U1370 ( .A(ctrlW[97]), .Z(n969));
Q_AN03 U1371 ( .A0(argTc[33]), .A1(n969), .A2(n967), .Z(n964));
Q_OA21 U1372 ( .A0(argTc[33]), .A1(n969), .B0(n967), .Z(n966));
Q_INV U1373 ( .A(ctrlW[96]), .Z(n968));
Q_AN03 U1374 ( .A0(argTc[32]), .A1(n968), .A2(n966), .Z(n965));
Q_OA21 U1375 ( .A0(argTc[32]), .A1(n968), .B0(n966), .Z(n960));
Q_OR03 U1376 ( .A0(n964), .A1(n965), .A2(n962), .Z(n961));
Q_INV U1377 ( .A(ctrlW[95]), .Z(n959));
Q_AO21 U1378 ( .A0(argTc[31]), .A1(n959), .B0(n950), .Z(n949));
Q_OR02 U1379 ( .A0(argTc[31]), .A1(n959), .Z(n958));
Q_INV U1380 ( .A(ctrlW[94]), .Z(n957));
Q_AN03 U1381 ( .A0(argTc[30]), .A1(n957), .A2(n958), .Z(n950));
Q_OA21 U1382 ( .A0(argTc[30]), .A1(n957), .B0(n958), .Z(n954));
Q_INV U1383 ( .A(ctrlW[93]), .Z(n956));
Q_AN03 U1384 ( .A0(argTc[29]), .A1(n956), .A2(n954), .Z(n951));
Q_OA21 U1385 ( .A0(argTc[29]), .A1(n956), .B0(n954), .Z(n953));
Q_INV U1386 ( .A(ctrlW[92]), .Z(n955));
Q_AN03 U1387 ( .A0(argTc[28]), .A1(n955), .A2(n953), .Z(n952));
Q_OA21 U1388 ( .A0(argTc[28]), .A1(n955), .B0(n953), .Z(n947));
Q_OR03 U1389 ( .A0(n951), .A1(n952), .A2(n949), .Z(n948));
Q_INV U1390 ( .A(ctrlW[91]), .Z(n946));
Q_AO21 U1391 ( .A0(argTc[27]), .A1(n946), .B0(n937), .Z(n936));
Q_OR02 U1392 ( .A0(argTc[27]), .A1(n946), .Z(n945));
Q_INV U1393 ( .A(ctrlW[90]), .Z(n944));
Q_AN03 U1394 ( .A0(argTc[26]), .A1(n944), .A2(n945), .Z(n937));
Q_OA21 U1395 ( .A0(argTc[26]), .A1(n944), .B0(n945), .Z(n941));
Q_INV U1396 ( .A(ctrlW[89]), .Z(n943));
Q_AN03 U1397 ( .A0(argTc[25]), .A1(n943), .A2(n941), .Z(n938));
Q_OA21 U1398 ( .A0(argTc[25]), .A1(n943), .B0(n941), .Z(n940));
Q_INV U1399 ( .A(ctrlW[88]), .Z(n942));
Q_AN03 U1400 ( .A0(argTc[24]), .A1(n942), .A2(n940), .Z(n939));
Q_OA21 U1401 ( .A0(argTc[24]), .A1(n942), .B0(n940), .Z(n934));
Q_OR03 U1402 ( .A0(n938), .A1(n939), .A2(n936), .Z(n935));
Q_INV U1403 ( .A(ctrlW[87]), .Z(n933));
Q_AO21 U1404 ( .A0(argTc[23]), .A1(n933), .B0(n924), .Z(n923));
Q_OR02 U1405 ( .A0(argTc[23]), .A1(n933), .Z(n932));
Q_INV U1406 ( .A(ctrlW[86]), .Z(n931));
Q_AN03 U1407 ( .A0(argTc[22]), .A1(n931), .A2(n932), .Z(n924));
Q_OA21 U1408 ( .A0(argTc[22]), .A1(n931), .B0(n932), .Z(n928));
Q_INV U1409 ( .A(ctrlW[85]), .Z(n930));
Q_AN03 U1410 ( .A0(argTc[21]), .A1(n930), .A2(n928), .Z(n925));
Q_OA21 U1411 ( .A0(argTc[21]), .A1(n930), .B0(n928), .Z(n927));
Q_INV U1412 ( .A(ctrlW[84]), .Z(n929));
Q_AN03 U1413 ( .A0(argTc[20]), .A1(n929), .A2(n927), .Z(n926));
Q_OA21 U1414 ( .A0(argTc[20]), .A1(n929), .B0(n927), .Z(n921));
Q_OR03 U1415 ( .A0(n925), .A1(n926), .A2(n923), .Z(n922));
Q_INV U1416 ( .A(ctrlW[83]), .Z(n920));
Q_AO21 U1417 ( .A0(argTc[19]), .A1(n920), .B0(n911), .Z(n910));
Q_OR02 U1418 ( .A0(argTc[19]), .A1(n920), .Z(n919));
Q_INV U1419 ( .A(ctrlW[82]), .Z(n918));
Q_AN03 U1420 ( .A0(argTc[18]), .A1(n918), .A2(n919), .Z(n911));
Q_OA21 U1421 ( .A0(argTc[18]), .A1(n918), .B0(n919), .Z(n915));
Q_INV U1422 ( .A(ctrlW[81]), .Z(n917));
Q_AN03 U1423 ( .A0(argTc[17]), .A1(n917), .A2(n915), .Z(n912));
Q_OA21 U1424 ( .A0(argTc[17]), .A1(n917), .B0(n915), .Z(n914));
Q_INV U1425 ( .A(ctrlW[80]), .Z(n916));
Q_AN03 U1426 ( .A0(argTc[16]), .A1(n916), .A2(n914), .Z(n913));
Q_OA21 U1427 ( .A0(argTc[16]), .A1(n916), .B0(n914), .Z(n908));
Q_OR03 U1428 ( .A0(n912), .A1(n913), .A2(n910), .Z(n909));
Q_INV U1429 ( .A(ctrlW[79]), .Z(n907));
Q_AO21 U1430 ( .A0(argTc[15]), .A1(n907), .B0(n898), .Z(n897));
Q_OR02 U1431 ( .A0(argTc[15]), .A1(n907), .Z(n906));
Q_INV U1432 ( .A(ctrlW[78]), .Z(n905));
Q_AN03 U1433 ( .A0(argTc[14]), .A1(n905), .A2(n906), .Z(n898));
Q_OA21 U1434 ( .A0(argTc[14]), .A1(n905), .B0(n906), .Z(n902));
Q_INV U1435 ( .A(ctrlW[77]), .Z(n904));
Q_AN03 U1436 ( .A0(argTc[13]), .A1(n904), .A2(n902), .Z(n899));
Q_OA21 U1437 ( .A0(argTc[13]), .A1(n904), .B0(n902), .Z(n901));
Q_INV U1438 ( .A(ctrlW[76]), .Z(n903));
Q_AN03 U1439 ( .A0(argTc[12]), .A1(n903), .A2(n901), .Z(n900));
Q_OA21 U1440 ( .A0(argTc[12]), .A1(n903), .B0(n901), .Z(n895));
Q_OR03 U1441 ( .A0(n899), .A1(n900), .A2(n897), .Z(n896));
Q_INV U1442 ( .A(ctrlW[75]), .Z(n894));
Q_AO21 U1443 ( .A0(argTc[11]), .A1(n894), .B0(n885), .Z(n884));
Q_OR02 U1444 ( .A0(argTc[11]), .A1(n894), .Z(n893));
Q_INV U1445 ( .A(ctrlW[74]), .Z(n892));
Q_AN03 U1446 ( .A0(argTc[10]), .A1(n892), .A2(n893), .Z(n885));
Q_OA21 U1447 ( .A0(argTc[10]), .A1(n892), .B0(n893), .Z(n889));
Q_INV U1448 ( .A(ctrlW[73]), .Z(n891));
Q_AN03 U1449 ( .A0(argTc[9]), .A1(n891), .A2(n889), .Z(n886));
Q_OA21 U1450 ( .A0(argTc[9]), .A1(n891), .B0(n889), .Z(n888));
Q_INV U1451 ( .A(ctrlW[72]), .Z(n890));
Q_AN03 U1452 ( .A0(argTc[8]), .A1(n890), .A2(n888), .Z(n887));
Q_OA21 U1453 ( .A0(argTc[8]), .A1(n890), .B0(n888), .Z(n882));
Q_OR03 U1454 ( .A0(n886), .A1(n887), .A2(n884), .Z(n883));
Q_INV U1455 ( .A(ctrlW[71]), .Z(n881));
Q_AO21 U1456 ( .A0(argTc[7]), .A1(n881), .B0(n872), .Z(n871));
Q_OR02 U1457 ( .A0(argTc[7]), .A1(n881), .Z(n880));
Q_INV U1458 ( .A(ctrlW[70]), .Z(n879));
Q_AN03 U1459 ( .A0(argTc[6]), .A1(n879), .A2(n880), .Z(n872));
Q_OA21 U1460 ( .A0(argTc[6]), .A1(n879), .B0(n880), .Z(n876));
Q_INV U1461 ( .A(ctrlW[69]), .Z(n878));
Q_AN03 U1462 ( .A0(argTc[5]), .A1(n878), .A2(n876), .Z(n873));
Q_OA21 U1463 ( .A0(argTc[5]), .A1(n878), .B0(n876), .Z(n875));
Q_INV U1464 ( .A(ctrlW[68]), .Z(n877));
Q_AN03 U1465 ( .A0(argTc[4]), .A1(n877), .A2(n875), .Z(n874));
Q_OA21 U1466 ( .A0(argTc[4]), .A1(n877), .B0(n875), .Z(n869));
Q_OR03 U1467 ( .A0(n873), .A1(n874), .A2(n871), .Z(n870));
Q_INV U1468 ( .A(ctrlW[67]), .Z(n868));
Q_AO21 U1469 ( .A0(argTc[3]), .A1(n868), .B0(n859), .Z(n858));
Q_OR02 U1470 ( .A0(argTc[3]), .A1(n868), .Z(n867));
Q_INV U1471 ( .A(ctrlW[66]), .Z(n866));
Q_AN03 U1472 ( .A0(argTc[2]), .A1(n866), .A2(n867), .Z(n859));
Q_OA21 U1473 ( .A0(argTc[2]), .A1(n866), .B0(n867), .Z(n863));
Q_INV U1474 ( .A(ctrlW[65]), .Z(n865));
Q_AN03 U1475 ( .A0(argTc[1]), .A1(n865), .A2(n863), .Z(n860));
Q_OA21 U1476 ( .A0(argTc[1]), .A1(n865), .B0(n863), .Z(n862));
Q_INV U1477 ( .A(ctrlW[64]), .Z(n864));
Q_AN03 U1478 ( .A0(argTc[0]), .A1(n864), .A2(n862), .Z(n861));
Q_OR03 U1479 ( .A0(n860), .A1(n861), .A2(n858), .Z(n857));
Q_AN02 U1480 ( .A0(n1051), .A1(n1038), .Z(n856));
Q_AN02 U1481 ( .A0(n856), .A1(n1025), .Z(n855));
Q_AO21 U1482 ( .A0(n855), .A1(n1013), .B0(n854), .Z(n853));
Q_AN02 U1483 ( .A0(n856), .A1(n1026), .Z(n854));
Q_AO21 U1484 ( .A0(n1051), .A1(n1039), .B0(n1052), .Z(n852));
Q_OR03 U1485 ( .A0(n852), .A1(n853), .A2(n832), .Z(n831));
Q_AN02 U1486 ( .A0(n855), .A1(n1012), .Z(n851));
Q_AN02 U1487 ( .A0(n999), .A1(n986), .Z(n850));
Q_AN02 U1488 ( .A0(n850), .A1(n973), .Z(n849));
Q_AO21 U1489 ( .A0(n849), .A1(n961), .B0(n848), .Z(n847));
Q_AN02 U1490 ( .A0(n850), .A1(n974), .Z(n848));
Q_AO21 U1491 ( .A0(n999), .A1(n987), .B0(n1000), .Z(n846));
Q_OA21 U1492 ( .A0(n846), .A1(n847), .B0(n851), .Z(n832));
Q_AN03 U1493 ( .A0(n849), .A1(n960), .A2(n851), .Z(n836));
Q_AN02 U1494 ( .A0(n947), .A1(n934), .Z(n845));
Q_AN02 U1495 ( .A0(n845), .A1(n921), .Z(n844));
Q_AO21 U1496 ( .A0(n844), .A1(n909), .B0(n843), .Z(n842));
Q_AN02 U1497 ( .A0(n845), .A1(n922), .Z(n843));
Q_AO21 U1498 ( .A0(n947), .A1(n935), .B0(n948), .Z(n841));
Q_OA21 U1499 ( .A0(n841), .A1(n842), .B0(n836), .Z(n833));
Q_AN03 U1500 ( .A0(n844), .A1(n908), .A2(n836), .Z(n835));
Q_AN02 U1501 ( .A0(n895), .A1(n882), .Z(n840));
Q_AN03 U1502 ( .A0(n840), .A1(n869), .A2(n857), .Z(n839));
Q_AO21 U1503 ( .A0(n840), .A1(n870), .B0(n839), .Z(n838));
Q_AO21 U1504 ( .A0(n895), .A1(n883), .B0(n896), .Z(n837));
Q_OA21 U1505 ( .A0(n837), .A1(n838), .B0(n835), .Z(n834));
Q_NR03 U1506 ( .A0(n833), .A1(n834), .A2(n831), .Z(n830));
Q_AN02 U1507 ( .A0(cmdR[1]), .A1(n830), .Z(hc));
Q_INV U1508 ( .A(xcva_top.xc_top.simTime[63]), .Z(n829));
Q_AO21 U1509 ( .A0(argTs[63]), .A1(n829), .B0(n820), .Z(n819));
Q_OR02 U1510 ( .A0(argTs[63]), .A1(n829), .Z(n828));
Q_INV U1511 ( .A(xcva_top.xc_top.simTime[62]), .Z(n827));
Q_AN03 U1512 ( .A0(argTs[62]), .A1(n827), .A2(n828), .Z(n820));
Q_OA21 U1513 ( .A0(argTs[62]), .A1(n827), .B0(n828), .Z(n824));
Q_INV U1514 ( .A(xcva_top.xc_top.simTime[61]), .Z(n826));
Q_AN03 U1515 ( .A0(argTs[61]), .A1(n826), .A2(n824), .Z(n821));
Q_OA21 U1516 ( .A0(argTs[61]), .A1(n826), .B0(n824), .Z(n823));
Q_INV U1517 ( .A(xcva_top.xc_top.simTime[60]), .Z(n825));
Q_AN03 U1518 ( .A0(argTs[60]), .A1(n825), .A2(n823), .Z(n822));
Q_OA21 U1519 ( .A0(argTs[60]), .A1(n825), .B0(n823), .Z(n817));
Q_OR03 U1520 ( .A0(n821), .A1(n822), .A2(n819), .Z(n818));
Q_INV U1521 ( .A(xcva_top.xc_top.simTime[59]), .Z(n816));
Q_AO21 U1522 ( .A0(argTs[59]), .A1(n816), .B0(n807), .Z(n806));
Q_OR02 U1523 ( .A0(argTs[59]), .A1(n816), .Z(n815));
Q_INV U1524 ( .A(xcva_top.xc_top.simTime[58]), .Z(n814));
Q_AN03 U1525 ( .A0(argTs[58]), .A1(n814), .A2(n815), .Z(n807));
Q_OA21 U1526 ( .A0(argTs[58]), .A1(n814), .B0(n815), .Z(n811));
Q_INV U1527 ( .A(xcva_top.xc_top.simTime[57]), .Z(n813));
Q_AN03 U1528 ( .A0(argTs[57]), .A1(n813), .A2(n811), .Z(n808));
Q_OA21 U1529 ( .A0(argTs[57]), .A1(n813), .B0(n811), .Z(n810));
Q_INV U1530 ( .A(xcva_top.xc_top.simTime[56]), .Z(n812));
Q_AN03 U1531 ( .A0(argTs[56]), .A1(n812), .A2(n810), .Z(n809));
Q_OA21 U1532 ( .A0(argTs[56]), .A1(n812), .B0(n810), .Z(n804));
Q_OR03 U1533 ( .A0(n808), .A1(n809), .A2(n806), .Z(n805));
Q_INV U1534 ( .A(xcva_top.xc_top.simTime[55]), .Z(n803));
Q_AO21 U1535 ( .A0(argTs[55]), .A1(n803), .B0(n794), .Z(n793));
Q_OR02 U1536 ( .A0(argTs[55]), .A1(n803), .Z(n802));
Q_INV U1537 ( .A(xcva_top.xc_top.simTime[54]), .Z(n801));
Q_AN03 U1538 ( .A0(argTs[54]), .A1(n801), .A2(n802), .Z(n794));
Q_OA21 U1539 ( .A0(argTs[54]), .A1(n801), .B0(n802), .Z(n798));
Q_INV U1540 ( .A(xcva_top.xc_top.simTime[53]), .Z(n800));
Q_AN03 U1541 ( .A0(argTs[53]), .A1(n800), .A2(n798), .Z(n795));
Q_OA21 U1542 ( .A0(argTs[53]), .A1(n800), .B0(n798), .Z(n797));
Q_INV U1543 ( .A(xcva_top.xc_top.simTime[52]), .Z(n799));
Q_AN03 U1544 ( .A0(argTs[52]), .A1(n799), .A2(n797), .Z(n796));
Q_OA21 U1545 ( .A0(argTs[52]), .A1(n799), .B0(n797), .Z(n791));
Q_OR03 U1546 ( .A0(n795), .A1(n796), .A2(n793), .Z(n792));
Q_INV U1547 ( .A(xcva_top.xc_top.simTime[51]), .Z(n790));
Q_AO21 U1548 ( .A0(argTs[51]), .A1(n790), .B0(n781), .Z(n780));
Q_OR02 U1549 ( .A0(argTs[51]), .A1(n790), .Z(n789));
Q_INV U1550 ( .A(xcva_top.xc_top.simTime[50]), .Z(n788));
Q_AN03 U1551 ( .A0(argTs[50]), .A1(n788), .A2(n789), .Z(n781));
Q_OA21 U1552 ( .A0(argTs[50]), .A1(n788), .B0(n789), .Z(n785));
Q_INV U1553 ( .A(xcva_top.xc_top.simTime[49]), .Z(n787));
Q_AN03 U1554 ( .A0(argTs[49]), .A1(n787), .A2(n785), .Z(n782));
Q_OA21 U1555 ( .A0(argTs[49]), .A1(n787), .B0(n785), .Z(n784));
Q_INV U1556 ( .A(xcva_top.xc_top.simTime[48]), .Z(n786));
Q_AN03 U1557 ( .A0(argTs[48]), .A1(n786), .A2(n784), .Z(n783));
Q_OA21 U1558 ( .A0(argTs[48]), .A1(n786), .B0(n784), .Z(n778));
Q_OR03 U1559 ( .A0(n782), .A1(n783), .A2(n780), .Z(n779));
Q_INV U1560 ( .A(xcva_top.xc_top.simTime[47]), .Z(n777));
Q_AO21 U1561 ( .A0(argTs[47]), .A1(n777), .B0(n768), .Z(n767));
Q_OR02 U1562 ( .A0(argTs[47]), .A1(n777), .Z(n776));
Q_INV U1563 ( .A(xcva_top.xc_top.simTime[46]), .Z(n775));
Q_AN03 U1564 ( .A0(argTs[46]), .A1(n775), .A2(n776), .Z(n768));
Q_OA21 U1565 ( .A0(argTs[46]), .A1(n775), .B0(n776), .Z(n772));
Q_INV U1566 ( .A(xcva_top.xc_top.simTime[45]), .Z(n774));
Q_AN03 U1567 ( .A0(argTs[45]), .A1(n774), .A2(n772), .Z(n769));
Q_OA21 U1568 ( .A0(argTs[45]), .A1(n774), .B0(n772), .Z(n771));
Q_INV U1569 ( .A(xcva_top.xc_top.simTime[44]), .Z(n773));
Q_AN03 U1570 ( .A0(argTs[44]), .A1(n773), .A2(n771), .Z(n770));
Q_OA21 U1571 ( .A0(argTs[44]), .A1(n773), .B0(n771), .Z(n765));
Q_OR03 U1572 ( .A0(n769), .A1(n770), .A2(n767), .Z(n766));
Q_INV U1573 ( .A(xcva_top.xc_top.simTime[43]), .Z(n764));
Q_AO21 U1574 ( .A0(argTs[43]), .A1(n764), .B0(n755), .Z(n754));
Q_OR02 U1575 ( .A0(argTs[43]), .A1(n764), .Z(n763));
Q_INV U1576 ( .A(xcva_top.xc_top.simTime[42]), .Z(n762));
Q_AN03 U1577 ( .A0(argTs[42]), .A1(n762), .A2(n763), .Z(n755));
Q_OA21 U1578 ( .A0(argTs[42]), .A1(n762), .B0(n763), .Z(n759));
Q_INV U1579 ( .A(xcva_top.xc_top.simTime[41]), .Z(n761));
Q_AN03 U1580 ( .A0(argTs[41]), .A1(n761), .A2(n759), .Z(n756));
Q_OA21 U1581 ( .A0(argTs[41]), .A1(n761), .B0(n759), .Z(n758));
Q_INV U1582 ( .A(xcva_top.xc_top.simTime[40]), .Z(n760));
Q_AN03 U1583 ( .A0(argTs[40]), .A1(n760), .A2(n758), .Z(n757));
Q_OA21 U1584 ( .A0(argTs[40]), .A1(n760), .B0(n758), .Z(n752));
Q_OR03 U1585 ( .A0(n756), .A1(n757), .A2(n754), .Z(n753));
Q_INV U1586 ( .A(xcva_top.xc_top.simTime[39]), .Z(n751));
Q_AO21 U1587 ( .A0(argTs[39]), .A1(n751), .B0(n742), .Z(n741));
Q_OR02 U1588 ( .A0(argTs[39]), .A1(n751), .Z(n750));
Q_INV U1589 ( .A(xcva_top.xc_top.simTime[38]), .Z(n749));
Q_AN03 U1590 ( .A0(argTs[38]), .A1(n749), .A2(n750), .Z(n742));
Q_OA21 U1591 ( .A0(argTs[38]), .A1(n749), .B0(n750), .Z(n746));
Q_INV U1592 ( .A(xcva_top.xc_top.simTime[37]), .Z(n748));
Q_AN03 U1593 ( .A0(argTs[37]), .A1(n748), .A2(n746), .Z(n743));
Q_OA21 U1594 ( .A0(argTs[37]), .A1(n748), .B0(n746), .Z(n745));
Q_INV U1595 ( .A(xcva_top.xc_top.simTime[36]), .Z(n747));
Q_AN03 U1596 ( .A0(argTs[36]), .A1(n747), .A2(n745), .Z(n744));
Q_OA21 U1597 ( .A0(argTs[36]), .A1(n747), .B0(n745), .Z(n739));
Q_OR03 U1598 ( .A0(n743), .A1(n744), .A2(n741), .Z(n740));
Q_INV U1599 ( .A(xcva_top.xc_top.simTime[35]), .Z(n738));
Q_AO21 U1600 ( .A0(argTs[35]), .A1(n738), .B0(n729), .Z(n728));
Q_OR02 U1601 ( .A0(argTs[35]), .A1(n738), .Z(n737));
Q_INV U1602 ( .A(xcva_top.xc_top.simTime[34]), .Z(n736));
Q_AN03 U1603 ( .A0(argTs[34]), .A1(n736), .A2(n737), .Z(n729));
Q_OA21 U1604 ( .A0(argTs[34]), .A1(n736), .B0(n737), .Z(n733));
Q_INV U1605 ( .A(xcva_top.xc_top.simTime[33]), .Z(n735));
Q_AN03 U1606 ( .A0(argTs[33]), .A1(n735), .A2(n733), .Z(n730));
Q_OA21 U1607 ( .A0(argTs[33]), .A1(n735), .B0(n733), .Z(n732));
Q_INV U1608 ( .A(xcva_top.xc_top.simTime[32]), .Z(n734));
Q_AN03 U1609 ( .A0(argTs[32]), .A1(n734), .A2(n732), .Z(n731));
Q_OA21 U1610 ( .A0(argTs[32]), .A1(n734), .B0(n732), .Z(n726));
Q_OR03 U1611 ( .A0(n730), .A1(n731), .A2(n728), .Z(n727));
Q_INV U1612 ( .A(xcva_top.xc_top.simTime[31]), .Z(n725));
Q_AO21 U1613 ( .A0(argTs[31]), .A1(n725), .B0(n716), .Z(n715));
Q_OR02 U1614 ( .A0(argTs[31]), .A1(n725), .Z(n724));
Q_INV U1615 ( .A(xcva_top.xc_top.simTime[30]), .Z(n723));
Q_AN03 U1616 ( .A0(argTs[30]), .A1(n723), .A2(n724), .Z(n716));
Q_OA21 U1617 ( .A0(argTs[30]), .A1(n723), .B0(n724), .Z(n720));
Q_INV U1618 ( .A(xcva_top.xc_top.simTime[29]), .Z(n722));
Q_AN03 U1619 ( .A0(argTs[29]), .A1(n722), .A2(n720), .Z(n717));
Q_OA21 U1620 ( .A0(argTs[29]), .A1(n722), .B0(n720), .Z(n719));
Q_INV U1621 ( .A(xcva_top.xc_top.simTime[28]), .Z(n721));
Q_AN03 U1622 ( .A0(argTs[28]), .A1(n721), .A2(n719), .Z(n718));
Q_OA21 U1623 ( .A0(argTs[28]), .A1(n721), .B0(n719), .Z(n713));
Q_OR03 U1624 ( .A0(n717), .A1(n718), .A2(n715), .Z(n714));
Q_INV U1625 ( .A(xcva_top.xc_top.simTime[27]), .Z(n712));
Q_AO21 U1626 ( .A0(argTs[27]), .A1(n712), .B0(n703), .Z(n702));
Q_OR02 U1627 ( .A0(argTs[27]), .A1(n712), .Z(n711));
Q_INV U1628 ( .A(xcva_top.xc_top.simTime[26]), .Z(n710));
Q_AN03 U1629 ( .A0(argTs[26]), .A1(n710), .A2(n711), .Z(n703));
Q_OA21 U1630 ( .A0(argTs[26]), .A1(n710), .B0(n711), .Z(n707));
Q_INV U1631 ( .A(xcva_top.xc_top.simTime[25]), .Z(n709));
Q_AN03 U1632 ( .A0(argTs[25]), .A1(n709), .A2(n707), .Z(n704));
Q_OA21 U1633 ( .A0(argTs[25]), .A1(n709), .B0(n707), .Z(n706));
Q_INV U1634 ( .A(xcva_top.xc_top.simTime[24]), .Z(n708));
Q_AN03 U1635 ( .A0(argTs[24]), .A1(n708), .A2(n706), .Z(n705));
Q_OA21 U1636 ( .A0(argTs[24]), .A1(n708), .B0(n706), .Z(n700));
Q_OR03 U1637 ( .A0(n704), .A1(n705), .A2(n702), .Z(n701));
Q_INV U1638 ( .A(xcva_top.xc_top.simTime[23]), .Z(n699));
Q_AO21 U1639 ( .A0(argTs[23]), .A1(n699), .B0(n690), .Z(n689));
Q_OR02 U1640 ( .A0(argTs[23]), .A1(n699), .Z(n698));
Q_INV U1641 ( .A(xcva_top.xc_top.simTime[22]), .Z(n697));
Q_AN03 U1642 ( .A0(argTs[22]), .A1(n697), .A2(n698), .Z(n690));
Q_OA21 U1643 ( .A0(argTs[22]), .A1(n697), .B0(n698), .Z(n694));
Q_INV U1644 ( .A(xcva_top.xc_top.simTime[21]), .Z(n696));
Q_AN03 U1645 ( .A0(argTs[21]), .A1(n696), .A2(n694), .Z(n691));
Q_OA21 U1646 ( .A0(argTs[21]), .A1(n696), .B0(n694), .Z(n693));
Q_INV U1647 ( .A(xcva_top.xc_top.simTime[20]), .Z(n695));
Q_AN03 U1648 ( .A0(argTs[20]), .A1(n695), .A2(n693), .Z(n692));
Q_OA21 U1649 ( .A0(argTs[20]), .A1(n695), .B0(n693), .Z(n687));
Q_OR03 U1650 ( .A0(n691), .A1(n692), .A2(n689), .Z(n688));
Q_INV U1651 ( .A(xcva_top.xc_top.simTime[19]), .Z(n686));
Q_AO21 U1652 ( .A0(argTs[19]), .A1(n686), .B0(n677), .Z(n676));
Q_OR02 U1653 ( .A0(argTs[19]), .A1(n686), .Z(n685));
Q_INV U1654 ( .A(xcva_top.xc_top.simTime[18]), .Z(n684));
Q_AN03 U1655 ( .A0(argTs[18]), .A1(n684), .A2(n685), .Z(n677));
Q_OA21 U1656 ( .A0(argTs[18]), .A1(n684), .B0(n685), .Z(n681));
Q_INV U1657 ( .A(xcva_top.xc_top.simTime[17]), .Z(n683));
Q_AN03 U1658 ( .A0(argTs[17]), .A1(n683), .A2(n681), .Z(n678));
Q_OA21 U1659 ( .A0(argTs[17]), .A1(n683), .B0(n681), .Z(n680));
Q_INV U1660 ( .A(xcva_top.xc_top.simTime[16]), .Z(n682));
Q_AN03 U1661 ( .A0(argTs[16]), .A1(n682), .A2(n680), .Z(n679));
Q_OA21 U1662 ( .A0(argTs[16]), .A1(n682), .B0(n680), .Z(n674));
Q_OR03 U1663 ( .A0(n678), .A1(n679), .A2(n676), .Z(n675));
Q_INV U1664 ( .A(xcva_top.xc_top.simTime[15]), .Z(n673));
Q_AO21 U1665 ( .A0(argTs[15]), .A1(n673), .B0(n664), .Z(n663));
Q_OR02 U1666 ( .A0(argTs[15]), .A1(n673), .Z(n672));
Q_INV U1667 ( .A(xcva_top.xc_top.simTime[14]), .Z(n671));
Q_AN03 U1668 ( .A0(argTs[14]), .A1(n671), .A2(n672), .Z(n664));
Q_OA21 U1669 ( .A0(argTs[14]), .A1(n671), .B0(n672), .Z(n668));
Q_INV U1670 ( .A(xcva_top.xc_top.simTime[13]), .Z(n670));
Q_AN03 U1671 ( .A0(argTs[13]), .A1(n670), .A2(n668), .Z(n665));
Q_OA21 U1672 ( .A0(argTs[13]), .A1(n670), .B0(n668), .Z(n667));
Q_INV U1673 ( .A(xcva_top.xc_top.simTime[12]), .Z(n669));
Q_AN03 U1674 ( .A0(argTs[12]), .A1(n669), .A2(n667), .Z(n666));
Q_OA21 U1675 ( .A0(argTs[12]), .A1(n669), .B0(n667), .Z(n661));
Q_OR03 U1676 ( .A0(n665), .A1(n666), .A2(n663), .Z(n662));
Q_INV U1677 ( .A(xcva_top.xc_top.simTime[11]), .Z(n660));
Q_AO21 U1678 ( .A0(argTs[11]), .A1(n660), .B0(n651), .Z(n650));
Q_OR02 U1679 ( .A0(argTs[11]), .A1(n660), .Z(n659));
Q_INV U1680 ( .A(xcva_top.xc_top.simTime[10]), .Z(n658));
Q_AN03 U1681 ( .A0(argTs[10]), .A1(n658), .A2(n659), .Z(n651));
Q_OA21 U1682 ( .A0(argTs[10]), .A1(n658), .B0(n659), .Z(n655));
Q_INV U1683 ( .A(xcva_top.xc_top.simTime[9]), .Z(n657));
Q_AN03 U1684 ( .A0(argTs[9]), .A1(n657), .A2(n655), .Z(n652));
Q_OA21 U1685 ( .A0(argTs[9]), .A1(n657), .B0(n655), .Z(n654));
Q_INV U1686 ( .A(xcva_top.xc_top.simTime[8]), .Z(n656));
Q_AN03 U1687 ( .A0(argTs[8]), .A1(n656), .A2(n654), .Z(n653));
Q_OA21 U1688 ( .A0(argTs[8]), .A1(n656), .B0(n654), .Z(n648));
Q_OR03 U1689 ( .A0(n652), .A1(n653), .A2(n650), .Z(n649));
Q_INV U1690 ( .A(xcva_top.xc_top.simTime[7]), .Z(n647));
Q_AO21 U1691 ( .A0(argTs[7]), .A1(n647), .B0(n638), .Z(n637));
Q_OR02 U1692 ( .A0(argTs[7]), .A1(n647), .Z(n646));
Q_INV U1693 ( .A(xcva_top.xc_top.simTime[6]), .Z(n645));
Q_AN03 U1694 ( .A0(argTs[6]), .A1(n645), .A2(n646), .Z(n638));
Q_OA21 U1695 ( .A0(argTs[6]), .A1(n645), .B0(n646), .Z(n642));
Q_INV U1696 ( .A(xcva_top.xc_top.simTime[5]), .Z(n644));
Q_AN03 U1697 ( .A0(argTs[5]), .A1(n644), .A2(n642), .Z(n639));
Q_OA21 U1698 ( .A0(argTs[5]), .A1(n644), .B0(n642), .Z(n641));
Q_INV U1699 ( .A(xcva_top.xc_top.simTime[4]), .Z(n643));
Q_AN03 U1700 ( .A0(argTs[4]), .A1(n643), .A2(n641), .Z(n640));
Q_OA21 U1701 ( .A0(argTs[4]), .A1(n643), .B0(n641), .Z(n635));
Q_OR03 U1702 ( .A0(n639), .A1(n640), .A2(n637), .Z(n636));
Q_INV U1703 ( .A(xcva_top.xc_top.simTime[3]), .Z(n634));
Q_AO21 U1704 ( .A0(argTs[3]), .A1(n634), .B0(n625), .Z(n624));
Q_OR02 U1705 ( .A0(argTs[3]), .A1(n634), .Z(n633));
Q_INV U1706 ( .A(xcva_top.xc_top.simTime[2]), .Z(n632));
Q_AN03 U1707 ( .A0(argTs[2]), .A1(n632), .A2(n633), .Z(n625));
Q_OA21 U1708 ( .A0(argTs[2]), .A1(n632), .B0(n633), .Z(n629));
Q_INV U1709 ( .A(xcva_top.xc_top.simTime[1]), .Z(n631));
Q_AN03 U1710 ( .A0(argTs[1]), .A1(n631), .A2(n629), .Z(n626));
Q_OA21 U1711 ( .A0(argTs[1]), .A1(n631), .B0(n629), .Z(n628));
Q_INV U1712 ( .A(xcva_top.xc_top.simTime[0]), .Z(n630));
Q_AN03 U1713 ( .A0(argTs[0]), .A1(n630), .A2(n628), .Z(n627));
Q_OR03 U1714 ( .A0(n626), .A1(n627), .A2(n624), .Z(n623));
Q_AN02 U1715 ( .A0(n817), .A1(n804), .Z(n622));
Q_AN02 U1716 ( .A0(n622), .A1(n791), .Z(n621));
Q_AO21 U1717 ( .A0(n621), .A1(n779), .B0(n620), .Z(n619));
Q_AN02 U1718 ( .A0(n622), .A1(n792), .Z(n620));
Q_AO21 U1719 ( .A0(n817), .A1(n805), .B0(n818), .Z(n618));
Q_OR03 U1720 ( .A0(n618), .A1(n619), .A2(n598), .Z(n597));
Q_AN02 U1721 ( .A0(n621), .A1(n778), .Z(n617));
Q_AN02 U1722 ( .A0(n765), .A1(n752), .Z(n616));
Q_AN02 U1723 ( .A0(n616), .A1(n739), .Z(n615));
Q_AO21 U1724 ( .A0(n615), .A1(n727), .B0(n614), .Z(n613));
Q_AN02 U1725 ( .A0(n616), .A1(n740), .Z(n614));
Q_AO21 U1726 ( .A0(n765), .A1(n753), .B0(n766), .Z(n612));
Q_OA21 U1727 ( .A0(n612), .A1(n613), .B0(n617), .Z(n598));
Q_AN03 U1728 ( .A0(n615), .A1(n726), .A2(n617), .Z(n602));
Q_AN02 U1729 ( .A0(n713), .A1(n700), .Z(n611));
Q_AN02 U1730 ( .A0(n611), .A1(n687), .Z(n610));
Q_AO21 U1731 ( .A0(n610), .A1(n675), .B0(n609), .Z(n608));
Q_AN02 U1732 ( .A0(n611), .A1(n688), .Z(n609));
Q_AO21 U1733 ( .A0(n713), .A1(n701), .B0(n714), .Z(n607));
Q_OA21 U1734 ( .A0(n607), .A1(n608), .B0(n602), .Z(n599));
Q_AN03 U1735 ( .A0(n610), .A1(n674), .A2(n602), .Z(n601));
Q_AN02 U1736 ( .A0(n661), .A1(n648), .Z(n606));
Q_AN03 U1737 ( .A0(n606), .A1(n635), .A2(n623), .Z(n605));
Q_AO21 U1738 ( .A0(n606), .A1(n636), .B0(n605), .Z(n604));
Q_AO21 U1739 ( .A0(n661), .A1(n649), .B0(n662), .Z(n603));
Q_OA21 U1740 ( .A0(n603), .A1(n604), .B0(n601), .Z(n600));
Q_NR03 U1741 ( .A0(n599), .A1(n600), .A2(n597), .Z(n596));
Q_AN02 U1742 ( .A0(cmdR[2]), .A1(n596), .Z(hs));
Q_OR03 U1743 ( .A0(sdlStopRply), .A1(cmdC[0]), .A2(hs), .Z(n595));
Q_OR02 U1744 ( .A0(n595), .A1(hc), .Z(holdEcm));
Q_FDP0 \ctrlR_REG[255] ( .CK(uclk), .D(n338), .Q(ctrlR[255]), .QN( ));
Q_FDP0 \ctrlR_REG[254] ( .CK(uclk), .D(n339), .Q(ctrlR[254]), .QN( ));
Q_FDP0 \ctrlR_REG[253] ( .CK(uclk), .D(n340), .Q(ctrlR[253]), .QN( ));
Q_FDP0 \ctrlR_REG[252] ( .CK(uclk), .D(n341), .Q(ctrlR[252]), .QN( ));
Q_FDP0 \ctrlR_REG[251] ( .CK(uclk), .D(n342), .Q(ctrlR[251]), .QN( ));
Q_FDP0 \ctrlR_REG[250] ( .CK(uclk), .D(n343), .Q(ctrlR[250]), .QN( ));
Q_FDP0 \ctrlR_REG[249] ( .CK(uclk), .D(n344), .Q(ctrlR[249]), .QN( ));
Q_FDP0 \ctrlR_REG[248] ( .CK(uclk), .D(n345), .Q(ctrlR[248]), .QN( ));
Q_FDP0 \ctrlR_REG[247] ( .CK(uclk), .D(n346), .Q(ctrlR[247]), .QN( ));
Q_FDP0 \ctrlR_REG[246] ( .CK(uclk), .D(n347), .Q(ctrlR[246]), .QN( ));
Q_FDP0 \ctrlR_REG[245] ( .CK(uclk), .D(n348), .Q(ctrlR[245]), .QN( ));
Q_FDP0 \ctrlR_REG[244] ( .CK(uclk), .D(n349), .Q(ctrlR[244]), .QN( ));
Q_FDP0 \ctrlR_REG[243] ( .CK(uclk), .D(n350), .Q(ctrlR[243]), .QN( ));
Q_FDP0 \ctrlR_REG[242] ( .CK(uclk), .D(n351), .Q(ctrlR[242]), .QN( ));
Q_FDP0 \ctrlR_REG[241] ( .CK(uclk), .D(n352), .Q(ctrlR[241]), .QN( ));
Q_FDP0 \ctrlR_REG[240] ( .CK(uclk), .D(n353), .Q(ctrlR[240]), .QN( ));
Q_FDP0 \ctrlR_REG[239] ( .CK(uclk), .D(n354), .Q(ctrlR[239]), .QN( ));
Q_FDP0 \ctrlR_REG[238] ( .CK(uclk), .D(n355), .Q(ctrlR[238]), .QN( ));
Q_FDP0 \ctrlR_REG[237] ( .CK(uclk), .D(n356), .Q(ctrlR[237]), .QN( ));
Q_FDP0 \ctrlR_REG[236] ( .CK(uclk), .D(n357), .Q(ctrlR[236]), .QN( ));
Q_FDP0 \ctrlR_REG[235] ( .CK(uclk), .D(n358), .Q(ctrlR[235]), .QN( ));
Q_FDP0 \ctrlR_REG[234] ( .CK(uclk), .D(n359), .Q(ctrlR[234]), .QN( ));
Q_FDP0 \ctrlR_REG[233] ( .CK(uclk), .D(n360), .Q(ctrlR[233]), .QN( ));
Q_FDP0 \ctrlR_REG[232] ( .CK(uclk), .D(n361), .Q(ctrlR[232]), .QN( ));
Q_FDP0 \ctrlR_REG[231] ( .CK(uclk), .D(n362), .Q(ctrlR[231]), .QN( ));
Q_FDP0 \ctrlR_REG[230] ( .CK(uclk), .D(n363), .Q(ctrlR[230]), .QN( ));
Q_FDP0 \ctrlR_REG[229] ( .CK(uclk), .D(n364), .Q(ctrlR[229]), .QN( ));
Q_FDP0 \ctrlR_REG[228] ( .CK(uclk), .D(n365), .Q(ctrlR[228]), .QN( ));
Q_FDP0 \ctrlR_REG[227] ( .CK(uclk), .D(n366), .Q(ctrlR[227]), .QN( ));
Q_FDP0 \ctrlR_REG[226] ( .CK(uclk), .D(n367), .Q(ctrlR[226]), .QN( ));
Q_FDP0 \ctrlR_REG[225] ( .CK(uclk), .D(n368), .Q(ctrlR[225]), .QN( ));
Q_FDP0 \ctrlR_REG[224] ( .CK(uclk), .D(n369), .Q(ctrlR[224]), .QN( ));
Q_FDP0 \ctrlR_REG[223] ( .CK(uclk), .D(n370), .Q(ctrlR[223]), .QN( ));
Q_FDP0 \ctrlR_REG[222] ( .CK(uclk), .D(n371), .Q(ctrlR[222]), .QN( ));
Q_FDP0 \ctrlR_REG[221] ( .CK(uclk), .D(n372), .Q(ctrlR[221]), .QN( ));
Q_FDP0 \ctrlR_REG[220] ( .CK(uclk), .D(n373), .Q(ctrlR[220]), .QN( ));
Q_FDP0 \ctrlR_REG[219] ( .CK(uclk), .D(n374), .Q(ctrlR[219]), .QN( ));
Q_FDP0 \ctrlR_REG[218] ( .CK(uclk), .D(n375), .Q(ctrlR[218]), .QN( ));
Q_FDP0 \ctrlR_REG[217] ( .CK(uclk), .D(n376), .Q(ctrlR[217]), .QN( ));
Q_FDP0 \ctrlR_REG[216] ( .CK(uclk), .D(n377), .Q(ctrlR[216]), .QN( ));
Q_FDP0 \ctrlR_REG[215] ( .CK(uclk), .D(n378), .Q(ctrlR[215]), .QN( ));
Q_FDP0 \ctrlR_REG[214] ( .CK(uclk), .D(n379), .Q(ctrlR[214]), .QN( ));
Q_FDP0 \ctrlR_REG[213] ( .CK(uclk), .D(n380), .Q(ctrlR[213]), .QN( ));
Q_FDP0 \ctrlR_REG[212] ( .CK(uclk), .D(n381), .Q(ctrlR[212]), .QN( ));
Q_FDP0 \ctrlR_REG[211] ( .CK(uclk), .D(n382), .Q(ctrlR[211]), .QN( ));
Q_FDP0 \ctrlR_REG[210] ( .CK(uclk), .D(n383), .Q(ctrlR[210]), .QN( ));
Q_FDP0 \ctrlR_REG[209] ( .CK(uclk), .D(n384), .Q(ctrlR[209]), .QN( ));
Q_FDP0 \ctrlR_REG[208] ( .CK(uclk), .D(n385), .Q(ctrlR[208]), .QN( ));
Q_FDP0 \ctrlR_REG[207] ( .CK(uclk), .D(n386), .Q(ctrlR[207]), .QN( ));
Q_FDP0 \ctrlR_REG[206] ( .CK(uclk), .D(n387), .Q(ctrlR[206]), .QN( ));
Q_FDP0 \ctrlR_REG[205] ( .CK(uclk), .D(n388), .Q(ctrlR[205]), .QN( ));
Q_FDP0 \ctrlR_REG[204] ( .CK(uclk), .D(n389), .Q(ctrlR[204]), .QN( ));
Q_FDP0 \ctrlR_REG[203] ( .CK(uclk), .D(n390), .Q(ctrlR[203]), .QN( ));
Q_FDP0 \ctrlR_REG[202] ( .CK(uclk), .D(n391), .Q(ctrlR[202]), .QN( ));
Q_FDP0 \ctrlR_REG[201] ( .CK(uclk), .D(n392), .Q(ctrlR[201]), .QN( ));
Q_FDP0 \ctrlR_REG[200] ( .CK(uclk), .D(n393), .Q(ctrlR[200]), .QN( ));
Q_FDP0 \ctrlR_REG[199] ( .CK(uclk), .D(n394), .Q(ctrlR[199]), .QN( ));
Q_FDP0 \ctrlR_REG[198] ( .CK(uclk), .D(n395), .Q(ctrlR[198]), .QN( ));
Q_FDP0 \ctrlR_REG[197] ( .CK(uclk), .D(n396), .Q(ctrlR[197]), .QN( ));
Q_FDP0 \ctrlR_REG[196] ( .CK(uclk), .D(n397), .Q(ctrlR[196]), .QN( ));
Q_FDP0 \ctrlR_REG[195] ( .CK(uclk), .D(n398), .Q(ctrlR[195]), .QN( ));
Q_FDP0 \ctrlR_REG[194] ( .CK(uclk), .D(n399), .Q(ctrlR[194]), .QN( ));
Q_FDP0 \ctrlR_REG[193] ( .CK(uclk), .D(n400), .Q(ctrlR[193]), .QN( ));
Q_FDP0 \ctrlR_REG[192] ( .CK(uclk), .D(n401), .Q(ctrlR[192]), .QN( ));
Q_FDP0 \ctrlR_REG[191] ( .CK(uclk), .D(n402), .Q(ctrlR[191]), .QN( ));
Q_FDP0 \ctrlR_REG[190] ( .CK(uclk), .D(n403), .Q(ctrlR[190]), .QN( ));
Q_FDP0 \ctrlR_REG[189] ( .CK(uclk), .D(n404), .Q(ctrlR[189]), .QN( ));
Q_FDP0 \ctrlR_REG[188] ( .CK(uclk), .D(n405), .Q(ctrlR[188]), .QN( ));
Q_FDP0 \ctrlR_REG[187] ( .CK(uclk), .D(n406), .Q(ctrlR[187]), .QN( ));
Q_FDP0 \ctrlR_REG[186] ( .CK(uclk), .D(n407), .Q(ctrlR[186]), .QN( ));
Q_FDP0 \ctrlR_REG[185] ( .CK(uclk), .D(n408), .Q(ctrlR[185]), .QN( ));
Q_FDP0 \ctrlR_REG[184] ( .CK(uclk), .D(n409), .Q(ctrlR[184]), .QN( ));
Q_FDP0 \ctrlR_REG[183] ( .CK(uclk), .D(n410), .Q(ctrlR[183]), .QN( ));
Q_FDP0 \ctrlR_REG[182] ( .CK(uclk), .D(n411), .Q(ctrlR[182]), .QN( ));
Q_FDP0 \ctrlR_REG[181] ( .CK(uclk), .D(n412), .Q(ctrlR[181]), .QN( ));
Q_FDP0 \ctrlR_REG[180] ( .CK(uclk), .D(n413), .Q(ctrlR[180]), .QN( ));
Q_FDP0 \ctrlR_REG[179] ( .CK(uclk), .D(n414), .Q(ctrlR[179]), .QN( ));
Q_FDP0 \ctrlR_REG[178] ( .CK(uclk), .D(n415), .Q(ctrlR[178]), .QN( ));
Q_FDP0 \ctrlR_REG[177] ( .CK(uclk), .D(n416), .Q(ctrlR[177]), .QN( ));
Q_FDP0 \ctrlR_REG[176] ( .CK(uclk), .D(n417), .Q(ctrlR[176]), .QN( ));
Q_FDP0 \ctrlR_REG[175] ( .CK(uclk), .D(n418), .Q(ctrlR[175]), .QN( ));
Q_FDP0 \ctrlR_REG[174] ( .CK(uclk), .D(n419), .Q(ctrlR[174]), .QN( ));
Q_FDP0 \ctrlR_REG[173] ( .CK(uclk), .D(n420), .Q(ctrlR[173]), .QN( ));
Q_FDP0 \ctrlR_REG[172] ( .CK(uclk), .D(n421), .Q(ctrlR[172]), .QN( ));
Q_FDP0 \ctrlR_REG[171] ( .CK(uclk), .D(n422), .Q(ctrlR[171]), .QN( ));
Q_FDP0 \ctrlR_REG[170] ( .CK(uclk), .D(n423), .Q(ctrlR[170]), .QN( ));
Q_FDP0 \ctrlR_REG[169] ( .CK(uclk), .D(n424), .Q(ctrlR[169]), .QN( ));
Q_FDP0 \ctrlR_REG[168] ( .CK(uclk), .D(n425), .Q(ctrlR[168]), .QN( ));
Q_FDP0 \ctrlR_REG[167] ( .CK(uclk), .D(n426), .Q(ctrlR[167]), .QN( ));
Q_FDP0 \ctrlR_REG[166] ( .CK(uclk), .D(n427), .Q(ctrlR[166]), .QN( ));
Q_FDP0 \ctrlR_REG[165] ( .CK(uclk), .D(n428), .Q(ctrlR[165]), .QN( ));
Q_FDP0 \ctrlR_REG[164] ( .CK(uclk), .D(n429), .Q(ctrlR[164]), .QN( ));
Q_FDP0 \ctrlR_REG[163] ( .CK(uclk), .D(n430), .Q(ctrlR[163]), .QN( ));
Q_FDP0 \ctrlR_REG[162] ( .CK(uclk), .D(n431), .Q(ctrlR[162]), .QN( ));
Q_FDP0 \ctrlR_REG[161] ( .CK(uclk), .D(n432), .Q(ctrlR[161]), .QN( ));
Q_FDP0 \ctrlR_REG[160] ( .CK(uclk), .D(n433), .Q(ctrlR[160]), .QN( ));
Q_FDP0 \ctrlR_REG[159] ( .CK(uclk), .D(n434), .Q(ctrlR[159]), .QN( ));
Q_FDP0 \ctrlR_REG[158] ( .CK(uclk), .D(n435), .Q(ctrlR[158]), .QN( ));
Q_FDP0 \ctrlR_REG[157] ( .CK(uclk), .D(n436), .Q(ctrlR[157]), .QN( ));
Q_FDP0 \ctrlR_REG[156] ( .CK(uclk), .D(n437), .Q(ctrlR[156]), .QN( ));
Q_FDP0 \ctrlR_REG[155] ( .CK(uclk), .D(n438), .Q(ctrlR[155]), .QN( ));
Q_FDP0 \ctrlR_REG[154] ( .CK(uclk), .D(n439), .Q(ctrlR[154]), .QN( ));
Q_FDP0 \ctrlR_REG[153] ( .CK(uclk), .D(n440), .Q(ctrlR[153]), .QN( ));
Q_FDP0 \ctrlR_REG[152] ( .CK(uclk), .D(n441), .Q(ctrlR[152]), .QN( ));
Q_FDP0 \ctrlR_REG[151] ( .CK(uclk), .D(n442), .Q(ctrlR[151]), .QN( ));
Q_FDP0 \ctrlR_REG[150] ( .CK(uclk), .D(n443), .Q(ctrlR[150]), .QN( ));
Q_FDP0 \ctrlR_REG[149] ( .CK(uclk), .D(n444), .Q(ctrlR[149]), .QN( ));
Q_FDP0 \ctrlR_REG[148] ( .CK(uclk), .D(n445), .Q(ctrlR[148]), .QN( ));
Q_FDP0 \ctrlR_REG[147] ( .CK(uclk), .D(n446), .Q(ctrlR[147]), .QN( ));
Q_FDP0 \ctrlR_REG[146] ( .CK(uclk), .D(n447), .Q(ctrlR[146]), .QN( ));
Q_FDP0 \ctrlR_REG[145] ( .CK(uclk), .D(n448), .Q(ctrlR[145]), .QN( ));
Q_FDP0 \ctrlR_REG[144] ( .CK(uclk), .D(n449), .Q(ctrlR[144]), .QN( ));
Q_FDP0 \ctrlR_REG[143] ( .CK(uclk), .D(n450), .Q(ctrlR[143]), .QN( ));
Q_FDP0 \ctrlR_REG[142] ( .CK(uclk), .D(n451), .Q(ctrlR[142]), .QN( ));
Q_FDP0 \ctrlR_REG[141] ( .CK(uclk), .D(n452), .Q(ctrlR[141]), .QN( ));
Q_FDP0 \ctrlR_REG[140] ( .CK(uclk), .D(n453), .Q(ctrlR[140]), .QN( ));
Q_FDP0 \ctrlR_REG[139] ( .CK(uclk), .D(n454), .Q(ctrlR[139]), .QN( ));
Q_FDP0 \ctrlR_REG[138] ( .CK(uclk), .D(n455), .Q(ctrlR[138]), .QN( ));
Q_FDP0 \ctrlR_REG[137] ( .CK(uclk), .D(n456), .Q(ctrlR[137]), .QN( ));
Q_FDP0 \ctrlR_REG[136] ( .CK(uclk), .D(n457), .Q(ctrlR[136]), .QN( ));
Q_FDP0 \ctrlR_REG[135] ( .CK(uclk), .D(n458), .Q(ctrlR[135]), .QN( ));
Q_FDP0 \ctrlR_REG[134] ( .CK(uclk), .D(n459), .Q(ctrlR[134]), .QN( ));
Q_FDP0 \ctrlR_REG[133] ( .CK(uclk), .D(n460), .Q(ctrlR[133]), .QN( ));
Q_FDP0 \ctrlR_REG[132] ( .CK(uclk), .D(n461), .Q(ctrlR[132]), .QN( ));
Q_FDP0 \ctrlR_REG[131] ( .CK(uclk), .D(n462), .Q(ctrlR[131]), .QN( ));
Q_FDP0 \ctrlR_REG[130] ( .CK(uclk), .D(n463), .Q(ctrlR[130]), .QN( ));
Q_FDP0 \ctrlR_REG[129] ( .CK(uclk), .D(n464), .Q(ctrlR[129]), .QN( ));
Q_FDP0 \ctrlR_REG[128] ( .CK(uclk), .D(n465), .Q(ctrlR[128]), .QN( ));
Q_FDP0 \ctrlR_REG[127] ( .CK(uclk), .D(n466), .Q(ctrlR[127]), .QN( ));
Q_FDP0 \ctrlR_REG[126] ( .CK(uclk), .D(n467), .Q(ctrlR[126]), .QN( ));
Q_FDP0 \ctrlR_REG[125] ( .CK(uclk), .D(n468), .Q(ctrlR[125]), .QN( ));
Q_FDP0 \ctrlR_REG[124] ( .CK(uclk), .D(n469), .Q(ctrlR[124]), .QN( ));
Q_FDP0 \ctrlR_REG[123] ( .CK(uclk), .D(n470), .Q(ctrlR[123]), .QN( ));
Q_FDP0 \ctrlR_REG[122] ( .CK(uclk), .D(n471), .Q(ctrlR[122]), .QN( ));
Q_FDP0 \ctrlR_REG[121] ( .CK(uclk), .D(n472), .Q(ctrlR[121]), .QN( ));
Q_FDP0 \ctrlR_REG[120] ( .CK(uclk), .D(n473), .Q(ctrlR[120]), .QN( ));
Q_FDP0 \ctrlR_REG[119] ( .CK(uclk), .D(n474), .Q(ctrlR[119]), .QN( ));
Q_FDP0 \ctrlR_REG[118] ( .CK(uclk), .D(n475), .Q(ctrlR[118]), .QN( ));
Q_FDP0 \ctrlR_REG[117] ( .CK(uclk), .D(n476), .Q(ctrlR[117]), .QN( ));
Q_FDP0 \ctrlR_REG[116] ( .CK(uclk), .D(n477), .Q(ctrlR[116]), .QN( ));
Q_FDP0 \ctrlR_REG[115] ( .CK(uclk), .D(n478), .Q(ctrlR[115]), .QN( ));
Q_FDP0 \ctrlR_REG[114] ( .CK(uclk), .D(n479), .Q(ctrlR[114]), .QN( ));
Q_FDP0 \ctrlR_REG[113] ( .CK(uclk), .D(n480), .Q(ctrlR[113]), .QN( ));
Q_FDP0 \ctrlR_REG[112] ( .CK(uclk), .D(n481), .Q(ctrlR[112]), .QN( ));
Q_FDP0 \ctrlR_REG[111] ( .CK(uclk), .D(n482), .Q(ctrlR[111]), .QN( ));
Q_FDP0 \ctrlR_REG[110] ( .CK(uclk), .D(n483), .Q(ctrlR[110]), .QN( ));
Q_FDP0 \ctrlR_REG[109] ( .CK(uclk), .D(n484), .Q(ctrlR[109]), .QN( ));
Q_FDP0 \ctrlR_REG[108] ( .CK(uclk), .D(n485), .Q(ctrlR[108]), .QN( ));
Q_FDP0 \ctrlR_REG[107] ( .CK(uclk), .D(n486), .Q(ctrlR[107]), .QN( ));
Q_FDP0 \ctrlR_REG[106] ( .CK(uclk), .D(n487), .Q(ctrlR[106]), .QN( ));
Q_FDP0 \ctrlR_REG[105] ( .CK(uclk), .D(n488), .Q(ctrlR[105]), .QN( ));
Q_FDP0 \ctrlR_REG[104] ( .CK(uclk), .D(n489), .Q(ctrlR[104]), .QN( ));
Q_FDP0 \ctrlR_REG[103] ( .CK(uclk), .D(n490), .Q(ctrlR[103]), .QN( ));
Q_FDP0 \ctrlR_REG[102] ( .CK(uclk), .D(n491), .Q(ctrlR[102]), .QN( ));
Q_FDP0 \ctrlR_REG[101] ( .CK(uclk), .D(n492), .Q(ctrlR[101]), .QN( ));
Q_FDP0 \ctrlR_REG[100] ( .CK(uclk), .D(n493), .Q(ctrlR[100]), .QN( ));
Q_FDP0 \ctrlR_REG[99] ( .CK(uclk), .D(n494), .Q(ctrlR[99]), .QN( ));
Q_FDP0 \ctrlR_REG[98] ( .CK(uclk), .D(n495), .Q(ctrlR[98]), .QN( ));
Q_FDP0 \ctrlR_REG[97] ( .CK(uclk), .D(n496), .Q(ctrlR[97]), .QN( ));
Q_FDP0 \ctrlR_REG[96] ( .CK(uclk), .D(n497), .Q(ctrlR[96]), .QN( ));
Q_FDP0 \ctrlR_REG[95] ( .CK(uclk), .D(n498), .Q(ctrlR[95]), .QN( ));
Q_FDP0 \ctrlR_REG[94] ( .CK(uclk), .D(n499), .Q(ctrlR[94]), .QN( ));
Q_FDP0 \ctrlR_REG[93] ( .CK(uclk), .D(n500), .Q(ctrlR[93]), .QN( ));
Q_FDP0 \ctrlR_REG[92] ( .CK(uclk), .D(n501), .Q(ctrlR[92]), .QN( ));
Q_FDP0 \ctrlR_REG[91] ( .CK(uclk), .D(n502), .Q(ctrlR[91]), .QN( ));
Q_FDP0 \ctrlR_REG[90] ( .CK(uclk), .D(n503), .Q(ctrlR[90]), .QN( ));
Q_FDP0 \ctrlR_REG[89] ( .CK(uclk), .D(n504), .Q(ctrlR[89]), .QN( ));
Q_FDP0 \ctrlR_REG[88] ( .CK(uclk), .D(n505), .Q(ctrlR[88]), .QN( ));
Q_FDP0 \ctrlR_REG[87] ( .CK(uclk), .D(n506), .Q(ctrlR[87]), .QN( ));
Q_FDP0 \ctrlR_REG[86] ( .CK(uclk), .D(n507), .Q(ctrlR[86]), .QN( ));
Q_FDP0 \ctrlR_REG[85] ( .CK(uclk), .D(n508), .Q(ctrlR[85]), .QN( ));
Q_FDP0 \ctrlR_REG[84] ( .CK(uclk), .D(n509), .Q(ctrlR[84]), .QN( ));
Q_FDP0 \ctrlR_REG[83] ( .CK(uclk), .D(n510), .Q(ctrlR[83]), .QN( ));
Q_FDP0 \ctrlR_REG[82] ( .CK(uclk), .D(n511), .Q(ctrlR[82]), .QN( ));
Q_FDP0 \ctrlR_REG[81] ( .CK(uclk), .D(n512), .Q(ctrlR[81]), .QN( ));
Q_FDP0 \ctrlR_REG[80] ( .CK(uclk), .D(n513), .Q(ctrlR[80]), .QN( ));
Q_FDP0 \ctrlR_REG[79] ( .CK(uclk), .D(n514), .Q(ctrlR[79]), .QN( ));
Q_FDP0 \ctrlR_REG[78] ( .CK(uclk), .D(n515), .Q(ctrlR[78]), .QN( ));
Q_FDP0 \ctrlR_REG[77] ( .CK(uclk), .D(n516), .Q(ctrlR[77]), .QN( ));
Q_FDP0 \ctrlR_REG[76] ( .CK(uclk), .D(n517), .Q(ctrlR[76]), .QN( ));
Q_FDP0 \ctrlR_REG[75] ( .CK(uclk), .D(n518), .Q(ctrlR[75]), .QN( ));
Q_FDP0 \ctrlR_REG[74] ( .CK(uclk), .D(n519), .Q(ctrlR[74]), .QN( ));
Q_FDP0 \ctrlR_REG[73] ( .CK(uclk), .D(n520), .Q(ctrlR[73]), .QN( ));
Q_FDP0 \ctrlR_REG[72] ( .CK(uclk), .D(n521), .Q(ctrlR[72]), .QN( ));
Q_FDP0 \ctrlR_REG[71] ( .CK(uclk), .D(n522), .Q(ctrlR[71]), .QN( ));
Q_FDP0 \ctrlR_REG[70] ( .CK(uclk), .D(n523), .Q(ctrlR[70]), .QN( ));
Q_FDP0 \ctrlR_REG[69] ( .CK(uclk), .D(n524), .Q(ctrlR[69]), .QN( ));
Q_FDP0 \ctrlR_REG[68] ( .CK(uclk), .D(n525), .Q(ctrlR[68]), .QN( ));
Q_FDP0 \ctrlR_REG[67] ( .CK(uclk), .D(n526), .Q(ctrlR[67]), .QN( ));
Q_FDP0 \ctrlR_REG[66] ( .CK(uclk), .D(n527), .Q(ctrlR[66]), .QN( ));
Q_FDP0 \ctrlR_REG[65] ( .CK(uclk), .D(n528), .Q(ctrlR[65]), .QN( ));
Q_FDP0 \ctrlR_REG[64] ( .CK(uclk), .D(n529), .Q(ctrlR[64]), .QN( ));
Q_FDP0 \ctrlR_REG[63] ( .CK(uclk), .D(n530), .Q(ctrlR[63]), .QN( ));
Q_FDP0 \ctrlR_REG[62] ( .CK(uclk), .D(n531), .Q(ctrlR[62]), .QN( ));
Q_FDP0 \ctrlR_REG[61] ( .CK(uclk), .D(n532), .Q(ctrlR[61]), .QN( ));
Q_FDP0 \ctrlR_REG[60] ( .CK(uclk), .D(n533), .Q(ctrlR[60]), .QN( ));
Q_FDP0 \ctrlR_REG[59] ( .CK(uclk), .D(n534), .Q(ctrlR[59]), .QN( ));
Q_FDP0 \ctrlR_REG[58] ( .CK(uclk), .D(n535), .Q(ctrlR[58]), .QN( ));
Q_FDP0 \ctrlR_REG[57] ( .CK(uclk), .D(n536), .Q(ctrlR[57]), .QN( ));
Q_FDP0 \ctrlR_REG[56] ( .CK(uclk), .D(n537), .Q(ctrlR[56]), .QN( ));
Q_FDP0 \ctrlR_REG[55] ( .CK(uclk), .D(n538), .Q(ctrlR[55]), .QN( ));
Q_FDP0 \ctrlR_REG[54] ( .CK(uclk), .D(n539), .Q(ctrlR[54]), .QN( ));
Q_FDP0 \ctrlR_REG[53] ( .CK(uclk), .D(n540), .Q(ctrlR[53]), .QN( ));
Q_FDP0 \ctrlR_REG[52] ( .CK(uclk), .D(n541), .Q(ctrlR[52]), .QN( ));
Q_FDP0 \ctrlR_REG[51] ( .CK(uclk), .D(n542), .Q(ctrlR[51]), .QN( ));
Q_FDP0 \ctrlR_REG[50] ( .CK(uclk), .D(n543), .Q(ctrlR[50]), .QN( ));
Q_FDP0 \ctrlR_REG[49] ( .CK(uclk), .D(n544), .Q(ctrlR[49]), .QN( ));
Q_FDP0 \ctrlR_REG[48] ( .CK(uclk), .D(n545), .Q(ctrlR[48]), .QN( ));
Q_FDP0 \ctrlR_REG[47] ( .CK(uclk), .D(n546), .Q(ctrlR[47]), .QN( ));
Q_FDP0 \ctrlR_REG[46] ( .CK(uclk), .D(n547), .Q(ctrlR[46]), .QN( ));
Q_FDP0 \ctrlR_REG[45] ( .CK(uclk), .D(n548), .Q(ctrlR[45]), .QN( ));
Q_FDP0 \ctrlR_REG[44] ( .CK(uclk), .D(n549), .Q(ctrlR[44]), .QN( ));
Q_FDP0 \ctrlR_REG[43] ( .CK(uclk), .D(n550), .Q(ctrlR[43]), .QN( ));
Q_FDP0 \ctrlR_REG[42] ( .CK(uclk), .D(n551), .Q(ctrlR[42]), .QN( ));
Q_FDP0 \ctrlR_REG[41] ( .CK(uclk), .D(n552), .Q(ctrlR[41]), .QN( ));
Q_FDP0 \ctrlR_REG[40] ( .CK(uclk), .D(n553), .Q(ctrlR[40]), .QN( ));
Q_FDP0 \ctrlR_REG[39] ( .CK(uclk), .D(n554), .Q(ctrlR[39]), .QN( ));
Q_FDP0 \ctrlR_REG[38] ( .CK(uclk), .D(n555), .Q(ctrlR[38]), .QN( ));
Q_FDP0 \ctrlR_REG[37] ( .CK(uclk), .D(n556), .Q(ctrlR[37]), .QN( ));
Q_FDP0 \ctrlR_REG[36] ( .CK(uclk), .D(n557), .Q(ctrlR[36]), .QN( ));
Q_FDP0 \ctrlR_REG[35] ( .CK(uclk), .D(n558), .Q(ctrlR[35]), .QN( ));
Q_FDP0 \ctrlR_REG[34] ( .CK(uclk), .D(n559), .Q(ctrlR[34]), .QN( ));
Q_FDP0 \ctrlR_REG[33] ( .CK(uclk), .D(n560), .Q(ctrlR[33]), .QN( ));
Q_FDP0 \ctrlR_REG[32] ( .CK(uclk), .D(n561), .Q(ctrlR[32]), .QN( ));
Q_FDP0 \ctrlR_REG[31] ( .CK(uclk), .D(n562), .Q(ctrlR[31]), .QN( ));
Q_FDP0 \ctrlR_REG[30] ( .CK(uclk), .D(n563), .Q(ctrlR[30]), .QN( ));
Q_FDP0 \ctrlR_REG[29] ( .CK(uclk), .D(n564), .Q(ctrlR[29]), .QN( ));
Q_FDP0 \ctrlR_REG[28] ( .CK(uclk), .D(n565), .Q(ctrlR[28]), .QN( ));
Q_FDP0 \ctrlR_REG[27] ( .CK(uclk), .D(n566), .Q(ctrlR[27]), .QN( ));
Q_FDP0 \ctrlR_REG[26] ( .CK(uclk), .D(n567), .Q(ctrlR[26]), .QN( ));
Q_FDP0 \ctrlR_REG[25] ( .CK(uclk), .D(n568), .Q(ctrlR[25]), .QN( ));
Q_FDP0 \ctrlR_REG[24] ( .CK(uclk), .D(n569), .Q(ctrlR[24]), .QN( ));
Q_FDP0 \ctrlR_REG[23] ( .CK(uclk), .D(n570), .Q(ctrlR[23]), .QN( ));
Q_FDP0 \ctrlR_REG[22] ( .CK(uclk), .D(n571), .Q(ctrlR[22]), .QN( ));
Q_FDP0 \ctrlR_REG[21] ( .CK(uclk), .D(n572), .Q(ctrlR[21]), .QN( ));
Q_FDP0 \ctrlR_REG[20] ( .CK(uclk), .D(n573), .Q(ctrlR[20]), .QN( ));
Q_FDP0 \ctrlR_REG[19] ( .CK(uclk), .D(n574), .Q(ctrlR[19]), .QN( ));
Q_FDP0 \ctrlR_REG[18] ( .CK(uclk), .D(n575), .Q(ctrlR[18]), .QN( ));
Q_FDP0 \ctrlR_REG[17] ( .CK(uclk), .D(n576), .Q(ctrlR[17]), .QN( ));
Q_FDP0 \ctrlR_REG[16] ( .CK(uclk), .D(n577), .Q(ctrlR[16]), .QN( ));
Q_FDP0 \ctrlR_REG[15] ( .CK(uclk), .D(n578), .Q(ctrlR[15]), .QN( ));
Q_FDP0 \ctrlR_REG[14] ( .CK(uclk), .D(n579), .Q(ctrlR[14]), .QN( ));
Q_FDP0 \ctrlR_REG[13] ( .CK(uclk), .D(n580), .Q(ctrlR[13]), .QN( ));
Q_FDP0 \ctrlR_REG[12] ( .CK(uclk), .D(n581), .Q(ctrlR[12]), .QN( ));
Q_FDP0 \ctrlR_REG[11] ( .CK(uclk), .D(n582), .Q(ctrlR[11]), .QN( ));
Q_FDP0 \ctrlR_REG[10] ( .CK(uclk), .D(n583), .Q(ctrlR[10]), .QN( ));
Q_FDP0 \ctrlR_REG[9] ( .CK(uclk), .D(n584), .Q(ctrlR[9]), .QN( ));
Q_FDP0 \ctrlR_REG[8] ( .CK(uclk), .D(n585), .Q(ctrlR[8]), .QN( ));
Q_FDP0 \ctrlR_REG[7] ( .CK(uclk), .D(n586), .Q(ctrlR[7]), .QN( ));
Q_FDP0 \ctrlR_REG[6] ( .CK(uclk), .D(n587), .Q(ctrlR[6]), .QN( ));
Q_FDP0 \ctrlR_REG[5] ( .CK(uclk), .D(n588), .Q(ctrlR[5]), .QN( ));
Q_FDP0 \ctrlR_REG[4] ( .CK(uclk), .D(n589), .Q(ctrlR[4]), .QN( ));
Q_FDP0 \ctrlR_REG[3] ( .CK(uclk), .D(n590), .Q(ctrlR[3]), .QN( ));
Q_FDP0 \ctrlR_REG[2] ( .CK(uclk), .D(n591), .Q(ctrlR[2]), .QN( ));
Q_FDP0 \ctrlR_REG[1] ( .CK(uclk), .D(n592), .Q(ctrlR[1]), .QN( ));
Q_FDP0 \ctrlR_REG[0] ( .CK(uclk), .D(n593), .Q(ctrlR[0]), .QN( ));
Q_BUFZP U2001 ( .OE(busyOn), .A(n337), .Z(xcva_top.xc_top.ecmHoldBusy));
Q_BUFZP U2002 ( .OE(holdEcm), .A(n337), .Z(xcva_top.xc_top.holdEcmTb));
Q_NOT_TOUCH _zzqnthw ( .sig());
ixc_uClkGen ukg ( uclk);
`ifdef CBV

reg [255:0] ctrl [0:3];
initial begin: U2005
  integer i;
  for (i=0; i<=3; i=i+1) ctrl[i] =
`ifdef CBV_MEM_INIT1
  {256{1'b1}};
`else
  256'b0;
`endif
end
reg [255:0] n1743;
assign {n338, n339, n340, n341, n342, n343, n344,
n345, n346, n347, n348, n349, n350, n351, n352,
n353, n354, n355, n356, n357, n358, n359, n360,
n361, n362, n363, n364, n365, n366, n367, n368,
n369, n370, n371, n372, n373, n374, n375, n376,
n377, n378, n379, n380, n381, n382, n383, n384,
n385, n386, n387, n388, n389, n390, n391, n392,
n393, n394, n395, n396, n397, n398, n399, n400,
n401, n402, n403, n404, n405, n406, n407, n408,
n409, n410, n411, n412, n413, n414, n415, n416,
n417, n418, n419, n420, n421, n422, n423, n424,
n425, n426, n427, n428, n429, n430, n431, n432,
n433, n434, n435, n436, n437, n438, n439, n440,
n441, n442, n443, n444, n445, n446, n447, n448,
n449, n450, n451, n452, n453, n454, n455, n456,
n457, n458, n459, n460, n461, n462, n463, n464,
n465, n466, n467, n468, n469, n470, n471, n472,
n473, n474, n475, n476, n477, n478, n479, n480,
n481, n482, n483, n484, n485, n486, n487, n488,
n489, n490, n491, n492, n493, n494, n495, n496,
n497, n498, n499, n500, n501, n502, n503, n504,
n505, n506, n507, n508, n509, n510, n511, n512,
n513, n514, n515, n516, n517, n518, n519, n520,
n521, n522, n523, n524, n525, n526, n527, n528,
n529, n530, n531, n532, n533, n534, n535, n536,
n537, n538, n539, n540, n541, n542, n543, n544,
n545, n546, n547, n548, n549, n550, n551, n552,
n553, n554, n555, n556, n557, n558, n559, n560,
n561, n562, n563, n564, n565, n566, n567, n568,
n569, n570, n571, n572, n573, n574, n575, n576,
n577, n578, n579, n580, n581, n582, n583, n584,
n585, n586, n587, n588, n589, n590, n591, n592,
n593} = n1743; 
always @(n594 or n1741 or n1740 or n1739 or n1738
 or n1737 or n1736 or n1735 or n1734 or n1733 or n1732 or n1731 or n1730
 or n1729 or n1728 or n1727 or n1726 or n1725 or n1724 or n1723 or n1722
 or n1721 or n1720 or n1719 or n1718 or n1717 or n1716 or n1715 or n1714
 or n1713 or n1712 or n1711 or n1710 or n1709 or n1708 or n1707 or n1706
 or n1705 or n1704 or n1703 or n1702 or n1701 or n1700 or n1699 or n1698
 or n1697 or n1696 or n1695 or n1694 or n1693 or n1692 or n1691 or n1690
 or n1689 or n1688 or n1687 or n1686 or n1685 or n1684 or n1683 or n1682
 or n1681 or n1680 or n1679 or n1678 or n1677 or n1676 or n1675 or n1674
 or n1673 or n1672 or n1671 or n1670 or n1669 or n1668 or n1667 or n1666
 or n1665 or n1664 or n1663 or n1662 or n1661 or n1660 or n1659 or n1658
 or n1657 or n1656 or n1655 or n1654 or n1653 or n1652 or n1651 or n1650
 or n1649 or n1648 or n1647 or n1646 or n1645 or n1644 or n1643 or n1642
 or n1641 or n1640 or n1639 or n1638 or n1637 or n1636 or n1635 or n1634
 or n1633 or n1632 or n1631 or n1630 or n1629 or n1628 or n1627 or n1626
 or n1625 or n1624 or n1623 or n1622 or n1621 or n1620 or n1619 or n1618
 or n1617 or n1616 or n1615 or n1614 or n1613 or n1612 or n1611 or n1610
 or n1609 or n1608 or n1607 or n1606 or n1605 or n1604 or n1603 or n1602
 or n1601 or n1600 or n1599 or n1598 or n1597 or n1596 or n1595 or n1594
 or n1593 or n1592 or n1591 or n1590 or n1589 or n1588 or n1587 or n1586
 or n1585 or n1584 or n1583 or n1582 or n1581 or n1580 or n1579 or n1578
 or n1577 or n1576 or n1575 or n1574 or n1573 or n1572 or n1571 or n1570
 or n1569 or n1568 or n1567 or n1566 or n1565 or n1564 or n1563 or n1562
 or n1561 or n1560 or n1559 or n1558 or n1557 or n1556 or n1555 or n1554
 or n1553 or n1552 or n1551 or n1550 or n1549 or n1548 or n1547 or n1546
 or n1545 or n1544 or n1543 or n1542 or n1541 or n1540 or n1539 or n1538
 or n1537 or n1536 or n1535 or n1534 or n1533 or n1532 or n1531 or n1530
 or n1529 or n1528 or n1527 or n1526 or n1525 or n1524 or n1523 or n1522
 or n1521 or n1520 or n1519 or n1518 or n1517 or n1516 or n1515 or n1514
 or n1513 or n1512 or n1511 or n1510 or n1509 or n1508 or n1507 or n1506
 or n1505 or n1504 or n1503 or n1502 or n1501 or n1500 or n1499 or n1498
 or n1497 or n1496 or n1495 or n1494 or n1493 or n1492 or n1491 or n1490
 or n1489 or n1488 or n1487 or n1486 or n1485 or n337)
#0 begin
if (n1485)
ctrl[{n594, n594}] =
{n1741, n1740, n1739, n1738, n1737,
 n1736, n1735, n1734, n1733, n1732, n1731, n1730, n1729,
 n1728, n1727, n1726, n1725, n1724, n1723, n1722, n1721,
 n1720, n1719, n1718, n1717, n1716, n1715, n1714, n1713,
 n1712, n1711, n1710, n1709, n1708, n1707, n1706, n1705,
 n1704, n1703, n1702, n1701, n1700, n1699, n1698, n1697,
 n1696, n1695, n1694, n1693, n1692, n1691, n1690, n1689,
 n1688, n1687, n1686, n1685, n1684, n1683, n1682, n1681,
 n1680, n1679, n1678, n1677, n1676, n1675, n1674, n1673,
 n1672, n1671, n1670, n1669, n1668, n1667, n1666, n1665,
 n1664, n1663, n1662, n1661, n1660, n1659, n1658, n1657,
 n1656, n1655, n1654, n1653, n1652, n1651, n1650, n1649,
 n1648, n1647, n1646, n1645, n1644, n1643, n1642, n1641,
 n1640, n1639, n1638, n1637, n1636, n1635, n1634, n1633,
 n1632, n1631, n1630, n1629, n1628, n1627, n1626, n1625,
 n1624, n1623, n1622, n1621, n1620, n1619, n1618, n1617,
 n1616, n1615, n1614, n1613, n1612, n1611, n1610, n1609,
 n1608, n1607, n1606, n1605, n1604, n1603, n1602, n1601,
 n1600, n1599, n1598, n1597, n1596, n1595, n1594, n1593,
 n1592, n1591, n1590, n1589, n1588, n1587, n1586, n1585,
 n1584, n1583, n1582, n1581, n1580, n1579, n1578, n1577,
 n1576, n1575, n1574, n1573, n1572, n1571, n1570, n1569,
 n1568, n1567, n1566, n1565, n1564, n1563, n1562, n1561,
 n1560, n1559, n1558, n1557, n1556, n1555, n1554, n1553,
 n1552, n1551, n1550, n1549, n1548, n1547, n1546, n1545,
 n1544, n1543, n1542, n1541, n1540, n1539, n1538, n1537,
 n1536, n1535, n1534, n1533, n1532, n1531, n1530, n1529,
 n1528, n1527, n1526, n1525, n1524, n1523, n1522, n1521,
 n1520, n1519, n1518, n1517, n1516, n1515, n1514, n1513,
 n1512, n1511, n1510, n1509, n1508, n1507, n1506, n1505,
 n1504, n1503, n1502, n1501, n1500, n1499, n1498, n1497,
 n1496, n1495, n1494, n1493, n1492, n1491, n1490, n1489,
 n1488, n1487, n1486};
n1743 = ctrl[{n594, n337}];
end
`else

MPW4X256 ctrl ( .A1(n594), .A0(n594), .DI255(n1741), .DI254(n1740), .DI253(n1739), .DI252(n1738),
 .DI251(n1737), .DI250(n1736), .DI249(n1735), .DI248(n1734), .DI247(n1733), .DI246(n1732), .DI245(n1731), .DI244(n1730),
 .DI243(n1729), .DI242(n1728), .DI241(n1727), .DI240(n1726), .DI239(n1725), .DI238(n1724), .DI237(n1723), .DI236(n1722),
 .DI235(n1721), .DI234(n1720), .DI233(n1719), .DI232(n1718), .DI231(n1717), .DI230(n1716), .DI229(n1715), .DI228(n1714),
 .DI227(n1713), .DI226(n1712), .DI225(n1711), .DI224(n1710), .DI223(n1709), .DI222(n1708), .DI221(n1707), .DI220(n1706),
 .DI219(n1705), .DI218(n1704), .DI217(n1703), .DI216(n1702), .DI215(n1701), .DI214(n1700), .DI213(n1699), .DI212(n1698),
 .DI211(n1697), .DI210(n1696), .DI209(n1695), .DI208(n1694), .DI207(n1693), .DI206(n1692), .DI205(n1691), .DI204(n1690),
 .DI203(n1689), .DI202(n1688), .DI201(n1687), .DI200(n1686), .DI199(n1685), .DI198(n1684), .DI197(n1683), .DI196(n1682),
 .DI195(n1681), .DI194(n1680), .DI193(n1679), .DI192(n1678), .DI191(n1677), .DI190(n1676), .DI189(n1675), .DI188(n1674),
 .DI187(n1673), .DI186(n1672), .DI185(n1671), .DI184(n1670), .DI183(n1669), .DI182(n1668), .DI181(n1667), .DI180(n1666),
 .DI179(n1665), .DI178(n1664), .DI177(n1663), .DI176(n1662), .DI175(n1661), .DI174(n1660), .DI173(n1659), .DI172(n1658),
 .DI171(n1657), .DI170(n1656), .DI169(n1655), .DI168(n1654), .DI167(n1653), .DI166(n1652), .DI165(n1651), .DI164(n1650),
 .DI163(n1649), .DI162(n1648), .DI161(n1647), .DI160(n1646), .DI159(n1645), .DI158(n1644), .DI157(n1643), .DI156(n1642),
 .DI155(n1641), .DI154(n1640), .DI153(n1639), .DI152(n1638), .DI151(n1637), .DI150(n1636), .DI149(n1635), .DI148(n1634),
 .DI147(n1633), .DI146(n1632), .DI145(n1631), .DI144(n1630), .DI143(n1629), .DI142(n1628), .DI141(n1627), .DI140(n1626),
 .DI139(n1625), .DI138(n1624), .DI137(n1623), .DI136(n1622), .DI135(n1621), .DI134(n1620), .DI133(n1619), .DI132(n1618),
 .DI131(n1617), .DI130(n1616), .DI129(n1615), .DI128(n1614), .DI127(n1613), .DI126(n1612), .DI125(n1611), .DI124(n1610),
 .DI123(n1609), .DI122(n1608), .DI121(n1607), .DI120(n1606), .DI119(n1605), .DI118(n1604), .DI117(n1603), .DI116(n1602),
 .DI115(n1601), .DI114(n1600), .DI113(n1599), .DI112(n1598), .DI111(n1597), .DI110(n1596), .DI109(n1595), .DI108(n1594),
 .DI107(n1593), .DI106(n1592), .DI105(n1591), .DI104(n1590), .DI103(n1589), .DI102(n1588), .DI101(n1587), .DI100(n1586),
 .DI99(n1585), .DI98(n1584), .DI97(n1583), .DI96(n1582), .DI95(n1581), .DI94(n1580), .DI93(n1579), .DI92(n1578),
 .DI91(n1577), .DI90(n1576), .DI89(n1575), .DI88(n1574), .DI87(n1573), .DI86(n1572), .DI85(n1571), .DI84(n1570),
 .DI83(n1569), .DI82(n1568), .DI81(n1567), .DI80(n1566), .DI79(n1565), .DI78(n1564), .DI77(n1563), .DI76(n1562),
 .DI75(n1561), .DI74(n1560), .DI73(n1559), .DI72(n1558), .DI71(n1557), .DI70(n1556), .DI69(n1555), .DI68(n1554),
 .DI67(n1553), .DI66(n1552), .DI65(n1551), .DI64(n1550), .DI63(n1549), .DI62(n1548), .DI61(n1547), .DI60(n1546),
 .DI59(n1545), .DI58(n1544), .DI57(n1543), .DI56(n1542), .DI55(n1541), .DI54(n1540), .DI53(n1539), .DI52(n1538),
 .DI51(n1537), .DI50(n1536), .DI49(n1535), .DI48(n1534), .DI47(n1533), .DI46(n1532), .DI45(n1531), .DI44(n1530),
 .DI43(n1529), .DI42(n1528), .DI41(n1527), .DI40(n1526), .DI39(n1525), .DI38(n1524), .DI37(n1523), .DI36(n1522),
 .DI35(n1521), .DI34(n1520), .DI33(n1519), .DI32(n1518), .DI31(n1517), .DI30(n1516), .DI29(n1515), .DI28(n1514),
 .DI27(n1513), .DI26(n1512), .DI25(n1511), .DI24(n1510), .DI23(n1509), .DI22(n1508), .DI21(n1507), .DI20(n1506),
 .DI19(n1505), .DI18(n1504), .DI17(n1503), .DI16(n1502), .DI15(n1501), .DI14(n1500), .DI13(n1499), .DI12(n1498),
 .DI11(n1497), .DI10(n1496), .DI9(n1495), .DI8(n1494), .DI7(n1493), .DI6(n1492), .DI5(n1491), .DI4(n1490),
 .DI3(n1489), .DI2(n1488), .DI1(n1487), .DI0(n1486), .WE(n1485), .SYNC_IN(n594), .SYNC_OUT(n1743));
// pragma CVASTRPROP INSTANCE "ctrl" HDL_MEMORY_DECL "1 255 0 0 3"
MPR4X256 U2006 ( .A1(n594), .A0(n337), .SYNC_IN(n1743), .DO255(n338), .DO254(n339), .DO253(n340),
 .DO252(n341), .DO251(n342), .DO250(n343), .DO249(n344), .DO248(n345), .DO247(n346), .DO246(n347), .DO245(n348),
 .DO244(n349), .DO243(n350), .DO242(n351), .DO241(n352), .DO240(n353), .DO239(n354), .DO238(n355), .DO237(n356),
 .DO236(n357), .DO235(n358), .DO234(n359), .DO233(n360), .DO232(n361), .DO231(n362), .DO230(n363), .DO229(n364),
 .DO228(n365), .DO227(n366), .DO226(n367), .DO225(n368), .DO224(n369), .DO223(n370), .DO222(n371), .DO221(n372),
 .DO220(n373), .DO219(n374), .DO218(n375), .DO217(n376), .DO216(n377), .DO215(n378), .DO214(n379), .DO213(n380),
 .DO212(n381), .DO211(n382), .DO210(n383), .DO209(n384), .DO208(n385), .DO207(n386), .DO206(n387), .DO205(n388),
 .DO204(n389), .DO203(n390), .DO202(n391), .DO201(n392), .DO200(n393), .DO199(n394), .DO198(n395), .DO197(n396),
 .DO196(n397), .DO195(n398), .DO194(n399), .DO193(n400), .DO192(n401), .DO191(n402), .DO190(n403), .DO189(n404),
 .DO188(n405), .DO187(n406), .DO186(n407), .DO185(n408), .DO184(n409), .DO183(n410), .DO182(n411), .DO181(n412),
 .DO180(n413), .DO179(n414), .DO178(n415), .DO177(n416), .DO176(n417), .DO175(n418), .DO174(n419), .DO173(n420),
 .DO172(n421), .DO171(n422), .DO170(n423), .DO169(n424), .DO168(n425), .DO167(n426), .DO166(n427), .DO165(n428),
 .DO164(n429), .DO163(n430), .DO162(n431), .DO161(n432), .DO160(n433), .DO159(n434), .DO158(n435), .DO157(n436),
 .DO156(n437), .DO155(n438), .DO154(n439), .DO153(n440), .DO152(n441), .DO151(n442), .DO150(n443), .DO149(n444),
 .DO148(n445), .DO147(n446), .DO146(n447), .DO145(n448), .DO144(n449), .DO143(n450), .DO142(n451), .DO141(n452),
 .DO140(n453), .DO139(n454), .DO138(n455), .DO137(n456), .DO136(n457), .DO135(n458), .DO134(n459), .DO133(n460),
 .DO132(n461), .DO131(n462), .DO130(n463), .DO129(n464), .DO128(n465), .DO127(n466), .DO126(n467), .DO125(n468),
 .DO124(n469), .DO123(n470), .DO122(n471), .DO121(n472), .DO120(n473), .DO119(n474), .DO118(n475), .DO117(n476),
 .DO116(n477), .DO115(n478), .DO114(n479), .DO113(n480), .DO112(n481), .DO111(n482), .DO110(n483), .DO109(n484),
 .DO108(n485), .DO107(n486), .DO106(n487), .DO105(n488), .DO104(n489), .DO103(n490), .DO102(n491), .DO101(n492),
 .DO100(n493), .DO99(n494), .DO98(n495), .DO97(n496), .DO96(n497), .DO95(n498), .DO94(n499), .DO93(n500),
 .DO92(n501), .DO91(n502), .DO90(n503), .DO89(n504), .DO88(n505), .DO87(n506), .DO86(n507), .DO85(n508),
 .DO84(n509), .DO83(n510), .DO82(n511), .DO81(n512), .DO80(n513), .DO79(n514), .DO78(n515), .DO77(n516),
 .DO76(n517), .DO75(n518), .DO74(n519), .DO73(n520), .DO72(n521), .DO71(n522), .DO70(n523), .DO69(n524),
 .DO68(n525), .DO67(n526), .DO66(n527), .DO65(n528), .DO64(n529), .DO63(n530), .DO62(n531), .DO61(n532),
 .DO60(n533), .DO59(n534), .DO58(n535), .DO57(n536), .DO56(n537), .DO55(n538), .DO54(n539), .DO53(n540),
 .DO52(n541), .DO51(n542), .DO50(n543), .DO49(n544), .DO48(n545), .DO47(n546), .DO46(n547), .DO45(n548),
 .DO44(n549), .DO43(n550), .DO42(n551), .DO41(n552), .DO40(n553), .DO39(n554), .DO38(n555), .DO37(n556),
 .DO36(n557), .DO35(n558), .DO34(n559), .DO33(n560), .DO32(n561), .DO31(n562), .DO30(n563), .DO29(n564),
 .DO28(n565), .DO27(n566), .DO26(n567), .DO25(n568), .DO24(n569), .DO23(n570), .DO22(n571), .DO21(n572),
 .DO20(n573), .DO19(n574), .DO18(n575), .DO17(n576), .DO16(n577), .DO15(n578), .DO14(n579), .DO13(n580),
 .DO12(n581), .DO11(n582), .DO10(n583), .DO9(n584), .DO8(n585), .DO7(n586), .DO6(n587), .DO5(n588),
 .DO4(n589), .DO3(n590), .DO2(n591), .DO1(n592), .DO0(n593), .SYNC_OUT( ));
`endif
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "ctrl 1 255 0 0 3"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "1"
// pragma CVASTRPROP MODULE HDLICE PROP_IXCOM_MOD TRUE
endmodule
`ifdef CBV
`else
`ifdef MPW4X256_MPR4X256
`else
module MPW4X256( A1, A0, DI255, DI254, DI253, DI252, DI251,
 DI250, DI249, DI248, DI247, DI246, DI245, DI244, DI243,
 DI242, DI241, DI240, DI239, DI238, DI237, DI236, DI235,
 DI234, DI233, DI232, DI231, DI230, DI229, DI228, DI227,
 DI226, DI225, DI224, DI223, DI222, DI221, DI220, DI219,
 DI218, DI217, DI216, DI215, DI214, DI213, DI212, DI211,
 DI210, DI209, DI208, DI207, DI206, DI205, DI204, DI203,
 DI202, DI201, DI200, DI199, DI198, DI197, DI196, DI195,
 DI194, DI193, DI192, DI191, DI190, DI189, DI188, DI187,
 DI186, DI185, DI184, DI183, DI182, DI181, DI180, DI179,
 DI178, DI177, DI176, DI175, DI174, DI173, DI172, DI171,
 DI170, DI169, DI168, DI167, DI166, DI165, DI164, DI163,
 DI162, DI161, DI160, DI159, DI158, DI157, DI156, DI155,
 DI154, DI153, DI152, DI151, DI150, DI149, DI148, DI147,
 DI146, DI145, DI144, DI143, DI142, DI141, DI140, DI139,
 DI138, DI137, DI136, DI135, DI134, DI133, DI132, DI131,
 DI130, DI129, DI128, DI127, DI126, DI125, DI124, DI123,
 DI122, DI121, DI120, DI119, DI118, DI117, DI116, DI115,
 DI114, DI113, DI112, DI111, DI110, DI109, DI108, DI107,
 DI106, DI105, DI104, DI103, DI102, DI101, DI100, DI99,
 DI98, DI97, DI96, DI95, DI94, DI93, DI92, DI91,
 DI90, DI89, DI88, DI87, DI86, DI85, DI84, DI83,
 DI82, DI81, DI80, DI79, DI78, DI77, DI76, DI75,
 DI74, DI73, DI72, DI71, DI70, DI69, DI68, DI67,
 DI66, DI65, DI64, DI63, DI62, DI61, DI60, DI59,
 DI58, DI57, DI56, DI55, DI54, DI53, DI52, DI51,
 DI50, DI49, DI48, DI47, DI46, DI45, DI44, DI43,
 DI42, DI41, DI40, DI39, DI38, DI37, DI36, DI35,
 DI34, DI33, DI32, DI31, DI30, DI29, DI28, DI27,
 DI26, DI25, DI24, DI23, DI22, DI21, DI20, DI19,
 DI18, DI17, DI16, DI15, DI14, DI13, DI12, DI11,
 DI10, DI9, DI8, DI7, DI6, DI5, DI4, DI3,
 DI2, DI1, DI0, WE, SYNC_IN, SYNC_OUT);
input  A1, A0, DI255, DI254, DI253, DI252, DI251, DI250,
 DI249, DI248, DI247, DI246, DI245, DI244, DI243, DI242, DI241, DI240,
 DI239, DI238, DI237, DI236, DI235, DI234, DI233, DI232, DI231, DI230,
 DI229, DI228, DI227, DI226, DI225, DI224, DI223, DI222, DI221, DI220,
 DI219, DI218, DI217, DI216, DI215, DI214, DI213, DI212, DI211, DI210,
 DI209, DI208, DI207, DI206, DI205, DI204, DI203, DI202, DI201, DI200,
 DI199, DI198, DI197, DI196, DI195, DI194, DI193, DI192, DI191, DI190,
 DI189, DI188, DI187, DI186, DI185, DI184, DI183, DI182, DI181, DI180,
 DI179, DI178, DI177, DI176, DI175, DI174, DI173, DI172, DI171, DI170,
 DI169, DI168, DI167, DI166, DI165, DI164, DI163, DI162, DI161, DI160,
 DI159, DI158, DI157, DI156, DI155, DI154, DI153, DI152, DI151, DI150,
 DI149, DI148, DI147, DI146, DI145, DI144, DI143, DI142, DI141, DI140,
 DI139, DI138, DI137, DI136, DI135, DI134, DI133, DI132, DI131, DI130,
 DI129, DI128, DI127, DI126, DI125, DI124, DI123, DI122, DI121, DI120,
 DI119, DI118, DI117, DI116, DI115, DI114, DI113, DI112, DI111, DI110,
 DI109, DI108, DI107, DI106, DI105, DI104, DI103, DI102, DI101, DI100,
 DI99, DI98, DI97, DI96, DI95, DI94, DI93, DI92, DI91, DI90,
 DI89, DI88, DI87, DI86, DI85, DI84, DI83, DI82, DI81, DI80,
 DI79, DI78, DI77, DI76, DI75, DI74, DI73, DI72, DI71, DI70,
 DI69, DI68, DI67, DI66, DI65, DI64, DI63, DI62, DI61, DI60,
 DI59, DI58, DI57, DI56, DI55, DI54, DI53, DI52, DI51, DI50,
 DI49, DI48, DI47, DI46, DI45, DI44, DI43, DI42, DI41, DI40,
 DI39, DI38, DI37, DI36, DI35, DI34, DI33, DI32, DI31, DI30,
 DI29, DI28, DI27, DI26, DI25, DI24, DI23, DI22, DI21, DI20,
 DI19, DI18, DI17, DI16, DI15, DI14, DI13, DI12, DI11, DI10,
 DI9, DI8, DI7, DI6, DI5, DI4, DI3, DI2, DI1, DI0,
 WE, SYNC_IN;
output  SYNC_OUT;
endmodule
`ifdef _MPR4X256_
`else
module MPR4X256( A1, A0, SYNC_IN, DO255, DO254, DO253, DO252,
 DO251, DO250, DO249, DO248, DO247, DO246, DO245, DO244,
 DO243, DO242, DO241, DO240, DO239, DO238, DO237, DO236,
 DO235, DO234, DO233, DO232, DO231, DO230, DO229, DO228,
 DO227, DO226, DO225, DO224, DO223, DO222, DO221, DO220,
 DO219, DO218, DO217, DO216, DO215, DO214, DO213, DO212,
 DO211, DO210, DO209, DO208, DO207, DO206, DO205, DO204,
 DO203, DO202, DO201, DO200, DO199, DO198, DO197, DO196,
 DO195, DO194, DO193, DO192, DO191, DO190, DO189, DO188,
 DO187, DO186, DO185, DO184, DO183, DO182, DO181, DO180,
 DO179, DO178, DO177, DO176, DO175, DO174, DO173, DO172,
 DO171, DO170, DO169, DO168, DO167, DO166, DO165, DO164,
 DO163, DO162, DO161, DO160, DO159, DO158, DO157, DO156,
 DO155, DO154, DO153, DO152, DO151, DO150, DO149, DO148,
 DO147, DO146, DO145, DO144, DO143, DO142, DO141, DO140,
 DO139, DO138, DO137, DO136, DO135, DO134, DO133, DO132,
 DO131, DO130, DO129, DO128, DO127, DO126, DO125, DO124,
 DO123, DO122, DO121, DO120, DO119, DO118, DO117, DO116,
 DO115, DO114, DO113, DO112, DO111, DO110, DO109, DO108,
 DO107, DO106, DO105, DO104, DO103, DO102, DO101, DO100,
 DO99, DO98, DO97, DO96, DO95, DO94, DO93, DO92,
 DO91, DO90, DO89, DO88, DO87, DO86, DO85, DO84,
 DO83, DO82, DO81, DO80, DO79, DO78, DO77, DO76,
 DO75, DO74, DO73, DO72, DO71, DO70, DO69, DO68,
 DO67, DO66, DO65, DO64, DO63, DO62, DO61, DO60,
 DO59, DO58, DO57, DO56, DO55, DO54, DO53, DO52,
 DO51, DO50, DO49, DO48, DO47, DO46, DO45, DO44,
 DO43, DO42, DO41, DO40, DO39, DO38, DO37, DO36,
 DO35, DO34, DO33, DO32, DO31, DO30, DO29, DO28,
 DO27, DO26, DO25, DO24, DO23, DO22, DO21, DO20,
 DO19, DO18, DO17, DO16, DO15, DO14, DO13, DO12,
 DO11, DO10, DO9, DO8, DO7, DO6, DO5, DO4,
 DO3, DO2, DO1, DO0, SYNC_OUT);
input  A1, A0, SYNC_IN;
output  DO255, DO254, DO253, DO252, DO251, DO250, DO249, DO248,
 DO247, DO246, DO245, DO244, DO243, DO242, DO241, DO240, DO239, DO238,
 DO237, DO236, DO235, DO234, DO233, DO232, DO231, DO230, DO229, DO228,
 DO227, DO226, DO225, DO224, DO223, DO222, DO221, DO220, DO219, DO218,
 DO217, DO216, DO215, DO214, DO213, DO212, DO211, DO210, DO209, DO208,
 DO207, DO206, DO205, DO204, DO203, DO202, DO201, DO200, DO199, DO198,
 DO197, DO196, DO195, DO194, DO193, DO192, DO191, DO190, DO189, DO188,
 DO187, DO186, DO185, DO184, DO183, DO182, DO181, DO180, DO179, DO178,
 DO177, DO176, DO175, DO174, DO173, DO172, DO171, DO170, DO169, DO168,
 DO167, DO166, DO165, DO164, DO163, DO162, DO161, DO160, DO159, DO158,
 DO157, DO156, DO155, DO154, DO153, DO152, DO151, DO150, DO149, DO148,
 DO147, DO146, DO145, DO144, DO143, DO142, DO141, DO140, DO139, DO138,
 DO137, DO136, DO135, DO134, DO133, DO132, DO131, DO130, DO129, DO128,
 DO127, DO126, DO125, DO124, DO123, DO122, DO121, DO120, DO119, DO118,
 DO117, DO116, DO115, DO114, DO113, DO112, DO111, DO110, DO109, DO108,
 DO107, DO106, DO105, DO104, DO103, DO102, DO101, DO100, DO99, DO98,
 DO97, DO96, DO95, DO94, DO93, DO92, DO91, DO90, DO89, DO88,
 DO87, DO86, DO85, DO84, DO83, DO82, DO81, DO80, DO79, DO78,
 DO77, DO76, DO75, DO74, DO73, DO72, DO71, DO70, DO69, DO68,
 DO67, DO66, DO65, DO64, DO63, DO62, DO61, DO60, DO59, DO58,
 DO57, DO56, DO55, DO54, DO53, DO52, DO51, DO50, DO49, DO48,
 DO47, DO46, DO45, DO44, DO43, DO42, DO41, DO40, DO39, DO38,
 DO37, DO36, DO35, DO34, DO33, DO32, DO31, DO30, DO29, DO28,
 DO27, DO26, DO25, DO24, DO23, DO22, DO21, DO20, DO19, DO18,
 DO17, DO16, DO15, DO14, DO13, DO12, DO11, DO10, DO9, DO8,
 DO7, DO6, DO5, DO4, DO3, DO2, DO1, DO0, SYNC_OUT;
endmodule
`define _MPR4X256_
`endif
`define MPW4X256_MPR4X256
`endif
`endif
