library ieee, quickturn ;
use ieee.std_logic_1164.all ;
use quickturn.verilog.all ;
entity _ixc_isc is
  attribute _2_state_: integer;
end _ixc_isc ;
