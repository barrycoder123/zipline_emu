library ieee, quickturn ;
use ieee.std_logic_1164.all ;
use quickturn.verilog.all ;
entity sfifo_conns_0 is
  attribute _2_state_: integer;
end sfifo_conns_0 ;
