
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
(* celldefine = 1 *) 
module nx_reg_indirect_access ( stat_code, stat_datawords, stat_addr, 
	capability_lst, capability_type, rd_dat, .mem_a( {\mem_a[0][31] , 
	\mem_a[0][30] , \mem_a[0][29] , \mem_a[0][28] , \mem_a[0][27] , 
	\mem_a[0][26] , \mem_a[0][25] , \mem_a[0][24] , \mem_a[0][23] , 
	\mem_a[0][22] , \mem_a[0][21] , \mem_a[0][20] , \mem_a[0][19] , 
	\mem_a[0][18] , \mem_a[0][17] , \mem_a[0][16] , \mem_a[0][15] , 
	\mem_a[0][14] , \mem_a[0][13] , \mem_a[0][12] , \mem_a[0][11] , 
	\mem_a[0][10] , \mem_a[0][9] , \mem_a[0][8] , \mem_a[0][7] , 
	\mem_a[0][6] , \mem_a[0][5] , \mem_a[0][4] , \mem_a[0][3] , 
	\mem_a[0][2] , \mem_a[0][1] , \mem_a[0][0] , \mem_a[1][31] , 
	\mem_a[1][30] , \mem_a[1][29] , \mem_a[1][28] , \mem_a[1][27] , 
	\mem_a[1][26] , \mem_a[1][25] , \mem_a[1][24] , \mem_a[1][23] , 
	\mem_a[1][22] , \mem_a[1][21] , \mem_a[1][20] , \mem_a[1][19] , 
	\mem_a[1][18] , \mem_a[1][17] , \mem_a[1][16] , \mem_a[1][15] , 
	\mem_a[1][14] , \mem_a[1][13] , \mem_a[1][12] , \mem_a[1][11] , 
	\mem_a[1][10] , \mem_a[1][9] , \mem_a[1][8] , \mem_a[1][7] , 
	\mem_a[1][6] , \mem_a[1][5] , \mem_a[1][4] , \mem_a[1][3] , 
	\mem_a[1][2] , \mem_a[1][1] , \mem_a[1][0] , \mem_a[2][31] , 
	\mem_a[2][30] , \mem_a[2][29] , \mem_a[2][28] , \mem_a[2][27] , 
	\mem_a[2][26] , \mem_a[2][25] , \mem_a[2][24] , \mem_a[2][23] , 
	\mem_a[2][22] , \mem_a[2][21] , \mem_a[2][20] , \mem_a[2][19] , 
	\mem_a[2][18] , \mem_a[2][17] , \mem_a[2][16] , \mem_a[2][15] , 
	\mem_a[2][14] , \mem_a[2][13] , \mem_a[2][12] , \mem_a[2][11] , 
	\mem_a[2][10] , \mem_a[2][9] , \mem_a[2][8] , \mem_a[2][7] , 
	\mem_a[2][6] , \mem_a[2][5] , \mem_a[2][4] , \mem_a[2][3] , 
	\mem_a[2][2] , \mem_a[2][1] , \mem_a[2][0] , \mem_a[3][31] , 
	\mem_a[3][30] , \mem_a[3][29] , \mem_a[3][28] , \mem_a[3][27] , 
	\mem_a[3][26] , \mem_a[3][25] , \mem_a[3][24] , \mem_a[3][23] , 
	\mem_a[3][22] , \mem_a[3][21] , \mem_a[3][20] , \mem_a[3][19] , 
	\mem_a[3][18] , \mem_a[3][17] , \mem_a[3][16] , \mem_a[3][15] , 
	\mem_a[3][14] , \mem_a[3][13] , \mem_a[3][12] , \mem_a[3][11] , 
	\mem_a[3][10] , \mem_a[3][9] , \mem_a[3][8] , \mem_a[3][7] , 
	\mem_a[3][6] , \mem_a[3][5] , \mem_a[3][4] , \mem_a[3][3] , 
	\mem_a[3][2] , \mem_a[3][1] , \mem_a[3][0] , \mem_a[4][31] , 
	\mem_a[4][30] , \mem_a[4][29] , \mem_a[4][28] , \mem_a[4][27] , 
	\mem_a[4][26] , \mem_a[4][25] , \mem_a[4][24] , \mem_a[4][23] , 
	\mem_a[4][22] , \mem_a[4][21] , \mem_a[4][20] , \mem_a[4][19] , 
	\mem_a[4][18] , \mem_a[4][17] , \mem_a[4][16] , \mem_a[4][15] , 
	\mem_a[4][14] , \mem_a[4][13] , \mem_a[4][12] , \mem_a[4][11] , 
	\mem_a[4][10] , \mem_a[4][9] , \mem_a[4][8] , \mem_a[4][7] , 
	\mem_a[4][6] , \mem_a[4][5] , \mem_a[4][4] , \mem_a[4][3] , 
	\mem_a[4][2] , \mem_a[4][1] , \mem_a[4][0] , \mem_a[5][31] , 
	\mem_a[5][30] , \mem_a[5][29] , \mem_a[5][28] , \mem_a[5][27] , 
	\mem_a[5][26] , \mem_a[5][25] , \mem_a[5][24] , \mem_a[5][23] , 
	\mem_a[5][22] , \mem_a[5][21] , \mem_a[5][20] , \mem_a[5][19] , 
	\mem_a[5][18] , \mem_a[5][17] , \mem_a[5][16] , \mem_a[5][15] , 
	\mem_a[5][14] , \mem_a[5][13] , \mem_a[5][12] , \mem_a[5][11] , 
	\mem_a[5][10] , \mem_a[5][9] , \mem_a[5][8] , \mem_a[5][7] , 
	\mem_a[5][6] , \mem_a[5][5] , \mem_a[5][4] , \mem_a[5][3] , 
	\mem_a[5][2] , \mem_a[5][1] , \mem_a[5][0] , \mem_a[6][31] , 
	\mem_a[6][30] , \mem_a[6][29] , \mem_a[6][28] , \mem_a[6][27] , 
	\mem_a[6][26] , \mem_a[6][25] , \mem_a[6][24] , \mem_a[6][23] , 
	\mem_a[6][22] , \mem_a[6][21] , \mem_a[6][20] , \mem_a[6][19] , 
	\mem_a[6][18] , \mem_a[6][17] , \mem_a[6][16] , \mem_a[6][15] , 
	\mem_a[6][14] , \mem_a[6][13] , \mem_a[6][12] , \mem_a[6][11] , 
	\mem_a[6][10] , \mem_a[6][9] , \mem_a[6][8] , \mem_a[6][7] , 
	\mem_a[6][6] , \mem_a[6][5] , \mem_a[6][4] , \mem_a[6][3] , 
	\mem_a[6][2] , \mem_a[6][1] , \mem_a[6][0] , \mem_a[7][31] , 
	\mem_a[7][30] , \mem_a[7][29] , \mem_a[7][28] , \mem_a[7][27] , 
	\mem_a[7][26] , \mem_a[7][25] , \mem_a[7][24] , \mem_a[7][23] , 
	\mem_a[7][22] , \mem_a[7][21] , \mem_a[7][20] , \mem_a[7][19] , 
	\mem_a[7][18] , \mem_a[7][17] , \mem_a[7][16] , \mem_a[7][15] , 
	\mem_a[7][14] , \mem_a[7][13] , \mem_a[7][12] , \mem_a[7][11] , 
	\mem_a[7][10] , \mem_a[7][9] , \mem_a[7][8] , \mem_a[7][7] , 
	\mem_a[7][6] , \mem_a[7][5] , \mem_a[7][4] , \mem_a[7][3] , 
	\mem_a[7][2] , \mem_a[7][1] , \mem_a[7][0] , \mem_a[8][31] , 
	\mem_a[8][30] , \mem_a[8][29] , \mem_a[8][28] , \mem_a[8][27] , 
	\mem_a[8][26] , \mem_a[8][25] , \mem_a[8][24] , \mem_a[8][23] , 
	\mem_a[8][22] , \mem_a[8][21] , \mem_a[8][20] , \mem_a[8][19] , 
	\mem_a[8][18] , \mem_a[8][17] , \mem_a[8][16] , \mem_a[8][15] , 
	\mem_a[8][14] , \mem_a[8][13] , \mem_a[8][12] , \mem_a[8][11] , 
	\mem_a[8][10] , \mem_a[8][9] , \mem_a[8][8] , \mem_a[8][7] , 
	\mem_a[8][6] , \mem_a[8][5] , \mem_a[8][4] , \mem_a[8][3] , 
	\mem_a[8][2] , \mem_a[8][1] , \mem_a[8][0] , \mem_a[9][31] , 
	\mem_a[9][30] , \mem_a[9][29] , \mem_a[9][28] , \mem_a[9][27] , 
	\mem_a[9][26] , \mem_a[9][25] , \mem_a[9][24] , \mem_a[9][23] , 
	\mem_a[9][22] , \mem_a[9][21] , \mem_a[9][20] , \mem_a[9][19] , 
	\mem_a[9][18] , \mem_a[9][17] , \mem_a[9][16] , \mem_a[9][15] , 
	\mem_a[9][14] , \mem_a[9][13] , \mem_a[9][12] , \mem_a[9][11] , 
	\mem_a[9][10] , \mem_a[9][9] , \mem_a[9][8] , \mem_a[9][7] , 
	\mem_a[9][6] , \mem_a[9][5] , \mem_a[9][4] , \mem_a[9][3] , 
	\mem_a[9][2] , \mem_a[9][1] , \mem_a[9][0] , \mem_a[10][31] , 
	\mem_a[10][30] , \mem_a[10][29] , \mem_a[10][28] , \mem_a[10][27] , 
	\mem_a[10][26] , \mem_a[10][25] , \mem_a[10][24] , \mem_a[10][23] , 
	\mem_a[10][22] , \mem_a[10][21] , \mem_a[10][20] , \mem_a[10][19] , 
	\mem_a[10][18] , \mem_a[10][17] , \mem_a[10][16] , \mem_a[10][15] , 
	\mem_a[10][14] , \mem_a[10][13] , \mem_a[10][12] , \mem_a[10][11] , 
	\mem_a[10][10] , \mem_a[10][9] , \mem_a[10][8] , \mem_a[10][7] , 
	\mem_a[10][6] , \mem_a[10][5] , \mem_a[10][4] , \mem_a[10][3] , 
	\mem_a[10][2] , \mem_a[10][1] , \mem_a[10][0] , \mem_a[11][31] , 
	\mem_a[11][30] , \mem_a[11][29] , \mem_a[11][28] , \mem_a[11][27] , 
	\mem_a[11][26] , \mem_a[11][25] , \mem_a[11][24] , \mem_a[11][23] , 
	\mem_a[11][22] , \mem_a[11][21] , \mem_a[11][20] , \mem_a[11][19] , 
	\mem_a[11][18] , \mem_a[11][17] , \mem_a[11][16] , \mem_a[11][15] , 
	\mem_a[11][14] , \mem_a[11][13] , \mem_a[11][12] , \mem_a[11][11] , 
	\mem_a[11][10] , \mem_a[11][9] , \mem_a[11][8] , \mem_a[11][7] , 
	\mem_a[11][6] , \mem_a[11][5] , \mem_a[11][4] , \mem_a[11][3] , 
	\mem_a[11][2] , \mem_a[11][1] , \mem_a[11][0] , \mem_a[12][31] , 
	\mem_a[12][30] , \mem_a[12][29] , \mem_a[12][28] , \mem_a[12][27] , 
	\mem_a[12][26] , \mem_a[12][25] , \mem_a[12][24] , \mem_a[12][23] , 
	\mem_a[12][22] , \mem_a[12][21] , \mem_a[12][20] , \mem_a[12][19] , 
	\mem_a[12][18] , \mem_a[12][17] , \mem_a[12][16] , \mem_a[12][15] , 
	\mem_a[12][14] , \mem_a[12][13] , \mem_a[12][12] , \mem_a[12][11] , 
	\mem_a[12][10] , \mem_a[12][9] , \mem_a[12][8] , \mem_a[12][7] , 
	\mem_a[12][6] , \mem_a[12][5] , \mem_a[12][4] , \mem_a[12][3] , 
	\mem_a[12][2] , \mem_a[12][1] , \mem_a[12][0] , \mem_a[13][31] , 
	\mem_a[13][30] , \mem_a[13][29] , \mem_a[13][28] , \mem_a[13][27] , 
	\mem_a[13][26] , \mem_a[13][25] , \mem_a[13][24] , \mem_a[13][23] , 
	\mem_a[13][22] , \mem_a[13][21] , \mem_a[13][20] , \mem_a[13][19] , 
	\mem_a[13][18] , \mem_a[13][17] , \mem_a[13][16] , \mem_a[13][15] , 
	\mem_a[13][14] , \mem_a[13][13] , \mem_a[13][12] , \mem_a[13][11] , 
	\mem_a[13][10] , \mem_a[13][9] , \mem_a[13][8] , \mem_a[13][7] , 
	\mem_a[13][6] , \mem_a[13][5] , \mem_a[13][4] , \mem_a[13][3] , 
	\mem_a[13][2] , \mem_a[13][1] , \mem_a[13][0] , \mem_a[14][31] , 
	\mem_a[14][30] , \mem_a[14][29] , \mem_a[14][28] , \mem_a[14][27] , 
	\mem_a[14][26] , \mem_a[14][25] , \mem_a[14][24] , \mem_a[14][23] , 
	\mem_a[14][22] , \mem_a[14][21] , \mem_a[14][20] , \mem_a[14][19] , 
	\mem_a[14][18] , \mem_a[14][17] , \mem_a[14][16] , \mem_a[14][15] , 
	\mem_a[14][14] , \mem_a[14][13] , \mem_a[14][12] , \mem_a[14][11] , 
	\mem_a[14][10] , \mem_a[14][9] , \mem_a[14][8] , \mem_a[14][7] , 
	\mem_a[14][6] , \mem_a[14][5] , \mem_a[14][4] , \mem_a[14][3] , 
	\mem_a[14][2] , \mem_a[14][1] , \mem_a[14][0] , \mem_a[15][31] , 
	\mem_a[15][30] , \mem_a[15][29] , \mem_a[15][28] , \mem_a[15][27] , 
	\mem_a[15][26] , \mem_a[15][25] , \mem_a[15][24] , \mem_a[15][23] , 
	\mem_a[15][22] , \mem_a[15][21] , \mem_a[15][20] , \mem_a[15][19] , 
	\mem_a[15][18] , \mem_a[15][17] , \mem_a[15][16] , \mem_a[15][15] , 
	\mem_a[15][14] , \mem_a[15][13] , \mem_a[15][12] , \mem_a[15][11] , 
	\mem_a[15][10] , \mem_a[15][9] , \mem_a[15][8] , \mem_a[15][7] , 
	\mem_a[15][6] , \mem_a[15][5] , \mem_a[15][4] , \mem_a[15][3] , 
	\mem_a[15][2] , \mem_a[15][1] , \mem_a[15][0] , \mem_a[16][31] , 
	\mem_a[16][30] , \mem_a[16][29] , \mem_a[16][28] , \mem_a[16][27] , 
	\mem_a[16][26] , \mem_a[16][25] , \mem_a[16][24] , \mem_a[16][23] , 
	\mem_a[16][22] , \mem_a[16][21] , \mem_a[16][20] , \mem_a[16][19] , 
	\mem_a[16][18] , \mem_a[16][17] , \mem_a[16][16] , \mem_a[16][15] , 
	\mem_a[16][14] , \mem_a[16][13] , \mem_a[16][12] , \mem_a[16][11] , 
	\mem_a[16][10] , \mem_a[16][9] , \mem_a[16][8] , \mem_a[16][7] , 
	\mem_a[16][6] , \mem_a[16][5] , \mem_a[16][4] , \mem_a[16][3] , 
	\mem_a[16][2] , \mem_a[16][1] , \mem_a[16][0] , \mem_a[17][31] , 
	\mem_a[17][30] , \mem_a[17][29] , \mem_a[17][28] , \mem_a[17][27] , 
	\mem_a[17][26] , \mem_a[17][25] , \mem_a[17][24] , \mem_a[17][23] , 
	\mem_a[17][22] , \mem_a[17][21] , \mem_a[17][20] , \mem_a[17][19] , 
	\mem_a[17][18] , \mem_a[17][17] , \mem_a[17][16] , \mem_a[17][15] , 
	\mem_a[17][14] , \mem_a[17][13] , \mem_a[17][12] , \mem_a[17][11] , 
	\mem_a[17][10] , \mem_a[17][9] , \mem_a[17][8] , \mem_a[17][7] , 
	\mem_a[17][6] , \mem_a[17][5] , \mem_a[17][4] , \mem_a[17][3] , 
	\mem_a[17][2] , \mem_a[17][1] , \mem_a[17][0] , \mem_a[18][31] , 
	\mem_a[18][30] , \mem_a[18][29] , \mem_a[18][28] , \mem_a[18][27] , 
	\mem_a[18][26] , \mem_a[18][25] , \mem_a[18][24] , \mem_a[18][23] , 
	\mem_a[18][22] , \mem_a[18][21] , \mem_a[18][20] , \mem_a[18][19] , 
	\mem_a[18][18] , \mem_a[18][17] , \mem_a[18][16] , \mem_a[18][15] , 
	\mem_a[18][14] , \mem_a[18][13] , \mem_a[18][12] , \mem_a[18][11] , 
	\mem_a[18][10] , \mem_a[18][9] , \mem_a[18][8] , \mem_a[18][7] , 
	\mem_a[18][6] , \mem_a[18][5] , \mem_a[18][4] , \mem_a[18][3] , 
	\mem_a[18][2] , \mem_a[18][1] , \mem_a[18][0] , \mem_a[19][31] , 
	\mem_a[19][30] , \mem_a[19][29] , \mem_a[19][28] , \mem_a[19][27] , 
	\mem_a[19][26] , \mem_a[19][25] , \mem_a[19][24] , \mem_a[19][23] , 
	\mem_a[19][22] , \mem_a[19][21] , \mem_a[19][20] , \mem_a[19][19] , 
	\mem_a[19][18] , \mem_a[19][17] , \mem_a[19][16] , \mem_a[19][15] , 
	\mem_a[19][14] , \mem_a[19][13] , \mem_a[19][12] , \mem_a[19][11] , 
	\mem_a[19][10] , \mem_a[19][9] , \mem_a[19][8] , \mem_a[19][7] , 
	\mem_a[19][6] , \mem_a[19][5] , \mem_a[19][4] , \mem_a[19][3] , 
	\mem_a[19][2] , \mem_a[19][1] , \mem_a[19][0] , \mem_a[20][31] , 
	\mem_a[20][30] , \mem_a[20][29] , \mem_a[20][28] , \mem_a[20][27] , 
	\mem_a[20][26] , \mem_a[20][25] , \mem_a[20][24] , \mem_a[20][23] , 
	\mem_a[20][22] , \mem_a[20][21] , \mem_a[20][20] , \mem_a[20][19] , 
	\mem_a[20][18] , \mem_a[20][17] , \mem_a[20][16] , \mem_a[20][15] , 
	\mem_a[20][14] , \mem_a[20][13] , \mem_a[20][12] , \mem_a[20][11] , 
	\mem_a[20][10] , \mem_a[20][9] , \mem_a[20][8] , \mem_a[20][7] , 
	\mem_a[20][6] , \mem_a[20][5] , \mem_a[20][4] , \mem_a[20][3] , 
	\mem_a[20][2] , \mem_a[20][1] , \mem_a[20][0] , \mem_a[21][31] , 
	\mem_a[21][30] , \mem_a[21][29] , \mem_a[21][28] , \mem_a[21][27] , 
	\mem_a[21][26] , \mem_a[21][25] , \mem_a[21][24] , \mem_a[21][23] , 
	\mem_a[21][22] , \mem_a[21][21] , \mem_a[21][20] , \mem_a[21][19] , 
	\mem_a[21][18] , \mem_a[21][17] , \mem_a[21][16] , \mem_a[21][15] , 
	\mem_a[21][14] , \mem_a[21][13] , \mem_a[21][12] , \mem_a[21][11] , 
	\mem_a[21][10] , \mem_a[21][9] , \mem_a[21][8] , \mem_a[21][7] , 
	\mem_a[21][6] , \mem_a[21][5] , \mem_a[21][4] , \mem_a[21][3] , 
	\mem_a[21][2] , \mem_a[21][1] , \mem_a[21][0] , \mem_a[22][31] , 
	\mem_a[22][30] , \mem_a[22][29] , \mem_a[22][28] , \mem_a[22][27] , 
	\mem_a[22][26] , \mem_a[22][25] , \mem_a[22][24] , \mem_a[22][23] , 
	\mem_a[22][22] , \mem_a[22][21] , \mem_a[22][20] , \mem_a[22][19] , 
	\mem_a[22][18] , \mem_a[22][17] , \mem_a[22][16] , \mem_a[22][15] , 
	\mem_a[22][14] , \mem_a[22][13] , \mem_a[22][12] , \mem_a[22][11] , 
	\mem_a[22][10] , \mem_a[22][9] , \mem_a[22][8] , \mem_a[22][7] , 
	\mem_a[22][6] , \mem_a[22][5] , \mem_a[22][4] , \mem_a[22][3] , 
	\mem_a[22][2] , \mem_a[22][1] , \mem_a[22][0] , \mem_a[23][31] , 
	\mem_a[23][30] , \mem_a[23][29] , \mem_a[23][28] , \mem_a[23][27] , 
	\mem_a[23][26] , \mem_a[23][25] , \mem_a[23][24] , \mem_a[23][23] , 
	\mem_a[23][22] , \mem_a[23][21] , \mem_a[23][20] , \mem_a[23][19] , 
	\mem_a[23][18] , \mem_a[23][17] , \mem_a[23][16] , \mem_a[23][15] , 
	\mem_a[23][14] , \mem_a[23][13] , \mem_a[23][12] , \mem_a[23][11] , 
	\mem_a[23][10] , \mem_a[23][9] , \mem_a[23][8] , \mem_a[23][7] , 
	\mem_a[23][6] , \mem_a[23][5] , \mem_a[23][4] , \mem_a[23][3] , 
	\mem_a[23][2] , \mem_a[23][1] , \mem_a[23][0] , \mem_a[24][31] , 
	\mem_a[24][30] , \mem_a[24][29] , \mem_a[24][28] , \mem_a[24][27] , 
	\mem_a[24][26] , \mem_a[24][25] , \mem_a[24][24] , \mem_a[24][23] , 
	\mem_a[24][22] , \mem_a[24][21] , \mem_a[24][20] , \mem_a[24][19] , 
	\mem_a[24][18] , \mem_a[24][17] , \mem_a[24][16] , \mem_a[24][15] , 
	\mem_a[24][14] , \mem_a[24][13] , \mem_a[24][12] , \mem_a[24][11] , 
	\mem_a[24][10] , \mem_a[24][9] , \mem_a[24][8] , \mem_a[24][7] , 
	\mem_a[24][6] , \mem_a[24][5] , \mem_a[24][4] , \mem_a[24][3] , 
	\mem_a[24][2] , \mem_a[24][1] , \mem_a[24][0] , \mem_a[25][31] , 
	\mem_a[25][30] , \mem_a[25][29] , \mem_a[25][28] , \mem_a[25][27] , 
	\mem_a[25][26] , \mem_a[25][25] , \mem_a[25][24] , \mem_a[25][23] , 
	\mem_a[25][22] , \mem_a[25][21] , \mem_a[25][20] , \mem_a[25][19] , 
	\mem_a[25][18] , \mem_a[25][17] , \mem_a[25][16] , \mem_a[25][15] , 
	\mem_a[25][14] , \mem_a[25][13] , \mem_a[25][12] , \mem_a[25][11] , 
	\mem_a[25][10] , \mem_a[25][9] , \mem_a[25][8] , \mem_a[25][7] , 
	\mem_a[25][6] , \mem_a[25][5] , \mem_a[25][4] , \mem_a[25][3] , 
	\mem_a[25][2] , \mem_a[25][1] , \mem_a[25][0] , \mem_a[26][31] , 
	\mem_a[26][30] , \mem_a[26][29] , \mem_a[26][28] , \mem_a[26][27] , 
	\mem_a[26][26] , \mem_a[26][25] , \mem_a[26][24] , \mem_a[26][23] , 
	\mem_a[26][22] , \mem_a[26][21] , \mem_a[26][20] , \mem_a[26][19] , 
	\mem_a[26][18] , \mem_a[26][17] , \mem_a[26][16] , \mem_a[26][15] , 
	\mem_a[26][14] , \mem_a[26][13] , \mem_a[26][12] , \mem_a[26][11] , 
	\mem_a[26][10] , \mem_a[26][9] , \mem_a[26][8] , \mem_a[26][7] , 
	\mem_a[26][6] , \mem_a[26][5] , \mem_a[26][4] , \mem_a[26][3] , 
	\mem_a[26][2] , \mem_a[26][1] , \mem_a[26][0] , \mem_a[27][31] , 
	\mem_a[27][30] , \mem_a[27][29] , \mem_a[27][28] , \mem_a[27][27] , 
	\mem_a[27][26] , \mem_a[27][25] , \mem_a[27][24] , \mem_a[27][23] , 
	\mem_a[27][22] , \mem_a[27][21] , \mem_a[27][20] , \mem_a[27][19] , 
	\mem_a[27][18] , \mem_a[27][17] , \mem_a[27][16] , \mem_a[27][15] , 
	\mem_a[27][14] , \mem_a[27][13] , \mem_a[27][12] , \mem_a[27][11] , 
	\mem_a[27][10] , \mem_a[27][9] , \mem_a[27][8] , \mem_a[27][7] , 
	\mem_a[27][6] , \mem_a[27][5] , \mem_a[27][4] , \mem_a[27][3] , 
	\mem_a[27][2] , \mem_a[27][1] , \mem_a[27][0] , \mem_a[28][31] , 
	\mem_a[28][30] , \mem_a[28][29] , \mem_a[28][28] , \mem_a[28][27] , 
	\mem_a[28][26] , \mem_a[28][25] , \mem_a[28][24] , \mem_a[28][23] , 
	\mem_a[28][22] , \mem_a[28][21] , \mem_a[28][20] , \mem_a[28][19] , 
	\mem_a[28][18] , \mem_a[28][17] , \mem_a[28][16] , \mem_a[28][15] , 
	\mem_a[28][14] , \mem_a[28][13] , \mem_a[28][12] , \mem_a[28][11] , 
	\mem_a[28][10] , \mem_a[28][9] , \mem_a[28][8] , \mem_a[28][7] , 
	\mem_a[28][6] , \mem_a[28][5] , \mem_a[28][4] , \mem_a[28][3] , 
	\mem_a[28][2] , \mem_a[28][1] , \mem_a[28][0] , \mem_a[29][31] , 
	\mem_a[29][30] , \mem_a[29][29] , \mem_a[29][28] , \mem_a[29][27] , 
	\mem_a[29][26] , \mem_a[29][25] , \mem_a[29][24] , \mem_a[29][23] , 
	\mem_a[29][22] , \mem_a[29][21] , \mem_a[29][20] , \mem_a[29][19] , 
	\mem_a[29][18] , \mem_a[29][17] , \mem_a[29][16] , \mem_a[29][15] , 
	\mem_a[29][14] , \mem_a[29][13] , \mem_a[29][12] , \mem_a[29][11] , 
	\mem_a[29][10] , \mem_a[29][9] , \mem_a[29][8] , \mem_a[29][7] , 
	\mem_a[29][6] , \mem_a[29][5] , \mem_a[29][4] , \mem_a[29][3] , 
	\mem_a[29][2] , \mem_a[29][1] , \mem_a[29][0] , \mem_a[30][31] , 
	\mem_a[30][30] , \mem_a[30][29] , \mem_a[30][28] , \mem_a[30][27] , 
	\mem_a[30][26] , \mem_a[30][25] , \mem_a[30][24] , \mem_a[30][23] , 
	\mem_a[30][22] , \mem_a[30][21] , \mem_a[30][20] , \mem_a[30][19] , 
	\mem_a[30][18] , \mem_a[30][17] , \mem_a[30][16] , \mem_a[30][15] , 
	\mem_a[30][14] , \mem_a[30][13] , \mem_a[30][12] , \mem_a[30][11] , 
	\mem_a[30][10] , \mem_a[30][9] , \mem_a[30][8] , \mem_a[30][7] , 
	\mem_a[30][6] , \mem_a[30][5] , \mem_a[30][4] , \mem_a[30][3] , 
	\mem_a[30][2] , \mem_a[30][1] , \mem_a[30][0] , \mem_a[31][31] , 
	\mem_a[31][30] , \mem_a[31][29] , \mem_a[31][28] , \mem_a[31][27] , 
	\mem_a[31][26] , \mem_a[31][25] , \mem_a[31][24] , \mem_a[31][23] , 
	\mem_a[31][22] , \mem_a[31][21] , \mem_a[31][20] , \mem_a[31][19] , 
	\mem_a[31][18] , \mem_a[31][17] , \mem_a[31][16] , \mem_a[31][15] , 
	\mem_a[31][14] , \mem_a[31][13] , \mem_a[31][12] , \mem_a[31][11] , 
	\mem_a[31][10] , \mem_a[31][9] , \mem_a[31][8] , \mem_a[31][7] , 
	\mem_a[31][6] , \mem_a[31][5] , \mem_a[31][4] , \mem_a[31][3] , 
	\mem_a[31][2] , \mem_a[31][1] , \mem_a[31][0] } ), clk, rst_n, addr, 
	cmnd_op, cmnd_addr, wr_stb, wr_dat, .rst_dat( {\rst_dat[0][31] , 
	\rst_dat[0][30] , \rst_dat[0][29] , \rst_dat[0][28] , 
	\rst_dat[0][27] , \rst_dat[0][26] , \rst_dat[0][25] , 
	\rst_dat[0][24] , \rst_dat[0][23] , \rst_dat[0][22] , 
	\rst_dat[0][21] , \rst_dat[0][20] , \rst_dat[0][19] , 
	\rst_dat[0][18] , \rst_dat[0][17] , \rst_dat[0][16] , 
	\rst_dat[0][15] , \rst_dat[0][14] , \rst_dat[0][13] , 
	\rst_dat[0][12] , \rst_dat[0][11] , \rst_dat[0][10] , 
	\rst_dat[0][9] , \rst_dat[0][8] , \rst_dat[0][7] , \rst_dat[0][6] , 
	\rst_dat[0][5] , \rst_dat[0][4] , \rst_dat[0][3] , \rst_dat[0][2] , 
	\rst_dat[0][1] , \rst_dat[0][0] , \rst_dat[1][31] , \rst_dat[1][30] , 
	\rst_dat[1][29] , \rst_dat[1][28] , \rst_dat[1][27] , 
	\rst_dat[1][26] , \rst_dat[1][25] , \rst_dat[1][24] , 
	\rst_dat[1][23] , \rst_dat[1][22] , \rst_dat[1][21] , 
	\rst_dat[1][20] , \rst_dat[1][19] , \rst_dat[1][18] , 
	\rst_dat[1][17] , \rst_dat[1][16] , \rst_dat[1][15] , 
	\rst_dat[1][14] , \rst_dat[1][13] , \rst_dat[1][12] , 
	\rst_dat[1][11] , \rst_dat[1][10] , \rst_dat[1][9] , \rst_dat[1][8] , 
	\rst_dat[1][7] , \rst_dat[1][6] , \rst_dat[1][5] , \rst_dat[1][4] , 
	\rst_dat[1][3] , \rst_dat[1][2] , \rst_dat[1][1] , \rst_dat[1][0] , 
	\rst_dat[2][31] , \rst_dat[2][30] , \rst_dat[2][29] , 
	\rst_dat[2][28] , \rst_dat[2][27] , \rst_dat[2][26] , 
	\rst_dat[2][25] , \rst_dat[2][24] , \rst_dat[2][23] , 
	\rst_dat[2][22] , \rst_dat[2][21] , \rst_dat[2][20] , 
	\rst_dat[2][19] , \rst_dat[2][18] , \rst_dat[2][17] , 
	\rst_dat[2][16] , \rst_dat[2][15] , \rst_dat[2][14] , 
	\rst_dat[2][13] , \rst_dat[2][12] , \rst_dat[2][11] , 
	\rst_dat[2][10] , \rst_dat[2][9] , \rst_dat[2][8] , \rst_dat[2][7] , 
	\rst_dat[2][6] , \rst_dat[2][5] , \rst_dat[2][4] , \rst_dat[2][3] , 
	\rst_dat[2][2] , \rst_dat[2][1] , \rst_dat[2][0] , \rst_dat[3][31] , 
	\rst_dat[3][30] , \rst_dat[3][29] , \rst_dat[3][28] , 
	\rst_dat[3][27] , \rst_dat[3][26] , \rst_dat[3][25] , 
	\rst_dat[3][24] , \rst_dat[3][23] , \rst_dat[3][22] , 
	\rst_dat[3][21] , \rst_dat[3][20] , \rst_dat[3][19] , 
	\rst_dat[3][18] , \rst_dat[3][17] , \rst_dat[3][16] , 
	\rst_dat[3][15] , \rst_dat[3][14] , \rst_dat[3][13] , 
	\rst_dat[3][12] , \rst_dat[3][11] , \rst_dat[3][10] , 
	\rst_dat[3][9] , \rst_dat[3][8] , \rst_dat[3][7] , \rst_dat[3][6] , 
	\rst_dat[3][5] , \rst_dat[3][4] , \rst_dat[3][3] , \rst_dat[3][2] , 
	\rst_dat[3][1] , \rst_dat[3][0] , \rst_dat[4][31] , \rst_dat[4][30] , 
	\rst_dat[4][29] , \rst_dat[4][28] , \rst_dat[4][27] , 
	\rst_dat[4][26] , \rst_dat[4][25] , \rst_dat[4][24] , 
	\rst_dat[4][23] , \rst_dat[4][22] , \rst_dat[4][21] , 
	\rst_dat[4][20] , \rst_dat[4][19] , \rst_dat[4][18] , 
	\rst_dat[4][17] , \rst_dat[4][16] , \rst_dat[4][15] , 
	\rst_dat[4][14] , \rst_dat[4][13] , \rst_dat[4][12] , 
	\rst_dat[4][11] , \rst_dat[4][10] , \rst_dat[4][9] , \rst_dat[4][8] , 
	\rst_dat[4][7] , \rst_dat[4][6] , \rst_dat[4][5] , \rst_dat[4][4] , 
	\rst_dat[4][3] , \rst_dat[4][2] , \rst_dat[4][1] , \rst_dat[4][0] , 
	\rst_dat[5][31] , \rst_dat[5][30] , \rst_dat[5][29] , 
	\rst_dat[5][28] , \rst_dat[5][27] , \rst_dat[5][26] , 
	\rst_dat[5][25] , \rst_dat[5][24] , \rst_dat[5][23] , 
	\rst_dat[5][22] , \rst_dat[5][21] , \rst_dat[5][20] , 
	\rst_dat[5][19] , \rst_dat[5][18] , \rst_dat[5][17] , 
	\rst_dat[5][16] , \rst_dat[5][15] , \rst_dat[5][14] , 
	\rst_dat[5][13] , \rst_dat[5][12] , \rst_dat[5][11] , 
	\rst_dat[5][10] , \rst_dat[5][9] , \rst_dat[5][8] , \rst_dat[5][7] , 
	\rst_dat[5][6] , \rst_dat[5][5] , \rst_dat[5][4] , \rst_dat[5][3] , 
	\rst_dat[5][2] , \rst_dat[5][1] , \rst_dat[5][0] , \rst_dat[6][31] , 
	\rst_dat[6][30] , \rst_dat[6][29] , \rst_dat[6][28] , 
	\rst_dat[6][27] , \rst_dat[6][26] , \rst_dat[6][25] , 
	\rst_dat[6][24] , \rst_dat[6][23] , \rst_dat[6][22] , 
	\rst_dat[6][21] , \rst_dat[6][20] , \rst_dat[6][19] , 
	\rst_dat[6][18] , \rst_dat[6][17] , \rst_dat[6][16] , 
	\rst_dat[6][15] , \rst_dat[6][14] , \rst_dat[6][13] , 
	\rst_dat[6][12] , \rst_dat[6][11] , \rst_dat[6][10] , 
	\rst_dat[6][9] , \rst_dat[6][8] , \rst_dat[6][7] , \rst_dat[6][6] , 
	\rst_dat[6][5] , \rst_dat[6][4] , \rst_dat[6][3] , \rst_dat[6][2] , 
	\rst_dat[6][1] , \rst_dat[6][0] , \rst_dat[7][31] , \rst_dat[7][30] , 
	\rst_dat[7][29] , \rst_dat[7][28] , \rst_dat[7][27] , 
	\rst_dat[7][26] , \rst_dat[7][25] , \rst_dat[7][24] , 
	\rst_dat[7][23] , \rst_dat[7][22] , \rst_dat[7][21] , 
	\rst_dat[7][20] , \rst_dat[7][19] , \rst_dat[7][18] , 
	\rst_dat[7][17] , \rst_dat[7][16] , \rst_dat[7][15] , 
	\rst_dat[7][14] , \rst_dat[7][13] , \rst_dat[7][12] , 
	\rst_dat[7][11] , \rst_dat[7][10] , \rst_dat[7][9] , \rst_dat[7][8] , 
	\rst_dat[7][7] , \rst_dat[7][6] , \rst_dat[7][5] , \rst_dat[7][4] , 
	\rst_dat[7][3] , \rst_dat[7][2] , \rst_dat[7][1] , \rst_dat[7][0] , 
	\rst_dat[8][31] , \rst_dat[8][30] , \rst_dat[8][29] , 
	\rst_dat[8][28] , \rst_dat[8][27] , \rst_dat[8][26] , 
	\rst_dat[8][25] , \rst_dat[8][24] , \rst_dat[8][23] , 
	\rst_dat[8][22] , \rst_dat[8][21] , \rst_dat[8][20] , 
	\rst_dat[8][19] , \rst_dat[8][18] , \rst_dat[8][17] , 
	\rst_dat[8][16] , \rst_dat[8][15] , \rst_dat[8][14] , 
	\rst_dat[8][13] , \rst_dat[8][12] , \rst_dat[8][11] , 
	\rst_dat[8][10] , \rst_dat[8][9] , \rst_dat[8][8] , \rst_dat[8][7] , 
	\rst_dat[8][6] , \rst_dat[8][5] , \rst_dat[8][4] , \rst_dat[8][3] , 
	\rst_dat[8][2] , \rst_dat[8][1] , \rst_dat[8][0] , \rst_dat[9][31] , 
	\rst_dat[9][30] , \rst_dat[9][29] , \rst_dat[9][28] , 
	\rst_dat[9][27] , \rst_dat[9][26] , \rst_dat[9][25] , 
	\rst_dat[9][24] , \rst_dat[9][23] , \rst_dat[9][22] , 
	\rst_dat[9][21] , \rst_dat[9][20] , \rst_dat[9][19] , 
	\rst_dat[9][18] , \rst_dat[9][17] , \rst_dat[9][16] , 
	\rst_dat[9][15] , \rst_dat[9][14] , \rst_dat[9][13] , 
	\rst_dat[9][12] , \rst_dat[9][11] , \rst_dat[9][10] , 
	\rst_dat[9][9] , \rst_dat[9][8] , \rst_dat[9][7] , \rst_dat[9][6] , 
	\rst_dat[9][5] , \rst_dat[9][4] , \rst_dat[9][3] , \rst_dat[9][2] , 
	\rst_dat[9][1] , \rst_dat[9][0] , \rst_dat[10][31] , 
	\rst_dat[10][30] , \rst_dat[10][29] , \rst_dat[10][28] , 
	\rst_dat[10][27] , \rst_dat[10][26] , \rst_dat[10][25] , 
	\rst_dat[10][24] , \rst_dat[10][23] , \rst_dat[10][22] , 
	\rst_dat[10][21] , \rst_dat[10][20] , \rst_dat[10][19] , 
	\rst_dat[10][18] , \rst_dat[10][17] , \rst_dat[10][16] , 
	\rst_dat[10][15] , \rst_dat[10][14] , \rst_dat[10][13] , 
	\rst_dat[10][12] , \rst_dat[10][11] , \rst_dat[10][10] , 
	\rst_dat[10][9] , \rst_dat[10][8] , \rst_dat[10][7] , 
	\rst_dat[10][6] , \rst_dat[10][5] , \rst_dat[10][4] , 
	\rst_dat[10][3] , \rst_dat[10][2] , \rst_dat[10][1] , 
	\rst_dat[10][0] , \rst_dat[11][31] , \rst_dat[11][30] , 
	\rst_dat[11][29] , \rst_dat[11][28] , \rst_dat[11][27] , 
	\rst_dat[11][26] , \rst_dat[11][25] , \rst_dat[11][24] , 
	\rst_dat[11][23] , \rst_dat[11][22] , \rst_dat[11][21] , 
	\rst_dat[11][20] , \rst_dat[11][19] , \rst_dat[11][18] , 
	\rst_dat[11][17] , \rst_dat[11][16] , \rst_dat[11][15] , 
	\rst_dat[11][14] , \rst_dat[11][13] , \rst_dat[11][12] , 
	\rst_dat[11][11] , \rst_dat[11][10] , \rst_dat[11][9] , 
	\rst_dat[11][8] , \rst_dat[11][7] , \rst_dat[11][6] , 
	\rst_dat[11][5] , \rst_dat[11][4] , \rst_dat[11][3] , 
	\rst_dat[11][2] , \rst_dat[11][1] , \rst_dat[11][0] , 
	\rst_dat[12][31] , \rst_dat[12][30] , \rst_dat[12][29] , 
	\rst_dat[12][28] , \rst_dat[12][27] , \rst_dat[12][26] , 
	\rst_dat[12][25] , \rst_dat[12][24] , \rst_dat[12][23] , 
	\rst_dat[12][22] , \rst_dat[12][21] , \rst_dat[12][20] , 
	\rst_dat[12][19] , \rst_dat[12][18] , \rst_dat[12][17] , 
	\rst_dat[12][16] , \rst_dat[12][15] , \rst_dat[12][14] , 
	\rst_dat[12][13] , \rst_dat[12][12] , \rst_dat[12][11] , 
	\rst_dat[12][10] , \rst_dat[12][9] , \rst_dat[12][8] , 
	\rst_dat[12][7] , \rst_dat[12][6] , \rst_dat[12][5] , 
	\rst_dat[12][4] , \rst_dat[12][3] , \rst_dat[12][2] , 
	\rst_dat[12][1] , \rst_dat[12][0] , \rst_dat[13][31] , 
	\rst_dat[13][30] , \rst_dat[13][29] , \rst_dat[13][28] , 
	\rst_dat[13][27] , \rst_dat[13][26] , \rst_dat[13][25] , 
	\rst_dat[13][24] , \rst_dat[13][23] , \rst_dat[13][22] , 
	\rst_dat[13][21] , \rst_dat[13][20] , \rst_dat[13][19] , 
	\rst_dat[13][18] , \rst_dat[13][17] , \rst_dat[13][16] , 
	\rst_dat[13][15] , \rst_dat[13][14] , \rst_dat[13][13] , 
	\rst_dat[13][12] , \rst_dat[13][11] , \rst_dat[13][10] , 
	\rst_dat[13][9] , \rst_dat[13][8] , \rst_dat[13][7] , 
	\rst_dat[13][6] , \rst_dat[13][5] , \rst_dat[13][4] , 
	\rst_dat[13][3] , \rst_dat[13][2] , \rst_dat[13][1] , 
	\rst_dat[13][0] , \rst_dat[14][31] , \rst_dat[14][30] , 
	\rst_dat[14][29] , \rst_dat[14][28] , \rst_dat[14][27] , 
	\rst_dat[14][26] , \rst_dat[14][25] , \rst_dat[14][24] , 
	\rst_dat[14][23] , \rst_dat[14][22] , \rst_dat[14][21] , 
	\rst_dat[14][20] , \rst_dat[14][19] , \rst_dat[14][18] , 
	\rst_dat[14][17] , \rst_dat[14][16] , \rst_dat[14][15] , 
	\rst_dat[14][14] , \rst_dat[14][13] , \rst_dat[14][12] , 
	\rst_dat[14][11] , \rst_dat[14][10] , \rst_dat[14][9] , 
	\rst_dat[14][8] , \rst_dat[14][7] , \rst_dat[14][6] , 
	\rst_dat[14][5] , \rst_dat[14][4] , \rst_dat[14][3] , 
	\rst_dat[14][2] , \rst_dat[14][1] , \rst_dat[14][0] , 
	\rst_dat[15][31] , \rst_dat[15][30] , \rst_dat[15][29] , 
	\rst_dat[15][28] , \rst_dat[15][27] , \rst_dat[15][26] , 
	\rst_dat[15][25] , \rst_dat[15][24] , \rst_dat[15][23] , 
	\rst_dat[15][22] , \rst_dat[15][21] , \rst_dat[15][20] , 
	\rst_dat[15][19] , \rst_dat[15][18] , \rst_dat[15][17] , 
	\rst_dat[15][16] , \rst_dat[15][15] , \rst_dat[15][14] , 
	\rst_dat[15][13] , \rst_dat[15][12] , \rst_dat[15][11] , 
	\rst_dat[15][10] , \rst_dat[15][9] , \rst_dat[15][8] , 
	\rst_dat[15][7] , \rst_dat[15][6] , \rst_dat[15][5] , 
	\rst_dat[15][4] , \rst_dat[15][3] , \rst_dat[15][2] , 
	\rst_dat[15][1] , \rst_dat[15][0] , \rst_dat[16][31] , 
	\rst_dat[16][30] , \rst_dat[16][29] , \rst_dat[16][28] , 
	\rst_dat[16][27] , \rst_dat[16][26] , \rst_dat[16][25] , 
	\rst_dat[16][24] , \rst_dat[16][23] , \rst_dat[16][22] , 
	\rst_dat[16][21] , \rst_dat[16][20] , \rst_dat[16][19] , 
	\rst_dat[16][18] , \rst_dat[16][17] , \rst_dat[16][16] , 
	\rst_dat[16][15] , \rst_dat[16][14] , \rst_dat[16][13] , 
	\rst_dat[16][12] , \rst_dat[16][11] , \rst_dat[16][10] , 
	\rst_dat[16][9] , \rst_dat[16][8] , \rst_dat[16][7] , 
	\rst_dat[16][6] , \rst_dat[16][5] , \rst_dat[16][4] , 
	\rst_dat[16][3] , \rst_dat[16][2] , \rst_dat[16][1] , 
	\rst_dat[16][0] , \rst_dat[17][31] , \rst_dat[17][30] , 
	\rst_dat[17][29] , \rst_dat[17][28] , \rst_dat[17][27] , 
	\rst_dat[17][26] , \rst_dat[17][25] , \rst_dat[17][24] , 
	\rst_dat[17][23] , \rst_dat[17][22] , \rst_dat[17][21] , 
	\rst_dat[17][20] , \rst_dat[17][19] , \rst_dat[17][18] , 
	\rst_dat[17][17] , \rst_dat[17][16] , \rst_dat[17][15] , 
	\rst_dat[17][14] , \rst_dat[17][13] , \rst_dat[17][12] , 
	\rst_dat[17][11] , \rst_dat[17][10] , \rst_dat[17][9] , 
	\rst_dat[17][8] , \rst_dat[17][7] , \rst_dat[17][6] , 
	\rst_dat[17][5] , \rst_dat[17][4] , \rst_dat[17][3] , 
	\rst_dat[17][2] , \rst_dat[17][1] , \rst_dat[17][0] , 
	\rst_dat[18][31] , \rst_dat[18][30] , \rst_dat[18][29] , 
	\rst_dat[18][28] , \rst_dat[18][27] , \rst_dat[18][26] , 
	\rst_dat[18][25] , \rst_dat[18][24] , \rst_dat[18][23] , 
	\rst_dat[18][22] , \rst_dat[18][21] , \rst_dat[18][20] , 
	\rst_dat[18][19] , \rst_dat[18][18] , \rst_dat[18][17] , 
	\rst_dat[18][16] , \rst_dat[18][15] , \rst_dat[18][14] , 
	\rst_dat[18][13] , \rst_dat[18][12] , \rst_dat[18][11] , 
	\rst_dat[18][10] , \rst_dat[18][9] , \rst_dat[18][8] , 
	\rst_dat[18][7] , \rst_dat[18][6] , \rst_dat[18][5] , 
	\rst_dat[18][4] , \rst_dat[18][3] , \rst_dat[18][2] , 
	\rst_dat[18][1] , \rst_dat[18][0] , \rst_dat[19][31] , 
	\rst_dat[19][30] , \rst_dat[19][29] , \rst_dat[19][28] , 
	\rst_dat[19][27] , \rst_dat[19][26] , \rst_dat[19][25] , 
	\rst_dat[19][24] , \rst_dat[19][23] , \rst_dat[19][22] , 
	\rst_dat[19][21] , \rst_dat[19][20] , \rst_dat[19][19] , 
	\rst_dat[19][18] , \rst_dat[19][17] , \rst_dat[19][16] , 
	\rst_dat[19][15] , \rst_dat[19][14] , \rst_dat[19][13] , 
	\rst_dat[19][12] , \rst_dat[19][11] , \rst_dat[19][10] , 
	\rst_dat[19][9] , \rst_dat[19][8] , \rst_dat[19][7] , 
	\rst_dat[19][6] , \rst_dat[19][5] , \rst_dat[19][4] , 
	\rst_dat[19][3] , \rst_dat[19][2] , \rst_dat[19][1] , 
	\rst_dat[19][0] , \rst_dat[20][31] , \rst_dat[20][30] , 
	\rst_dat[20][29] , \rst_dat[20][28] , \rst_dat[20][27] , 
	\rst_dat[20][26] , \rst_dat[20][25] , \rst_dat[20][24] , 
	\rst_dat[20][23] , \rst_dat[20][22] , \rst_dat[20][21] , 
	\rst_dat[20][20] , \rst_dat[20][19] , \rst_dat[20][18] , 
	\rst_dat[20][17] , \rst_dat[20][16] , \rst_dat[20][15] , 
	\rst_dat[20][14] , \rst_dat[20][13] , \rst_dat[20][12] , 
	\rst_dat[20][11] , \rst_dat[20][10] , \rst_dat[20][9] , 
	\rst_dat[20][8] , \rst_dat[20][7] , \rst_dat[20][6] , 
	\rst_dat[20][5] , \rst_dat[20][4] , \rst_dat[20][3] , 
	\rst_dat[20][2] , \rst_dat[20][1] , \rst_dat[20][0] , 
	\rst_dat[21][31] , \rst_dat[21][30] , \rst_dat[21][29] , 
	\rst_dat[21][28] , \rst_dat[21][27] , \rst_dat[21][26] , 
	\rst_dat[21][25] , \rst_dat[21][24] , \rst_dat[21][23] , 
	\rst_dat[21][22] , \rst_dat[21][21] , \rst_dat[21][20] , 
	\rst_dat[21][19] , \rst_dat[21][18] , \rst_dat[21][17] , 
	\rst_dat[21][16] , \rst_dat[21][15] , \rst_dat[21][14] , 
	\rst_dat[21][13] , \rst_dat[21][12] , \rst_dat[21][11] , 
	\rst_dat[21][10] , \rst_dat[21][9] , \rst_dat[21][8] , 
	\rst_dat[21][7] , \rst_dat[21][6] , \rst_dat[21][5] , 
	\rst_dat[21][4] , \rst_dat[21][3] , \rst_dat[21][2] , 
	\rst_dat[21][1] , \rst_dat[21][0] , \rst_dat[22][31] , 
	\rst_dat[22][30] , \rst_dat[22][29] , \rst_dat[22][28] , 
	\rst_dat[22][27] , \rst_dat[22][26] , \rst_dat[22][25] , 
	\rst_dat[22][24] , \rst_dat[22][23] , \rst_dat[22][22] , 
	\rst_dat[22][21] , \rst_dat[22][20] , \rst_dat[22][19] , 
	\rst_dat[22][18] , \rst_dat[22][17] , \rst_dat[22][16] , 
	\rst_dat[22][15] , \rst_dat[22][14] , \rst_dat[22][13] , 
	\rst_dat[22][12] , \rst_dat[22][11] , \rst_dat[22][10] , 
	\rst_dat[22][9] , \rst_dat[22][8] , \rst_dat[22][7] , 
	\rst_dat[22][6] , \rst_dat[22][5] , \rst_dat[22][4] , 
	\rst_dat[22][3] , \rst_dat[22][2] , \rst_dat[22][1] , 
	\rst_dat[22][0] , \rst_dat[23][31] , \rst_dat[23][30] , 
	\rst_dat[23][29] , \rst_dat[23][28] , \rst_dat[23][27] , 
	\rst_dat[23][26] , \rst_dat[23][25] , \rst_dat[23][24] , 
	\rst_dat[23][23] , \rst_dat[23][22] , \rst_dat[23][21] , 
	\rst_dat[23][20] , \rst_dat[23][19] , \rst_dat[23][18] , 
	\rst_dat[23][17] , \rst_dat[23][16] , \rst_dat[23][15] , 
	\rst_dat[23][14] , \rst_dat[23][13] , \rst_dat[23][12] , 
	\rst_dat[23][11] , \rst_dat[23][10] , \rst_dat[23][9] , 
	\rst_dat[23][8] , \rst_dat[23][7] , \rst_dat[23][6] , 
	\rst_dat[23][5] , \rst_dat[23][4] , \rst_dat[23][3] , 
	\rst_dat[23][2] , \rst_dat[23][1] , \rst_dat[23][0] , 
	\rst_dat[24][31] , \rst_dat[24][30] , \rst_dat[24][29] , 
	\rst_dat[24][28] , \rst_dat[24][27] , \rst_dat[24][26] , 
	\rst_dat[24][25] , \rst_dat[24][24] , \rst_dat[24][23] , 
	\rst_dat[24][22] , \rst_dat[24][21] , \rst_dat[24][20] , 
	\rst_dat[24][19] , \rst_dat[24][18] , \rst_dat[24][17] , 
	\rst_dat[24][16] , \rst_dat[24][15] , \rst_dat[24][14] , 
	\rst_dat[24][13] , \rst_dat[24][12] , \rst_dat[24][11] , 
	\rst_dat[24][10] , \rst_dat[24][9] , \rst_dat[24][8] , 
	\rst_dat[24][7] , \rst_dat[24][6] , \rst_dat[24][5] , 
	\rst_dat[24][4] , \rst_dat[24][3] , \rst_dat[24][2] , 
	\rst_dat[24][1] , \rst_dat[24][0] , \rst_dat[25][31] , 
	\rst_dat[25][30] , \rst_dat[25][29] , \rst_dat[25][28] , 
	\rst_dat[25][27] , \rst_dat[25][26] , \rst_dat[25][25] , 
	\rst_dat[25][24] , \rst_dat[25][23] , \rst_dat[25][22] , 
	\rst_dat[25][21] , \rst_dat[25][20] , \rst_dat[25][19] , 
	\rst_dat[25][18] , \rst_dat[25][17] , \rst_dat[25][16] , 
	\rst_dat[25][15] , \rst_dat[25][14] , \rst_dat[25][13] , 
	\rst_dat[25][12] , \rst_dat[25][11] , \rst_dat[25][10] , 
	\rst_dat[25][9] , \rst_dat[25][8] , \rst_dat[25][7] , 
	\rst_dat[25][6] , \rst_dat[25][5] , \rst_dat[25][4] , 
	\rst_dat[25][3] , \rst_dat[25][2] , \rst_dat[25][1] , 
	\rst_dat[25][0] , \rst_dat[26][31] , \rst_dat[26][30] , 
	\rst_dat[26][29] , \rst_dat[26][28] , \rst_dat[26][27] , 
	\rst_dat[26][26] , \rst_dat[26][25] , \rst_dat[26][24] , 
	\rst_dat[26][23] , \rst_dat[26][22] , \rst_dat[26][21] , 
	\rst_dat[26][20] , \rst_dat[26][19] , \rst_dat[26][18] , 
	\rst_dat[26][17] , \rst_dat[26][16] , \rst_dat[26][15] , 
	\rst_dat[26][14] , \rst_dat[26][13] , \rst_dat[26][12] , 
	\rst_dat[26][11] , \rst_dat[26][10] , \rst_dat[26][9] , 
	\rst_dat[26][8] , \rst_dat[26][7] , \rst_dat[26][6] , 
	\rst_dat[26][5] , \rst_dat[26][4] , \rst_dat[26][3] , 
	\rst_dat[26][2] , \rst_dat[26][1] , \rst_dat[26][0] , 
	\rst_dat[27][31] , \rst_dat[27][30] , \rst_dat[27][29] , 
	\rst_dat[27][28] , \rst_dat[27][27] , \rst_dat[27][26] , 
	\rst_dat[27][25] , \rst_dat[27][24] , \rst_dat[27][23] , 
	\rst_dat[27][22] , \rst_dat[27][21] , \rst_dat[27][20] , 
	\rst_dat[27][19] , \rst_dat[27][18] , \rst_dat[27][17] , 
	\rst_dat[27][16] , \rst_dat[27][15] , \rst_dat[27][14] , 
	\rst_dat[27][13] , \rst_dat[27][12] , \rst_dat[27][11] , 
	\rst_dat[27][10] , \rst_dat[27][9] , \rst_dat[27][8] , 
	\rst_dat[27][7] , \rst_dat[27][6] , \rst_dat[27][5] , 
	\rst_dat[27][4] , \rst_dat[27][3] , \rst_dat[27][2] , 
	\rst_dat[27][1] , \rst_dat[27][0] , \rst_dat[28][31] , 
	\rst_dat[28][30] , \rst_dat[28][29] , \rst_dat[28][28] , 
	\rst_dat[28][27] , \rst_dat[28][26] , \rst_dat[28][25] , 
	\rst_dat[28][24] , \rst_dat[28][23] , \rst_dat[28][22] , 
	\rst_dat[28][21] , \rst_dat[28][20] , \rst_dat[28][19] , 
	\rst_dat[28][18] , \rst_dat[28][17] , \rst_dat[28][16] , 
	\rst_dat[28][15] , \rst_dat[28][14] , \rst_dat[28][13] , 
	\rst_dat[28][12] , \rst_dat[28][11] , \rst_dat[28][10] , 
	\rst_dat[28][9] , \rst_dat[28][8] , \rst_dat[28][7] , 
	\rst_dat[28][6] , \rst_dat[28][5] , \rst_dat[28][4] , 
	\rst_dat[28][3] , \rst_dat[28][2] , \rst_dat[28][1] , 
	\rst_dat[28][0] , \rst_dat[29][31] , \rst_dat[29][30] , 
	\rst_dat[29][29] , \rst_dat[29][28] , \rst_dat[29][27] , 
	\rst_dat[29][26] , \rst_dat[29][25] , \rst_dat[29][24] , 
	\rst_dat[29][23] , \rst_dat[29][22] , \rst_dat[29][21] , 
	\rst_dat[29][20] , \rst_dat[29][19] , \rst_dat[29][18] , 
	\rst_dat[29][17] , \rst_dat[29][16] , \rst_dat[29][15] , 
	\rst_dat[29][14] , \rst_dat[29][13] , \rst_dat[29][12] , 
	\rst_dat[29][11] , \rst_dat[29][10] , \rst_dat[29][9] , 
	\rst_dat[29][8] , \rst_dat[29][7] , \rst_dat[29][6] , 
	\rst_dat[29][5] , \rst_dat[29][4] , \rst_dat[29][3] , 
	\rst_dat[29][2] , \rst_dat[29][1] , \rst_dat[29][0] , 
	\rst_dat[30][31] , \rst_dat[30][30] , \rst_dat[30][29] , 
	\rst_dat[30][28] , \rst_dat[30][27] , \rst_dat[30][26] , 
	\rst_dat[30][25] , \rst_dat[30][24] , \rst_dat[30][23] , 
	\rst_dat[30][22] , \rst_dat[30][21] , \rst_dat[30][20] , 
	\rst_dat[30][19] , \rst_dat[30][18] , \rst_dat[30][17] , 
	\rst_dat[30][16] , \rst_dat[30][15] , \rst_dat[30][14] , 
	\rst_dat[30][13] , \rst_dat[30][12] , \rst_dat[30][11] , 
	\rst_dat[30][10] , \rst_dat[30][9] , \rst_dat[30][8] , 
	\rst_dat[30][7] , \rst_dat[30][6] , \rst_dat[30][5] , 
	\rst_dat[30][4] , \rst_dat[30][3] , \rst_dat[30][2] , 
	\rst_dat[30][1] , \rst_dat[30][0] , \rst_dat[31][31] , 
	\rst_dat[31][30] , \rst_dat[31][29] , \rst_dat[31][28] , 
	\rst_dat[31][27] , \rst_dat[31][26] , \rst_dat[31][25] , 
	\rst_dat[31][24] , \rst_dat[31][23] , \rst_dat[31][22] , 
	\rst_dat[31][21] , \rst_dat[31][20] , \rst_dat[31][19] , 
	\rst_dat[31][18] , \rst_dat[31][17] , \rst_dat[31][16] , 
	\rst_dat[31][15] , \rst_dat[31][14] , \rst_dat[31][13] , 
	\rst_dat[31][12] , \rst_dat[31][11] , \rst_dat[31][10] , 
	\rst_dat[31][9] , \rst_dat[31][8] , \rst_dat[31][7] , 
	\rst_dat[31][6] , \rst_dat[31][5] , \rst_dat[31][4] , 
	\rst_dat[31][3] , \rst_dat[31][2] , \rst_dat[31][1] , 
	\rst_dat[31][0] } ));
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output [2:0] stat_code;
output [4:0] stat_datawords;
output [4:0] stat_addr;
output [15:0] capability_lst;
output [3:0] capability_type;
output [31:0] rd_dat;
output \mem_a[0][31] ;
output \mem_a[0][30] ;
output \mem_a[0][29] ;
output \mem_a[0][28] ;
output \mem_a[0][27] ;
output \mem_a[0][26] ;
output \mem_a[0][25] ;
output \mem_a[0][24] ;
output \mem_a[0][23] ;
output \mem_a[0][22] ;
output \mem_a[0][21] ;
output \mem_a[0][20] ;
output \mem_a[0][19] ;
output \mem_a[0][18] ;
output \mem_a[0][17] ;
output \mem_a[0][16] ;
output \mem_a[0][15] ;
output \mem_a[0][14] ;
output \mem_a[0][13] ;
output \mem_a[0][12] ;
output \mem_a[0][11] ;
output \mem_a[0][10] ;
output \mem_a[0][9] ;
output \mem_a[0][8] ;
output \mem_a[0][7] ;
output \mem_a[0][6] ;
output \mem_a[0][5] ;
output \mem_a[0][4] ;
output \mem_a[0][3] ;
output \mem_a[0][2] ;
output \mem_a[0][1] ;
output \mem_a[0][0] ;
output \mem_a[1][31] ;
output \mem_a[1][30] ;
output \mem_a[1][29] ;
output \mem_a[1][28] ;
output \mem_a[1][27] ;
output \mem_a[1][26] ;
output \mem_a[1][25] ;
output \mem_a[1][24] ;
output \mem_a[1][23] ;
output \mem_a[1][22] ;
output \mem_a[1][21] ;
output \mem_a[1][20] ;
output \mem_a[1][19] ;
output \mem_a[1][18] ;
output \mem_a[1][17] ;
output \mem_a[1][16] ;
output \mem_a[1][15] ;
output \mem_a[1][14] ;
output \mem_a[1][13] ;
output \mem_a[1][12] ;
output \mem_a[1][11] ;
output \mem_a[1][10] ;
output \mem_a[1][9] ;
output \mem_a[1][8] ;
output \mem_a[1][7] ;
output \mem_a[1][6] ;
output \mem_a[1][5] ;
output \mem_a[1][4] ;
output \mem_a[1][3] ;
output \mem_a[1][2] ;
output \mem_a[1][1] ;
output \mem_a[1][0] ;
output \mem_a[2][31] ;
output \mem_a[2][30] ;
output \mem_a[2][29] ;
output \mem_a[2][28] ;
output \mem_a[2][27] ;
output \mem_a[2][26] ;
output \mem_a[2][25] ;
output \mem_a[2][24] ;
output \mem_a[2][23] ;
output \mem_a[2][22] ;
output \mem_a[2][21] ;
output \mem_a[2][20] ;
output \mem_a[2][19] ;
output \mem_a[2][18] ;
output \mem_a[2][17] ;
output \mem_a[2][16] ;
output \mem_a[2][15] ;
output \mem_a[2][14] ;
output \mem_a[2][13] ;
output \mem_a[2][12] ;
output \mem_a[2][11] ;
output \mem_a[2][10] ;
output \mem_a[2][9] ;
output \mem_a[2][8] ;
output \mem_a[2][7] ;
output \mem_a[2][6] ;
output \mem_a[2][5] ;
output \mem_a[2][4] ;
output \mem_a[2][3] ;
output \mem_a[2][2] ;
output \mem_a[2][1] ;
output \mem_a[2][0] ;
output \mem_a[3][31] ;
output \mem_a[3][30] ;
output \mem_a[3][29] ;
output \mem_a[3][28] ;
output \mem_a[3][27] ;
output \mem_a[3][26] ;
output \mem_a[3][25] ;
output \mem_a[3][24] ;
output \mem_a[3][23] ;
output \mem_a[3][22] ;
output \mem_a[3][21] ;
output \mem_a[3][20] ;
output \mem_a[3][19] ;
output \mem_a[3][18] ;
output \mem_a[3][17] ;
output \mem_a[3][16] ;
output \mem_a[3][15] ;
output \mem_a[3][14] ;
output \mem_a[3][13] ;
output \mem_a[3][12] ;
output \mem_a[3][11] ;
output \mem_a[3][10] ;
output \mem_a[3][9] ;
output \mem_a[3][8] ;
output \mem_a[3][7] ;
output \mem_a[3][6] ;
output \mem_a[3][5] ;
output \mem_a[3][4] ;
output \mem_a[3][3] ;
output \mem_a[3][2] ;
output \mem_a[3][1] ;
output \mem_a[3][0] ;
output \mem_a[4][31] ;
output \mem_a[4][30] ;
output \mem_a[4][29] ;
output \mem_a[4][28] ;
output \mem_a[4][27] ;
output \mem_a[4][26] ;
output \mem_a[4][25] ;
output \mem_a[4][24] ;
output \mem_a[4][23] ;
output \mem_a[4][22] ;
output \mem_a[4][21] ;
output \mem_a[4][20] ;
output \mem_a[4][19] ;
output \mem_a[4][18] ;
output \mem_a[4][17] ;
output \mem_a[4][16] ;
output \mem_a[4][15] ;
output \mem_a[4][14] ;
output \mem_a[4][13] ;
output \mem_a[4][12] ;
output \mem_a[4][11] ;
output \mem_a[4][10] ;
output \mem_a[4][9] ;
output \mem_a[4][8] ;
output \mem_a[4][7] ;
output \mem_a[4][6] ;
output \mem_a[4][5] ;
output \mem_a[4][4] ;
output \mem_a[4][3] ;
output \mem_a[4][2] ;
output \mem_a[4][1] ;
output \mem_a[4][0] ;
output \mem_a[5][31] ;
output \mem_a[5][30] ;
output \mem_a[5][29] ;
output \mem_a[5][28] ;
output \mem_a[5][27] ;
output \mem_a[5][26] ;
output \mem_a[5][25] ;
output \mem_a[5][24] ;
output \mem_a[5][23] ;
output \mem_a[5][22] ;
output \mem_a[5][21] ;
output \mem_a[5][20] ;
output \mem_a[5][19] ;
output \mem_a[5][18] ;
output \mem_a[5][17] ;
output \mem_a[5][16] ;
output \mem_a[5][15] ;
output \mem_a[5][14] ;
output \mem_a[5][13] ;
output \mem_a[5][12] ;
output \mem_a[5][11] ;
output \mem_a[5][10] ;
output \mem_a[5][9] ;
output \mem_a[5][8] ;
output \mem_a[5][7] ;
output \mem_a[5][6] ;
output \mem_a[5][5] ;
output \mem_a[5][4] ;
output \mem_a[5][3] ;
output \mem_a[5][2] ;
output \mem_a[5][1] ;
output \mem_a[5][0] ;
output \mem_a[6][31] ;
output \mem_a[6][30] ;
output \mem_a[6][29] ;
output \mem_a[6][28] ;
output \mem_a[6][27] ;
output \mem_a[6][26] ;
output \mem_a[6][25] ;
output \mem_a[6][24] ;
output \mem_a[6][23] ;
output \mem_a[6][22] ;
output \mem_a[6][21] ;
output \mem_a[6][20] ;
output \mem_a[6][19] ;
output \mem_a[6][18] ;
output \mem_a[6][17] ;
output \mem_a[6][16] ;
output \mem_a[6][15] ;
output \mem_a[6][14] ;
output \mem_a[6][13] ;
output \mem_a[6][12] ;
output \mem_a[6][11] ;
output \mem_a[6][10] ;
output \mem_a[6][9] ;
output \mem_a[6][8] ;
output \mem_a[6][7] ;
output \mem_a[6][6] ;
output \mem_a[6][5] ;
output \mem_a[6][4] ;
output \mem_a[6][3] ;
output \mem_a[6][2] ;
output \mem_a[6][1] ;
output \mem_a[6][0] ;
output \mem_a[7][31] ;
output \mem_a[7][30] ;
output \mem_a[7][29] ;
output \mem_a[7][28] ;
output \mem_a[7][27] ;
output \mem_a[7][26] ;
output \mem_a[7][25] ;
output \mem_a[7][24] ;
output \mem_a[7][23] ;
output \mem_a[7][22] ;
output \mem_a[7][21] ;
output \mem_a[7][20] ;
output \mem_a[7][19] ;
output \mem_a[7][18] ;
output \mem_a[7][17] ;
output \mem_a[7][16] ;
output \mem_a[7][15] ;
output \mem_a[7][14] ;
output \mem_a[7][13] ;
output \mem_a[7][12] ;
output \mem_a[7][11] ;
output \mem_a[7][10] ;
output \mem_a[7][9] ;
output \mem_a[7][8] ;
output \mem_a[7][7] ;
output \mem_a[7][6] ;
output \mem_a[7][5] ;
output \mem_a[7][4] ;
output \mem_a[7][3] ;
output \mem_a[7][2] ;
output \mem_a[7][1] ;
output \mem_a[7][0] ;
output \mem_a[8][31] ;
output \mem_a[8][30] ;
output \mem_a[8][29] ;
output \mem_a[8][28] ;
output \mem_a[8][27] ;
output \mem_a[8][26] ;
output \mem_a[8][25] ;
output \mem_a[8][24] ;
output \mem_a[8][23] ;
output \mem_a[8][22] ;
output \mem_a[8][21] ;
output \mem_a[8][20] ;
output \mem_a[8][19] ;
output \mem_a[8][18] ;
output \mem_a[8][17] ;
output \mem_a[8][16] ;
output \mem_a[8][15] ;
output \mem_a[8][14] ;
output \mem_a[8][13] ;
output \mem_a[8][12] ;
output \mem_a[8][11] ;
output \mem_a[8][10] ;
output \mem_a[8][9] ;
output \mem_a[8][8] ;
output \mem_a[8][7] ;
output \mem_a[8][6] ;
output \mem_a[8][5] ;
output \mem_a[8][4] ;
output \mem_a[8][3] ;
output \mem_a[8][2] ;
output \mem_a[8][1] ;
output \mem_a[8][0] ;
output \mem_a[9][31] ;
output \mem_a[9][30] ;
output \mem_a[9][29] ;
output \mem_a[9][28] ;
output \mem_a[9][27] ;
output \mem_a[9][26] ;
output \mem_a[9][25] ;
output \mem_a[9][24] ;
output \mem_a[9][23] ;
output \mem_a[9][22] ;
output \mem_a[9][21] ;
output \mem_a[9][20] ;
output \mem_a[9][19] ;
output \mem_a[9][18] ;
output \mem_a[9][17] ;
output \mem_a[9][16] ;
output \mem_a[9][15] ;
output \mem_a[9][14] ;
output \mem_a[9][13] ;
output \mem_a[9][12] ;
output \mem_a[9][11] ;
output \mem_a[9][10] ;
output \mem_a[9][9] ;
output \mem_a[9][8] ;
output \mem_a[9][7] ;
output \mem_a[9][6] ;
output \mem_a[9][5] ;
output \mem_a[9][4] ;
output \mem_a[9][3] ;
output \mem_a[9][2] ;
output \mem_a[9][1] ;
output \mem_a[9][0] ;
output \mem_a[10][31] ;
output \mem_a[10][30] ;
output \mem_a[10][29] ;
output \mem_a[10][28] ;
output \mem_a[10][27] ;
output \mem_a[10][26] ;
output \mem_a[10][25] ;
output \mem_a[10][24] ;
output \mem_a[10][23] ;
output \mem_a[10][22] ;
output \mem_a[10][21] ;
output \mem_a[10][20] ;
output \mem_a[10][19] ;
output \mem_a[10][18] ;
output \mem_a[10][17] ;
output \mem_a[10][16] ;
output \mem_a[10][15] ;
output \mem_a[10][14] ;
output \mem_a[10][13] ;
output \mem_a[10][12] ;
output \mem_a[10][11] ;
output \mem_a[10][10] ;
output \mem_a[10][9] ;
output \mem_a[10][8] ;
output \mem_a[10][7] ;
output \mem_a[10][6] ;
output \mem_a[10][5] ;
output \mem_a[10][4] ;
output \mem_a[10][3] ;
output \mem_a[10][2] ;
output \mem_a[10][1] ;
output \mem_a[10][0] ;
output \mem_a[11][31] ;
output \mem_a[11][30] ;
output \mem_a[11][29] ;
output \mem_a[11][28] ;
output \mem_a[11][27] ;
output \mem_a[11][26] ;
output \mem_a[11][25] ;
output \mem_a[11][24] ;
output \mem_a[11][23] ;
output \mem_a[11][22] ;
output \mem_a[11][21] ;
output \mem_a[11][20] ;
output \mem_a[11][19] ;
output \mem_a[11][18] ;
output \mem_a[11][17] ;
output \mem_a[11][16] ;
output \mem_a[11][15] ;
output \mem_a[11][14] ;
output \mem_a[11][13] ;
output \mem_a[11][12] ;
output \mem_a[11][11] ;
output \mem_a[11][10] ;
output \mem_a[11][9] ;
output \mem_a[11][8] ;
output \mem_a[11][7] ;
output \mem_a[11][6] ;
output \mem_a[11][5] ;
output \mem_a[11][4] ;
output \mem_a[11][3] ;
output \mem_a[11][2] ;
output \mem_a[11][1] ;
output \mem_a[11][0] ;
output \mem_a[12][31] ;
output \mem_a[12][30] ;
output \mem_a[12][29] ;
output \mem_a[12][28] ;
output \mem_a[12][27] ;
output \mem_a[12][26] ;
output \mem_a[12][25] ;
output \mem_a[12][24] ;
output \mem_a[12][23] ;
output \mem_a[12][22] ;
output \mem_a[12][21] ;
output \mem_a[12][20] ;
output \mem_a[12][19] ;
output \mem_a[12][18] ;
output \mem_a[12][17] ;
output \mem_a[12][16] ;
output \mem_a[12][15] ;
output \mem_a[12][14] ;
output \mem_a[12][13] ;
output \mem_a[12][12] ;
output \mem_a[12][11] ;
output \mem_a[12][10] ;
output \mem_a[12][9] ;
output \mem_a[12][8] ;
output \mem_a[12][7] ;
output \mem_a[12][6] ;
output \mem_a[12][5] ;
output \mem_a[12][4] ;
output \mem_a[12][3] ;
output \mem_a[12][2] ;
output \mem_a[12][1] ;
output \mem_a[12][0] ;
output \mem_a[13][31] ;
output \mem_a[13][30] ;
output \mem_a[13][29] ;
output \mem_a[13][28] ;
output \mem_a[13][27] ;
output \mem_a[13][26] ;
output \mem_a[13][25] ;
output \mem_a[13][24] ;
output \mem_a[13][23] ;
output \mem_a[13][22] ;
output \mem_a[13][21] ;
output \mem_a[13][20] ;
output \mem_a[13][19] ;
output \mem_a[13][18] ;
output \mem_a[13][17] ;
output \mem_a[13][16] ;
output \mem_a[13][15] ;
output \mem_a[13][14] ;
output \mem_a[13][13] ;
output \mem_a[13][12] ;
output \mem_a[13][11] ;
output \mem_a[13][10] ;
output \mem_a[13][9] ;
output \mem_a[13][8] ;
output \mem_a[13][7] ;
output \mem_a[13][6] ;
output \mem_a[13][5] ;
output \mem_a[13][4] ;
output \mem_a[13][3] ;
output \mem_a[13][2] ;
output \mem_a[13][1] ;
output \mem_a[13][0] ;
output \mem_a[14][31] ;
output \mem_a[14][30] ;
output \mem_a[14][29] ;
output \mem_a[14][28] ;
output \mem_a[14][27] ;
output \mem_a[14][26] ;
output \mem_a[14][25] ;
output \mem_a[14][24] ;
output \mem_a[14][23] ;
output \mem_a[14][22] ;
output \mem_a[14][21] ;
output \mem_a[14][20] ;
output \mem_a[14][19] ;
output \mem_a[14][18] ;
output \mem_a[14][17] ;
output \mem_a[14][16] ;
output \mem_a[14][15] ;
output \mem_a[14][14] ;
output \mem_a[14][13] ;
output \mem_a[14][12] ;
output \mem_a[14][11] ;
output \mem_a[14][10] ;
output \mem_a[14][9] ;
output \mem_a[14][8] ;
output \mem_a[14][7] ;
output \mem_a[14][6] ;
output \mem_a[14][5] ;
output \mem_a[14][4] ;
output \mem_a[14][3] ;
output \mem_a[14][2] ;
output \mem_a[14][1] ;
output \mem_a[14][0] ;
output \mem_a[15][31] ;
output \mem_a[15][30] ;
output \mem_a[15][29] ;
output \mem_a[15][28] ;
output \mem_a[15][27] ;
output \mem_a[15][26] ;
output \mem_a[15][25] ;
output \mem_a[15][24] ;
output \mem_a[15][23] ;
output \mem_a[15][22] ;
output \mem_a[15][21] ;
output \mem_a[15][20] ;
output \mem_a[15][19] ;
output \mem_a[15][18] ;
output \mem_a[15][17] ;
output \mem_a[15][16] ;
output \mem_a[15][15] ;
output \mem_a[15][14] ;
output \mem_a[15][13] ;
output \mem_a[15][12] ;
output \mem_a[15][11] ;
output \mem_a[15][10] ;
output \mem_a[15][9] ;
output \mem_a[15][8] ;
output \mem_a[15][7] ;
output \mem_a[15][6] ;
output \mem_a[15][5] ;
output \mem_a[15][4] ;
output \mem_a[15][3] ;
output \mem_a[15][2] ;
output \mem_a[15][1] ;
output \mem_a[15][0] ;
output \mem_a[16][31] ;
output \mem_a[16][30] ;
output \mem_a[16][29] ;
output \mem_a[16][28] ;
output \mem_a[16][27] ;
output \mem_a[16][26] ;
output \mem_a[16][25] ;
output \mem_a[16][24] ;
output \mem_a[16][23] ;
output \mem_a[16][22] ;
output \mem_a[16][21] ;
output \mem_a[16][20] ;
output \mem_a[16][19] ;
output \mem_a[16][18] ;
output \mem_a[16][17] ;
output \mem_a[16][16] ;
output \mem_a[16][15] ;
output \mem_a[16][14] ;
output \mem_a[16][13] ;
output \mem_a[16][12] ;
output \mem_a[16][11] ;
output \mem_a[16][10] ;
output \mem_a[16][9] ;
output \mem_a[16][8] ;
output \mem_a[16][7] ;
output \mem_a[16][6] ;
output \mem_a[16][5] ;
output \mem_a[16][4] ;
output \mem_a[16][3] ;
output \mem_a[16][2] ;
output \mem_a[16][1] ;
output \mem_a[16][0] ;
output \mem_a[17][31] ;
output \mem_a[17][30] ;
output \mem_a[17][29] ;
output \mem_a[17][28] ;
output \mem_a[17][27] ;
output \mem_a[17][26] ;
output \mem_a[17][25] ;
output \mem_a[17][24] ;
output \mem_a[17][23] ;
output \mem_a[17][22] ;
output \mem_a[17][21] ;
output \mem_a[17][20] ;
output \mem_a[17][19] ;
output \mem_a[17][18] ;
output \mem_a[17][17] ;
output \mem_a[17][16] ;
output \mem_a[17][15] ;
output \mem_a[17][14] ;
output \mem_a[17][13] ;
output \mem_a[17][12] ;
output \mem_a[17][11] ;
output \mem_a[17][10] ;
output \mem_a[17][9] ;
output \mem_a[17][8] ;
output \mem_a[17][7] ;
output \mem_a[17][6] ;
output \mem_a[17][5] ;
output \mem_a[17][4] ;
output \mem_a[17][3] ;
output \mem_a[17][2] ;
output \mem_a[17][1] ;
output \mem_a[17][0] ;
output \mem_a[18][31] ;
output \mem_a[18][30] ;
output \mem_a[18][29] ;
output \mem_a[18][28] ;
output \mem_a[18][27] ;
output \mem_a[18][26] ;
output \mem_a[18][25] ;
output \mem_a[18][24] ;
output \mem_a[18][23] ;
output \mem_a[18][22] ;
output \mem_a[18][21] ;
output \mem_a[18][20] ;
output \mem_a[18][19] ;
output \mem_a[18][18] ;
output \mem_a[18][17] ;
output \mem_a[18][16] ;
output \mem_a[18][15] ;
output \mem_a[18][14] ;
output \mem_a[18][13] ;
output \mem_a[18][12] ;
output \mem_a[18][11] ;
output \mem_a[18][10] ;
output \mem_a[18][9] ;
output \mem_a[18][8] ;
output \mem_a[18][7] ;
output \mem_a[18][6] ;
output \mem_a[18][5] ;
output \mem_a[18][4] ;
output \mem_a[18][3] ;
output \mem_a[18][2] ;
output \mem_a[18][1] ;
output \mem_a[18][0] ;
output \mem_a[19][31] ;
output \mem_a[19][30] ;
output \mem_a[19][29] ;
output \mem_a[19][28] ;
output \mem_a[19][27] ;
output \mem_a[19][26] ;
output \mem_a[19][25] ;
output \mem_a[19][24] ;
output \mem_a[19][23] ;
output \mem_a[19][22] ;
output \mem_a[19][21] ;
output \mem_a[19][20] ;
output \mem_a[19][19] ;
output \mem_a[19][18] ;
output \mem_a[19][17] ;
output \mem_a[19][16] ;
output \mem_a[19][15] ;
output \mem_a[19][14] ;
output \mem_a[19][13] ;
output \mem_a[19][12] ;
output \mem_a[19][11] ;
output \mem_a[19][10] ;
output \mem_a[19][9] ;
output \mem_a[19][8] ;
output \mem_a[19][7] ;
output \mem_a[19][6] ;
output \mem_a[19][5] ;
output \mem_a[19][4] ;
output \mem_a[19][3] ;
output \mem_a[19][2] ;
output \mem_a[19][1] ;
output \mem_a[19][0] ;
output \mem_a[20][31] ;
output \mem_a[20][30] ;
output \mem_a[20][29] ;
output \mem_a[20][28] ;
output \mem_a[20][27] ;
output \mem_a[20][26] ;
output \mem_a[20][25] ;
output \mem_a[20][24] ;
output \mem_a[20][23] ;
output \mem_a[20][22] ;
output \mem_a[20][21] ;
output \mem_a[20][20] ;
output \mem_a[20][19] ;
output \mem_a[20][18] ;
output \mem_a[20][17] ;
output \mem_a[20][16] ;
output \mem_a[20][15] ;
output \mem_a[20][14] ;
output \mem_a[20][13] ;
output \mem_a[20][12] ;
output \mem_a[20][11] ;
output \mem_a[20][10] ;
output \mem_a[20][9] ;
output \mem_a[20][8] ;
output \mem_a[20][7] ;
output \mem_a[20][6] ;
output \mem_a[20][5] ;
output \mem_a[20][4] ;
output \mem_a[20][3] ;
output \mem_a[20][2] ;
output \mem_a[20][1] ;
output \mem_a[20][0] ;
output \mem_a[21][31] ;
output \mem_a[21][30] ;
output \mem_a[21][29] ;
output \mem_a[21][28] ;
output \mem_a[21][27] ;
output \mem_a[21][26] ;
output \mem_a[21][25] ;
output \mem_a[21][24] ;
output \mem_a[21][23] ;
output \mem_a[21][22] ;
output \mem_a[21][21] ;
output \mem_a[21][20] ;
output \mem_a[21][19] ;
output \mem_a[21][18] ;
output \mem_a[21][17] ;
output \mem_a[21][16] ;
output \mem_a[21][15] ;
output \mem_a[21][14] ;
output \mem_a[21][13] ;
output \mem_a[21][12] ;
output \mem_a[21][11] ;
output \mem_a[21][10] ;
output \mem_a[21][9] ;
output \mem_a[21][8] ;
output \mem_a[21][7] ;
output \mem_a[21][6] ;
output \mem_a[21][5] ;
output \mem_a[21][4] ;
output \mem_a[21][3] ;
output \mem_a[21][2] ;
output \mem_a[21][1] ;
output \mem_a[21][0] ;
output \mem_a[22][31] ;
output \mem_a[22][30] ;
output \mem_a[22][29] ;
output \mem_a[22][28] ;
output \mem_a[22][27] ;
output \mem_a[22][26] ;
output \mem_a[22][25] ;
output \mem_a[22][24] ;
output \mem_a[22][23] ;
output \mem_a[22][22] ;
output \mem_a[22][21] ;
output \mem_a[22][20] ;
output \mem_a[22][19] ;
output \mem_a[22][18] ;
output \mem_a[22][17] ;
output \mem_a[22][16] ;
output \mem_a[22][15] ;
output \mem_a[22][14] ;
output \mem_a[22][13] ;
output \mem_a[22][12] ;
output \mem_a[22][11] ;
output \mem_a[22][10] ;
output \mem_a[22][9] ;
output \mem_a[22][8] ;
output \mem_a[22][7] ;
output \mem_a[22][6] ;
output \mem_a[22][5] ;
output \mem_a[22][4] ;
output \mem_a[22][3] ;
output \mem_a[22][2] ;
output \mem_a[22][1] ;
output \mem_a[22][0] ;
output \mem_a[23][31] ;
output \mem_a[23][30] ;
output \mem_a[23][29] ;
output \mem_a[23][28] ;
output \mem_a[23][27] ;
output \mem_a[23][26] ;
output \mem_a[23][25] ;
output \mem_a[23][24] ;
output \mem_a[23][23] ;
output \mem_a[23][22] ;
output \mem_a[23][21] ;
output \mem_a[23][20] ;
output \mem_a[23][19] ;
output \mem_a[23][18] ;
output \mem_a[23][17] ;
output \mem_a[23][16] ;
output \mem_a[23][15] ;
output \mem_a[23][14] ;
output \mem_a[23][13] ;
output \mem_a[23][12] ;
output \mem_a[23][11] ;
output \mem_a[23][10] ;
output \mem_a[23][9] ;
output \mem_a[23][8] ;
output \mem_a[23][7] ;
output \mem_a[23][6] ;
output \mem_a[23][5] ;
output \mem_a[23][4] ;
output \mem_a[23][3] ;
output \mem_a[23][2] ;
output \mem_a[23][1] ;
output \mem_a[23][0] ;
output \mem_a[24][31] ;
output \mem_a[24][30] ;
output \mem_a[24][29] ;
output \mem_a[24][28] ;
output \mem_a[24][27] ;
output \mem_a[24][26] ;
output \mem_a[24][25] ;
output \mem_a[24][24] ;
output \mem_a[24][23] ;
output \mem_a[24][22] ;
output \mem_a[24][21] ;
output \mem_a[24][20] ;
output \mem_a[24][19] ;
output \mem_a[24][18] ;
output \mem_a[24][17] ;
output \mem_a[24][16] ;
output \mem_a[24][15] ;
output \mem_a[24][14] ;
output \mem_a[24][13] ;
output \mem_a[24][12] ;
output \mem_a[24][11] ;
output \mem_a[24][10] ;
output \mem_a[24][9] ;
output \mem_a[24][8] ;
output \mem_a[24][7] ;
output \mem_a[24][6] ;
output \mem_a[24][5] ;
output \mem_a[24][4] ;
output \mem_a[24][3] ;
output \mem_a[24][2] ;
output \mem_a[24][1] ;
output \mem_a[24][0] ;
output \mem_a[25][31] ;
output \mem_a[25][30] ;
output \mem_a[25][29] ;
output \mem_a[25][28] ;
output \mem_a[25][27] ;
output \mem_a[25][26] ;
output \mem_a[25][25] ;
output \mem_a[25][24] ;
output \mem_a[25][23] ;
output \mem_a[25][22] ;
output \mem_a[25][21] ;
output \mem_a[25][20] ;
output \mem_a[25][19] ;
output \mem_a[25][18] ;
output \mem_a[25][17] ;
output \mem_a[25][16] ;
output \mem_a[25][15] ;
output \mem_a[25][14] ;
output \mem_a[25][13] ;
output \mem_a[25][12] ;
output \mem_a[25][11] ;
output \mem_a[25][10] ;
output \mem_a[25][9] ;
output \mem_a[25][8] ;
output \mem_a[25][7] ;
output \mem_a[25][6] ;
output \mem_a[25][5] ;
output \mem_a[25][4] ;
output \mem_a[25][3] ;
output \mem_a[25][2] ;
output \mem_a[25][1] ;
output \mem_a[25][0] ;
output \mem_a[26][31] ;
output \mem_a[26][30] ;
output \mem_a[26][29] ;
output \mem_a[26][28] ;
output \mem_a[26][27] ;
output \mem_a[26][26] ;
output \mem_a[26][25] ;
output \mem_a[26][24] ;
output \mem_a[26][23] ;
output \mem_a[26][22] ;
output \mem_a[26][21] ;
output \mem_a[26][20] ;
output \mem_a[26][19] ;
output \mem_a[26][18] ;
output \mem_a[26][17] ;
output \mem_a[26][16] ;
output \mem_a[26][15] ;
output \mem_a[26][14] ;
output \mem_a[26][13] ;
output \mem_a[26][12] ;
output \mem_a[26][11] ;
output \mem_a[26][10] ;
output \mem_a[26][9] ;
output \mem_a[26][8] ;
output \mem_a[26][7] ;
output \mem_a[26][6] ;
output \mem_a[26][5] ;
output \mem_a[26][4] ;
output \mem_a[26][3] ;
output \mem_a[26][2] ;
output \mem_a[26][1] ;
output \mem_a[26][0] ;
output \mem_a[27][31] ;
output \mem_a[27][30] ;
output \mem_a[27][29] ;
output \mem_a[27][28] ;
output \mem_a[27][27] ;
output \mem_a[27][26] ;
output \mem_a[27][25] ;
output \mem_a[27][24] ;
output \mem_a[27][23] ;
output \mem_a[27][22] ;
output \mem_a[27][21] ;
output \mem_a[27][20] ;
output \mem_a[27][19] ;
output \mem_a[27][18] ;
output \mem_a[27][17] ;
output \mem_a[27][16] ;
output \mem_a[27][15] ;
output \mem_a[27][14] ;
output \mem_a[27][13] ;
output \mem_a[27][12] ;
output \mem_a[27][11] ;
output \mem_a[27][10] ;
output \mem_a[27][9] ;
output \mem_a[27][8] ;
output \mem_a[27][7] ;
output \mem_a[27][6] ;
output \mem_a[27][5] ;
output \mem_a[27][4] ;
output \mem_a[27][3] ;
output \mem_a[27][2] ;
output \mem_a[27][1] ;
output \mem_a[27][0] ;
output \mem_a[28][31] ;
output \mem_a[28][30] ;
output \mem_a[28][29] ;
output \mem_a[28][28] ;
output \mem_a[28][27] ;
output \mem_a[28][26] ;
output \mem_a[28][25] ;
output \mem_a[28][24] ;
output \mem_a[28][23] ;
output \mem_a[28][22] ;
output \mem_a[28][21] ;
output \mem_a[28][20] ;
output \mem_a[28][19] ;
output \mem_a[28][18] ;
output \mem_a[28][17] ;
output \mem_a[28][16] ;
output \mem_a[28][15] ;
output \mem_a[28][14] ;
output \mem_a[28][13] ;
output \mem_a[28][12] ;
output \mem_a[28][11] ;
output \mem_a[28][10] ;
output \mem_a[28][9] ;
output \mem_a[28][8] ;
output \mem_a[28][7] ;
output \mem_a[28][6] ;
output \mem_a[28][5] ;
output \mem_a[28][4] ;
output \mem_a[28][3] ;
output \mem_a[28][2] ;
output \mem_a[28][1] ;
output \mem_a[28][0] ;
output \mem_a[29][31] ;
output \mem_a[29][30] ;
output \mem_a[29][29] ;
output \mem_a[29][28] ;
output \mem_a[29][27] ;
output \mem_a[29][26] ;
output \mem_a[29][25] ;
output \mem_a[29][24] ;
output \mem_a[29][23] ;
output \mem_a[29][22] ;
output \mem_a[29][21] ;
output \mem_a[29][20] ;
output \mem_a[29][19] ;
output \mem_a[29][18] ;
output \mem_a[29][17] ;
output \mem_a[29][16] ;
output \mem_a[29][15] ;
output \mem_a[29][14] ;
output \mem_a[29][13] ;
output \mem_a[29][12] ;
output \mem_a[29][11] ;
output \mem_a[29][10] ;
output \mem_a[29][9] ;
output \mem_a[29][8] ;
output \mem_a[29][7] ;
output \mem_a[29][6] ;
output \mem_a[29][5] ;
output \mem_a[29][4] ;
output \mem_a[29][3] ;
output \mem_a[29][2] ;
output \mem_a[29][1] ;
output \mem_a[29][0] ;
output \mem_a[30][31] ;
output \mem_a[30][30] ;
output \mem_a[30][29] ;
output \mem_a[30][28] ;
output \mem_a[30][27] ;
output \mem_a[30][26] ;
output \mem_a[30][25] ;
output \mem_a[30][24] ;
output \mem_a[30][23] ;
output \mem_a[30][22] ;
output \mem_a[30][21] ;
output \mem_a[30][20] ;
output \mem_a[30][19] ;
output \mem_a[30][18] ;
output \mem_a[30][17] ;
output \mem_a[30][16] ;
output \mem_a[30][15] ;
output \mem_a[30][14] ;
output \mem_a[30][13] ;
output \mem_a[30][12] ;
output \mem_a[30][11] ;
output \mem_a[30][10] ;
output \mem_a[30][9] ;
output \mem_a[30][8] ;
output \mem_a[30][7] ;
output \mem_a[30][6] ;
output \mem_a[30][5] ;
output \mem_a[30][4] ;
output \mem_a[30][3] ;
output \mem_a[30][2] ;
output \mem_a[30][1] ;
output \mem_a[30][0] ;
output \mem_a[31][31] ;
output \mem_a[31][30] ;
output \mem_a[31][29] ;
output \mem_a[31][28] ;
output \mem_a[31][27] ;
output \mem_a[31][26] ;
output \mem_a[31][25] ;
output \mem_a[31][24] ;
output \mem_a[31][23] ;
output \mem_a[31][22] ;
output \mem_a[31][21] ;
output \mem_a[31][20] ;
output \mem_a[31][19] ;
output \mem_a[31][18] ;
output \mem_a[31][17] ;
output \mem_a[31][16] ;
output \mem_a[31][15] ;
output \mem_a[31][14] ;
output \mem_a[31][13] ;
output \mem_a[31][12] ;
output \mem_a[31][11] ;
output \mem_a[31][10] ;
output \mem_a[31][9] ;
output \mem_a[31][8] ;
output \mem_a[31][7] ;
output \mem_a[31][6] ;
output \mem_a[31][5] ;
output \mem_a[31][4] ;
output \mem_a[31][3] ;
output \mem_a[31][2] ;
output \mem_a[31][1] ;
output \mem_a[31][0] ;
input clk;
input rst_n;
input [10:0] addr;
input [3:0] cmnd_op;
input [4:0] cmnd_addr;
input wr_stb;
input [31:0] wr_dat;
input \rst_dat[0][31] ;
input \rst_dat[0][30] ;
input \rst_dat[0][29] ;
input \rst_dat[0][28] ;
input \rst_dat[0][27] ;
input \rst_dat[0][26] ;
input \rst_dat[0][25] ;
input \rst_dat[0][24] ;
input \rst_dat[0][23] ;
input \rst_dat[0][22] ;
input \rst_dat[0][21] ;
input \rst_dat[0][20] ;
input \rst_dat[0][19] ;
input \rst_dat[0][18] ;
input \rst_dat[0][17] ;
input \rst_dat[0][16] ;
input \rst_dat[0][15] ;
input \rst_dat[0][14] ;
input \rst_dat[0][13] ;
input \rst_dat[0][12] ;
input \rst_dat[0][11] ;
input \rst_dat[0][10] ;
input \rst_dat[0][9] ;
input \rst_dat[0][8] ;
input \rst_dat[0][7] ;
input \rst_dat[0][6] ;
input \rst_dat[0][5] ;
input \rst_dat[0][4] ;
input \rst_dat[0][3] ;
input \rst_dat[0][2] ;
input \rst_dat[0][1] ;
input \rst_dat[0][0] ;
input \rst_dat[1][31] ;
input \rst_dat[1][30] ;
input \rst_dat[1][29] ;
input \rst_dat[1][28] ;
input \rst_dat[1][27] ;
input \rst_dat[1][26] ;
input \rst_dat[1][25] ;
input \rst_dat[1][24] ;
input \rst_dat[1][23] ;
input \rst_dat[1][22] ;
input \rst_dat[1][21] ;
input \rst_dat[1][20] ;
input \rst_dat[1][19] ;
input \rst_dat[1][18] ;
input \rst_dat[1][17] ;
input \rst_dat[1][16] ;
input \rst_dat[1][15] ;
input \rst_dat[1][14] ;
input \rst_dat[1][13] ;
input \rst_dat[1][12] ;
input \rst_dat[1][11] ;
input \rst_dat[1][10] ;
input \rst_dat[1][9] ;
input \rst_dat[1][8] ;
input \rst_dat[1][7] ;
input \rst_dat[1][6] ;
input \rst_dat[1][5] ;
input \rst_dat[1][4] ;
input \rst_dat[1][3] ;
input \rst_dat[1][2] ;
input \rst_dat[1][1] ;
input \rst_dat[1][0] ;
input \rst_dat[2][31] ;
input \rst_dat[2][30] ;
input \rst_dat[2][29] ;
input \rst_dat[2][28] ;
input \rst_dat[2][27] ;
input \rst_dat[2][26] ;
input \rst_dat[2][25] ;
input \rst_dat[2][24] ;
input \rst_dat[2][23] ;
input \rst_dat[2][22] ;
input \rst_dat[2][21] ;
input \rst_dat[2][20] ;
input \rst_dat[2][19] ;
input \rst_dat[2][18] ;
input \rst_dat[2][17] ;
input \rst_dat[2][16] ;
input \rst_dat[2][15] ;
input \rst_dat[2][14] ;
input \rst_dat[2][13] ;
input \rst_dat[2][12] ;
input \rst_dat[2][11] ;
input \rst_dat[2][10] ;
input \rst_dat[2][9] ;
input \rst_dat[2][8] ;
input \rst_dat[2][7] ;
input \rst_dat[2][6] ;
input \rst_dat[2][5] ;
input \rst_dat[2][4] ;
input \rst_dat[2][3] ;
input \rst_dat[2][2] ;
input \rst_dat[2][1] ;
input \rst_dat[2][0] ;
input \rst_dat[3][31] ;
input \rst_dat[3][30] ;
input \rst_dat[3][29] ;
input \rst_dat[3][28] ;
input \rst_dat[3][27] ;
input \rst_dat[3][26] ;
input \rst_dat[3][25] ;
input \rst_dat[3][24] ;
input \rst_dat[3][23] ;
input \rst_dat[3][22] ;
input \rst_dat[3][21] ;
input \rst_dat[3][20] ;
input \rst_dat[3][19] ;
input \rst_dat[3][18] ;
input \rst_dat[3][17] ;
input \rst_dat[3][16] ;
input \rst_dat[3][15] ;
input \rst_dat[3][14] ;
input \rst_dat[3][13] ;
input \rst_dat[3][12] ;
input \rst_dat[3][11] ;
input \rst_dat[3][10] ;
input \rst_dat[3][9] ;
input \rst_dat[3][8] ;
input \rst_dat[3][7] ;
input \rst_dat[3][6] ;
input \rst_dat[3][5] ;
input \rst_dat[3][4] ;
input \rst_dat[3][3] ;
input \rst_dat[3][2] ;
input \rst_dat[3][1] ;
input \rst_dat[3][0] ;
input \rst_dat[4][31] ;
input \rst_dat[4][30] ;
input \rst_dat[4][29] ;
input \rst_dat[4][28] ;
input \rst_dat[4][27] ;
input \rst_dat[4][26] ;
input \rst_dat[4][25] ;
input \rst_dat[4][24] ;
input \rst_dat[4][23] ;
input \rst_dat[4][22] ;
input \rst_dat[4][21] ;
input \rst_dat[4][20] ;
input \rst_dat[4][19] ;
input \rst_dat[4][18] ;
input \rst_dat[4][17] ;
input \rst_dat[4][16] ;
input \rst_dat[4][15] ;
input \rst_dat[4][14] ;
input \rst_dat[4][13] ;
input \rst_dat[4][12] ;
input \rst_dat[4][11] ;
input \rst_dat[4][10] ;
input \rst_dat[4][9] ;
input \rst_dat[4][8] ;
input \rst_dat[4][7] ;
input \rst_dat[4][6] ;
input \rst_dat[4][5] ;
input \rst_dat[4][4] ;
input \rst_dat[4][3] ;
input \rst_dat[4][2] ;
input \rst_dat[4][1] ;
input \rst_dat[4][0] ;
input \rst_dat[5][31] ;
input \rst_dat[5][30] ;
input \rst_dat[5][29] ;
input \rst_dat[5][28] ;
input \rst_dat[5][27] ;
input \rst_dat[5][26] ;
input \rst_dat[5][25] ;
input \rst_dat[5][24] ;
input \rst_dat[5][23] ;
input \rst_dat[5][22] ;
input \rst_dat[5][21] ;
input \rst_dat[5][20] ;
input \rst_dat[5][19] ;
input \rst_dat[5][18] ;
input \rst_dat[5][17] ;
input \rst_dat[5][16] ;
input \rst_dat[5][15] ;
input \rst_dat[5][14] ;
input \rst_dat[5][13] ;
input \rst_dat[5][12] ;
input \rst_dat[5][11] ;
input \rst_dat[5][10] ;
input \rst_dat[5][9] ;
input \rst_dat[5][8] ;
input \rst_dat[5][7] ;
input \rst_dat[5][6] ;
input \rst_dat[5][5] ;
input \rst_dat[5][4] ;
input \rst_dat[5][3] ;
input \rst_dat[5][2] ;
input \rst_dat[5][1] ;
input \rst_dat[5][0] ;
input \rst_dat[6][31] ;
input \rst_dat[6][30] ;
input \rst_dat[6][29] ;
input \rst_dat[6][28] ;
input \rst_dat[6][27] ;
input \rst_dat[6][26] ;
input \rst_dat[6][25] ;
input \rst_dat[6][24] ;
input \rst_dat[6][23] ;
input \rst_dat[6][22] ;
input \rst_dat[6][21] ;
input \rst_dat[6][20] ;
input \rst_dat[6][19] ;
input \rst_dat[6][18] ;
input \rst_dat[6][17] ;
input \rst_dat[6][16] ;
input \rst_dat[6][15] ;
input \rst_dat[6][14] ;
input \rst_dat[6][13] ;
input \rst_dat[6][12] ;
input \rst_dat[6][11] ;
input \rst_dat[6][10] ;
input \rst_dat[6][9] ;
input \rst_dat[6][8] ;
input \rst_dat[6][7] ;
input \rst_dat[6][6] ;
input \rst_dat[6][5] ;
input \rst_dat[6][4] ;
input \rst_dat[6][3] ;
input \rst_dat[6][2] ;
input \rst_dat[6][1] ;
input \rst_dat[6][0] ;
input \rst_dat[7][31] ;
input \rst_dat[7][30] ;
input \rst_dat[7][29] ;
input \rst_dat[7][28] ;
input \rst_dat[7][27] ;
input \rst_dat[7][26] ;
input \rst_dat[7][25] ;
input \rst_dat[7][24] ;
input \rst_dat[7][23] ;
input \rst_dat[7][22] ;
input \rst_dat[7][21] ;
input \rst_dat[7][20] ;
input \rst_dat[7][19] ;
input \rst_dat[7][18] ;
input \rst_dat[7][17] ;
input \rst_dat[7][16] ;
input \rst_dat[7][15] ;
input \rst_dat[7][14] ;
input \rst_dat[7][13] ;
input \rst_dat[7][12] ;
input \rst_dat[7][11] ;
input \rst_dat[7][10] ;
input \rst_dat[7][9] ;
input \rst_dat[7][8] ;
input \rst_dat[7][7] ;
input \rst_dat[7][6] ;
input \rst_dat[7][5] ;
input \rst_dat[7][4] ;
input \rst_dat[7][3] ;
input \rst_dat[7][2] ;
input \rst_dat[7][1] ;
input \rst_dat[7][0] ;
input \rst_dat[8][31] ;
input \rst_dat[8][30] ;
input \rst_dat[8][29] ;
input \rst_dat[8][28] ;
input \rst_dat[8][27] ;
input \rst_dat[8][26] ;
input \rst_dat[8][25] ;
input \rst_dat[8][24] ;
input \rst_dat[8][23] ;
input \rst_dat[8][22] ;
input \rst_dat[8][21] ;
input \rst_dat[8][20] ;
input \rst_dat[8][19] ;
input \rst_dat[8][18] ;
input \rst_dat[8][17] ;
input \rst_dat[8][16] ;
input \rst_dat[8][15] ;
input \rst_dat[8][14] ;
input \rst_dat[8][13] ;
input \rst_dat[8][12] ;
input \rst_dat[8][11] ;
input \rst_dat[8][10] ;
input \rst_dat[8][9] ;
input \rst_dat[8][8] ;
input \rst_dat[8][7] ;
input \rst_dat[8][6] ;
input \rst_dat[8][5] ;
input \rst_dat[8][4] ;
input \rst_dat[8][3] ;
input \rst_dat[8][2] ;
input \rst_dat[8][1] ;
input \rst_dat[8][0] ;
input \rst_dat[9][31] ;
input \rst_dat[9][30] ;
input \rst_dat[9][29] ;
input \rst_dat[9][28] ;
input \rst_dat[9][27] ;
input \rst_dat[9][26] ;
input \rst_dat[9][25] ;
input \rst_dat[9][24] ;
input \rst_dat[9][23] ;
input \rst_dat[9][22] ;
input \rst_dat[9][21] ;
input \rst_dat[9][20] ;
input \rst_dat[9][19] ;
input \rst_dat[9][18] ;
input \rst_dat[9][17] ;
input \rst_dat[9][16] ;
input \rst_dat[9][15] ;
input \rst_dat[9][14] ;
input \rst_dat[9][13] ;
input \rst_dat[9][12] ;
input \rst_dat[9][11] ;
input \rst_dat[9][10] ;
input \rst_dat[9][9] ;
input \rst_dat[9][8] ;
input \rst_dat[9][7] ;
input \rst_dat[9][6] ;
input \rst_dat[9][5] ;
input \rst_dat[9][4] ;
input \rst_dat[9][3] ;
input \rst_dat[9][2] ;
input \rst_dat[9][1] ;
input \rst_dat[9][0] ;
input \rst_dat[10][31] ;
input \rst_dat[10][30] ;
input \rst_dat[10][29] ;
input \rst_dat[10][28] ;
input \rst_dat[10][27] ;
input \rst_dat[10][26] ;
input \rst_dat[10][25] ;
input \rst_dat[10][24] ;
input \rst_dat[10][23] ;
input \rst_dat[10][22] ;
input \rst_dat[10][21] ;
input \rst_dat[10][20] ;
input \rst_dat[10][19] ;
input \rst_dat[10][18] ;
input \rst_dat[10][17] ;
input \rst_dat[10][16] ;
input \rst_dat[10][15] ;
input \rst_dat[10][14] ;
input \rst_dat[10][13] ;
input \rst_dat[10][12] ;
input \rst_dat[10][11] ;
input \rst_dat[10][10] ;
input \rst_dat[10][9] ;
input \rst_dat[10][8] ;
input \rst_dat[10][7] ;
input \rst_dat[10][6] ;
input \rst_dat[10][5] ;
input \rst_dat[10][4] ;
input \rst_dat[10][3] ;
input \rst_dat[10][2] ;
input \rst_dat[10][1] ;
input \rst_dat[10][0] ;
input \rst_dat[11][31] ;
input \rst_dat[11][30] ;
input \rst_dat[11][29] ;
input \rst_dat[11][28] ;
input \rst_dat[11][27] ;
input \rst_dat[11][26] ;
input \rst_dat[11][25] ;
input \rst_dat[11][24] ;
input \rst_dat[11][23] ;
input \rst_dat[11][22] ;
input \rst_dat[11][21] ;
input \rst_dat[11][20] ;
input \rst_dat[11][19] ;
input \rst_dat[11][18] ;
input \rst_dat[11][17] ;
input \rst_dat[11][16] ;
input \rst_dat[11][15] ;
input \rst_dat[11][14] ;
input \rst_dat[11][13] ;
input \rst_dat[11][12] ;
input \rst_dat[11][11] ;
input \rst_dat[11][10] ;
input \rst_dat[11][9] ;
input \rst_dat[11][8] ;
input \rst_dat[11][7] ;
input \rst_dat[11][6] ;
input \rst_dat[11][5] ;
input \rst_dat[11][4] ;
input \rst_dat[11][3] ;
input \rst_dat[11][2] ;
input \rst_dat[11][1] ;
input \rst_dat[11][0] ;
input \rst_dat[12][31] ;
input \rst_dat[12][30] ;
input \rst_dat[12][29] ;
input \rst_dat[12][28] ;
input \rst_dat[12][27] ;
input \rst_dat[12][26] ;
input \rst_dat[12][25] ;
input \rst_dat[12][24] ;
input \rst_dat[12][23] ;
input \rst_dat[12][22] ;
input \rst_dat[12][21] ;
input \rst_dat[12][20] ;
input \rst_dat[12][19] ;
input \rst_dat[12][18] ;
input \rst_dat[12][17] ;
input \rst_dat[12][16] ;
input \rst_dat[12][15] ;
input \rst_dat[12][14] ;
input \rst_dat[12][13] ;
input \rst_dat[12][12] ;
input \rst_dat[12][11] ;
input \rst_dat[12][10] ;
input \rst_dat[12][9] ;
input \rst_dat[12][8] ;
input \rst_dat[12][7] ;
input \rst_dat[12][6] ;
input \rst_dat[12][5] ;
input \rst_dat[12][4] ;
input \rst_dat[12][3] ;
input \rst_dat[12][2] ;
input \rst_dat[12][1] ;
input \rst_dat[12][0] ;
input \rst_dat[13][31] ;
input \rst_dat[13][30] ;
input \rst_dat[13][29] ;
input \rst_dat[13][28] ;
input \rst_dat[13][27] ;
input \rst_dat[13][26] ;
input \rst_dat[13][25] ;
input \rst_dat[13][24] ;
input \rst_dat[13][23] ;
input \rst_dat[13][22] ;
input \rst_dat[13][21] ;
input \rst_dat[13][20] ;
input \rst_dat[13][19] ;
input \rst_dat[13][18] ;
input \rst_dat[13][17] ;
input \rst_dat[13][16] ;
input \rst_dat[13][15] ;
input \rst_dat[13][14] ;
input \rst_dat[13][13] ;
input \rst_dat[13][12] ;
input \rst_dat[13][11] ;
input \rst_dat[13][10] ;
input \rst_dat[13][9] ;
input \rst_dat[13][8] ;
input \rst_dat[13][7] ;
input \rst_dat[13][6] ;
input \rst_dat[13][5] ;
input \rst_dat[13][4] ;
input \rst_dat[13][3] ;
input \rst_dat[13][2] ;
input \rst_dat[13][1] ;
input \rst_dat[13][0] ;
input \rst_dat[14][31] ;
input \rst_dat[14][30] ;
input \rst_dat[14][29] ;
input \rst_dat[14][28] ;
input \rst_dat[14][27] ;
input \rst_dat[14][26] ;
input \rst_dat[14][25] ;
input \rst_dat[14][24] ;
input \rst_dat[14][23] ;
input \rst_dat[14][22] ;
input \rst_dat[14][21] ;
input \rst_dat[14][20] ;
input \rst_dat[14][19] ;
input \rst_dat[14][18] ;
input \rst_dat[14][17] ;
input \rst_dat[14][16] ;
input \rst_dat[14][15] ;
input \rst_dat[14][14] ;
input \rst_dat[14][13] ;
input \rst_dat[14][12] ;
input \rst_dat[14][11] ;
input \rst_dat[14][10] ;
input \rst_dat[14][9] ;
input \rst_dat[14][8] ;
input \rst_dat[14][7] ;
input \rst_dat[14][6] ;
input \rst_dat[14][5] ;
input \rst_dat[14][4] ;
input \rst_dat[14][3] ;
input \rst_dat[14][2] ;
input \rst_dat[14][1] ;
input \rst_dat[14][0] ;
input \rst_dat[15][31] ;
input \rst_dat[15][30] ;
input \rst_dat[15][29] ;
input \rst_dat[15][28] ;
input \rst_dat[15][27] ;
input \rst_dat[15][26] ;
input \rst_dat[15][25] ;
input \rst_dat[15][24] ;
input \rst_dat[15][23] ;
input \rst_dat[15][22] ;
input \rst_dat[15][21] ;
input \rst_dat[15][20] ;
input \rst_dat[15][19] ;
input \rst_dat[15][18] ;
input \rst_dat[15][17] ;
input \rst_dat[15][16] ;
input \rst_dat[15][15] ;
input \rst_dat[15][14] ;
input \rst_dat[15][13] ;
input \rst_dat[15][12] ;
input \rst_dat[15][11] ;
input \rst_dat[15][10] ;
input \rst_dat[15][9] ;
input \rst_dat[15][8] ;
input \rst_dat[15][7] ;
input \rst_dat[15][6] ;
input \rst_dat[15][5] ;
input \rst_dat[15][4] ;
input \rst_dat[15][3] ;
input \rst_dat[15][2] ;
input \rst_dat[15][1] ;
input \rst_dat[15][0] ;
input \rst_dat[16][31] ;
input \rst_dat[16][30] ;
input \rst_dat[16][29] ;
input \rst_dat[16][28] ;
input \rst_dat[16][27] ;
input \rst_dat[16][26] ;
input \rst_dat[16][25] ;
input \rst_dat[16][24] ;
input \rst_dat[16][23] ;
input \rst_dat[16][22] ;
input \rst_dat[16][21] ;
input \rst_dat[16][20] ;
input \rst_dat[16][19] ;
input \rst_dat[16][18] ;
input \rst_dat[16][17] ;
input \rst_dat[16][16] ;
input \rst_dat[16][15] ;
input \rst_dat[16][14] ;
input \rst_dat[16][13] ;
input \rst_dat[16][12] ;
input \rst_dat[16][11] ;
input \rst_dat[16][10] ;
input \rst_dat[16][9] ;
input \rst_dat[16][8] ;
input \rst_dat[16][7] ;
input \rst_dat[16][6] ;
input \rst_dat[16][5] ;
input \rst_dat[16][4] ;
input \rst_dat[16][3] ;
input \rst_dat[16][2] ;
input \rst_dat[16][1] ;
input \rst_dat[16][0] ;
input \rst_dat[17][31] ;
input \rst_dat[17][30] ;
input \rst_dat[17][29] ;
input \rst_dat[17][28] ;
input \rst_dat[17][27] ;
input \rst_dat[17][26] ;
input \rst_dat[17][25] ;
input \rst_dat[17][24] ;
input \rst_dat[17][23] ;
input \rst_dat[17][22] ;
input \rst_dat[17][21] ;
input \rst_dat[17][20] ;
input \rst_dat[17][19] ;
input \rst_dat[17][18] ;
input \rst_dat[17][17] ;
input \rst_dat[17][16] ;
input \rst_dat[17][15] ;
input \rst_dat[17][14] ;
input \rst_dat[17][13] ;
input \rst_dat[17][12] ;
input \rst_dat[17][11] ;
input \rst_dat[17][10] ;
input \rst_dat[17][9] ;
input \rst_dat[17][8] ;
input \rst_dat[17][7] ;
input \rst_dat[17][6] ;
input \rst_dat[17][5] ;
input \rst_dat[17][4] ;
input \rst_dat[17][3] ;
input \rst_dat[17][2] ;
input \rst_dat[17][1] ;
input \rst_dat[17][0] ;
input \rst_dat[18][31] ;
input \rst_dat[18][30] ;
input \rst_dat[18][29] ;
input \rst_dat[18][28] ;
input \rst_dat[18][27] ;
input \rst_dat[18][26] ;
input \rst_dat[18][25] ;
input \rst_dat[18][24] ;
input \rst_dat[18][23] ;
input \rst_dat[18][22] ;
input \rst_dat[18][21] ;
input \rst_dat[18][20] ;
input \rst_dat[18][19] ;
input \rst_dat[18][18] ;
input \rst_dat[18][17] ;
input \rst_dat[18][16] ;
input \rst_dat[18][15] ;
input \rst_dat[18][14] ;
input \rst_dat[18][13] ;
input \rst_dat[18][12] ;
input \rst_dat[18][11] ;
input \rst_dat[18][10] ;
input \rst_dat[18][9] ;
input \rst_dat[18][8] ;
input \rst_dat[18][7] ;
input \rst_dat[18][6] ;
input \rst_dat[18][5] ;
input \rst_dat[18][4] ;
input \rst_dat[18][3] ;
input \rst_dat[18][2] ;
input \rst_dat[18][1] ;
input \rst_dat[18][0] ;
input \rst_dat[19][31] ;
input \rst_dat[19][30] ;
input \rst_dat[19][29] ;
input \rst_dat[19][28] ;
input \rst_dat[19][27] ;
input \rst_dat[19][26] ;
input \rst_dat[19][25] ;
input \rst_dat[19][24] ;
input \rst_dat[19][23] ;
input \rst_dat[19][22] ;
input \rst_dat[19][21] ;
input \rst_dat[19][20] ;
input \rst_dat[19][19] ;
input \rst_dat[19][18] ;
input \rst_dat[19][17] ;
input \rst_dat[19][16] ;
input \rst_dat[19][15] ;
input \rst_dat[19][14] ;
input \rst_dat[19][13] ;
input \rst_dat[19][12] ;
input \rst_dat[19][11] ;
input \rst_dat[19][10] ;
input \rst_dat[19][9] ;
input \rst_dat[19][8] ;
input \rst_dat[19][7] ;
input \rst_dat[19][6] ;
input \rst_dat[19][5] ;
input \rst_dat[19][4] ;
input \rst_dat[19][3] ;
input \rst_dat[19][2] ;
input \rst_dat[19][1] ;
input \rst_dat[19][0] ;
input \rst_dat[20][31] ;
input \rst_dat[20][30] ;
input \rst_dat[20][29] ;
input \rst_dat[20][28] ;
input \rst_dat[20][27] ;
input \rst_dat[20][26] ;
input \rst_dat[20][25] ;
input \rst_dat[20][24] ;
input \rst_dat[20][23] ;
input \rst_dat[20][22] ;
input \rst_dat[20][21] ;
input \rst_dat[20][20] ;
input \rst_dat[20][19] ;
input \rst_dat[20][18] ;
input \rst_dat[20][17] ;
input \rst_dat[20][16] ;
input \rst_dat[20][15] ;
input \rst_dat[20][14] ;
input \rst_dat[20][13] ;
input \rst_dat[20][12] ;
input \rst_dat[20][11] ;
input \rst_dat[20][10] ;
input \rst_dat[20][9] ;
input \rst_dat[20][8] ;
input \rst_dat[20][7] ;
input \rst_dat[20][6] ;
input \rst_dat[20][5] ;
input \rst_dat[20][4] ;
input \rst_dat[20][3] ;
input \rst_dat[20][2] ;
input \rst_dat[20][1] ;
input \rst_dat[20][0] ;
input \rst_dat[21][31] ;
input \rst_dat[21][30] ;
input \rst_dat[21][29] ;
input \rst_dat[21][28] ;
input \rst_dat[21][27] ;
input \rst_dat[21][26] ;
input \rst_dat[21][25] ;
input \rst_dat[21][24] ;
input \rst_dat[21][23] ;
input \rst_dat[21][22] ;
input \rst_dat[21][21] ;
input \rst_dat[21][20] ;
input \rst_dat[21][19] ;
input \rst_dat[21][18] ;
input \rst_dat[21][17] ;
input \rst_dat[21][16] ;
input \rst_dat[21][15] ;
input \rst_dat[21][14] ;
input \rst_dat[21][13] ;
input \rst_dat[21][12] ;
input \rst_dat[21][11] ;
input \rst_dat[21][10] ;
input \rst_dat[21][9] ;
input \rst_dat[21][8] ;
input \rst_dat[21][7] ;
input \rst_dat[21][6] ;
input \rst_dat[21][5] ;
input \rst_dat[21][4] ;
input \rst_dat[21][3] ;
input \rst_dat[21][2] ;
input \rst_dat[21][1] ;
input \rst_dat[21][0] ;
input \rst_dat[22][31] ;
input \rst_dat[22][30] ;
input \rst_dat[22][29] ;
input \rst_dat[22][28] ;
input \rst_dat[22][27] ;
input \rst_dat[22][26] ;
input \rst_dat[22][25] ;
input \rst_dat[22][24] ;
input \rst_dat[22][23] ;
input \rst_dat[22][22] ;
input \rst_dat[22][21] ;
input \rst_dat[22][20] ;
input \rst_dat[22][19] ;
input \rst_dat[22][18] ;
input \rst_dat[22][17] ;
input \rst_dat[22][16] ;
input \rst_dat[22][15] ;
input \rst_dat[22][14] ;
input \rst_dat[22][13] ;
input \rst_dat[22][12] ;
input \rst_dat[22][11] ;
input \rst_dat[22][10] ;
input \rst_dat[22][9] ;
input \rst_dat[22][8] ;
input \rst_dat[22][7] ;
input \rst_dat[22][6] ;
input \rst_dat[22][5] ;
input \rst_dat[22][4] ;
input \rst_dat[22][3] ;
input \rst_dat[22][2] ;
input \rst_dat[22][1] ;
input \rst_dat[22][0] ;
input \rst_dat[23][31] ;
input \rst_dat[23][30] ;
input \rst_dat[23][29] ;
input \rst_dat[23][28] ;
input \rst_dat[23][27] ;
input \rst_dat[23][26] ;
input \rst_dat[23][25] ;
input \rst_dat[23][24] ;
input \rst_dat[23][23] ;
input \rst_dat[23][22] ;
input \rst_dat[23][21] ;
input \rst_dat[23][20] ;
input \rst_dat[23][19] ;
input \rst_dat[23][18] ;
input \rst_dat[23][17] ;
input \rst_dat[23][16] ;
input \rst_dat[23][15] ;
input \rst_dat[23][14] ;
input \rst_dat[23][13] ;
input \rst_dat[23][12] ;
input \rst_dat[23][11] ;
input \rst_dat[23][10] ;
input \rst_dat[23][9] ;
input \rst_dat[23][8] ;
input \rst_dat[23][7] ;
input \rst_dat[23][6] ;
input \rst_dat[23][5] ;
input \rst_dat[23][4] ;
input \rst_dat[23][3] ;
input \rst_dat[23][2] ;
input \rst_dat[23][1] ;
input \rst_dat[23][0] ;
input \rst_dat[24][31] ;
input \rst_dat[24][30] ;
input \rst_dat[24][29] ;
input \rst_dat[24][28] ;
input \rst_dat[24][27] ;
input \rst_dat[24][26] ;
input \rst_dat[24][25] ;
input \rst_dat[24][24] ;
input \rst_dat[24][23] ;
input \rst_dat[24][22] ;
input \rst_dat[24][21] ;
input \rst_dat[24][20] ;
input \rst_dat[24][19] ;
input \rst_dat[24][18] ;
input \rst_dat[24][17] ;
input \rst_dat[24][16] ;
input \rst_dat[24][15] ;
input \rst_dat[24][14] ;
input \rst_dat[24][13] ;
input \rst_dat[24][12] ;
input \rst_dat[24][11] ;
input \rst_dat[24][10] ;
input \rst_dat[24][9] ;
input \rst_dat[24][8] ;
input \rst_dat[24][7] ;
input \rst_dat[24][6] ;
input \rst_dat[24][5] ;
input \rst_dat[24][4] ;
input \rst_dat[24][3] ;
input \rst_dat[24][2] ;
input \rst_dat[24][1] ;
input \rst_dat[24][0] ;
input \rst_dat[25][31] ;
input \rst_dat[25][30] ;
input \rst_dat[25][29] ;
input \rst_dat[25][28] ;
input \rst_dat[25][27] ;
input \rst_dat[25][26] ;
input \rst_dat[25][25] ;
input \rst_dat[25][24] ;
input \rst_dat[25][23] ;
input \rst_dat[25][22] ;
input \rst_dat[25][21] ;
input \rst_dat[25][20] ;
input \rst_dat[25][19] ;
input \rst_dat[25][18] ;
input \rst_dat[25][17] ;
input \rst_dat[25][16] ;
input \rst_dat[25][15] ;
input \rst_dat[25][14] ;
input \rst_dat[25][13] ;
input \rst_dat[25][12] ;
input \rst_dat[25][11] ;
input \rst_dat[25][10] ;
input \rst_dat[25][9] ;
input \rst_dat[25][8] ;
input \rst_dat[25][7] ;
input \rst_dat[25][6] ;
input \rst_dat[25][5] ;
input \rst_dat[25][4] ;
input \rst_dat[25][3] ;
input \rst_dat[25][2] ;
input \rst_dat[25][1] ;
input \rst_dat[25][0] ;
input \rst_dat[26][31] ;
input \rst_dat[26][30] ;
input \rst_dat[26][29] ;
input \rst_dat[26][28] ;
input \rst_dat[26][27] ;
input \rst_dat[26][26] ;
input \rst_dat[26][25] ;
input \rst_dat[26][24] ;
input \rst_dat[26][23] ;
input \rst_dat[26][22] ;
input \rst_dat[26][21] ;
input \rst_dat[26][20] ;
input \rst_dat[26][19] ;
input \rst_dat[26][18] ;
input \rst_dat[26][17] ;
input \rst_dat[26][16] ;
input \rst_dat[26][15] ;
input \rst_dat[26][14] ;
input \rst_dat[26][13] ;
input \rst_dat[26][12] ;
input \rst_dat[26][11] ;
input \rst_dat[26][10] ;
input \rst_dat[26][9] ;
input \rst_dat[26][8] ;
input \rst_dat[26][7] ;
input \rst_dat[26][6] ;
input \rst_dat[26][5] ;
input \rst_dat[26][4] ;
input \rst_dat[26][3] ;
input \rst_dat[26][2] ;
input \rst_dat[26][1] ;
input \rst_dat[26][0] ;
input \rst_dat[27][31] ;
input \rst_dat[27][30] ;
input \rst_dat[27][29] ;
input \rst_dat[27][28] ;
input \rst_dat[27][27] ;
input \rst_dat[27][26] ;
input \rst_dat[27][25] ;
input \rst_dat[27][24] ;
input \rst_dat[27][23] ;
input \rst_dat[27][22] ;
input \rst_dat[27][21] ;
input \rst_dat[27][20] ;
input \rst_dat[27][19] ;
input \rst_dat[27][18] ;
input \rst_dat[27][17] ;
input \rst_dat[27][16] ;
input \rst_dat[27][15] ;
input \rst_dat[27][14] ;
input \rst_dat[27][13] ;
input \rst_dat[27][12] ;
input \rst_dat[27][11] ;
input \rst_dat[27][10] ;
input \rst_dat[27][9] ;
input \rst_dat[27][8] ;
input \rst_dat[27][7] ;
input \rst_dat[27][6] ;
input \rst_dat[27][5] ;
input \rst_dat[27][4] ;
input \rst_dat[27][3] ;
input \rst_dat[27][2] ;
input \rst_dat[27][1] ;
input \rst_dat[27][0] ;
input \rst_dat[28][31] ;
input \rst_dat[28][30] ;
input \rst_dat[28][29] ;
input \rst_dat[28][28] ;
input \rst_dat[28][27] ;
input \rst_dat[28][26] ;
input \rst_dat[28][25] ;
input \rst_dat[28][24] ;
input \rst_dat[28][23] ;
input \rst_dat[28][22] ;
input \rst_dat[28][21] ;
input \rst_dat[28][20] ;
input \rst_dat[28][19] ;
input \rst_dat[28][18] ;
input \rst_dat[28][17] ;
input \rst_dat[28][16] ;
input \rst_dat[28][15] ;
input \rst_dat[28][14] ;
input \rst_dat[28][13] ;
input \rst_dat[28][12] ;
input \rst_dat[28][11] ;
input \rst_dat[28][10] ;
input \rst_dat[28][9] ;
input \rst_dat[28][8] ;
input \rst_dat[28][7] ;
input \rst_dat[28][6] ;
input \rst_dat[28][5] ;
input \rst_dat[28][4] ;
input \rst_dat[28][3] ;
input \rst_dat[28][2] ;
input \rst_dat[28][1] ;
input \rst_dat[28][0] ;
input \rst_dat[29][31] ;
input \rst_dat[29][30] ;
input \rst_dat[29][29] ;
input \rst_dat[29][28] ;
input \rst_dat[29][27] ;
input \rst_dat[29][26] ;
input \rst_dat[29][25] ;
input \rst_dat[29][24] ;
input \rst_dat[29][23] ;
input \rst_dat[29][22] ;
input \rst_dat[29][21] ;
input \rst_dat[29][20] ;
input \rst_dat[29][19] ;
input \rst_dat[29][18] ;
input \rst_dat[29][17] ;
input \rst_dat[29][16] ;
input \rst_dat[29][15] ;
input \rst_dat[29][14] ;
input \rst_dat[29][13] ;
input \rst_dat[29][12] ;
input \rst_dat[29][11] ;
input \rst_dat[29][10] ;
input \rst_dat[29][9] ;
input \rst_dat[29][8] ;
input \rst_dat[29][7] ;
input \rst_dat[29][6] ;
input \rst_dat[29][5] ;
input \rst_dat[29][4] ;
input \rst_dat[29][3] ;
input \rst_dat[29][2] ;
input \rst_dat[29][1] ;
input \rst_dat[29][0] ;
input \rst_dat[30][31] ;
input \rst_dat[30][30] ;
input \rst_dat[30][29] ;
input \rst_dat[30][28] ;
input \rst_dat[30][27] ;
input \rst_dat[30][26] ;
input \rst_dat[30][25] ;
input \rst_dat[30][24] ;
input \rst_dat[30][23] ;
input \rst_dat[30][22] ;
input \rst_dat[30][21] ;
input \rst_dat[30][20] ;
input \rst_dat[30][19] ;
input \rst_dat[30][18] ;
input \rst_dat[30][17] ;
input \rst_dat[30][16] ;
input \rst_dat[30][15] ;
input \rst_dat[30][14] ;
input \rst_dat[30][13] ;
input \rst_dat[30][12] ;
input \rst_dat[30][11] ;
input \rst_dat[30][10] ;
input \rst_dat[30][9] ;
input \rst_dat[30][8] ;
input \rst_dat[30][7] ;
input \rst_dat[30][6] ;
input \rst_dat[30][5] ;
input \rst_dat[30][4] ;
input \rst_dat[30][3] ;
input \rst_dat[30][2] ;
input \rst_dat[30][1] ;
input \rst_dat[30][0] ;
input \rst_dat[31][31] ;
input \rst_dat[31][30] ;
input \rst_dat[31][29] ;
input \rst_dat[31][28] ;
input \rst_dat[31][27] ;
input \rst_dat[31][26] ;
input \rst_dat[31][25] ;
input \rst_dat[31][24] ;
input \rst_dat[31][23] ;
input \rst_dat[31][22] ;
input \rst_dat[31][21] ;
input \rst_dat[31][20] ;
input \rst_dat[31][19] ;
input \rst_dat[31][18] ;
input \rst_dat[31][17] ;
input \rst_dat[31][16] ;
input \rst_dat[31][15] ;
input \rst_dat[31][14] ;
input \rst_dat[31][13] ;
input \rst_dat[31][12] ;
input \rst_dat[31][11] ;
input \rst_dat[31][10] ;
input \rst_dat[31][9] ;
input \rst_dat[31][8] ;
input \rst_dat[31][7] ;
input \rst_dat[31][6] ;
input \rst_dat[31][5] ;
input \rst_dat[31][4] ;
input \rst_dat[31][3] ;
input \rst_dat[31][2] ;
input \rst_dat[31][1] ;
input \rst_dat[31][0] ;
wire [0:2] _zy_simnet_stat_code_0_w$;
wire [0:4] _zy_simnet_stat_datawords_1_w$;
wire [0:4] _zy_simnet_stat_addr_2_w$;
wire [0:15] _zy_simnet_capability_lst_3_w$;
wire [0:3] _zy_simnet_capability_type_4_w$;
wire [0:31] _zy_simnet_rd_dat_5_w$;
wire _zy_simnet_cio_6;
wire [0:2] _zy_simnet_stat_code_7_w$;
wire [0:4] _zy_simnet_stat_datawords_8_w$;
wire [0:4] _zy_simnet_stat_addr_9_w$;
wire _zy_simnet_dio_10;
wire [0:15] _zy_simnet_capability_lst_11_w$;
wire [0:3] _zy_simnet_capability_type_12_w$;
wire _zy_simnet_dio_13;
wire [0:4] _zy_simnet_addr_limit_14_w$;
wire [0:31] _zy_simnet_rd_dat_15_w$;
wire _zy_simnet_sw_cs_16_w$;
wire _zy_simnet_dio_17;
wire _zy_simnet_sw_we_18_w$;
wire [0:4] _zy_simnet_sw_add_19_w$;
wire [0:31] _zy_simnet_sw_wdat_20_w$;
wire [0:31] _zy_simnet_sw_rdat_21_w$;
wire _zy_simnet_cio_22;
wire [0:3] _zy_simnet_cio_23;
wire _zy_simnet_cio_24;
wire _zy_simnet_dio_25;
wire _zy_simnet_reset_26_w$;
wire [1023:0] _zyixc_ctx_wdata_1;
wire _zzM132L132_bcMevClk0;
wire _zzM132L132_bcReq0;
wire _zzM132L132_bcBusy0;
wire _zzM132L132_bcWait0;
wire _zz_zy_simnet_sw_cs_16_w$_M132_bcSv1;
wire _zz_zy_simnet_sw_we_18_w$_M132_bcSv2;
wire [0:4] _zz_zy_simnet_sw_add_19_w$_M132_bcSv3;
wire [0:31] _zz_zy_simnet_sw_wdat_20_w$_M132_bcSv4;
wire _zz_zy_simnet_reset_26_w$_M132_bcSv5;
wire _zzM132_bcBehEvalClk;
wire _zzM132_bcBehHalt;
wire reset;
wire [4:0] sw_add;
wire sw_cs;
wire [31:0] sw_wdat;
wire [31:0] sw_rdat;
wire sw_we;
wire [4:0] addr_limit;
wire [31:0] _zzM132_bcBehEval;
supply1 n1;
supply1 n5;
supply1 n6;
supply0 n7;
supply0 n8;
supply0 n9;
Q_BUF U0 ( .A(n1), .Z(_zy_simnet_cio_24));
Q_BUF U1 ( .A(n9), .Z(_zy_simnet_cio_23[3]));
Q_BUF U2 ( .A(n9), .Z(_zy_simnet_cio_23[2]));
Q_BUF U3 ( .A(n9), .Z(_zy_simnet_cio_23[1]));
Q_BUF U4 ( .A(n9), .Z(_zy_simnet_cio_23[0]));
Q_BUF U5 ( .A(n9), .Z(_zy_simnet_cio_22));
Q_BUF U6 ( .A(n9), .Z(_zy_simnet_cio_6));
Q_BUF U7 ( .A(n1), .Z(addr_limit[0]));
Q_BUF U8 ( .A(n1), .Z(addr_limit[1]));
Q_BUF U9 ( .A(n1), .Z(addr_limit[2]));
Q_BUF U10 ( .A(n1), .Z(addr_limit[3]));
Q_BUF U11 ( .A(n1), .Z(addr_limit[4]));
Q_BUF U12 ( .A(n9), .Z(n2));
Q_AN02 U13 ( .A0(n183), .A1(n184), .Z(n3));
nx_indirect_access_cntrl_xcm111 u_cntrl ( clk, rst_n, wr_stb, addr[10:0], 
	cmnd_op[3:0], cmnd_addr[4:0], _zy_simnet_cio_6, 
	_zy_simnet_stat_code_7_w$[0:2], _zy_simnet_stat_datawords_8_w$[0:4], 
	_zy_simnet_stat_addr_9_w$[0:4], _zy_simnet_dio_10, 
	_zy_simnet_capability_lst_11_w$[0:15], 
	_zy_simnet_capability_type_12_w$[0:3], _zy_simnet_dio_13, 
	_zy_simnet_addr_limit_14_w$[0:4], wr_dat[31:0], 
	_zy_simnet_rd_dat_15_w$[0:31], _zy_simnet_sw_cs_16_w$, 
	_zy_simnet_dio_17, _zy_simnet_sw_we_18_w$, 
	_zy_simnet_sw_add_19_w$[0:4], _zy_simnet_sw_wdat_20_w$[0:31], 
	_zy_simnet_sw_rdat_21_w$[0:31], _zy_simnet_cio_22, 
	_zy_simnet_cio_23[0:3], _zy_simnet_cio_24, _zy_simnet_dio_25, 
	_zy_simnet_reset_26_w$);
ixc_capLoopXp _zzM132L34_bcBehEvalP0 ( _zzM132_bcBehEvalClk, n2,, 
	_zzM132_bcBehHalt);
ixc_sample_logic _zz_zy_simnet_reset_26_w$_M132_bcSp5 ( 
	_zz_zy_simnet_reset_26_w$_M132_bcSv5, _zy_simnet_reset_26_w$);
ixc_sample_logic_32 _zz_zy_simnet_sw_wdat_20_w$_M132_bcSp4 ( 
	_zz_zy_simnet_sw_wdat_20_w$_M132_bcSv4[0:31], 
	_zy_simnet_sw_wdat_20_w$[0:31]);
ixc_sample_logic_5 _zz_zy_simnet_sw_add_19_w$_M132_bcSp3 ( 
	_zz_zy_simnet_sw_add_19_w$_M132_bcSv3[0:4], 
	_zy_simnet_sw_add_19_w$[0:4]);
ixc_sample_logic _zz_zy_simnet_sw_we_18_w$_M132_bcSp2 ( 
	_zz_zy_simnet_sw_we_18_w$_M132_bcSv2, _zy_simnet_sw_we_18_w$);
ixc_sample_logic _zz_zy_simnet_sw_cs_16_w$_M132_bcSp1 ( 
	_zz_zy_simnet_sw_cs_16_w$_M132_bcSv1, _zy_simnet_sw_cs_16_w$);
ixc_mevClk_2_0_0_3_1_0_1 _zzM132L132_bcMevClkP0 ( _zzM132L132_bcMevClk0, { 
	clk, rst_n}, { n5, n6}, n7, n8, _zzM132L132_bcReq0, 
	_zzM132L132_bcBusy0, _zzM132L132_bcWait0);
ixc_context_write_1024 _zzixc_ctxwr_1 ( { \mem_a[0][31] , \mem_a[0][30] , 
	\mem_a[0][29] , \mem_a[0][28] , \mem_a[0][27] , \mem_a[0][26] , 
	\mem_a[0][25] , \mem_a[0][24] , \mem_a[0][23] , \mem_a[0][22] , 
	\mem_a[0][21] , \mem_a[0][20] , \mem_a[0][19] , \mem_a[0][18] , 
	\mem_a[0][17] , \mem_a[0][16] , \mem_a[0][15] , \mem_a[0][14] , 
	\mem_a[0][13] , \mem_a[0][12] , \mem_a[0][11] , \mem_a[0][10] , 
	\mem_a[0][9] , \mem_a[0][8] , \mem_a[0][7] , \mem_a[0][6] , 
	\mem_a[0][5] , \mem_a[0][4] , \mem_a[0][3] , \mem_a[0][2] , 
	\mem_a[0][1] , \mem_a[0][0] , \mem_a[1][31] , \mem_a[1][30] , 
	\mem_a[1][29] , \mem_a[1][28] , \mem_a[1][27] , \mem_a[1][26] , 
	\mem_a[1][25] , \mem_a[1][24] , \mem_a[1][23] , \mem_a[1][22] , 
	\mem_a[1][21] , \mem_a[1][20] , \mem_a[1][19] , \mem_a[1][18] , 
	\mem_a[1][17] , \mem_a[1][16] , \mem_a[1][15] , \mem_a[1][14] , 
	\mem_a[1][13] , \mem_a[1][12] , \mem_a[1][11] , \mem_a[1][10] , 
	\mem_a[1][9] , \mem_a[1][8] , \mem_a[1][7] , \mem_a[1][6] , 
	\mem_a[1][5] , \mem_a[1][4] , \mem_a[1][3] , \mem_a[1][2] , 
	\mem_a[1][1] , \mem_a[1][0] , \mem_a[2][31] , \mem_a[2][30] , 
	\mem_a[2][29] , \mem_a[2][28] , \mem_a[2][27] , \mem_a[2][26] , 
	\mem_a[2][25] , \mem_a[2][24] , \mem_a[2][23] , \mem_a[2][22] , 
	\mem_a[2][21] , \mem_a[2][20] , \mem_a[2][19] , \mem_a[2][18] , 
	\mem_a[2][17] , \mem_a[2][16] , \mem_a[2][15] , \mem_a[2][14] , 
	\mem_a[2][13] , \mem_a[2][12] , \mem_a[2][11] , \mem_a[2][10] , 
	\mem_a[2][9] , \mem_a[2][8] , \mem_a[2][7] , \mem_a[2][6] , 
	\mem_a[2][5] , \mem_a[2][4] , \mem_a[2][3] , \mem_a[2][2] , 
	\mem_a[2][1] , \mem_a[2][0] , \mem_a[3][31] , \mem_a[3][30] , 
	\mem_a[3][29] , \mem_a[3][28] , \mem_a[3][27] , \mem_a[3][26] , 
	\mem_a[3][25] , \mem_a[3][24] , \mem_a[3][23] , \mem_a[3][22] , 
	\mem_a[3][21] , \mem_a[3][20] , \mem_a[3][19] , \mem_a[3][18] , 
	\mem_a[3][17] , \mem_a[3][16] , \mem_a[3][15] , \mem_a[3][14] , 
	\mem_a[3][13] , \mem_a[3][12] , \mem_a[3][11] , \mem_a[3][10] , 
	\mem_a[3][9] , \mem_a[3][8] , \mem_a[3][7] , \mem_a[3][6] , 
	\mem_a[3][5] , \mem_a[3][4] , \mem_a[3][3] , \mem_a[3][2] , 
	\mem_a[3][1] , \mem_a[3][0] , \mem_a[4][31] , \mem_a[4][30] , 
	\mem_a[4][29] , \mem_a[4][28] , \mem_a[4][27] , \mem_a[4][26] , 
	\mem_a[4][25] , \mem_a[4][24] , \mem_a[4][23] , \mem_a[4][22] , 
	\mem_a[4][21] , \mem_a[4][20] , \mem_a[4][19] , \mem_a[4][18] , 
	\mem_a[4][17] , \mem_a[4][16] , \mem_a[4][15] , \mem_a[4][14] , 
	\mem_a[4][13] , \mem_a[4][12] , \mem_a[4][11] , \mem_a[4][10] , 
	\mem_a[4][9] , \mem_a[4][8] , \mem_a[4][7] , \mem_a[4][6] , 
	\mem_a[4][5] , \mem_a[4][4] , \mem_a[4][3] , \mem_a[4][2] , 
	\mem_a[4][1] , \mem_a[4][0] , \mem_a[5][31] , \mem_a[5][30] , 
	\mem_a[5][29] , \mem_a[5][28] , \mem_a[5][27] , \mem_a[5][26] , 
	\mem_a[5][25] , \mem_a[5][24] , \mem_a[5][23] , \mem_a[5][22] , 
	\mem_a[5][21] , \mem_a[5][20] , \mem_a[5][19] , \mem_a[5][18] , 
	\mem_a[5][17] , \mem_a[5][16] , \mem_a[5][15] , \mem_a[5][14] , 
	\mem_a[5][13] , \mem_a[5][12] , \mem_a[5][11] , \mem_a[5][10] , 
	\mem_a[5][9] , \mem_a[5][8] , \mem_a[5][7] , \mem_a[5][6] , 
	\mem_a[5][5] , \mem_a[5][4] , \mem_a[5][3] , \mem_a[5][2] , 
	\mem_a[5][1] , \mem_a[5][0] , \mem_a[6][31] , \mem_a[6][30] , 
	\mem_a[6][29] , \mem_a[6][28] , \mem_a[6][27] , \mem_a[6][26] , 
	\mem_a[6][25] , \mem_a[6][24] , \mem_a[6][23] , \mem_a[6][22] , 
	\mem_a[6][21] , \mem_a[6][20] , \mem_a[6][19] , \mem_a[6][18] , 
	\mem_a[6][17] , \mem_a[6][16] , \mem_a[6][15] , \mem_a[6][14] , 
	\mem_a[6][13] , \mem_a[6][12] , \mem_a[6][11] , \mem_a[6][10] , 
	\mem_a[6][9] , \mem_a[6][8] , \mem_a[6][7] , \mem_a[6][6] , 
	\mem_a[6][5] , \mem_a[6][4] , \mem_a[6][3] , \mem_a[6][2] , 
	\mem_a[6][1] , \mem_a[6][0] , \mem_a[7][31] , \mem_a[7][30] , 
	\mem_a[7][29] , \mem_a[7][28] , \mem_a[7][27] , \mem_a[7][26] , 
	\mem_a[7][25] , \mem_a[7][24] , \mem_a[7][23] , \mem_a[7][22] , 
	\mem_a[7][21] , \mem_a[7][20] , \mem_a[7][19] , \mem_a[7][18] , 
	\mem_a[7][17] , \mem_a[7][16] , \mem_a[7][15] , \mem_a[7][14] , 
	\mem_a[7][13] , \mem_a[7][12] , \mem_a[7][11] , \mem_a[7][10] , 
	\mem_a[7][9] , \mem_a[7][8] , \mem_a[7][7] , \mem_a[7][6] , 
	\mem_a[7][5] , \mem_a[7][4] , \mem_a[7][3] , \mem_a[7][2] , 
	\mem_a[7][1] , \mem_a[7][0] , \mem_a[8][31] , \mem_a[8][30] , 
	\mem_a[8][29] , \mem_a[8][28] , \mem_a[8][27] , \mem_a[8][26] , 
	\mem_a[8][25] , \mem_a[8][24] , \mem_a[8][23] , \mem_a[8][22] , 
	\mem_a[8][21] , \mem_a[8][20] , \mem_a[8][19] , \mem_a[8][18] , 
	\mem_a[8][17] , \mem_a[8][16] , \mem_a[8][15] , \mem_a[8][14] , 
	\mem_a[8][13] , \mem_a[8][12] , \mem_a[8][11] , \mem_a[8][10] , 
	\mem_a[8][9] , \mem_a[8][8] , \mem_a[8][7] , \mem_a[8][6] , 
	\mem_a[8][5] , \mem_a[8][4] , \mem_a[8][3] , \mem_a[8][2] , 
	\mem_a[8][1] , \mem_a[8][0] , \mem_a[9][31] , \mem_a[9][30] , 
	\mem_a[9][29] , \mem_a[9][28] , \mem_a[9][27] , \mem_a[9][26] , 
	\mem_a[9][25] , \mem_a[9][24] , \mem_a[9][23] , \mem_a[9][22] , 
	\mem_a[9][21] , \mem_a[9][20] , \mem_a[9][19] , \mem_a[9][18] , 
	\mem_a[9][17] , \mem_a[9][16] , \mem_a[9][15] , \mem_a[9][14] , 
	\mem_a[9][13] , \mem_a[9][12] , \mem_a[9][11] , \mem_a[9][10] , 
	\mem_a[9][9] , \mem_a[9][8] , \mem_a[9][7] , \mem_a[9][6] , 
	\mem_a[9][5] , \mem_a[9][4] , \mem_a[9][3] , \mem_a[9][2] , 
	\mem_a[9][1] , \mem_a[9][0] , \mem_a[10][31] , \mem_a[10][30] , 
	\mem_a[10][29] , \mem_a[10][28] , \mem_a[10][27] , \mem_a[10][26] , 
	\mem_a[10][25] , \mem_a[10][24] , \mem_a[10][23] , \mem_a[10][22] , 
	\mem_a[10][21] , \mem_a[10][20] , \mem_a[10][19] , \mem_a[10][18] , 
	\mem_a[10][17] , \mem_a[10][16] , \mem_a[10][15] , \mem_a[10][14] , 
	\mem_a[10][13] , \mem_a[10][12] , \mem_a[10][11] , \mem_a[10][10] , 
	\mem_a[10][9] , \mem_a[10][8] , \mem_a[10][7] , \mem_a[10][6] , 
	\mem_a[10][5] , \mem_a[10][4] , \mem_a[10][3] , \mem_a[10][2] , 
	\mem_a[10][1] , \mem_a[10][0] , \mem_a[11][31] , \mem_a[11][30] , 
	\mem_a[11][29] , \mem_a[11][28] , \mem_a[11][27] , \mem_a[11][26] , 
	\mem_a[11][25] , \mem_a[11][24] , \mem_a[11][23] , \mem_a[11][22] , 
	\mem_a[11][21] , \mem_a[11][20] , \mem_a[11][19] , \mem_a[11][18] , 
	\mem_a[11][17] , \mem_a[11][16] , \mem_a[11][15] , \mem_a[11][14] , 
	\mem_a[11][13] , \mem_a[11][12] , \mem_a[11][11] , \mem_a[11][10] , 
	\mem_a[11][9] , \mem_a[11][8] , \mem_a[11][7] , \mem_a[11][6] , 
	\mem_a[11][5] , \mem_a[11][4] , \mem_a[11][3] , \mem_a[11][2] , 
	\mem_a[11][1] , \mem_a[11][0] , \mem_a[12][31] , \mem_a[12][30] , 
	\mem_a[12][29] , \mem_a[12][28] , \mem_a[12][27] , \mem_a[12][26] , 
	\mem_a[12][25] , \mem_a[12][24] , \mem_a[12][23] , \mem_a[12][22] , 
	\mem_a[12][21] , \mem_a[12][20] , \mem_a[12][19] , \mem_a[12][18] , 
	\mem_a[12][17] , \mem_a[12][16] , \mem_a[12][15] , \mem_a[12][14] , 
	\mem_a[12][13] , \mem_a[12][12] , \mem_a[12][11] , \mem_a[12][10] , 
	\mem_a[12][9] , \mem_a[12][8] , \mem_a[12][7] , \mem_a[12][6] , 
	\mem_a[12][5] , \mem_a[12][4] , \mem_a[12][3] , \mem_a[12][2] , 
	\mem_a[12][1] , \mem_a[12][0] , \mem_a[13][31] , \mem_a[13][30] , 
	\mem_a[13][29] , \mem_a[13][28] , \mem_a[13][27] , \mem_a[13][26] , 
	\mem_a[13][25] , \mem_a[13][24] , \mem_a[13][23] , \mem_a[13][22] , 
	\mem_a[13][21] , \mem_a[13][20] , \mem_a[13][19] , \mem_a[13][18] , 
	\mem_a[13][17] , \mem_a[13][16] , \mem_a[13][15] , \mem_a[13][14] , 
	\mem_a[13][13] , \mem_a[13][12] , \mem_a[13][11] , \mem_a[13][10] , 
	\mem_a[13][9] , \mem_a[13][8] , \mem_a[13][7] , \mem_a[13][6] , 
	\mem_a[13][5] , \mem_a[13][4] , \mem_a[13][3] , \mem_a[13][2] , 
	\mem_a[13][1] , \mem_a[13][0] , \mem_a[14][31] , \mem_a[14][30] , 
	\mem_a[14][29] , \mem_a[14][28] , \mem_a[14][27] , \mem_a[14][26] , 
	\mem_a[14][25] , \mem_a[14][24] , \mem_a[14][23] , \mem_a[14][22] , 
	\mem_a[14][21] , \mem_a[14][20] , \mem_a[14][19] , \mem_a[14][18] , 
	\mem_a[14][17] , \mem_a[14][16] , \mem_a[14][15] , \mem_a[14][14] , 
	\mem_a[14][13] , \mem_a[14][12] , \mem_a[14][11] , \mem_a[14][10] , 
	\mem_a[14][9] , \mem_a[14][8] , \mem_a[14][7] , \mem_a[14][6] , 
	\mem_a[14][5] , \mem_a[14][4] , \mem_a[14][3] , \mem_a[14][2] , 
	\mem_a[14][1] , \mem_a[14][0] , \mem_a[15][31] , \mem_a[15][30] , 
	\mem_a[15][29] , \mem_a[15][28] , \mem_a[15][27] , \mem_a[15][26] , 
	\mem_a[15][25] , \mem_a[15][24] , \mem_a[15][23] , \mem_a[15][22] , 
	\mem_a[15][21] , \mem_a[15][20] , \mem_a[15][19] , \mem_a[15][18] , 
	\mem_a[15][17] , \mem_a[15][16] , \mem_a[15][15] , \mem_a[15][14] , 
	\mem_a[15][13] , \mem_a[15][12] , \mem_a[15][11] , \mem_a[15][10] , 
	\mem_a[15][9] , \mem_a[15][8] , \mem_a[15][7] , \mem_a[15][6] , 
	\mem_a[15][5] , \mem_a[15][4] , \mem_a[15][3] , \mem_a[15][2] , 
	\mem_a[15][1] , \mem_a[15][0] , \mem_a[16][31] , \mem_a[16][30] , 
	\mem_a[16][29] , \mem_a[16][28] , \mem_a[16][27] , \mem_a[16][26] , 
	\mem_a[16][25] , \mem_a[16][24] , \mem_a[16][23] , \mem_a[16][22] , 
	\mem_a[16][21] , \mem_a[16][20] , \mem_a[16][19] , \mem_a[16][18] , 
	\mem_a[16][17] , \mem_a[16][16] , \mem_a[16][15] , \mem_a[16][14] , 
	\mem_a[16][13] , \mem_a[16][12] , \mem_a[16][11] , \mem_a[16][10] , 
	\mem_a[16][9] , \mem_a[16][8] , \mem_a[16][7] , \mem_a[16][6] , 
	\mem_a[16][5] , \mem_a[16][4] , \mem_a[16][3] , \mem_a[16][2] , 
	\mem_a[16][1] , \mem_a[16][0] , \mem_a[17][31] , \mem_a[17][30] , 
	\mem_a[17][29] , \mem_a[17][28] , \mem_a[17][27] , \mem_a[17][26] , 
	\mem_a[17][25] , \mem_a[17][24] , \mem_a[17][23] , \mem_a[17][22] , 
	\mem_a[17][21] , \mem_a[17][20] , \mem_a[17][19] , \mem_a[17][18] , 
	\mem_a[17][17] , \mem_a[17][16] , \mem_a[17][15] , \mem_a[17][14] , 
	\mem_a[17][13] , \mem_a[17][12] , \mem_a[17][11] , \mem_a[17][10] , 
	\mem_a[17][9] , \mem_a[17][8] , \mem_a[17][7] , \mem_a[17][6] , 
	\mem_a[17][5] , \mem_a[17][4] , \mem_a[17][3] , \mem_a[17][2] , 
	\mem_a[17][1] , \mem_a[17][0] , \mem_a[18][31] , \mem_a[18][30] , 
	\mem_a[18][29] , \mem_a[18][28] , \mem_a[18][27] , \mem_a[18][26] , 
	\mem_a[18][25] , \mem_a[18][24] , \mem_a[18][23] , \mem_a[18][22] , 
	\mem_a[18][21] , \mem_a[18][20] , \mem_a[18][19] , \mem_a[18][18] , 
	\mem_a[18][17] , \mem_a[18][16] , \mem_a[18][15] , \mem_a[18][14] , 
	\mem_a[18][13] , \mem_a[18][12] , \mem_a[18][11] , \mem_a[18][10] , 
	\mem_a[18][9] , \mem_a[18][8] , \mem_a[18][7] , \mem_a[18][6] , 
	\mem_a[18][5] , \mem_a[18][4] , \mem_a[18][3] , \mem_a[18][2] , 
	\mem_a[18][1] , \mem_a[18][0] , \mem_a[19][31] , \mem_a[19][30] , 
	\mem_a[19][29] , \mem_a[19][28] , \mem_a[19][27] , \mem_a[19][26] , 
	\mem_a[19][25] , \mem_a[19][24] , \mem_a[19][23] , \mem_a[19][22] , 
	\mem_a[19][21] , \mem_a[19][20] , \mem_a[19][19] , \mem_a[19][18] , 
	\mem_a[19][17] , \mem_a[19][16] , \mem_a[19][15] , \mem_a[19][14] , 
	\mem_a[19][13] , \mem_a[19][12] , \mem_a[19][11] , \mem_a[19][10] , 
	\mem_a[19][9] , \mem_a[19][8] , \mem_a[19][7] , \mem_a[19][6] , 
	\mem_a[19][5] , \mem_a[19][4] , \mem_a[19][3] , \mem_a[19][2] , 
	\mem_a[19][1] , \mem_a[19][0] , \mem_a[20][31] , \mem_a[20][30] , 
	\mem_a[20][29] , \mem_a[20][28] , \mem_a[20][27] , \mem_a[20][26] , 
	\mem_a[20][25] , \mem_a[20][24] , \mem_a[20][23] , \mem_a[20][22] , 
	\mem_a[20][21] , \mem_a[20][20] , \mem_a[20][19] , \mem_a[20][18] , 
	\mem_a[20][17] , \mem_a[20][16] , \mem_a[20][15] , \mem_a[20][14] , 
	\mem_a[20][13] , \mem_a[20][12] , \mem_a[20][11] , \mem_a[20][10] , 
	\mem_a[20][9] , \mem_a[20][8] , \mem_a[20][7] , \mem_a[20][6] , 
	\mem_a[20][5] , \mem_a[20][4] , \mem_a[20][3] , \mem_a[20][2] , 
	\mem_a[20][1] , \mem_a[20][0] , \mem_a[21][31] , \mem_a[21][30] , 
	\mem_a[21][29] , \mem_a[21][28] , \mem_a[21][27] , \mem_a[21][26] , 
	\mem_a[21][25] , \mem_a[21][24] , \mem_a[21][23] , \mem_a[21][22] , 
	\mem_a[21][21] , \mem_a[21][20] , \mem_a[21][19] , \mem_a[21][18] , 
	\mem_a[21][17] , \mem_a[21][16] , \mem_a[21][15] , \mem_a[21][14] , 
	\mem_a[21][13] , \mem_a[21][12] , \mem_a[21][11] , \mem_a[21][10] , 
	\mem_a[21][9] , \mem_a[21][8] , \mem_a[21][7] , \mem_a[21][6] , 
	\mem_a[21][5] , \mem_a[21][4] , \mem_a[21][3] , \mem_a[21][2] , 
	\mem_a[21][1] , \mem_a[21][0] , \mem_a[22][31] , \mem_a[22][30] , 
	\mem_a[22][29] , \mem_a[22][28] , \mem_a[22][27] , \mem_a[22][26] , 
	\mem_a[22][25] , \mem_a[22][24] , \mem_a[22][23] , \mem_a[22][22] , 
	\mem_a[22][21] , \mem_a[22][20] , \mem_a[22][19] , \mem_a[22][18] , 
	\mem_a[22][17] , \mem_a[22][16] , \mem_a[22][15] , \mem_a[22][14] , 
	\mem_a[22][13] , \mem_a[22][12] , \mem_a[22][11] , \mem_a[22][10] , 
	\mem_a[22][9] , \mem_a[22][8] , \mem_a[22][7] , \mem_a[22][6] , 
	\mem_a[22][5] , \mem_a[22][4] , \mem_a[22][3] , \mem_a[22][2] , 
	\mem_a[22][1] , \mem_a[22][0] , \mem_a[23][31] , \mem_a[23][30] , 
	\mem_a[23][29] , \mem_a[23][28] , \mem_a[23][27] , \mem_a[23][26] , 
	\mem_a[23][25] , \mem_a[23][24] , \mem_a[23][23] , \mem_a[23][22] , 
	\mem_a[23][21] , \mem_a[23][20] , \mem_a[23][19] , \mem_a[23][18] , 
	\mem_a[23][17] , \mem_a[23][16] , \mem_a[23][15] , \mem_a[23][14] , 
	\mem_a[23][13] , \mem_a[23][12] , \mem_a[23][11] , \mem_a[23][10] , 
	\mem_a[23][9] , \mem_a[23][8] , \mem_a[23][7] , \mem_a[23][6] , 
	\mem_a[23][5] , \mem_a[23][4] , \mem_a[23][3] , \mem_a[23][2] , 
	\mem_a[23][1] , \mem_a[23][0] , \mem_a[24][31] , \mem_a[24][30] , 
	\mem_a[24][29] , \mem_a[24][28] , \mem_a[24][27] , \mem_a[24][26] , 
	\mem_a[24][25] , \mem_a[24][24] , \mem_a[24][23] , \mem_a[24][22] , 
	\mem_a[24][21] , \mem_a[24][20] , \mem_a[24][19] , \mem_a[24][18] , 
	\mem_a[24][17] , \mem_a[24][16] , \mem_a[24][15] , \mem_a[24][14] , 
	\mem_a[24][13] , \mem_a[24][12] , \mem_a[24][11] , \mem_a[24][10] , 
	\mem_a[24][9] , \mem_a[24][8] , \mem_a[24][7] , \mem_a[24][6] , 
	\mem_a[24][5] , \mem_a[24][4] , \mem_a[24][3] , \mem_a[24][2] , 
	\mem_a[24][1] , \mem_a[24][0] , \mem_a[25][31] , \mem_a[25][30] , 
	\mem_a[25][29] , \mem_a[25][28] , \mem_a[25][27] , \mem_a[25][26] , 
	\mem_a[25][25] , \mem_a[25][24] , \mem_a[25][23] , \mem_a[25][22] , 
	\mem_a[25][21] , \mem_a[25][20] , \mem_a[25][19] , \mem_a[25][18] , 
	\mem_a[25][17] , \mem_a[25][16] , \mem_a[25][15] , \mem_a[25][14] , 
	\mem_a[25][13] , \mem_a[25][12] , \mem_a[25][11] , \mem_a[25][10] , 
	\mem_a[25][9] , \mem_a[25][8] , \mem_a[25][7] , \mem_a[25][6] , 
	\mem_a[25][5] , \mem_a[25][4] , \mem_a[25][3] , \mem_a[25][2] , 
	\mem_a[25][1] , \mem_a[25][0] , \mem_a[26][31] , \mem_a[26][30] , 
	\mem_a[26][29] , \mem_a[26][28] , \mem_a[26][27] , \mem_a[26][26] , 
	\mem_a[26][25] , \mem_a[26][24] , \mem_a[26][23] , \mem_a[26][22] , 
	\mem_a[26][21] , \mem_a[26][20] , \mem_a[26][19] , \mem_a[26][18] , 
	\mem_a[26][17] , \mem_a[26][16] , \mem_a[26][15] , \mem_a[26][14] , 
	\mem_a[26][13] , \mem_a[26][12] , \mem_a[26][11] , \mem_a[26][10] , 
	\mem_a[26][9] , \mem_a[26][8] , \mem_a[26][7] , \mem_a[26][6] , 
	\mem_a[26][5] , \mem_a[26][4] , \mem_a[26][3] , \mem_a[26][2] , 
	\mem_a[26][1] , \mem_a[26][0] , \mem_a[27][31] , \mem_a[27][30] , 
	\mem_a[27][29] , \mem_a[27][28] , \mem_a[27][27] , \mem_a[27][26] , 
	\mem_a[27][25] , \mem_a[27][24] , \mem_a[27][23] , \mem_a[27][22] , 
	\mem_a[27][21] , \mem_a[27][20] , \mem_a[27][19] , \mem_a[27][18] , 
	\mem_a[27][17] , \mem_a[27][16] , \mem_a[27][15] , \mem_a[27][14] , 
	\mem_a[27][13] , \mem_a[27][12] , \mem_a[27][11] , \mem_a[27][10] , 
	\mem_a[27][9] , \mem_a[27][8] , \mem_a[27][7] , \mem_a[27][6] , 
	\mem_a[27][5] , \mem_a[27][4] , \mem_a[27][3] , \mem_a[27][2] , 
	\mem_a[27][1] , \mem_a[27][0] , \mem_a[28][31] , \mem_a[28][30] , 
	\mem_a[28][29] , \mem_a[28][28] , \mem_a[28][27] , \mem_a[28][26] , 
	\mem_a[28][25] , \mem_a[28][24] , \mem_a[28][23] , \mem_a[28][22] , 
	\mem_a[28][21] , \mem_a[28][20] , \mem_a[28][19] , \mem_a[28][18] , 
	\mem_a[28][17] , \mem_a[28][16] , \mem_a[28][15] , \mem_a[28][14] , 
	\mem_a[28][13] , \mem_a[28][12] , \mem_a[28][11] , \mem_a[28][10] , 
	\mem_a[28][9] , \mem_a[28][8] , \mem_a[28][7] , \mem_a[28][6] , 
	\mem_a[28][5] , \mem_a[28][4] , \mem_a[28][3] , \mem_a[28][2] , 
	\mem_a[28][1] , \mem_a[28][0] , \mem_a[29][31] , \mem_a[29][30] , 
	\mem_a[29][29] , \mem_a[29][28] , \mem_a[29][27] , \mem_a[29][26] , 
	\mem_a[29][25] , \mem_a[29][24] , \mem_a[29][23] , \mem_a[29][22] , 
	\mem_a[29][21] , \mem_a[29][20] , \mem_a[29][19] , \mem_a[29][18] , 
	\mem_a[29][17] , \mem_a[29][16] , \mem_a[29][15] , \mem_a[29][14] , 
	\mem_a[29][13] , \mem_a[29][12] , \mem_a[29][11] , \mem_a[29][10] , 
	\mem_a[29][9] , \mem_a[29][8] , \mem_a[29][7] , \mem_a[29][6] , 
	\mem_a[29][5] , \mem_a[29][4] , \mem_a[29][3] , \mem_a[29][2] , 
	\mem_a[29][1] , \mem_a[29][0] , \mem_a[30][31] , \mem_a[30][30] , 
	\mem_a[30][29] , \mem_a[30][28] , \mem_a[30][27] , \mem_a[30][26] , 
	\mem_a[30][25] , \mem_a[30][24] , \mem_a[30][23] , \mem_a[30][22] , 
	\mem_a[30][21] , \mem_a[30][20] , \mem_a[30][19] , \mem_a[30][18] , 
	\mem_a[30][17] , \mem_a[30][16] , \mem_a[30][15] , \mem_a[30][14] , 
	\mem_a[30][13] , \mem_a[30][12] , \mem_a[30][11] , \mem_a[30][10] , 
	\mem_a[30][9] , \mem_a[30][8] , \mem_a[30][7] , \mem_a[30][6] , 
	\mem_a[30][5] , \mem_a[30][4] , \mem_a[30][3] , \mem_a[30][2] , 
	\mem_a[30][1] , \mem_a[30][0] , \mem_a[31][31] , \mem_a[31][30] , 
	\mem_a[31][29] , \mem_a[31][28] , \mem_a[31][27] , \mem_a[31][26] , 
	\mem_a[31][25] , \mem_a[31][24] , \mem_a[31][23] , \mem_a[31][22] , 
	\mem_a[31][21] , \mem_a[31][20] , \mem_a[31][19] , \mem_a[31][18] , 
	\mem_a[31][17] , \mem_a[31][16] , \mem_a[31][15] , \mem_a[31][14] , 
	\mem_a[31][13] , \mem_a[31][12] , \mem_a[31][11] , \mem_a[31][10] , 
	\mem_a[31][9] , \mem_a[31][8] , \mem_a[31][7] , \mem_a[31][6] , 
	\mem_a[31][5] , \mem_a[31][4] , \mem_a[31][3] , \mem_a[31][2] , 
	\mem_a[31][1] , \mem_a[31][0] });
ixc_context_read_1024 _zzixc_ctxrd_0 ( { \mem_a[0][31] , \mem_a[0][30] , 
	\mem_a[0][29] , \mem_a[0][28] , \mem_a[0][27] , \mem_a[0][26] , 
	\mem_a[0][25] , \mem_a[0][24] , \mem_a[0][23] , \mem_a[0][22] , 
	\mem_a[0][21] , \mem_a[0][20] , \mem_a[0][19] , \mem_a[0][18] , 
	\mem_a[0][17] , \mem_a[0][16] , \mem_a[0][15] , \mem_a[0][14] , 
	\mem_a[0][13] , \mem_a[0][12] , \mem_a[0][11] , \mem_a[0][10] , 
	\mem_a[0][9] , \mem_a[0][8] , \mem_a[0][7] , \mem_a[0][6] , 
	\mem_a[0][5] , \mem_a[0][4] , \mem_a[0][3] , \mem_a[0][2] , 
	\mem_a[0][1] , \mem_a[0][0] , \mem_a[1][31] , \mem_a[1][30] , 
	\mem_a[1][29] , \mem_a[1][28] , \mem_a[1][27] , \mem_a[1][26] , 
	\mem_a[1][25] , \mem_a[1][24] , \mem_a[1][23] , \mem_a[1][22] , 
	\mem_a[1][21] , \mem_a[1][20] , \mem_a[1][19] , \mem_a[1][18] , 
	\mem_a[1][17] , \mem_a[1][16] , \mem_a[1][15] , \mem_a[1][14] , 
	\mem_a[1][13] , \mem_a[1][12] , \mem_a[1][11] , \mem_a[1][10] , 
	\mem_a[1][9] , \mem_a[1][8] , \mem_a[1][7] , \mem_a[1][6] , 
	\mem_a[1][5] , \mem_a[1][4] , \mem_a[1][3] , \mem_a[1][2] , 
	\mem_a[1][1] , \mem_a[1][0] , \mem_a[2][31] , \mem_a[2][30] , 
	\mem_a[2][29] , \mem_a[2][28] , \mem_a[2][27] , \mem_a[2][26] , 
	\mem_a[2][25] , \mem_a[2][24] , \mem_a[2][23] , \mem_a[2][22] , 
	\mem_a[2][21] , \mem_a[2][20] , \mem_a[2][19] , \mem_a[2][18] , 
	\mem_a[2][17] , \mem_a[2][16] , \mem_a[2][15] , \mem_a[2][14] , 
	\mem_a[2][13] , \mem_a[2][12] , \mem_a[2][11] , \mem_a[2][10] , 
	\mem_a[2][9] , \mem_a[2][8] , \mem_a[2][7] , \mem_a[2][6] , 
	\mem_a[2][5] , \mem_a[2][4] , \mem_a[2][3] , \mem_a[2][2] , 
	\mem_a[2][1] , \mem_a[2][0] , \mem_a[3][31] , \mem_a[3][30] , 
	\mem_a[3][29] , \mem_a[3][28] , \mem_a[3][27] , \mem_a[3][26] , 
	\mem_a[3][25] , \mem_a[3][24] , \mem_a[3][23] , \mem_a[3][22] , 
	\mem_a[3][21] , \mem_a[3][20] , \mem_a[3][19] , \mem_a[3][18] , 
	\mem_a[3][17] , \mem_a[3][16] , \mem_a[3][15] , \mem_a[3][14] , 
	\mem_a[3][13] , \mem_a[3][12] , \mem_a[3][11] , \mem_a[3][10] , 
	\mem_a[3][9] , \mem_a[3][8] , \mem_a[3][7] , \mem_a[3][6] , 
	\mem_a[3][5] , \mem_a[3][4] , \mem_a[3][3] , \mem_a[3][2] , 
	\mem_a[3][1] , \mem_a[3][0] , \mem_a[4][31] , \mem_a[4][30] , 
	\mem_a[4][29] , \mem_a[4][28] , \mem_a[4][27] , \mem_a[4][26] , 
	\mem_a[4][25] , \mem_a[4][24] , \mem_a[4][23] , \mem_a[4][22] , 
	\mem_a[4][21] , \mem_a[4][20] , \mem_a[4][19] , \mem_a[4][18] , 
	\mem_a[4][17] , \mem_a[4][16] , \mem_a[4][15] , \mem_a[4][14] , 
	\mem_a[4][13] , \mem_a[4][12] , \mem_a[4][11] , \mem_a[4][10] , 
	\mem_a[4][9] , \mem_a[4][8] , \mem_a[4][7] , \mem_a[4][6] , 
	\mem_a[4][5] , \mem_a[4][4] , \mem_a[4][3] , \mem_a[4][2] , 
	\mem_a[4][1] , \mem_a[4][0] , \mem_a[5][31] , \mem_a[5][30] , 
	\mem_a[5][29] , \mem_a[5][28] , \mem_a[5][27] , \mem_a[5][26] , 
	\mem_a[5][25] , \mem_a[5][24] , \mem_a[5][23] , \mem_a[5][22] , 
	\mem_a[5][21] , \mem_a[5][20] , \mem_a[5][19] , \mem_a[5][18] , 
	\mem_a[5][17] , \mem_a[5][16] , \mem_a[5][15] , \mem_a[5][14] , 
	\mem_a[5][13] , \mem_a[5][12] , \mem_a[5][11] , \mem_a[5][10] , 
	\mem_a[5][9] , \mem_a[5][8] , \mem_a[5][7] , \mem_a[5][6] , 
	\mem_a[5][5] , \mem_a[5][4] , \mem_a[5][3] , \mem_a[5][2] , 
	\mem_a[5][1] , \mem_a[5][0] , \mem_a[6][31] , \mem_a[6][30] , 
	\mem_a[6][29] , \mem_a[6][28] , \mem_a[6][27] , \mem_a[6][26] , 
	\mem_a[6][25] , \mem_a[6][24] , \mem_a[6][23] , \mem_a[6][22] , 
	\mem_a[6][21] , \mem_a[6][20] , \mem_a[6][19] , \mem_a[6][18] , 
	\mem_a[6][17] , \mem_a[6][16] , \mem_a[6][15] , \mem_a[6][14] , 
	\mem_a[6][13] , \mem_a[6][12] , \mem_a[6][11] , \mem_a[6][10] , 
	\mem_a[6][9] , \mem_a[6][8] , \mem_a[6][7] , \mem_a[6][6] , 
	\mem_a[6][5] , \mem_a[6][4] , \mem_a[6][3] , \mem_a[6][2] , 
	\mem_a[6][1] , \mem_a[6][0] , \mem_a[7][31] , \mem_a[7][30] , 
	\mem_a[7][29] , \mem_a[7][28] , \mem_a[7][27] , \mem_a[7][26] , 
	\mem_a[7][25] , \mem_a[7][24] , \mem_a[7][23] , \mem_a[7][22] , 
	\mem_a[7][21] , \mem_a[7][20] , \mem_a[7][19] , \mem_a[7][18] , 
	\mem_a[7][17] , \mem_a[7][16] , \mem_a[7][15] , \mem_a[7][14] , 
	\mem_a[7][13] , \mem_a[7][12] , \mem_a[7][11] , \mem_a[7][10] , 
	\mem_a[7][9] , \mem_a[7][8] , \mem_a[7][7] , \mem_a[7][6] , 
	\mem_a[7][5] , \mem_a[7][4] , \mem_a[7][3] , \mem_a[7][2] , 
	\mem_a[7][1] , \mem_a[7][0] , \mem_a[8][31] , \mem_a[8][30] , 
	\mem_a[8][29] , \mem_a[8][28] , \mem_a[8][27] , \mem_a[8][26] , 
	\mem_a[8][25] , \mem_a[8][24] , \mem_a[8][23] , \mem_a[8][22] , 
	\mem_a[8][21] , \mem_a[8][20] , \mem_a[8][19] , \mem_a[8][18] , 
	\mem_a[8][17] , \mem_a[8][16] , \mem_a[8][15] , \mem_a[8][14] , 
	\mem_a[8][13] , \mem_a[8][12] , \mem_a[8][11] , \mem_a[8][10] , 
	\mem_a[8][9] , \mem_a[8][8] , \mem_a[8][7] , \mem_a[8][6] , 
	\mem_a[8][5] , \mem_a[8][4] , \mem_a[8][3] , \mem_a[8][2] , 
	\mem_a[8][1] , \mem_a[8][0] , \mem_a[9][31] , \mem_a[9][30] , 
	\mem_a[9][29] , \mem_a[9][28] , \mem_a[9][27] , \mem_a[9][26] , 
	\mem_a[9][25] , \mem_a[9][24] , \mem_a[9][23] , \mem_a[9][22] , 
	\mem_a[9][21] , \mem_a[9][20] , \mem_a[9][19] , \mem_a[9][18] , 
	\mem_a[9][17] , \mem_a[9][16] , \mem_a[9][15] , \mem_a[9][14] , 
	\mem_a[9][13] , \mem_a[9][12] , \mem_a[9][11] , \mem_a[9][10] , 
	\mem_a[9][9] , \mem_a[9][8] , \mem_a[9][7] , \mem_a[9][6] , 
	\mem_a[9][5] , \mem_a[9][4] , \mem_a[9][3] , \mem_a[9][2] , 
	\mem_a[9][1] , \mem_a[9][0] , \mem_a[10][31] , \mem_a[10][30] , 
	\mem_a[10][29] , \mem_a[10][28] , \mem_a[10][27] , \mem_a[10][26] , 
	\mem_a[10][25] , \mem_a[10][24] , \mem_a[10][23] , \mem_a[10][22] , 
	\mem_a[10][21] , \mem_a[10][20] , \mem_a[10][19] , \mem_a[10][18] , 
	\mem_a[10][17] , \mem_a[10][16] , \mem_a[10][15] , \mem_a[10][14] , 
	\mem_a[10][13] , \mem_a[10][12] , \mem_a[10][11] , \mem_a[10][10] , 
	\mem_a[10][9] , \mem_a[10][8] , \mem_a[10][7] , \mem_a[10][6] , 
	\mem_a[10][5] , \mem_a[10][4] , \mem_a[10][3] , \mem_a[10][2] , 
	\mem_a[10][1] , \mem_a[10][0] , \mem_a[11][31] , \mem_a[11][30] , 
	\mem_a[11][29] , \mem_a[11][28] , \mem_a[11][27] , \mem_a[11][26] , 
	\mem_a[11][25] , \mem_a[11][24] , \mem_a[11][23] , \mem_a[11][22] , 
	\mem_a[11][21] , \mem_a[11][20] , \mem_a[11][19] , \mem_a[11][18] , 
	\mem_a[11][17] , \mem_a[11][16] , \mem_a[11][15] , \mem_a[11][14] , 
	\mem_a[11][13] , \mem_a[11][12] , \mem_a[11][11] , \mem_a[11][10] , 
	\mem_a[11][9] , \mem_a[11][8] , \mem_a[11][7] , \mem_a[11][6] , 
	\mem_a[11][5] , \mem_a[11][4] , \mem_a[11][3] , \mem_a[11][2] , 
	\mem_a[11][1] , \mem_a[11][0] , \mem_a[12][31] , \mem_a[12][30] , 
	\mem_a[12][29] , \mem_a[12][28] , \mem_a[12][27] , \mem_a[12][26] , 
	\mem_a[12][25] , \mem_a[12][24] , \mem_a[12][23] , \mem_a[12][22] , 
	\mem_a[12][21] , \mem_a[12][20] , \mem_a[12][19] , \mem_a[12][18] , 
	\mem_a[12][17] , \mem_a[12][16] , \mem_a[12][15] , \mem_a[12][14] , 
	\mem_a[12][13] , \mem_a[12][12] , \mem_a[12][11] , \mem_a[12][10] , 
	\mem_a[12][9] , \mem_a[12][8] , \mem_a[12][7] , \mem_a[12][6] , 
	\mem_a[12][5] , \mem_a[12][4] , \mem_a[12][3] , \mem_a[12][2] , 
	\mem_a[12][1] , \mem_a[12][0] , \mem_a[13][31] , \mem_a[13][30] , 
	\mem_a[13][29] , \mem_a[13][28] , \mem_a[13][27] , \mem_a[13][26] , 
	\mem_a[13][25] , \mem_a[13][24] , \mem_a[13][23] , \mem_a[13][22] , 
	\mem_a[13][21] , \mem_a[13][20] , \mem_a[13][19] , \mem_a[13][18] , 
	\mem_a[13][17] , \mem_a[13][16] , \mem_a[13][15] , \mem_a[13][14] , 
	\mem_a[13][13] , \mem_a[13][12] , \mem_a[13][11] , \mem_a[13][10] , 
	\mem_a[13][9] , \mem_a[13][8] , \mem_a[13][7] , \mem_a[13][6] , 
	\mem_a[13][5] , \mem_a[13][4] , \mem_a[13][3] , \mem_a[13][2] , 
	\mem_a[13][1] , \mem_a[13][0] , \mem_a[14][31] , \mem_a[14][30] , 
	\mem_a[14][29] , \mem_a[14][28] , \mem_a[14][27] , \mem_a[14][26] , 
	\mem_a[14][25] , \mem_a[14][24] , \mem_a[14][23] , \mem_a[14][22] , 
	\mem_a[14][21] , \mem_a[14][20] , \mem_a[14][19] , \mem_a[14][18] , 
	\mem_a[14][17] , \mem_a[14][16] , \mem_a[14][15] , \mem_a[14][14] , 
	\mem_a[14][13] , \mem_a[14][12] , \mem_a[14][11] , \mem_a[14][10] , 
	\mem_a[14][9] , \mem_a[14][8] , \mem_a[14][7] , \mem_a[14][6] , 
	\mem_a[14][5] , \mem_a[14][4] , \mem_a[14][3] , \mem_a[14][2] , 
	\mem_a[14][1] , \mem_a[14][0] , \mem_a[15][31] , \mem_a[15][30] , 
	\mem_a[15][29] , \mem_a[15][28] , \mem_a[15][27] , \mem_a[15][26] , 
	\mem_a[15][25] , \mem_a[15][24] , \mem_a[15][23] , \mem_a[15][22] , 
	\mem_a[15][21] , \mem_a[15][20] , \mem_a[15][19] , \mem_a[15][18] , 
	\mem_a[15][17] , \mem_a[15][16] , \mem_a[15][15] , \mem_a[15][14] , 
	\mem_a[15][13] , \mem_a[15][12] , \mem_a[15][11] , \mem_a[15][10] , 
	\mem_a[15][9] , \mem_a[15][8] , \mem_a[15][7] , \mem_a[15][6] , 
	\mem_a[15][5] , \mem_a[15][4] , \mem_a[15][3] , \mem_a[15][2] , 
	\mem_a[15][1] , \mem_a[15][0] , \mem_a[16][31] , \mem_a[16][30] , 
	\mem_a[16][29] , \mem_a[16][28] , \mem_a[16][27] , \mem_a[16][26] , 
	\mem_a[16][25] , \mem_a[16][24] , \mem_a[16][23] , \mem_a[16][22] , 
	\mem_a[16][21] , \mem_a[16][20] , \mem_a[16][19] , \mem_a[16][18] , 
	\mem_a[16][17] , \mem_a[16][16] , \mem_a[16][15] , \mem_a[16][14] , 
	\mem_a[16][13] , \mem_a[16][12] , \mem_a[16][11] , \mem_a[16][10] , 
	\mem_a[16][9] , \mem_a[16][8] , \mem_a[16][7] , \mem_a[16][6] , 
	\mem_a[16][5] , \mem_a[16][4] , \mem_a[16][3] , \mem_a[16][2] , 
	\mem_a[16][1] , \mem_a[16][0] , \mem_a[17][31] , \mem_a[17][30] , 
	\mem_a[17][29] , \mem_a[17][28] , \mem_a[17][27] , \mem_a[17][26] , 
	\mem_a[17][25] , \mem_a[17][24] , \mem_a[17][23] , \mem_a[17][22] , 
	\mem_a[17][21] , \mem_a[17][20] , \mem_a[17][19] , \mem_a[17][18] , 
	\mem_a[17][17] , \mem_a[17][16] , \mem_a[17][15] , \mem_a[17][14] , 
	\mem_a[17][13] , \mem_a[17][12] , \mem_a[17][11] , \mem_a[17][10] , 
	\mem_a[17][9] , \mem_a[17][8] , \mem_a[17][7] , \mem_a[17][6] , 
	\mem_a[17][5] , \mem_a[17][4] , \mem_a[17][3] , \mem_a[17][2] , 
	\mem_a[17][1] , \mem_a[17][0] , \mem_a[18][31] , \mem_a[18][30] , 
	\mem_a[18][29] , \mem_a[18][28] , \mem_a[18][27] , \mem_a[18][26] , 
	\mem_a[18][25] , \mem_a[18][24] , \mem_a[18][23] , \mem_a[18][22] , 
	\mem_a[18][21] , \mem_a[18][20] , \mem_a[18][19] , \mem_a[18][18] , 
	\mem_a[18][17] , \mem_a[18][16] , \mem_a[18][15] , \mem_a[18][14] , 
	\mem_a[18][13] , \mem_a[18][12] , \mem_a[18][11] , \mem_a[18][10] , 
	\mem_a[18][9] , \mem_a[18][8] , \mem_a[18][7] , \mem_a[18][6] , 
	\mem_a[18][5] , \mem_a[18][4] , \mem_a[18][3] , \mem_a[18][2] , 
	\mem_a[18][1] , \mem_a[18][0] , \mem_a[19][31] , \mem_a[19][30] , 
	\mem_a[19][29] , \mem_a[19][28] , \mem_a[19][27] , \mem_a[19][26] , 
	\mem_a[19][25] , \mem_a[19][24] , \mem_a[19][23] , \mem_a[19][22] , 
	\mem_a[19][21] , \mem_a[19][20] , \mem_a[19][19] , \mem_a[19][18] , 
	\mem_a[19][17] , \mem_a[19][16] , \mem_a[19][15] , \mem_a[19][14] , 
	\mem_a[19][13] , \mem_a[19][12] , \mem_a[19][11] , \mem_a[19][10] , 
	\mem_a[19][9] , \mem_a[19][8] , \mem_a[19][7] , \mem_a[19][6] , 
	\mem_a[19][5] , \mem_a[19][4] , \mem_a[19][3] , \mem_a[19][2] , 
	\mem_a[19][1] , \mem_a[19][0] , \mem_a[20][31] , \mem_a[20][30] , 
	\mem_a[20][29] , \mem_a[20][28] , \mem_a[20][27] , \mem_a[20][26] , 
	\mem_a[20][25] , \mem_a[20][24] , \mem_a[20][23] , \mem_a[20][22] , 
	\mem_a[20][21] , \mem_a[20][20] , \mem_a[20][19] , \mem_a[20][18] , 
	\mem_a[20][17] , \mem_a[20][16] , \mem_a[20][15] , \mem_a[20][14] , 
	\mem_a[20][13] , \mem_a[20][12] , \mem_a[20][11] , \mem_a[20][10] , 
	\mem_a[20][9] , \mem_a[20][8] , \mem_a[20][7] , \mem_a[20][6] , 
	\mem_a[20][5] , \mem_a[20][4] , \mem_a[20][3] , \mem_a[20][2] , 
	\mem_a[20][1] , \mem_a[20][0] , \mem_a[21][31] , \mem_a[21][30] , 
	\mem_a[21][29] , \mem_a[21][28] , \mem_a[21][27] , \mem_a[21][26] , 
	\mem_a[21][25] , \mem_a[21][24] , \mem_a[21][23] , \mem_a[21][22] , 
	\mem_a[21][21] , \mem_a[21][20] , \mem_a[21][19] , \mem_a[21][18] , 
	\mem_a[21][17] , \mem_a[21][16] , \mem_a[21][15] , \mem_a[21][14] , 
	\mem_a[21][13] , \mem_a[21][12] , \mem_a[21][11] , \mem_a[21][10] , 
	\mem_a[21][9] , \mem_a[21][8] , \mem_a[21][7] , \mem_a[21][6] , 
	\mem_a[21][5] , \mem_a[21][4] , \mem_a[21][3] , \mem_a[21][2] , 
	\mem_a[21][1] , \mem_a[21][0] , \mem_a[22][31] , \mem_a[22][30] , 
	\mem_a[22][29] , \mem_a[22][28] , \mem_a[22][27] , \mem_a[22][26] , 
	\mem_a[22][25] , \mem_a[22][24] , \mem_a[22][23] , \mem_a[22][22] , 
	\mem_a[22][21] , \mem_a[22][20] , \mem_a[22][19] , \mem_a[22][18] , 
	\mem_a[22][17] , \mem_a[22][16] , \mem_a[22][15] , \mem_a[22][14] , 
	\mem_a[22][13] , \mem_a[22][12] , \mem_a[22][11] , \mem_a[22][10] , 
	\mem_a[22][9] , \mem_a[22][8] , \mem_a[22][7] , \mem_a[22][6] , 
	\mem_a[22][5] , \mem_a[22][4] , \mem_a[22][3] , \mem_a[22][2] , 
	\mem_a[22][1] , \mem_a[22][0] , \mem_a[23][31] , \mem_a[23][30] , 
	\mem_a[23][29] , \mem_a[23][28] , \mem_a[23][27] , \mem_a[23][26] , 
	\mem_a[23][25] , \mem_a[23][24] , \mem_a[23][23] , \mem_a[23][22] , 
	\mem_a[23][21] , \mem_a[23][20] , \mem_a[23][19] , \mem_a[23][18] , 
	\mem_a[23][17] , \mem_a[23][16] , \mem_a[23][15] , \mem_a[23][14] , 
	\mem_a[23][13] , \mem_a[23][12] , \mem_a[23][11] , \mem_a[23][10] , 
	\mem_a[23][9] , \mem_a[23][8] , \mem_a[23][7] , \mem_a[23][6] , 
	\mem_a[23][5] , \mem_a[23][4] , \mem_a[23][3] , \mem_a[23][2] , 
	\mem_a[23][1] , \mem_a[23][0] , \mem_a[24][31] , \mem_a[24][30] , 
	\mem_a[24][29] , \mem_a[24][28] , \mem_a[24][27] , \mem_a[24][26] , 
	\mem_a[24][25] , \mem_a[24][24] , \mem_a[24][23] , \mem_a[24][22] , 
	\mem_a[24][21] , \mem_a[24][20] , \mem_a[24][19] , \mem_a[24][18] , 
	\mem_a[24][17] , \mem_a[24][16] , \mem_a[24][15] , \mem_a[24][14] , 
	\mem_a[24][13] , \mem_a[24][12] , \mem_a[24][11] , \mem_a[24][10] , 
	\mem_a[24][9] , \mem_a[24][8] , \mem_a[24][7] , \mem_a[24][6] , 
	\mem_a[24][5] , \mem_a[24][4] , \mem_a[24][3] , \mem_a[24][2] , 
	\mem_a[24][1] , \mem_a[24][0] , \mem_a[25][31] , \mem_a[25][30] , 
	\mem_a[25][29] , \mem_a[25][28] , \mem_a[25][27] , \mem_a[25][26] , 
	\mem_a[25][25] , \mem_a[25][24] , \mem_a[25][23] , \mem_a[25][22] , 
	\mem_a[25][21] , \mem_a[25][20] , \mem_a[25][19] , \mem_a[25][18] , 
	\mem_a[25][17] , \mem_a[25][16] , \mem_a[25][15] , \mem_a[25][14] , 
	\mem_a[25][13] , \mem_a[25][12] , \mem_a[25][11] , \mem_a[25][10] , 
	\mem_a[25][9] , \mem_a[25][8] , \mem_a[25][7] , \mem_a[25][6] , 
	\mem_a[25][5] , \mem_a[25][4] , \mem_a[25][3] , \mem_a[25][2] , 
	\mem_a[25][1] , \mem_a[25][0] , \mem_a[26][31] , \mem_a[26][30] , 
	\mem_a[26][29] , \mem_a[26][28] , \mem_a[26][27] , \mem_a[26][26] , 
	\mem_a[26][25] , \mem_a[26][24] , \mem_a[26][23] , \mem_a[26][22] , 
	\mem_a[26][21] , \mem_a[26][20] , \mem_a[26][19] , \mem_a[26][18] , 
	\mem_a[26][17] , \mem_a[26][16] , \mem_a[26][15] , \mem_a[26][14] , 
	\mem_a[26][13] , \mem_a[26][12] , \mem_a[26][11] , \mem_a[26][10] , 
	\mem_a[26][9] , \mem_a[26][8] , \mem_a[26][7] , \mem_a[26][6] , 
	\mem_a[26][5] , \mem_a[26][4] , \mem_a[26][3] , \mem_a[26][2] , 
	\mem_a[26][1] , \mem_a[26][0] , \mem_a[27][31] , \mem_a[27][30] , 
	\mem_a[27][29] , \mem_a[27][28] , \mem_a[27][27] , \mem_a[27][26] , 
	\mem_a[27][25] , \mem_a[27][24] , \mem_a[27][23] , \mem_a[27][22] , 
	\mem_a[27][21] , \mem_a[27][20] , \mem_a[27][19] , \mem_a[27][18] , 
	\mem_a[27][17] , \mem_a[27][16] , \mem_a[27][15] , \mem_a[27][14] , 
	\mem_a[27][13] , \mem_a[27][12] , \mem_a[27][11] , \mem_a[27][10] , 
	\mem_a[27][9] , \mem_a[27][8] , \mem_a[27][7] , \mem_a[27][6] , 
	\mem_a[27][5] , \mem_a[27][4] , \mem_a[27][3] , \mem_a[27][2] , 
	\mem_a[27][1] , \mem_a[27][0] , \mem_a[28][31] , \mem_a[28][30] , 
	\mem_a[28][29] , \mem_a[28][28] , \mem_a[28][27] , \mem_a[28][26] , 
	\mem_a[28][25] , \mem_a[28][24] , \mem_a[28][23] , \mem_a[28][22] , 
	\mem_a[28][21] , \mem_a[28][20] , \mem_a[28][19] , \mem_a[28][18] , 
	\mem_a[28][17] , \mem_a[28][16] , \mem_a[28][15] , \mem_a[28][14] , 
	\mem_a[28][13] , \mem_a[28][12] , \mem_a[28][11] , \mem_a[28][10] , 
	\mem_a[28][9] , \mem_a[28][8] , \mem_a[28][7] , \mem_a[28][6] , 
	\mem_a[28][5] , \mem_a[28][4] , \mem_a[28][3] , \mem_a[28][2] , 
	\mem_a[28][1] , \mem_a[28][0] , \mem_a[29][31] , \mem_a[29][30] , 
	\mem_a[29][29] , \mem_a[29][28] , \mem_a[29][27] , \mem_a[29][26] , 
	\mem_a[29][25] , \mem_a[29][24] , \mem_a[29][23] , \mem_a[29][22] , 
	\mem_a[29][21] , \mem_a[29][20] , \mem_a[29][19] , \mem_a[29][18] , 
	\mem_a[29][17] , \mem_a[29][16] , \mem_a[29][15] , \mem_a[29][14] , 
	\mem_a[29][13] , \mem_a[29][12] , \mem_a[29][11] , \mem_a[29][10] , 
	\mem_a[29][9] , \mem_a[29][8] , \mem_a[29][7] , \mem_a[29][6] , 
	\mem_a[29][5] , \mem_a[29][4] , \mem_a[29][3] , \mem_a[29][2] , 
	\mem_a[29][1] , \mem_a[29][0] , \mem_a[30][31] , \mem_a[30][30] , 
	\mem_a[30][29] , \mem_a[30][28] , \mem_a[30][27] , \mem_a[30][26] , 
	\mem_a[30][25] , \mem_a[30][24] , \mem_a[30][23] , \mem_a[30][22] , 
	\mem_a[30][21] , \mem_a[30][20] , \mem_a[30][19] , \mem_a[30][18] , 
	\mem_a[30][17] , \mem_a[30][16] , \mem_a[30][15] , \mem_a[30][14] , 
	\mem_a[30][13] , \mem_a[30][12] , \mem_a[30][11] , \mem_a[30][10] , 
	\mem_a[30][9] , \mem_a[30][8] , \mem_a[30][7] , \mem_a[30][6] , 
	\mem_a[30][5] , \mem_a[30][4] , \mem_a[30][3] , \mem_a[30][2] , 
	\mem_a[30][1] , \mem_a[30][0] , \mem_a[31][31] , \mem_a[31][30] , 
	\mem_a[31][29] , \mem_a[31][28] , \mem_a[31][27] , \mem_a[31][26] , 
	\mem_a[31][25] , \mem_a[31][24] , \mem_a[31][23] , \mem_a[31][22] , 
	\mem_a[31][21] , \mem_a[31][20] , \mem_a[31][19] , \mem_a[31][18] , 
	\mem_a[31][17] , \mem_a[31][16] , \mem_a[31][15] , \mem_a[31][14] , 
	\mem_a[31][13] , \mem_a[31][12] , \mem_a[31][11] , \mem_a[31][10] , 
	\mem_a[31][9] , \mem_a[31][8] , \mem_a[31][7] , \mem_a[31][6] , 
	\mem_a[31][5] , \mem_a[31][4] , \mem_a[31][3] , \mem_a[31][2] , 
	\mem_a[31][1] , \mem_a[31][0] });
ixc_assign _zz_strnp_18 ( reset, _zz_zy_simnet_reset_26_w$_M132_bcSv5);
ixc_assign_32 _zz_strnp_17 ( _zy_simnet_sw_rdat_21_w$[0:31], sw_rdat[31:0]);
ixc_assign_32 _zz_strnp_16 ( sw_wdat[31:0], 
	_zz_zy_simnet_sw_wdat_20_w$_M132_bcSv4[0:31]);
ixc_assign_5 _zz_strnp_15 ( sw_add[4:0], 
	_zz_zy_simnet_sw_add_19_w$_M132_bcSv3[0:4]);
ixc_assign _zz_strnp_14 ( sw_we, _zz_zy_simnet_sw_we_18_w$_M132_bcSv2);
ixc_assign _zz_strnp_13 ( sw_cs, _zz_zy_simnet_sw_cs_16_w$_M132_bcSv1);
ixc_assign_32 _zz_strnp_12 ( rd_dat[31:0], _zy_simnet_rd_dat_15_w$[0:31]);
ixc_assign_5 _zz_strnp_11 ( _zy_simnet_addr_limit_14_w$[0:4], addr_limit[4:0]);
ixc_assign_4 _zz_strnp_10 ( capability_type[3:0], 
	_zy_simnet_capability_type_12_w$[0:3]);
ixc_assign_16 _zz_strnp_9 ( capability_lst[15:0], 
	_zy_simnet_capability_lst_11_w$[0:15]);
ixc_assign_5 _zz_strnp_8 ( stat_addr[4:0], _zy_simnet_stat_addr_9_w$[0:4]);
ixc_assign_5 _zz_strnp_7 ( stat_datawords[4:0], 
	_zy_simnet_stat_datawords_8_w$[0:4]);
ixc_assign_3 _zz_strnp_6 ( stat_code[2:0], _zy_simnet_stat_code_7_w$[0:2]);
ixc_assign_32 _zz_strnp_5 ( _zy_simnet_rd_dat_5_w$[0:31], rd_dat[31:0]);
ixc_assign_4 _zz_strnp_4 ( _zy_simnet_capability_type_4_w$[0:3], 
	capability_type[3:0]);
ixc_assign_16 _zz_strnp_3 ( _zy_simnet_capability_lst_3_w$[0:15], 
	capability_lst[15:0]);
ixc_assign_5 _zz_strnp_2 ( _zy_simnet_stat_addr_2_w$[0:4], stat_addr[4:0]);
ixc_assign_5 _zz_strnp_1 ( _zy_simnet_stat_datawords_1_w$[0:4], 
	stat_datawords[4:0]);
ixc_assign_3 _zz_strnp_0 ( _zy_simnet_stat_code_0_w$[0:2], stat_code[2:0]);
Q_NOT_TOUCH _zzqnt ( .sig());
Q_AN03 U44 ( .A0(n45), .A1(sw_add[0]), .A2(n42), .Z(n185));
Q_AN03 U45 ( .A0(n45), .A1(sw_add[1]), .A2(n42), .Z(n186));
Q_AN03 U46 ( .A0(n45), .A1(sw_add[2]), .A2(n42), .Z(n187));
Q_AN03 U47 ( .A0(n45), .A1(sw_add[3]), .A2(n42), .Z(n188));
Q_AN03 U48 ( .A0(n45), .A1(sw_add[4]), .A2(n42), .Z(n189));
Q_MX02 U49 ( .S(n45), .A0(\rst_dat[0][0] ), .A1(sw_wdat[0]), .Z(n10));
Q_MX02 U50 ( .S(n45), .A0(\rst_dat[0][1] ), .A1(sw_wdat[1]), .Z(n11));
Q_MX02 U51 ( .S(n45), .A0(\rst_dat[0][2] ), .A1(sw_wdat[2]), .Z(n12));
Q_MX02 U52 ( .S(n45), .A0(\rst_dat[0][3] ), .A1(sw_wdat[3]), .Z(n13));
Q_MX02 U53 ( .S(n45), .A0(\rst_dat[0][4] ), .A1(sw_wdat[4]), .Z(n14));
Q_MX02 U54 ( .S(n45), .A0(\rst_dat[0][5] ), .A1(sw_wdat[5]), .Z(n15));
Q_MX02 U55 ( .S(n45), .A0(\rst_dat[0][6] ), .A1(sw_wdat[6]), .Z(n16));
Q_MX02 U56 ( .S(n45), .A0(\rst_dat[0][7] ), .A1(sw_wdat[7]), .Z(n17));
Q_MX02 U57 ( .S(n45), .A0(\rst_dat[0][8] ), .A1(sw_wdat[8]), .Z(n18));
Q_MX02 U58 ( .S(n45), .A0(\rst_dat[0][9] ), .A1(sw_wdat[9]), .Z(n19));
Q_MX02 U59 ( .S(n45), .A0(\rst_dat[0][10] ), .A1(sw_wdat[10]), .Z(n20));
Q_MX02 U60 ( .S(n45), .A0(\rst_dat[0][11] ), .A1(sw_wdat[11]), .Z(n21));
Q_MX02 U61 ( .S(n45), .A0(\rst_dat[0][12] ), .A1(sw_wdat[12]), .Z(n22));
Q_MX02 U62 ( .S(n45), .A0(\rst_dat[0][13] ), .A1(sw_wdat[13]), .Z(n23));
Q_MX02 U63 ( .S(n45), .A0(\rst_dat[0][14] ), .A1(sw_wdat[14]), .Z(n24));
Q_MX02 U64 ( .S(n45), .A0(\rst_dat[0][15] ), .A1(sw_wdat[15]), .Z(n25));
Q_MX02 U65 ( .S(n45), .A0(\rst_dat[0][16] ), .A1(sw_wdat[16]), .Z(n26));
Q_MX02 U66 ( .S(n45), .A0(\rst_dat[0][17] ), .A1(sw_wdat[17]), .Z(n27));
Q_MX02 U67 ( .S(n45), .A0(\rst_dat[0][18] ), .A1(sw_wdat[18]), .Z(n28));
Q_MX02 U68 ( .S(n45), .A0(\rst_dat[0][19] ), .A1(sw_wdat[19]), .Z(n29));
Q_MX02 U69 ( .S(n45), .A0(\rst_dat[0][20] ), .A1(sw_wdat[20]), .Z(n30));
Q_MX02 U70 ( .S(n45), .A0(\rst_dat[0][21] ), .A1(sw_wdat[21]), .Z(n31));
Q_MX02 U71 ( .S(n45), .A0(\rst_dat[0][22] ), .A1(sw_wdat[22]), .Z(n32));
Q_MX02 U72 ( .S(n45), .A0(\rst_dat[0][23] ), .A1(sw_wdat[23]), .Z(n33));
Q_MX02 U73 ( .S(n45), .A0(\rst_dat[0][24] ), .A1(sw_wdat[24]), .Z(n34));
Q_MX02 U74 ( .S(n45), .A0(\rst_dat[0][25] ), .A1(sw_wdat[25]), .Z(n35));
Q_MX02 U75 ( .S(n45), .A0(\rst_dat[0][26] ), .A1(sw_wdat[26]), .Z(n36));
Q_MX02 U76 ( .S(n45), .A0(\rst_dat[0][27] ), .A1(sw_wdat[27]), .Z(n37));
Q_MX02 U77 ( .S(n45), .A0(\rst_dat[0][28] ), .A1(sw_wdat[28]), .Z(n38));
Q_MX02 U78 ( .S(n45), .A0(\rst_dat[0][29] ), .A1(sw_wdat[29]), .Z(n39));
Q_MX02 U79 ( .S(n45), .A0(\rst_dat[0][30] ), .A1(sw_wdat[30]), .Z(n40));
Q_MX02 U80 ( .S(n45), .A0(\rst_dat[0][31] ), .A1(sw_wdat[31]), .Z(n41));
Q_INV U81 ( .A(n45), .Z(n46));
Q_ND02 U82 ( .A0(n45), .A1(n43), .Z(n42));
Q_AN02 U83 ( .A0(rst_n), .A1(n44), .Z(n45));
Q_INV U84 ( .A(reset), .Z(n44));
Q_ND02 U85 ( .A0(sw_cs), .A1(sw_we), .Z(n43));
Q_MX02 U86 ( .S(sw_we), .A0(n110), .A1(sw_wdat[0]), .Z(n47));
Q_MX02 U87 ( .S(sw_we), .A0(n109), .A1(sw_wdat[1]), .Z(n48));
Q_MX02 U88 ( .S(sw_we), .A0(n108), .A1(sw_wdat[2]), .Z(n49));
Q_MX02 U89 ( .S(sw_we), .A0(n107), .A1(sw_wdat[3]), .Z(n50));
Q_MX02 U90 ( .S(sw_we), .A0(n106), .A1(sw_wdat[4]), .Z(n51));
Q_MX02 U91 ( .S(sw_we), .A0(n105), .A1(sw_wdat[5]), .Z(n52));
Q_MX02 U92 ( .S(sw_we), .A0(n104), .A1(sw_wdat[6]), .Z(n53));
Q_MX02 U93 ( .S(sw_we), .A0(n103), .A1(sw_wdat[7]), .Z(n54));
Q_MX02 U94 ( .S(sw_we), .A0(n102), .A1(sw_wdat[8]), .Z(n55));
Q_MX02 U95 ( .S(sw_we), .A0(n101), .A1(sw_wdat[9]), .Z(n56));
Q_MX02 U96 ( .S(sw_we), .A0(n100), .A1(sw_wdat[10]), .Z(n57));
Q_MX02 U97 ( .S(sw_we), .A0(n99), .A1(sw_wdat[11]), .Z(n58));
Q_MX02 U98 ( .S(sw_we), .A0(n98), .A1(sw_wdat[12]), .Z(n59));
Q_MX02 U99 ( .S(sw_we), .A0(n97), .A1(sw_wdat[13]), .Z(n60));
Q_MX02 U100 ( .S(sw_we), .A0(n96), .A1(sw_wdat[14]), .Z(n61));
Q_MX02 U101 ( .S(sw_we), .A0(n95), .A1(sw_wdat[15]), .Z(n62));
Q_MX02 U102 ( .S(sw_we), .A0(n94), .A1(sw_wdat[16]), .Z(n63));
Q_MX02 U103 ( .S(sw_we), .A0(n93), .A1(sw_wdat[17]), .Z(n64));
Q_MX02 U104 ( .S(sw_we), .A0(n92), .A1(sw_wdat[18]), .Z(n65));
Q_MX02 U105 ( .S(sw_we), .A0(n91), .A1(sw_wdat[19]), .Z(n66));
Q_MX02 U106 ( .S(sw_we), .A0(n90), .A1(sw_wdat[20]), .Z(n67));
Q_MX02 U107 ( .S(sw_we), .A0(n89), .A1(sw_wdat[21]), .Z(n68));
Q_MX02 U108 ( .S(sw_we), .A0(n88), .A1(sw_wdat[22]), .Z(n69));
Q_MX02 U109 ( .S(sw_we), .A0(n87), .A1(sw_wdat[23]), .Z(n70));
Q_MX02 U110 ( .S(sw_we), .A0(n86), .A1(sw_wdat[24]), .Z(n71));
Q_MX02 U111 ( .S(sw_we), .A0(n85), .A1(sw_wdat[25]), .Z(n72));
Q_MX02 U112 ( .S(sw_we), .A0(n84), .A1(sw_wdat[26]), .Z(n73));
Q_MX02 U113 ( .S(sw_we), .A0(n83), .A1(sw_wdat[27]), .Z(n74));
Q_MX02 U114 ( .S(sw_we), .A0(n82), .A1(sw_wdat[28]), .Z(n75));
Q_MX02 U115 ( .S(sw_we), .A0(n81), .A1(sw_wdat[29]), .Z(n76));
Q_MX02 U116 ( .S(sw_we), .A0(n80), .A1(sw_wdat[30]), .Z(n77));
Q_MX02 U117 ( .S(sw_we), .A0(n79), .A1(sw_wdat[31]), .Z(n78));
Q_AN03 U118 ( .A0(_zzM132_bcBehEval[30]), .A1(_zzM132_bcBehEval[29]), .A2(_zzM132_bcBehEval[28]), .Z(n111));
Q_AN03 U119 ( .A0(_zzM132_bcBehEval[27]), .A1(_zzM132_bcBehEval[26]), .A2(_zzM132_bcBehEval[25]), .Z(n112));
Q_AN03 U120 ( .A0(_zzM132_bcBehEval[24]), .A1(_zzM132_bcBehEval[23]), .A2(_zzM132_bcBehEval[22]), .Z(n113));
Q_AN03 U121 ( .A0(_zzM132_bcBehEval[21]), .A1(_zzM132_bcBehEval[20]), .A2(_zzM132_bcBehEval[19]), .Z(n114));
Q_AN03 U122 ( .A0(_zzM132_bcBehEval[18]), .A1(_zzM132_bcBehEval[17]), .A2(_zzM132_bcBehEval[16]), .Z(n115));
Q_AN03 U123 ( .A0(_zzM132_bcBehEval[15]), .A1(_zzM132_bcBehEval[14]), .A2(_zzM132_bcBehEval[13]), .Z(n116));
Q_AN03 U124 ( .A0(_zzM132_bcBehEval[12]), .A1(_zzM132_bcBehEval[11]), .A2(_zzM132_bcBehEval[10]), .Z(n117));
Q_AN03 U125 ( .A0(_zzM132_bcBehEval[9]), .A1(_zzM132_bcBehEval[8]), .A2(_zzM132_bcBehEval[7]), .Z(n118));
Q_AN03 U126 ( .A0(_zzM132_bcBehEval[6]), .A1(_zzM132_bcBehEval[5]), .A2(_zzM132_bcBehEval[4]), .Z(n119));
Q_AN03 U127 ( .A0(_zzM132_bcBehEval[3]), .A1(_zzM132_bcBehEval[2]), .A2(_zzM132_bcBehEval[1]), .Z(n120));
Q_AN03 U128 ( .A0(_zzM132_bcBehEval[0]), .A1(n111), .A2(n112), .Z(n121));
Q_AN03 U129 ( .A0(n113), .A1(n114), .A2(n115), .Z(n122));
Q_AN03 U130 ( .A0(n116), .A1(n117), .A2(n118), .Z(n123));
Q_AN03 U131 ( .A0(n119), .A1(n120), .A2(n121), .Z(n124));
Q_ND03 U132 ( .A0(n122), .A1(n123), .A2(n124), .Z(n125));
Q_AD01HF U133 ( .A0(_zzM132_bcBehEval[1]), .B0(_zzM132_bcBehEval[0]), .S(n126), .CO(n127));
Q_AD01HF U134 ( .A0(_zzM132_bcBehEval[2]), .B0(n127), .S(n128), .CO(n129));
Q_AD01HF U135 ( .A0(_zzM132_bcBehEval[3]), .B0(n129), .S(n130), .CO(n131));
Q_AD01HF U136 ( .A0(_zzM132_bcBehEval[4]), .B0(n131), .S(n132), .CO(n133));
Q_AD01HF U137 ( .A0(_zzM132_bcBehEval[5]), .B0(n133), .S(n134), .CO(n135));
Q_AD01HF U138 ( .A0(_zzM132_bcBehEval[6]), .B0(n135), .S(n136), .CO(n137));
Q_AD01HF U139 ( .A0(_zzM132_bcBehEval[7]), .B0(n137), .S(n138), .CO(n139));
Q_AD01HF U140 ( .A0(_zzM132_bcBehEval[8]), .B0(n139), .S(n140), .CO(n141));
Q_AD01HF U141 ( .A0(_zzM132_bcBehEval[9]), .B0(n141), .S(n142), .CO(n143));
Q_AD01HF U142 ( .A0(_zzM132_bcBehEval[10]), .B0(n143), .S(n144), .CO(n145));
Q_AD01HF U143 ( .A0(_zzM132_bcBehEval[11]), .B0(n145), .S(n146), .CO(n147));
Q_AD01HF U144 ( .A0(_zzM132_bcBehEval[12]), .B0(n147), .S(n148), .CO(n149));
Q_AD01HF U145 ( .A0(_zzM132_bcBehEval[13]), .B0(n149), .S(n150), .CO(n151));
Q_AD01HF U146 ( .A0(_zzM132_bcBehEval[14]), .B0(n151), .S(n152), .CO(n153));
Q_AD01HF U147 ( .A0(_zzM132_bcBehEval[15]), .B0(n153), .S(n154), .CO(n155));
Q_AD01HF U148 ( .A0(_zzM132_bcBehEval[16]), .B0(n155), .S(n156), .CO(n157));
Q_AD01HF U149 ( .A0(_zzM132_bcBehEval[17]), .B0(n157), .S(n158), .CO(n159));
Q_AD01HF U150 ( .A0(_zzM132_bcBehEval[18]), .B0(n159), .S(n160), .CO(n161));
Q_AD01HF U151 ( .A0(_zzM132_bcBehEval[19]), .B0(n161), .S(n162), .CO(n163));
Q_AD01HF U152 ( .A0(_zzM132_bcBehEval[20]), .B0(n163), .S(n164), .CO(n165));
Q_AD01HF U153 ( .A0(_zzM132_bcBehEval[21]), .B0(n165), .S(n166), .CO(n167));
Q_AD01HF U154 ( .A0(_zzM132_bcBehEval[22]), .B0(n167), .S(n168), .CO(n169));
Q_AD01HF U155 ( .A0(_zzM132_bcBehEval[23]), .B0(n169), .S(n170), .CO(n171));
Q_AD01HF U156 ( .A0(_zzM132_bcBehEval[24]), .B0(n171), .S(n172), .CO(n173));
Q_AD01HF U157 ( .A0(_zzM132_bcBehEval[25]), .B0(n173), .S(n174), .CO(n175));
Q_AD01HF U158 ( .A0(_zzM132_bcBehEval[26]), .B0(n175), .S(n176), .CO(n177));
Q_AD01HF U159 ( .A0(_zzM132_bcBehEval[27]), .B0(n177), .S(n178), .CO(n179));
Q_AD01HF U160 ( .A0(_zzM132_bcBehEval[28]), .B0(n179), .S(n180), .CO(n181));
Q_AD01HF U161 ( .A0(_zzM132_bcBehEval[29]), .B0(n181), .S(n182), .CO(n183));
Q_AN02 U162 ( .A0(_zzM132L132_bcWait0), .A1(n125), .Z(n184));
Q_INV U163 ( .A(n185), .Z(n190));
Q_INV U164 ( .A(n186), .Z(n191));
Q_NR02 U165 ( .A0(n186), .A1(n185), .Z(n192));
Q_AN02 U166 ( .A0(n191), .A1(n185), .Z(n193));
Q_AN02 U167 ( .A0(n186), .A1(n190), .Z(n194));
Q_AN02 U168 ( .A0(n186), .A1(n185), .Z(n195));
Q_INV U169 ( .A(n187), .Z(n196));
Q_INV U170 ( .A(n188), .Z(n197));
Q_INV U171 ( .A(n189), .Z(n198));
Q_NR02 U172 ( .A0(n189), .A1(n188), .Z(n199));
Q_AN02 U173 ( .A0(n198), .A1(n188), .Z(n200));
Q_AN02 U174 ( .A0(n189), .A1(n197), .Z(n201));
Q_AN02 U175 ( .A0(n189), .A1(n188), .Z(n202));
Q_AN02 U176 ( .A0(n199), .A1(n196), .Z(n203));
Q_AN02 U177 ( .A0(n199), .A1(n187), .Z(n204));
Q_AN02 U178 ( .A0(n200), .A1(n196), .Z(n205));
Q_AN02 U179 ( .A0(n200), .A1(n187), .Z(n206));
Q_AN02 U180 ( .A0(n201), .A1(n196), .Z(n207));
Q_AN02 U181 ( .A0(n201), .A1(n187), .Z(n208));
Q_AN02 U182 ( .A0(n202), .A1(n196), .Z(n209));
Q_AN02 U183 ( .A0(n202), .A1(n187), .Z(n210));
Q_AN03 U184 ( .A0(n203), .A1(n192), .A2(n42), .Z(n211));
Q_AO21 U185 ( .A0(n203), .A1(n193), .B0(n46), .Z(n212));
Q_AO21 U186 ( .A0(n203), .A1(n194), .B0(n46), .Z(n245));
Q_AO21 U187 ( .A0(n203), .A1(n195), .B0(n46), .Z(n278));
Q_AO21 U188 ( .A0(n204), .A1(n192), .B0(n46), .Z(n311));
Q_AO21 U189 ( .A0(n204), .A1(n193), .B0(n46), .Z(n344));
Q_AO21 U190 ( .A0(n204), .A1(n194), .B0(n46), .Z(n377));
Q_AO21 U191 ( .A0(n204), .A1(n195), .B0(n46), .Z(n410));
Q_AO21 U192 ( .A0(n205), .A1(n192), .B0(n46), .Z(n443));
Q_AO21 U193 ( .A0(n205), .A1(n193), .B0(n46), .Z(n476));
Q_AO21 U194 ( .A0(n205), .A1(n194), .B0(n46), .Z(n509));
Q_AO21 U195 ( .A0(n205), .A1(n195), .B0(n46), .Z(n542));
Q_AO21 U196 ( .A0(n206), .A1(n192), .B0(n46), .Z(n575));
Q_AO21 U197 ( .A0(n206), .A1(n193), .B0(n46), .Z(n608));
Q_AO21 U198 ( .A0(n206), .A1(n194), .B0(n46), .Z(n641));
Q_AO21 U199 ( .A0(n206), .A1(n195), .B0(n46), .Z(n674));
Q_AO21 U200 ( .A0(n207), .A1(n192), .B0(n46), .Z(n707));
Q_AO21 U201 ( .A0(n207), .A1(n193), .B0(n46), .Z(n740));
Q_AO21 U202 ( .A0(n207), .A1(n194), .B0(n46), .Z(n773));
Q_AO21 U203 ( .A0(n207), .A1(n195), .B0(n46), .Z(n806));
Q_AO21 U204 ( .A0(n208), .A1(n192), .B0(n46), .Z(n839));
Q_AO21 U205 ( .A0(n208), .A1(n193), .B0(n46), .Z(n872));
Q_AO21 U206 ( .A0(n208), .A1(n194), .B0(n46), .Z(n905));
Q_AO21 U207 ( .A0(n208), .A1(n195), .B0(n46), .Z(n938));
Q_AO21 U208 ( .A0(n209), .A1(n192), .B0(n46), .Z(n971));
Q_AO21 U209 ( .A0(n209), .A1(n193), .B0(n46), .Z(n1004));
Q_AO21 U210 ( .A0(n209), .A1(n194), .B0(n46), .Z(n1037));
Q_AO21 U211 ( .A0(n209), .A1(n195), .B0(n46), .Z(n1070));
Q_AO21 U212 ( .A0(n210), .A1(n192), .B0(n46), .Z(n1103));
Q_AO21 U213 ( .A0(n210), .A1(n193), .B0(n46), .Z(n1136));
Q_AO21 U214 ( .A0(n210), .A1(n194), .B0(n46), .Z(n1169));
Q_AO21 U215 ( .A0(n210), .A1(n195), .B0(n46), .Z(n1202));
Q_MX02 U216 ( .S(n45), .A0(\rst_dat[1][0] ), .A1(n10), .Z(n213));
Q_MX02 U217 ( .S(n45), .A0(\rst_dat[1][1] ), .A1(n11), .Z(n214));
Q_MX02 U218 ( .S(n45), .A0(\rst_dat[1][2] ), .A1(n12), .Z(n215));
Q_MX02 U219 ( .S(n45), .A0(\rst_dat[1][3] ), .A1(n13), .Z(n216));
Q_MX02 U220 ( .S(n45), .A0(\rst_dat[1][4] ), .A1(n14), .Z(n217));
Q_MX02 U221 ( .S(n45), .A0(\rst_dat[1][5] ), .A1(n15), .Z(n218));
Q_MX02 U222 ( .S(n45), .A0(\rst_dat[1][6] ), .A1(n16), .Z(n219));
Q_MX02 U223 ( .S(n45), .A0(\rst_dat[1][7] ), .A1(n17), .Z(n220));
Q_MX02 U224 ( .S(n45), .A0(\rst_dat[1][8] ), .A1(n18), .Z(n221));
Q_MX02 U225 ( .S(n45), .A0(\rst_dat[1][9] ), .A1(n19), .Z(n222));
Q_MX02 U226 ( .S(n45), .A0(\rst_dat[1][10] ), .A1(n20), .Z(n223));
Q_MX02 U227 ( .S(n45), .A0(\rst_dat[1][11] ), .A1(n21), .Z(n224));
Q_MX02 U228 ( .S(n45), .A0(\rst_dat[1][12] ), .A1(n22), .Z(n225));
Q_MX02 U229 ( .S(n45), .A0(\rst_dat[1][13] ), .A1(n23), .Z(n226));
Q_MX02 U230 ( .S(n45), .A0(\rst_dat[1][14] ), .A1(n24), .Z(n227));
Q_MX02 U231 ( .S(n45), .A0(\rst_dat[1][15] ), .A1(n25), .Z(n228));
Q_MX02 U232 ( .S(n45), .A0(\rst_dat[1][16] ), .A1(n26), .Z(n229));
Q_MX02 U233 ( .S(n45), .A0(\rst_dat[1][17] ), .A1(n27), .Z(n230));
Q_MX02 U234 ( .S(n45), .A0(\rst_dat[1][18] ), .A1(n28), .Z(n231));
Q_MX02 U235 ( .S(n45), .A0(\rst_dat[1][19] ), .A1(n29), .Z(n232));
Q_MX02 U236 ( .S(n45), .A0(\rst_dat[1][20] ), .A1(n30), .Z(n233));
Q_MX02 U237 ( .S(n45), .A0(\rst_dat[1][21] ), .A1(n31), .Z(n234));
Q_MX02 U238 ( .S(n45), .A0(\rst_dat[1][22] ), .A1(n32), .Z(n235));
Q_MX02 U239 ( .S(n45), .A0(\rst_dat[1][23] ), .A1(n33), .Z(n236));
Q_MX02 U240 ( .S(n45), .A0(\rst_dat[1][24] ), .A1(n34), .Z(n237));
Q_MX02 U241 ( .S(n45), .A0(\rst_dat[1][25] ), .A1(n35), .Z(n238));
Q_MX02 U242 ( .S(n45), .A0(\rst_dat[1][26] ), .A1(n36), .Z(n239));
Q_MX02 U243 ( .S(n45), .A0(\rst_dat[1][27] ), .A1(n37), .Z(n240));
Q_MX02 U244 ( .S(n45), .A0(\rst_dat[1][28] ), .A1(n38), .Z(n241));
Q_MX02 U245 ( .S(n45), .A0(\rst_dat[1][29] ), .A1(n39), .Z(n242));
Q_MX02 U246 ( .S(n45), .A0(\rst_dat[1][30] ), .A1(n40), .Z(n243));
Q_MX02 U247 ( .S(n45), .A0(\rst_dat[1][31] ), .A1(n41), .Z(n244));
Q_MX02 U248 ( .S(n45), .A0(\rst_dat[2][0] ), .A1(n10), .Z(n246));
Q_MX02 U249 ( .S(n45), .A0(\rst_dat[2][1] ), .A1(n11), .Z(n247));
Q_MX02 U250 ( .S(n45), .A0(\rst_dat[2][2] ), .A1(n12), .Z(n248));
Q_MX02 U251 ( .S(n45), .A0(\rst_dat[2][3] ), .A1(n13), .Z(n249));
Q_MX02 U252 ( .S(n45), .A0(\rst_dat[2][4] ), .A1(n14), .Z(n250));
Q_MX02 U253 ( .S(n45), .A0(\rst_dat[2][5] ), .A1(n15), .Z(n251));
Q_MX02 U254 ( .S(n45), .A0(\rst_dat[2][6] ), .A1(n16), .Z(n252));
Q_MX02 U255 ( .S(n45), .A0(\rst_dat[2][7] ), .A1(n17), .Z(n253));
Q_MX02 U256 ( .S(n45), .A0(\rst_dat[2][8] ), .A1(n18), .Z(n254));
Q_MX02 U257 ( .S(n45), .A0(\rst_dat[2][9] ), .A1(n19), .Z(n255));
Q_MX02 U258 ( .S(n45), .A0(\rst_dat[2][10] ), .A1(n20), .Z(n256));
Q_MX02 U259 ( .S(n45), .A0(\rst_dat[2][11] ), .A1(n21), .Z(n257));
Q_MX02 U260 ( .S(n45), .A0(\rst_dat[2][12] ), .A1(n22), .Z(n258));
Q_MX02 U261 ( .S(n45), .A0(\rst_dat[2][13] ), .A1(n23), .Z(n259));
Q_MX02 U262 ( .S(n45), .A0(\rst_dat[2][14] ), .A1(n24), .Z(n260));
Q_MX02 U263 ( .S(n45), .A0(\rst_dat[2][15] ), .A1(n25), .Z(n261));
Q_MX02 U264 ( .S(n45), .A0(\rst_dat[2][16] ), .A1(n26), .Z(n262));
Q_MX02 U265 ( .S(n45), .A0(\rst_dat[2][17] ), .A1(n27), .Z(n263));
Q_MX02 U266 ( .S(n45), .A0(\rst_dat[2][18] ), .A1(n28), .Z(n264));
Q_MX02 U267 ( .S(n45), .A0(\rst_dat[2][19] ), .A1(n29), .Z(n265));
Q_MX02 U268 ( .S(n45), .A0(\rst_dat[2][20] ), .A1(n30), .Z(n266));
Q_MX02 U269 ( .S(n45), .A0(\rst_dat[2][21] ), .A1(n31), .Z(n267));
Q_MX02 U270 ( .S(n45), .A0(\rst_dat[2][22] ), .A1(n32), .Z(n268));
Q_MX02 U271 ( .S(n45), .A0(\rst_dat[2][23] ), .A1(n33), .Z(n269));
Q_MX02 U272 ( .S(n45), .A0(\rst_dat[2][24] ), .A1(n34), .Z(n270));
Q_MX02 U273 ( .S(n45), .A0(\rst_dat[2][25] ), .A1(n35), .Z(n271));
Q_MX02 U274 ( .S(n45), .A0(\rst_dat[2][26] ), .A1(n36), .Z(n272));
Q_MX02 U275 ( .S(n45), .A0(\rst_dat[2][27] ), .A1(n37), .Z(n273));
Q_MX02 U276 ( .S(n45), .A0(\rst_dat[2][28] ), .A1(n38), .Z(n274));
Q_MX02 U277 ( .S(n45), .A0(\rst_dat[2][29] ), .A1(n39), .Z(n275));
Q_MX02 U278 ( .S(n45), .A0(\rst_dat[2][30] ), .A1(n40), .Z(n276));
Q_MX02 U279 ( .S(n45), .A0(\rst_dat[2][31] ), .A1(n41), .Z(n277));
Q_MX02 U280 ( .S(n45), .A0(\rst_dat[3][0] ), .A1(n10), .Z(n279));
Q_MX02 U281 ( .S(n45), .A0(\rst_dat[3][1] ), .A1(n11), .Z(n280));
Q_MX02 U282 ( .S(n45), .A0(\rst_dat[3][2] ), .A1(n12), .Z(n281));
Q_MX02 U283 ( .S(n45), .A0(\rst_dat[3][3] ), .A1(n13), .Z(n282));
Q_MX02 U284 ( .S(n45), .A0(\rst_dat[3][4] ), .A1(n14), .Z(n283));
Q_MX02 U285 ( .S(n45), .A0(\rst_dat[3][5] ), .A1(n15), .Z(n284));
Q_MX02 U286 ( .S(n45), .A0(\rst_dat[3][6] ), .A1(n16), .Z(n285));
Q_MX02 U287 ( .S(n45), .A0(\rst_dat[3][7] ), .A1(n17), .Z(n286));
Q_MX02 U288 ( .S(n45), .A0(\rst_dat[3][8] ), .A1(n18), .Z(n287));
Q_MX02 U289 ( .S(n45), .A0(\rst_dat[3][9] ), .A1(n19), .Z(n288));
Q_MX02 U290 ( .S(n45), .A0(\rst_dat[3][10] ), .A1(n20), .Z(n289));
Q_MX02 U291 ( .S(n45), .A0(\rst_dat[3][11] ), .A1(n21), .Z(n290));
Q_MX02 U292 ( .S(n45), .A0(\rst_dat[3][12] ), .A1(n22), .Z(n291));
Q_MX02 U293 ( .S(n45), .A0(\rst_dat[3][13] ), .A1(n23), .Z(n292));
Q_MX02 U294 ( .S(n45), .A0(\rst_dat[3][14] ), .A1(n24), .Z(n293));
Q_MX02 U295 ( .S(n45), .A0(\rst_dat[3][15] ), .A1(n25), .Z(n294));
Q_MX02 U296 ( .S(n45), .A0(\rst_dat[3][16] ), .A1(n26), .Z(n295));
Q_MX02 U297 ( .S(n45), .A0(\rst_dat[3][17] ), .A1(n27), .Z(n296));
Q_MX02 U298 ( .S(n45), .A0(\rst_dat[3][18] ), .A1(n28), .Z(n297));
Q_MX02 U299 ( .S(n45), .A0(\rst_dat[3][19] ), .A1(n29), .Z(n298));
Q_MX02 U300 ( .S(n45), .A0(\rst_dat[3][20] ), .A1(n30), .Z(n299));
Q_MX02 U301 ( .S(n45), .A0(\rst_dat[3][21] ), .A1(n31), .Z(n300));
Q_MX02 U302 ( .S(n45), .A0(\rst_dat[3][22] ), .A1(n32), .Z(n301));
Q_MX02 U303 ( .S(n45), .A0(\rst_dat[3][23] ), .A1(n33), .Z(n302));
Q_MX02 U304 ( .S(n45), .A0(\rst_dat[3][24] ), .A1(n34), .Z(n303));
Q_MX02 U305 ( .S(n45), .A0(\rst_dat[3][25] ), .A1(n35), .Z(n304));
Q_MX02 U306 ( .S(n45), .A0(\rst_dat[3][26] ), .A1(n36), .Z(n305));
Q_MX02 U307 ( .S(n45), .A0(\rst_dat[3][27] ), .A1(n37), .Z(n306));
Q_MX02 U308 ( .S(n45), .A0(\rst_dat[3][28] ), .A1(n38), .Z(n307));
Q_MX02 U309 ( .S(n45), .A0(\rst_dat[3][29] ), .A1(n39), .Z(n308));
Q_MX02 U310 ( .S(n45), .A0(\rst_dat[3][30] ), .A1(n40), .Z(n309));
Q_MX02 U311 ( .S(n45), .A0(\rst_dat[3][31] ), .A1(n41), .Z(n310));
Q_MX02 U312 ( .S(n45), .A0(\rst_dat[4][0] ), .A1(n10), .Z(n312));
Q_MX02 U313 ( .S(n45), .A0(\rst_dat[4][1] ), .A1(n11), .Z(n313));
Q_MX02 U314 ( .S(n45), .A0(\rst_dat[4][2] ), .A1(n12), .Z(n314));
Q_MX02 U315 ( .S(n45), .A0(\rst_dat[4][3] ), .A1(n13), .Z(n315));
Q_MX02 U316 ( .S(n45), .A0(\rst_dat[4][4] ), .A1(n14), .Z(n316));
Q_MX02 U317 ( .S(n45), .A0(\rst_dat[4][5] ), .A1(n15), .Z(n317));
Q_MX02 U318 ( .S(n45), .A0(\rst_dat[4][6] ), .A1(n16), .Z(n318));
Q_MX02 U319 ( .S(n45), .A0(\rst_dat[4][7] ), .A1(n17), .Z(n319));
Q_MX02 U320 ( .S(n45), .A0(\rst_dat[4][8] ), .A1(n18), .Z(n320));
Q_MX02 U321 ( .S(n45), .A0(\rst_dat[4][9] ), .A1(n19), .Z(n321));
Q_MX02 U322 ( .S(n45), .A0(\rst_dat[4][10] ), .A1(n20), .Z(n322));
Q_MX02 U323 ( .S(n45), .A0(\rst_dat[4][11] ), .A1(n21), .Z(n323));
Q_MX02 U324 ( .S(n45), .A0(\rst_dat[4][12] ), .A1(n22), .Z(n324));
Q_MX02 U325 ( .S(n45), .A0(\rst_dat[4][13] ), .A1(n23), .Z(n325));
Q_MX02 U326 ( .S(n45), .A0(\rst_dat[4][14] ), .A1(n24), .Z(n326));
Q_MX02 U327 ( .S(n45), .A0(\rst_dat[4][15] ), .A1(n25), .Z(n327));
Q_MX02 U328 ( .S(n45), .A0(\rst_dat[4][16] ), .A1(n26), .Z(n328));
Q_MX02 U329 ( .S(n45), .A0(\rst_dat[4][17] ), .A1(n27), .Z(n329));
Q_MX02 U330 ( .S(n45), .A0(\rst_dat[4][18] ), .A1(n28), .Z(n330));
Q_MX02 U331 ( .S(n45), .A0(\rst_dat[4][19] ), .A1(n29), .Z(n331));
Q_MX02 U332 ( .S(n45), .A0(\rst_dat[4][20] ), .A1(n30), .Z(n332));
Q_MX02 U333 ( .S(n45), .A0(\rst_dat[4][21] ), .A1(n31), .Z(n333));
Q_MX02 U334 ( .S(n45), .A0(\rst_dat[4][22] ), .A1(n32), .Z(n334));
Q_MX02 U335 ( .S(n45), .A0(\rst_dat[4][23] ), .A1(n33), .Z(n335));
Q_MX02 U336 ( .S(n45), .A0(\rst_dat[4][24] ), .A1(n34), .Z(n336));
Q_MX02 U337 ( .S(n45), .A0(\rst_dat[4][25] ), .A1(n35), .Z(n337));
Q_MX02 U338 ( .S(n45), .A0(\rst_dat[4][26] ), .A1(n36), .Z(n338));
Q_MX02 U339 ( .S(n45), .A0(\rst_dat[4][27] ), .A1(n37), .Z(n339));
Q_MX02 U340 ( .S(n45), .A0(\rst_dat[4][28] ), .A1(n38), .Z(n340));
Q_MX02 U341 ( .S(n45), .A0(\rst_dat[4][29] ), .A1(n39), .Z(n341));
Q_MX02 U342 ( .S(n45), .A0(\rst_dat[4][30] ), .A1(n40), .Z(n342));
Q_MX02 U343 ( .S(n45), .A0(\rst_dat[4][31] ), .A1(n41), .Z(n343));
Q_MX02 U344 ( .S(n45), .A0(\rst_dat[5][0] ), .A1(n10), .Z(n345));
Q_MX02 U345 ( .S(n45), .A0(\rst_dat[5][1] ), .A1(n11), .Z(n346));
Q_MX02 U346 ( .S(n45), .A0(\rst_dat[5][2] ), .A1(n12), .Z(n347));
Q_MX02 U347 ( .S(n45), .A0(\rst_dat[5][3] ), .A1(n13), .Z(n348));
Q_MX02 U348 ( .S(n45), .A0(\rst_dat[5][4] ), .A1(n14), .Z(n349));
Q_MX02 U349 ( .S(n45), .A0(\rst_dat[5][5] ), .A1(n15), .Z(n350));
Q_MX02 U350 ( .S(n45), .A0(\rst_dat[5][6] ), .A1(n16), .Z(n351));
Q_MX02 U351 ( .S(n45), .A0(\rst_dat[5][7] ), .A1(n17), .Z(n352));
Q_MX02 U352 ( .S(n45), .A0(\rst_dat[5][8] ), .A1(n18), .Z(n353));
Q_MX02 U353 ( .S(n45), .A0(\rst_dat[5][9] ), .A1(n19), .Z(n354));
Q_MX02 U354 ( .S(n45), .A0(\rst_dat[5][10] ), .A1(n20), .Z(n355));
Q_MX02 U355 ( .S(n45), .A0(\rst_dat[5][11] ), .A1(n21), .Z(n356));
Q_MX02 U356 ( .S(n45), .A0(\rst_dat[5][12] ), .A1(n22), .Z(n357));
Q_MX02 U357 ( .S(n45), .A0(\rst_dat[5][13] ), .A1(n23), .Z(n358));
Q_MX02 U358 ( .S(n45), .A0(\rst_dat[5][14] ), .A1(n24), .Z(n359));
Q_MX02 U359 ( .S(n45), .A0(\rst_dat[5][15] ), .A1(n25), .Z(n360));
Q_MX02 U360 ( .S(n45), .A0(\rst_dat[5][16] ), .A1(n26), .Z(n361));
Q_MX02 U361 ( .S(n45), .A0(\rst_dat[5][17] ), .A1(n27), .Z(n362));
Q_MX02 U362 ( .S(n45), .A0(\rst_dat[5][18] ), .A1(n28), .Z(n363));
Q_MX02 U363 ( .S(n45), .A0(\rst_dat[5][19] ), .A1(n29), .Z(n364));
Q_MX02 U364 ( .S(n45), .A0(\rst_dat[5][20] ), .A1(n30), .Z(n365));
Q_MX02 U365 ( .S(n45), .A0(\rst_dat[5][21] ), .A1(n31), .Z(n366));
Q_MX02 U366 ( .S(n45), .A0(\rst_dat[5][22] ), .A1(n32), .Z(n367));
Q_MX02 U367 ( .S(n45), .A0(\rst_dat[5][23] ), .A1(n33), .Z(n368));
Q_MX02 U368 ( .S(n45), .A0(\rst_dat[5][24] ), .A1(n34), .Z(n369));
Q_MX02 U369 ( .S(n45), .A0(\rst_dat[5][25] ), .A1(n35), .Z(n370));
Q_MX02 U370 ( .S(n45), .A0(\rst_dat[5][26] ), .A1(n36), .Z(n371));
Q_MX02 U371 ( .S(n45), .A0(\rst_dat[5][27] ), .A1(n37), .Z(n372));
Q_MX02 U372 ( .S(n45), .A0(\rst_dat[5][28] ), .A1(n38), .Z(n373));
Q_MX02 U373 ( .S(n45), .A0(\rst_dat[5][29] ), .A1(n39), .Z(n374));
Q_MX02 U374 ( .S(n45), .A0(\rst_dat[5][30] ), .A1(n40), .Z(n375));
Q_MX02 U375 ( .S(n45), .A0(\rst_dat[5][31] ), .A1(n41), .Z(n376));
Q_MX02 U376 ( .S(n45), .A0(\rst_dat[6][0] ), .A1(n10), .Z(n378));
Q_MX02 U377 ( .S(n45), .A0(\rst_dat[6][1] ), .A1(n11), .Z(n379));
Q_MX02 U378 ( .S(n45), .A0(\rst_dat[6][2] ), .A1(n12), .Z(n380));
Q_MX02 U379 ( .S(n45), .A0(\rst_dat[6][3] ), .A1(n13), .Z(n381));
Q_MX02 U380 ( .S(n45), .A0(\rst_dat[6][4] ), .A1(n14), .Z(n382));
Q_MX02 U381 ( .S(n45), .A0(\rst_dat[6][5] ), .A1(n15), .Z(n383));
Q_MX02 U382 ( .S(n45), .A0(\rst_dat[6][6] ), .A1(n16), .Z(n384));
Q_MX02 U383 ( .S(n45), .A0(\rst_dat[6][7] ), .A1(n17), .Z(n385));
Q_MX02 U384 ( .S(n45), .A0(\rst_dat[6][8] ), .A1(n18), .Z(n386));
Q_MX02 U385 ( .S(n45), .A0(\rst_dat[6][9] ), .A1(n19), .Z(n387));
Q_MX02 U386 ( .S(n45), .A0(\rst_dat[6][10] ), .A1(n20), .Z(n388));
Q_MX02 U387 ( .S(n45), .A0(\rst_dat[6][11] ), .A1(n21), .Z(n389));
Q_MX02 U388 ( .S(n45), .A0(\rst_dat[6][12] ), .A1(n22), .Z(n390));
Q_MX02 U389 ( .S(n45), .A0(\rst_dat[6][13] ), .A1(n23), .Z(n391));
Q_MX02 U390 ( .S(n45), .A0(\rst_dat[6][14] ), .A1(n24), .Z(n392));
Q_MX02 U391 ( .S(n45), .A0(\rst_dat[6][15] ), .A1(n25), .Z(n393));
Q_MX02 U392 ( .S(n45), .A0(\rst_dat[6][16] ), .A1(n26), .Z(n394));
Q_MX02 U393 ( .S(n45), .A0(\rst_dat[6][17] ), .A1(n27), .Z(n395));
Q_MX02 U394 ( .S(n45), .A0(\rst_dat[6][18] ), .A1(n28), .Z(n396));
Q_MX02 U395 ( .S(n45), .A0(\rst_dat[6][19] ), .A1(n29), .Z(n397));
Q_MX02 U396 ( .S(n45), .A0(\rst_dat[6][20] ), .A1(n30), .Z(n398));
Q_MX02 U397 ( .S(n45), .A0(\rst_dat[6][21] ), .A1(n31), .Z(n399));
Q_MX02 U398 ( .S(n45), .A0(\rst_dat[6][22] ), .A1(n32), .Z(n400));
Q_MX02 U399 ( .S(n45), .A0(\rst_dat[6][23] ), .A1(n33), .Z(n401));
Q_MX02 U400 ( .S(n45), .A0(\rst_dat[6][24] ), .A1(n34), .Z(n402));
Q_MX02 U401 ( .S(n45), .A0(\rst_dat[6][25] ), .A1(n35), .Z(n403));
Q_MX02 U402 ( .S(n45), .A0(\rst_dat[6][26] ), .A1(n36), .Z(n404));
Q_MX02 U403 ( .S(n45), .A0(\rst_dat[6][27] ), .A1(n37), .Z(n405));
Q_MX02 U404 ( .S(n45), .A0(\rst_dat[6][28] ), .A1(n38), .Z(n406));
Q_MX02 U405 ( .S(n45), .A0(\rst_dat[6][29] ), .A1(n39), .Z(n407));
Q_MX02 U406 ( .S(n45), .A0(\rst_dat[6][30] ), .A1(n40), .Z(n408));
Q_MX02 U407 ( .S(n45), .A0(\rst_dat[6][31] ), .A1(n41), .Z(n409));
Q_MX02 U408 ( .S(n45), .A0(\rst_dat[7][0] ), .A1(n10), .Z(n411));
Q_MX02 U409 ( .S(n45), .A0(\rst_dat[7][1] ), .A1(n11), .Z(n412));
Q_MX02 U410 ( .S(n45), .A0(\rst_dat[7][2] ), .A1(n12), .Z(n413));
Q_MX02 U411 ( .S(n45), .A0(\rst_dat[7][3] ), .A1(n13), .Z(n414));
Q_MX02 U412 ( .S(n45), .A0(\rst_dat[7][4] ), .A1(n14), .Z(n415));
Q_MX02 U413 ( .S(n45), .A0(\rst_dat[7][5] ), .A1(n15), .Z(n416));
Q_MX02 U414 ( .S(n45), .A0(\rst_dat[7][6] ), .A1(n16), .Z(n417));
Q_MX02 U415 ( .S(n45), .A0(\rst_dat[7][7] ), .A1(n17), .Z(n418));
Q_MX02 U416 ( .S(n45), .A0(\rst_dat[7][8] ), .A1(n18), .Z(n419));
Q_MX02 U417 ( .S(n45), .A0(\rst_dat[7][9] ), .A1(n19), .Z(n420));
Q_MX02 U418 ( .S(n45), .A0(\rst_dat[7][10] ), .A1(n20), .Z(n421));
Q_MX02 U419 ( .S(n45), .A0(\rst_dat[7][11] ), .A1(n21), .Z(n422));
Q_MX02 U420 ( .S(n45), .A0(\rst_dat[7][12] ), .A1(n22), .Z(n423));
Q_MX02 U421 ( .S(n45), .A0(\rst_dat[7][13] ), .A1(n23), .Z(n424));
Q_MX02 U422 ( .S(n45), .A0(\rst_dat[7][14] ), .A1(n24), .Z(n425));
Q_MX02 U423 ( .S(n45), .A0(\rst_dat[7][15] ), .A1(n25), .Z(n426));
Q_MX02 U424 ( .S(n45), .A0(\rst_dat[7][16] ), .A1(n26), .Z(n427));
Q_MX02 U425 ( .S(n45), .A0(\rst_dat[7][17] ), .A1(n27), .Z(n428));
Q_MX02 U426 ( .S(n45), .A0(\rst_dat[7][18] ), .A1(n28), .Z(n429));
Q_MX02 U427 ( .S(n45), .A0(\rst_dat[7][19] ), .A1(n29), .Z(n430));
Q_MX02 U428 ( .S(n45), .A0(\rst_dat[7][20] ), .A1(n30), .Z(n431));
Q_MX02 U429 ( .S(n45), .A0(\rst_dat[7][21] ), .A1(n31), .Z(n432));
Q_MX02 U430 ( .S(n45), .A0(\rst_dat[7][22] ), .A1(n32), .Z(n433));
Q_MX02 U431 ( .S(n45), .A0(\rst_dat[7][23] ), .A1(n33), .Z(n434));
Q_MX02 U432 ( .S(n45), .A0(\rst_dat[7][24] ), .A1(n34), .Z(n435));
Q_MX02 U433 ( .S(n45), .A0(\rst_dat[7][25] ), .A1(n35), .Z(n436));
Q_MX02 U434 ( .S(n45), .A0(\rst_dat[7][26] ), .A1(n36), .Z(n437));
Q_MX02 U435 ( .S(n45), .A0(\rst_dat[7][27] ), .A1(n37), .Z(n438));
Q_MX02 U436 ( .S(n45), .A0(\rst_dat[7][28] ), .A1(n38), .Z(n439));
Q_MX02 U437 ( .S(n45), .A0(\rst_dat[7][29] ), .A1(n39), .Z(n440));
Q_MX02 U438 ( .S(n45), .A0(\rst_dat[7][30] ), .A1(n40), .Z(n441));
Q_MX02 U439 ( .S(n45), .A0(\rst_dat[7][31] ), .A1(n41), .Z(n442));
Q_MX02 U440 ( .S(n45), .A0(\rst_dat[8][0] ), .A1(n10), .Z(n444));
Q_MX02 U441 ( .S(n45), .A0(\rst_dat[8][1] ), .A1(n11), .Z(n445));
Q_MX02 U442 ( .S(n45), .A0(\rst_dat[8][2] ), .A1(n12), .Z(n446));
Q_MX02 U443 ( .S(n45), .A0(\rst_dat[8][3] ), .A1(n13), .Z(n447));
Q_MX02 U444 ( .S(n45), .A0(\rst_dat[8][4] ), .A1(n14), .Z(n448));
Q_MX02 U445 ( .S(n45), .A0(\rst_dat[8][5] ), .A1(n15), .Z(n449));
Q_MX02 U446 ( .S(n45), .A0(\rst_dat[8][6] ), .A1(n16), .Z(n450));
Q_MX02 U447 ( .S(n45), .A0(\rst_dat[8][7] ), .A1(n17), .Z(n451));
Q_MX02 U448 ( .S(n45), .A0(\rst_dat[8][8] ), .A1(n18), .Z(n452));
Q_MX02 U449 ( .S(n45), .A0(\rst_dat[8][9] ), .A1(n19), .Z(n453));
Q_MX02 U450 ( .S(n45), .A0(\rst_dat[8][10] ), .A1(n20), .Z(n454));
Q_MX02 U451 ( .S(n45), .A0(\rst_dat[8][11] ), .A1(n21), .Z(n455));
Q_MX02 U452 ( .S(n45), .A0(\rst_dat[8][12] ), .A1(n22), .Z(n456));
Q_MX02 U453 ( .S(n45), .A0(\rst_dat[8][13] ), .A1(n23), .Z(n457));
Q_MX02 U454 ( .S(n45), .A0(\rst_dat[8][14] ), .A1(n24), .Z(n458));
Q_MX02 U455 ( .S(n45), .A0(\rst_dat[8][15] ), .A1(n25), .Z(n459));
Q_MX02 U456 ( .S(n45), .A0(\rst_dat[8][16] ), .A1(n26), .Z(n460));
Q_MX02 U457 ( .S(n45), .A0(\rst_dat[8][17] ), .A1(n27), .Z(n461));
Q_MX02 U458 ( .S(n45), .A0(\rst_dat[8][18] ), .A1(n28), .Z(n462));
Q_MX02 U459 ( .S(n45), .A0(\rst_dat[8][19] ), .A1(n29), .Z(n463));
Q_MX02 U460 ( .S(n45), .A0(\rst_dat[8][20] ), .A1(n30), .Z(n464));
Q_MX02 U461 ( .S(n45), .A0(\rst_dat[8][21] ), .A1(n31), .Z(n465));
Q_MX02 U462 ( .S(n45), .A0(\rst_dat[8][22] ), .A1(n32), .Z(n466));
Q_MX02 U463 ( .S(n45), .A0(\rst_dat[8][23] ), .A1(n33), .Z(n467));
Q_MX02 U464 ( .S(n45), .A0(\rst_dat[8][24] ), .A1(n34), .Z(n468));
Q_MX02 U465 ( .S(n45), .A0(\rst_dat[8][25] ), .A1(n35), .Z(n469));
Q_MX02 U466 ( .S(n45), .A0(\rst_dat[8][26] ), .A1(n36), .Z(n470));
Q_MX02 U467 ( .S(n45), .A0(\rst_dat[8][27] ), .A1(n37), .Z(n471));
Q_MX02 U468 ( .S(n45), .A0(\rst_dat[8][28] ), .A1(n38), .Z(n472));
Q_MX02 U469 ( .S(n45), .A0(\rst_dat[8][29] ), .A1(n39), .Z(n473));
Q_MX02 U470 ( .S(n45), .A0(\rst_dat[8][30] ), .A1(n40), .Z(n474));
Q_MX02 U471 ( .S(n45), .A0(\rst_dat[8][31] ), .A1(n41), .Z(n475));
Q_MX02 U472 ( .S(n45), .A0(\rst_dat[9][0] ), .A1(n10), .Z(n477));
Q_MX02 U473 ( .S(n45), .A0(\rst_dat[9][1] ), .A1(n11), .Z(n478));
Q_MX02 U474 ( .S(n45), .A0(\rst_dat[9][2] ), .A1(n12), .Z(n479));
Q_MX02 U475 ( .S(n45), .A0(\rst_dat[9][3] ), .A1(n13), .Z(n480));
Q_MX02 U476 ( .S(n45), .A0(\rst_dat[9][4] ), .A1(n14), .Z(n481));
Q_MX02 U477 ( .S(n45), .A0(\rst_dat[9][5] ), .A1(n15), .Z(n482));
Q_MX02 U478 ( .S(n45), .A0(\rst_dat[9][6] ), .A1(n16), .Z(n483));
Q_MX02 U479 ( .S(n45), .A0(\rst_dat[9][7] ), .A1(n17), .Z(n484));
Q_MX02 U480 ( .S(n45), .A0(\rst_dat[9][8] ), .A1(n18), .Z(n485));
Q_MX02 U481 ( .S(n45), .A0(\rst_dat[9][9] ), .A1(n19), .Z(n486));
Q_MX02 U482 ( .S(n45), .A0(\rst_dat[9][10] ), .A1(n20), .Z(n487));
Q_MX02 U483 ( .S(n45), .A0(\rst_dat[9][11] ), .A1(n21), .Z(n488));
Q_MX02 U484 ( .S(n45), .A0(\rst_dat[9][12] ), .A1(n22), .Z(n489));
Q_MX02 U485 ( .S(n45), .A0(\rst_dat[9][13] ), .A1(n23), .Z(n490));
Q_MX02 U486 ( .S(n45), .A0(\rst_dat[9][14] ), .A1(n24), .Z(n491));
Q_MX02 U487 ( .S(n45), .A0(\rst_dat[9][15] ), .A1(n25), .Z(n492));
Q_MX02 U488 ( .S(n45), .A0(\rst_dat[9][16] ), .A1(n26), .Z(n493));
Q_MX02 U489 ( .S(n45), .A0(\rst_dat[9][17] ), .A1(n27), .Z(n494));
Q_MX02 U490 ( .S(n45), .A0(\rst_dat[9][18] ), .A1(n28), .Z(n495));
Q_MX02 U491 ( .S(n45), .A0(\rst_dat[9][19] ), .A1(n29), .Z(n496));
Q_MX02 U492 ( .S(n45), .A0(\rst_dat[9][20] ), .A1(n30), .Z(n497));
Q_MX02 U493 ( .S(n45), .A0(\rst_dat[9][21] ), .A1(n31), .Z(n498));
Q_MX02 U494 ( .S(n45), .A0(\rst_dat[9][22] ), .A1(n32), .Z(n499));
Q_MX02 U495 ( .S(n45), .A0(\rst_dat[9][23] ), .A1(n33), .Z(n500));
Q_MX02 U496 ( .S(n45), .A0(\rst_dat[9][24] ), .A1(n34), .Z(n501));
Q_MX02 U497 ( .S(n45), .A0(\rst_dat[9][25] ), .A1(n35), .Z(n502));
Q_MX02 U498 ( .S(n45), .A0(\rst_dat[9][26] ), .A1(n36), .Z(n503));
Q_MX02 U499 ( .S(n45), .A0(\rst_dat[9][27] ), .A1(n37), .Z(n504));
Q_MX02 U500 ( .S(n45), .A0(\rst_dat[9][28] ), .A1(n38), .Z(n505));
Q_MX02 U501 ( .S(n45), .A0(\rst_dat[9][29] ), .A1(n39), .Z(n506));
Q_MX02 U502 ( .S(n45), .A0(\rst_dat[9][30] ), .A1(n40), .Z(n507));
Q_MX02 U503 ( .S(n45), .A0(\rst_dat[9][31] ), .A1(n41), .Z(n508));
Q_MX02 U504 ( .S(n45), .A0(\rst_dat[10][0] ), .A1(n10), .Z(n510));
Q_MX02 U505 ( .S(n45), .A0(\rst_dat[10][1] ), .A1(n11), .Z(n511));
Q_MX02 U506 ( .S(n45), .A0(\rst_dat[10][2] ), .A1(n12), .Z(n512));
Q_MX02 U507 ( .S(n45), .A0(\rst_dat[10][3] ), .A1(n13), .Z(n513));
Q_MX02 U508 ( .S(n45), .A0(\rst_dat[10][4] ), .A1(n14), .Z(n514));
Q_MX02 U509 ( .S(n45), .A0(\rst_dat[10][5] ), .A1(n15), .Z(n515));
Q_MX02 U510 ( .S(n45), .A0(\rst_dat[10][6] ), .A1(n16), .Z(n516));
Q_MX02 U511 ( .S(n45), .A0(\rst_dat[10][7] ), .A1(n17), .Z(n517));
Q_MX02 U512 ( .S(n45), .A0(\rst_dat[10][8] ), .A1(n18), .Z(n518));
Q_MX02 U513 ( .S(n45), .A0(\rst_dat[10][9] ), .A1(n19), .Z(n519));
Q_MX02 U514 ( .S(n45), .A0(\rst_dat[10][10] ), .A1(n20), .Z(n520));
Q_MX02 U515 ( .S(n45), .A0(\rst_dat[10][11] ), .A1(n21), .Z(n521));
Q_MX02 U516 ( .S(n45), .A0(\rst_dat[10][12] ), .A1(n22), .Z(n522));
Q_MX02 U517 ( .S(n45), .A0(\rst_dat[10][13] ), .A1(n23), .Z(n523));
Q_MX02 U518 ( .S(n45), .A0(\rst_dat[10][14] ), .A1(n24), .Z(n524));
Q_MX02 U519 ( .S(n45), .A0(\rst_dat[10][15] ), .A1(n25), .Z(n525));
Q_MX02 U520 ( .S(n45), .A0(\rst_dat[10][16] ), .A1(n26), .Z(n526));
Q_MX02 U521 ( .S(n45), .A0(\rst_dat[10][17] ), .A1(n27), .Z(n527));
Q_MX02 U522 ( .S(n45), .A0(\rst_dat[10][18] ), .A1(n28), .Z(n528));
Q_MX02 U523 ( .S(n45), .A0(\rst_dat[10][19] ), .A1(n29), .Z(n529));
Q_MX02 U524 ( .S(n45), .A0(\rst_dat[10][20] ), .A1(n30), .Z(n530));
Q_MX02 U525 ( .S(n45), .A0(\rst_dat[10][21] ), .A1(n31), .Z(n531));
Q_MX02 U526 ( .S(n45), .A0(\rst_dat[10][22] ), .A1(n32), .Z(n532));
Q_MX02 U527 ( .S(n45), .A0(\rst_dat[10][23] ), .A1(n33), .Z(n533));
Q_MX02 U528 ( .S(n45), .A0(\rst_dat[10][24] ), .A1(n34), .Z(n534));
Q_MX02 U529 ( .S(n45), .A0(\rst_dat[10][25] ), .A1(n35), .Z(n535));
Q_MX02 U530 ( .S(n45), .A0(\rst_dat[10][26] ), .A1(n36), .Z(n536));
Q_MX02 U531 ( .S(n45), .A0(\rst_dat[10][27] ), .A1(n37), .Z(n537));
Q_MX02 U532 ( .S(n45), .A0(\rst_dat[10][28] ), .A1(n38), .Z(n538));
Q_MX02 U533 ( .S(n45), .A0(\rst_dat[10][29] ), .A1(n39), .Z(n539));
Q_MX02 U534 ( .S(n45), .A0(\rst_dat[10][30] ), .A1(n40), .Z(n540));
Q_MX02 U535 ( .S(n45), .A0(\rst_dat[10][31] ), .A1(n41), .Z(n541));
Q_MX02 U536 ( .S(n45), .A0(\rst_dat[11][0] ), .A1(n10), .Z(n543));
Q_MX02 U537 ( .S(n45), .A0(\rst_dat[11][1] ), .A1(n11), .Z(n544));
Q_MX02 U538 ( .S(n45), .A0(\rst_dat[11][2] ), .A1(n12), .Z(n545));
Q_MX02 U539 ( .S(n45), .A0(\rst_dat[11][3] ), .A1(n13), .Z(n546));
Q_MX02 U540 ( .S(n45), .A0(\rst_dat[11][4] ), .A1(n14), .Z(n547));
Q_MX02 U541 ( .S(n45), .A0(\rst_dat[11][5] ), .A1(n15), .Z(n548));
Q_MX02 U542 ( .S(n45), .A0(\rst_dat[11][6] ), .A1(n16), .Z(n549));
Q_MX02 U543 ( .S(n45), .A0(\rst_dat[11][7] ), .A1(n17), .Z(n550));
Q_MX02 U544 ( .S(n45), .A0(\rst_dat[11][8] ), .A1(n18), .Z(n551));
Q_MX02 U545 ( .S(n45), .A0(\rst_dat[11][9] ), .A1(n19), .Z(n552));
Q_MX02 U546 ( .S(n45), .A0(\rst_dat[11][10] ), .A1(n20), .Z(n553));
Q_MX02 U547 ( .S(n45), .A0(\rst_dat[11][11] ), .A1(n21), .Z(n554));
Q_MX02 U548 ( .S(n45), .A0(\rst_dat[11][12] ), .A1(n22), .Z(n555));
Q_MX02 U549 ( .S(n45), .A0(\rst_dat[11][13] ), .A1(n23), .Z(n556));
Q_MX02 U550 ( .S(n45), .A0(\rst_dat[11][14] ), .A1(n24), .Z(n557));
Q_MX02 U551 ( .S(n45), .A0(\rst_dat[11][15] ), .A1(n25), .Z(n558));
Q_MX02 U552 ( .S(n45), .A0(\rst_dat[11][16] ), .A1(n26), .Z(n559));
Q_MX02 U553 ( .S(n45), .A0(\rst_dat[11][17] ), .A1(n27), .Z(n560));
Q_MX02 U554 ( .S(n45), .A0(\rst_dat[11][18] ), .A1(n28), .Z(n561));
Q_MX02 U555 ( .S(n45), .A0(\rst_dat[11][19] ), .A1(n29), .Z(n562));
Q_MX02 U556 ( .S(n45), .A0(\rst_dat[11][20] ), .A1(n30), .Z(n563));
Q_MX02 U557 ( .S(n45), .A0(\rst_dat[11][21] ), .A1(n31), .Z(n564));
Q_MX02 U558 ( .S(n45), .A0(\rst_dat[11][22] ), .A1(n32), .Z(n565));
Q_MX02 U559 ( .S(n45), .A0(\rst_dat[11][23] ), .A1(n33), .Z(n566));
Q_MX02 U560 ( .S(n45), .A0(\rst_dat[11][24] ), .A1(n34), .Z(n567));
Q_MX02 U561 ( .S(n45), .A0(\rst_dat[11][25] ), .A1(n35), .Z(n568));
Q_MX02 U562 ( .S(n45), .A0(\rst_dat[11][26] ), .A1(n36), .Z(n569));
Q_MX02 U563 ( .S(n45), .A0(\rst_dat[11][27] ), .A1(n37), .Z(n570));
Q_MX02 U564 ( .S(n45), .A0(\rst_dat[11][28] ), .A1(n38), .Z(n571));
Q_MX02 U565 ( .S(n45), .A0(\rst_dat[11][29] ), .A1(n39), .Z(n572));
Q_MX02 U566 ( .S(n45), .A0(\rst_dat[11][30] ), .A1(n40), .Z(n573));
Q_MX02 U567 ( .S(n45), .A0(\rst_dat[11][31] ), .A1(n41), .Z(n574));
Q_MX02 U568 ( .S(n45), .A0(\rst_dat[12][0] ), .A1(n10), .Z(n576));
Q_MX02 U569 ( .S(n45), .A0(\rst_dat[12][1] ), .A1(n11), .Z(n577));
Q_MX02 U570 ( .S(n45), .A0(\rst_dat[12][2] ), .A1(n12), .Z(n578));
Q_MX02 U571 ( .S(n45), .A0(\rst_dat[12][3] ), .A1(n13), .Z(n579));
Q_MX02 U572 ( .S(n45), .A0(\rst_dat[12][4] ), .A1(n14), .Z(n580));
Q_MX02 U573 ( .S(n45), .A0(\rst_dat[12][5] ), .A1(n15), .Z(n581));
Q_MX02 U574 ( .S(n45), .A0(\rst_dat[12][6] ), .A1(n16), .Z(n582));
Q_MX02 U575 ( .S(n45), .A0(\rst_dat[12][7] ), .A1(n17), .Z(n583));
Q_MX02 U576 ( .S(n45), .A0(\rst_dat[12][8] ), .A1(n18), .Z(n584));
Q_MX02 U577 ( .S(n45), .A0(\rst_dat[12][9] ), .A1(n19), .Z(n585));
Q_MX02 U578 ( .S(n45), .A0(\rst_dat[12][10] ), .A1(n20), .Z(n586));
Q_MX02 U579 ( .S(n45), .A0(\rst_dat[12][11] ), .A1(n21), .Z(n587));
Q_MX02 U580 ( .S(n45), .A0(\rst_dat[12][12] ), .A1(n22), .Z(n588));
Q_MX02 U581 ( .S(n45), .A0(\rst_dat[12][13] ), .A1(n23), .Z(n589));
Q_MX02 U582 ( .S(n45), .A0(\rst_dat[12][14] ), .A1(n24), .Z(n590));
Q_MX02 U583 ( .S(n45), .A0(\rst_dat[12][15] ), .A1(n25), .Z(n591));
Q_MX02 U584 ( .S(n45), .A0(\rst_dat[12][16] ), .A1(n26), .Z(n592));
Q_MX02 U585 ( .S(n45), .A0(\rst_dat[12][17] ), .A1(n27), .Z(n593));
Q_MX02 U586 ( .S(n45), .A0(\rst_dat[12][18] ), .A1(n28), .Z(n594));
Q_MX02 U587 ( .S(n45), .A0(\rst_dat[12][19] ), .A1(n29), .Z(n595));
Q_MX02 U588 ( .S(n45), .A0(\rst_dat[12][20] ), .A1(n30), .Z(n596));
Q_MX02 U589 ( .S(n45), .A0(\rst_dat[12][21] ), .A1(n31), .Z(n597));
Q_MX02 U590 ( .S(n45), .A0(\rst_dat[12][22] ), .A1(n32), .Z(n598));
Q_MX02 U591 ( .S(n45), .A0(\rst_dat[12][23] ), .A1(n33), .Z(n599));
Q_MX02 U592 ( .S(n45), .A0(\rst_dat[12][24] ), .A1(n34), .Z(n600));
Q_MX02 U593 ( .S(n45), .A0(\rst_dat[12][25] ), .A1(n35), .Z(n601));
Q_MX02 U594 ( .S(n45), .A0(\rst_dat[12][26] ), .A1(n36), .Z(n602));
Q_MX02 U595 ( .S(n45), .A0(\rst_dat[12][27] ), .A1(n37), .Z(n603));
Q_MX02 U596 ( .S(n45), .A0(\rst_dat[12][28] ), .A1(n38), .Z(n604));
Q_MX02 U597 ( .S(n45), .A0(\rst_dat[12][29] ), .A1(n39), .Z(n605));
Q_MX02 U598 ( .S(n45), .A0(\rst_dat[12][30] ), .A1(n40), .Z(n606));
Q_MX02 U599 ( .S(n45), .A0(\rst_dat[12][31] ), .A1(n41), .Z(n607));
Q_MX02 U600 ( .S(n45), .A0(\rst_dat[13][0] ), .A1(n10), .Z(n609));
Q_MX02 U601 ( .S(n45), .A0(\rst_dat[13][1] ), .A1(n11), .Z(n610));
Q_MX02 U602 ( .S(n45), .A0(\rst_dat[13][2] ), .A1(n12), .Z(n611));
Q_MX02 U603 ( .S(n45), .A0(\rst_dat[13][3] ), .A1(n13), .Z(n612));
Q_MX02 U604 ( .S(n45), .A0(\rst_dat[13][4] ), .A1(n14), .Z(n613));
Q_MX02 U605 ( .S(n45), .A0(\rst_dat[13][5] ), .A1(n15), .Z(n614));
Q_MX02 U606 ( .S(n45), .A0(\rst_dat[13][6] ), .A1(n16), .Z(n615));
Q_MX02 U607 ( .S(n45), .A0(\rst_dat[13][7] ), .A1(n17), .Z(n616));
Q_MX02 U608 ( .S(n45), .A0(\rst_dat[13][8] ), .A1(n18), .Z(n617));
Q_MX02 U609 ( .S(n45), .A0(\rst_dat[13][9] ), .A1(n19), .Z(n618));
Q_MX02 U610 ( .S(n45), .A0(\rst_dat[13][10] ), .A1(n20), .Z(n619));
Q_MX02 U611 ( .S(n45), .A0(\rst_dat[13][11] ), .A1(n21), .Z(n620));
Q_MX02 U612 ( .S(n45), .A0(\rst_dat[13][12] ), .A1(n22), .Z(n621));
Q_MX02 U613 ( .S(n45), .A0(\rst_dat[13][13] ), .A1(n23), .Z(n622));
Q_MX02 U614 ( .S(n45), .A0(\rst_dat[13][14] ), .A1(n24), .Z(n623));
Q_MX02 U615 ( .S(n45), .A0(\rst_dat[13][15] ), .A1(n25), .Z(n624));
Q_MX02 U616 ( .S(n45), .A0(\rst_dat[13][16] ), .A1(n26), .Z(n625));
Q_MX02 U617 ( .S(n45), .A0(\rst_dat[13][17] ), .A1(n27), .Z(n626));
Q_MX02 U618 ( .S(n45), .A0(\rst_dat[13][18] ), .A1(n28), .Z(n627));
Q_MX02 U619 ( .S(n45), .A0(\rst_dat[13][19] ), .A1(n29), .Z(n628));
Q_MX02 U620 ( .S(n45), .A0(\rst_dat[13][20] ), .A1(n30), .Z(n629));
Q_MX02 U621 ( .S(n45), .A0(\rst_dat[13][21] ), .A1(n31), .Z(n630));
Q_MX02 U622 ( .S(n45), .A0(\rst_dat[13][22] ), .A1(n32), .Z(n631));
Q_MX02 U623 ( .S(n45), .A0(\rst_dat[13][23] ), .A1(n33), .Z(n632));
Q_MX02 U624 ( .S(n45), .A0(\rst_dat[13][24] ), .A1(n34), .Z(n633));
Q_MX02 U625 ( .S(n45), .A0(\rst_dat[13][25] ), .A1(n35), .Z(n634));
Q_MX02 U626 ( .S(n45), .A0(\rst_dat[13][26] ), .A1(n36), .Z(n635));
Q_MX02 U627 ( .S(n45), .A0(\rst_dat[13][27] ), .A1(n37), .Z(n636));
Q_MX02 U628 ( .S(n45), .A0(\rst_dat[13][28] ), .A1(n38), .Z(n637));
Q_MX02 U629 ( .S(n45), .A0(\rst_dat[13][29] ), .A1(n39), .Z(n638));
Q_MX02 U630 ( .S(n45), .A0(\rst_dat[13][30] ), .A1(n40), .Z(n639));
Q_MX02 U631 ( .S(n45), .A0(\rst_dat[13][31] ), .A1(n41), .Z(n640));
Q_MX02 U632 ( .S(n45), .A0(\rst_dat[14][0] ), .A1(n10), .Z(n642));
Q_MX02 U633 ( .S(n45), .A0(\rst_dat[14][1] ), .A1(n11), .Z(n643));
Q_MX02 U634 ( .S(n45), .A0(\rst_dat[14][2] ), .A1(n12), .Z(n644));
Q_MX02 U635 ( .S(n45), .A0(\rst_dat[14][3] ), .A1(n13), .Z(n645));
Q_MX02 U636 ( .S(n45), .A0(\rst_dat[14][4] ), .A1(n14), .Z(n646));
Q_MX02 U637 ( .S(n45), .A0(\rst_dat[14][5] ), .A1(n15), .Z(n647));
Q_MX02 U638 ( .S(n45), .A0(\rst_dat[14][6] ), .A1(n16), .Z(n648));
Q_MX02 U639 ( .S(n45), .A0(\rst_dat[14][7] ), .A1(n17), .Z(n649));
Q_MX02 U640 ( .S(n45), .A0(\rst_dat[14][8] ), .A1(n18), .Z(n650));
Q_MX02 U641 ( .S(n45), .A0(\rst_dat[14][9] ), .A1(n19), .Z(n651));
Q_MX02 U642 ( .S(n45), .A0(\rst_dat[14][10] ), .A1(n20), .Z(n652));
Q_MX02 U643 ( .S(n45), .A0(\rst_dat[14][11] ), .A1(n21), .Z(n653));
Q_MX02 U644 ( .S(n45), .A0(\rst_dat[14][12] ), .A1(n22), .Z(n654));
Q_MX02 U645 ( .S(n45), .A0(\rst_dat[14][13] ), .A1(n23), .Z(n655));
Q_MX02 U646 ( .S(n45), .A0(\rst_dat[14][14] ), .A1(n24), .Z(n656));
Q_MX02 U647 ( .S(n45), .A0(\rst_dat[14][15] ), .A1(n25), .Z(n657));
Q_MX02 U648 ( .S(n45), .A0(\rst_dat[14][16] ), .A1(n26), .Z(n658));
Q_MX02 U649 ( .S(n45), .A0(\rst_dat[14][17] ), .A1(n27), .Z(n659));
Q_MX02 U650 ( .S(n45), .A0(\rst_dat[14][18] ), .A1(n28), .Z(n660));
Q_MX02 U651 ( .S(n45), .A0(\rst_dat[14][19] ), .A1(n29), .Z(n661));
Q_MX02 U652 ( .S(n45), .A0(\rst_dat[14][20] ), .A1(n30), .Z(n662));
Q_MX02 U653 ( .S(n45), .A0(\rst_dat[14][21] ), .A1(n31), .Z(n663));
Q_MX02 U654 ( .S(n45), .A0(\rst_dat[14][22] ), .A1(n32), .Z(n664));
Q_MX02 U655 ( .S(n45), .A0(\rst_dat[14][23] ), .A1(n33), .Z(n665));
Q_MX02 U656 ( .S(n45), .A0(\rst_dat[14][24] ), .A1(n34), .Z(n666));
Q_MX02 U657 ( .S(n45), .A0(\rst_dat[14][25] ), .A1(n35), .Z(n667));
Q_MX02 U658 ( .S(n45), .A0(\rst_dat[14][26] ), .A1(n36), .Z(n668));
Q_MX02 U659 ( .S(n45), .A0(\rst_dat[14][27] ), .A1(n37), .Z(n669));
Q_MX02 U660 ( .S(n45), .A0(\rst_dat[14][28] ), .A1(n38), .Z(n670));
Q_MX02 U661 ( .S(n45), .A0(\rst_dat[14][29] ), .A1(n39), .Z(n671));
Q_MX02 U662 ( .S(n45), .A0(\rst_dat[14][30] ), .A1(n40), .Z(n672));
Q_MX02 U663 ( .S(n45), .A0(\rst_dat[14][31] ), .A1(n41), .Z(n673));
Q_MX02 U664 ( .S(n45), .A0(\rst_dat[15][0] ), .A1(n10), .Z(n675));
Q_MX02 U665 ( .S(n45), .A0(\rst_dat[15][1] ), .A1(n11), .Z(n676));
Q_MX02 U666 ( .S(n45), .A0(\rst_dat[15][2] ), .A1(n12), .Z(n677));
Q_MX02 U667 ( .S(n45), .A0(\rst_dat[15][3] ), .A1(n13), .Z(n678));
Q_MX02 U668 ( .S(n45), .A0(\rst_dat[15][4] ), .A1(n14), .Z(n679));
Q_MX02 U669 ( .S(n45), .A0(\rst_dat[15][5] ), .A1(n15), .Z(n680));
Q_MX02 U670 ( .S(n45), .A0(\rst_dat[15][6] ), .A1(n16), .Z(n681));
Q_MX02 U671 ( .S(n45), .A0(\rst_dat[15][7] ), .A1(n17), .Z(n682));
Q_MX02 U672 ( .S(n45), .A0(\rst_dat[15][8] ), .A1(n18), .Z(n683));
Q_MX02 U673 ( .S(n45), .A0(\rst_dat[15][9] ), .A1(n19), .Z(n684));
Q_MX02 U674 ( .S(n45), .A0(\rst_dat[15][10] ), .A1(n20), .Z(n685));
Q_MX02 U675 ( .S(n45), .A0(\rst_dat[15][11] ), .A1(n21), .Z(n686));
Q_MX02 U676 ( .S(n45), .A0(\rst_dat[15][12] ), .A1(n22), .Z(n687));
Q_MX02 U677 ( .S(n45), .A0(\rst_dat[15][13] ), .A1(n23), .Z(n688));
Q_MX02 U678 ( .S(n45), .A0(\rst_dat[15][14] ), .A1(n24), .Z(n689));
Q_MX02 U679 ( .S(n45), .A0(\rst_dat[15][15] ), .A1(n25), .Z(n690));
Q_MX02 U680 ( .S(n45), .A0(\rst_dat[15][16] ), .A1(n26), .Z(n691));
Q_MX02 U681 ( .S(n45), .A0(\rst_dat[15][17] ), .A1(n27), .Z(n692));
Q_MX02 U682 ( .S(n45), .A0(\rst_dat[15][18] ), .A1(n28), .Z(n693));
Q_MX02 U683 ( .S(n45), .A0(\rst_dat[15][19] ), .A1(n29), .Z(n694));
Q_MX02 U684 ( .S(n45), .A0(\rst_dat[15][20] ), .A1(n30), .Z(n695));
Q_MX02 U685 ( .S(n45), .A0(\rst_dat[15][21] ), .A1(n31), .Z(n696));
Q_MX02 U686 ( .S(n45), .A0(\rst_dat[15][22] ), .A1(n32), .Z(n697));
Q_MX02 U687 ( .S(n45), .A0(\rst_dat[15][23] ), .A1(n33), .Z(n698));
Q_MX02 U688 ( .S(n45), .A0(\rst_dat[15][24] ), .A1(n34), .Z(n699));
Q_MX02 U689 ( .S(n45), .A0(\rst_dat[15][25] ), .A1(n35), .Z(n700));
Q_MX02 U690 ( .S(n45), .A0(\rst_dat[15][26] ), .A1(n36), .Z(n701));
Q_MX02 U691 ( .S(n45), .A0(\rst_dat[15][27] ), .A1(n37), .Z(n702));
Q_MX02 U692 ( .S(n45), .A0(\rst_dat[15][28] ), .A1(n38), .Z(n703));
Q_MX02 U693 ( .S(n45), .A0(\rst_dat[15][29] ), .A1(n39), .Z(n704));
Q_MX02 U694 ( .S(n45), .A0(\rst_dat[15][30] ), .A1(n40), .Z(n705));
Q_MX02 U695 ( .S(n45), .A0(\rst_dat[15][31] ), .A1(n41), .Z(n706));
Q_MX02 U696 ( .S(n45), .A0(\rst_dat[16][0] ), .A1(n10), .Z(n708));
Q_MX02 U697 ( .S(n45), .A0(\rst_dat[16][1] ), .A1(n11), .Z(n709));
Q_MX02 U698 ( .S(n45), .A0(\rst_dat[16][2] ), .A1(n12), .Z(n710));
Q_MX02 U699 ( .S(n45), .A0(\rst_dat[16][3] ), .A1(n13), .Z(n711));
Q_MX02 U700 ( .S(n45), .A0(\rst_dat[16][4] ), .A1(n14), .Z(n712));
Q_MX02 U701 ( .S(n45), .A0(\rst_dat[16][5] ), .A1(n15), .Z(n713));
Q_MX02 U702 ( .S(n45), .A0(\rst_dat[16][6] ), .A1(n16), .Z(n714));
Q_MX02 U703 ( .S(n45), .A0(\rst_dat[16][7] ), .A1(n17), .Z(n715));
Q_MX02 U704 ( .S(n45), .A0(\rst_dat[16][8] ), .A1(n18), .Z(n716));
Q_MX02 U705 ( .S(n45), .A0(\rst_dat[16][9] ), .A1(n19), .Z(n717));
Q_MX02 U706 ( .S(n45), .A0(\rst_dat[16][10] ), .A1(n20), .Z(n718));
Q_MX02 U707 ( .S(n45), .A0(\rst_dat[16][11] ), .A1(n21), .Z(n719));
Q_MX02 U708 ( .S(n45), .A0(\rst_dat[16][12] ), .A1(n22), .Z(n720));
Q_MX02 U709 ( .S(n45), .A0(\rst_dat[16][13] ), .A1(n23), .Z(n721));
Q_MX02 U710 ( .S(n45), .A0(\rst_dat[16][14] ), .A1(n24), .Z(n722));
Q_MX02 U711 ( .S(n45), .A0(\rst_dat[16][15] ), .A1(n25), .Z(n723));
Q_MX02 U712 ( .S(n45), .A0(\rst_dat[16][16] ), .A1(n26), .Z(n724));
Q_MX02 U713 ( .S(n45), .A0(\rst_dat[16][17] ), .A1(n27), .Z(n725));
Q_MX02 U714 ( .S(n45), .A0(\rst_dat[16][18] ), .A1(n28), .Z(n726));
Q_MX02 U715 ( .S(n45), .A0(\rst_dat[16][19] ), .A1(n29), .Z(n727));
Q_MX02 U716 ( .S(n45), .A0(\rst_dat[16][20] ), .A1(n30), .Z(n728));
Q_MX02 U717 ( .S(n45), .A0(\rst_dat[16][21] ), .A1(n31), .Z(n729));
Q_MX02 U718 ( .S(n45), .A0(\rst_dat[16][22] ), .A1(n32), .Z(n730));
Q_MX02 U719 ( .S(n45), .A0(\rst_dat[16][23] ), .A1(n33), .Z(n731));
Q_MX02 U720 ( .S(n45), .A0(\rst_dat[16][24] ), .A1(n34), .Z(n732));
Q_MX02 U721 ( .S(n45), .A0(\rst_dat[16][25] ), .A1(n35), .Z(n733));
Q_MX02 U722 ( .S(n45), .A0(\rst_dat[16][26] ), .A1(n36), .Z(n734));
Q_MX02 U723 ( .S(n45), .A0(\rst_dat[16][27] ), .A1(n37), .Z(n735));
Q_MX02 U724 ( .S(n45), .A0(\rst_dat[16][28] ), .A1(n38), .Z(n736));
Q_MX02 U725 ( .S(n45), .A0(\rst_dat[16][29] ), .A1(n39), .Z(n737));
Q_MX02 U726 ( .S(n45), .A0(\rst_dat[16][30] ), .A1(n40), .Z(n738));
Q_MX02 U727 ( .S(n45), .A0(\rst_dat[16][31] ), .A1(n41), .Z(n739));
Q_MX02 U728 ( .S(n45), .A0(\rst_dat[17][0] ), .A1(n10), .Z(n741));
Q_MX02 U729 ( .S(n45), .A0(\rst_dat[17][1] ), .A1(n11), .Z(n742));
Q_MX02 U730 ( .S(n45), .A0(\rst_dat[17][2] ), .A1(n12), .Z(n743));
Q_MX02 U731 ( .S(n45), .A0(\rst_dat[17][3] ), .A1(n13), .Z(n744));
Q_MX02 U732 ( .S(n45), .A0(\rst_dat[17][4] ), .A1(n14), .Z(n745));
Q_MX02 U733 ( .S(n45), .A0(\rst_dat[17][5] ), .A1(n15), .Z(n746));
Q_MX02 U734 ( .S(n45), .A0(\rst_dat[17][6] ), .A1(n16), .Z(n747));
Q_MX02 U735 ( .S(n45), .A0(\rst_dat[17][7] ), .A1(n17), .Z(n748));
Q_MX02 U736 ( .S(n45), .A0(\rst_dat[17][8] ), .A1(n18), .Z(n749));
Q_MX02 U737 ( .S(n45), .A0(\rst_dat[17][9] ), .A1(n19), .Z(n750));
Q_MX02 U738 ( .S(n45), .A0(\rst_dat[17][10] ), .A1(n20), .Z(n751));
Q_MX02 U739 ( .S(n45), .A0(\rst_dat[17][11] ), .A1(n21), .Z(n752));
Q_MX02 U740 ( .S(n45), .A0(\rst_dat[17][12] ), .A1(n22), .Z(n753));
Q_MX02 U741 ( .S(n45), .A0(\rst_dat[17][13] ), .A1(n23), .Z(n754));
Q_MX02 U742 ( .S(n45), .A0(\rst_dat[17][14] ), .A1(n24), .Z(n755));
Q_MX02 U743 ( .S(n45), .A0(\rst_dat[17][15] ), .A1(n25), .Z(n756));
Q_MX02 U744 ( .S(n45), .A0(\rst_dat[17][16] ), .A1(n26), .Z(n757));
Q_MX02 U745 ( .S(n45), .A0(\rst_dat[17][17] ), .A1(n27), .Z(n758));
Q_MX02 U746 ( .S(n45), .A0(\rst_dat[17][18] ), .A1(n28), .Z(n759));
Q_MX02 U747 ( .S(n45), .A0(\rst_dat[17][19] ), .A1(n29), .Z(n760));
Q_MX02 U748 ( .S(n45), .A0(\rst_dat[17][20] ), .A1(n30), .Z(n761));
Q_MX02 U749 ( .S(n45), .A0(\rst_dat[17][21] ), .A1(n31), .Z(n762));
Q_MX02 U750 ( .S(n45), .A0(\rst_dat[17][22] ), .A1(n32), .Z(n763));
Q_MX02 U751 ( .S(n45), .A0(\rst_dat[17][23] ), .A1(n33), .Z(n764));
Q_MX02 U752 ( .S(n45), .A0(\rst_dat[17][24] ), .A1(n34), .Z(n765));
Q_MX02 U753 ( .S(n45), .A0(\rst_dat[17][25] ), .A1(n35), .Z(n766));
Q_MX02 U754 ( .S(n45), .A0(\rst_dat[17][26] ), .A1(n36), .Z(n767));
Q_MX02 U755 ( .S(n45), .A0(\rst_dat[17][27] ), .A1(n37), .Z(n768));
Q_MX02 U756 ( .S(n45), .A0(\rst_dat[17][28] ), .A1(n38), .Z(n769));
Q_MX02 U757 ( .S(n45), .A0(\rst_dat[17][29] ), .A1(n39), .Z(n770));
Q_MX02 U758 ( .S(n45), .A0(\rst_dat[17][30] ), .A1(n40), .Z(n771));
Q_MX02 U759 ( .S(n45), .A0(\rst_dat[17][31] ), .A1(n41), .Z(n772));
Q_MX02 U760 ( .S(n45), .A0(\rst_dat[18][0] ), .A1(n10), .Z(n774));
Q_MX02 U761 ( .S(n45), .A0(\rst_dat[18][1] ), .A1(n11), .Z(n775));
Q_MX02 U762 ( .S(n45), .A0(\rst_dat[18][2] ), .A1(n12), .Z(n776));
Q_MX02 U763 ( .S(n45), .A0(\rst_dat[18][3] ), .A1(n13), .Z(n777));
Q_MX02 U764 ( .S(n45), .A0(\rst_dat[18][4] ), .A1(n14), .Z(n778));
Q_MX02 U765 ( .S(n45), .A0(\rst_dat[18][5] ), .A1(n15), .Z(n779));
Q_MX02 U766 ( .S(n45), .A0(\rst_dat[18][6] ), .A1(n16), .Z(n780));
Q_MX02 U767 ( .S(n45), .A0(\rst_dat[18][7] ), .A1(n17), .Z(n781));
Q_MX02 U768 ( .S(n45), .A0(\rst_dat[18][8] ), .A1(n18), .Z(n782));
Q_MX02 U769 ( .S(n45), .A0(\rst_dat[18][9] ), .A1(n19), .Z(n783));
Q_MX02 U770 ( .S(n45), .A0(\rst_dat[18][10] ), .A1(n20), .Z(n784));
Q_MX02 U771 ( .S(n45), .A0(\rst_dat[18][11] ), .A1(n21), .Z(n785));
Q_MX02 U772 ( .S(n45), .A0(\rst_dat[18][12] ), .A1(n22), .Z(n786));
Q_MX02 U773 ( .S(n45), .A0(\rst_dat[18][13] ), .A1(n23), .Z(n787));
Q_MX02 U774 ( .S(n45), .A0(\rst_dat[18][14] ), .A1(n24), .Z(n788));
Q_MX02 U775 ( .S(n45), .A0(\rst_dat[18][15] ), .A1(n25), .Z(n789));
Q_MX02 U776 ( .S(n45), .A0(\rst_dat[18][16] ), .A1(n26), .Z(n790));
Q_MX02 U777 ( .S(n45), .A0(\rst_dat[18][17] ), .A1(n27), .Z(n791));
Q_MX02 U778 ( .S(n45), .A0(\rst_dat[18][18] ), .A1(n28), .Z(n792));
Q_MX02 U779 ( .S(n45), .A0(\rst_dat[18][19] ), .A1(n29), .Z(n793));
Q_MX02 U780 ( .S(n45), .A0(\rst_dat[18][20] ), .A1(n30), .Z(n794));
Q_MX02 U781 ( .S(n45), .A0(\rst_dat[18][21] ), .A1(n31), .Z(n795));
Q_MX02 U782 ( .S(n45), .A0(\rst_dat[18][22] ), .A1(n32), .Z(n796));
Q_MX02 U783 ( .S(n45), .A0(\rst_dat[18][23] ), .A1(n33), .Z(n797));
Q_MX02 U784 ( .S(n45), .A0(\rst_dat[18][24] ), .A1(n34), .Z(n798));
Q_MX02 U785 ( .S(n45), .A0(\rst_dat[18][25] ), .A1(n35), .Z(n799));
Q_MX02 U786 ( .S(n45), .A0(\rst_dat[18][26] ), .A1(n36), .Z(n800));
Q_MX02 U787 ( .S(n45), .A0(\rst_dat[18][27] ), .A1(n37), .Z(n801));
Q_MX02 U788 ( .S(n45), .A0(\rst_dat[18][28] ), .A1(n38), .Z(n802));
Q_MX02 U789 ( .S(n45), .A0(\rst_dat[18][29] ), .A1(n39), .Z(n803));
Q_MX02 U790 ( .S(n45), .A0(\rst_dat[18][30] ), .A1(n40), .Z(n804));
Q_MX02 U791 ( .S(n45), .A0(\rst_dat[18][31] ), .A1(n41), .Z(n805));
Q_MX02 U792 ( .S(n45), .A0(\rst_dat[19][0] ), .A1(n10), .Z(n807));
Q_MX02 U793 ( .S(n45), .A0(\rst_dat[19][1] ), .A1(n11), .Z(n808));
Q_MX02 U794 ( .S(n45), .A0(\rst_dat[19][2] ), .A1(n12), .Z(n809));
Q_MX02 U795 ( .S(n45), .A0(\rst_dat[19][3] ), .A1(n13), .Z(n810));
Q_MX02 U796 ( .S(n45), .A0(\rst_dat[19][4] ), .A1(n14), .Z(n811));
Q_MX02 U797 ( .S(n45), .A0(\rst_dat[19][5] ), .A1(n15), .Z(n812));
Q_MX02 U798 ( .S(n45), .A0(\rst_dat[19][6] ), .A1(n16), .Z(n813));
Q_MX02 U799 ( .S(n45), .A0(\rst_dat[19][7] ), .A1(n17), .Z(n814));
Q_MX02 U800 ( .S(n45), .A0(\rst_dat[19][8] ), .A1(n18), .Z(n815));
Q_MX02 U801 ( .S(n45), .A0(\rst_dat[19][9] ), .A1(n19), .Z(n816));
Q_MX02 U802 ( .S(n45), .A0(\rst_dat[19][10] ), .A1(n20), .Z(n817));
Q_MX02 U803 ( .S(n45), .A0(\rst_dat[19][11] ), .A1(n21), .Z(n818));
Q_MX02 U804 ( .S(n45), .A0(\rst_dat[19][12] ), .A1(n22), .Z(n819));
Q_MX02 U805 ( .S(n45), .A0(\rst_dat[19][13] ), .A1(n23), .Z(n820));
Q_MX02 U806 ( .S(n45), .A0(\rst_dat[19][14] ), .A1(n24), .Z(n821));
Q_MX02 U807 ( .S(n45), .A0(\rst_dat[19][15] ), .A1(n25), .Z(n822));
Q_MX02 U808 ( .S(n45), .A0(\rst_dat[19][16] ), .A1(n26), .Z(n823));
Q_MX02 U809 ( .S(n45), .A0(\rst_dat[19][17] ), .A1(n27), .Z(n824));
Q_MX02 U810 ( .S(n45), .A0(\rst_dat[19][18] ), .A1(n28), .Z(n825));
Q_MX02 U811 ( .S(n45), .A0(\rst_dat[19][19] ), .A1(n29), .Z(n826));
Q_MX02 U812 ( .S(n45), .A0(\rst_dat[19][20] ), .A1(n30), .Z(n827));
Q_MX02 U813 ( .S(n45), .A0(\rst_dat[19][21] ), .A1(n31), .Z(n828));
Q_MX02 U814 ( .S(n45), .A0(\rst_dat[19][22] ), .A1(n32), .Z(n829));
Q_MX02 U815 ( .S(n45), .A0(\rst_dat[19][23] ), .A1(n33), .Z(n830));
Q_MX02 U816 ( .S(n45), .A0(\rst_dat[19][24] ), .A1(n34), .Z(n831));
Q_MX02 U817 ( .S(n45), .A0(\rst_dat[19][25] ), .A1(n35), .Z(n832));
Q_MX02 U818 ( .S(n45), .A0(\rst_dat[19][26] ), .A1(n36), .Z(n833));
Q_MX02 U819 ( .S(n45), .A0(\rst_dat[19][27] ), .A1(n37), .Z(n834));
Q_MX02 U820 ( .S(n45), .A0(\rst_dat[19][28] ), .A1(n38), .Z(n835));
Q_MX02 U821 ( .S(n45), .A0(\rst_dat[19][29] ), .A1(n39), .Z(n836));
Q_MX02 U822 ( .S(n45), .A0(\rst_dat[19][30] ), .A1(n40), .Z(n837));
Q_MX02 U823 ( .S(n45), .A0(\rst_dat[19][31] ), .A1(n41), .Z(n838));
Q_MX02 U824 ( .S(n45), .A0(\rst_dat[20][0] ), .A1(n10), .Z(n840));
Q_MX02 U825 ( .S(n45), .A0(\rst_dat[20][1] ), .A1(n11), .Z(n841));
Q_MX02 U826 ( .S(n45), .A0(\rst_dat[20][2] ), .A1(n12), .Z(n842));
Q_MX02 U827 ( .S(n45), .A0(\rst_dat[20][3] ), .A1(n13), .Z(n843));
Q_MX02 U828 ( .S(n45), .A0(\rst_dat[20][4] ), .A1(n14), .Z(n844));
Q_MX02 U829 ( .S(n45), .A0(\rst_dat[20][5] ), .A1(n15), .Z(n845));
Q_MX02 U830 ( .S(n45), .A0(\rst_dat[20][6] ), .A1(n16), .Z(n846));
Q_MX02 U831 ( .S(n45), .A0(\rst_dat[20][7] ), .A1(n17), .Z(n847));
Q_MX02 U832 ( .S(n45), .A0(\rst_dat[20][8] ), .A1(n18), .Z(n848));
Q_MX02 U833 ( .S(n45), .A0(\rst_dat[20][9] ), .A1(n19), .Z(n849));
Q_MX02 U834 ( .S(n45), .A0(\rst_dat[20][10] ), .A1(n20), .Z(n850));
Q_MX02 U835 ( .S(n45), .A0(\rst_dat[20][11] ), .A1(n21), .Z(n851));
Q_MX02 U836 ( .S(n45), .A0(\rst_dat[20][12] ), .A1(n22), .Z(n852));
Q_MX02 U837 ( .S(n45), .A0(\rst_dat[20][13] ), .A1(n23), .Z(n853));
Q_MX02 U838 ( .S(n45), .A0(\rst_dat[20][14] ), .A1(n24), .Z(n854));
Q_MX02 U839 ( .S(n45), .A0(\rst_dat[20][15] ), .A1(n25), .Z(n855));
Q_MX02 U840 ( .S(n45), .A0(\rst_dat[20][16] ), .A1(n26), .Z(n856));
Q_MX02 U841 ( .S(n45), .A0(\rst_dat[20][17] ), .A1(n27), .Z(n857));
Q_MX02 U842 ( .S(n45), .A0(\rst_dat[20][18] ), .A1(n28), .Z(n858));
Q_MX02 U843 ( .S(n45), .A0(\rst_dat[20][19] ), .A1(n29), .Z(n859));
Q_MX02 U844 ( .S(n45), .A0(\rst_dat[20][20] ), .A1(n30), .Z(n860));
Q_MX02 U845 ( .S(n45), .A0(\rst_dat[20][21] ), .A1(n31), .Z(n861));
Q_MX02 U846 ( .S(n45), .A0(\rst_dat[20][22] ), .A1(n32), .Z(n862));
Q_MX02 U847 ( .S(n45), .A0(\rst_dat[20][23] ), .A1(n33), .Z(n863));
Q_MX02 U848 ( .S(n45), .A0(\rst_dat[20][24] ), .A1(n34), .Z(n864));
Q_MX02 U849 ( .S(n45), .A0(\rst_dat[20][25] ), .A1(n35), .Z(n865));
Q_MX02 U850 ( .S(n45), .A0(\rst_dat[20][26] ), .A1(n36), .Z(n866));
Q_MX02 U851 ( .S(n45), .A0(\rst_dat[20][27] ), .A1(n37), .Z(n867));
Q_MX02 U852 ( .S(n45), .A0(\rst_dat[20][28] ), .A1(n38), .Z(n868));
Q_MX02 U853 ( .S(n45), .A0(\rst_dat[20][29] ), .A1(n39), .Z(n869));
Q_MX02 U854 ( .S(n45), .A0(\rst_dat[20][30] ), .A1(n40), .Z(n870));
Q_MX02 U855 ( .S(n45), .A0(\rst_dat[20][31] ), .A1(n41), .Z(n871));
Q_MX02 U856 ( .S(n45), .A0(\rst_dat[21][0] ), .A1(n10), .Z(n873));
Q_MX02 U857 ( .S(n45), .A0(\rst_dat[21][1] ), .A1(n11), .Z(n874));
Q_MX02 U858 ( .S(n45), .A0(\rst_dat[21][2] ), .A1(n12), .Z(n875));
Q_MX02 U859 ( .S(n45), .A0(\rst_dat[21][3] ), .A1(n13), .Z(n876));
Q_MX02 U860 ( .S(n45), .A0(\rst_dat[21][4] ), .A1(n14), .Z(n877));
Q_MX02 U861 ( .S(n45), .A0(\rst_dat[21][5] ), .A1(n15), .Z(n878));
Q_MX02 U862 ( .S(n45), .A0(\rst_dat[21][6] ), .A1(n16), .Z(n879));
Q_MX02 U863 ( .S(n45), .A0(\rst_dat[21][7] ), .A1(n17), .Z(n880));
Q_MX02 U864 ( .S(n45), .A0(\rst_dat[21][8] ), .A1(n18), .Z(n881));
Q_MX02 U865 ( .S(n45), .A0(\rst_dat[21][9] ), .A1(n19), .Z(n882));
Q_MX02 U866 ( .S(n45), .A0(\rst_dat[21][10] ), .A1(n20), .Z(n883));
Q_MX02 U867 ( .S(n45), .A0(\rst_dat[21][11] ), .A1(n21), .Z(n884));
Q_MX02 U868 ( .S(n45), .A0(\rst_dat[21][12] ), .A1(n22), .Z(n885));
Q_MX02 U869 ( .S(n45), .A0(\rst_dat[21][13] ), .A1(n23), .Z(n886));
Q_MX02 U870 ( .S(n45), .A0(\rst_dat[21][14] ), .A1(n24), .Z(n887));
Q_MX02 U871 ( .S(n45), .A0(\rst_dat[21][15] ), .A1(n25), .Z(n888));
Q_MX02 U872 ( .S(n45), .A0(\rst_dat[21][16] ), .A1(n26), .Z(n889));
Q_MX02 U873 ( .S(n45), .A0(\rst_dat[21][17] ), .A1(n27), .Z(n890));
Q_MX02 U874 ( .S(n45), .A0(\rst_dat[21][18] ), .A1(n28), .Z(n891));
Q_MX02 U875 ( .S(n45), .A0(\rst_dat[21][19] ), .A1(n29), .Z(n892));
Q_MX02 U876 ( .S(n45), .A0(\rst_dat[21][20] ), .A1(n30), .Z(n893));
Q_MX02 U877 ( .S(n45), .A0(\rst_dat[21][21] ), .A1(n31), .Z(n894));
Q_MX02 U878 ( .S(n45), .A0(\rst_dat[21][22] ), .A1(n32), .Z(n895));
Q_MX02 U879 ( .S(n45), .A0(\rst_dat[21][23] ), .A1(n33), .Z(n896));
Q_MX02 U880 ( .S(n45), .A0(\rst_dat[21][24] ), .A1(n34), .Z(n897));
Q_MX02 U881 ( .S(n45), .A0(\rst_dat[21][25] ), .A1(n35), .Z(n898));
Q_MX02 U882 ( .S(n45), .A0(\rst_dat[21][26] ), .A1(n36), .Z(n899));
Q_MX02 U883 ( .S(n45), .A0(\rst_dat[21][27] ), .A1(n37), .Z(n900));
Q_MX02 U884 ( .S(n45), .A0(\rst_dat[21][28] ), .A1(n38), .Z(n901));
Q_MX02 U885 ( .S(n45), .A0(\rst_dat[21][29] ), .A1(n39), .Z(n902));
Q_MX02 U886 ( .S(n45), .A0(\rst_dat[21][30] ), .A1(n40), .Z(n903));
Q_MX02 U887 ( .S(n45), .A0(\rst_dat[21][31] ), .A1(n41), .Z(n904));
Q_MX02 U888 ( .S(n45), .A0(\rst_dat[22][0] ), .A1(n10), .Z(n906));
Q_MX02 U889 ( .S(n45), .A0(\rst_dat[22][1] ), .A1(n11), .Z(n907));
Q_MX02 U890 ( .S(n45), .A0(\rst_dat[22][2] ), .A1(n12), .Z(n908));
Q_MX02 U891 ( .S(n45), .A0(\rst_dat[22][3] ), .A1(n13), .Z(n909));
Q_MX02 U892 ( .S(n45), .A0(\rst_dat[22][4] ), .A1(n14), .Z(n910));
Q_MX02 U893 ( .S(n45), .A0(\rst_dat[22][5] ), .A1(n15), .Z(n911));
Q_MX02 U894 ( .S(n45), .A0(\rst_dat[22][6] ), .A1(n16), .Z(n912));
Q_MX02 U895 ( .S(n45), .A0(\rst_dat[22][7] ), .A1(n17), .Z(n913));
Q_MX02 U896 ( .S(n45), .A0(\rst_dat[22][8] ), .A1(n18), .Z(n914));
Q_MX02 U897 ( .S(n45), .A0(\rst_dat[22][9] ), .A1(n19), .Z(n915));
Q_MX02 U898 ( .S(n45), .A0(\rst_dat[22][10] ), .A1(n20), .Z(n916));
Q_MX02 U899 ( .S(n45), .A0(\rst_dat[22][11] ), .A1(n21), .Z(n917));
Q_MX02 U900 ( .S(n45), .A0(\rst_dat[22][12] ), .A1(n22), .Z(n918));
Q_MX02 U901 ( .S(n45), .A0(\rst_dat[22][13] ), .A1(n23), .Z(n919));
Q_MX02 U902 ( .S(n45), .A0(\rst_dat[22][14] ), .A1(n24), .Z(n920));
Q_MX02 U903 ( .S(n45), .A0(\rst_dat[22][15] ), .A1(n25), .Z(n921));
Q_MX02 U904 ( .S(n45), .A0(\rst_dat[22][16] ), .A1(n26), .Z(n922));
Q_MX02 U905 ( .S(n45), .A0(\rst_dat[22][17] ), .A1(n27), .Z(n923));
Q_MX02 U906 ( .S(n45), .A0(\rst_dat[22][18] ), .A1(n28), .Z(n924));
Q_MX02 U907 ( .S(n45), .A0(\rst_dat[22][19] ), .A1(n29), .Z(n925));
Q_MX02 U908 ( .S(n45), .A0(\rst_dat[22][20] ), .A1(n30), .Z(n926));
Q_MX02 U909 ( .S(n45), .A0(\rst_dat[22][21] ), .A1(n31), .Z(n927));
Q_MX02 U910 ( .S(n45), .A0(\rst_dat[22][22] ), .A1(n32), .Z(n928));
Q_MX02 U911 ( .S(n45), .A0(\rst_dat[22][23] ), .A1(n33), .Z(n929));
Q_MX02 U912 ( .S(n45), .A0(\rst_dat[22][24] ), .A1(n34), .Z(n930));
Q_MX02 U913 ( .S(n45), .A0(\rst_dat[22][25] ), .A1(n35), .Z(n931));
Q_MX02 U914 ( .S(n45), .A0(\rst_dat[22][26] ), .A1(n36), .Z(n932));
Q_MX02 U915 ( .S(n45), .A0(\rst_dat[22][27] ), .A1(n37), .Z(n933));
Q_MX02 U916 ( .S(n45), .A0(\rst_dat[22][28] ), .A1(n38), .Z(n934));
Q_MX02 U917 ( .S(n45), .A0(\rst_dat[22][29] ), .A1(n39), .Z(n935));
Q_MX02 U918 ( .S(n45), .A0(\rst_dat[22][30] ), .A1(n40), .Z(n936));
Q_MX02 U919 ( .S(n45), .A0(\rst_dat[22][31] ), .A1(n41), .Z(n937));
Q_MX02 U920 ( .S(n45), .A0(\rst_dat[23][0] ), .A1(n10), .Z(n939));
Q_MX02 U921 ( .S(n45), .A0(\rst_dat[23][1] ), .A1(n11), .Z(n940));
Q_MX02 U922 ( .S(n45), .A0(\rst_dat[23][2] ), .A1(n12), .Z(n941));
Q_MX02 U923 ( .S(n45), .A0(\rst_dat[23][3] ), .A1(n13), .Z(n942));
Q_MX02 U924 ( .S(n45), .A0(\rst_dat[23][4] ), .A1(n14), .Z(n943));
Q_MX02 U925 ( .S(n45), .A0(\rst_dat[23][5] ), .A1(n15), .Z(n944));
Q_MX02 U926 ( .S(n45), .A0(\rst_dat[23][6] ), .A1(n16), .Z(n945));
Q_MX02 U927 ( .S(n45), .A0(\rst_dat[23][7] ), .A1(n17), .Z(n946));
Q_MX02 U928 ( .S(n45), .A0(\rst_dat[23][8] ), .A1(n18), .Z(n947));
Q_MX02 U929 ( .S(n45), .A0(\rst_dat[23][9] ), .A1(n19), .Z(n948));
Q_MX02 U930 ( .S(n45), .A0(\rst_dat[23][10] ), .A1(n20), .Z(n949));
Q_MX02 U931 ( .S(n45), .A0(\rst_dat[23][11] ), .A1(n21), .Z(n950));
Q_MX02 U932 ( .S(n45), .A0(\rst_dat[23][12] ), .A1(n22), .Z(n951));
Q_MX02 U933 ( .S(n45), .A0(\rst_dat[23][13] ), .A1(n23), .Z(n952));
Q_MX02 U934 ( .S(n45), .A0(\rst_dat[23][14] ), .A1(n24), .Z(n953));
Q_MX02 U935 ( .S(n45), .A0(\rst_dat[23][15] ), .A1(n25), .Z(n954));
Q_MX02 U936 ( .S(n45), .A0(\rst_dat[23][16] ), .A1(n26), .Z(n955));
Q_MX02 U937 ( .S(n45), .A0(\rst_dat[23][17] ), .A1(n27), .Z(n956));
Q_MX02 U938 ( .S(n45), .A0(\rst_dat[23][18] ), .A1(n28), .Z(n957));
Q_MX02 U939 ( .S(n45), .A0(\rst_dat[23][19] ), .A1(n29), .Z(n958));
Q_MX02 U940 ( .S(n45), .A0(\rst_dat[23][20] ), .A1(n30), .Z(n959));
Q_MX02 U941 ( .S(n45), .A0(\rst_dat[23][21] ), .A1(n31), .Z(n960));
Q_MX02 U942 ( .S(n45), .A0(\rst_dat[23][22] ), .A1(n32), .Z(n961));
Q_MX02 U943 ( .S(n45), .A0(\rst_dat[23][23] ), .A1(n33), .Z(n962));
Q_MX02 U944 ( .S(n45), .A0(\rst_dat[23][24] ), .A1(n34), .Z(n963));
Q_MX02 U945 ( .S(n45), .A0(\rst_dat[23][25] ), .A1(n35), .Z(n964));
Q_MX02 U946 ( .S(n45), .A0(\rst_dat[23][26] ), .A1(n36), .Z(n965));
Q_MX02 U947 ( .S(n45), .A0(\rst_dat[23][27] ), .A1(n37), .Z(n966));
Q_MX02 U948 ( .S(n45), .A0(\rst_dat[23][28] ), .A1(n38), .Z(n967));
Q_MX02 U949 ( .S(n45), .A0(\rst_dat[23][29] ), .A1(n39), .Z(n968));
Q_MX02 U950 ( .S(n45), .A0(\rst_dat[23][30] ), .A1(n40), .Z(n969));
Q_MX02 U951 ( .S(n45), .A0(\rst_dat[23][31] ), .A1(n41), .Z(n970));
Q_MX02 U952 ( .S(n45), .A0(\rst_dat[24][0] ), .A1(n10), .Z(n972));
Q_MX02 U953 ( .S(n45), .A0(\rst_dat[24][1] ), .A1(n11), .Z(n973));
Q_MX02 U954 ( .S(n45), .A0(\rst_dat[24][2] ), .A1(n12), .Z(n974));
Q_MX02 U955 ( .S(n45), .A0(\rst_dat[24][3] ), .A1(n13), .Z(n975));
Q_MX02 U956 ( .S(n45), .A0(\rst_dat[24][4] ), .A1(n14), .Z(n976));
Q_MX02 U957 ( .S(n45), .A0(\rst_dat[24][5] ), .A1(n15), .Z(n977));
Q_MX02 U958 ( .S(n45), .A0(\rst_dat[24][6] ), .A1(n16), .Z(n978));
Q_MX02 U959 ( .S(n45), .A0(\rst_dat[24][7] ), .A1(n17), .Z(n979));
Q_MX02 U960 ( .S(n45), .A0(\rst_dat[24][8] ), .A1(n18), .Z(n980));
Q_MX02 U961 ( .S(n45), .A0(\rst_dat[24][9] ), .A1(n19), .Z(n981));
Q_MX02 U962 ( .S(n45), .A0(\rst_dat[24][10] ), .A1(n20), .Z(n982));
Q_MX02 U963 ( .S(n45), .A0(\rst_dat[24][11] ), .A1(n21), .Z(n983));
Q_MX02 U964 ( .S(n45), .A0(\rst_dat[24][12] ), .A1(n22), .Z(n984));
Q_MX02 U965 ( .S(n45), .A0(\rst_dat[24][13] ), .A1(n23), .Z(n985));
Q_MX02 U966 ( .S(n45), .A0(\rst_dat[24][14] ), .A1(n24), .Z(n986));
Q_MX02 U967 ( .S(n45), .A0(\rst_dat[24][15] ), .A1(n25), .Z(n987));
Q_MX02 U968 ( .S(n45), .A0(\rst_dat[24][16] ), .A1(n26), .Z(n988));
Q_MX02 U969 ( .S(n45), .A0(\rst_dat[24][17] ), .A1(n27), .Z(n989));
Q_MX02 U970 ( .S(n45), .A0(\rst_dat[24][18] ), .A1(n28), .Z(n990));
Q_MX02 U971 ( .S(n45), .A0(\rst_dat[24][19] ), .A1(n29), .Z(n991));
Q_MX02 U972 ( .S(n45), .A0(\rst_dat[24][20] ), .A1(n30), .Z(n992));
Q_MX02 U973 ( .S(n45), .A0(\rst_dat[24][21] ), .A1(n31), .Z(n993));
Q_MX02 U974 ( .S(n45), .A0(\rst_dat[24][22] ), .A1(n32), .Z(n994));
Q_MX02 U975 ( .S(n45), .A0(\rst_dat[24][23] ), .A1(n33), .Z(n995));
Q_MX02 U976 ( .S(n45), .A0(\rst_dat[24][24] ), .A1(n34), .Z(n996));
Q_MX02 U977 ( .S(n45), .A0(\rst_dat[24][25] ), .A1(n35), .Z(n997));
Q_MX02 U978 ( .S(n45), .A0(\rst_dat[24][26] ), .A1(n36), .Z(n998));
Q_MX02 U979 ( .S(n45), .A0(\rst_dat[24][27] ), .A1(n37), .Z(n999));
Q_MX02 U980 ( .S(n45), .A0(\rst_dat[24][28] ), .A1(n38), .Z(n1000));
Q_MX02 U981 ( .S(n45), .A0(\rst_dat[24][29] ), .A1(n39), .Z(n1001));
Q_MX02 U982 ( .S(n45), .A0(\rst_dat[24][30] ), .A1(n40), .Z(n1002));
Q_MX02 U983 ( .S(n45), .A0(\rst_dat[24][31] ), .A1(n41), .Z(n1003));
Q_MX02 U984 ( .S(n45), .A0(\rst_dat[25][0] ), .A1(n10), .Z(n1005));
Q_MX02 U985 ( .S(n45), .A0(\rst_dat[25][1] ), .A1(n11), .Z(n1006));
Q_MX02 U986 ( .S(n45), .A0(\rst_dat[25][2] ), .A1(n12), .Z(n1007));
Q_MX02 U987 ( .S(n45), .A0(\rst_dat[25][3] ), .A1(n13), .Z(n1008));
Q_MX02 U988 ( .S(n45), .A0(\rst_dat[25][4] ), .A1(n14), .Z(n1009));
Q_MX02 U989 ( .S(n45), .A0(\rst_dat[25][5] ), .A1(n15), .Z(n1010));
Q_MX02 U990 ( .S(n45), .A0(\rst_dat[25][6] ), .A1(n16), .Z(n1011));
Q_MX02 U991 ( .S(n45), .A0(\rst_dat[25][7] ), .A1(n17), .Z(n1012));
Q_MX02 U992 ( .S(n45), .A0(\rst_dat[25][8] ), .A1(n18), .Z(n1013));
Q_MX02 U993 ( .S(n45), .A0(\rst_dat[25][9] ), .A1(n19), .Z(n1014));
Q_MX02 U994 ( .S(n45), .A0(\rst_dat[25][10] ), .A1(n20), .Z(n1015));
Q_MX02 U995 ( .S(n45), .A0(\rst_dat[25][11] ), .A1(n21), .Z(n1016));
Q_MX02 U996 ( .S(n45), .A0(\rst_dat[25][12] ), .A1(n22), .Z(n1017));
Q_MX02 U997 ( .S(n45), .A0(\rst_dat[25][13] ), .A1(n23), .Z(n1018));
Q_MX02 U998 ( .S(n45), .A0(\rst_dat[25][14] ), .A1(n24), .Z(n1019));
Q_MX02 U999 ( .S(n45), .A0(\rst_dat[25][15] ), .A1(n25), .Z(n1020));
Q_MX02 U1000 ( .S(n45), .A0(\rst_dat[25][16] ), .A1(n26), .Z(n1021));
Q_MX02 U1001 ( .S(n45), .A0(\rst_dat[25][17] ), .A1(n27), .Z(n1022));
Q_MX02 U1002 ( .S(n45), .A0(\rst_dat[25][18] ), .A1(n28), .Z(n1023));
Q_MX02 U1003 ( .S(n45), .A0(\rst_dat[25][19] ), .A1(n29), .Z(n1024));
Q_MX02 U1004 ( .S(n45), .A0(\rst_dat[25][20] ), .A1(n30), .Z(n1025));
Q_MX02 U1005 ( .S(n45), .A0(\rst_dat[25][21] ), .A1(n31), .Z(n1026));
Q_MX02 U1006 ( .S(n45), .A0(\rst_dat[25][22] ), .A1(n32), .Z(n1027));
Q_MX02 U1007 ( .S(n45), .A0(\rst_dat[25][23] ), .A1(n33), .Z(n1028));
Q_MX02 U1008 ( .S(n45), .A0(\rst_dat[25][24] ), .A1(n34), .Z(n1029));
Q_MX02 U1009 ( .S(n45), .A0(\rst_dat[25][25] ), .A1(n35), .Z(n1030));
Q_MX02 U1010 ( .S(n45), .A0(\rst_dat[25][26] ), .A1(n36), .Z(n1031));
Q_MX02 U1011 ( .S(n45), .A0(\rst_dat[25][27] ), .A1(n37), .Z(n1032));
Q_MX02 U1012 ( .S(n45), .A0(\rst_dat[25][28] ), .A1(n38), .Z(n1033));
Q_MX02 U1013 ( .S(n45), .A0(\rst_dat[25][29] ), .A1(n39), .Z(n1034));
Q_MX02 U1014 ( .S(n45), .A0(\rst_dat[25][30] ), .A1(n40), .Z(n1035));
Q_MX02 U1015 ( .S(n45), .A0(\rst_dat[25][31] ), .A1(n41), .Z(n1036));
Q_MX02 U1016 ( .S(n45), .A0(\rst_dat[26][0] ), .A1(n10), .Z(n1038));
Q_MX02 U1017 ( .S(n45), .A0(\rst_dat[26][1] ), .A1(n11), .Z(n1039));
Q_MX02 U1018 ( .S(n45), .A0(\rst_dat[26][2] ), .A1(n12), .Z(n1040));
Q_MX02 U1019 ( .S(n45), .A0(\rst_dat[26][3] ), .A1(n13), .Z(n1041));
Q_MX02 U1020 ( .S(n45), .A0(\rst_dat[26][4] ), .A1(n14), .Z(n1042));
Q_MX02 U1021 ( .S(n45), .A0(\rst_dat[26][5] ), .A1(n15), .Z(n1043));
Q_MX02 U1022 ( .S(n45), .A0(\rst_dat[26][6] ), .A1(n16), .Z(n1044));
Q_MX02 U1023 ( .S(n45), .A0(\rst_dat[26][7] ), .A1(n17), .Z(n1045));
Q_MX02 U1024 ( .S(n45), .A0(\rst_dat[26][8] ), .A1(n18), .Z(n1046));
Q_MX02 U1025 ( .S(n45), .A0(\rst_dat[26][9] ), .A1(n19), .Z(n1047));
Q_MX02 U1026 ( .S(n45), .A0(\rst_dat[26][10] ), .A1(n20), .Z(n1048));
Q_MX02 U1027 ( .S(n45), .A0(\rst_dat[26][11] ), .A1(n21), .Z(n1049));
Q_MX02 U1028 ( .S(n45), .A0(\rst_dat[26][12] ), .A1(n22), .Z(n1050));
Q_MX02 U1029 ( .S(n45), .A0(\rst_dat[26][13] ), .A1(n23), .Z(n1051));
Q_MX02 U1030 ( .S(n45), .A0(\rst_dat[26][14] ), .A1(n24), .Z(n1052));
Q_MX02 U1031 ( .S(n45), .A0(\rst_dat[26][15] ), .A1(n25), .Z(n1053));
Q_MX02 U1032 ( .S(n45), .A0(\rst_dat[26][16] ), .A1(n26), .Z(n1054));
Q_MX02 U1033 ( .S(n45), .A0(\rst_dat[26][17] ), .A1(n27), .Z(n1055));
Q_MX02 U1034 ( .S(n45), .A0(\rst_dat[26][18] ), .A1(n28), .Z(n1056));
Q_MX02 U1035 ( .S(n45), .A0(\rst_dat[26][19] ), .A1(n29), .Z(n1057));
Q_MX02 U1036 ( .S(n45), .A0(\rst_dat[26][20] ), .A1(n30), .Z(n1058));
Q_MX02 U1037 ( .S(n45), .A0(\rst_dat[26][21] ), .A1(n31), .Z(n1059));
Q_MX02 U1038 ( .S(n45), .A0(\rst_dat[26][22] ), .A1(n32), .Z(n1060));
Q_MX02 U1039 ( .S(n45), .A0(\rst_dat[26][23] ), .A1(n33), .Z(n1061));
Q_MX02 U1040 ( .S(n45), .A0(\rst_dat[26][24] ), .A1(n34), .Z(n1062));
Q_MX02 U1041 ( .S(n45), .A0(\rst_dat[26][25] ), .A1(n35), .Z(n1063));
Q_MX02 U1042 ( .S(n45), .A0(\rst_dat[26][26] ), .A1(n36), .Z(n1064));
Q_MX02 U1043 ( .S(n45), .A0(\rst_dat[26][27] ), .A1(n37), .Z(n1065));
Q_MX02 U1044 ( .S(n45), .A0(\rst_dat[26][28] ), .A1(n38), .Z(n1066));
Q_MX02 U1045 ( .S(n45), .A0(\rst_dat[26][29] ), .A1(n39), .Z(n1067));
Q_MX02 U1046 ( .S(n45), .A0(\rst_dat[26][30] ), .A1(n40), .Z(n1068));
Q_MX02 U1047 ( .S(n45), .A0(\rst_dat[26][31] ), .A1(n41), .Z(n1069));
Q_MX02 U1048 ( .S(n45), .A0(\rst_dat[27][0] ), .A1(n10), .Z(n1071));
Q_MX02 U1049 ( .S(n45), .A0(\rst_dat[27][1] ), .A1(n11), .Z(n1072));
Q_MX02 U1050 ( .S(n45), .A0(\rst_dat[27][2] ), .A1(n12), .Z(n1073));
Q_MX02 U1051 ( .S(n45), .A0(\rst_dat[27][3] ), .A1(n13), .Z(n1074));
Q_MX02 U1052 ( .S(n45), .A0(\rst_dat[27][4] ), .A1(n14), .Z(n1075));
Q_MX02 U1053 ( .S(n45), .A0(\rst_dat[27][5] ), .A1(n15), .Z(n1076));
Q_MX02 U1054 ( .S(n45), .A0(\rst_dat[27][6] ), .A1(n16), .Z(n1077));
Q_MX02 U1055 ( .S(n45), .A0(\rst_dat[27][7] ), .A1(n17), .Z(n1078));
Q_MX02 U1056 ( .S(n45), .A0(\rst_dat[27][8] ), .A1(n18), .Z(n1079));
Q_MX02 U1057 ( .S(n45), .A0(\rst_dat[27][9] ), .A1(n19), .Z(n1080));
Q_MX02 U1058 ( .S(n45), .A0(\rst_dat[27][10] ), .A1(n20), .Z(n1081));
Q_MX02 U1059 ( .S(n45), .A0(\rst_dat[27][11] ), .A1(n21), .Z(n1082));
Q_MX02 U1060 ( .S(n45), .A0(\rst_dat[27][12] ), .A1(n22), .Z(n1083));
Q_MX02 U1061 ( .S(n45), .A0(\rst_dat[27][13] ), .A1(n23), .Z(n1084));
Q_MX02 U1062 ( .S(n45), .A0(\rst_dat[27][14] ), .A1(n24), .Z(n1085));
Q_MX02 U1063 ( .S(n45), .A0(\rst_dat[27][15] ), .A1(n25), .Z(n1086));
Q_MX02 U1064 ( .S(n45), .A0(\rst_dat[27][16] ), .A1(n26), .Z(n1087));
Q_MX02 U1065 ( .S(n45), .A0(\rst_dat[27][17] ), .A1(n27), .Z(n1088));
Q_MX02 U1066 ( .S(n45), .A0(\rst_dat[27][18] ), .A1(n28), .Z(n1089));
Q_MX02 U1067 ( .S(n45), .A0(\rst_dat[27][19] ), .A1(n29), .Z(n1090));
Q_MX02 U1068 ( .S(n45), .A0(\rst_dat[27][20] ), .A1(n30), .Z(n1091));
Q_MX02 U1069 ( .S(n45), .A0(\rst_dat[27][21] ), .A1(n31), .Z(n1092));
Q_MX02 U1070 ( .S(n45), .A0(\rst_dat[27][22] ), .A1(n32), .Z(n1093));
Q_MX02 U1071 ( .S(n45), .A0(\rst_dat[27][23] ), .A1(n33), .Z(n1094));
Q_MX02 U1072 ( .S(n45), .A0(\rst_dat[27][24] ), .A1(n34), .Z(n1095));
Q_MX02 U1073 ( .S(n45), .A0(\rst_dat[27][25] ), .A1(n35), .Z(n1096));
Q_MX02 U1074 ( .S(n45), .A0(\rst_dat[27][26] ), .A1(n36), .Z(n1097));
Q_MX02 U1075 ( .S(n45), .A0(\rst_dat[27][27] ), .A1(n37), .Z(n1098));
Q_MX02 U1076 ( .S(n45), .A0(\rst_dat[27][28] ), .A1(n38), .Z(n1099));
Q_MX02 U1077 ( .S(n45), .A0(\rst_dat[27][29] ), .A1(n39), .Z(n1100));
Q_MX02 U1078 ( .S(n45), .A0(\rst_dat[27][30] ), .A1(n40), .Z(n1101));
Q_MX02 U1079 ( .S(n45), .A0(\rst_dat[27][31] ), .A1(n41), .Z(n1102));
Q_MX02 U1080 ( .S(n45), .A0(\rst_dat[28][0] ), .A1(n10), .Z(n1104));
Q_MX02 U1081 ( .S(n45), .A0(\rst_dat[28][1] ), .A1(n11), .Z(n1105));
Q_MX02 U1082 ( .S(n45), .A0(\rst_dat[28][2] ), .A1(n12), .Z(n1106));
Q_MX02 U1083 ( .S(n45), .A0(\rst_dat[28][3] ), .A1(n13), .Z(n1107));
Q_MX02 U1084 ( .S(n45), .A0(\rst_dat[28][4] ), .A1(n14), .Z(n1108));
Q_MX02 U1085 ( .S(n45), .A0(\rst_dat[28][5] ), .A1(n15), .Z(n1109));
Q_MX02 U1086 ( .S(n45), .A0(\rst_dat[28][6] ), .A1(n16), .Z(n1110));
Q_MX02 U1087 ( .S(n45), .A0(\rst_dat[28][7] ), .A1(n17), .Z(n1111));
Q_MX02 U1088 ( .S(n45), .A0(\rst_dat[28][8] ), .A1(n18), .Z(n1112));
Q_MX02 U1089 ( .S(n45), .A0(\rst_dat[28][9] ), .A1(n19), .Z(n1113));
Q_MX02 U1090 ( .S(n45), .A0(\rst_dat[28][10] ), .A1(n20), .Z(n1114));
Q_MX02 U1091 ( .S(n45), .A0(\rst_dat[28][11] ), .A1(n21), .Z(n1115));
Q_MX02 U1092 ( .S(n45), .A0(\rst_dat[28][12] ), .A1(n22), .Z(n1116));
Q_MX02 U1093 ( .S(n45), .A0(\rst_dat[28][13] ), .A1(n23), .Z(n1117));
Q_MX02 U1094 ( .S(n45), .A0(\rst_dat[28][14] ), .A1(n24), .Z(n1118));
Q_MX02 U1095 ( .S(n45), .A0(\rst_dat[28][15] ), .A1(n25), .Z(n1119));
Q_MX02 U1096 ( .S(n45), .A0(\rst_dat[28][16] ), .A1(n26), .Z(n1120));
Q_MX02 U1097 ( .S(n45), .A0(\rst_dat[28][17] ), .A1(n27), .Z(n1121));
Q_MX02 U1098 ( .S(n45), .A0(\rst_dat[28][18] ), .A1(n28), .Z(n1122));
Q_MX02 U1099 ( .S(n45), .A0(\rst_dat[28][19] ), .A1(n29), .Z(n1123));
Q_MX02 U1100 ( .S(n45), .A0(\rst_dat[28][20] ), .A1(n30), .Z(n1124));
Q_MX02 U1101 ( .S(n45), .A0(\rst_dat[28][21] ), .A1(n31), .Z(n1125));
Q_MX02 U1102 ( .S(n45), .A0(\rst_dat[28][22] ), .A1(n32), .Z(n1126));
Q_MX02 U1103 ( .S(n45), .A0(\rst_dat[28][23] ), .A1(n33), .Z(n1127));
Q_MX02 U1104 ( .S(n45), .A0(\rst_dat[28][24] ), .A1(n34), .Z(n1128));
Q_MX02 U1105 ( .S(n45), .A0(\rst_dat[28][25] ), .A1(n35), .Z(n1129));
Q_MX02 U1106 ( .S(n45), .A0(\rst_dat[28][26] ), .A1(n36), .Z(n1130));
Q_MX02 U1107 ( .S(n45), .A0(\rst_dat[28][27] ), .A1(n37), .Z(n1131));
Q_MX02 U1108 ( .S(n45), .A0(\rst_dat[28][28] ), .A1(n38), .Z(n1132));
Q_MX02 U1109 ( .S(n45), .A0(\rst_dat[28][29] ), .A1(n39), .Z(n1133));
Q_MX02 U1110 ( .S(n45), .A0(\rst_dat[28][30] ), .A1(n40), .Z(n1134));
Q_MX02 U1111 ( .S(n45), .A0(\rst_dat[28][31] ), .A1(n41), .Z(n1135));
Q_MX02 U1112 ( .S(n45), .A0(\rst_dat[29][0] ), .A1(n10), .Z(n1137));
Q_MX02 U1113 ( .S(n45), .A0(\rst_dat[29][1] ), .A1(n11), .Z(n1138));
Q_MX02 U1114 ( .S(n45), .A0(\rst_dat[29][2] ), .A1(n12), .Z(n1139));
Q_MX02 U1115 ( .S(n45), .A0(\rst_dat[29][3] ), .A1(n13), .Z(n1140));
Q_MX02 U1116 ( .S(n45), .A0(\rst_dat[29][4] ), .A1(n14), .Z(n1141));
Q_MX02 U1117 ( .S(n45), .A0(\rst_dat[29][5] ), .A1(n15), .Z(n1142));
Q_MX02 U1118 ( .S(n45), .A0(\rst_dat[29][6] ), .A1(n16), .Z(n1143));
Q_MX02 U1119 ( .S(n45), .A0(\rst_dat[29][7] ), .A1(n17), .Z(n1144));
Q_MX02 U1120 ( .S(n45), .A0(\rst_dat[29][8] ), .A1(n18), .Z(n1145));
Q_MX02 U1121 ( .S(n45), .A0(\rst_dat[29][9] ), .A1(n19), .Z(n1146));
Q_MX02 U1122 ( .S(n45), .A0(\rst_dat[29][10] ), .A1(n20), .Z(n1147));
Q_MX02 U1123 ( .S(n45), .A0(\rst_dat[29][11] ), .A1(n21), .Z(n1148));
Q_MX02 U1124 ( .S(n45), .A0(\rst_dat[29][12] ), .A1(n22), .Z(n1149));
Q_MX02 U1125 ( .S(n45), .A0(\rst_dat[29][13] ), .A1(n23), .Z(n1150));
Q_MX02 U1126 ( .S(n45), .A0(\rst_dat[29][14] ), .A1(n24), .Z(n1151));
Q_MX02 U1127 ( .S(n45), .A0(\rst_dat[29][15] ), .A1(n25), .Z(n1152));
Q_MX02 U1128 ( .S(n45), .A0(\rst_dat[29][16] ), .A1(n26), .Z(n1153));
Q_MX02 U1129 ( .S(n45), .A0(\rst_dat[29][17] ), .A1(n27), .Z(n1154));
Q_MX02 U1130 ( .S(n45), .A0(\rst_dat[29][18] ), .A1(n28), .Z(n1155));
Q_MX02 U1131 ( .S(n45), .A0(\rst_dat[29][19] ), .A1(n29), .Z(n1156));
Q_MX02 U1132 ( .S(n45), .A0(\rst_dat[29][20] ), .A1(n30), .Z(n1157));
Q_MX02 U1133 ( .S(n45), .A0(\rst_dat[29][21] ), .A1(n31), .Z(n1158));
Q_MX02 U1134 ( .S(n45), .A0(\rst_dat[29][22] ), .A1(n32), .Z(n1159));
Q_MX02 U1135 ( .S(n45), .A0(\rst_dat[29][23] ), .A1(n33), .Z(n1160));
Q_MX02 U1136 ( .S(n45), .A0(\rst_dat[29][24] ), .A1(n34), .Z(n1161));
Q_MX02 U1137 ( .S(n45), .A0(\rst_dat[29][25] ), .A1(n35), .Z(n1162));
Q_MX02 U1138 ( .S(n45), .A0(\rst_dat[29][26] ), .A1(n36), .Z(n1163));
Q_MX02 U1139 ( .S(n45), .A0(\rst_dat[29][27] ), .A1(n37), .Z(n1164));
Q_MX02 U1140 ( .S(n45), .A0(\rst_dat[29][28] ), .A1(n38), .Z(n1165));
Q_MX02 U1141 ( .S(n45), .A0(\rst_dat[29][29] ), .A1(n39), .Z(n1166));
Q_MX02 U1142 ( .S(n45), .A0(\rst_dat[29][30] ), .A1(n40), .Z(n1167));
Q_MX02 U1143 ( .S(n45), .A0(\rst_dat[29][31] ), .A1(n41), .Z(n1168));
Q_MX02 U1144 ( .S(n45), .A0(\rst_dat[30][0] ), .A1(n10), .Z(n1170));
Q_MX02 U1145 ( .S(n45), .A0(\rst_dat[30][1] ), .A1(n11), .Z(n1171));
Q_MX02 U1146 ( .S(n45), .A0(\rst_dat[30][2] ), .A1(n12), .Z(n1172));
Q_MX02 U1147 ( .S(n45), .A0(\rst_dat[30][3] ), .A1(n13), .Z(n1173));
Q_MX02 U1148 ( .S(n45), .A0(\rst_dat[30][4] ), .A1(n14), .Z(n1174));
Q_MX02 U1149 ( .S(n45), .A0(\rst_dat[30][5] ), .A1(n15), .Z(n1175));
Q_MX02 U1150 ( .S(n45), .A0(\rst_dat[30][6] ), .A1(n16), .Z(n1176));
Q_MX02 U1151 ( .S(n45), .A0(\rst_dat[30][7] ), .A1(n17), .Z(n1177));
Q_MX02 U1152 ( .S(n45), .A0(\rst_dat[30][8] ), .A1(n18), .Z(n1178));
Q_MX02 U1153 ( .S(n45), .A0(\rst_dat[30][9] ), .A1(n19), .Z(n1179));
Q_MX02 U1154 ( .S(n45), .A0(\rst_dat[30][10] ), .A1(n20), .Z(n1180));
Q_MX02 U1155 ( .S(n45), .A0(\rst_dat[30][11] ), .A1(n21), .Z(n1181));
Q_MX02 U1156 ( .S(n45), .A0(\rst_dat[30][12] ), .A1(n22), .Z(n1182));
Q_MX02 U1157 ( .S(n45), .A0(\rst_dat[30][13] ), .A1(n23), .Z(n1183));
Q_MX02 U1158 ( .S(n45), .A0(\rst_dat[30][14] ), .A1(n24), .Z(n1184));
Q_MX02 U1159 ( .S(n45), .A0(\rst_dat[30][15] ), .A1(n25), .Z(n1185));
Q_MX02 U1160 ( .S(n45), .A0(\rst_dat[30][16] ), .A1(n26), .Z(n1186));
Q_MX02 U1161 ( .S(n45), .A0(\rst_dat[30][17] ), .A1(n27), .Z(n1187));
Q_MX02 U1162 ( .S(n45), .A0(\rst_dat[30][18] ), .A1(n28), .Z(n1188));
Q_MX02 U1163 ( .S(n45), .A0(\rst_dat[30][19] ), .A1(n29), .Z(n1189));
Q_MX02 U1164 ( .S(n45), .A0(\rst_dat[30][20] ), .A1(n30), .Z(n1190));
Q_MX02 U1165 ( .S(n45), .A0(\rst_dat[30][21] ), .A1(n31), .Z(n1191));
Q_MX02 U1166 ( .S(n45), .A0(\rst_dat[30][22] ), .A1(n32), .Z(n1192));
Q_MX02 U1167 ( .S(n45), .A0(\rst_dat[30][23] ), .A1(n33), .Z(n1193));
Q_MX02 U1168 ( .S(n45), .A0(\rst_dat[30][24] ), .A1(n34), .Z(n1194));
Q_MX02 U1169 ( .S(n45), .A0(\rst_dat[30][25] ), .A1(n35), .Z(n1195));
Q_MX02 U1170 ( .S(n45), .A0(\rst_dat[30][26] ), .A1(n36), .Z(n1196));
Q_MX02 U1171 ( .S(n45), .A0(\rst_dat[30][27] ), .A1(n37), .Z(n1197));
Q_MX02 U1172 ( .S(n45), .A0(\rst_dat[30][28] ), .A1(n38), .Z(n1198));
Q_MX02 U1173 ( .S(n45), .A0(\rst_dat[30][29] ), .A1(n39), .Z(n1199));
Q_MX02 U1174 ( .S(n45), .A0(\rst_dat[30][30] ), .A1(n40), .Z(n1200));
Q_MX02 U1175 ( .S(n45), .A0(\rst_dat[30][31] ), .A1(n41), .Z(n1201));
Q_MX02 U1176 ( .S(n45), .A0(\rst_dat[31][0] ), .A1(n10), .Z(n1203));
Q_MX02 U1177 ( .S(n45), .A0(\rst_dat[31][1] ), .A1(n11), .Z(n1204));
Q_MX02 U1178 ( .S(n45), .A0(\rst_dat[31][2] ), .A1(n12), .Z(n1205));
Q_MX02 U1179 ( .S(n45), .A0(\rst_dat[31][3] ), .A1(n13), .Z(n1206));
Q_MX02 U1180 ( .S(n45), .A0(\rst_dat[31][4] ), .A1(n14), .Z(n1207));
Q_MX02 U1181 ( .S(n45), .A0(\rst_dat[31][5] ), .A1(n15), .Z(n1208));
Q_MX02 U1182 ( .S(n45), .A0(\rst_dat[31][6] ), .A1(n16), .Z(n1209));
Q_MX02 U1183 ( .S(n45), .A0(\rst_dat[31][7] ), .A1(n17), .Z(n1210));
Q_MX02 U1184 ( .S(n45), .A0(\rst_dat[31][8] ), .A1(n18), .Z(n1211));
Q_MX02 U1185 ( .S(n45), .A0(\rst_dat[31][9] ), .A1(n19), .Z(n1212));
Q_MX02 U1186 ( .S(n45), .A0(\rst_dat[31][10] ), .A1(n20), .Z(n1213));
Q_MX02 U1187 ( .S(n45), .A0(\rst_dat[31][11] ), .A1(n21), .Z(n1214));
Q_MX02 U1188 ( .S(n45), .A0(\rst_dat[31][12] ), .A1(n22), .Z(n1215));
Q_MX02 U1189 ( .S(n45), .A0(\rst_dat[31][13] ), .A1(n23), .Z(n1216));
Q_MX02 U1190 ( .S(n45), .A0(\rst_dat[31][14] ), .A1(n24), .Z(n1217));
Q_MX02 U1191 ( .S(n45), .A0(\rst_dat[31][15] ), .A1(n25), .Z(n1218));
Q_MX02 U1192 ( .S(n45), .A0(\rst_dat[31][16] ), .A1(n26), .Z(n1219));
Q_MX02 U1193 ( .S(n45), .A0(\rst_dat[31][17] ), .A1(n27), .Z(n1220));
Q_MX02 U1194 ( .S(n45), .A0(\rst_dat[31][18] ), .A1(n28), .Z(n1221));
Q_MX02 U1195 ( .S(n45), .A0(\rst_dat[31][19] ), .A1(n29), .Z(n1222));
Q_MX02 U1196 ( .S(n45), .A0(\rst_dat[31][20] ), .A1(n30), .Z(n1223));
Q_MX02 U1197 ( .S(n45), .A0(\rst_dat[31][21] ), .A1(n31), .Z(n1224));
Q_MX02 U1198 ( .S(n45), .A0(\rst_dat[31][22] ), .A1(n32), .Z(n1225));
Q_MX02 U1199 ( .S(n45), .A0(\rst_dat[31][23] ), .A1(n33), .Z(n1226));
Q_MX02 U1200 ( .S(n45), .A0(\rst_dat[31][24] ), .A1(n34), .Z(n1227));
Q_MX02 U1201 ( .S(n45), .A0(\rst_dat[31][25] ), .A1(n35), .Z(n1228));
Q_MX02 U1202 ( .S(n45), .A0(\rst_dat[31][26] ), .A1(n36), .Z(n1229));
Q_MX02 U1203 ( .S(n45), .A0(\rst_dat[31][27] ), .A1(n37), .Z(n1230));
Q_MX02 U1204 ( .S(n45), .A0(\rst_dat[31][28] ), .A1(n38), .Z(n1231));
Q_MX02 U1205 ( .S(n45), .A0(\rst_dat[31][29] ), .A1(n39), .Z(n1232));
Q_MX02 U1206 ( .S(n45), .A0(\rst_dat[31][30] ), .A1(n40), .Z(n1233));
Q_MX02 U1207 ( .S(n45), .A0(\rst_dat[31][31] ), .A1(n41), .Z(n1234));
Q_MX08 U1208 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][0] ), .A1(\mem_a[25][0] ), .A2(\mem_a[26][0] ), .A3(\mem_a[27][0] ), .A4(\mem_a[28][0] ), .A5(\mem_a[29][0] ), .A6(\mem_a[30][0] ), .A7(\mem_a[31][0] ), .Z(n1235));
Q_MX08 U1209 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][0] ), .A1(\mem_a[17][0] ), .A2(\mem_a[18][0] ), .A3(\mem_a[19][0] ), .A4(\mem_a[20][0] ), .A5(\mem_a[21][0] ), .A6(\mem_a[22][0] ), .A7(\mem_a[23][0] ), .Z(n1236));
Q_MX08 U1210 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][0] ), .A1(\mem_a[9][0] ), .A2(\mem_a[10][0] ), .A3(\mem_a[11][0] ), .A4(\mem_a[12][0] ), .A5(\mem_a[13][0] ), .A6(\mem_a[14][0] ), .A7(\mem_a[15][0] ), .Z(n1237));
Q_MX08 U1211 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][0] ), .A1(\mem_a[1][0] ), .A2(\mem_a[2][0] ), .A3(\mem_a[3][0] ), .A4(\mem_a[4][0] ), .A5(\mem_a[5][0] ), .A6(\mem_a[6][0] ), .A7(\mem_a[7][0] ), .Z(n1238));
Q_MX04 U1212 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1238), .A1(n1237), .A2(n1236), .A3(n1235), .Z(n110));
Q_MX08 U1213 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][1] ), .A1(\mem_a[25][1] ), .A2(\mem_a[26][1] ), .A3(\mem_a[27][1] ), .A4(\mem_a[28][1] ), .A5(\mem_a[29][1] ), .A6(\mem_a[30][1] ), .A7(\mem_a[31][1] ), .Z(n1239));
Q_MX08 U1214 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][1] ), .A1(\mem_a[17][1] ), .A2(\mem_a[18][1] ), .A3(\mem_a[19][1] ), .A4(\mem_a[20][1] ), .A5(\mem_a[21][1] ), .A6(\mem_a[22][1] ), .A7(\mem_a[23][1] ), .Z(n1240));
Q_MX08 U1215 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][1] ), .A1(\mem_a[9][1] ), .A2(\mem_a[10][1] ), .A3(\mem_a[11][1] ), .A4(\mem_a[12][1] ), .A5(\mem_a[13][1] ), .A6(\mem_a[14][1] ), .A7(\mem_a[15][1] ), .Z(n1241));
Q_MX08 U1216 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][1] ), .A1(\mem_a[1][1] ), .A2(\mem_a[2][1] ), .A3(\mem_a[3][1] ), .A4(\mem_a[4][1] ), .A5(\mem_a[5][1] ), .A6(\mem_a[6][1] ), .A7(\mem_a[7][1] ), .Z(n1242));
Q_MX04 U1217 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1242), .A1(n1241), .A2(n1240), .A3(n1239), .Z(n109));
Q_MX08 U1218 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][2] ), .A1(\mem_a[25][2] ), .A2(\mem_a[26][2] ), .A3(\mem_a[27][2] ), .A4(\mem_a[28][2] ), .A5(\mem_a[29][2] ), .A6(\mem_a[30][2] ), .A7(\mem_a[31][2] ), .Z(n1243));
Q_MX08 U1219 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][2] ), .A1(\mem_a[17][2] ), .A2(\mem_a[18][2] ), .A3(\mem_a[19][2] ), .A4(\mem_a[20][2] ), .A5(\mem_a[21][2] ), .A6(\mem_a[22][2] ), .A7(\mem_a[23][2] ), .Z(n1244));
Q_MX08 U1220 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][2] ), .A1(\mem_a[9][2] ), .A2(\mem_a[10][2] ), .A3(\mem_a[11][2] ), .A4(\mem_a[12][2] ), .A5(\mem_a[13][2] ), .A6(\mem_a[14][2] ), .A7(\mem_a[15][2] ), .Z(n1245));
Q_MX08 U1221 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][2] ), .A1(\mem_a[1][2] ), .A2(\mem_a[2][2] ), .A3(\mem_a[3][2] ), .A4(\mem_a[4][2] ), .A5(\mem_a[5][2] ), .A6(\mem_a[6][2] ), .A7(\mem_a[7][2] ), .Z(n1246));
Q_MX04 U1222 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1246), .A1(n1245), .A2(n1244), .A3(n1243), .Z(n108));
Q_MX08 U1223 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][3] ), .A1(\mem_a[25][3] ), .A2(\mem_a[26][3] ), .A3(\mem_a[27][3] ), .A4(\mem_a[28][3] ), .A5(\mem_a[29][3] ), .A6(\mem_a[30][3] ), .A7(\mem_a[31][3] ), .Z(n1247));
Q_MX08 U1224 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][3] ), .A1(\mem_a[17][3] ), .A2(\mem_a[18][3] ), .A3(\mem_a[19][3] ), .A4(\mem_a[20][3] ), .A5(\mem_a[21][3] ), .A6(\mem_a[22][3] ), .A7(\mem_a[23][3] ), .Z(n1248));
Q_MX08 U1225 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][3] ), .A1(\mem_a[9][3] ), .A2(\mem_a[10][3] ), .A3(\mem_a[11][3] ), .A4(\mem_a[12][3] ), .A5(\mem_a[13][3] ), .A6(\mem_a[14][3] ), .A7(\mem_a[15][3] ), .Z(n1249));
Q_MX08 U1226 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][3] ), .A1(\mem_a[1][3] ), .A2(\mem_a[2][3] ), .A3(\mem_a[3][3] ), .A4(\mem_a[4][3] ), .A5(\mem_a[5][3] ), .A6(\mem_a[6][3] ), .A7(\mem_a[7][3] ), .Z(n1250));
Q_MX04 U1227 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1250), .A1(n1249), .A2(n1248), .A3(n1247), .Z(n107));
Q_MX08 U1228 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][4] ), .A1(\mem_a[25][4] ), .A2(\mem_a[26][4] ), .A3(\mem_a[27][4] ), .A4(\mem_a[28][4] ), .A5(\mem_a[29][4] ), .A6(\mem_a[30][4] ), .A7(\mem_a[31][4] ), .Z(n1251));
Q_MX08 U1229 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][4] ), .A1(\mem_a[17][4] ), .A2(\mem_a[18][4] ), .A3(\mem_a[19][4] ), .A4(\mem_a[20][4] ), .A5(\mem_a[21][4] ), .A6(\mem_a[22][4] ), .A7(\mem_a[23][4] ), .Z(n1252));
Q_MX08 U1230 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][4] ), .A1(\mem_a[9][4] ), .A2(\mem_a[10][4] ), .A3(\mem_a[11][4] ), .A4(\mem_a[12][4] ), .A5(\mem_a[13][4] ), .A6(\mem_a[14][4] ), .A7(\mem_a[15][4] ), .Z(n1253));
Q_MX08 U1231 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][4] ), .A1(\mem_a[1][4] ), .A2(\mem_a[2][4] ), .A3(\mem_a[3][4] ), .A4(\mem_a[4][4] ), .A5(\mem_a[5][4] ), .A6(\mem_a[6][4] ), .A7(\mem_a[7][4] ), .Z(n1254));
Q_MX04 U1232 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1254), .A1(n1253), .A2(n1252), .A3(n1251), .Z(n106));
Q_MX08 U1233 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][5] ), .A1(\mem_a[25][5] ), .A2(\mem_a[26][5] ), .A3(\mem_a[27][5] ), .A4(\mem_a[28][5] ), .A5(\mem_a[29][5] ), .A6(\mem_a[30][5] ), .A7(\mem_a[31][5] ), .Z(n1255));
Q_MX08 U1234 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][5] ), .A1(\mem_a[17][5] ), .A2(\mem_a[18][5] ), .A3(\mem_a[19][5] ), .A4(\mem_a[20][5] ), .A5(\mem_a[21][5] ), .A6(\mem_a[22][5] ), .A7(\mem_a[23][5] ), .Z(n1256));
Q_MX08 U1235 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][5] ), .A1(\mem_a[9][5] ), .A2(\mem_a[10][5] ), .A3(\mem_a[11][5] ), .A4(\mem_a[12][5] ), .A5(\mem_a[13][5] ), .A6(\mem_a[14][5] ), .A7(\mem_a[15][5] ), .Z(n1257));
Q_MX08 U1236 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][5] ), .A1(\mem_a[1][5] ), .A2(\mem_a[2][5] ), .A3(\mem_a[3][5] ), .A4(\mem_a[4][5] ), .A5(\mem_a[5][5] ), .A6(\mem_a[6][5] ), .A7(\mem_a[7][5] ), .Z(n1258));
Q_MX04 U1237 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1258), .A1(n1257), .A2(n1256), .A3(n1255), .Z(n105));
Q_MX08 U1238 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][6] ), .A1(\mem_a[25][6] ), .A2(\mem_a[26][6] ), .A3(\mem_a[27][6] ), .A4(\mem_a[28][6] ), .A5(\mem_a[29][6] ), .A6(\mem_a[30][6] ), .A7(\mem_a[31][6] ), .Z(n1259));
Q_MX08 U1239 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][6] ), .A1(\mem_a[17][6] ), .A2(\mem_a[18][6] ), .A3(\mem_a[19][6] ), .A4(\mem_a[20][6] ), .A5(\mem_a[21][6] ), .A6(\mem_a[22][6] ), .A7(\mem_a[23][6] ), .Z(n1260));
Q_MX08 U1240 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][6] ), .A1(\mem_a[9][6] ), .A2(\mem_a[10][6] ), .A3(\mem_a[11][6] ), .A4(\mem_a[12][6] ), .A5(\mem_a[13][6] ), .A6(\mem_a[14][6] ), .A7(\mem_a[15][6] ), .Z(n1261));
Q_MX08 U1241 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][6] ), .A1(\mem_a[1][6] ), .A2(\mem_a[2][6] ), .A3(\mem_a[3][6] ), .A4(\mem_a[4][6] ), .A5(\mem_a[5][6] ), .A6(\mem_a[6][6] ), .A7(\mem_a[7][6] ), .Z(n1262));
Q_MX04 U1242 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1262), .A1(n1261), .A2(n1260), .A3(n1259), .Z(n104));
Q_MX08 U1243 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][7] ), .A1(\mem_a[25][7] ), .A2(\mem_a[26][7] ), .A3(\mem_a[27][7] ), .A4(\mem_a[28][7] ), .A5(\mem_a[29][7] ), .A6(\mem_a[30][7] ), .A7(\mem_a[31][7] ), .Z(n1263));
Q_MX08 U1244 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][7] ), .A1(\mem_a[17][7] ), .A2(\mem_a[18][7] ), .A3(\mem_a[19][7] ), .A4(\mem_a[20][7] ), .A5(\mem_a[21][7] ), .A6(\mem_a[22][7] ), .A7(\mem_a[23][7] ), .Z(n1264));
Q_MX08 U1245 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][7] ), .A1(\mem_a[9][7] ), .A2(\mem_a[10][7] ), .A3(\mem_a[11][7] ), .A4(\mem_a[12][7] ), .A5(\mem_a[13][7] ), .A6(\mem_a[14][7] ), .A7(\mem_a[15][7] ), .Z(n1265));
Q_MX08 U1246 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][7] ), .A1(\mem_a[1][7] ), .A2(\mem_a[2][7] ), .A3(\mem_a[3][7] ), .A4(\mem_a[4][7] ), .A5(\mem_a[5][7] ), .A6(\mem_a[6][7] ), .A7(\mem_a[7][7] ), .Z(n1266));
Q_MX04 U1247 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1266), .A1(n1265), .A2(n1264), .A3(n1263), .Z(n103));
Q_MX08 U1248 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][8] ), .A1(\mem_a[25][8] ), .A2(\mem_a[26][8] ), .A3(\mem_a[27][8] ), .A4(\mem_a[28][8] ), .A5(\mem_a[29][8] ), .A6(\mem_a[30][8] ), .A7(\mem_a[31][8] ), .Z(n1267));
Q_MX08 U1249 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][8] ), .A1(\mem_a[17][8] ), .A2(\mem_a[18][8] ), .A3(\mem_a[19][8] ), .A4(\mem_a[20][8] ), .A5(\mem_a[21][8] ), .A6(\mem_a[22][8] ), .A7(\mem_a[23][8] ), .Z(n1268));
Q_MX08 U1250 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][8] ), .A1(\mem_a[9][8] ), .A2(\mem_a[10][8] ), .A3(\mem_a[11][8] ), .A4(\mem_a[12][8] ), .A5(\mem_a[13][8] ), .A6(\mem_a[14][8] ), .A7(\mem_a[15][8] ), .Z(n1269));
Q_MX08 U1251 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][8] ), .A1(\mem_a[1][8] ), .A2(\mem_a[2][8] ), .A3(\mem_a[3][8] ), .A4(\mem_a[4][8] ), .A5(\mem_a[5][8] ), .A6(\mem_a[6][8] ), .A7(\mem_a[7][8] ), .Z(n1270));
Q_MX04 U1252 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1270), .A1(n1269), .A2(n1268), .A3(n1267), .Z(n102));
Q_MX08 U1253 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][9] ), .A1(\mem_a[25][9] ), .A2(\mem_a[26][9] ), .A3(\mem_a[27][9] ), .A4(\mem_a[28][9] ), .A5(\mem_a[29][9] ), .A6(\mem_a[30][9] ), .A7(\mem_a[31][9] ), .Z(n1271));
Q_MX08 U1254 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][9] ), .A1(\mem_a[17][9] ), .A2(\mem_a[18][9] ), .A3(\mem_a[19][9] ), .A4(\mem_a[20][9] ), .A5(\mem_a[21][9] ), .A6(\mem_a[22][9] ), .A7(\mem_a[23][9] ), .Z(n1272));
Q_MX08 U1255 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][9] ), .A1(\mem_a[9][9] ), .A2(\mem_a[10][9] ), .A3(\mem_a[11][9] ), .A4(\mem_a[12][9] ), .A5(\mem_a[13][9] ), .A6(\mem_a[14][9] ), .A7(\mem_a[15][9] ), .Z(n1273));
Q_MX08 U1256 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][9] ), .A1(\mem_a[1][9] ), .A2(\mem_a[2][9] ), .A3(\mem_a[3][9] ), .A4(\mem_a[4][9] ), .A5(\mem_a[5][9] ), .A6(\mem_a[6][9] ), .A7(\mem_a[7][9] ), .Z(n1274));
Q_MX04 U1257 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1274), .A1(n1273), .A2(n1272), .A3(n1271), .Z(n101));
Q_MX08 U1258 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][10] ), .A1(\mem_a[25][10] ), .A2(\mem_a[26][10] ), .A3(\mem_a[27][10] ), .A4(\mem_a[28][10] ), .A5(\mem_a[29][10] ), .A6(\mem_a[30][10] ), .A7(\mem_a[31][10] ), .Z(n1275));
Q_MX08 U1259 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][10] ), .A1(\mem_a[17][10] ), .A2(\mem_a[18][10] ), .A3(\mem_a[19][10] ), .A4(\mem_a[20][10] ), .A5(\mem_a[21][10] ), .A6(\mem_a[22][10] ), .A7(\mem_a[23][10] ), .Z(n1276));
Q_MX08 U1260 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][10] ), .A1(\mem_a[9][10] ), .A2(\mem_a[10][10] ), .A3(\mem_a[11][10] ), .A4(\mem_a[12][10] ), .A5(\mem_a[13][10] ), .A6(\mem_a[14][10] ), .A7(\mem_a[15][10] ), .Z(n1277));
Q_MX08 U1261 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][10] ), .A1(\mem_a[1][10] ), .A2(\mem_a[2][10] ), .A3(\mem_a[3][10] ), .A4(\mem_a[4][10] ), .A5(\mem_a[5][10] ), .A6(\mem_a[6][10] ), .A7(\mem_a[7][10] ), .Z(n1278));
Q_MX04 U1262 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1278), .A1(n1277), .A2(n1276), .A3(n1275), .Z(n100));
Q_MX08 U1263 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][11] ), .A1(\mem_a[25][11] ), .A2(\mem_a[26][11] ), .A3(\mem_a[27][11] ), .A4(\mem_a[28][11] ), .A5(\mem_a[29][11] ), .A6(\mem_a[30][11] ), .A7(\mem_a[31][11] ), .Z(n1279));
Q_MX08 U1264 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][11] ), .A1(\mem_a[17][11] ), .A2(\mem_a[18][11] ), .A3(\mem_a[19][11] ), .A4(\mem_a[20][11] ), .A5(\mem_a[21][11] ), .A6(\mem_a[22][11] ), .A7(\mem_a[23][11] ), .Z(n1280));
Q_MX08 U1265 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][11] ), .A1(\mem_a[9][11] ), .A2(\mem_a[10][11] ), .A3(\mem_a[11][11] ), .A4(\mem_a[12][11] ), .A5(\mem_a[13][11] ), .A6(\mem_a[14][11] ), .A7(\mem_a[15][11] ), .Z(n1281));
Q_MX08 U1266 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][11] ), .A1(\mem_a[1][11] ), .A2(\mem_a[2][11] ), .A3(\mem_a[3][11] ), .A4(\mem_a[4][11] ), .A5(\mem_a[5][11] ), .A6(\mem_a[6][11] ), .A7(\mem_a[7][11] ), .Z(n1282));
Q_MX04 U1267 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1282), .A1(n1281), .A2(n1280), .A3(n1279), .Z(n99));
Q_MX08 U1268 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][12] ), .A1(\mem_a[25][12] ), .A2(\mem_a[26][12] ), .A3(\mem_a[27][12] ), .A4(\mem_a[28][12] ), .A5(\mem_a[29][12] ), .A6(\mem_a[30][12] ), .A7(\mem_a[31][12] ), .Z(n1283));
Q_MX08 U1269 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][12] ), .A1(\mem_a[17][12] ), .A2(\mem_a[18][12] ), .A3(\mem_a[19][12] ), .A4(\mem_a[20][12] ), .A5(\mem_a[21][12] ), .A6(\mem_a[22][12] ), .A7(\mem_a[23][12] ), .Z(n1284));
Q_MX08 U1270 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][12] ), .A1(\mem_a[9][12] ), .A2(\mem_a[10][12] ), .A3(\mem_a[11][12] ), .A4(\mem_a[12][12] ), .A5(\mem_a[13][12] ), .A6(\mem_a[14][12] ), .A7(\mem_a[15][12] ), .Z(n1285));
Q_MX08 U1271 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][12] ), .A1(\mem_a[1][12] ), .A2(\mem_a[2][12] ), .A3(\mem_a[3][12] ), .A4(\mem_a[4][12] ), .A5(\mem_a[5][12] ), .A6(\mem_a[6][12] ), .A7(\mem_a[7][12] ), .Z(n1286));
Q_MX04 U1272 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1286), .A1(n1285), .A2(n1284), .A3(n1283), .Z(n98));
Q_MX08 U1273 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][13] ), .A1(\mem_a[25][13] ), .A2(\mem_a[26][13] ), .A3(\mem_a[27][13] ), .A4(\mem_a[28][13] ), .A5(\mem_a[29][13] ), .A6(\mem_a[30][13] ), .A7(\mem_a[31][13] ), .Z(n1287));
Q_MX08 U1274 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][13] ), .A1(\mem_a[17][13] ), .A2(\mem_a[18][13] ), .A3(\mem_a[19][13] ), .A4(\mem_a[20][13] ), .A5(\mem_a[21][13] ), .A6(\mem_a[22][13] ), .A7(\mem_a[23][13] ), .Z(n1288));
Q_MX08 U1275 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][13] ), .A1(\mem_a[9][13] ), .A2(\mem_a[10][13] ), .A3(\mem_a[11][13] ), .A4(\mem_a[12][13] ), .A5(\mem_a[13][13] ), .A6(\mem_a[14][13] ), .A7(\mem_a[15][13] ), .Z(n1289));
Q_MX08 U1276 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][13] ), .A1(\mem_a[1][13] ), .A2(\mem_a[2][13] ), .A3(\mem_a[3][13] ), .A4(\mem_a[4][13] ), .A5(\mem_a[5][13] ), .A6(\mem_a[6][13] ), .A7(\mem_a[7][13] ), .Z(n1290));
Q_MX04 U1277 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1290), .A1(n1289), .A2(n1288), .A3(n1287), .Z(n97));
Q_MX08 U1278 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][14] ), .A1(\mem_a[25][14] ), .A2(\mem_a[26][14] ), .A3(\mem_a[27][14] ), .A4(\mem_a[28][14] ), .A5(\mem_a[29][14] ), .A6(\mem_a[30][14] ), .A7(\mem_a[31][14] ), .Z(n1291));
Q_MX08 U1279 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][14] ), .A1(\mem_a[17][14] ), .A2(\mem_a[18][14] ), .A3(\mem_a[19][14] ), .A4(\mem_a[20][14] ), .A5(\mem_a[21][14] ), .A6(\mem_a[22][14] ), .A7(\mem_a[23][14] ), .Z(n1292));
Q_MX08 U1280 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][14] ), .A1(\mem_a[9][14] ), .A2(\mem_a[10][14] ), .A3(\mem_a[11][14] ), .A4(\mem_a[12][14] ), .A5(\mem_a[13][14] ), .A6(\mem_a[14][14] ), .A7(\mem_a[15][14] ), .Z(n1293));
Q_MX08 U1281 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][14] ), .A1(\mem_a[1][14] ), .A2(\mem_a[2][14] ), .A3(\mem_a[3][14] ), .A4(\mem_a[4][14] ), .A5(\mem_a[5][14] ), .A6(\mem_a[6][14] ), .A7(\mem_a[7][14] ), .Z(n1294));
Q_MX04 U1282 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1294), .A1(n1293), .A2(n1292), .A3(n1291), .Z(n96));
Q_MX08 U1283 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][15] ), .A1(\mem_a[25][15] ), .A2(\mem_a[26][15] ), .A3(\mem_a[27][15] ), .A4(\mem_a[28][15] ), .A5(\mem_a[29][15] ), .A6(\mem_a[30][15] ), .A7(\mem_a[31][15] ), .Z(n1295));
Q_MX08 U1284 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][15] ), .A1(\mem_a[17][15] ), .A2(\mem_a[18][15] ), .A3(\mem_a[19][15] ), .A4(\mem_a[20][15] ), .A5(\mem_a[21][15] ), .A6(\mem_a[22][15] ), .A7(\mem_a[23][15] ), .Z(n1296));
Q_MX08 U1285 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][15] ), .A1(\mem_a[9][15] ), .A2(\mem_a[10][15] ), .A3(\mem_a[11][15] ), .A4(\mem_a[12][15] ), .A5(\mem_a[13][15] ), .A6(\mem_a[14][15] ), .A7(\mem_a[15][15] ), .Z(n1297));
Q_MX08 U1286 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][15] ), .A1(\mem_a[1][15] ), .A2(\mem_a[2][15] ), .A3(\mem_a[3][15] ), .A4(\mem_a[4][15] ), .A5(\mem_a[5][15] ), .A6(\mem_a[6][15] ), .A7(\mem_a[7][15] ), .Z(n1298));
Q_MX04 U1287 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1298), .A1(n1297), .A2(n1296), .A3(n1295), .Z(n95));
Q_MX08 U1288 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][16] ), .A1(\mem_a[25][16] ), .A2(\mem_a[26][16] ), .A3(\mem_a[27][16] ), .A4(\mem_a[28][16] ), .A5(\mem_a[29][16] ), .A6(\mem_a[30][16] ), .A7(\mem_a[31][16] ), .Z(n1299));
Q_MX08 U1289 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][16] ), .A1(\mem_a[17][16] ), .A2(\mem_a[18][16] ), .A3(\mem_a[19][16] ), .A4(\mem_a[20][16] ), .A5(\mem_a[21][16] ), .A6(\mem_a[22][16] ), .A7(\mem_a[23][16] ), .Z(n1300));
Q_MX08 U1290 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][16] ), .A1(\mem_a[9][16] ), .A2(\mem_a[10][16] ), .A3(\mem_a[11][16] ), .A4(\mem_a[12][16] ), .A5(\mem_a[13][16] ), .A6(\mem_a[14][16] ), .A7(\mem_a[15][16] ), .Z(n1301));
Q_MX08 U1291 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][16] ), .A1(\mem_a[1][16] ), .A2(\mem_a[2][16] ), .A3(\mem_a[3][16] ), .A4(\mem_a[4][16] ), .A5(\mem_a[5][16] ), .A6(\mem_a[6][16] ), .A7(\mem_a[7][16] ), .Z(n1302));
Q_MX04 U1292 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1302), .A1(n1301), .A2(n1300), .A3(n1299), .Z(n94));
Q_MX08 U1293 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][17] ), .A1(\mem_a[25][17] ), .A2(\mem_a[26][17] ), .A3(\mem_a[27][17] ), .A4(\mem_a[28][17] ), .A5(\mem_a[29][17] ), .A6(\mem_a[30][17] ), .A7(\mem_a[31][17] ), .Z(n1303));
Q_MX08 U1294 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][17] ), .A1(\mem_a[17][17] ), .A2(\mem_a[18][17] ), .A3(\mem_a[19][17] ), .A4(\mem_a[20][17] ), .A5(\mem_a[21][17] ), .A6(\mem_a[22][17] ), .A7(\mem_a[23][17] ), .Z(n1304));
Q_MX08 U1295 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][17] ), .A1(\mem_a[9][17] ), .A2(\mem_a[10][17] ), .A3(\mem_a[11][17] ), .A4(\mem_a[12][17] ), .A5(\mem_a[13][17] ), .A6(\mem_a[14][17] ), .A7(\mem_a[15][17] ), .Z(n1305));
Q_MX08 U1296 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][17] ), .A1(\mem_a[1][17] ), .A2(\mem_a[2][17] ), .A3(\mem_a[3][17] ), .A4(\mem_a[4][17] ), .A5(\mem_a[5][17] ), .A6(\mem_a[6][17] ), .A7(\mem_a[7][17] ), .Z(n1306));
Q_MX04 U1297 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1306), .A1(n1305), .A2(n1304), .A3(n1303), .Z(n93));
Q_MX08 U1298 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][18] ), .A1(\mem_a[25][18] ), .A2(\mem_a[26][18] ), .A3(\mem_a[27][18] ), .A4(\mem_a[28][18] ), .A5(\mem_a[29][18] ), .A6(\mem_a[30][18] ), .A7(\mem_a[31][18] ), .Z(n1307));
Q_MX08 U1299 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][18] ), .A1(\mem_a[17][18] ), .A2(\mem_a[18][18] ), .A3(\mem_a[19][18] ), .A4(\mem_a[20][18] ), .A5(\mem_a[21][18] ), .A6(\mem_a[22][18] ), .A7(\mem_a[23][18] ), .Z(n1308));
Q_MX08 U1300 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][18] ), .A1(\mem_a[9][18] ), .A2(\mem_a[10][18] ), .A3(\mem_a[11][18] ), .A4(\mem_a[12][18] ), .A5(\mem_a[13][18] ), .A6(\mem_a[14][18] ), .A7(\mem_a[15][18] ), .Z(n1309));
Q_MX08 U1301 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][18] ), .A1(\mem_a[1][18] ), .A2(\mem_a[2][18] ), .A3(\mem_a[3][18] ), .A4(\mem_a[4][18] ), .A5(\mem_a[5][18] ), .A6(\mem_a[6][18] ), .A7(\mem_a[7][18] ), .Z(n1310));
Q_MX04 U1302 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1310), .A1(n1309), .A2(n1308), .A3(n1307), .Z(n92));
Q_MX08 U1303 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][19] ), .A1(\mem_a[25][19] ), .A2(\mem_a[26][19] ), .A3(\mem_a[27][19] ), .A4(\mem_a[28][19] ), .A5(\mem_a[29][19] ), .A6(\mem_a[30][19] ), .A7(\mem_a[31][19] ), .Z(n1311));
Q_MX08 U1304 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][19] ), .A1(\mem_a[17][19] ), .A2(\mem_a[18][19] ), .A3(\mem_a[19][19] ), .A4(\mem_a[20][19] ), .A5(\mem_a[21][19] ), .A6(\mem_a[22][19] ), .A7(\mem_a[23][19] ), .Z(n1312));
Q_MX08 U1305 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][19] ), .A1(\mem_a[9][19] ), .A2(\mem_a[10][19] ), .A3(\mem_a[11][19] ), .A4(\mem_a[12][19] ), .A5(\mem_a[13][19] ), .A6(\mem_a[14][19] ), .A7(\mem_a[15][19] ), .Z(n1313));
Q_MX08 U1306 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][19] ), .A1(\mem_a[1][19] ), .A2(\mem_a[2][19] ), .A3(\mem_a[3][19] ), .A4(\mem_a[4][19] ), .A5(\mem_a[5][19] ), .A6(\mem_a[6][19] ), .A7(\mem_a[7][19] ), .Z(n1314));
Q_MX04 U1307 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1314), .A1(n1313), .A2(n1312), .A3(n1311), .Z(n91));
Q_MX08 U1308 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][20] ), .A1(\mem_a[25][20] ), .A2(\mem_a[26][20] ), .A3(\mem_a[27][20] ), .A4(\mem_a[28][20] ), .A5(\mem_a[29][20] ), .A6(\mem_a[30][20] ), .A7(\mem_a[31][20] ), .Z(n1315));
Q_MX08 U1309 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][20] ), .A1(\mem_a[17][20] ), .A2(\mem_a[18][20] ), .A3(\mem_a[19][20] ), .A4(\mem_a[20][20] ), .A5(\mem_a[21][20] ), .A6(\mem_a[22][20] ), .A7(\mem_a[23][20] ), .Z(n1316));
Q_MX08 U1310 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][20] ), .A1(\mem_a[9][20] ), .A2(\mem_a[10][20] ), .A3(\mem_a[11][20] ), .A4(\mem_a[12][20] ), .A5(\mem_a[13][20] ), .A6(\mem_a[14][20] ), .A7(\mem_a[15][20] ), .Z(n1317));
Q_MX08 U1311 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][20] ), .A1(\mem_a[1][20] ), .A2(\mem_a[2][20] ), .A3(\mem_a[3][20] ), .A4(\mem_a[4][20] ), .A5(\mem_a[5][20] ), .A6(\mem_a[6][20] ), .A7(\mem_a[7][20] ), .Z(n1318));
Q_MX04 U1312 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1318), .A1(n1317), .A2(n1316), .A3(n1315), .Z(n90));
Q_MX08 U1313 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][21] ), .A1(\mem_a[25][21] ), .A2(\mem_a[26][21] ), .A3(\mem_a[27][21] ), .A4(\mem_a[28][21] ), .A5(\mem_a[29][21] ), .A6(\mem_a[30][21] ), .A7(\mem_a[31][21] ), .Z(n1319));
Q_MX08 U1314 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][21] ), .A1(\mem_a[17][21] ), .A2(\mem_a[18][21] ), .A3(\mem_a[19][21] ), .A4(\mem_a[20][21] ), .A5(\mem_a[21][21] ), .A6(\mem_a[22][21] ), .A7(\mem_a[23][21] ), .Z(n1320));
Q_MX08 U1315 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][21] ), .A1(\mem_a[9][21] ), .A2(\mem_a[10][21] ), .A3(\mem_a[11][21] ), .A4(\mem_a[12][21] ), .A5(\mem_a[13][21] ), .A6(\mem_a[14][21] ), .A7(\mem_a[15][21] ), .Z(n1321));
Q_MX08 U1316 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][21] ), .A1(\mem_a[1][21] ), .A2(\mem_a[2][21] ), .A3(\mem_a[3][21] ), .A4(\mem_a[4][21] ), .A5(\mem_a[5][21] ), .A6(\mem_a[6][21] ), .A7(\mem_a[7][21] ), .Z(n1322));
Q_MX04 U1317 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1322), .A1(n1321), .A2(n1320), .A3(n1319), .Z(n89));
Q_MX08 U1318 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][22] ), .A1(\mem_a[25][22] ), .A2(\mem_a[26][22] ), .A3(\mem_a[27][22] ), .A4(\mem_a[28][22] ), .A5(\mem_a[29][22] ), .A6(\mem_a[30][22] ), .A7(\mem_a[31][22] ), .Z(n1323));
Q_MX08 U1319 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][22] ), .A1(\mem_a[17][22] ), .A2(\mem_a[18][22] ), .A3(\mem_a[19][22] ), .A4(\mem_a[20][22] ), .A5(\mem_a[21][22] ), .A6(\mem_a[22][22] ), .A7(\mem_a[23][22] ), .Z(n1324));
Q_MX08 U1320 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][22] ), .A1(\mem_a[9][22] ), .A2(\mem_a[10][22] ), .A3(\mem_a[11][22] ), .A4(\mem_a[12][22] ), .A5(\mem_a[13][22] ), .A6(\mem_a[14][22] ), .A7(\mem_a[15][22] ), .Z(n1325));
Q_MX08 U1321 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][22] ), .A1(\mem_a[1][22] ), .A2(\mem_a[2][22] ), .A3(\mem_a[3][22] ), .A4(\mem_a[4][22] ), .A5(\mem_a[5][22] ), .A6(\mem_a[6][22] ), .A7(\mem_a[7][22] ), .Z(n1326));
Q_MX04 U1322 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1326), .A1(n1325), .A2(n1324), .A3(n1323), .Z(n88));
Q_MX08 U1323 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][23] ), .A1(\mem_a[25][23] ), .A2(\mem_a[26][23] ), .A3(\mem_a[27][23] ), .A4(\mem_a[28][23] ), .A5(\mem_a[29][23] ), .A6(\mem_a[30][23] ), .A7(\mem_a[31][23] ), .Z(n1327));
Q_MX08 U1324 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][23] ), .A1(\mem_a[17][23] ), .A2(\mem_a[18][23] ), .A3(\mem_a[19][23] ), .A4(\mem_a[20][23] ), .A5(\mem_a[21][23] ), .A6(\mem_a[22][23] ), .A7(\mem_a[23][23] ), .Z(n1328));
Q_MX08 U1325 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][23] ), .A1(\mem_a[9][23] ), .A2(\mem_a[10][23] ), .A3(\mem_a[11][23] ), .A4(\mem_a[12][23] ), .A5(\mem_a[13][23] ), .A6(\mem_a[14][23] ), .A7(\mem_a[15][23] ), .Z(n1329));
Q_MX08 U1326 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][23] ), .A1(\mem_a[1][23] ), .A2(\mem_a[2][23] ), .A3(\mem_a[3][23] ), .A4(\mem_a[4][23] ), .A5(\mem_a[5][23] ), .A6(\mem_a[6][23] ), .A7(\mem_a[7][23] ), .Z(n1330));
Q_MX04 U1327 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1330), .A1(n1329), .A2(n1328), .A3(n1327), .Z(n87));
Q_MX08 U1328 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][24] ), .A1(\mem_a[25][24] ), .A2(\mem_a[26][24] ), .A3(\mem_a[27][24] ), .A4(\mem_a[28][24] ), .A5(\mem_a[29][24] ), .A6(\mem_a[30][24] ), .A7(\mem_a[31][24] ), .Z(n1331));
Q_MX08 U1329 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][24] ), .A1(\mem_a[17][24] ), .A2(\mem_a[18][24] ), .A3(\mem_a[19][24] ), .A4(\mem_a[20][24] ), .A5(\mem_a[21][24] ), .A6(\mem_a[22][24] ), .A7(\mem_a[23][24] ), .Z(n1332));
Q_MX08 U1330 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][24] ), .A1(\mem_a[9][24] ), .A2(\mem_a[10][24] ), .A3(\mem_a[11][24] ), .A4(\mem_a[12][24] ), .A5(\mem_a[13][24] ), .A6(\mem_a[14][24] ), .A7(\mem_a[15][24] ), .Z(n1333));
Q_MX08 U1331 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][24] ), .A1(\mem_a[1][24] ), .A2(\mem_a[2][24] ), .A3(\mem_a[3][24] ), .A4(\mem_a[4][24] ), .A5(\mem_a[5][24] ), .A6(\mem_a[6][24] ), .A7(\mem_a[7][24] ), .Z(n1334));
Q_MX04 U1332 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1334), .A1(n1333), .A2(n1332), .A3(n1331), .Z(n86));
Q_MX08 U1333 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][25] ), .A1(\mem_a[25][25] ), .A2(\mem_a[26][25] ), .A3(\mem_a[27][25] ), .A4(\mem_a[28][25] ), .A5(\mem_a[29][25] ), .A6(\mem_a[30][25] ), .A7(\mem_a[31][25] ), .Z(n1335));
Q_MX08 U1334 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][25] ), .A1(\mem_a[17][25] ), .A2(\mem_a[18][25] ), .A3(\mem_a[19][25] ), .A4(\mem_a[20][25] ), .A5(\mem_a[21][25] ), .A6(\mem_a[22][25] ), .A7(\mem_a[23][25] ), .Z(n1336));
Q_MX08 U1335 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][25] ), .A1(\mem_a[9][25] ), .A2(\mem_a[10][25] ), .A3(\mem_a[11][25] ), .A4(\mem_a[12][25] ), .A5(\mem_a[13][25] ), .A6(\mem_a[14][25] ), .A7(\mem_a[15][25] ), .Z(n1337));
Q_MX08 U1336 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][25] ), .A1(\mem_a[1][25] ), .A2(\mem_a[2][25] ), .A3(\mem_a[3][25] ), .A4(\mem_a[4][25] ), .A5(\mem_a[5][25] ), .A6(\mem_a[6][25] ), .A7(\mem_a[7][25] ), .Z(n1338));
Q_MX04 U1337 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1338), .A1(n1337), .A2(n1336), .A3(n1335), .Z(n85));
Q_MX08 U1338 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][26] ), .A1(\mem_a[25][26] ), .A2(\mem_a[26][26] ), .A3(\mem_a[27][26] ), .A4(\mem_a[28][26] ), .A5(\mem_a[29][26] ), .A6(\mem_a[30][26] ), .A7(\mem_a[31][26] ), .Z(n1339));
Q_MX08 U1339 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][26] ), .A1(\mem_a[17][26] ), .A2(\mem_a[18][26] ), .A3(\mem_a[19][26] ), .A4(\mem_a[20][26] ), .A5(\mem_a[21][26] ), .A6(\mem_a[22][26] ), .A7(\mem_a[23][26] ), .Z(n1340));
Q_MX08 U1340 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][26] ), .A1(\mem_a[9][26] ), .A2(\mem_a[10][26] ), .A3(\mem_a[11][26] ), .A4(\mem_a[12][26] ), .A5(\mem_a[13][26] ), .A6(\mem_a[14][26] ), .A7(\mem_a[15][26] ), .Z(n1341));
Q_MX08 U1341 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][26] ), .A1(\mem_a[1][26] ), .A2(\mem_a[2][26] ), .A3(\mem_a[3][26] ), .A4(\mem_a[4][26] ), .A5(\mem_a[5][26] ), .A6(\mem_a[6][26] ), .A7(\mem_a[7][26] ), .Z(n1342));
Q_MX04 U1342 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1342), .A1(n1341), .A2(n1340), .A3(n1339), .Z(n84));
Q_MX08 U1343 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][27] ), .A1(\mem_a[25][27] ), .A2(\mem_a[26][27] ), .A3(\mem_a[27][27] ), .A4(\mem_a[28][27] ), .A5(\mem_a[29][27] ), .A6(\mem_a[30][27] ), .A7(\mem_a[31][27] ), .Z(n1343));
Q_MX08 U1344 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][27] ), .A1(\mem_a[17][27] ), .A2(\mem_a[18][27] ), .A3(\mem_a[19][27] ), .A4(\mem_a[20][27] ), .A5(\mem_a[21][27] ), .A6(\mem_a[22][27] ), .A7(\mem_a[23][27] ), .Z(n1344));
Q_MX08 U1345 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][27] ), .A1(\mem_a[9][27] ), .A2(\mem_a[10][27] ), .A3(\mem_a[11][27] ), .A4(\mem_a[12][27] ), .A5(\mem_a[13][27] ), .A6(\mem_a[14][27] ), .A7(\mem_a[15][27] ), .Z(n1345));
Q_MX08 U1346 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][27] ), .A1(\mem_a[1][27] ), .A2(\mem_a[2][27] ), .A3(\mem_a[3][27] ), .A4(\mem_a[4][27] ), .A5(\mem_a[5][27] ), .A6(\mem_a[6][27] ), .A7(\mem_a[7][27] ), .Z(n1346));
Q_MX04 U1347 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1346), .A1(n1345), .A2(n1344), .A3(n1343), .Z(n83));
Q_MX08 U1348 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][28] ), .A1(\mem_a[25][28] ), .A2(\mem_a[26][28] ), .A3(\mem_a[27][28] ), .A4(\mem_a[28][28] ), .A5(\mem_a[29][28] ), .A6(\mem_a[30][28] ), .A7(\mem_a[31][28] ), .Z(n1347));
Q_MX08 U1349 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][28] ), .A1(\mem_a[17][28] ), .A2(\mem_a[18][28] ), .A3(\mem_a[19][28] ), .A4(\mem_a[20][28] ), .A5(\mem_a[21][28] ), .A6(\mem_a[22][28] ), .A7(\mem_a[23][28] ), .Z(n1348));
Q_MX08 U1350 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][28] ), .A1(\mem_a[9][28] ), .A2(\mem_a[10][28] ), .A3(\mem_a[11][28] ), .A4(\mem_a[12][28] ), .A5(\mem_a[13][28] ), .A6(\mem_a[14][28] ), .A7(\mem_a[15][28] ), .Z(n1349));
Q_MX08 U1351 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][28] ), .A1(\mem_a[1][28] ), .A2(\mem_a[2][28] ), .A3(\mem_a[3][28] ), .A4(\mem_a[4][28] ), .A5(\mem_a[5][28] ), .A6(\mem_a[6][28] ), .A7(\mem_a[7][28] ), .Z(n1350));
Q_MX04 U1352 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1350), .A1(n1349), .A2(n1348), .A3(n1347), .Z(n82));
Q_MX08 U1353 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][29] ), .A1(\mem_a[25][29] ), .A2(\mem_a[26][29] ), .A3(\mem_a[27][29] ), .A4(\mem_a[28][29] ), .A5(\mem_a[29][29] ), .A6(\mem_a[30][29] ), .A7(\mem_a[31][29] ), .Z(n1351));
Q_MX08 U1354 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][29] ), .A1(\mem_a[17][29] ), .A2(\mem_a[18][29] ), .A3(\mem_a[19][29] ), .A4(\mem_a[20][29] ), .A5(\mem_a[21][29] ), .A6(\mem_a[22][29] ), .A7(\mem_a[23][29] ), .Z(n1352));
Q_MX08 U1355 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][29] ), .A1(\mem_a[9][29] ), .A2(\mem_a[10][29] ), .A3(\mem_a[11][29] ), .A4(\mem_a[12][29] ), .A5(\mem_a[13][29] ), .A6(\mem_a[14][29] ), .A7(\mem_a[15][29] ), .Z(n1353));
Q_MX08 U1356 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][29] ), .A1(\mem_a[1][29] ), .A2(\mem_a[2][29] ), .A3(\mem_a[3][29] ), .A4(\mem_a[4][29] ), .A5(\mem_a[5][29] ), .A6(\mem_a[6][29] ), .A7(\mem_a[7][29] ), .Z(n1354));
Q_MX04 U1357 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1354), .A1(n1353), .A2(n1352), .A3(n1351), .Z(n81));
Q_MX08 U1358 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][30] ), .A1(\mem_a[25][30] ), .A2(\mem_a[26][30] ), .A3(\mem_a[27][30] ), .A4(\mem_a[28][30] ), .A5(\mem_a[29][30] ), .A6(\mem_a[30][30] ), .A7(\mem_a[31][30] ), .Z(n1355));
Q_MX08 U1359 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][30] ), .A1(\mem_a[17][30] ), .A2(\mem_a[18][30] ), .A3(\mem_a[19][30] ), .A4(\mem_a[20][30] ), .A5(\mem_a[21][30] ), .A6(\mem_a[22][30] ), .A7(\mem_a[23][30] ), .Z(n1356));
Q_MX08 U1360 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][30] ), .A1(\mem_a[9][30] ), .A2(\mem_a[10][30] ), .A3(\mem_a[11][30] ), .A4(\mem_a[12][30] ), .A5(\mem_a[13][30] ), .A6(\mem_a[14][30] ), .A7(\mem_a[15][30] ), .Z(n1357));
Q_MX08 U1361 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][30] ), .A1(\mem_a[1][30] ), .A2(\mem_a[2][30] ), .A3(\mem_a[3][30] ), .A4(\mem_a[4][30] ), .A5(\mem_a[5][30] ), .A6(\mem_a[6][30] ), .A7(\mem_a[7][30] ), .Z(n1358));
Q_MX04 U1362 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1358), .A1(n1357), .A2(n1356), .A3(n1355), .Z(n80));
Q_MX08 U1363 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][31] ), .A1(\mem_a[25][31] ), .A2(\mem_a[26][31] ), .A3(\mem_a[27][31] ), .A4(\mem_a[28][31] ), .A5(\mem_a[29][31] ), .A6(\mem_a[30][31] ), .A7(\mem_a[31][31] ), .Z(n1359));
Q_MX08 U1364 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][31] ), .A1(\mem_a[17][31] ), .A2(\mem_a[18][31] ), .A3(\mem_a[19][31] ), .A4(\mem_a[20][31] ), .A5(\mem_a[21][31] ), .A6(\mem_a[22][31] ), .A7(\mem_a[23][31] ), .Z(n1360));
Q_MX08 U1365 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][31] ), .A1(\mem_a[9][31] ), .A2(\mem_a[10][31] ), .A3(\mem_a[11][31] ), .A4(\mem_a[12][31] ), .A5(\mem_a[13][31] ), .A6(\mem_a[14][31] ), .A7(\mem_a[15][31] ), .Z(n1361));
Q_MX08 U1366 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][31] ), .A1(\mem_a[1][31] ), .A2(\mem_a[2][31] ), .A3(\mem_a[3][31] ), .A4(\mem_a[4][31] ), .A5(\mem_a[5][31] ), .A6(\mem_a[6][31] ), .A7(\mem_a[7][31] ), .Z(n1362));
Q_MX04 U1367 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n1362), .A1(n1361), .A2(n1360), .A3(n1359), .Z(n79));
Q_FDP4EP \mem_a_REG[31][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1234), .Q(\mem_a[31][31] ));
Q_FDP4EP \mem_a_REG[31][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1233), .Q(\mem_a[31][30] ));
Q_FDP4EP \mem_a_REG[31][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1232), .Q(\mem_a[31][29] ));
Q_FDP4EP \mem_a_REG[31][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1231), .Q(\mem_a[31][28] ));
Q_FDP4EP \mem_a_REG[31][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1230), .Q(\mem_a[31][27] ));
Q_FDP4EP \mem_a_REG[31][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1229), .Q(\mem_a[31][26] ));
Q_FDP4EP \mem_a_REG[31][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1228), .Q(\mem_a[31][25] ));
Q_FDP4EP \mem_a_REG[31][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1227), .Q(\mem_a[31][24] ));
Q_FDP4EP \mem_a_REG[31][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1226), .Q(\mem_a[31][23] ));
Q_FDP4EP \mem_a_REG[31][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1225), .Q(\mem_a[31][22] ));
Q_FDP4EP \mem_a_REG[31][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1224), .Q(\mem_a[31][21] ));
Q_FDP4EP \mem_a_REG[31][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1223), .Q(\mem_a[31][20] ));
Q_FDP4EP \mem_a_REG[31][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1222), .Q(\mem_a[31][19] ));
Q_FDP4EP \mem_a_REG[31][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1221), .Q(\mem_a[31][18] ));
Q_FDP4EP \mem_a_REG[31][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1220), .Q(\mem_a[31][17] ));
Q_FDP4EP \mem_a_REG[31][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1219), .Q(\mem_a[31][16] ));
Q_FDP4EP \mem_a_REG[31][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1218), .Q(\mem_a[31][15] ));
Q_FDP4EP \mem_a_REG[31][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1217), .Q(\mem_a[31][14] ));
Q_FDP4EP \mem_a_REG[31][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1216), .Q(\mem_a[31][13] ));
Q_FDP4EP \mem_a_REG[31][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1215), .Q(\mem_a[31][12] ));
Q_FDP4EP \mem_a_REG[31][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1214), .Q(\mem_a[31][11] ));
Q_FDP4EP \mem_a_REG[31][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1213), .Q(\mem_a[31][10] ));
Q_FDP4EP \mem_a_REG[31][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1212), .Q(\mem_a[31][9] ));
Q_FDP4EP \mem_a_REG[31][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1211), .Q(\mem_a[31][8] ));
Q_FDP4EP \mem_a_REG[31][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1210), .Q(\mem_a[31][7] ));
Q_FDP4EP \mem_a_REG[31][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1209), .Q(\mem_a[31][6] ));
Q_FDP4EP \mem_a_REG[31][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1208), .Q(\mem_a[31][5] ));
Q_FDP4EP \mem_a_REG[31][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1207), .Q(\mem_a[31][4] ));
Q_FDP4EP \mem_a_REG[31][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1206), .Q(\mem_a[31][3] ));
Q_FDP4EP \mem_a_REG[31][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1205), .Q(\mem_a[31][2] ));
Q_FDP4EP \mem_a_REG[31][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1204), .Q(\mem_a[31][1] ));
Q_FDP4EP \mem_a_REG[31][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n1202), .R(n9), .D(n1203), .Q(\mem_a[31][0] ));
Q_FDP4EP \mem_a_REG[30][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1201), .Q(\mem_a[30][31] ));
Q_FDP4EP \mem_a_REG[30][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1200), .Q(\mem_a[30][30] ));
Q_FDP4EP \mem_a_REG[30][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1199), .Q(\mem_a[30][29] ));
Q_FDP4EP \mem_a_REG[30][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1198), .Q(\mem_a[30][28] ));
Q_FDP4EP \mem_a_REG[30][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1197), .Q(\mem_a[30][27] ));
Q_FDP4EP \mem_a_REG[30][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1196), .Q(\mem_a[30][26] ));
Q_FDP4EP \mem_a_REG[30][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1195), .Q(\mem_a[30][25] ));
Q_FDP4EP \mem_a_REG[30][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1194), .Q(\mem_a[30][24] ));
Q_FDP4EP \mem_a_REG[30][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1193), .Q(\mem_a[30][23] ));
Q_FDP4EP \mem_a_REG[30][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1192), .Q(\mem_a[30][22] ));
Q_FDP4EP \mem_a_REG[30][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1191), .Q(\mem_a[30][21] ));
Q_FDP4EP \mem_a_REG[30][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1190), .Q(\mem_a[30][20] ));
Q_FDP4EP \mem_a_REG[30][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1189), .Q(\mem_a[30][19] ));
Q_FDP4EP \mem_a_REG[30][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1188), .Q(\mem_a[30][18] ));
Q_FDP4EP \mem_a_REG[30][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1187), .Q(\mem_a[30][17] ));
Q_FDP4EP \mem_a_REG[30][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1186), .Q(\mem_a[30][16] ));
Q_FDP4EP \mem_a_REG[30][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1185), .Q(\mem_a[30][15] ));
Q_FDP4EP \mem_a_REG[30][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1184), .Q(\mem_a[30][14] ));
Q_FDP4EP \mem_a_REG[30][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1183), .Q(\mem_a[30][13] ));
Q_FDP4EP \mem_a_REG[30][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1182), .Q(\mem_a[30][12] ));
Q_FDP4EP \mem_a_REG[30][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1181), .Q(\mem_a[30][11] ));
Q_FDP4EP \mem_a_REG[30][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1180), .Q(\mem_a[30][10] ));
Q_FDP4EP \mem_a_REG[30][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1179), .Q(\mem_a[30][9] ));
Q_FDP4EP \mem_a_REG[30][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1178), .Q(\mem_a[30][8] ));
Q_FDP4EP \mem_a_REG[30][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1177), .Q(\mem_a[30][7] ));
Q_FDP4EP \mem_a_REG[30][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1176), .Q(\mem_a[30][6] ));
Q_FDP4EP \mem_a_REG[30][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1175), .Q(\mem_a[30][5] ));
Q_FDP4EP \mem_a_REG[30][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1174), .Q(\mem_a[30][4] ));
Q_FDP4EP \mem_a_REG[30][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1173), .Q(\mem_a[30][3] ));
Q_FDP4EP \mem_a_REG[30][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1172), .Q(\mem_a[30][2] ));
Q_FDP4EP \mem_a_REG[30][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1171), .Q(\mem_a[30][1] ));
Q_FDP4EP \mem_a_REG[30][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n1169), .R(n9), .D(n1170), .Q(\mem_a[30][0] ));
Q_FDP4EP \mem_a_REG[29][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1168), .Q(\mem_a[29][31] ));
Q_FDP4EP \mem_a_REG[29][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1167), .Q(\mem_a[29][30] ));
Q_FDP4EP \mem_a_REG[29][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1166), .Q(\mem_a[29][29] ));
Q_FDP4EP \mem_a_REG[29][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1165), .Q(\mem_a[29][28] ));
Q_FDP4EP \mem_a_REG[29][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1164), .Q(\mem_a[29][27] ));
Q_FDP4EP \mem_a_REG[29][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1163), .Q(\mem_a[29][26] ));
Q_FDP4EP \mem_a_REG[29][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1162), .Q(\mem_a[29][25] ));
Q_FDP4EP \mem_a_REG[29][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1161), .Q(\mem_a[29][24] ));
Q_FDP4EP \mem_a_REG[29][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1160), .Q(\mem_a[29][23] ));
Q_FDP4EP \mem_a_REG[29][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1159), .Q(\mem_a[29][22] ));
Q_FDP4EP \mem_a_REG[29][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1158), .Q(\mem_a[29][21] ));
Q_FDP4EP \mem_a_REG[29][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1157), .Q(\mem_a[29][20] ));
Q_FDP4EP \mem_a_REG[29][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1156), .Q(\mem_a[29][19] ));
Q_FDP4EP \mem_a_REG[29][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1155), .Q(\mem_a[29][18] ));
Q_FDP4EP \mem_a_REG[29][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1154), .Q(\mem_a[29][17] ));
Q_FDP4EP \mem_a_REG[29][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1153), .Q(\mem_a[29][16] ));
Q_FDP4EP \mem_a_REG[29][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1152), .Q(\mem_a[29][15] ));
Q_FDP4EP \mem_a_REG[29][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1151), .Q(\mem_a[29][14] ));
Q_FDP4EP \mem_a_REG[29][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1150), .Q(\mem_a[29][13] ));
Q_FDP4EP \mem_a_REG[29][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1149), .Q(\mem_a[29][12] ));
Q_FDP4EP \mem_a_REG[29][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1148), .Q(\mem_a[29][11] ));
Q_FDP4EP \mem_a_REG[29][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1147), .Q(\mem_a[29][10] ));
Q_FDP4EP \mem_a_REG[29][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1146), .Q(\mem_a[29][9] ));
Q_FDP4EP \mem_a_REG[29][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1145), .Q(\mem_a[29][8] ));
Q_FDP4EP \mem_a_REG[29][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1144), .Q(\mem_a[29][7] ));
Q_FDP4EP \mem_a_REG[29][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1143), .Q(\mem_a[29][6] ));
Q_FDP4EP \mem_a_REG[29][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1142), .Q(\mem_a[29][5] ));
Q_FDP4EP \mem_a_REG[29][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1141), .Q(\mem_a[29][4] ));
Q_FDP4EP \mem_a_REG[29][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1140), .Q(\mem_a[29][3] ));
Q_FDP4EP \mem_a_REG[29][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1139), .Q(\mem_a[29][2] ));
Q_FDP4EP \mem_a_REG[29][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1138), .Q(\mem_a[29][1] ));
Q_FDP4EP \mem_a_REG[29][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n1136), .R(n9), .D(n1137), .Q(\mem_a[29][0] ));
Q_FDP4EP \mem_a_REG[28][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1135), .Q(\mem_a[28][31] ));
Q_FDP4EP \mem_a_REG[28][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1134), .Q(\mem_a[28][30] ));
Q_FDP4EP \mem_a_REG[28][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1133), .Q(\mem_a[28][29] ));
Q_FDP4EP \mem_a_REG[28][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1132), .Q(\mem_a[28][28] ));
Q_FDP4EP \mem_a_REG[28][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1131), .Q(\mem_a[28][27] ));
Q_FDP4EP \mem_a_REG[28][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1130), .Q(\mem_a[28][26] ));
Q_FDP4EP \mem_a_REG[28][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1129), .Q(\mem_a[28][25] ));
Q_FDP4EP \mem_a_REG[28][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1128), .Q(\mem_a[28][24] ));
Q_FDP4EP \mem_a_REG[28][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1127), .Q(\mem_a[28][23] ));
Q_FDP4EP \mem_a_REG[28][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1126), .Q(\mem_a[28][22] ));
Q_FDP4EP \mem_a_REG[28][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1125), .Q(\mem_a[28][21] ));
Q_FDP4EP \mem_a_REG[28][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1124), .Q(\mem_a[28][20] ));
Q_FDP4EP \mem_a_REG[28][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1123), .Q(\mem_a[28][19] ));
Q_FDP4EP \mem_a_REG[28][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1122), .Q(\mem_a[28][18] ));
Q_FDP4EP \mem_a_REG[28][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1121), .Q(\mem_a[28][17] ));
Q_FDP4EP \mem_a_REG[28][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1120), .Q(\mem_a[28][16] ));
Q_FDP4EP \mem_a_REG[28][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1119), .Q(\mem_a[28][15] ));
Q_FDP4EP \mem_a_REG[28][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1118), .Q(\mem_a[28][14] ));
Q_FDP4EP \mem_a_REG[28][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1117), .Q(\mem_a[28][13] ));
Q_FDP4EP \mem_a_REG[28][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1116), .Q(\mem_a[28][12] ));
Q_FDP4EP \mem_a_REG[28][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1115), .Q(\mem_a[28][11] ));
Q_FDP4EP \mem_a_REG[28][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1114), .Q(\mem_a[28][10] ));
Q_FDP4EP \mem_a_REG[28][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1113), .Q(\mem_a[28][9] ));
Q_FDP4EP \mem_a_REG[28][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1112), .Q(\mem_a[28][8] ));
Q_FDP4EP \mem_a_REG[28][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1111), .Q(\mem_a[28][7] ));
Q_FDP4EP \mem_a_REG[28][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1110), .Q(\mem_a[28][6] ));
Q_FDP4EP \mem_a_REG[28][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1109), .Q(\mem_a[28][5] ));
Q_FDP4EP \mem_a_REG[28][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1108), .Q(\mem_a[28][4] ));
Q_FDP4EP \mem_a_REG[28][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1107), .Q(\mem_a[28][3] ));
Q_FDP4EP \mem_a_REG[28][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1106), .Q(\mem_a[28][2] ));
Q_FDP4EP \mem_a_REG[28][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1105), .Q(\mem_a[28][1] ));
Q_FDP4EP \mem_a_REG[28][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n1103), .R(n9), .D(n1104), .Q(\mem_a[28][0] ));
Q_FDP4EP \mem_a_REG[27][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1102), .Q(\mem_a[27][31] ));
Q_FDP4EP \mem_a_REG[27][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1101), .Q(\mem_a[27][30] ));
Q_FDP4EP \mem_a_REG[27][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1100), .Q(\mem_a[27][29] ));
Q_FDP4EP \mem_a_REG[27][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1099), .Q(\mem_a[27][28] ));
Q_FDP4EP \mem_a_REG[27][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1098), .Q(\mem_a[27][27] ));
Q_FDP4EP \mem_a_REG[27][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1097), .Q(\mem_a[27][26] ));
Q_FDP4EP \mem_a_REG[27][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1096), .Q(\mem_a[27][25] ));
Q_FDP4EP \mem_a_REG[27][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1095), .Q(\mem_a[27][24] ));
Q_FDP4EP \mem_a_REG[27][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1094), .Q(\mem_a[27][23] ));
Q_FDP4EP \mem_a_REG[27][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1093), .Q(\mem_a[27][22] ));
Q_FDP4EP \mem_a_REG[27][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1092), .Q(\mem_a[27][21] ));
Q_FDP4EP \mem_a_REG[27][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1091), .Q(\mem_a[27][20] ));
Q_FDP4EP \mem_a_REG[27][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1090), .Q(\mem_a[27][19] ));
Q_FDP4EP \mem_a_REG[27][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1089), .Q(\mem_a[27][18] ));
Q_FDP4EP \mem_a_REG[27][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1088), .Q(\mem_a[27][17] ));
Q_FDP4EP \mem_a_REG[27][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1087), .Q(\mem_a[27][16] ));
Q_FDP4EP \mem_a_REG[27][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1086), .Q(\mem_a[27][15] ));
Q_FDP4EP \mem_a_REG[27][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1085), .Q(\mem_a[27][14] ));
Q_FDP4EP \mem_a_REG[27][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1084), .Q(\mem_a[27][13] ));
Q_FDP4EP \mem_a_REG[27][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1083), .Q(\mem_a[27][12] ));
Q_FDP4EP \mem_a_REG[27][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1082), .Q(\mem_a[27][11] ));
Q_FDP4EP \mem_a_REG[27][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1081), .Q(\mem_a[27][10] ));
Q_FDP4EP \mem_a_REG[27][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1080), .Q(\mem_a[27][9] ));
Q_FDP4EP \mem_a_REG[27][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1079), .Q(\mem_a[27][8] ));
Q_FDP4EP \mem_a_REG[27][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1078), .Q(\mem_a[27][7] ));
Q_FDP4EP \mem_a_REG[27][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1077), .Q(\mem_a[27][6] ));
Q_FDP4EP \mem_a_REG[27][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1076), .Q(\mem_a[27][5] ));
Q_FDP4EP \mem_a_REG[27][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1075), .Q(\mem_a[27][4] ));
Q_FDP4EP \mem_a_REG[27][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1074), .Q(\mem_a[27][3] ));
Q_FDP4EP \mem_a_REG[27][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1073), .Q(\mem_a[27][2] ));
Q_FDP4EP \mem_a_REG[27][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1072), .Q(\mem_a[27][1] ));
Q_FDP4EP \mem_a_REG[27][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n1070), .R(n9), .D(n1071), .Q(\mem_a[27][0] ));
Q_FDP4EP \mem_a_REG[26][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1069), .Q(\mem_a[26][31] ));
Q_FDP4EP \mem_a_REG[26][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1068), .Q(\mem_a[26][30] ));
Q_FDP4EP \mem_a_REG[26][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1067), .Q(\mem_a[26][29] ));
Q_FDP4EP \mem_a_REG[26][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1066), .Q(\mem_a[26][28] ));
Q_FDP4EP \mem_a_REG[26][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1065), .Q(\mem_a[26][27] ));
Q_FDP4EP \mem_a_REG[26][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1064), .Q(\mem_a[26][26] ));
Q_FDP4EP \mem_a_REG[26][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1063), .Q(\mem_a[26][25] ));
Q_FDP4EP \mem_a_REG[26][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1062), .Q(\mem_a[26][24] ));
Q_FDP4EP \mem_a_REG[26][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1061), .Q(\mem_a[26][23] ));
Q_FDP4EP \mem_a_REG[26][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1060), .Q(\mem_a[26][22] ));
Q_FDP4EP \mem_a_REG[26][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1059), .Q(\mem_a[26][21] ));
Q_FDP4EP \mem_a_REG[26][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1058), .Q(\mem_a[26][20] ));
Q_FDP4EP \mem_a_REG[26][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1057), .Q(\mem_a[26][19] ));
Q_FDP4EP \mem_a_REG[26][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1056), .Q(\mem_a[26][18] ));
Q_FDP4EP \mem_a_REG[26][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1055), .Q(\mem_a[26][17] ));
Q_FDP4EP \mem_a_REG[26][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1054), .Q(\mem_a[26][16] ));
Q_FDP4EP \mem_a_REG[26][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1053), .Q(\mem_a[26][15] ));
Q_FDP4EP \mem_a_REG[26][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1052), .Q(\mem_a[26][14] ));
Q_FDP4EP \mem_a_REG[26][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1051), .Q(\mem_a[26][13] ));
Q_FDP4EP \mem_a_REG[26][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1050), .Q(\mem_a[26][12] ));
Q_FDP4EP \mem_a_REG[26][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1049), .Q(\mem_a[26][11] ));
Q_FDP4EP \mem_a_REG[26][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1048), .Q(\mem_a[26][10] ));
Q_FDP4EP \mem_a_REG[26][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1047), .Q(\mem_a[26][9] ));
Q_FDP4EP \mem_a_REG[26][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1046), .Q(\mem_a[26][8] ));
Q_FDP4EP \mem_a_REG[26][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1045), .Q(\mem_a[26][7] ));
Q_FDP4EP \mem_a_REG[26][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1044), .Q(\mem_a[26][6] ));
Q_FDP4EP \mem_a_REG[26][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1043), .Q(\mem_a[26][5] ));
Q_FDP4EP \mem_a_REG[26][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1042), .Q(\mem_a[26][4] ));
Q_FDP4EP \mem_a_REG[26][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1041), .Q(\mem_a[26][3] ));
Q_FDP4EP \mem_a_REG[26][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1040), .Q(\mem_a[26][2] ));
Q_FDP4EP \mem_a_REG[26][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1039), .Q(\mem_a[26][1] ));
Q_FDP4EP \mem_a_REG[26][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n1037), .R(n9), .D(n1038), .Q(\mem_a[26][0] ));
Q_FDP4EP \mem_a_REG[25][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1036), .Q(\mem_a[25][31] ));
Q_FDP4EP \mem_a_REG[25][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1035), .Q(\mem_a[25][30] ));
Q_FDP4EP \mem_a_REG[25][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1034), .Q(\mem_a[25][29] ));
Q_FDP4EP \mem_a_REG[25][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1033), .Q(\mem_a[25][28] ));
Q_FDP4EP \mem_a_REG[25][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1032), .Q(\mem_a[25][27] ));
Q_FDP4EP \mem_a_REG[25][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1031), .Q(\mem_a[25][26] ));
Q_FDP4EP \mem_a_REG[25][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1030), .Q(\mem_a[25][25] ));
Q_FDP4EP \mem_a_REG[25][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1029), .Q(\mem_a[25][24] ));
Q_FDP4EP \mem_a_REG[25][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1028), .Q(\mem_a[25][23] ));
Q_FDP4EP \mem_a_REG[25][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1027), .Q(\mem_a[25][22] ));
Q_FDP4EP \mem_a_REG[25][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1026), .Q(\mem_a[25][21] ));
Q_FDP4EP \mem_a_REG[25][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1025), .Q(\mem_a[25][20] ));
Q_FDP4EP \mem_a_REG[25][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1024), .Q(\mem_a[25][19] ));
Q_FDP4EP \mem_a_REG[25][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1023), .Q(\mem_a[25][18] ));
Q_FDP4EP \mem_a_REG[25][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1022), .Q(\mem_a[25][17] ));
Q_FDP4EP \mem_a_REG[25][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1021), .Q(\mem_a[25][16] ));
Q_FDP4EP \mem_a_REG[25][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1020), .Q(\mem_a[25][15] ));
Q_FDP4EP \mem_a_REG[25][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1019), .Q(\mem_a[25][14] ));
Q_FDP4EP \mem_a_REG[25][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1018), .Q(\mem_a[25][13] ));
Q_FDP4EP \mem_a_REG[25][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1017), .Q(\mem_a[25][12] ));
Q_FDP4EP \mem_a_REG[25][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1016), .Q(\mem_a[25][11] ));
Q_FDP4EP \mem_a_REG[25][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1015), .Q(\mem_a[25][10] ));
Q_FDP4EP \mem_a_REG[25][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1014), .Q(\mem_a[25][9] ));
Q_FDP4EP \mem_a_REG[25][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1013), .Q(\mem_a[25][8] ));
Q_FDP4EP \mem_a_REG[25][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1012), .Q(\mem_a[25][7] ));
Q_FDP4EP \mem_a_REG[25][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1011), .Q(\mem_a[25][6] ));
Q_FDP4EP \mem_a_REG[25][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1010), .Q(\mem_a[25][5] ));
Q_FDP4EP \mem_a_REG[25][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1009), .Q(\mem_a[25][4] ));
Q_FDP4EP \mem_a_REG[25][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1008), .Q(\mem_a[25][3] ));
Q_FDP4EP \mem_a_REG[25][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1007), .Q(\mem_a[25][2] ));
Q_FDP4EP \mem_a_REG[25][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1006), .Q(\mem_a[25][1] ));
Q_FDP4EP \mem_a_REG[25][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n1004), .R(n9), .D(n1005), .Q(\mem_a[25][0] ));
Q_FDP4EP \mem_a_REG[24][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n1003), .Q(\mem_a[24][31] ));
Q_FDP4EP \mem_a_REG[24][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n1002), .Q(\mem_a[24][30] ));
Q_FDP4EP \mem_a_REG[24][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n1001), .Q(\mem_a[24][29] ));
Q_FDP4EP \mem_a_REG[24][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n1000), .Q(\mem_a[24][28] ));
Q_FDP4EP \mem_a_REG[24][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n999), .Q(\mem_a[24][27] ));
Q_FDP4EP \mem_a_REG[24][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n998), .Q(\mem_a[24][26] ));
Q_FDP4EP \mem_a_REG[24][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n997), .Q(\mem_a[24][25] ));
Q_FDP4EP \mem_a_REG[24][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n996), .Q(\mem_a[24][24] ));
Q_FDP4EP \mem_a_REG[24][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n995), .Q(\mem_a[24][23] ));
Q_FDP4EP \mem_a_REG[24][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n994), .Q(\mem_a[24][22] ));
Q_FDP4EP \mem_a_REG[24][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n993), .Q(\mem_a[24][21] ));
Q_FDP4EP \mem_a_REG[24][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n992), .Q(\mem_a[24][20] ));
Q_FDP4EP \mem_a_REG[24][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n991), .Q(\mem_a[24][19] ));
Q_FDP4EP \mem_a_REG[24][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n990), .Q(\mem_a[24][18] ));
Q_FDP4EP \mem_a_REG[24][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n989), .Q(\mem_a[24][17] ));
Q_FDP4EP \mem_a_REG[24][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n988), .Q(\mem_a[24][16] ));
Q_FDP4EP \mem_a_REG[24][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n987), .Q(\mem_a[24][15] ));
Q_FDP4EP \mem_a_REG[24][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n986), .Q(\mem_a[24][14] ));
Q_FDP4EP \mem_a_REG[24][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n985), .Q(\mem_a[24][13] ));
Q_FDP4EP \mem_a_REG[24][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n984), .Q(\mem_a[24][12] ));
Q_FDP4EP \mem_a_REG[24][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n983), .Q(\mem_a[24][11] ));
Q_FDP4EP \mem_a_REG[24][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n982), .Q(\mem_a[24][10] ));
Q_FDP4EP \mem_a_REG[24][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n981), .Q(\mem_a[24][9] ));
Q_FDP4EP \mem_a_REG[24][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n980), .Q(\mem_a[24][8] ));
Q_FDP4EP \mem_a_REG[24][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n979), .Q(\mem_a[24][7] ));
Q_FDP4EP \mem_a_REG[24][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n978), .Q(\mem_a[24][6] ));
Q_FDP4EP \mem_a_REG[24][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n977), .Q(\mem_a[24][5] ));
Q_FDP4EP \mem_a_REG[24][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n976), .Q(\mem_a[24][4] ));
Q_FDP4EP \mem_a_REG[24][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n975), .Q(\mem_a[24][3] ));
Q_FDP4EP \mem_a_REG[24][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n974), .Q(\mem_a[24][2] ));
Q_FDP4EP \mem_a_REG[24][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n973), .Q(\mem_a[24][1] ));
Q_FDP4EP \mem_a_REG[24][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n971), .R(n9), .D(n972), .Q(\mem_a[24][0] ));
Q_FDP4EP \mem_a_REG[23][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n970), .Q(\mem_a[23][31] ));
Q_FDP4EP \mem_a_REG[23][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n969), .Q(\mem_a[23][30] ));
Q_FDP4EP \mem_a_REG[23][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n968), .Q(\mem_a[23][29] ));
Q_FDP4EP \mem_a_REG[23][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n967), .Q(\mem_a[23][28] ));
Q_FDP4EP \mem_a_REG[23][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n966), .Q(\mem_a[23][27] ));
Q_FDP4EP \mem_a_REG[23][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n965), .Q(\mem_a[23][26] ));
Q_FDP4EP \mem_a_REG[23][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n964), .Q(\mem_a[23][25] ));
Q_FDP4EP \mem_a_REG[23][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n963), .Q(\mem_a[23][24] ));
Q_FDP4EP \mem_a_REG[23][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n962), .Q(\mem_a[23][23] ));
Q_FDP4EP \mem_a_REG[23][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n961), .Q(\mem_a[23][22] ));
Q_FDP4EP \mem_a_REG[23][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n960), .Q(\mem_a[23][21] ));
Q_FDP4EP \mem_a_REG[23][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n959), .Q(\mem_a[23][20] ));
Q_FDP4EP \mem_a_REG[23][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n958), .Q(\mem_a[23][19] ));
Q_FDP4EP \mem_a_REG[23][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n957), .Q(\mem_a[23][18] ));
Q_FDP4EP \mem_a_REG[23][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n956), .Q(\mem_a[23][17] ));
Q_FDP4EP \mem_a_REG[23][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n955), .Q(\mem_a[23][16] ));
Q_FDP4EP \mem_a_REG[23][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n954), .Q(\mem_a[23][15] ));
Q_FDP4EP \mem_a_REG[23][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n953), .Q(\mem_a[23][14] ));
Q_FDP4EP \mem_a_REG[23][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n952), .Q(\mem_a[23][13] ));
Q_FDP4EP \mem_a_REG[23][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n951), .Q(\mem_a[23][12] ));
Q_FDP4EP \mem_a_REG[23][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n950), .Q(\mem_a[23][11] ));
Q_FDP4EP \mem_a_REG[23][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n949), .Q(\mem_a[23][10] ));
Q_FDP4EP \mem_a_REG[23][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n948), .Q(\mem_a[23][9] ));
Q_FDP4EP \mem_a_REG[23][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n947), .Q(\mem_a[23][8] ));
Q_FDP4EP \mem_a_REG[23][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n946), .Q(\mem_a[23][7] ));
Q_FDP4EP \mem_a_REG[23][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n945), .Q(\mem_a[23][6] ));
Q_FDP4EP \mem_a_REG[23][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n944), .Q(\mem_a[23][5] ));
Q_FDP4EP \mem_a_REG[23][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n943), .Q(\mem_a[23][4] ));
Q_FDP4EP \mem_a_REG[23][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n942), .Q(\mem_a[23][3] ));
Q_FDP4EP \mem_a_REG[23][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n941), .Q(\mem_a[23][2] ));
Q_FDP4EP \mem_a_REG[23][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n940), .Q(\mem_a[23][1] ));
Q_FDP4EP \mem_a_REG[23][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n938), .R(n9), .D(n939), .Q(\mem_a[23][0] ));
Q_FDP4EP \mem_a_REG[22][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n937), .Q(\mem_a[22][31] ));
Q_FDP4EP \mem_a_REG[22][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n936), .Q(\mem_a[22][30] ));
Q_FDP4EP \mem_a_REG[22][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n935), .Q(\mem_a[22][29] ));
Q_FDP4EP \mem_a_REG[22][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n934), .Q(\mem_a[22][28] ));
Q_FDP4EP \mem_a_REG[22][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n933), .Q(\mem_a[22][27] ));
Q_FDP4EP \mem_a_REG[22][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n932), .Q(\mem_a[22][26] ));
Q_FDP4EP \mem_a_REG[22][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n931), .Q(\mem_a[22][25] ));
Q_FDP4EP \mem_a_REG[22][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n930), .Q(\mem_a[22][24] ));
Q_FDP4EP \mem_a_REG[22][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n929), .Q(\mem_a[22][23] ));
Q_FDP4EP \mem_a_REG[22][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n928), .Q(\mem_a[22][22] ));
Q_FDP4EP \mem_a_REG[22][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n927), .Q(\mem_a[22][21] ));
Q_FDP4EP \mem_a_REG[22][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n926), .Q(\mem_a[22][20] ));
Q_FDP4EP \mem_a_REG[22][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n925), .Q(\mem_a[22][19] ));
Q_FDP4EP \mem_a_REG[22][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n924), .Q(\mem_a[22][18] ));
Q_FDP4EP \mem_a_REG[22][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n923), .Q(\mem_a[22][17] ));
Q_FDP4EP \mem_a_REG[22][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n922), .Q(\mem_a[22][16] ));
Q_FDP4EP \mem_a_REG[22][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n921), .Q(\mem_a[22][15] ));
Q_FDP4EP \mem_a_REG[22][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n920), .Q(\mem_a[22][14] ));
Q_FDP4EP \mem_a_REG[22][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n919), .Q(\mem_a[22][13] ));
Q_FDP4EP \mem_a_REG[22][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n918), .Q(\mem_a[22][12] ));
Q_FDP4EP \mem_a_REG[22][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n917), .Q(\mem_a[22][11] ));
Q_FDP4EP \mem_a_REG[22][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n916), .Q(\mem_a[22][10] ));
Q_FDP4EP \mem_a_REG[22][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n915), .Q(\mem_a[22][9] ));
Q_FDP4EP \mem_a_REG[22][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n914), .Q(\mem_a[22][8] ));
Q_FDP4EP \mem_a_REG[22][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n913), .Q(\mem_a[22][7] ));
Q_FDP4EP \mem_a_REG[22][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n912), .Q(\mem_a[22][6] ));
Q_FDP4EP \mem_a_REG[22][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n911), .Q(\mem_a[22][5] ));
Q_FDP4EP \mem_a_REG[22][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n910), .Q(\mem_a[22][4] ));
Q_FDP4EP \mem_a_REG[22][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n909), .Q(\mem_a[22][3] ));
Q_FDP4EP \mem_a_REG[22][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n908), .Q(\mem_a[22][2] ));
Q_FDP4EP \mem_a_REG[22][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n907), .Q(\mem_a[22][1] ));
Q_FDP4EP \mem_a_REG[22][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n905), .R(n9), .D(n906), .Q(\mem_a[22][0] ));
Q_FDP4EP \mem_a_REG[21][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n904), .Q(\mem_a[21][31] ));
Q_FDP4EP \mem_a_REG[21][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n903), .Q(\mem_a[21][30] ));
Q_FDP4EP \mem_a_REG[21][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n902), .Q(\mem_a[21][29] ));
Q_FDP4EP \mem_a_REG[21][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n901), .Q(\mem_a[21][28] ));
Q_FDP4EP \mem_a_REG[21][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n900), .Q(\mem_a[21][27] ));
Q_FDP4EP \mem_a_REG[21][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n899), .Q(\mem_a[21][26] ));
Q_FDP4EP \mem_a_REG[21][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n898), .Q(\mem_a[21][25] ));
Q_FDP4EP \mem_a_REG[21][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n897), .Q(\mem_a[21][24] ));
Q_FDP4EP \mem_a_REG[21][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n896), .Q(\mem_a[21][23] ));
Q_FDP4EP \mem_a_REG[21][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n895), .Q(\mem_a[21][22] ));
Q_FDP4EP \mem_a_REG[21][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n894), .Q(\mem_a[21][21] ));
Q_FDP4EP \mem_a_REG[21][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n893), .Q(\mem_a[21][20] ));
Q_FDP4EP \mem_a_REG[21][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n892), .Q(\mem_a[21][19] ));
Q_FDP4EP \mem_a_REG[21][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n891), .Q(\mem_a[21][18] ));
Q_FDP4EP \mem_a_REG[21][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n890), .Q(\mem_a[21][17] ));
Q_FDP4EP \mem_a_REG[21][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n889), .Q(\mem_a[21][16] ));
Q_FDP4EP \mem_a_REG[21][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n888), .Q(\mem_a[21][15] ));
Q_FDP4EP \mem_a_REG[21][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n887), .Q(\mem_a[21][14] ));
Q_FDP4EP \mem_a_REG[21][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n886), .Q(\mem_a[21][13] ));
Q_FDP4EP \mem_a_REG[21][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n885), .Q(\mem_a[21][12] ));
Q_FDP4EP \mem_a_REG[21][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n884), .Q(\mem_a[21][11] ));
Q_FDP4EP \mem_a_REG[21][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n883), .Q(\mem_a[21][10] ));
Q_FDP4EP \mem_a_REG[21][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n882), .Q(\mem_a[21][9] ));
Q_FDP4EP \mem_a_REG[21][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n881), .Q(\mem_a[21][8] ));
Q_FDP4EP \mem_a_REG[21][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n880), .Q(\mem_a[21][7] ));
Q_FDP4EP \mem_a_REG[21][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n879), .Q(\mem_a[21][6] ));
Q_FDP4EP \mem_a_REG[21][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n878), .Q(\mem_a[21][5] ));
Q_FDP4EP \mem_a_REG[21][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n877), .Q(\mem_a[21][4] ));
Q_FDP4EP \mem_a_REG[21][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n876), .Q(\mem_a[21][3] ));
Q_FDP4EP \mem_a_REG[21][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n875), .Q(\mem_a[21][2] ));
Q_FDP4EP \mem_a_REG[21][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n874), .Q(\mem_a[21][1] ));
Q_FDP4EP \mem_a_REG[21][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n872), .R(n9), .D(n873), .Q(\mem_a[21][0] ));
Q_FDP4EP \mem_a_REG[20][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n871), .Q(\mem_a[20][31] ));
Q_FDP4EP \mem_a_REG[20][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n870), .Q(\mem_a[20][30] ));
Q_FDP4EP \mem_a_REG[20][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n869), .Q(\mem_a[20][29] ));
Q_FDP4EP \mem_a_REG[20][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n868), .Q(\mem_a[20][28] ));
Q_FDP4EP \mem_a_REG[20][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n867), .Q(\mem_a[20][27] ));
Q_FDP4EP \mem_a_REG[20][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n866), .Q(\mem_a[20][26] ));
Q_FDP4EP \mem_a_REG[20][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n865), .Q(\mem_a[20][25] ));
Q_FDP4EP \mem_a_REG[20][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n864), .Q(\mem_a[20][24] ));
Q_FDP4EP \mem_a_REG[20][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n863), .Q(\mem_a[20][23] ));
Q_FDP4EP \mem_a_REG[20][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n862), .Q(\mem_a[20][22] ));
Q_FDP4EP \mem_a_REG[20][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n861), .Q(\mem_a[20][21] ));
Q_FDP4EP \mem_a_REG[20][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n860), .Q(\mem_a[20][20] ));
Q_FDP4EP \mem_a_REG[20][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n859), .Q(\mem_a[20][19] ));
Q_FDP4EP \mem_a_REG[20][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n858), .Q(\mem_a[20][18] ));
Q_FDP4EP \mem_a_REG[20][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n857), .Q(\mem_a[20][17] ));
Q_FDP4EP \mem_a_REG[20][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n856), .Q(\mem_a[20][16] ));
Q_FDP4EP \mem_a_REG[20][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n855), .Q(\mem_a[20][15] ));
Q_FDP4EP \mem_a_REG[20][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n854), .Q(\mem_a[20][14] ));
Q_FDP4EP \mem_a_REG[20][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n853), .Q(\mem_a[20][13] ));
Q_FDP4EP \mem_a_REG[20][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n852), .Q(\mem_a[20][12] ));
Q_FDP4EP \mem_a_REG[20][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n851), .Q(\mem_a[20][11] ));
Q_FDP4EP \mem_a_REG[20][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n850), .Q(\mem_a[20][10] ));
Q_FDP4EP \mem_a_REG[20][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n849), .Q(\mem_a[20][9] ));
Q_FDP4EP \mem_a_REG[20][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n848), .Q(\mem_a[20][8] ));
Q_FDP4EP \mem_a_REG[20][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n847), .Q(\mem_a[20][7] ));
Q_FDP4EP \mem_a_REG[20][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n846), .Q(\mem_a[20][6] ));
Q_FDP4EP \mem_a_REG[20][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n845), .Q(\mem_a[20][5] ));
Q_FDP4EP \mem_a_REG[20][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n844), .Q(\mem_a[20][4] ));
Q_FDP4EP \mem_a_REG[20][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n843), .Q(\mem_a[20][3] ));
Q_FDP4EP \mem_a_REG[20][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n842), .Q(\mem_a[20][2] ));
Q_FDP4EP \mem_a_REG[20][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n841), .Q(\mem_a[20][1] ));
Q_FDP4EP \mem_a_REG[20][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n839), .R(n9), .D(n840), .Q(\mem_a[20][0] ));
Q_FDP4EP \mem_a_REG[19][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n838), .Q(\mem_a[19][31] ));
Q_FDP4EP \mem_a_REG[19][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n837), .Q(\mem_a[19][30] ));
Q_FDP4EP \mem_a_REG[19][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n836), .Q(\mem_a[19][29] ));
Q_FDP4EP \mem_a_REG[19][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n835), .Q(\mem_a[19][28] ));
Q_FDP4EP \mem_a_REG[19][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n834), .Q(\mem_a[19][27] ));
Q_FDP4EP \mem_a_REG[19][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n833), .Q(\mem_a[19][26] ));
Q_FDP4EP \mem_a_REG[19][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n832), .Q(\mem_a[19][25] ));
Q_FDP4EP \mem_a_REG[19][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n831), .Q(\mem_a[19][24] ));
Q_FDP4EP \mem_a_REG[19][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n830), .Q(\mem_a[19][23] ));
Q_FDP4EP \mem_a_REG[19][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n829), .Q(\mem_a[19][22] ));
Q_FDP4EP \mem_a_REG[19][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n828), .Q(\mem_a[19][21] ));
Q_FDP4EP \mem_a_REG[19][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n827), .Q(\mem_a[19][20] ));
Q_FDP4EP \mem_a_REG[19][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n826), .Q(\mem_a[19][19] ));
Q_FDP4EP \mem_a_REG[19][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n825), .Q(\mem_a[19][18] ));
Q_FDP4EP \mem_a_REG[19][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n824), .Q(\mem_a[19][17] ));
Q_FDP4EP \mem_a_REG[19][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n823), .Q(\mem_a[19][16] ));
Q_FDP4EP \mem_a_REG[19][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n822), .Q(\mem_a[19][15] ));
Q_FDP4EP \mem_a_REG[19][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n821), .Q(\mem_a[19][14] ));
Q_FDP4EP \mem_a_REG[19][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n820), .Q(\mem_a[19][13] ));
Q_FDP4EP \mem_a_REG[19][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n819), .Q(\mem_a[19][12] ));
Q_FDP4EP \mem_a_REG[19][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n818), .Q(\mem_a[19][11] ));
Q_FDP4EP \mem_a_REG[19][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n817), .Q(\mem_a[19][10] ));
Q_FDP4EP \mem_a_REG[19][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n816), .Q(\mem_a[19][9] ));
Q_FDP4EP \mem_a_REG[19][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n815), .Q(\mem_a[19][8] ));
Q_FDP4EP \mem_a_REG[19][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n814), .Q(\mem_a[19][7] ));
Q_FDP4EP \mem_a_REG[19][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n813), .Q(\mem_a[19][6] ));
Q_FDP4EP \mem_a_REG[19][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n812), .Q(\mem_a[19][5] ));
Q_FDP4EP \mem_a_REG[19][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n811), .Q(\mem_a[19][4] ));
Q_FDP4EP \mem_a_REG[19][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n810), .Q(\mem_a[19][3] ));
Q_FDP4EP \mem_a_REG[19][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n809), .Q(\mem_a[19][2] ));
Q_FDP4EP \mem_a_REG[19][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n808), .Q(\mem_a[19][1] ));
Q_FDP4EP \mem_a_REG[19][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n806), .R(n9), .D(n807), .Q(\mem_a[19][0] ));
Q_FDP4EP \mem_a_REG[18][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n805), .Q(\mem_a[18][31] ));
Q_FDP4EP \mem_a_REG[18][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n804), .Q(\mem_a[18][30] ));
Q_FDP4EP \mem_a_REG[18][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n803), .Q(\mem_a[18][29] ));
Q_FDP4EP \mem_a_REG[18][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n802), .Q(\mem_a[18][28] ));
Q_FDP4EP \mem_a_REG[18][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n801), .Q(\mem_a[18][27] ));
Q_FDP4EP \mem_a_REG[18][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n800), .Q(\mem_a[18][26] ));
Q_FDP4EP \mem_a_REG[18][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n799), .Q(\mem_a[18][25] ));
Q_FDP4EP \mem_a_REG[18][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n798), .Q(\mem_a[18][24] ));
Q_FDP4EP \mem_a_REG[18][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n797), .Q(\mem_a[18][23] ));
Q_FDP4EP \mem_a_REG[18][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n796), .Q(\mem_a[18][22] ));
Q_FDP4EP \mem_a_REG[18][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n795), .Q(\mem_a[18][21] ));
Q_FDP4EP \mem_a_REG[18][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n794), .Q(\mem_a[18][20] ));
Q_FDP4EP \mem_a_REG[18][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n793), .Q(\mem_a[18][19] ));
Q_FDP4EP \mem_a_REG[18][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n792), .Q(\mem_a[18][18] ));
Q_FDP4EP \mem_a_REG[18][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n791), .Q(\mem_a[18][17] ));
Q_FDP4EP \mem_a_REG[18][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n790), .Q(\mem_a[18][16] ));
Q_FDP4EP \mem_a_REG[18][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n789), .Q(\mem_a[18][15] ));
Q_FDP4EP \mem_a_REG[18][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n788), .Q(\mem_a[18][14] ));
Q_FDP4EP \mem_a_REG[18][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n787), .Q(\mem_a[18][13] ));
Q_FDP4EP \mem_a_REG[18][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n786), .Q(\mem_a[18][12] ));
Q_FDP4EP \mem_a_REG[18][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n785), .Q(\mem_a[18][11] ));
Q_FDP4EP \mem_a_REG[18][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n784), .Q(\mem_a[18][10] ));
Q_FDP4EP \mem_a_REG[18][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n783), .Q(\mem_a[18][9] ));
Q_FDP4EP \mem_a_REG[18][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n782), .Q(\mem_a[18][8] ));
Q_FDP4EP \mem_a_REG[18][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n781), .Q(\mem_a[18][7] ));
Q_FDP4EP \mem_a_REG[18][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n780), .Q(\mem_a[18][6] ));
Q_FDP4EP \mem_a_REG[18][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n779), .Q(\mem_a[18][5] ));
Q_FDP4EP \mem_a_REG[18][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n778), .Q(\mem_a[18][4] ));
Q_FDP4EP \mem_a_REG[18][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n777), .Q(\mem_a[18][3] ));
Q_FDP4EP \mem_a_REG[18][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n776), .Q(\mem_a[18][2] ));
Q_FDP4EP \mem_a_REG[18][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n775), .Q(\mem_a[18][1] ));
Q_FDP4EP \mem_a_REG[18][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n773), .R(n9), .D(n774), .Q(\mem_a[18][0] ));
Q_FDP4EP \mem_a_REG[17][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n772), .Q(\mem_a[17][31] ));
Q_FDP4EP \mem_a_REG[17][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n771), .Q(\mem_a[17][30] ));
Q_FDP4EP \mem_a_REG[17][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n770), .Q(\mem_a[17][29] ));
Q_FDP4EP \mem_a_REG[17][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n769), .Q(\mem_a[17][28] ));
Q_FDP4EP \mem_a_REG[17][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n768), .Q(\mem_a[17][27] ));
Q_FDP4EP \mem_a_REG[17][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n767), .Q(\mem_a[17][26] ));
Q_FDP4EP \mem_a_REG[17][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n766), .Q(\mem_a[17][25] ));
Q_FDP4EP \mem_a_REG[17][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n765), .Q(\mem_a[17][24] ));
Q_FDP4EP \mem_a_REG[17][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n764), .Q(\mem_a[17][23] ));
Q_FDP4EP \mem_a_REG[17][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n763), .Q(\mem_a[17][22] ));
Q_FDP4EP \mem_a_REG[17][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n762), .Q(\mem_a[17][21] ));
Q_FDP4EP \mem_a_REG[17][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n761), .Q(\mem_a[17][20] ));
Q_FDP4EP \mem_a_REG[17][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n760), .Q(\mem_a[17][19] ));
Q_FDP4EP \mem_a_REG[17][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n759), .Q(\mem_a[17][18] ));
Q_FDP4EP \mem_a_REG[17][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n758), .Q(\mem_a[17][17] ));
Q_FDP4EP \mem_a_REG[17][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n757), .Q(\mem_a[17][16] ));
Q_FDP4EP \mem_a_REG[17][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n756), .Q(\mem_a[17][15] ));
Q_FDP4EP \mem_a_REG[17][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n755), .Q(\mem_a[17][14] ));
Q_FDP4EP \mem_a_REG[17][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n754), .Q(\mem_a[17][13] ));
Q_FDP4EP \mem_a_REG[17][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n753), .Q(\mem_a[17][12] ));
Q_FDP4EP \mem_a_REG[17][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n752), .Q(\mem_a[17][11] ));
Q_FDP4EP \mem_a_REG[17][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n751), .Q(\mem_a[17][10] ));
Q_FDP4EP \mem_a_REG[17][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n750), .Q(\mem_a[17][9] ));
Q_FDP4EP \mem_a_REG[17][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n749), .Q(\mem_a[17][8] ));
Q_FDP4EP \mem_a_REG[17][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n748), .Q(\mem_a[17][7] ));
Q_FDP4EP \mem_a_REG[17][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n747), .Q(\mem_a[17][6] ));
Q_FDP4EP \mem_a_REG[17][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n746), .Q(\mem_a[17][5] ));
Q_FDP4EP \mem_a_REG[17][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n745), .Q(\mem_a[17][4] ));
Q_FDP4EP \mem_a_REG[17][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n744), .Q(\mem_a[17][3] ));
Q_FDP4EP \mem_a_REG[17][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n743), .Q(\mem_a[17][2] ));
Q_FDP4EP \mem_a_REG[17][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n742), .Q(\mem_a[17][1] ));
Q_FDP4EP \mem_a_REG[17][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n740), .R(n9), .D(n741), .Q(\mem_a[17][0] ));
Q_FDP4EP \mem_a_REG[16][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n739), .Q(\mem_a[16][31] ));
Q_FDP4EP \mem_a_REG[16][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n738), .Q(\mem_a[16][30] ));
Q_FDP4EP \mem_a_REG[16][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n737), .Q(\mem_a[16][29] ));
Q_FDP4EP \mem_a_REG[16][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n736), .Q(\mem_a[16][28] ));
Q_FDP4EP \mem_a_REG[16][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n735), .Q(\mem_a[16][27] ));
Q_FDP4EP \mem_a_REG[16][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n734), .Q(\mem_a[16][26] ));
Q_FDP4EP \mem_a_REG[16][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n733), .Q(\mem_a[16][25] ));
Q_FDP4EP \mem_a_REG[16][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n732), .Q(\mem_a[16][24] ));
Q_FDP4EP \mem_a_REG[16][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n731), .Q(\mem_a[16][23] ));
Q_FDP4EP \mem_a_REG[16][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n730), .Q(\mem_a[16][22] ));
Q_FDP4EP \mem_a_REG[16][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n729), .Q(\mem_a[16][21] ));
Q_FDP4EP \mem_a_REG[16][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n728), .Q(\mem_a[16][20] ));
Q_FDP4EP \mem_a_REG[16][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n727), .Q(\mem_a[16][19] ));
Q_FDP4EP \mem_a_REG[16][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n726), .Q(\mem_a[16][18] ));
Q_FDP4EP \mem_a_REG[16][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n725), .Q(\mem_a[16][17] ));
Q_FDP4EP \mem_a_REG[16][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n724), .Q(\mem_a[16][16] ));
Q_FDP4EP \mem_a_REG[16][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n723), .Q(\mem_a[16][15] ));
Q_FDP4EP \mem_a_REG[16][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n722), .Q(\mem_a[16][14] ));
Q_FDP4EP \mem_a_REG[16][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n721), .Q(\mem_a[16][13] ));
Q_FDP4EP \mem_a_REG[16][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n720), .Q(\mem_a[16][12] ));
Q_FDP4EP \mem_a_REG[16][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n719), .Q(\mem_a[16][11] ));
Q_FDP4EP \mem_a_REG[16][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n718), .Q(\mem_a[16][10] ));
Q_FDP4EP \mem_a_REG[16][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n717), .Q(\mem_a[16][9] ));
Q_FDP4EP \mem_a_REG[16][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n716), .Q(\mem_a[16][8] ));
Q_FDP4EP \mem_a_REG[16][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n715), .Q(\mem_a[16][7] ));
Q_FDP4EP \mem_a_REG[16][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n714), .Q(\mem_a[16][6] ));
Q_FDP4EP \mem_a_REG[16][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n713), .Q(\mem_a[16][5] ));
Q_FDP4EP \mem_a_REG[16][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n712), .Q(\mem_a[16][4] ));
Q_FDP4EP \mem_a_REG[16][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n711), .Q(\mem_a[16][3] ));
Q_FDP4EP \mem_a_REG[16][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n710), .Q(\mem_a[16][2] ));
Q_FDP4EP \mem_a_REG[16][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n709), .Q(\mem_a[16][1] ));
Q_FDP4EP \mem_a_REG[16][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n707), .R(n9), .D(n708), .Q(\mem_a[16][0] ));
Q_FDP4EP \mem_a_REG[15][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n706), .Q(\mem_a[15][31] ));
Q_FDP4EP \mem_a_REG[15][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n705), .Q(\mem_a[15][30] ));
Q_FDP4EP \mem_a_REG[15][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n704), .Q(\mem_a[15][29] ));
Q_FDP4EP \mem_a_REG[15][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n703), .Q(\mem_a[15][28] ));
Q_FDP4EP \mem_a_REG[15][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n702), .Q(\mem_a[15][27] ));
Q_FDP4EP \mem_a_REG[15][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n701), .Q(\mem_a[15][26] ));
Q_FDP4EP \mem_a_REG[15][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n700), .Q(\mem_a[15][25] ));
Q_FDP4EP \mem_a_REG[15][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n699), .Q(\mem_a[15][24] ));
Q_FDP4EP \mem_a_REG[15][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n698), .Q(\mem_a[15][23] ));
Q_FDP4EP \mem_a_REG[15][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n697), .Q(\mem_a[15][22] ));
Q_FDP4EP \mem_a_REG[15][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n696), .Q(\mem_a[15][21] ));
Q_FDP4EP \mem_a_REG[15][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n695), .Q(\mem_a[15][20] ));
Q_FDP4EP \mem_a_REG[15][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n694), .Q(\mem_a[15][19] ));
Q_FDP4EP \mem_a_REG[15][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n693), .Q(\mem_a[15][18] ));
Q_FDP4EP \mem_a_REG[15][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n692), .Q(\mem_a[15][17] ));
Q_FDP4EP \mem_a_REG[15][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n691), .Q(\mem_a[15][16] ));
Q_FDP4EP \mem_a_REG[15][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n690), .Q(\mem_a[15][15] ));
Q_FDP4EP \mem_a_REG[15][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n689), .Q(\mem_a[15][14] ));
Q_FDP4EP \mem_a_REG[15][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n688), .Q(\mem_a[15][13] ));
Q_FDP4EP \mem_a_REG[15][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n687), .Q(\mem_a[15][12] ));
Q_FDP4EP \mem_a_REG[15][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n686), .Q(\mem_a[15][11] ));
Q_FDP4EP \mem_a_REG[15][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n685), .Q(\mem_a[15][10] ));
Q_FDP4EP \mem_a_REG[15][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n684), .Q(\mem_a[15][9] ));
Q_FDP4EP \mem_a_REG[15][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n683), .Q(\mem_a[15][8] ));
Q_FDP4EP \mem_a_REG[15][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n682), .Q(\mem_a[15][7] ));
Q_FDP4EP \mem_a_REG[15][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n681), .Q(\mem_a[15][6] ));
Q_FDP4EP \mem_a_REG[15][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n680), .Q(\mem_a[15][5] ));
Q_FDP4EP \mem_a_REG[15][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n679), .Q(\mem_a[15][4] ));
Q_FDP4EP \mem_a_REG[15][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n678), .Q(\mem_a[15][3] ));
Q_FDP4EP \mem_a_REG[15][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n677), .Q(\mem_a[15][2] ));
Q_FDP4EP \mem_a_REG[15][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n676), .Q(\mem_a[15][1] ));
Q_FDP4EP \mem_a_REG[15][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n674), .R(n9), .D(n675), .Q(\mem_a[15][0] ));
Q_FDP4EP \mem_a_REG[14][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n673), .Q(\mem_a[14][31] ));
Q_FDP4EP \mem_a_REG[14][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n672), .Q(\mem_a[14][30] ));
Q_FDP4EP \mem_a_REG[14][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n671), .Q(\mem_a[14][29] ));
Q_FDP4EP \mem_a_REG[14][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n670), .Q(\mem_a[14][28] ));
Q_FDP4EP \mem_a_REG[14][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n669), .Q(\mem_a[14][27] ));
Q_FDP4EP \mem_a_REG[14][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n668), .Q(\mem_a[14][26] ));
Q_FDP4EP \mem_a_REG[14][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n667), .Q(\mem_a[14][25] ));
Q_FDP4EP \mem_a_REG[14][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n666), .Q(\mem_a[14][24] ));
Q_FDP4EP \mem_a_REG[14][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n665), .Q(\mem_a[14][23] ));
Q_FDP4EP \mem_a_REG[14][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n664), .Q(\mem_a[14][22] ));
Q_FDP4EP \mem_a_REG[14][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n663), .Q(\mem_a[14][21] ));
Q_FDP4EP \mem_a_REG[14][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n662), .Q(\mem_a[14][20] ));
Q_FDP4EP \mem_a_REG[14][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n661), .Q(\mem_a[14][19] ));
Q_FDP4EP \mem_a_REG[14][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n660), .Q(\mem_a[14][18] ));
Q_FDP4EP \mem_a_REG[14][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n659), .Q(\mem_a[14][17] ));
Q_FDP4EP \mem_a_REG[14][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n658), .Q(\mem_a[14][16] ));
Q_FDP4EP \mem_a_REG[14][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n657), .Q(\mem_a[14][15] ));
Q_FDP4EP \mem_a_REG[14][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n656), .Q(\mem_a[14][14] ));
Q_FDP4EP \mem_a_REG[14][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n655), .Q(\mem_a[14][13] ));
Q_FDP4EP \mem_a_REG[14][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n654), .Q(\mem_a[14][12] ));
Q_FDP4EP \mem_a_REG[14][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n653), .Q(\mem_a[14][11] ));
Q_FDP4EP \mem_a_REG[14][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n652), .Q(\mem_a[14][10] ));
Q_FDP4EP \mem_a_REG[14][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n651), .Q(\mem_a[14][9] ));
Q_FDP4EP \mem_a_REG[14][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n650), .Q(\mem_a[14][8] ));
Q_FDP4EP \mem_a_REG[14][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n649), .Q(\mem_a[14][7] ));
Q_FDP4EP \mem_a_REG[14][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n648), .Q(\mem_a[14][6] ));
Q_FDP4EP \mem_a_REG[14][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n647), .Q(\mem_a[14][5] ));
Q_FDP4EP \mem_a_REG[14][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n646), .Q(\mem_a[14][4] ));
Q_FDP4EP \mem_a_REG[14][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n645), .Q(\mem_a[14][3] ));
Q_FDP4EP \mem_a_REG[14][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n644), .Q(\mem_a[14][2] ));
Q_FDP4EP \mem_a_REG[14][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n643), .Q(\mem_a[14][1] ));
Q_FDP4EP \mem_a_REG[14][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n641), .R(n9), .D(n642), .Q(\mem_a[14][0] ));
Q_FDP4EP \mem_a_REG[13][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n640), .Q(\mem_a[13][31] ));
Q_FDP4EP \mem_a_REG[13][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n639), .Q(\mem_a[13][30] ));
Q_FDP4EP \mem_a_REG[13][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n638), .Q(\mem_a[13][29] ));
Q_FDP4EP \mem_a_REG[13][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n637), .Q(\mem_a[13][28] ));
Q_FDP4EP \mem_a_REG[13][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n636), .Q(\mem_a[13][27] ));
Q_FDP4EP \mem_a_REG[13][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n635), .Q(\mem_a[13][26] ));
Q_FDP4EP \mem_a_REG[13][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n634), .Q(\mem_a[13][25] ));
Q_FDP4EP \mem_a_REG[13][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n633), .Q(\mem_a[13][24] ));
Q_FDP4EP \mem_a_REG[13][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n632), .Q(\mem_a[13][23] ));
Q_FDP4EP \mem_a_REG[13][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n631), .Q(\mem_a[13][22] ));
Q_FDP4EP \mem_a_REG[13][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n630), .Q(\mem_a[13][21] ));
Q_FDP4EP \mem_a_REG[13][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n629), .Q(\mem_a[13][20] ));
Q_FDP4EP \mem_a_REG[13][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n628), .Q(\mem_a[13][19] ));
Q_FDP4EP \mem_a_REG[13][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n627), .Q(\mem_a[13][18] ));
Q_FDP4EP \mem_a_REG[13][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n626), .Q(\mem_a[13][17] ));
Q_FDP4EP \mem_a_REG[13][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n625), .Q(\mem_a[13][16] ));
Q_FDP4EP \mem_a_REG[13][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n624), .Q(\mem_a[13][15] ));
Q_FDP4EP \mem_a_REG[13][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n623), .Q(\mem_a[13][14] ));
Q_FDP4EP \mem_a_REG[13][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n622), .Q(\mem_a[13][13] ));
Q_FDP4EP \mem_a_REG[13][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n621), .Q(\mem_a[13][12] ));
Q_FDP4EP \mem_a_REG[13][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n620), .Q(\mem_a[13][11] ));
Q_FDP4EP \mem_a_REG[13][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n619), .Q(\mem_a[13][10] ));
Q_FDP4EP \mem_a_REG[13][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n618), .Q(\mem_a[13][9] ));
Q_FDP4EP \mem_a_REG[13][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n617), .Q(\mem_a[13][8] ));
Q_FDP4EP \mem_a_REG[13][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n616), .Q(\mem_a[13][7] ));
Q_FDP4EP \mem_a_REG[13][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n615), .Q(\mem_a[13][6] ));
Q_FDP4EP \mem_a_REG[13][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n614), .Q(\mem_a[13][5] ));
Q_FDP4EP \mem_a_REG[13][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n613), .Q(\mem_a[13][4] ));
Q_FDP4EP \mem_a_REG[13][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n612), .Q(\mem_a[13][3] ));
Q_FDP4EP \mem_a_REG[13][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n611), .Q(\mem_a[13][2] ));
Q_FDP4EP \mem_a_REG[13][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n610), .Q(\mem_a[13][1] ));
Q_FDP4EP \mem_a_REG[13][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n608), .R(n9), .D(n609), .Q(\mem_a[13][0] ));
Q_FDP4EP \mem_a_REG[12][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n607), .Q(\mem_a[12][31] ));
Q_FDP4EP \mem_a_REG[12][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n606), .Q(\mem_a[12][30] ));
Q_FDP4EP \mem_a_REG[12][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n605), .Q(\mem_a[12][29] ));
Q_FDP4EP \mem_a_REG[12][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n604), .Q(\mem_a[12][28] ));
Q_FDP4EP \mem_a_REG[12][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n603), .Q(\mem_a[12][27] ));
Q_FDP4EP \mem_a_REG[12][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n602), .Q(\mem_a[12][26] ));
Q_FDP4EP \mem_a_REG[12][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n601), .Q(\mem_a[12][25] ));
Q_FDP4EP \mem_a_REG[12][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n600), .Q(\mem_a[12][24] ));
Q_FDP4EP \mem_a_REG[12][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n599), .Q(\mem_a[12][23] ));
Q_FDP4EP \mem_a_REG[12][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n598), .Q(\mem_a[12][22] ));
Q_FDP4EP \mem_a_REG[12][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n597), .Q(\mem_a[12][21] ));
Q_FDP4EP \mem_a_REG[12][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n596), .Q(\mem_a[12][20] ));
Q_FDP4EP \mem_a_REG[12][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n595), .Q(\mem_a[12][19] ));
Q_FDP4EP \mem_a_REG[12][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n594), .Q(\mem_a[12][18] ));
Q_FDP4EP \mem_a_REG[12][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n593), .Q(\mem_a[12][17] ));
Q_FDP4EP \mem_a_REG[12][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n592), .Q(\mem_a[12][16] ));
Q_FDP4EP \mem_a_REG[12][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n591), .Q(\mem_a[12][15] ));
Q_FDP4EP \mem_a_REG[12][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n590), .Q(\mem_a[12][14] ));
Q_FDP4EP \mem_a_REG[12][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n589), .Q(\mem_a[12][13] ));
Q_FDP4EP \mem_a_REG[12][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n588), .Q(\mem_a[12][12] ));
Q_FDP4EP \mem_a_REG[12][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n587), .Q(\mem_a[12][11] ));
Q_FDP4EP \mem_a_REG[12][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n586), .Q(\mem_a[12][10] ));
Q_FDP4EP \mem_a_REG[12][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n585), .Q(\mem_a[12][9] ));
Q_FDP4EP \mem_a_REG[12][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n584), .Q(\mem_a[12][8] ));
Q_FDP4EP \mem_a_REG[12][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n583), .Q(\mem_a[12][7] ));
Q_FDP4EP \mem_a_REG[12][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n582), .Q(\mem_a[12][6] ));
Q_FDP4EP \mem_a_REG[12][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n581), .Q(\mem_a[12][5] ));
Q_FDP4EP \mem_a_REG[12][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n580), .Q(\mem_a[12][4] ));
Q_FDP4EP \mem_a_REG[12][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n579), .Q(\mem_a[12][3] ));
Q_FDP4EP \mem_a_REG[12][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n578), .Q(\mem_a[12][2] ));
Q_FDP4EP \mem_a_REG[12][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n577), .Q(\mem_a[12][1] ));
Q_FDP4EP \mem_a_REG[12][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n575), .R(n9), .D(n576), .Q(\mem_a[12][0] ));
Q_FDP4EP \mem_a_REG[11][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n574), .Q(\mem_a[11][31] ));
Q_FDP4EP \mem_a_REG[11][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n573), .Q(\mem_a[11][30] ));
Q_FDP4EP \mem_a_REG[11][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n572), .Q(\mem_a[11][29] ));
Q_FDP4EP \mem_a_REG[11][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n571), .Q(\mem_a[11][28] ));
Q_FDP4EP \mem_a_REG[11][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n570), .Q(\mem_a[11][27] ));
Q_FDP4EP \mem_a_REG[11][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n569), .Q(\mem_a[11][26] ));
Q_FDP4EP \mem_a_REG[11][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n568), .Q(\mem_a[11][25] ));
Q_FDP4EP \mem_a_REG[11][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n567), .Q(\mem_a[11][24] ));
Q_FDP4EP \mem_a_REG[11][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n566), .Q(\mem_a[11][23] ));
Q_FDP4EP \mem_a_REG[11][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n565), .Q(\mem_a[11][22] ));
Q_FDP4EP \mem_a_REG[11][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n564), .Q(\mem_a[11][21] ));
Q_FDP4EP \mem_a_REG[11][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n563), .Q(\mem_a[11][20] ));
Q_FDP4EP \mem_a_REG[11][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n562), .Q(\mem_a[11][19] ));
Q_FDP4EP \mem_a_REG[11][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n561), .Q(\mem_a[11][18] ));
Q_FDP4EP \mem_a_REG[11][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n560), .Q(\mem_a[11][17] ));
Q_FDP4EP \mem_a_REG[11][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n559), .Q(\mem_a[11][16] ));
Q_FDP4EP \mem_a_REG[11][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n558), .Q(\mem_a[11][15] ));
Q_FDP4EP \mem_a_REG[11][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n557), .Q(\mem_a[11][14] ));
Q_FDP4EP \mem_a_REG[11][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n556), .Q(\mem_a[11][13] ));
Q_FDP4EP \mem_a_REG[11][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n555), .Q(\mem_a[11][12] ));
Q_FDP4EP \mem_a_REG[11][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n554), .Q(\mem_a[11][11] ));
Q_FDP4EP \mem_a_REG[11][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n553), .Q(\mem_a[11][10] ));
Q_FDP4EP \mem_a_REG[11][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n552), .Q(\mem_a[11][9] ));
Q_FDP4EP \mem_a_REG[11][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n551), .Q(\mem_a[11][8] ));
Q_FDP4EP \mem_a_REG[11][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n550), .Q(\mem_a[11][7] ));
Q_FDP4EP \mem_a_REG[11][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n549), .Q(\mem_a[11][6] ));
Q_FDP4EP \mem_a_REG[11][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n548), .Q(\mem_a[11][5] ));
Q_FDP4EP \mem_a_REG[11][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n547), .Q(\mem_a[11][4] ));
Q_FDP4EP \mem_a_REG[11][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n546), .Q(\mem_a[11][3] ));
Q_FDP4EP \mem_a_REG[11][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n545), .Q(\mem_a[11][2] ));
Q_FDP4EP \mem_a_REG[11][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n544), .Q(\mem_a[11][1] ));
Q_FDP4EP \mem_a_REG[11][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n542), .R(n9), .D(n543), .Q(\mem_a[11][0] ));
Q_FDP4EP \mem_a_REG[10][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n541), .Q(\mem_a[10][31] ));
Q_FDP4EP \mem_a_REG[10][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n540), .Q(\mem_a[10][30] ));
Q_FDP4EP \mem_a_REG[10][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n539), .Q(\mem_a[10][29] ));
Q_FDP4EP \mem_a_REG[10][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n538), .Q(\mem_a[10][28] ));
Q_FDP4EP \mem_a_REG[10][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n537), .Q(\mem_a[10][27] ));
Q_FDP4EP \mem_a_REG[10][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n536), .Q(\mem_a[10][26] ));
Q_FDP4EP \mem_a_REG[10][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n535), .Q(\mem_a[10][25] ));
Q_FDP4EP \mem_a_REG[10][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n534), .Q(\mem_a[10][24] ));
Q_FDP4EP \mem_a_REG[10][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n533), .Q(\mem_a[10][23] ));
Q_FDP4EP \mem_a_REG[10][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n532), .Q(\mem_a[10][22] ));
Q_FDP4EP \mem_a_REG[10][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n531), .Q(\mem_a[10][21] ));
Q_FDP4EP \mem_a_REG[10][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n530), .Q(\mem_a[10][20] ));
Q_FDP4EP \mem_a_REG[10][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n529), .Q(\mem_a[10][19] ));
Q_FDP4EP \mem_a_REG[10][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n528), .Q(\mem_a[10][18] ));
Q_FDP4EP \mem_a_REG[10][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n527), .Q(\mem_a[10][17] ));
Q_FDP4EP \mem_a_REG[10][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n526), .Q(\mem_a[10][16] ));
Q_FDP4EP \mem_a_REG[10][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n525), .Q(\mem_a[10][15] ));
Q_FDP4EP \mem_a_REG[10][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n524), .Q(\mem_a[10][14] ));
Q_FDP4EP \mem_a_REG[10][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n523), .Q(\mem_a[10][13] ));
Q_FDP4EP \mem_a_REG[10][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n522), .Q(\mem_a[10][12] ));
Q_FDP4EP \mem_a_REG[10][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n521), .Q(\mem_a[10][11] ));
Q_FDP4EP \mem_a_REG[10][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n520), .Q(\mem_a[10][10] ));
Q_FDP4EP \mem_a_REG[10][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n519), .Q(\mem_a[10][9] ));
Q_FDP4EP \mem_a_REG[10][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n518), .Q(\mem_a[10][8] ));
Q_FDP4EP \mem_a_REG[10][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n517), .Q(\mem_a[10][7] ));
Q_FDP4EP \mem_a_REG[10][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n516), .Q(\mem_a[10][6] ));
Q_FDP4EP \mem_a_REG[10][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n515), .Q(\mem_a[10][5] ));
Q_FDP4EP \mem_a_REG[10][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n514), .Q(\mem_a[10][4] ));
Q_FDP4EP \mem_a_REG[10][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n513), .Q(\mem_a[10][3] ));
Q_FDP4EP \mem_a_REG[10][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n512), .Q(\mem_a[10][2] ));
Q_FDP4EP \mem_a_REG[10][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n511), .Q(\mem_a[10][1] ));
Q_FDP4EP \mem_a_REG[10][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n509), .R(n9), .D(n510), .Q(\mem_a[10][0] ));
Q_FDP4EP \mem_a_REG[9][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n508), .Q(\mem_a[9][31] ));
Q_FDP4EP \mem_a_REG[9][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n507), .Q(\mem_a[9][30] ));
Q_FDP4EP \mem_a_REG[9][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n506), .Q(\mem_a[9][29] ));
Q_FDP4EP \mem_a_REG[9][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n505), .Q(\mem_a[9][28] ));
Q_FDP4EP \mem_a_REG[9][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n504), .Q(\mem_a[9][27] ));
Q_FDP4EP \mem_a_REG[9][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n503), .Q(\mem_a[9][26] ));
Q_FDP4EP \mem_a_REG[9][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n502), .Q(\mem_a[9][25] ));
Q_FDP4EP \mem_a_REG[9][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n501), .Q(\mem_a[9][24] ));
Q_FDP4EP \mem_a_REG[9][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n500), .Q(\mem_a[9][23] ));
Q_FDP4EP \mem_a_REG[9][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n499), .Q(\mem_a[9][22] ));
Q_FDP4EP \mem_a_REG[9][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n498), .Q(\mem_a[9][21] ));
Q_FDP4EP \mem_a_REG[9][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n497), .Q(\mem_a[9][20] ));
Q_FDP4EP \mem_a_REG[9][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n496), .Q(\mem_a[9][19] ));
Q_FDP4EP \mem_a_REG[9][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n495), .Q(\mem_a[9][18] ));
Q_FDP4EP \mem_a_REG[9][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n494), .Q(\mem_a[9][17] ));
Q_FDP4EP \mem_a_REG[9][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n493), .Q(\mem_a[9][16] ));
Q_FDP4EP \mem_a_REG[9][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n492), .Q(\mem_a[9][15] ));
Q_FDP4EP \mem_a_REG[9][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n491), .Q(\mem_a[9][14] ));
Q_FDP4EP \mem_a_REG[9][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n490), .Q(\mem_a[9][13] ));
Q_FDP4EP \mem_a_REG[9][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n489), .Q(\mem_a[9][12] ));
Q_FDP4EP \mem_a_REG[9][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n488), .Q(\mem_a[9][11] ));
Q_FDP4EP \mem_a_REG[9][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n487), .Q(\mem_a[9][10] ));
Q_FDP4EP \mem_a_REG[9][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n486), .Q(\mem_a[9][9] ));
Q_FDP4EP \mem_a_REG[9][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n485), .Q(\mem_a[9][8] ));
Q_FDP4EP \mem_a_REG[9][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n484), .Q(\mem_a[9][7] ));
Q_FDP4EP \mem_a_REG[9][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n483), .Q(\mem_a[9][6] ));
Q_FDP4EP \mem_a_REG[9][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n482), .Q(\mem_a[9][5] ));
Q_FDP4EP \mem_a_REG[9][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n481), .Q(\mem_a[9][4] ));
Q_FDP4EP \mem_a_REG[9][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n480), .Q(\mem_a[9][3] ));
Q_FDP4EP \mem_a_REG[9][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n479), .Q(\mem_a[9][2] ));
Q_FDP4EP \mem_a_REG[9][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n478), .Q(\mem_a[9][1] ));
Q_FDP4EP \mem_a_REG[9][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n476), .R(n9), .D(n477), .Q(\mem_a[9][0] ));
Q_FDP4EP \mem_a_REG[8][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n475), .Q(\mem_a[8][31] ));
Q_FDP4EP \mem_a_REG[8][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n474), .Q(\mem_a[8][30] ));
Q_FDP4EP \mem_a_REG[8][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n473), .Q(\mem_a[8][29] ));
Q_FDP4EP \mem_a_REG[8][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n472), .Q(\mem_a[8][28] ));
Q_FDP4EP \mem_a_REG[8][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n471), .Q(\mem_a[8][27] ));
Q_FDP4EP \mem_a_REG[8][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n470), .Q(\mem_a[8][26] ));
Q_FDP4EP \mem_a_REG[8][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n469), .Q(\mem_a[8][25] ));
Q_FDP4EP \mem_a_REG[8][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n468), .Q(\mem_a[8][24] ));
Q_FDP4EP \mem_a_REG[8][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n467), .Q(\mem_a[8][23] ));
Q_FDP4EP \mem_a_REG[8][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n466), .Q(\mem_a[8][22] ));
Q_FDP4EP \mem_a_REG[8][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n465), .Q(\mem_a[8][21] ));
Q_FDP4EP \mem_a_REG[8][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n464), .Q(\mem_a[8][20] ));
Q_FDP4EP \mem_a_REG[8][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n463), .Q(\mem_a[8][19] ));
Q_FDP4EP \mem_a_REG[8][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n462), .Q(\mem_a[8][18] ));
Q_FDP4EP \mem_a_REG[8][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n461), .Q(\mem_a[8][17] ));
Q_FDP4EP \mem_a_REG[8][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n460), .Q(\mem_a[8][16] ));
Q_FDP4EP \mem_a_REG[8][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n459), .Q(\mem_a[8][15] ));
Q_FDP4EP \mem_a_REG[8][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n458), .Q(\mem_a[8][14] ));
Q_FDP4EP \mem_a_REG[8][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n457), .Q(\mem_a[8][13] ));
Q_FDP4EP \mem_a_REG[8][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n456), .Q(\mem_a[8][12] ));
Q_FDP4EP \mem_a_REG[8][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n455), .Q(\mem_a[8][11] ));
Q_FDP4EP \mem_a_REG[8][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n454), .Q(\mem_a[8][10] ));
Q_FDP4EP \mem_a_REG[8][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n453), .Q(\mem_a[8][9] ));
Q_FDP4EP \mem_a_REG[8][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n452), .Q(\mem_a[8][8] ));
Q_FDP4EP \mem_a_REG[8][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n451), .Q(\mem_a[8][7] ));
Q_FDP4EP \mem_a_REG[8][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n450), .Q(\mem_a[8][6] ));
Q_FDP4EP \mem_a_REG[8][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n449), .Q(\mem_a[8][5] ));
Q_FDP4EP \mem_a_REG[8][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n448), .Q(\mem_a[8][4] ));
Q_FDP4EP \mem_a_REG[8][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n447), .Q(\mem_a[8][3] ));
Q_FDP4EP \mem_a_REG[8][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n446), .Q(\mem_a[8][2] ));
Q_FDP4EP \mem_a_REG[8][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n445), .Q(\mem_a[8][1] ));
Q_FDP4EP \mem_a_REG[8][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n443), .R(n9), .D(n444), .Q(\mem_a[8][0] ));
Q_FDP4EP \mem_a_REG[7][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n442), .Q(\mem_a[7][31] ));
Q_FDP4EP \mem_a_REG[7][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n441), .Q(\mem_a[7][30] ));
Q_FDP4EP \mem_a_REG[7][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n440), .Q(\mem_a[7][29] ));
Q_FDP4EP \mem_a_REG[7][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n439), .Q(\mem_a[7][28] ));
Q_FDP4EP \mem_a_REG[7][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n438), .Q(\mem_a[7][27] ));
Q_FDP4EP \mem_a_REG[7][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n437), .Q(\mem_a[7][26] ));
Q_FDP4EP \mem_a_REG[7][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n436), .Q(\mem_a[7][25] ));
Q_FDP4EP \mem_a_REG[7][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n435), .Q(\mem_a[7][24] ));
Q_FDP4EP \mem_a_REG[7][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n434), .Q(\mem_a[7][23] ));
Q_FDP4EP \mem_a_REG[7][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n433), .Q(\mem_a[7][22] ));
Q_FDP4EP \mem_a_REG[7][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n432), .Q(\mem_a[7][21] ));
Q_FDP4EP \mem_a_REG[7][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n431), .Q(\mem_a[7][20] ));
Q_FDP4EP \mem_a_REG[7][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n430), .Q(\mem_a[7][19] ));
Q_FDP4EP \mem_a_REG[7][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n429), .Q(\mem_a[7][18] ));
Q_FDP4EP \mem_a_REG[7][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n428), .Q(\mem_a[7][17] ));
Q_FDP4EP \mem_a_REG[7][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n427), .Q(\mem_a[7][16] ));
Q_FDP4EP \mem_a_REG[7][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n426), .Q(\mem_a[7][15] ));
Q_FDP4EP \mem_a_REG[7][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n425), .Q(\mem_a[7][14] ));
Q_FDP4EP \mem_a_REG[7][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n424), .Q(\mem_a[7][13] ));
Q_FDP4EP \mem_a_REG[7][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n423), .Q(\mem_a[7][12] ));
Q_FDP4EP \mem_a_REG[7][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n422), .Q(\mem_a[7][11] ));
Q_FDP4EP \mem_a_REG[7][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n421), .Q(\mem_a[7][10] ));
Q_FDP4EP \mem_a_REG[7][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n420), .Q(\mem_a[7][9] ));
Q_FDP4EP \mem_a_REG[7][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n419), .Q(\mem_a[7][8] ));
Q_FDP4EP \mem_a_REG[7][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n418), .Q(\mem_a[7][7] ));
Q_FDP4EP \mem_a_REG[7][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n417), .Q(\mem_a[7][6] ));
Q_FDP4EP \mem_a_REG[7][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n416), .Q(\mem_a[7][5] ));
Q_FDP4EP \mem_a_REG[7][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n415), .Q(\mem_a[7][4] ));
Q_FDP4EP \mem_a_REG[7][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n414), .Q(\mem_a[7][3] ));
Q_FDP4EP \mem_a_REG[7][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n413), .Q(\mem_a[7][2] ));
Q_FDP4EP \mem_a_REG[7][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n412), .Q(\mem_a[7][1] ));
Q_FDP4EP \mem_a_REG[7][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n410), .R(n9), .D(n411), .Q(\mem_a[7][0] ));
Q_FDP4EP \mem_a_REG[6][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n409), .Q(\mem_a[6][31] ));
Q_FDP4EP \mem_a_REG[6][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n408), .Q(\mem_a[6][30] ));
Q_FDP4EP \mem_a_REG[6][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n407), .Q(\mem_a[6][29] ));
Q_FDP4EP \mem_a_REG[6][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n406), .Q(\mem_a[6][28] ));
Q_FDP4EP \mem_a_REG[6][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n405), .Q(\mem_a[6][27] ));
Q_FDP4EP \mem_a_REG[6][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n404), .Q(\mem_a[6][26] ));
Q_FDP4EP \mem_a_REG[6][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n403), .Q(\mem_a[6][25] ));
Q_FDP4EP \mem_a_REG[6][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n402), .Q(\mem_a[6][24] ));
Q_FDP4EP \mem_a_REG[6][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n401), .Q(\mem_a[6][23] ));
Q_FDP4EP \mem_a_REG[6][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n400), .Q(\mem_a[6][22] ));
Q_FDP4EP \mem_a_REG[6][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n399), .Q(\mem_a[6][21] ));
Q_FDP4EP \mem_a_REG[6][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n398), .Q(\mem_a[6][20] ));
Q_FDP4EP \mem_a_REG[6][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n397), .Q(\mem_a[6][19] ));
Q_FDP4EP \mem_a_REG[6][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n396), .Q(\mem_a[6][18] ));
Q_FDP4EP \mem_a_REG[6][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n395), .Q(\mem_a[6][17] ));
Q_FDP4EP \mem_a_REG[6][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n394), .Q(\mem_a[6][16] ));
Q_FDP4EP \mem_a_REG[6][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n393), .Q(\mem_a[6][15] ));
Q_FDP4EP \mem_a_REG[6][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n392), .Q(\mem_a[6][14] ));
Q_FDP4EP \mem_a_REG[6][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n391), .Q(\mem_a[6][13] ));
Q_FDP4EP \mem_a_REG[6][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n390), .Q(\mem_a[6][12] ));
Q_FDP4EP \mem_a_REG[6][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n389), .Q(\mem_a[6][11] ));
Q_FDP4EP \mem_a_REG[6][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n388), .Q(\mem_a[6][10] ));
Q_FDP4EP \mem_a_REG[6][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n387), .Q(\mem_a[6][9] ));
Q_FDP4EP \mem_a_REG[6][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n386), .Q(\mem_a[6][8] ));
Q_FDP4EP \mem_a_REG[6][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n385), .Q(\mem_a[6][7] ));
Q_FDP4EP \mem_a_REG[6][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n384), .Q(\mem_a[6][6] ));
Q_FDP4EP \mem_a_REG[6][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n383), .Q(\mem_a[6][5] ));
Q_FDP4EP \mem_a_REG[6][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n382), .Q(\mem_a[6][4] ));
Q_FDP4EP \mem_a_REG[6][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n381), .Q(\mem_a[6][3] ));
Q_FDP4EP \mem_a_REG[6][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n380), .Q(\mem_a[6][2] ));
Q_FDP4EP \mem_a_REG[6][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n379), .Q(\mem_a[6][1] ));
Q_FDP4EP \mem_a_REG[6][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n377), .R(n9), .D(n378), .Q(\mem_a[6][0] ));
Q_FDP4EP \mem_a_REG[5][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n376), .Q(\mem_a[5][31] ));
Q_FDP4EP \mem_a_REG[5][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n375), .Q(\mem_a[5][30] ));
Q_FDP4EP \mem_a_REG[5][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n374), .Q(\mem_a[5][29] ));
Q_FDP4EP \mem_a_REG[5][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n373), .Q(\mem_a[5][28] ));
Q_FDP4EP \mem_a_REG[5][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n372), .Q(\mem_a[5][27] ));
Q_FDP4EP \mem_a_REG[5][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n371), .Q(\mem_a[5][26] ));
Q_FDP4EP \mem_a_REG[5][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n370), .Q(\mem_a[5][25] ));
Q_FDP4EP \mem_a_REG[5][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n369), .Q(\mem_a[5][24] ));
Q_FDP4EP \mem_a_REG[5][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n368), .Q(\mem_a[5][23] ));
Q_FDP4EP \mem_a_REG[5][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n367), .Q(\mem_a[5][22] ));
Q_FDP4EP \mem_a_REG[5][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n366), .Q(\mem_a[5][21] ));
Q_FDP4EP \mem_a_REG[5][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n365), .Q(\mem_a[5][20] ));
Q_FDP4EP \mem_a_REG[5][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n364), .Q(\mem_a[5][19] ));
Q_FDP4EP \mem_a_REG[5][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n363), .Q(\mem_a[5][18] ));
Q_FDP4EP \mem_a_REG[5][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n362), .Q(\mem_a[5][17] ));
Q_FDP4EP \mem_a_REG[5][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n361), .Q(\mem_a[5][16] ));
Q_FDP4EP \mem_a_REG[5][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n360), .Q(\mem_a[5][15] ));
Q_FDP4EP \mem_a_REG[5][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n359), .Q(\mem_a[5][14] ));
Q_FDP4EP \mem_a_REG[5][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n358), .Q(\mem_a[5][13] ));
Q_FDP4EP \mem_a_REG[5][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n357), .Q(\mem_a[5][12] ));
Q_FDP4EP \mem_a_REG[5][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n356), .Q(\mem_a[5][11] ));
Q_FDP4EP \mem_a_REG[5][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n355), .Q(\mem_a[5][10] ));
Q_FDP4EP \mem_a_REG[5][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n354), .Q(\mem_a[5][9] ));
Q_FDP4EP \mem_a_REG[5][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n353), .Q(\mem_a[5][8] ));
Q_FDP4EP \mem_a_REG[5][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n352), .Q(\mem_a[5][7] ));
Q_FDP4EP \mem_a_REG[5][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n351), .Q(\mem_a[5][6] ));
Q_FDP4EP \mem_a_REG[5][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n350), .Q(\mem_a[5][5] ));
Q_FDP4EP \mem_a_REG[5][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n349), .Q(\mem_a[5][4] ));
Q_FDP4EP \mem_a_REG[5][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n348), .Q(\mem_a[5][3] ));
Q_FDP4EP \mem_a_REG[5][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n347), .Q(\mem_a[5][2] ));
Q_FDP4EP \mem_a_REG[5][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n346), .Q(\mem_a[5][1] ));
Q_FDP4EP \mem_a_REG[5][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n344), .R(n9), .D(n345), .Q(\mem_a[5][0] ));
Q_FDP4EP \mem_a_REG[4][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n343), .Q(\mem_a[4][31] ));
Q_FDP4EP \mem_a_REG[4][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n342), .Q(\mem_a[4][30] ));
Q_FDP4EP \mem_a_REG[4][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n341), .Q(\mem_a[4][29] ));
Q_FDP4EP \mem_a_REG[4][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n340), .Q(\mem_a[4][28] ));
Q_FDP4EP \mem_a_REG[4][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n339), .Q(\mem_a[4][27] ));
Q_FDP4EP \mem_a_REG[4][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n338), .Q(\mem_a[4][26] ));
Q_FDP4EP \mem_a_REG[4][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n337), .Q(\mem_a[4][25] ));
Q_FDP4EP \mem_a_REG[4][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n336), .Q(\mem_a[4][24] ));
Q_FDP4EP \mem_a_REG[4][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n335), .Q(\mem_a[4][23] ));
Q_FDP4EP \mem_a_REG[4][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n334), .Q(\mem_a[4][22] ));
Q_FDP4EP \mem_a_REG[4][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n333), .Q(\mem_a[4][21] ));
Q_FDP4EP \mem_a_REG[4][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n332), .Q(\mem_a[4][20] ));
Q_FDP4EP \mem_a_REG[4][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n331), .Q(\mem_a[4][19] ));
Q_FDP4EP \mem_a_REG[4][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n330), .Q(\mem_a[4][18] ));
Q_FDP4EP \mem_a_REG[4][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n329), .Q(\mem_a[4][17] ));
Q_FDP4EP \mem_a_REG[4][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n328), .Q(\mem_a[4][16] ));
Q_FDP4EP \mem_a_REG[4][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n327), .Q(\mem_a[4][15] ));
Q_FDP4EP \mem_a_REG[4][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n326), .Q(\mem_a[4][14] ));
Q_FDP4EP \mem_a_REG[4][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n325), .Q(\mem_a[4][13] ));
Q_FDP4EP \mem_a_REG[4][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n324), .Q(\mem_a[4][12] ));
Q_FDP4EP \mem_a_REG[4][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n323), .Q(\mem_a[4][11] ));
Q_FDP4EP \mem_a_REG[4][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n322), .Q(\mem_a[4][10] ));
Q_FDP4EP \mem_a_REG[4][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n321), .Q(\mem_a[4][9] ));
Q_FDP4EP \mem_a_REG[4][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n320), .Q(\mem_a[4][8] ));
Q_FDP4EP \mem_a_REG[4][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n319), .Q(\mem_a[4][7] ));
Q_FDP4EP \mem_a_REG[4][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n318), .Q(\mem_a[4][6] ));
Q_FDP4EP \mem_a_REG[4][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n317), .Q(\mem_a[4][5] ));
Q_FDP4EP \mem_a_REG[4][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n316), .Q(\mem_a[4][4] ));
Q_FDP4EP \mem_a_REG[4][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n315), .Q(\mem_a[4][3] ));
Q_FDP4EP \mem_a_REG[4][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n314), .Q(\mem_a[4][2] ));
Q_FDP4EP \mem_a_REG[4][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n313), .Q(\mem_a[4][1] ));
Q_FDP4EP \mem_a_REG[4][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n311), .R(n9), .D(n312), .Q(\mem_a[4][0] ));
Q_FDP4EP \mem_a_REG[3][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n310), .Q(\mem_a[3][31] ));
Q_FDP4EP \mem_a_REG[3][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n309), .Q(\mem_a[3][30] ));
Q_FDP4EP \mem_a_REG[3][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n308), .Q(\mem_a[3][29] ));
Q_FDP4EP \mem_a_REG[3][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n307), .Q(\mem_a[3][28] ));
Q_FDP4EP \mem_a_REG[3][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n306), .Q(\mem_a[3][27] ));
Q_FDP4EP \mem_a_REG[3][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n305), .Q(\mem_a[3][26] ));
Q_FDP4EP \mem_a_REG[3][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n304), .Q(\mem_a[3][25] ));
Q_FDP4EP \mem_a_REG[3][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n303), .Q(\mem_a[3][24] ));
Q_FDP4EP \mem_a_REG[3][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n302), .Q(\mem_a[3][23] ));
Q_FDP4EP \mem_a_REG[3][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n301), .Q(\mem_a[3][22] ));
Q_FDP4EP \mem_a_REG[3][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n300), .Q(\mem_a[3][21] ));
Q_FDP4EP \mem_a_REG[3][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n299), .Q(\mem_a[3][20] ));
Q_FDP4EP \mem_a_REG[3][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n298), .Q(\mem_a[3][19] ));
Q_FDP4EP \mem_a_REG[3][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n297), .Q(\mem_a[3][18] ));
Q_FDP4EP \mem_a_REG[3][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n296), .Q(\mem_a[3][17] ));
Q_FDP4EP \mem_a_REG[3][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n295), .Q(\mem_a[3][16] ));
Q_FDP4EP \mem_a_REG[3][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n294), .Q(\mem_a[3][15] ));
Q_FDP4EP \mem_a_REG[3][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n293), .Q(\mem_a[3][14] ));
Q_FDP4EP \mem_a_REG[3][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n292), .Q(\mem_a[3][13] ));
Q_FDP4EP \mem_a_REG[3][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n291), .Q(\mem_a[3][12] ));
Q_FDP4EP \mem_a_REG[3][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n290), .Q(\mem_a[3][11] ));
Q_FDP4EP \mem_a_REG[3][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n289), .Q(\mem_a[3][10] ));
Q_FDP4EP \mem_a_REG[3][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n288), .Q(\mem_a[3][9] ));
Q_FDP4EP \mem_a_REG[3][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n287), .Q(\mem_a[3][8] ));
Q_FDP4EP \mem_a_REG[3][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n286), .Q(\mem_a[3][7] ));
Q_FDP4EP \mem_a_REG[3][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n285), .Q(\mem_a[3][6] ));
Q_FDP4EP \mem_a_REG[3][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n284), .Q(\mem_a[3][5] ));
Q_FDP4EP \mem_a_REG[3][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n283), .Q(\mem_a[3][4] ));
Q_FDP4EP \mem_a_REG[3][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n282), .Q(\mem_a[3][3] ));
Q_FDP4EP \mem_a_REG[3][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n281), .Q(\mem_a[3][2] ));
Q_FDP4EP \mem_a_REG[3][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n280), .Q(\mem_a[3][1] ));
Q_FDP4EP \mem_a_REG[3][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n278), .R(n9), .D(n279), .Q(\mem_a[3][0] ));
Q_FDP4EP \mem_a_REG[2][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n277), .Q(\mem_a[2][31] ));
Q_FDP4EP \mem_a_REG[2][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n276), .Q(\mem_a[2][30] ));
Q_FDP4EP \mem_a_REG[2][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n275), .Q(\mem_a[2][29] ));
Q_FDP4EP \mem_a_REG[2][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n274), .Q(\mem_a[2][28] ));
Q_FDP4EP \mem_a_REG[2][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n273), .Q(\mem_a[2][27] ));
Q_FDP4EP \mem_a_REG[2][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n272), .Q(\mem_a[2][26] ));
Q_FDP4EP \mem_a_REG[2][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n271), .Q(\mem_a[2][25] ));
Q_FDP4EP \mem_a_REG[2][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n270), .Q(\mem_a[2][24] ));
Q_FDP4EP \mem_a_REG[2][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n269), .Q(\mem_a[2][23] ));
Q_FDP4EP \mem_a_REG[2][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n268), .Q(\mem_a[2][22] ));
Q_FDP4EP \mem_a_REG[2][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n267), .Q(\mem_a[2][21] ));
Q_FDP4EP \mem_a_REG[2][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n266), .Q(\mem_a[2][20] ));
Q_FDP4EP \mem_a_REG[2][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n265), .Q(\mem_a[2][19] ));
Q_FDP4EP \mem_a_REG[2][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n264), .Q(\mem_a[2][18] ));
Q_FDP4EP \mem_a_REG[2][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n263), .Q(\mem_a[2][17] ));
Q_FDP4EP \mem_a_REG[2][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n262), .Q(\mem_a[2][16] ));
Q_FDP4EP \mem_a_REG[2][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n261), .Q(\mem_a[2][15] ));
Q_FDP4EP \mem_a_REG[2][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n260), .Q(\mem_a[2][14] ));
Q_FDP4EP \mem_a_REG[2][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n259), .Q(\mem_a[2][13] ));
Q_FDP4EP \mem_a_REG[2][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n258), .Q(\mem_a[2][12] ));
Q_FDP4EP \mem_a_REG[2][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n257), .Q(\mem_a[2][11] ));
Q_FDP4EP \mem_a_REG[2][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n256), .Q(\mem_a[2][10] ));
Q_FDP4EP \mem_a_REG[2][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n255), .Q(\mem_a[2][9] ));
Q_FDP4EP \mem_a_REG[2][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n254), .Q(\mem_a[2][8] ));
Q_FDP4EP \mem_a_REG[2][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n253), .Q(\mem_a[2][7] ));
Q_FDP4EP \mem_a_REG[2][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n252), .Q(\mem_a[2][6] ));
Q_FDP4EP \mem_a_REG[2][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n251), .Q(\mem_a[2][5] ));
Q_FDP4EP \mem_a_REG[2][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n250), .Q(\mem_a[2][4] ));
Q_FDP4EP \mem_a_REG[2][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n249), .Q(\mem_a[2][3] ));
Q_FDP4EP \mem_a_REG[2][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n248), .Q(\mem_a[2][2] ));
Q_FDP4EP \mem_a_REG[2][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n247), .Q(\mem_a[2][1] ));
Q_FDP4EP \mem_a_REG[2][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n245), .R(n9), .D(n246), .Q(\mem_a[2][0] ));
Q_FDP4EP \mem_a_REG[1][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n244), .Q(\mem_a[1][31] ));
Q_FDP4EP \mem_a_REG[1][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n243), .Q(\mem_a[1][30] ));
Q_FDP4EP \mem_a_REG[1][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n242), .Q(\mem_a[1][29] ));
Q_FDP4EP \mem_a_REG[1][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n241), .Q(\mem_a[1][28] ));
Q_FDP4EP \mem_a_REG[1][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n240), .Q(\mem_a[1][27] ));
Q_FDP4EP \mem_a_REG[1][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n239), .Q(\mem_a[1][26] ));
Q_FDP4EP \mem_a_REG[1][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n238), .Q(\mem_a[1][25] ));
Q_FDP4EP \mem_a_REG[1][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n237), .Q(\mem_a[1][24] ));
Q_FDP4EP \mem_a_REG[1][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n236), .Q(\mem_a[1][23] ));
Q_FDP4EP \mem_a_REG[1][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n235), .Q(\mem_a[1][22] ));
Q_FDP4EP \mem_a_REG[1][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n234), .Q(\mem_a[1][21] ));
Q_FDP4EP \mem_a_REG[1][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n233), .Q(\mem_a[1][20] ));
Q_FDP4EP \mem_a_REG[1][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n232), .Q(\mem_a[1][19] ));
Q_FDP4EP \mem_a_REG[1][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n231), .Q(\mem_a[1][18] ));
Q_FDP4EP \mem_a_REG[1][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n230), .Q(\mem_a[1][17] ));
Q_FDP4EP \mem_a_REG[1][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n229), .Q(\mem_a[1][16] ));
Q_FDP4EP \mem_a_REG[1][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n228), .Q(\mem_a[1][15] ));
Q_FDP4EP \mem_a_REG[1][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n227), .Q(\mem_a[1][14] ));
Q_FDP4EP \mem_a_REG[1][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n226), .Q(\mem_a[1][13] ));
Q_FDP4EP \mem_a_REG[1][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n225), .Q(\mem_a[1][12] ));
Q_FDP4EP \mem_a_REG[1][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n224), .Q(\mem_a[1][11] ));
Q_FDP4EP \mem_a_REG[1][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n223), .Q(\mem_a[1][10] ));
Q_FDP4EP \mem_a_REG[1][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n222), .Q(\mem_a[1][9] ));
Q_FDP4EP \mem_a_REG[1][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n221), .Q(\mem_a[1][8] ));
Q_FDP4EP \mem_a_REG[1][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n220), .Q(\mem_a[1][7] ));
Q_FDP4EP \mem_a_REG[1][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n219), .Q(\mem_a[1][6] ));
Q_FDP4EP \mem_a_REG[1][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n218), .Q(\mem_a[1][5] ));
Q_FDP4EP \mem_a_REG[1][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n217), .Q(\mem_a[1][4] ));
Q_FDP4EP \mem_a_REG[1][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n216), .Q(\mem_a[1][3] ));
Q_FDP4EP \mem_a_REG[1][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n215), .Q(\mem_a[1][2] ));
Q_FDP4EP \mem_a_REG[1][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n214), .Q(\mem_a[1][1] ));
Q_FDP4EP \mem_a_REG[1][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n212), .R(n9), .D(n213), .Q(\mem_a[1][0] ));
Q_FDP4EP \mem_a_REG[0][31] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n41), .Q(\mem_a[0][31] ));
Q_FDP4EP \mem_a_REG[0][30] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n40), .Q(\mem_a[0][30] ));
Q_FDP4EP \mem_a_REG[0][29] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n39), .Q(\mem_a[0][29] ));
Q_FDP4EP \mem_a_REG[0][28] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n38), .Q(\mem_a[0][28] ));
Q_FDP4EP \mem_a_REG[0][27] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n37), .Q(\mem_a[0][27] ));
Q_FDP4EP \mem_a_REG[0][26] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n36), .Q(\mem_a[0][26] ));
Q_FDP4EP \mem_a_REG[0][25] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n35), .Q(\mem_a[0][25] ));
Q_FDP4EP \mem_a_REG[0][24] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n34), .Q(\mem_a[0][24] ));
Q_FDP4EP \mem_a_REG[0][23] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n33), .Q(\mem_a[0][23] ));
Q_FDP4EP \mem_a_REG[0][22] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n32), .Q(\mem_a[0][22] ));
Q_FDP4EP \mem_a_REG[0][21] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n31), .Q(\mem_a[0][21] ));
Q_FDP4EP \mem_a_REG[0][20] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n30), .Q(\mem_a[0][20] ));
Q_FDP4EP \mem_a_REG[0][19] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n29), .Q(\mem_a[0][19] ));
Q_FDP4EP \mem_a_REG[0][18] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n28), .Q(\mem_a[0][18] ));
Q_FDP4EP \mem_a_REG[0][17] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n27), .Q(\mem_a[0][17] ));
Q_FDP4EP \mem_a_REG[0][16] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n26), .Q(\mem_a[0][16] ));
Q_FDP4EP \mem_a_REG[0][15] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n25), .Q(\mem_a[0][15] ));
Q_FDP4EP \mem_a_REG[0][14] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n24), .Q(\mem_a[0][14] ));
Q_FDP4EP \mem_a_REG[0][13] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n23), .Q(\mem_a[0][13] ));
Q_FDP4EP \mem_a_REG[0][12] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n22), .Q(\mem_a[0][12] ));
Q_FDP4EP \mem_a_REG[0][11] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n21), .Q(\mem_a[0][11] ));
Q_FDP4EP \mem_a_REG[0][10] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n20), .Q(\mem_a[0][10] ));
Q_FDP4EP \mem_a_REG[0][9] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n19), .Q(\mem_a[0][9] ));
Q_FDP4EP \mem_a_REG[0][8] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n18), .Q(\mem_a[0][8] ));
Q_FDP4EP \mem_a_REG[0][7] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n17), .Q(\mem_a[0][7] ));
Q_FDP4EP \mem_a_REG[0][6] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n16), .Q(\mem_a[0][6] ));
Q_FDP4EP \mem_a_REG[0][5] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n15), .Q(\mem_a[0][5] ));
Q_FDP4EP \mem_a_REG[0][4] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n14), .Q(\mem_a[0][4] ));
Q_FDP4EP \mem_a_REG[0][3] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n13), .Q(\mem_a[0][3] ));
Q_FDP4EP \mem_a_REG[0][2] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n12), .Q(\mem_a[0][2] ));
Q_FDP4EP \mem_a_REG[0][1] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n11), .Q(\mem_a[0][1] ));
Q_FDP4EP \mem_a_REG[0][0] ( .CK(_zzM132L132_bcMevClk0), .CE(n211), .R(n9), .D(n10), .Q(\mem_a[0][0] ));
Q_INV U2392 ( .A(_zzM132_bcBehEval[0]), .Z(n1363));
Q_FDP4EP \_zzM132_bcBehEval_REG[0] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n1363), .Q(_zzM132_bcBehEval[0]));
Q_FDP4EP \_zzM132_bcBehEval_REG[1] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n126), .Q(_zzM132_bcBehEval[1]));
Q_FDP4EP \_zzM132_bcBehEval_REG[2] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n128), .Q(_zzM132_bcBehEval[2]));
Q_FDP4EP \_zzM132_bcBehEval_REG[3] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n130), .Q(_zzM132_bcBehEval[3]));
Q_FDP4EP \_zzM132_bcBehEval_REG[4] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n132), .Q(_zzM132_bcBehEval[4]));
Q_FDP4EP \_zzM132_bcBehEval_REG[5] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n134), .Q(_zzM132_bcBehEval[5]));
Q_FDP4EP \_zzM132_bcBehEval_REG[6] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n136), .Q(_zzM132_bcBehEval[6]));
Q_FDP4EP \_zzM132_bcBehEval_REG[7] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n138), .Q(_zzM132_bcBehEval[7]));
Q_FDP4EP \_zzM132_bcBehEval_REG[8] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n140), .Q(_zzM132_bcBehEval[8]));
Q_FDP4EP \_zzM132_bcBehEval_REG[9] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n142), .Q(_zzM132_bcBehEval[9]));
Q_FDP4EP \_zzM132_bcBehEval_REG[10] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n144), .Q(_zzM132_bcBehEval[10]));
Q_FDP4EP \_zzM132_bcBehEval_REG[11] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n146), .Q(_zzM132_bcBehEval[11]));
Q_FDP4EP \_zzM132_bcBehEval_REG[12] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n148), .Q(_zzM132_bcBehEval[12]));
Q_FDP4EP \_zzM132_bcBehEval_REG[13] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n150), .Q(_zzM132_bcBehEval[13]));
Q_FDP4EP \_zzM132_bcBehEval_REG[14] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n152), .Q(_zzM132_bcBehEval[14]));
Q_FDP4EP \_zzM132_bcBehEval_REG[15] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n154), .Q(_zzM132_bcBehEval[15]));
Q_FDP4EP \_zzM132_bcBehEval_REG[16] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n156), .Q(_zzM132_bcBehEval[16]));
Q_FDP4EP \_zzM132_bcBehEval_REG[17] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n158), .Q(_zzM132_bcBehEval[17]));
Q_FDP4EP \_zzM132_bcBehEval_REG[18] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n160), .Q(_zzM132_bcBehEval[18]));
Q_FDP4EP \_zzM132_bcBehEval_REG[19] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n162), .Q(_zzM132_bcBehEval[19]));
Q_FDP4EP \_zzM132_bcBehEval_REG[20] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n164), .Q(_zzM132_bcBehEval[20]));
Q_FDP4EP \_zzM132_bcBehEval_REG[21] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n166), .Q(_zzM132_bcBehEval[21]));
Q_FDP4EP \_zzM132_bcBehEval_REG[22] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n168), .Q(_zzM132_bcBehEval[22]));
Q_FDP4EP \_zzM132_bcBehEval_REG[23] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n170), .Q(_zzM132_bcBehEval[23]));
Q_FDP4EP \_zzM132_bcBehEval_REG[24] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n172), .Q(_zzM132_bcBehEval[24]));
Q_FDP4EP \_zzM132_bcBehEval_REG[25] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n174), .Q(_zzM132_bcBehEval[25]));
Q_FDP4EP \_zzM132_bcBehEval_REG[26] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n176), .Q(_zzM132_bcBehEval[26]));
Q_FDP4EP \_zzM132_bcBehEval_REG[27] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n178), .Q(_zzM132_bcBehEval[27]));
Q_FDP4EP \_zzM132_bcBehEval_REG[28] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n180), .Q(_zzM132_bcBehEval[28]));
Q_FDP4EP \_zzM132_bcBehEval_REG[29] ( .CK(_zzM132_bcBehEvalClk), .CE(n184), .R(n9), .D(n182), .Q(_zzM132_bcBehEval[29]));
Q_INV U2423 ( .A(_zzM132_bcBehEval[30]), .Z(n1364));
Q_FDP4EP \_zzM132_bcBehEval_REG[30] ( .CK(_zzM132_bcBehEvalClk), .CE(n3), .R(n9), .D(n1364), .Q(_zzM132_bcBehEval[30]));
Q_FDP4EP \_zzM132_bcBehEval_REG[31] ( .CK(_zzM132_bcBehEvalClk), .CE(_zzM132L132_bcWait0), .R(n9), .D(_zzM132_bcBehHalt), .Q(_zzM132_bcBehEval[31]));
Q_FDP4EP \sw_rdat_REG[0] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n47), .Q(sw_rdat[0]));
Q_INV U2427 ( .A(rst_n), .Z(n1365));
Q_FDP4EP \sw_rdat_REG[1] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n48), .Q(sw_rdat[1]));
Q_FDP4EP \sw_rdat_REG[2] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n49), .Q(sw_rdat[2]));
Q_FDP4EP \sw_rdat_REG[3] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n50), .Q(sw_rdat[3]));
Q_FDP4EP \sw_rdat_REG[4] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n51), .Q(sw_rdat[4]));
Q_FDP4EP \sw_rdat_REG[5] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n52), .Q(sw_rdat[5]));
Q_FDP4EP \sw_rdat_REG[6] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n53), .Q(sw_rdat[6]));
Q_FDP4EP \sw_rdat_REG[7] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n54), .Q(sw_rdat[7]));
Q_FDP4EP \sw_rdat_REG[8] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n55), .Q(sw_rdat[8]));
Q_FDP4EP \sw_rdat_REG[9] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n56), .Q(sw_rdat[9]));
Q_FDP4EP \sw_rdat_REG[10] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n57), .Q(sw_rdat[10]));
Q_FDP4EP \sw_rdat_REG[11] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n58), .Q(sw_rdat[11]));
Q_FDP4EP \sw_rdat_REG[12] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n59), .Q(sw_rdat[12]));
Q_FDP4EP \sw_rdat_REG[13] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n60), .Q(sw_rdat[13]));
Q_FDP4EP \sw_rdat_REG[14] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n61), .Q(sw_rdat[14]));
Q_FDP4EP \sw_rdat_REG[15] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n62), .Q(sw_rdat[15]));
Q_FDP4EP \sw_rdat_REG[16] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n63), .Q(sw_rdat[16]));
Q_FDP4EP \sw_rdat_REG[17] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n64), .Q(sw_rdat[17]));
Q_FDP4EP \sw_rdat_REG[18] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n65), .Q(sw_rdat[18]));
Q_FDP4EP \sw_rdat_REG[19] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n66), .Q(sw_rdat[19]));
Q_FDP4EP \sw_rdat_REG[20] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n67), .Q(sw_rdat[20]));
Q_FDP4EP \sw_rdat_REG[21] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n68), .Q(sw_rdat[21]));
Q_FDP4EP \sw_rdat_REG[22] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n69), .Q(sw_rdat[22]));
Q_FDP4EP \sw_rdat_REG[23] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n70), .Q(sw_rdat[23]));
Q_FDP4EP \sw_rdat_REG[24] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n71), .Q(sw_rdat[24]));
Q_FDP4EP \sw_rdat_REG[25] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n72), .Q(sw_rdat[25]));
Q_FDP4EP \sw_rdat_REG[26] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n73), .Q(sw_rdat[26]));
Q_FDP4EP \sw_rdat_REG[27] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n74), .Q(sw_rdat[27]));
Q_FDP4EP \sw_rdat_REG[28] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n75), .Q(sw_rdat[28]));
Q_FDP4EP \sw_rdat_REG[29] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n76), .Q(sw_rdat[29]));
Q_FDP4EP \sw_rdat_REG[30] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n77), .Q(sw_rdat[30]));
Q_FDP4EP \sw_rdat_REG[31] ( .CK(clk), .CE(sw_cs), .R(n1365), .D(n78), .Q(sw_rdat[31]));
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m1 "mem_a 1 31 0 0 31"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_NON_CMM "1"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "rst_dat 1 31 0 0 31"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "1"
// pragma CVASTRPROP MODULE HDLICE PROP_RANOFF TRUE
endmodule
