
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
(* celldefine = 1 *) 
module nx_fifo_ctrl_ram_1r1w_xcm18 ( mem_wen, mem_waddr, mem_wdata, mem_ren, 
	mem_raddr, empty, full, used_slots, free_slots, rerr, rdata, 
	underflow, overflow, clk, rst_n, mem_rdata, mem_ecc_error, wen, 
	wdata, ren, clear);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output mem_wen;
output [7:0] mem_waddr;
output [82:0] mem_wdata;
output mem_ren;
output [7:0] mem_raddr;
output empty;
output full;
output [7:0] used_slots;
output [7:0] free_slots;
output rerr;
output [82:0] rdata;
output underflow;
output overflow;
input clk;
input rst_n;
input [82:0] mem_rdata;
input mem_ecc_error;
input wen;
input [82:0] wdata;
input ren;
input clear;
wire _zy_simnet_mem_wen_0_w$;
wire [0:7] _zy_simnet_mem_waddr_1_w$;
wire [0:82] _zy_simnet_mem_wdata_2_w$;
wire _zy_simnet_mem_ren_3_w$;
wire [0:7] _zy_simnet_mem_raddr_4_w$;
wire _zy_simnet_empty_5_w$;
wire _zy_simnet_full_6_w$;
wire [0:7] _zy_simnet_used_slots_7_w$;
wire [0:7] _zy_simnet_free_slots_8_w$;
wire _zy_simnet_rerr_9_w$;
wire [0:82] _zy_simnet_rdata_10_w$;
wire _zy_simnet_underflow_11_w$;
wire _zy_simnet_overflow_12_w$;
wire _zy_sva__asrtLbl279_1_reset_or;
wire _zy_sva_sf1hot_0;
wire _zyixc_port_1_0_s2hW;
wire [7:0] r_used_slots;
wire [7:0] c_used_slots;
wire [7:0] r_free_slots;
wire [7:0] c_free_slots;
wire [2:0] r_mem_ren_dly;
wire [2:0] c_mem_ren_dly;
wire [7:0] r_mem_wptr;
wire [7:0] c_mem_wptr;
wire [7:0] r_mem_rptr;
wire [7:0] c_mem_rptr;
wire r_mem_empty;
wire c_mem_empty;
wire r_mem_full;
wire c_mem_full;
wire [2:0] r_prefetch_wptr;
wire [2:0] c_prefetch_wptr;
wire [1:0] r_prefetch_rptr;
wire [1:0] c_prefetch_rptr;
wire [1:0] r_prefetch_depth;
wire [1:0] c_prefetch_depth;
wire r_prefetch_empty;
wire c_prefetch_empty;
wire r_prefetch_full;
wire c_prefetch_full;
wire prefetch_wen;
wire [2:0] prefetch_lden_bypass;
wire [2:0] prefetch_lden_mem;
`_2_ wire [2:0] _zy_sva_b0;
`_2_ wire [0:0] _zy_sva__asrtLbl279_1_1_fail;
`_2_ wire _zyixc_port_1_0_req;
`_2_ wire _zyixc_port_1_0_ack;
`_2_ wire _zyixc_port_1_0_isf;
`_2_ wire _zyixc_port_1_0_osf;
supply0 n845;
supply0 n846;
supply0 n847;
Q_BUF U0 ( .A(r_prefetch_wptr[2]), .Z(\c_mem_prefetch_wptr_dly[0][2] ));
Q_BUF U1 ( .A(r_prefetch_wptr[1]), .Z(\c_mem_prefetch_wptr_dly[0][1] ));
Q_BUF U2 ( .A(r_prefetch_wptr[0]), .Z(\c_mem_prefetch_wptr_dly[0][0] ));
Q_BUF U3 ( .A(\r_mem_prefetch_wptr_dly[0][0] ), .Z(\c_mem_prefetch_wptr_dly[1][0] ));
Q_BUF U4 ( .A(\r_mem_prefetch_wptr_dly[0][1] ), .Z(\c_mem_prefetch_wptr_dly[1][1] ));
Q_BUF U5 ( .A(\r_mem_prefetch_wptr_dly[0][2] ), .Z(\c_mem_prefetch_wptr_dly[1][2] ));
Q_BUF U6 ( .A(\r_mem_prefetch_wptr_dly[1][0] ), .Z(\c_mem_prefetch_wptr_dly[2][0] ));
Q_BUF U7 ( .A(\r_mem_prefetch_wptr_dly[1][1] ), .Z(\c_mem_prefetch_wptr_dly[2][1] ));
Q_BUF U8 ( .A(\r_mem_prefetch_wptr_dly[1][2] ), .Z(\c_mem_prefetch_wptr_dly[2][2] ));
Q_BUF U9 ( .A(n845), .Z(n1));
Q_MX03 U10 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][83] ), .A1(\r_prefetch_data[1][83] ), .A2(\r_prefetch_data[2][83] ), .Z(n2));
Q_MX03 U11 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][82] ), .A1(\r_prefetch_data[1][82] ), .A2(\r_prefetch_data[2][82] ), .Z(n3));
Q_MX03 U12 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][81] ), .A1(\r_prefetch_data[1][81] ), .A2(\r_prefetch_data[2][81] ), .Z(n4));
Q_MX03 U13 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][80] ), .A1(\r_prefetch_data[1][80] ), .A2(\r_prefetch_data[2][80] ), .Z(n5));
Q_MX03 U14 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][79] ), .A1(\r_prefetch_data[1][79] ), .A2(\r_prefetch_data[2][79] ), .Z(n6));
Q_MX03 U15 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][78] ), .A1(\r_prefetch_data[1][78] ), .A2(\r_prefetch_data[2][78] ), .Z(n7));
Q_MX03 U16 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][77] ), .A1(\r_prefetch_data[1][77] ), .A2(\r_prefetch_data[2][77] ), .Z(n8));
Q_MX03 U17 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][76] ), .A1(\r_prefetch_data[1][76] ), .A2(\r_prefetch_data[2][76] ), .Z(n9));
Q_MX03 U18 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][75] ), .A1(\r_prefetch_data[1][75] ), .A2(\r_prefetch_data[2][75] ), .Z(n10));
Q_MX03 U19 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][74] ), .A1(\r_prefetch_data[1][74] ), .A2(\r_prefetch_data[2][74] ), .Z(n11));
Q_MX03 U20 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][73] ), .A1(\r_prefetch_data[1][73] ), .A2(\r_prefetch_data[2][73] ), .Z(n12));
Q_MX03 U21 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][72] ), .A1(\r_prefetch_data[1][72] ), .A2(\r_prefetch_data[2][72] ), .Z(n13));
Q_MX03 U22 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][71] ), .A1(\r_prefetch_data[1][71] ), .A2(\r_prefetch_data[2][71] ), .Z(n14));
Q_MX03 U23 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][70] ), .A1(\r_prefetch_data[1][70] ), .A2(\r_prefetch_data[2][70] ), .Z(n15));
Q_MX03 U24 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][69] ), .A1(\r_prefetch_data[1][69] ), .A2(\r_prefetch_data[2][69] ), .Z(n16));
Q_MX03 U25 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][68] ), .A1(\r_prefetch_data[1][68] ), .A2(\r_prefetch_data[2][68] ), .Z(n17));
Q_MX03 U26 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][67] ), .A1(\r_prefetch_data[1][67] ), .A2(\r_prefetch_data[2][67] ), .Z(n18));
Q_MX03 U27 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][66] ), .A1(\r_prefetch_data[1][66] ), .A2(\r_prefetch_data[2][66] ), .Z(n19));
Q_MX03 U28 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][65] ), .A1(\r_prefetch_data[1][65] ), .A2(\r_prefetch_data[2][65] ), .Z(n20));
Q_MX03 U29 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][64] ), .A1(\r_prefetch_data[1][64] ), .A2(\r_prefetch_data[2][64] ), .Z(n21));
Q_MX03 U30 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][63] ), .A1(\r_prefetch_data[1][63] ), .A2(\r_prefetch_data[2][63] ), .Z(n22));
Q_MX03 U31 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][62] ), .A1(\r_prefetch_data[1][62] ), .A2(\r_prefetch_data[2][62] ), .Z(n23));
Q_MX03 U32 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][61] ), .A1(\r_prefetch_data[1][61] ), .A2(\r_prefetch_data[2][61] ), .Z(n24));
Q_MX03 U33 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][60] ), .A1(\r_prefetch_data[1][60] ), .A2(\r_prefetch_data[2][60] ), .Z(n25));
Q_MX03 U34 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][59] ), .A1(\r_prefetch_data[1][59] ), .A2(\r_prefetch_data[2][59] ), .Z(n26));
Q_MX03 U35 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][58] ), .A1(\r_prefetch_data[1][58] ), .A2(\r_prefetch_data[2][58] ), .Z(n27));
Q_MX03 U36 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][57] ), .A1(\r_prefetch_data[1][57] ), .A2(\r_prefetch_data[2][57] ), .Z(n28));
Q_MX03 U37 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][56] ), .A1(\r_prefetch_data[1][56] ), .A2(\r_prefetch_data[2][56] ), .Z(n29));
Q_MX03 U38 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][55] ), .A1(\r_prefetch_data[1][55] ), .A2(\r_prefetch_data[2][55] ), .Z(n30));
Q_MX03 U39 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][54] ), .A1(\r_prefetch_data[1][54] ), .A2(\r_prefetch_data[2][54] ), .Z(n31));
Q_MX03 U40 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][53] ), .A1(\r_prefetch_data[1][53] ), .A2(\r_prefetch_data[2][53] ), .Z(n32));
Q_MX03 U41 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][52] ), .A1(\r_prefetch_data[1][52] ), .A2(\r_prefetch_data[2][52] ), .Z(n33));
Q_MX03 U42 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][51] ), .A1(\r_prefetch_data[1][51] ), .A2(\r_prefetch_data[2][51] ), .Z(n34));
Q_MX03 U43 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][50] ), .A1(\r_prefetch_data[1][50] ), .A2(\r_prefetch_data[2][50] ), .Z(n35));
Q_MX03 U44 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][49] ), .A1(\r_prefetch_data[1][49] ), .A2(\r_prefetch_data[2][49] ), .Z(n36));
Q_MX03 U45 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][48] ), .A1(\r_prefetch_data[1][48] ), .A2(\r_prefetch_data[2][48] ), .Z(n37));
Q_MX03 U46 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][47] ), .A1(\r_prefetch_data[1][47] ), .A2(\r_prefetch_data[2][47] ), .Z(n38));
Q_MX03 U47 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][46] ), .A1(\r_prefetch_data[1][46] ), .A2(\r_prefetch_data[2][46] ), .Z(n39));
Q_MX03 U48 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][45] ), .A1(\r_prefetch_data[1][45] ), .A2(\r_prefetch_data[2][45] ), .Z(n40));
Q_MX03 U49 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][44] ), .A1(\r_prefetch_data[1][44] ), .A2(\r_prefetch_data[2][44] ), .Z(n41));
Q_MX03 U50 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][43] ), .A1(\r_prefetch_data[1][43] ), .A2(\r_prefetch_data[2][43] ), .Z(n42));
Q_MX03 U51 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][42] ), .A1(\r_prefetch_data[1][42] ), .A2(\r_prefetch_data[2][42] ), .Z(n43));
Q_MX03 U52 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][41] ), .A1(\r_prefetch_data[1][41] ), .A2(\r_prefetch_data[2][41] ), .Z(n44));
Q_MX03 U53 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][40] ), .A1(\r_prefetch_data[1][40] ), .A2(\r_prefetch_data[2][40] ), .Z(n45));
Q_MX03 U54 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][39] ), .A1(\r_prefetch_data[1][39] ), .A2(\r_prefetch_data[2][39] ), .Z(n46));
Q_MX03 U55 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][38] ), .A1(\r_prefetch_data[1][38] ), .A2(\r_prefetch_data[2][38] ), .Z(n47));
Q_MX03 U56 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][37] ), .A1(\r_prefetch_data[1][37] ), .A2(\r_prefetch_data[2][37] ), .Z(n48));
Q_MX03 U57 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][36] ), .A1(\r_prefetch_data[1][36] ), .A2(\r_prefetch_data[2][36] ), .Z(n49));
Q_MX03 U58 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][35] ), .A1(\r_prefetch_data[1][35] ), .A2(\r_prefetch_data[2][35] ), .Z(n50));
Q_MX03 U59 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][34] ), .A1(\r_prefetch_data[1][34] ), .A2(\r_prefetch_data[2][34] ), .Z(n51));
Q_MX03 U60 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][33] ), .A1(\r_prefetch_data[1][33] ), .A2(\r_prefetch_data[2][33] ), .Z(n52));
Q_MX03 U61 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][32] ), .A1(\r_prefetch_data[1][32] ), .A2(\r_prefetch_data[2][32] ), .Z(n53));
Q_MX03 U62 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][31] ), .A1(\r_prefetch_data[1][31] ), .A2(\r_prefetch_data[2][31] ), .Z(n54));
Q_MX03 U63 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][30] ), .A1(\r_prefetch_data[1][30] ), .A2(\r_prefetch_data[2][30] ), .Z(n55));
Q_MX03 U64 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][29] ), .A1(\r_prefetch_data[1][29] ), .A2(\r_prefetch_data[2][29] ), .Z(n56));
Q_MX03 U65 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][28] ), .A1(\r_prefetch_data[1][28] ), .A2(\r_prefetch_data[2][28] ), .Z(n57));
Q_MX03 U66 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][27] ), .A1(\r_prefetch_data[1][27] ), .A2(\r_prefetch_data[2][27] ), .Z(n58));
Q_MX03 U67 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][26] ), .A1(\r_prefetch_data[1][26] ), .A2(\r_prefetch_data[2][26] ), .Z(n59));
Q_MX03 U68 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][25] ), .A1(\r_prefetch_data[1][25] ), .A2(\r_prefetch_data[2][25] ), .Z(n60));
Q_MX03 U69 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][24] ), .A1(\r_prefetch_data[1][24] ), .A2(\r_prefetch_data[2][24] ), .Z(n61));
Q_MX03 U70 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][23] ), .A1(\r_prefetch_data[1][23] ), .A2(\r_prefetch_data[2][23] ), .Z(n62));
Q_MX03 U71 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][22] ), .A1(\r_prefetch_data[1][22] ), .A2(\r_prefetch_data[2][22] ), .Z(n63));
Q_MX03 U72 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][21] ), .A1(\r_prefetch_data[1][21] ), .A2(\r_prefetch_data[2][21] ), .Z(n64));
Q_MX03 U73 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][20] ), .A1(\r_prefetch_data[1][20] ), .A2(\r_prefetch_data[2][20] ), .Z(n65));
Q_MX03 U74 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][19] ), .A1(\r_prefetch_data[1][19] ), .A2(\r_prefetch_data[2][19] ), .Z(n66));
Q_MX03 U75 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][18] ), .A1(\r_prefetch_data[1][18] ), .A2(\r_prefetch_data[2][18] ), .Z(n67));
Q_MX03 U76 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][17] ), .A1(\r_prefetch_data[1][17] ), .A2(\r_prefetch_data[2][17] ), .Z(n68));
Q_MX03 U77 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][16] ), .A1(\r_prefetch_data[1][16] ), .A2(\r_prefetch_data[2][16] ), .Z(n69));
Q_MX03 U78 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][15] ), .A1(\r_prefetch_data[1][15] ), .A2(\r_prefetch_data[2][15] ), .Z(n70));
Q_MX03 U79 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][14] ), .A1(\r_prefetch_data[1][14] ), .A2(\r_prefetch_data[2][14] ), .Z(n71));
Q_MX03 U80 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][13] ), .A1(\r_prefetch_data[1][13] ), .A2(\r_prefetch_data[2][13] ), .Z(n72));
Q_MX03 U81 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][12] ), .A1(\r_prefetch_data[1][12] ), .A2(\r_prefetch_data[2][12] ), .Z(n73));
Q_MX03 U82 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][11] ), .A1(\r_prefetch_data[1][11] ), .A2(\r_prefetch_data[2][11] ), .Z(n74));
Q_MX03 U83 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][10] ), .A1(\r_prefetch_data[1][10] ), .A2(\r_prefetch_data[2][10] ), .Z(n75));
Q_MX03 U84 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][9] ), .A1(\r_prefetch_data[1][9] ), .A2(\r_prefetch_data[2][9] ), .Z(n76));
Q_MX03 U85 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][8] ), .A1(\r_prefetch_data[1][8] ), .A2(\r_prefetch_data[2][8] ), .Z(n77));
Q_MX03 U86 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][7] ), .A1(\r_prefetch_data[1][7] ), .A2(\r_prefetch_data[2][7] ), .Z(n78));
Q_MX03 U87 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][6] ), .A1(\r_prefetch_data[1][6] ), .A2(\r_prefetch_data[2][6] ), .Z(n79));
Q_MX03 U88 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][5] ), .A1(\r_prefetch_data[1][5] ), .A2(\r_prefetch_data[2][5] ), .Z(n80));
Q_MX03 U89 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][4] ), .A1(\r_prefetch_data[1][4] ), .A2(\r_prefetch_data[2][4] ), .Z(n81));
Q_MX03 U90 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][3] ), .A1(\r_prefetch_data[1][3] ), .A2(\r_prefetch_data[2][3] ), .Z(n82));
Q_MX03 U91 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][2] ), .A1(\r_prefetch_data[1][2] ), .A2(\r_prefetch_data[2][2] ), .Z(n83));
Q_MX03 U92 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][1] ), .A1(\r_prefetch_data[1][1] ), .A2(\r_prefetch_data[2][1] ), .Z(n84));
Q_MX03 U93 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][0] ), .A1(\r_prefetch_data[1][0] ), .A2(\r_prefetch_data[2][0] ), .Z(n85));
Q_FDP0 \r_mem_prefetch_wptr_dly_REG[2][2] ( .CK(clk), .D(\c_mem_prefetch_wptr_dly[2][2] ), .Q(\r_mem_prefetch_wptr_dly[2][2] ), .QN( ));
Q_FDP0 \r_mem_prefetch_wptr_dly_REG[2][1] ( .CK(clk), .D(\c_mem_prefetch_wptr_dly[2][1] ), .Q(\r_mem_prefetch_wptr_dly[2][1] ), .QN( ));
Q_FDP0 \r_mem_prefetch_wptr_dly_REG[2][0] ( .CK(clk), .D(\c_mem_prefetch_wptr_dly[2][0] ), .Q(\r_mem_prefetch_wptr_dly[2][0] ), .QN( ));
Q_FDP0 \r_mem_prefetch_wptr_dly_REG[1][2] ( .CK(clk), .D(\c_mem_prefetch_wptr_dly[1][2] ), .Q(\r_mem_prefetch_wptr_dly[1][2] ), .QN( ));
Q_FDP0 \r_mem_prefetch_wptr_dly_REG[1][1] ( .CK(clk), .D(\c_mem_prefetch_wptr_dly[1][1] ), .Q(\r_mem_prefetch_wptr_dly[1][1] ), .QN( ));
Q_FDP0 \r_mem_prefetch_wptr_dly_REG[1][0] ( .CK(clk), .D(\c_mem_prefetch_wptr_dly[1][0] ), .Q(\r_mem_prefetch_wptr_dly[1][0] ), .QN( ));
Q_FDP0 \r_mem_prefetch_wptr_dly_REG[0][2] ( .CK(clk), .D(\c_mem_prefetch_wptr_dly[0][2] ), .Q(\r_mem_prefetch_wptr_dly[0][2] ), .QN( ));
Q_FDP0 \r_mem_prefetch_wptr_dly_REG[0][1] ( .CK(clk), .D(\c_mem_prefetch_wptr_dly[0][1] ), .Q(\r_mem_prefetch_wptr_dly[0][1] ), .QN( ));
Q_FDP0 \r_mem_prefetch_wptr_dly_REG[0][0] ( .CK(clk), .D(\c_mem_prefetch_wptr_dly[0][0] ), .Q(\r_mem_prefetch_wptr_dly[0][0] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][83] ( .CK(clk), .D(\c_prefetch_data[2][83] ), .Q(\r_prefetch_data[2][83] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][82] ( .CK(clk), .D(\c_prefetch_data[2][82] ), .Q(\r_prefetch_data[2][82] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][81] ( .CK(clk), .D(\c_prefetch_data[2][81] ), .Q(\r_prefetch_data[2][81] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][80] ( .CK(clk), .D(\c_prefetch_data[2][80] ), .Q(\r_prefetch_data[2][80] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][79] ( .CK(clk), .D(\c_prefetch_data[2][79] ), .Q(\r_prefetch_data[2][79] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][78] ( .CK(clk), .D(\c_prefetch_data[2][78] ), .Q(\r_prefetch_data[2][78] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][77] ( .CK(clk), .D(\c_prefetch_data[2][77] ), .Q(\r_prefetch_data[2][77] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][76] ( .CK(clk), .D(\c_prefetch_data[2][76] ), .Q(\r_prefetch_data[2][76] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][75] ( .CK(clk), .D(\c_prefetch_data[2][75] ), .Q(\r_prefetch_data[2][75] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][74] ( .CK(clk), .D(\c_prefetch_data[2][74] ), .Q(\r_prefetch_data[2][74] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][73] ( .CK(clk), .D(\c_prefetch_data[2][73] ), .Q(\r_prefetch_data[2][73] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][72] ( .CK(clk), .D(\c_prefetch_data[2][72] ), .Q(\r_prefetch_data[2][72] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][71] ( .CK(clk), .D(\c_prefetch_data[2][71] ), .Q(\r_prefetch_data[2][71] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][70] ( .CK(clk), .D(\c_prefetch_data[2][70] ), .Q(\r_prefetch_data[2][70] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][69] ( .CK(clk), .D(\c_prefetch_data[2][69] ), .Q(\r_prefetch_data[2][69] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][68] ( .CK(clk), .D(\c_prefetch_data[2][68] ), .Q(\r_prefetch_data[2][68] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][67] ( .CK(clk), .D(\c_prefetch_data[2][67] ), .Q(\r_prefetch_data[2][67] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][66] ( .CK(clk), .D(\c_prefetch_data[2][66] ), .Q(\r_prefetch_data[2][66] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][65] ( .CK(clk), .D(\c_prefetch_data[2][65] ), .Q(\r_prefetch_data[2][65] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][64] ( .CK(clk), .D(\c_prefetch_data[2][64] ), .Q(\r_prefetch_data[2][64] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][63] ( .CK(clk), .D(\c_prefetch_data[2][63] ), .Q(\r_prefetch_data[2][63] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][62] ( .CK(clk), .D(\c_prefetch_data[2][62] ), .Q(\r_prefetch_data[2][62] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][61] ( .CK(clk), .D(\c_prefetch_data[2][61] ), .Q(\r_prefetch_data[2][61] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][60] ( .CK(clk), .D(\c_prefetch_data[2][60] ), .Q(\r_prefetch_data[2][60] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][59] ( .CK(clk), .D(\c_prefetch_data[2][59] ), .Q(\r_prefetch_data[2][59] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][58] ( .CK(clk), .D(\c_prefetch_data[2][58] ), .Q(\r_prefetch_data[2][58] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][57] ( .CK(clk), .D(\c_prefetch_data[2][57] ), .Q(\r_prefetch_data[2][57] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][56] ( .CK(clk), .D(\c_prefetch_data[2][56] ), .Q(\r_prefetch_data[2][56] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][55] ( .CK(clk), .D(\c_prefetch_data[2][55] ), .Q(\r_prefetch_data[2][55] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][54] ( .CK(clk), .D(\c_prefetch_data[2][54] ), .Q(\r_prefetch_data[2][54] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][53] ( .CK(clk), .D(\c_prefetch_data[2][53] ), .Q(\r_prefetch_data[2][53] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][52] ( .CK(clk), .D(\c_prefetch_data[2][52] ), .Q(\r_prefetch_data[2][52] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][51] ( .CK(clk), .D(\c_prefetch_data[2][51] ), .Q(\r_prefetch_data[2][51] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][50] ( .CK(clk), .D(\c_prefetch_data[2][50] ), .Q(\r_prefetch_data[2][50] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][49] ( .CK(clk), .D(\c_prefetch_data[2][49] ), .Q(\r_prefetch_data[2][49] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][48] ( .CK(clk), .D(\c_prefetch_data[2][48] ), .Q(\r_prefetch_data[2][48] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][47] ( .CK(clk), .D(\c_prefetch_data[2][47] ), .Q(\r_prefetch_data[2][47] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][46] ( .CK(clk), .D(\c_prefetch_data[2][46] ), .Q(\r_prefetch_data[2][46] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][45] ( .CK(clk), .D(\c_prefetch_data[2][45] ), .Q(\r_prefetch_data[2][45] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][44] ( .CK(clk), .D(\c_prefetch_data[2][44] ), .Q(\r_prefetch_data[2][44] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][43] ( .CK(clk), .D(\c_prefetch_data[2][43] ), .Q(\r_prefetch_data[2][43] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][42] ( .CK(clk), .D(\c_prefetch_data[2][42] ), .Q(\r_prefetch_data[2][42] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][41] ( .CK(clk), .D(\c_prefetch_data[2][41] ), .Q(\r_prefetch_data[2][41] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][40] ( .CK(clk), .D(\c_prefetch_data[2][40] ), .Q(\r_prefetch_data[2][40] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][39] ( .CK(clk), .D(\c_prefetch_data[2][39] ), .Q(\r_prefetch_data[2][39] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][38] ( .CK(clk), .D(\c_prefetch_data[2][38] ), .Q(\r_prefetch_data[2][38] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][37] ( .CK(clk), .D(\c_prefetch_data[2][37] ), .Q(\r_prefetch_data[2][37] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][36] ( .CK(clk), .D(\c_prefetch_data[2][36] ), .Q(\r_prefetch_data[2][36] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][35] ( .CK(clk), .D(\c_prefetch_data[2][35] ), .Q(\r_prefetch_data[2][35] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][34] ( .CK(clk), .D(\c_prefetch_data[2][34] ), .Q(\r_prefetch_data[2][34] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][33] ( .CK(clk), .D(\c_prefetch_data[2][33] ), .Q(\r_prefetch_data[2][33] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][32] ( .CK(clk), .D(\c_prefetch_data[2][32] ), .Q(\r_prefetch_data[2][32] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][31] ( .CK(clk), .D(\c_prefetch_data[2][31] ), .Q(\r_prefetch_data[2][31] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][30] ( .CK(clk), .D(\c_prefetch_data[2][30] ), .Q(\r_prefetch_data[2][30] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][29] ( .CK(clk), .D(\c_prefetch_data[2][29] ), .Q(\r_prefetch_data[2][29] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][28] ( .CK(clk), .D(\c_prefetch_data[2][28] ), .Q(\r_prefetch_data[2][28] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][27] ( .CK(clk), .D(\c_prefetch_data[2][27] ), .Q(\r_prefetch_data[2][27] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][26] ( .CK(clk), .D(\c_prefetch_data[2][26] ), .Q(\r_prefetch_data[2][26] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][25] ( .CK(clk), .D(\c_prefetch_data[2][25] ), .Q(\r_prefetch_data[2][25] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][24] ( .CK(clk), .D(\c_prefetch_data[2][24] ), .Q(\r_prefetch_data[2][24] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][23] ( .CK(clk), .D(\c_prefetch_data[2][23] ), .Q(\r_prefetch_data[2][23] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][22] ( .CK(clk), .D(\c_prefetch_data[2][22] ), .Q(\r_prefetch_data[2][22] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][21] ( .CK(clk), .D(\c_prefetch_data[2][21] ), .Q(\r_prefetch_data[2][21] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][20] ( .CK(clk), .D(\c_prefetch_data[2][20] ), .Q(\r_prefetch_data[2][20] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][19] ( .CK(clk), .D(\c_prefetch_data[2][19] ), .Q(\r_prefetch_data[2][19] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][18] ( .CK(clk), .D(\c_prefetch_data[2][18] ), .Q(\r_prefetch_data[2][18] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][17] ( .CK(clk), .D(\c_prefetch_data[2][17] ), .Q(\r_prefetch_data[2][17] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][16] ( .CK(clk), .D(\c_prefetch_data[2][16] ), .Q(\r_prefetch_data[2][16] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][15] ( .CK(clk), .D(\c_prefetch_data[2][15] ), .Q(\r_prefetch_data[2][15] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][14] ( .CK(clk), .D(\c_prefetch_data[2][14] ), .Q(\r_prefetch_data[2][14] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][13] ( .CK(clk), .D(\c_prefetch_data[2][13] ), .Q(\r_prefetch_data[2][13] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][12] ( .CK(clk), .D(\c_prefetch_data[2][12] ), .Q(\r_prefetch_data[2][12] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][11] ( .CK(clk), .D(\c_prefetch_data[2][11] ), .Q(\r_prefetch_data[2][11] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][10] ( .CK(clk), .D(\c_prefetch_data[2][10] ), .Q(\r_prefetch_data[2][10] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][9] ( .CK(clk), .D(\c_prefetch_data[2][9] ), .Q(\r_prefetch_data[2][9] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][8] ( .CK(clk), .D(\c_prefetch_data[2][8] ), .Q(\r_prefetch_data[2][8] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][7] ( .CK(clk), .D(\c_prefetch_data[2][7] ), .Q(\r_prefetch_data[2][7] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][6] ( .CK(clk), .D(\c_prefetch_data[2][6] ), .Q(\r_prefetch_data[2][6] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][5] ( .CK(clk), .D(\c_prefetch_data[2][5] ), .Q(\r_prefetch_data[2][5] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][4] ( .CK(clk), .D(\c_prefetch_data[2][4] ), .Q(\r_prefetch_data[2][4] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][3] ( .CK(clk), .D(\c_prefetch_data[2][3] ), .Q(\r_prefetch_data[2][3] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][2] ( .CK(clk), .D(\c_prefetch_data[2][2] ), .Q(\r_prefetch_data[2][2] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][1] ( .CK(clk), .D(\c_prefetch_data[2][1] ), .Q(\r_prefetch_data[2][1] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][0] ( .CK(clk), .D(\c_prefetch_data[2][0] ), .Q(\r_prefetch_data[2][0] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][83] ( .CK(clk), .D(\c_prefetch_data[1][83] ), .Q(\r_prefetch_data[1][83] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][82] ( .CK(clk), .D(\c_prefetch_data[1][82] ), .Q(\r_prefetch_data[1][82] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][81] ( .CK(clk), .D(\c_prefetch_data[1][81] ), .Q(\r_prefetch_data[1][81] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][80] ( .CK(clk), .D(\c_prefetch_data[1][80] ), .Q(\r_prefetch_data[1][80] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][79] ( .CK(clk), .D(\c_prefetch_data[1][79] ), .Q(\r_prefetch_data[1][79] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][78] ( .CK(clk), .D(\c_prefetch_data[1][78] ), .Q(\r_prefetch_data[1][78] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][77] ( .CK(clk), .D(\c_prefetch_data[1][77] ), .Q(\r_prefetch_data[1][77] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][76] ( .CK(clk), .D(\c_prefetch_data[1][76] ), .Q(\r_prefetch_data[1][76] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][75] ( .CK(clk), .D(\c_prefetch_data[1][75] ), .Q(\r_prefetch_data[1][75] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][74] ( .CK(clk), .D(\c_prefetch_data[1][74] ), .Q(\r_prefetch_data[1][74] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][73] ( .CK(clk), .D(\c_prefetch_data[1][73] ), .Q(\r_prefetch_data[1][73] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][72] ( .CK(clk), .D(\c_prefetch_data[1][72] ), .Q(\r_prefetch_data[1][72] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][71] ( .CK(clk), .D(\c_prefetch_data[1][71] ), .Q(\r_prefetch_data[1][71] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][70] ( .CK(clk), .D(\c_prefetch_data[1][70] ), .Q(\r_prefetch_data[1][70] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][69] ( .CK(clk), .D(\c_prefetch_data[1][69] ), .Q(\r_prefetch_data[1][69] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][68] ( .CK(clk), .D(\c_prefetch_data[1][68] ), .Q(\r_prefetch_data[1][68] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][67] ( .CK(clk), .D(\c_prefetch_data[1][67] ), .Q(\r_prefetch_data[1][67] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][66] ( .CK(clk), .D(\c_prefetch_data[1][66] ), .Q(\r_prefetch_data[1][66] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][65] ( .CK(clk), .D(\c_prefetch_data[1][65] ), .Q(\r_prefetch_data[1][65] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][64] ( .CK(clk), .D(\c_prefetch_data[1][64] ), .Q(\r_prefetch_data[1][64] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][63] ( .CK(clk), .D(\c_prefetch_data[1][63] ), .Q(\r_prefetch_data[1][63] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][62] ( .CK(clk), .D(\c_prefetch_data[1][62] ), .Q(\r_prefetch_data[1][62] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][61] ( .CK(clk), .D(\c_prefetch_data[1][61] ), .Q(\r_prefetch_data[1][61] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][60] ( .CK(clk), .D(\c_prefetch_data[1][60] ), .Q(\r_prefetch_data[1][60] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][59] ( .CK(clk), .D(\c_prefetch_data[1][59] ), .Q(\r_prefetch_data[1][59] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][58] ( .CK(clk), .D(\c_prefetch_data[1][58] ), .Q(\r_prefetch_data[1][58] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][57] ( .CK(clk), .D(\c_prefetch_data[1][57] ), .Q(\r_prefetch_data[1][57] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][56] ( .CK(clk), .D(\c_prefetch_data[1][56] ), .Q(\r_prefetch_data[1][56] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][55] ( .CK(clk), .D(\c_prefetch_data[1][55] ), .Q(\r_prefetch_data[1][55] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][54] ( .CK(clk), .D(\c_prefetch_data[1][54] ), .Q(\r_prefetch_data[1][54] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][53] ( .CK(clk), .D(\c_prefetch_data[1][53] ), .Q(\r_prefetch_data[1][53] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][52] ( .CK(clk), .D(\c_prefetch_data[1][52] ), .Q(\r_prefetch_data[1][52] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][51] ( .CK(clk), .D(\c_prefetch_data[1][51] ), .Q(\r_prefetch_data[1][51] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][50] ( .CK(clk), .D(\c_prefetch_data[1][50] ), .Q(\r_prefetch_data[1][50] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][49] ( .CK(clk), .D(\c_prefetch_data[1][49] ), .Q(\r_prefetch_data[1][49] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][48] ( .CK(clk), .D(\c_prefetch_data[1][48] ), .Q(\r_prefetch_data[1][48] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][47] ( .CK(clk), .D(\c_prefetch_data[1][47] ), .Q(\r_prefetch_data[1][47] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][46] ( .CK(clk), .D(\c_prefetch_data[1][46] ), .Q(\r_prefetch_data[1][46] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][45] ( .CK(clk), .D(\c_prefetch_data[1][45] ), .Q(\r_prefetch_data[1][45] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][44] ( .CK(clk), .D(\c_prefetch_data[1][44] ), .Q(\r_prefetch_data[1][44] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][43] ( .CK(clk), .D(\c_prefetch_data[1][43] ), .Q(\r_prefetch_data[1][43] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][42] ( .CK(clk), .D(\c_prefetch_data[1][42] ), .Q(\r_prefetch_data[1][42] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][41] ( .CK(clk), .D(\c_prefetch_data[1][41] ), .Q(\r_prefetch_data[1][41] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][40] ( .CK(clk), .D(\c_prefetch_data[1][40] ), .Q(\r_prefetch_data[1][40] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][39] ( .CK(clk), .D(\c_prefetch_data[1][39] ), .Q(\r_prefetch_data[1][39] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][38] ( .CK(clk), .D(\c_prefetch_data[1][38] ), .Q(\r_prefetch_data[1][38] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][37] ( .CK(clk), .D(\c_prefetch_data[1][37] ), .Q(\r_prefetch_data[1][37] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][36] ( .CK(clk), .D(\c_prefetch_data[1][36] ), .Q(\r_prefetch_data[1][36] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][35] ( .CK(clk), .D(\c_prefetch_data[1][35] ), .Q(\r_prefetch_data[1][35] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][34] ( .CK(clk), .D(\c_prefetch_data[1][34] ), .Q(\r_prefetch_data[1][34] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][33] ( .CK(clk), .D(\c_prefetch_data[1][33] ), .Q(\r_prefetch_data[1][33] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][32] ( .CK(clk), .D(\c_prefetch_data[1][32] ), .Q(\r_prefetch_data[1][32] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][31] ( .CK(clk), .D(\c_prefetch_data[1][31] ), .Q(\r_prefetch_data[1][31] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][30] ( .CK(clk), .D(\c_prefetch_data[1][30] ), .Q(\r_prefetch_data[1][30] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][29] ( .CK(clk), .D(\c_prefetch_data[1][29] ), .Q(\r_prefetch_data[1][29] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][28] ( .CK(clk), .D(\c_prefetch_data[1][28] ), .Q(\r_prefetch_data[1][28] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][27] ( .CK(clk), .D(\c_prefetch_data[1][27] ), .Q(\r_prefetch_data[1][27] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][26] ( .CK(clk), .D(\c_prefetch_data[1][26] ), .Q(\r_prefetch_data[1][26] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][25] ( .CK(clk), .D(\c_prefetch_data[1][25] ), .Q(\r_prefetch_data[1][25] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][24] ( .CK(clk), .D(\c_prefetch_data[1][24] ), .Q(\r_prefetch_data[1][24] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][23] ( .CK(clk), .D(\c_prefetch_data[1][23] ), .Q(\r_prefetch_data[1][23] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][22] ( .CK(clk), .D(\c_prefetch_data[1][22] ), .Q(\r_prefetch_data[1][22] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][21] ( .CK(clk), .D(\c_prefetch_data[1][21] ), .Q(\r_prefetch_data[1][21] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][20] ( .CK(clk), .D(\c_prefetch_data[1][20] ), .Q(\r_prefetch_data[1][20] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][19] ( .CK(clk), .D(\c_prefetch_data[1][19] ), .Q(\r_prefetch_data[1][19] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][18] ( .CK(clk), .D(\c_prefetch_data[1][18] ), .Q(\r_prefetch_data[1][18] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][17] ( .CK(clk), .D(\c_prefetch_data[1][17] ), .Q(\r_prefetch_data[1][17] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][16] ( .CK(clk), .D(\c_prefetch_data[1][16] ), .Q(\r_prefetch_data[1][16] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][15] ( .CK(clk), .D(\c_prefetch_data[1][15] ), .Q(\r_prefetch_data[1][15] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][14] ( .CK(clk), .D(\c_prefetch_data[1][14] ), .Q(\r_prefetch_data[1][14] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][13] ( .CK(clk), .D(\c_prefetch_data[1][13] ), .Q(\r_prefetch_data[1][13] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][12] ( .CK(clk), .D(\c_prefetch_data[1][12] ), .Q(\r_prefetch_data[1][12] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][11] ( .CK(clk), .D(\c_prefetch_data[1][11] ), .Q(\r_prefetch_data[1][11] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][10] ( .CK(clk), .D(\c_prefetch_data[1][10] ), .Q(\r_prefetch_data[1][10] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][9] ( .CK(clk), .D(\c_prefetch_data[1][9] ), .Q(\r_prefetch_data[1][9] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][8] ( .CK(clk), .D(\c_prefetch_data[1][8] ), .Q(\r_prefetch_data[1][8] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][7] ( .CK(clk), .D(\c_prefetch_data[1][7] ), .Q(\r_prefetch_data[1][7] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][6] ( .CK(clk), .D(\c_prefetch_data[1][6] ), .Q(\r_prefetch_data[1][6] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][5] ( .CK(clk), .D(\c_prefetch_data[1][5] ), .Q(\r_prefetch_data[1][5] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][4] ( .CK(clk), .D(\c_prefetch_data[1][4] ), .Q(\r_prefetch_data[1][4] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][3] ( .CK(clk), .D(\c_prefetch_data[1][3] ), .Q(\r_prefetch_data[1][3] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][2] ( .CK(clk), .D(\c_prefetch_data[1][2] ), .Q(\r_prefetch_data[1][2] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][1] ( .CK(clk), .D(\c_prefetch_data[1][1] ), .Q(\r_prefetch_data[1][1] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][0] ( .CK(clk), .D(\c_prefetch_data[1][0] ), .Q(\r_prefetch_data[1][0] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][83] ( .CK(clk), .D(\c_prefetch_data[0][83] ), .Q(\r_prefetch_data[0][83] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][82] ( .CK(clk), .D(\c_prefetch_data[0][82] ), .Q(\r_prefetch_data[0][82] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][81] ( .CK(clk), .D(\c_prefetch_data[0][81] ), .Q(\r_prefetch_data[0][81] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][80] ( .CK(clk), .D(\c_prefetch_data[0][80] ), .Q(\r_prefetch_data[0][80] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][79] ( .CK(clk), .D(\c_prefetch_data[0][79] ), .Q(\r_prefetch_data[0][79] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][78] ( .CK(clk), .D(\c_prefetch_data[0][78] ), .Q(\r_prefetch_data[0][78] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][77] ( .CK(clk), .D(\c_prefetch_data[0][77] ), .Q(\r_prefetch_data[0][77] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][76] ( .CK(clk), .D(\c_prefetch_data[0][76] ), .Q(\r_prefetch_data[0][76] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][75] ( .CK(clk), .D(\c_prefetch_data[0][75] ), .Q(\r_prefetch_data[0][75] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][74] ( .CK(clk), .D(\c_prefetch_data[0][74] ), .Q(\r_prefetch_data[0][74] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][73] ( .CK(clk), .D(\c_prefetch_data[0][73] ), .Q(\r_prefetch_data[0][73] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][72] ( .CK(clk), .D(\c_prefetch_data[0][72] ), .Q(\r_prefetch_data[0][72] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][71] ( .CK(clk), .D(\c_prefetch_data[0][71] ), .Q(\r_prefetch_data[0][71] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][70] ( .CK(clk), .D(\c_prefetch_data[0][70] ), .Q(\r_prefetch_data[0][70] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][69] ( .CK(clk), .D(\c_prefetch_data[0][69] ), .Q(\r_prefetch_data[0][69] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][68] ( .CK(clk), .D(\c_prefetch_data[0][68] ), .Q(\r_prefetch_data[0][68] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][67] ( .CK(clk), .D(\c_prefetch_data[0][67] ), .Q(\r_prefetch_data[0][67] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][66] ( .CK(clk), .D(\c_prefetch_data[0][66] ), .Q(\r_prefetch_data[0][66] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][65] ( .CK(clk), .D(\c_prefetch_data[0][65] ), .Q(\r_prefetch_data[0][65] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][64] ( .CK(clk), .D(\c_prefetch_data[0][64] ), .Q(\r_prefetch_data[0][64] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][63] ( .CK(clk), .D(\c_prefetch_data[0][63] ), .Q(\r_prefetch_data[0][63] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][62] ( .CK(clk), .D(\c_prefetch_data[0][62] ), .Q(\r_prefetch_data[0][62] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][61] ( .CK(clk), .D(\c_prefetch_data[0][61] ), .Q(\r_prefetch_data[0][61] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][60] ( .CK(clk), .D(\c_prefetch_data[0][60] ), .Q(\r_prefetch_data[0][60] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][59] ( .CK(clk), .D(\c_prefetch_data[0][59] ), .Q(\r_prefetch_data[0][59] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][58] ( .CK(clk), .D(\c_prefetch_data[0][58] ), .Q(\r_prefetch_data[0][58] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][57] ( .CK(clk), .D(\c_prefetch_data[0][57] ), .Q(\r_prefetch_data[0][57] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][56] ( .CK(clk), .D(\c_prefetch_data[0][56] ), .Q(\r_prefetch_data[0][56] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][55] ( .CK(clk), .D(\c_prefetch_data[0][55] ), .Q(\r_prefetch_data[0][55] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][54] ( .CK(clk), .D(\c_prefetch_data[0][54] ), .Q(\r_prefetch_data[0][54] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][53] ( .CK(clk), .D(\c_prefetch_data[0][53] ), .Q(\r_prefetch_data[0][53] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][52] ( .CK(clk), .D(\c_prefetch_data[0][52] ), .Q(\r_prefetch_data[0][52] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][51] ( .CK(clk), .D(\c_prefetch_data[0][51] ), .Q(\r_prefetch_data[0][51] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][50] ( .CK(clk), .D(\c_prefetch_data[0][50] ), .Q(\r_prefetch_data[0][50] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][49] ( .CK(clk), .D(\c_prefetch_data[0][49] ), .Q(\r_prefetch_data[0][49] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][48] ( .CK(clk), .D(\c_prefetch_data[0][48] ), .Q(\r_prefetch_data[0][48] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][47] ( .CK(clk), .D(\c_prefetch_data[0][47] ), .Q(\r_prefetch_data[0][47] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][46] ( .CK(clk), .D(\c_prefetch_data[0][46] ), .Q(\r_prefetch_data[0][46] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][45] ( .CK(clk), .D(\c_prefetch_data[0][45] ), .Q(\r_prefetch_data[0][45] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][44] ( .CK(clk), .D(\c_prefetch_data[0][44] ), .Q(\r_prefetch_data[0][44] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][43] ( .CK(clk), .D(\c_prefetch_data[0][43] ), .Q(\r_prefetch_data[0][43] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][42] ( .CK(clk), .D(\c_prefetch_data[0][42] ), .Q(\r_prefetch_data[0][42] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][41] ( .CK(clk), .D(\c_prefetch_data[0][41] ), .Q(\r_prefetch_data[0][41] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][40] ( .CK(clk), .D(\c_prefetch_data[0][40] ), .Q(\r_prefetch_data[0][40] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][39] ( .CK(clk), .D(\c_prefetch_data[0][39] ), .Q(\r_prefetch_data[0][39] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][38] ( .CK(clk), .D(\c_prefetch_data[0][38] ), .Q(\r_prefetch_data[0][38] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][37] ( .CK(clk), .D(\c_prefetch_data[0][37] ), .Q(\r_prefetch_data[0][37] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][36] ( .CK(clk), .D(\c_prefetch_data[0][36] ), .Q(\r_prefetch_data[0][36] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][35] ( .CK(clk), .D(\c_prefetch_data[0][35] ), .Q(\r_prefetch_data[0][35] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][34] ( .CK(clk), .D(\c_prefetch_data[0][34] ), .Q(\r_prefetch_data[0][34] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][33] ( .CK(clk), .D(\c_prefetch_data[0][33] ), .Q(\r_prefetch_data[0][33] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][32] ( .CK(clk), .D(\c_prefetch_data[0][32] ), .Q(\r_prefetch_data[0][32] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][31] ( .CK(clk), .D(\c_prefetch_data[0][31] ), .Q(\r_prefetch_data[0][31] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][30] ( .CK(clk), .D(\c_prefetch_data[0][30] ), .Q(\r_prefetch_data[0][30] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][29] ( .CK(clk), .D(\c_prefetch_data[0][29] ), .Q(\r_prefetch_data[0][29] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][28] ( .CK(clk), .D(\c_prefetch_data[0][28] ), .Q(\r_prefetch_data[0][28] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][27] ( .CK(clk), .D(\c_prefetch_data[0][27] ), .Q(\r_prefetch_data[0][27] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][26] ( .CK(clk), .D(\c_prefetch_data[0][26] ), .Q(\r_prefetch_data[0][26] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][25] ( .CK(clk), .D(\c_prefetch_data[0][25] ), .Q(\r_prefetch_data[0][25] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][24] ( .CK(clk), .D(\c_prefetch_data[0][24] ), .Q(\r_prefetch_data[0][24] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][23] ( .CK(clk), .D(\c_prefetch_data[0][23] ), .Q(\r_prefetch_data[0][23] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][22] ( .CK(clk), .D(\c_prefetch_data[0][22] ), .Q(\r_prefetch_data[0][22] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][21] ( .CK(clk), .D(\c_prefetch_data[0][21] ), .Q(\r_prefetch_data[0][21] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][20] ( .CK(clk), .D(\c_prefetch_data[0][20] ), .Q(\r_prefetch_data[0][20] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][19] ( .CK(clk), .D(\c_prefetch_data[0][19] ), .Q(\r_prefetch_data[0][19] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][18] ( .CK(clk), .D(\c_prefetch_data[0][18] ), .Q(\r_prefetch_data[0][18] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][17] ( .CK(clk), .D(\c_prefetch_data[0][17] ), .Q(\r_prefetch_data[0][17] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][16] ( .CK(clk), .D(\c_prefetch_data[0][16] ), .Q(\r_prefetch_data[0][16] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][15] ( .CK(clk), .D(\c_prefetch_data[0][15] ), .Q(\r_prefetch_data[0][15] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][14] ( .CK(clk), .D(\c_prefetch_data[0][14] ), .Q(\r_prefetch_data[0][14] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][13] ( .CK(clk), .D(\c_prefetch_data[0][13] ), .Q(\r_prefetch_data[0][13] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][12] ( .CK(clk), .D(\c_prefetch_data[0][12] ), .Q(\r_prefetch_data[0][12] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][11] ( .CK(clk), .D(\c_prefetch_data[0][11] ), .Q(\r_prefetch_data[0][11] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][10] ( .CK(clk), .D(\c_prefetch_data[0][10] ), .Q(\r_prefetch_data[0][10] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][9] ( .CK(clk), .D(\c_prefetch_data[0][9] ), .Q(\r_prefetch_data[0][9] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][8] ( .CK(clk), .D(\c_prefetch_data[0][8] ), .Q(\r_prefetch_data[0][8] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][7] ( .CK(clk), .D(\c_prefetch_data[0][7] ), .Q(\r_prefetch_data[0][7] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][6] ( .CK(clk), .D(\c_prefetch_data[0][6] ), .Q(\r_prefetch_data[0][6] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][5] ( .CK(clk), .D(\c_prefetch_data[0][5] ), .Q(\r_prefetch_data[0][5] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][4] ( .CK(clk), .D(\c_prefetch_data[0][4] ), .Q(\r_prefetch_data[0][4] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][3] ( .CK(clk), .D(\c_prefetch_data[0][3] ), .Q(\r_prefetch_data[0][3] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][2] ( .CK(clk), .D(\c_prefetch_data[0][2] ), .Q(\r_prefetch_data[0][2] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][1] ( .CK(clk), .D(\c_prefetch_data[0][1] ), .Q(\r_prefetch_data[0][1] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][0] ( .CK(clk), .D(\c_prefetch_data[0][0] ), .Q(\r_prefetch_data[0][0] ), .QN( ));
Q_FDP1 \r_mem_ren_dly_REG[2] ( .CK(clk), .R(rst_n), .D(c_mem_ren_dly[2]), .Q(r_mem_ren_dly[2]), .QN( ));
Q_FDP1 \r_mem_ren_dly_REG[1] ( .CK(clk), .R(rst_n), .D(c_mem_ren_dly[1]), .Q(r_mem_ren_dly[1]), .QN( ));
Q_FDP1 \r_mem_ren_dly_REG[0] ( .CK(clk), .R(rst_n), .D(c_mem_ren_dly[0]), .Q(r_mem_ren_dly[0]), .QN( ));
Q_FDP2 r_mem_empty_REG  ( .CK(clk), .S(rst_n), .D(c_mem_empty), .Q(r_mem_empty), .QN(n151));
Q_FDP1 r_mem_full_REG  ( .CK(clk), .R(rst_n), .D(c_mem_full), .Q(r_mem_full), .QN(n111));
Q_FDP1 \r_mem_wptr_REG[7] ( .CK(clk), .R(rst_n), .D(c_mem_wptr[7]), .Q(r_mem_wptr[7]), .QN( ));
Q_FDP1 \r_mem_wptr_REG[6] ( .CK(clk), .R(rst_n), .D(c_mem_wptr[6]), .Q(r_mem_wptr[6]), .QN(n833));
Q_FDP1 \r_mem_wptr_REG[5] ( .CK(clk), .R(rst_n), .D(c_mem_wptr[5]), .Q(r_mem_wptr[5]), .QN( ));
Q_FDP1 \r_mem_wptr_REG[4] ( .CK(clk), .R(rst_n), .D(c_mem_wptr[4]), .Q(r_mem_wptr[4]), .QN(n834));
Q_FDP1 \r_mem_wptr_REG[3] ( .CK(clk), .R(rst_n), .D(c_mem_wptr[3]), .Q(r_mem_wptr[3]), .QN(n835));
Q_FDP1 \r_mem_wptr_REG[2] ( .CK(clk), .R(rst_n), .D(c_mem_wptr[2]), .Q(r_mem_wptr[2]), .QN( ));
Q_FDP1 \r_mem_wptr_REG[1] ( .CK(clk), .R(rst_n), .D(c_mem_wptr[1]), .Q(r_mem_wptr[1]), .QN( ));
Q_FDP1 \r_mem_wptr_REG[0] ( .CK(clk), .R(rst_n), .D(c_mem_wptr[0]), .Q(r_mem_wptr[0]), .QN(n273));
Q_FDP1 \r_mem_rptr_REG[7] ( .CK(clk), .R(rst_n), .D(c_mem_rptr[7]), .Q(r_mem_rptr[7]), .QN( ));
Q_FDP1 \r_mem_rptr_REG[6] ( .CK(clk), .R(rst_n), .D(c_mem_rptr[6]), .Q(r_mem_rptr[6]), .QN(n839));
Q_FDP1 \r_mem_rptr_REG[5] ( .CK(clk), .R(rst_n), .D(c_mem_rptr[5]), .Q(r_mem_rptr[5]), .QN( ));
Q_FDP1 \r_mem_rptr_REG[4] ( .CK(clk), .R(rst_n), .D(c_mem_rptr[4]), .Q(r_mem_rptr[4]), .QN(n840));
Q_FDP1 \r_mem_rptr_REG[3] ( .CK(clk), .R(rst_n), .D(c_mem_rptr[3]), .Q(r_mem_rptr[3]), .QN(n841));
Q_FDP1 \r_mem_rptr_REG[2] ( .CK(clk), .R(rst_n), .D(c_mem_rptr[2]), .Q(r_mem_rptr[2]), .QN( ));
Q_FDP1 \r_mem_rptr_REG[1] ( .CK(clk), .R(rst_n), .D(c_mem_rptr[1]), .Q(r_mem_rptr[1]), .QN( ));
Q_FDP1 \r_mem_rptr_REG[0] ( .CK(clk), .R(rst_n), .D(c_mem_rptr[0]), .Q(r_mem_rptr[0]), .QN( ));
Q_FDP2 r_prefetch_empty_REG  ( .CK(clk), .S(rst_n), .D(c_prefetch_empty), .Q(r_prefetch_empty), .QN( ));
Q_FDP1 r_prefetch_full_REG  ( .CK(clk), .R(rst_n), .D(c_prefetch_full), .Q(r_prefetch_full), .QN( ));
Q_FDP1 \r_prefetch_wptr_REG[2] ( .CK(clk), .R(rst_n), .D(c_prefetch_wptr[2]), .Q(r_prefetch_wptr[2]), .QN( ));
Q_FDP1 \r_prefetch_wptr_REG[1] ( .CK(clk), .R(rst_n), .D(c_prefetch_wptr[1]), .Q(r_prefetch_wptr[1]), .QN( ));
Q_FDP2 \r_prefetch_wptr_REG[0] ( .CK(clk), .S(rst_n), .D(c_prefetch_wptr[0]), .Q(r_prefetch_wptr[0]), .QN( ));
Q_FDP1 \r_prefetch_rptr_REG[1] ( .CK(clk), .R(rst_n), .D(c_prefetch_rptr[1]), .Q(r_prefetch_rptr[1]), .QN( ));
Q_FDP1 \r_prefetch_rptr_REG[0] ( .CK(clk), .R(rst_n), .D(c_prefetch_rptr[0]), .Q(r_prefetch_rptr[0]), .QN(n842));
Q_FDP1 \r_prefetch_depth_REG[1] ( .CK(clk), .R(rst_n), .D(c_prefetch_depth[1]), .Q(r_prefetch_depth[1]), .QN(n192));
Q_FDP1 \r_prefetch_depth_REG[0] ( .CK(clk), .R(rst_n), .D(c_prefetch_depth[0]), .Q(r_prefetch_depth[0]), .QN(n193));
Q_FDP1 \r_used_slots_REG[7] ( .CK(clk), .R(rst_n), .D(c_used_slots[7]), .Q(r_used_slots[7]), .QN( ));
Q_FDP1 \r_used_slots_REG[6] ( .CK(clk), .R(rst_n), .D(c_used_slots[6]), .Q(r_used_slots[6]), .QN( ));
Q_FDP1 \r_used_slots_REG[5] ( .CK(clk), .R(rst_n), .D(c_used_slots[5]), .Q(r_used_slots[5]), .QN( ));
Q_FDP1 \r_used_slots_REG[4] ( .CK(clk), .R(rst_n), .D(c_used_slots[4]), .Q(r_used_slots[4]), .QN( ));
Q_FDP1 \r_used_slots_REG[3] ( .CK(clk), .R(rst_n), .D(c_used_slots[3]), .Q(r_used_slots[3]), .QN( ));
Q_FDP1 \r_used_slots_REG[2] ( .CK(clk), .R(rst_n), .D(c_used_slots[2]), .Q(r_used_slots[2]), .QN( ));
Q_FDP1 \r_used_slots_REG[1] ( .CK(clk), .R(rst_n), .D(c_used_slots[1]), .Q(r_used_slots[1]), .QN( ));
Q_FDP1 \r_used_slots_REG[0] ( .CK(clk), .R(rst_n), .D(c_used_slots[0]), .Q(r_used_slots[0]), .QN(n311));
Q_FDP2 \r_free_slots_REG[7] ( .CK(clk), .S(rst_n), .D(c_free_slots[7]), .Q(r_free_slots[7]), .QN( ));
Q_FDP1 \r_free_slots_REG[6] ( .CK(clk), .R(rst_n), .D(c_free_slots[6]), .Q(r_free_slots[6]), .QN( ));
Q_FDP2 \r_free_slots_REG[5] ( .CK(clk), .S(rst_n), .D(c_free_slots[5]), .Q(r_free_slots[5]), .QN( ));
Q_FDP1 \r_free_slots_REG[4] ( .CK(clk), .R(rst_n), .D(c_free_slots[4]), .Q(r_free_slots[4]), .QN( ));
Q_FDP2 \r_free_slots_REG[3] ( .CK(clk), .S(rst_n), .D(c_free_slots[3]), .Q(r_free_slots[3]), .QN( ));
Q_FDP1 \r_free_slots_REG[2] ( .CK(clk), .R(rst_n), .D(c_free_slots[2]), .Q(r_free_slots[2]), .QN( ));
Q_FDP2 \r_free_slots_REG[1] ( .CK(clk), .S(rst_n), .D(c_free_slots[1]), .Q(r_free_slots[1]), .QN( ));
Q_FDP2 \r_free_slots_REG[0] ( .CK(clk), .S(rst_n), .D(c_free_slots[0]), .Q(r_free_slots[0]), .QN(n324));
Q_OR02 U401 ( .A0(n151), .A1(n86), .Z(n124));
Q_AN02 U402 ( .A0(wen), .A1(n111), .Z(n147));
Q_AN02 U403 ( .A0(n147), .A1(n124), .Z(mem_wen));
Q_AN02 U404 ( .A0(ren), .A1(empty), .Z(underflow));
Q_AN02 U405 ( .A0(wen), .A1(r_mem_full), .Z(overflow));
Q_INV U406 ( .A(wen), .Z(n121));
Q_INV U407 ( .A(ren), .Z(n110));
Q_OR02 U408 ( .A0(n110), .A1(empty), .Z(n128));
Q_INV U409 ( .A(n128), .Z(n141));
Q_INV U410 ( .A(clear), .Z(n107));
Q_AN02 U411 ( .A0(n107), .A1(n112), .Z(n92));
Q_AN02 U412 ( .A0(n147), .A1(n107), .Z(n119));
Q_AN02 U413 ( .A0(n128), .A1(n119), .Z(n113));
Q_NR02 U414 ( .A0(n113), .A1(clear), .Z(n114));
Q_NR02 U415 ( .A0(n147), .A1(clear), .Z(n115));
Q_AO21 U416 ( .A0(n141), .A1(n115), .B0(clear), .Z(n116));
Q_INV U417 ( .A(n116), .Z(n93));
Q_INV U418 ( .A(n86), .Z(n152));
Q_NR02 U419 ( .A0(n147), .A1(n86), .Z(n118));
Q_AO21 U420 ( .A0(n118), .A1(n117), .B0(clear), .Z(n94));
Q_AN02 U421 ( .A0(n124), .A1(n119), .Z(n108));
Q_NR02 U422 ( .A0(n108), .A1(n94), .Z(n120));
Q_OR03 U423 ( .A0(n88), .A1(r_mem_full), .A2(n121), .Z(n123));
Q_INV U424 ( .A(n124), .Z(n148));
Q_AN02 U425 ( .A0(n123), .A1(n86), .Z(n122));
Q_OA21 U426 ( .A0(n148), .A1(n122), .B0(n107), .Z(n95));
Q_INV U427 ( .A(n123), .Z(n125));
Q_AN03 U428 ( .A0(n107), .A1(n124), .A2(n125), .Z(n96));
Q_OR02 U429 ( .A0(n151), .A1(n147), .Z(n142));
Q_NR02 U430 ( .A0(n86), .A1(clear), .Z(n145));
Q_AN02 U431 ( .A0(n145), .A1(n142), .Z(n97));
Q_OR02 U432 ( .A0(n97), .A1(clear), .Z(n126));
Q_INV U433 ( .A(n126), .Z(n98));
Q_NR02 U434 ( .A0(n91), .A1(clear), .Z(n127));
Q_AN02 U435 ( .A0(n141), .A1(n127), .Z(n99));
Q_AN02 U436 ( .A0(n107), .A1(n128), .Z(n100));
Q_INV U437 ( .A(n142), .Z(n129));
Q_OR02 U438 ( .A0(n86), .A1(n129), .Z(n150));
Q_OA21 U439 ( .A0(n110), .A1(empty), .B0(n142), .Z(n140));
Q_AN02 U440 ( .A0(n150), .A1(n141), .Z(n131));
Q_AN02 U441 ( .A0(n140), .A1(n152), .Z(n130));
Q_OA21 U442 ( .A0(n131), .A1(n130), .B0(n107), .Z(n101));
Q_AN02 U443 ( .A0(n140), .A1(n145), .Z(n132));
Q_NR02 U444 ( .A0(n132), .A1(clear), .Z(n133));
Q_AN03 U445 ( .A0(n192), .A1(r_prefetch_depth[0]), .A2(n141), .Z(n134));
Q_AO21 U446 ( .A0(n150), .A1(n134), .B0(clear), .Z(n102));
Q_NR02 U447 ( .A0(n97), .A1(n102), .Z(n135));
Q_NR02 U448 ( .A0(r_prefetch_depth[0]), .A1(n86), .Z(n136));
Q_AN02 U449 ( .A0(r_prefetch_depth[1]), .A1(n107), .Z(n137));
Q_AN03 U450 ( .A0(n137), .A1(n136), .A2(n140), .Z(n138));
Q_NR02 U451 ( .A0(n138), .A1(clear), .Z(n139));
Q_AN03 U452 ( .A0(r_prefetch_depth[1]), .A1(n193), .A2(n140), .Z(n144));
Q_AN02 U453 ( .A0(n142), .A1(n141), .Z(n143));
Q_OA21 U454 ( .A0(n144), .A1(n143), .B0(n145), .Z(n106));
Q_NR02 U455 ( .A0(n108), .A1(clear), .Z(n146));
Q_AN02 U456 ( .A0(n148), .A1(n147), .Z(n109));
Q_ND02 U457 ( .A0(ren), .A1(n87), .Z(n149));
Q_INV U458 ( .A(n150), .Z(prefetch_wen));
Q_NR02 U459 ( .A0(n86), .A1(r_mem_empty), .Z(mem_ren));
Q_AN02 U460 ( .A0(n107), .A1(r_mem_ren_dly[1]), .Z(c_mem_ren_dly[2]));
Q_AN02 U461 ( .A0(n107), .A1(r_mem_ren_dly[0]), .Z(c_mem_ren_dly[1]));
Q_AN02 U462 ( .A0(n107), .A1(mem_ren), .Z(c_mem_ren_dly[0]));
Q_MX02 U463 ( .S(n87), .A0(n2), .A1(mem_ecc_error), .Z(rerr));
Q_MX02 U464 ( .S(n87), .A0(n3), .A1(mem_rdata[82]), .Z(rdata[82]));
Q_MX02 U465 ( .S(n87), .A0(n4), .A1(mem_rdata[81]), .Z(rdata[81]));
Q_MX02 U466 ( .S(n87), .A0(n5), .A1(mem_rdata[80]), .Z(rdata[80]));
Q_MX02 U467 ( .S(n87), .A0(n6), .A1(mem_rdata[79]), .Z(rdata[79]));
Q_MX02 U468 ( .S(n87), .A0(n7), .A1(mem_rdata[78]), .Z(rdata[78]));
Q_MX02 U469 ( .S(n87), .A0(n8), .A1(mem_rdata[77]), .Z(rdata[77]));
Q_MX02 U470 ( .S(n87), .A0(n9), .A1(mem_rdata[76]), .Z(rdata[76]));
Q_MX02 U471 ( .S(n87), .A0(n10), .A1(mem_rdata[75]), .Z(rdata[75]));
Q_MX02 U472 ( .S(n87), .A0(n11), .A1(mem_rdata[74]), .Z(rdata[74]));
Q_MX02 U473 ( .S(n87), .A0(n12), .A1(mem_rdata[73]), .Z(rdata[73]));
Q_MX02 U474 ( .S(n87), .A0(n13), .A1(mem_rdata[72]), .Z(rdata[72]));
Q_MX02 U475 ( .S(n87), .A0(n14), .A1(mem_rdata[71]), .Z(rdata[71]));
Q_MX02 U476 ( .S(n87), .A0(n15), .A1(mem_rdata[70]), .Z(rdata[70]));
Q_MX02 U477 ( .S(n87), .A0(n16), .A1(mem_rdata[69]), .Z(rdata[69]));
Q_MX02 U478 ( .S(n87), .A0(n17), .A1(mem_rdata[68]), .Z(rdata[68]));
Q_MX02 U479 ( .S(n87), .A0(n18), .A1(mem_rdata[67]), .Z(rdata[67]));
Q_MX02 U480 ( .S(n87), .A0(n19), .A1(mem_rdata[66]), .Z(rdata[66]));
Q_MX02 U481 ( .S(n87), .A0(n20), .A1(mem_rdata[65]), .Z(rdata[65]));
Q_MX02 U482 ( .S(n87), .A0(n21), .A1(mem_rdata[64]), .Z(rdata[64]));
Q_MX02 U483 ( .S(n87), .A0(n22), .A1(mem_rdata[63]), .Z(rdata[63]));
Q_MX02 U484 ( .S(n87), .A0(n23), .A1(mem_rdata[62]), .Z(rdata[62]));
Q_MX02 U485 ( .S(n87), .A0(n24), .A1(mem_rdata[61]), .Z(rdata[61]));
Q_MX02 U486 ( .S(n87), .A0(n25), .A1(mem_rdata[60]), .Z(rdata[60]));
Q_MX02 U487 ( .S(n87), .A0(n26), .A1(mem_rdata[59]), .Z(rdata[59]));
Q_MX02 U488 ( .S(n87), .A0(n27), .A1(mem_rdata[58]), .Z(rdata[58]));
Q_MX02 U489 ( .S(n87), .A0(n28), .A1(mem_rdata[57]), .Z(rdata[57]));
Q_MX02 U490 ( .S(n87), .A0(n29), .A1(mem_rdata[56]), .Z(rdata[56]));
Q_MX02 U491 ( .S(n87), .A0(n30), .A1(mem_rdata[55]), .Z(rdata[55]));
Q_MX02 U492 ( .S(n87), .A0(n31), .A1(mem_rdata[54]), .Z(rdata[54]));
Q_MX02 U493 ( .S(n87), .A0(n32), .A1(mem_rdata[53]), .Z(rdata[53]));
Q_MX02 U494 ( .S(n87), .A0(n33), .A1(mem_rdata[52]), .Z(rdata[52]));
Q_MX02 U495 ( .S(n87), .A0(n34), .A1(mem_rdata[51]), .Z(rdata[51]));
Q_MX02 U496 ( .S(n87), .A0(n35), .A1(mem_rdata[50]), .Z(rdata[50]));
Q_MX02 U497 ( .S(n87), .A0(n36), .A1(mem_rdata[49]), .Z(rdata[49]));
Q_MX02 U498 ( .S(n87), .A0(n37), .A1(mem_rdata[48]), .Z(rdata[48]));
Q_MX02 U499 ( .S(n87), .A0(n38), .A1(mem_rdata[47]), .Z(rdata[47]));
Q_MX02 U500 ( .S(n87), .A0(n39), .A1(mem_rdata[46]), .Z(rdata[46]));
Q_MX02 U501 ( .S(n87), .A0(n40), .A1(mem_rdata[45]), .Z(rdata[45]));
Q_MX02 U502 ( .S(n87), .A0(n41), .A1(mem_rdata[44]), .Z(rdata[44]));
Q_MX02 U503 ( .S(n87), .A0(n42), .A1(mem_rdata[43]), .Z(rdata[43]));
Q_MX02 U504 ( .S(n87), .A0(n43), .A1(mem_rdata[42]), .Z(rdata[42]));
Q_MX02 U505 ( .S(n87), .A0(n44), .A1(mem_rdata[41]), .Z(rdata[41]));
Q_MX02 U506 ( .S(n87), .A0(n45), .A1(mem_rdata[40]), .Z(rdata[40]));
Q_MX02 U507 ( .S(n87), .A0(n46), .A1(mem_rdata[39]), .Z(rdata[39]));
Q_MX02 U508 ( .S(n87), .A0(n47), .A1(mem_rdata[38]), .Z(rdata[38]));
Q_MX02 U509 ( .S(n87), .A0(n48), .A1(mem_rdata[37]), .Z(rdata[37]));
Q_MX02 U510 ( .S(n87), .A0(n49), .A1(mem_rdata[36]), .Z(rdata[36]));
Q_MX02 U511 ( .S(n87), .A0(n50), .A1(mem_rdata[35]), .Z(rdata[35]));
Q_MX02 U512 ( .S(n87), .A0(n51), .A1(mem_rdata[34]), .Z(rdata[34]));
Q_MX02 U513 ( .S(n87), .A0(n52), .A1(mem_rdata[33]), .Z(rdata[33]));
Q_MX02 U514 ( .S(n87), .A0(n53), .A1(mem_rdata[32]), .Z(rdata[32]));
Q_MX02 U515 ( .S(n87), .A0(n54), .A1(mem_rdata[31]), .Z(rdata[31]));
Q_MX02 U516 ( .S(n87), .A0(n55), .A1(mem_rdata[30]), .Z(rdata[30]));
Q_MX02 U517 ( .S(n87), .A0(n56), .A1(mem_rdata[29]), .Z(rdata[29]));
Q_MX02 U518 ( .S(n87), .A0(n57), .A1(mem_rdata[28]), .Z(rdata[28]));
Q_MX02 U519 ( .S(n87), .A0(n58), .A1(mem_rdata[27]), .Z(rdata[27]));
Q_MX02 U520 ( .S(n87), .A0(n59), .A1(mem_rdata[26]), .Z(rdata[26]));
Q_MX02 U521 ( .S(n87), .A0(n60), .A1(mem_rdata[25]), .Z(rdata[25]));
Q_MX02 U522 ( .S(n87), .A0(n61), .A1(mem_rdata[24]), .Z(rdata[24]));
Q_MX02 U523 ( .S(n87), .A0(n62), .A1(mem_rdata[23]), .Z(rdata[23]));
Q_MX02 U524 ( .S(n87), .A0(n63), .A1(mem_rdata[22]), .Z(rdata[22]));
Q_MX02 U525 ( .S(n87), .A0(n64), .A1(mem_rdata[21]), .Z(rdata[21]));
Q_MX02 U526 ( .S(n87), .A0(n65), .A1(mem_rdata[20]), .Z(rdata[20]));
Q_MX02 U527 ( .S(n87), .A0(n66), .A1(mem_rdata[19]), .Z(rdata[19]));
Q_MX02 U528 ( .S(n87), .A0(n67), .A1(mem_rdata[18]), .Z(rdata[18]));
Q_MX02 U529 ( .S(n87), .A0(n68), .A1(mem_rdata[17]), .Z(rdata[17]));
Q_MX02 U530 ( .S(n87), .A0(n69), .A1(mem_rdata[16]), .Z(rdata[16]));
Q_MX02 U531 ( .S(n87), .A0(n70), .A1(mem_rdata[15]), .Z(rdata[15]));
Q_MX02 U532 ( .S(n87), .A0(n71), .A1(mem_rdata[14]), .Z(rdata[14]));
Q_MX02 U533 ( .S(n87), .A0(n72), .A1(mem_rdata[13]), .Z(rdata[13]));
Q_MX02 U534 ( .S(n87), .A0(n73), .A1(mem_rdata[12]), .Z(rdata[12]));
Q_MX02 U535 ( .S(n87), .A0(n74), .A1(mem_rdata[11]), .Z(rdata[11]));
Q_MX02 U536 ( .S(n87), .A0(n75), .A1(mem_rdata[10]), .Z(rdata[10]));
Q_MX02 U537 ( .S(n87), .A0(n76), .A1(mem_rdata[9]), .Z(rdata[9]));
Q_MX02 U538 ( .S(n87), .A0(n77), .A1(mem_rdata[8]), .Z(rdata[8]));
Q_MX02 U539 ( .S(n87), .A0(n78), .A1(mem_rdata[7]), .Z(rdata[7]));
Q_MX02 U540 ( .S(n87), .A0(n79), .A1(mem_rdata[6]), .Z(rdata[6]));
Q_MX02 U541 ( .S(n87), .A0(n80), .A1(mem_rdata[5]), .Z(rdata[5]));
Q_MX02 U542 ( .S(n87), .A0(n81), .A1(mem_rdata[4]), .Z(rdata[4]));
Q_MX02 U543 ( .S(n87), .A0(n82), .A1(mem_rdata[3]), .Z(rdata[3]));
Q_MX02 U544 ( .S(n87), .A0(n83), .A1(mem_rdata[2]), .Z(rdata[2]));
Q_MX02 U545 ( .S(n87), .A0(n84), .A1(mem_rdata[1]), .Z(rdata[1]));
Q_MX02 U546 ( .S(n87), .A0(n85), .A1(mem_rdata[0]), .Z(rdata[0]));
Q_MX02 U547 ( .S(n92), .A0(n153), .A1(n154), .Z(c_used_slots[7]));
Q_AN02 U548 ( .A0(n114), .A1(r_used_slots[7]), .Z(n153));
Q_MX02 U549 ( .S(n114), .A0(n299), .A1(n286), .Z(n154));
Q_MX02 U550 ( .S(n92), .A0(n155), .A1(n156), .Z(c_used_slots[6]));
Q_AN02 U551 ( .A0(n114), .A1(r_used_slots[6]), .Z(n155));
Q_MX02 U552 ( .S(n114), .A0(n301), .A1(n288), .Z(n156));
Q_MX02 U553 ( .S(n92), .A0(n157), .A1(n158), .Z(c_used_slots[5]));
Q_AN02 U554 ( .A0(n114), .A1(r_used_slots[5]), .Z(n157));
Q_MX02 U555 ( .S(n114), .A0(n303), .A1(n290), .Z(n158));
Q_MX02 U556 ( .S(n92), .A0(n159), .A1(n160), .Z(c_used_slots[4]));
Q_AN02 U557 ( .A0(n114), .A1(r_used_slots[4]), .Z(n159));
Q_MX02 U558 ( .S(n114), .A0(n305), .A1(n292), .Z(n160));
Q_MX02 U559 ( .S(n92), .A0(n161), .A1(n162), .Z(c_used_slots[3]));
Q_AN02 U560 ( .A0(n114), .A1(r_used_slots[3]), .Z(n161));
Q_MX02 U561 ( .S(n114), .A0(n307), .A1(n294), .Z(n162));
Q_MX02 U562 ( .S(n92), .A0(n163), .A1(n164), .Z(c_used_slots[2]));
Q_AN02 U563 ( .A0(n114), .A1(r_used_slots[2]), .Z(n163));
Q_MX02 U564 ( .S(n114), .A0(n309), .A1(n296), .Z(n164));
Q_MX02 U565 ( .S(n92), .A0(n165), .A1(n166), .Z(c_used_slots[1]));
Q_AN02 U566 ( .A0(n114), .A1(r_used_slots[1]), .Z(n165));
Q_MX02 U567 ( .S(n92), .A0(n167), .A1(n311), .Z(c_used_slots[0]));
Q_AN02 U568 ( .A0(n114), .A1(r_used_slots[0]), .Z(n167));
Q_MX02 U569 ( .S(n92), .A0(n168), .A1(n169), .Z(c_free_slots[7]));
Q_OR02 U570 ( .A0(n116), .A1(r_free_slots[7]), .Z(n168));
Q_MX02 U571 ( .S(n116), .A0(n274), .A1(n312), .Z(n169));
Q_MX02 U572 ( .S(n92), .A0(n170), .A1(n171), .Z(c_free_slots[6]));
Q_AN02 U573 ( .A0(n93), .A1(r_free_slots[6]), .Z(n170));
Q_MX02 U574 ( .S(n116), .A0(n276), .A1(n314), .Z(n171));
Q_MX02 U575 ( .S(n92), .A0(n172), .A1(n173), .Z(c_free_slots[5]));
Q_OR02 U576 ( .A0(n116), .A1(r_free_slots[5]), .Z(n172));
Q_MX02 U577 ( .S(n116), .A0(n278), .A1(n316), .Z(n173));
Q_MX02 U578 ( .S(n92), .A0(n174), .A1(n175), .Z(c_free_slots[4]));
Q_AN02 U579 ( .A0(n93), .A1(r_free_slots[4]), .Z(n174));
Q_MX02 U580 ( .S(n116), .A0(n280), .A1(n318), .Z(n175));
Q_MX02 U581 ( .S(n92), .A0(n176), .A1(n177), .Z(c_free_slots[3]));
Q_OR02 U582 ( .A0(n116), .A1(r_free_slots[3]), .Z(n176));
Q_MX02 U583 ( .S(n116), .A0(n282), .A1(n320), .Z(n177));
Q_MX02 U584 ( .S(n92), .A0(n178), .A1(n179), .Z(c_free_slots[2]));
Q_AN02 U585 ( .A0(n93), .A1(r_free_slots[2]), .Z(n178));
Q_MX02 U586 ( .S(n116), .A0(n284), .A1(n322), .Z(n179));
Q_MX02 U587 ( .S(n92), .A0(n180), .A1(n181), .Z(c_free_slots[1]));
Q_OR02 U588 ( .A0(n116), .A1(r_free_slots[1]), .Z(n180));
Q_MX02 U589 ( .S(n92), .A0(n182), .A1(n324), .Z(c_free_slots[0]));
Q_OR02 U590 ( .A0(n116), .A1(r_free_slots[0]), .Z(n182));
Q_MX02 U591 ( .S(n120), .A0(n94), .A1(r_mem_empty), .Z(c_mem_empty));
Q_MX02 U592 ( .S(n95), .A0(n96), .A1(r_mem_full), .Z(c_mem_full));
Q_MX02 U593 ( .S(n97), .A0(n183), .A1(\c_mem_prefetch_wptr_dly[0][1] ), .Z(c_prefetch_wptr[2]));
Q_AN02 U594 ( .A0(n98), .A1(\c_mem_prefetch_wptr_dly[0][2] ), .Z(n183));
Q_MX02 U595 ( .S(n97), .A0(n184), .A1(\c_mem_prefetch_wptr_dly[0][0] ), .Z(c_prefetch_wptr[1]));
Q_AN02 U596 ( .A0(n98), .A1(\c_mem_prefetch_wptr_dly[0][1] ), .Z(n184));
Q_MX02 U597 ( .S(n97), .A0(n185), .A1(\c_mem_prefetch_wptr_dly[0][2] ), .Z(c_prefetch_wptr[0]));
Q_OR02 U598 ( .A0(n126), .A1(\c_mem_prefetch_wptr_dly[0][0] ), .Z(n185));
Q_MX02 U599 ( .S(n99), .A0(n186), .A1(n194), .Z(c_prefetch_rptr[1]));
Q_AN02 U600 ( .A0(n100), .A1(r_prefetch_rptr[1]), .Z(n186));
Q_MX02 U601 ( .S(n99), .A0(n187), .A1(n842), .Z(c_prefetch_rptr[0]));
Q_AN02 U602 ( .A0(n100), .A1(r_prefetch_rptr[0]), .Z(n187));
Q_MX02 U603 ( .S(n101), .A0(n188), .A1(n189), .Z(c_prefetch_depth[1]));
Q_AN02 U604 ( .A0(n133), .A1(r_prefetch_depth[1]), .Z(n188));
Q_MX02 U605 ( .S(n101), .A0(n190), .A1(n193), .Z(c_prefetch_depth[0]));
Q_AN02 U606 ( .A0(n133), .A1(r_prefetch_depth[0]), .Z(n190));
Q_MX02 U607 ( .S(n135), .A0(n102), .A1(r_prefetch_empty), .Z(c_prefetch_empty));
Q_XOR2 U608 ( .A0(r_prefetch_depth[0]), .A1(n192), .Z(n191));
Q_XOR2 U609 ( .A0(r_prefetch_rptr[1]), .A1(r_prefetch_rptr[0]), .Z(n194));
Q_AN02 U610 ( .A0(n107), .A1(n206), .Z(c_mem_rptr[7]));
Q_AN02 U611 ( .A0(n107), .A1(n207), .Z(c_mem_rptr[6]));
Q_AN02 U612 ( .A0(n107), .A1(n208), .Z(c_mem_rptr[5]));
Q_AN02 U613 ( .A0(n107), .A1(n209), .Z(c_mem_rptr[4]));
Q_AN02 U614 ( .A0(n107), .A1(n210), .Z(c_mem_rptr[3]));
Q_AN02 U615 ( .A0(n107), .A1(n211), .Z(c_mem_rptr[2]));
Q_AN02 U616 ( .A0(n107), .A1(n212), .Z(c_mem_rptr[1]));
Q_AN02 U617 ( .A0(n107), .A1(n213), .Z(c_mem_rptr[0]));
Q_ND02 U618 ( .A0(n196), .A1(n195), .Z(n88));
Q_AN03 U619 ( .A0(n199), .A1(n198), .A2(n197), .Z(n195));
Q_AN03 U620 ( .A0(n202), .A1(n201), .A2(n200), .Z(n196));
Q_AN03 U621 ( .A0(n205), .A1(n204), .A2(n203), .Z(n197));
Q_XNR2 U622 ( .A0(n253), .A1(n206), .Z(n198));
Q_XNR2 U623 ( .A0(n254), .A1(n207), .Z(n199));
Q_XNR2 U624 ( .A0(n255), .A1(n208), .Z(n200));
Q_XNR2 U625 ( .A0(n256), .A1(n209), .Z(n201));
Q_XNR2 U626 ( .A0(n257), .A1(n210), .Z(n202));
Q_XNR2 U627 ( .A0(n258), .A1(n211), .Z(n203));
Q_XNR2 U628 ( .A0(n259), .A1(n212), .Z(n204));
Q_XNR2 U629 ( .A0(n273), .A1(n213), .Z(n205));
Q_MX02 U630 ( .S(mem_ren), .A0(r_mem_rptr[7]), .A1(n225), .Z(n206));
Q_MX02 U631 ( .S(mem_ren), .A0(r_mem_rptr[6]), .A1(n226), .Z(n207));
Q_MX02 U632 ( .S(mem_ren), .A0(r_mem_rptr[5]), .A1(n227), .Z(n208));
Q_MX02 U633 ( .S(mem_ren), .A0(r_mem_rptr[4]), .A1(n228), .Z(n209));
Q_MX02 U634 ( .S(mem_ren), .A0(r_mem_rptr[3]), .A1(n229), .Z(n210));
Q_MX02 U635 ( .S(mem_ren), .A0(r_mem_rptr[2]), .A1(n230), .Z(n211));
Q_MX02 U636 ( .S(mem_ren), .A0(r_mem_rptr[1]), .A1(n231), .Z(n212));
Q_AN03 U637 ( .A0(n215), .A1(n214), .A2(n151), .Z(n117));
Q_AN03 U638 ( .A0(n218), .A1(n217), .A2(n216), .Z(n214));
Q_AN03 U639 ( .A0(n221), .A1(n220), .A2(n219), .Z(n215));
Q_AN03 U640 ( .A0(n224), .A1(n223), .A2(n222), .Z(n216));
Q_XNR2 U641 ( .A0(n225), .A1(r_mem_wptr[7]), .Z(n217));
Q_XNR2 U642 ( .A0(n226), .A1(r_mem_wptr[6]), .Z(n218));
Q_XNR2 U643 ( .A0(n227), .A1(r_mem_wptr[5]), .Z(n219));
Q_XNR2 U644 ( .A0(n228), .A1(r_mem_wptr[4]), .Z(n220));
Q_XNR2 U645 ( .A0(n229), .A1(r_mem_wptr[3]), .Z(n221));
Q_XNR2 U646 ( .A0(n230), .A1(r_mem_wptr[2]), .Z(n222));
Q_XNR2 U647 ( .A0(n231), .A1(r_mem_wptr[1]), .Z(n223));
Q_XOR2 U648 ( .A0(r_mem_rptr[0]), .A1(r_mem_wptr[0]), .Z(n224));
Q_AN02 U649 ( .A0(n90), .A1(n232), .Z(n225));
Q_AN02 U650 ( .A0(n90), .A1(n234), .Z(n226));
Q_AN02 U651 ( .A0(n90), .A1(n236), .Z(n227));
Q_AN02 U652 ( .A0(n90), .A1(n238), .Z(n228));
Q_AN02 U653 ( .A0(n90), .A1(n240), .Z(n229));
Q_AN02 U654 ( .A0(n90), .A1(n242), .Z(n230));
Q_AN02 U655 ( .A0(n90), .A1(n244), .Z(n231));
Q_XOR2 U656 ( .A0(r_mem_rptr[7]), .A1(n233), .Z(n232));
Q_AD01HF U657 ( .A0(r_mem_rptr[6]), .B0(n235), .S(n234), .CO(n233));
Q_AD01HF U658 ( .A0(r_mem_rptr[5]), .B0(n237), .S(n236), .CO(n235));
Q_AD01HF U659 ( .A0(r_mem_rptr[4]), .B0(n239), .S(n238), .CO(n237));
Q_AD01HF U660 ( .A0(r_mem_rptr[3]), .B0(n241), .S(n240), .CO(n239));
Q_AD01HF U661 ( .A0(r_mem_rptr[2]), .B0(n243), .S(n242), .CO(n241));
Q_AD01HF U662 ( .A0(r_mem_rptr[1]), .B0(r_mem_rptr[0]), .S(n244), .CO(n243));
Q_MX02 U663 ( .S(n108), .A0(n245), .A1(n253), .Z(c_mem_wptr[7]));
Q_AN02 U664 ( .A0(n146), .A1(r_mem_wptr[7]), .Z(n245));
Q_MX02 U665 ( .S(n108), .A0(n246), .A1(n254), .Z(c_mem_wptr[6]));
Q_AN02 U666 ( .A0(n146), .A1(r_mem_wptr[6]), .Z(n246));
Q_MX02 U667 ( .S(n108), .A0(n247), .A1(n255), .Z(c_mem_wptr[5]));
Q_AN02 U668 ( .A0(n146), .A1(r_mem_wptr[5]), .Z(n247));
Q_MX02 U669 ( .S(n108), .A0(n248), .A1(n256), .Z(c_mem_wptr[4]));
Q_AN02 U670 ( .A0(n146), .A1(r_mem_wptr[4]), .Z(n248));
Q_MX02 U671 ( .S(n108), .A0(n249), .A1(n257), .Z(c_mem_wptr[3]));
Q_AN02 U672 ( .A0(n146), .A1(r_mem_wptr[3]), .Z(n249));
Q_MX02 U673 ( .S(n108), .A0(n250), .A1(n258), .Z(c_mem_wptr[2]));
Q_AN02 U674 ( .A0(n146), .A1(r_mem_wptr[2]), .Z(n250));
Q_MX02 U675 ( .S(n108), .A0(n251), .A1(n259), .Z(c_mem_wptr[1]));
Q_AN02 U676 ( .A0(n146), .A1(r_mem_wptr[1]), .Z(n251));
Q_MX02 U677 ( .S(n108), .A0(n252), .A1(n273), .Z(c_mem_wptr[0]));
Q_AN02 U678 ( .A0(n146), .A1(r_mem_wptr[0]), .Z(n252));
Q_AN02 U679 ( .A0(n89), .A1(n260), .Z(n253));
Q_AN02 U680 ( .A0(n89), .A1(n262), .Z(n254));
Q_AN02 U681 ( .A0(n89), .A1(n264), .Z(n255));
Q_AN02 U682 ( .A0(n89), .A1(n266), .Z(n256));
Q_AN02 U683 ( .A0(n89), .A1(n268), .Z(n257));
Q_AN02 U684 ( .A0(n89), .A1(n270), .Z(n258));
Q_AN02 U685 ( .A0(n89), .A1(n272), .Z(n259));
Q_XOR2 U686 ( .A0(r_mem_wptr[7]), .A1(n261), .Z(n260));
Q_AD01HF U687 ( .A0(r_mem_wptr[6]), .B0(n263), .S(n262), .CO(n261));
Q_AD01HF U688 ( .A0(r_mem_wptr[5]), .B0(n265), .S(n264), .CO(n263));
Q_AD01HF U689 ( .A0(r_mem_wptr[4]), .B0(n267), .S(n266), .CO(n265));
Q_AD01HF U690 ( .A0(r_mem_wptr[3]), .B0(n269), .S(n268), .CO(n267));
Q_AD01HF U691 ( .A0(r_mem_wptr[2]), .B0(n271), .S(n270), .CO(n269));
Q_AD01HF U692 ( .A0(r_mem_wptr[1]), .B0(r_mem_wptr[0]), .S(n272), .CO(n271));
Q_XNR2 U693 ( .A0(r_free_slots[7]), .A1(n275), .Z(n274));
Q_OR02 U694 ( .A0(r_free_slots[6]), .A1(n277), .Z(n275));
Q_XNR2 U695 ( .A0(r_free_slots[6]), .A1(n277), .Z(n276));
Q_OR02 U696 ( .A0(r_free_slots[5]), .A1(n279), .Z(n277));
Q_XNR2 U697 ( .A0(r_free_slots[5]), .A1(n279), .Z(n278));
Q_OR02 U698 ( .A0(r_free_slots[4]), .A1(n281), .Z(n279));
Q_XNR2 U699 ( .A0(r_free_slots[4]), .A1(n281), .Z(n280));
Q_OR02 U700 ( .A0(r_free_slots[3]), .A1(n283), .Z(n281));
Q_XNR2 U701 ( .A0(r_free_slots[3]), .A1(n283), .Z(n282));
Q_OR02 U702 ( .A0(r_free_slots[2]), .A1(n285), .Z(n283));
Q_XNR2 U703 ( .A0(r_free_slots[2]), .A1(n285), .Z(n284));
Q_OR02 U704 ( .A0(r_free_slots[1]), .A1(r_free_slots[0]), .Z(n285));
Q_XNR3 U705 ( .A0(r_free_slots[1]), .A1(r_free_slots[0]), .A2(n116), .Z(n181));
Q_XNR2 U706 ( .A0(r_used_slots[7]), .A1(n287), .Z(n286));
Q_OR02 U707 ( .A0(r_used_slots[6]), .A1(n289), .Z(n287));
Q_XNR2 U708 ( .A0(r_used_slots[6]), .A1(n289), .Z(n288));
Q_OR02 U709 ( .A0(r_used_slots[5]), .A1(n291), .Z(n289));
Q_XNR2 U710 ( .A0(r_used_slots[5]), .A1(n291), .Z(n290));
Q_OR02 U711 ( .A0(r_used_slots[4]), .A1(n293), .Z(n291));
Q_XNR2 U712 ( .A0(r_used_slots[4]), .A1(n293), .Z(n292));
Q_OR02 U713 ( .A0(r_used_slots[3]), .A1(n295), .Z(n293));
Q_XNR2 U714 ( .A0(r_used_slots[3]), .A1(n295), .Z(n294));
Q_OR02 U715 ( .A0(r_used_slots[2]), .A1(n297), .Z(n295));
Q_XNR2 U716 ( .A0(r_used_slots[2]), .A1(n297), .Z(n296));
Q_OR02 U717 ( .A0(r_used_slots[1]), .A1(r_used_slots[0]), .Z(n297));
Q_XNR2 U718 ( .A0(r_used_slots[1]), .A1(r_used_slots[0]), .Z(n298));
Q_XOR2 U719 ( .A0(r_used_slots[7]), .A1(n300), .Z(n299));
Q_AD01HF U720 ( .A0(r_used_slots[6]), .B0(n302), .S(n301), .CO(n300));
Q_AD01HF U721 ( .A0(r_used_slots[5]), .B0(n304), .S(n303), .CO(n302));
Q_AD01HF U722 ( .A0(r_used_slots[4]), .B0(n306), .S(n305), .CO(n304));
Q_AD01HF U723 ( .A0(r_used_slots[3]), .B0(n308), .S(n307), .CO(n306));
Q_AD01HF U724 ( .A0(r_used_slots[2]), .B0(n310), .S(n309), .CO(n308));
Q_XOR2 U725 ( .A0(r_free_slots[7]), .A1(n313), .Z(n312));
Q_AD01HF U726 ( .A0(r_free_slots[6]), .B0(n315), .S(n314), .CO(n313));
Q_AD01HF U727 ( .A0(r_free_slots[5]), .B0(n317), .S(n316), .CO(n315));
Q_AD01HF U728 ( .A0(r_free_slots[4]), .B0(n319), .S(n318), .CO(n317));
Q_AD01HF U729 ( .A0(r_free_slots[3]), .B0(n321), .S(n320), .CO(n319));
Q_AD01HF U730 ( .A0(r_free_slots[2]), .B0(n323), .S(n322), .CO(n321));
Q_MX02 U731 ( .S(n103), .A0(\r_prefetch_data[0][83] ), .A1(n743), .Z(\c_prefetch_data[0][83] ));
Q_MX02 U732 ( .S(n103), .A0(\r_prefetch_data[0][82] ), .A1(n660), .Z(\c_prefetch_data[0][82] ));
Q_MX02 U733 ( .S(n103), .A0(\r_prefetch_data[0][81] ), .A1(n661), .Z(\c_prefetch_data[0][81] ));
Q_MX02 U734 ( .S(n103), .A0(\r_prefetch_data[0][80] ), .A1(n662), .Z(\c_prefetch_data[0][80] ));
Q_MX02 U735 ( .S(n103), .A0(\r_prefetch_data[0][79] ), .A1(n663), .Z(\c_prefetch_data[0][79] ));
Q_MX02 U736 ( .S(n103), .A0(\r_prefetch_data[0][78] ), .A1(n664), .Z(\c_prefetch_data[0][78] ));
Q_MX02 U737 ( .S(n103), .A0(\r_prefetch_data[0][77] ), .A1(n665), .Z(\c_prefetch_data[0][77] ));
Q_MX02 U738 ( .S(n103), .A0(\r_prefetch_data[0][76] ), .A1(n666), .Z(\c_prefetch_data[0][76] ));
Q_MX02 U739 ( .S(n103), .A0(\r_prefetch_data[0][75] ), .A1(n667), .Z(\c_prefetch_data[0][75] ));
Q_MX02 U740 ( .S(n103), .A0(\r_prefetch_data[0][74] ), .A1(n668), .Z(\c_prefetch_data[0][74] ));
Q_MX02 U741 ( .S(n103), .A0(\r_prefetch_data[0][73] ), .A1(n669), .Z(\c_prefetch_data[0][73] ));
Q_MX02 U742 ( .S(n103), .A0(\r_prefetch_data[0][72] ), .A1(n670), .Z(\c_prefetch_data[0][72] ));
Q_MX02 U743 ( .S(n103), .A0(\r_prefetch_data[0][71] ), .A1(n671), .Z(\c_prefetch_data[0][71] ));
Q_MX02 U744 ( .S(n103), .A0(\r_prefetch_data[0][70] ), .A1(n672), .Z(\c_prefetch_data[0][70] ));
Q_MX02 U745 ( .S(n103), .A0(\r_prefetch_data[0][69] ), .A1(n673), .Z(\c_prefetch_data[0][69] ));
Q_MX02 U746 ( .S(n103), .A0(\r_prefetch_data[0][68] ), .A1(n674), .Z(\c_prefetch_data[0][68] ));
Q_MX02 U747 ( .S(n103), .A0(\r_prefetch_data[0][67] ), .A1(n675), .Z(\c_prefetch_data[0][67] ));
Q_MX02 U748 ( .S(n103), .A0(\r_prefetch_data[0][66] ), .A1(n676), .Z(\c_prefetch_data[0][66] ));
Q_MX02 U749 ( .S(n103), .A0(\r_prefetch_data[0][65] ), .A1(n677), .Z(\c_prefetch_data[0][65] ));
Q_MX02 U750 ( .S(n103), .A0(\r_prefetch_data[0][64] ), .A1(n678), .Z(\c_prefetch_data[0][64] ));
Q_MX02 U751 ( .S(n103), .A0(\r_prefetch_data[0][63] ), .A1(n679), .Z(\c_prefetch_data[0][63] ));
Q_MX02 U752 ( .S(n103), .A0(\r_prefetch_data[0][62] ), .A1(n680), .Z(\c_prefetch_data[0][62] ));
Q_MX02 U753 ( .S(n103), .A0(\r_prefetch_data[0][61] ), .A1(n681), .Z(\c_prefetch_data[0][61] ));
Q_MX02 U754 ( .S(n103), .A0(\r_prefetch_data[0][60] ), .A1(n682), .Z(\c_prefetch_data[0][60] ));
Q_MX02 U755 ( .S(n103), .A0(\r_prefetch_data[0][59] ), .A1(n683), .Z(\c_prefetch_data[0][59] ));
Q_MX02 U756 ( .S(n103), .A0(\r_prefetch_data[0][58] ), .A1(n684), .Z(\c_prefetch_data[0][58] ));
Q_MX02 U757 ( .S(n103), .A0(\r_prefetch_data[0][57] ), .A1(n685), .Z(\c_prefetch_data[0][57] ));
Q_MX02 U758 ( .S(n103), .A0(\r_prefetch_data[0][56] ), .A1(n686), .Z(\c_prefetch_data[0][56] ));
Q_MX02 U759 ( .S(n103), .A0(\r_prefetch_data[0][55] ), .A1(n687), .Z(\c_prefetch_data[0][55] ));
Q_MX02 U760 ( .S(n103), .A0(\r_prefetch_data[0][54] ), .A1(n688), .Z(\c_prefetch_data[0][54] ));
Q_MX02 U761 ( .S(n103), .A0(\r_prefetch_data[0][53] ), .A1(n689), .Z(\c_prefetch_data[0][53] ));
Q_MX02 U762 ( .S(n103), .A0(\r_prefetch_data[0][52] ), .A1(n690), .Z(\c_prefetch_data[0][52] ));
Q_MX02 U763 ( .S(n103), .A0(\r_prefetch_data[0][51] ), .A1(n691), .Z(\c_prefetch_data[0][51] ));
Q_MX02 U764 ( .S(n103), .A0(\r_prefetch_data[0][50] ), .A1(n692), .Z(\c_prefetch_data[0][50] ));
Q_MX02 U765 ( .S(n103), .A0(\r_prefetch_data[0][49] ), .A1(n693), .Z(\c_prefetch_data[0][49] ));
Q_MX02 U766 ( .S(n103), .A0(\r_prefetch_data[0][48] ), .A1(n694), .Z(\c_prefetch_data[0][48] ));
Q_MX02 U767 ( .S(n103), .A0(\r_prefetch_data[0][47] ), .A1(n695), .Z(\c_prefetch_data[0][47] ));
Q_MX02 U768 ( .S(n103), .A0(\r_prefetch_data[0][46] ), .A1(n696), .Z(\c_prefetch_data[0][46] ));
Q_MX02 U769 ( .S(n103), .A0(\r_prefetch_data[0][45] ), .A1(n697), .Z(\c_prefetch_data[0][45] ));
Q_MX02 U770 ( .S(n103), .A0(\r_prefetch_data[0][44] ), .A1(n698), .Z(\c_prefetch_data[0][44] ));
Q_MX02 U771 ( .S(n103), .A0(\r_prefetch_data[0][43] ), .A1(n699), .Z(\c_prefetch_data[0][43] ));
Q_MX02 U772 ( .S(n103), .A0(\r_prefetch_data[0][42] ), .A1(n700), .Z(\c_prefetch_data[0][42] ));
Q_MX02 U773 ( .S(n103), .A0(\r_prefetch_data[0][41] ), .A1(n701), .Z(\c_prefetch_data[0][41] ));
Q_MX02 U774 ( .S(n103), .A0(\r_prefetch_data[0][40] ), .A1(n702), .Z(\c_prefetch_data[0][40] ));
Q_MX02 U775 ( .S(n103), .A0(\r_prefetch_data[0][39] ), .A1(n703), .Z(\c_prefetch_data[0][39] ));
Q_MX02 U776 ( .S(n103), .A0(\r_prefetch_data[0][38] ), .A1(n704), .Z(\c_prefetch_data[0][38] ));
Q_MX02 U777 ( .S(n103), .A0(\r_prefetch_data[0][37] ), .A1(n705), .Z(\c_prefetch_data[0][37] ));
Q_MX02 U778 ( .S(n103), .A0(\r_prefetch_data[0][36] ), .A1(n706), .Z(\c_prefetch_data[0][36] ));
Q_MX02 U779 ( .S(n103), .A0(\r_prefetch_data[0][35] ), .A1(n707), .Z(\c_prefetch_data[0][35] ));
Q_MX02 U780 ( .S(n103), .A0(\r_prefetch_data[0][34] ), .A1(n708), .Z(\c_prefetch_data[0][34] ));
Q_MX02 U781 ( .S(n103), .A0(\r_prefetch_data[0][33] ), .A1(n709), .Z(\c_prefetch_data[0][33] ));
Q_MX02 U782 ( .S(n103), .A0(\r_prefetch_data[0][32] ), .A1(n710), .Z(\c_prefetch_data[0][32] ));
Q_MX02 U783 ( .S(n103), .A0(\r_prefetch_data[0][31] ), .A1(n711), .Z(\c_prefetch_data[0][31] ));
Q_MX02 U784 ( .S(n103), .A0(\r_prefetch_data[0][30] ), .A1(n712), .Z(\c_prefetch_data[0][30] ));
Q_MX02 U785 ( .S(n103), .A0(\r_prefetch_data[0][29] ), .A1(n713), .Z(\c_prefetch_data[0][29] ));
Q_MX02 U786 ( .S(n103), .A0(\r_prefetch_data[0][28] ), .A1(n714), .Z(\c_prefetch_data[0][28] ));
Q_MX02 U787 ( .S(n103), .A0(\r_prefetch_data[0][27] ), .A1(n715), .Z(\c_prefetch_data[0][27] ));
Q_MX02 U788 ( .S(n103), .A0(\r_prefetch_data[0][26] ), .A1(n716), .Z(\c_prefetch_data[0][26] ));
Q_MX02 U789 ( .S(n103), .A0(\r_prefetch_data[0][25] ), .A1(n717), .Z(\c_prefetch_data[0][25] ));
Q_MX02 U790 ( .S(n103), .A0(\r_prefetch_data[0][24] ), .A1(n718), .Z(\c_prefetch_data[0][24] ));
Q_MX02 U791 ( .S(n103), .A0(\r_prefetch_data[0][23] ), .A1(n719), .Z(\c_prefetch_data[0][23] ));
Q_MX02 U792 ( .S(n103), .A0(\r_prefetch_data[0][22] ), .A1(n720), .Z(\c_prefetch_data[0][22] ));
Q_MX02 U793 ( .S(n103), .A0(\r_prefetch_data[0][21] ), .A1(n721), .Z(\c_prefetch_data[0][21] ));
Q_MX02 U794 ( .S(n103), .A0(\r_prefetch_data[0][20] ), .A1(n722), .Z(\c_prefetch_data[0][20] ));
Q_MX02 U795 ( .S(n103), .A0(\r_prefetch_data[0][19] ), .A1(n723), .Z(\c_prefetch_data[0][19] ));
Q_MX02 U796 ( .S(n103), .A0(\r_prefetch_data[0][18] ), .A1(n724), .Z(\c_prefetch_data[0][18] ));
Q_MX02 U797 ( .S(n103), .A0(\r_prefetch_data[0][17] ), .A1(n725), .Z(\c_prefetch_data[0][17] ));
Q_MX02 U798 ( .S(n103), .A0(\r_prefetch_data[0][16] ), .A1(n726), .Z(\c_prefetch_data[0][16] ));
Q_MX02 U799 ( .S(n103), .A0(\r_prefetch_data[0][15] ), .A1(n727), .Z(\c_prefetch_data[0][15] ));
Q_MX02 U800 ( .S(n103), .A0(\r_prefetch_data[0][14] ), .A1(n728), .Z(\c_prefetch_data[0][14] ));
Q_MX02 U801 ( .S(n103), .A0(\r_prefetch_data[0][13] ), .A1(n729), .Z(\c_prefetch_data[0][13] ));
Q_MX02 U802 ( .S(n103), .A0(\r_prefetch_data[0][12] ), .A1(n730), .Z(\c_prefetch_data[0][12] ));
Q_MX02 U803 ( .S(n103), .A0(\r_prefetch_data[0][11] ), .A1(n731), .Z(\c_prefetch_data[0][11] ));
Q_MX02 U804 ( .S(n103), .A0(\r_prefetch_data[0][10] ), .A1(n732), .Z(\c_prefetch_data[0][10] ));
Q_MX02 U805 ( .S(n103), .A0(\r_prefetch_data[0][9] ), .A1(n733), .Z(\c_prefetch_data[0][9] ));
Q_MX02 U806 ( .S(n103), .A0(\r_prefetch_data[0][8] ), .A1(n734), .Z(\c_prefetch_data[0][8] ));
Q_MX02 U807 ( .S(n103), .A0(\r_prefetch_data[0][7] ), .A1(n735), .Z(\c_prefetch_data[0][7] ));
Q_MX02 U808 ( .S(n103), .A0(\r_prefetch_data[0][6] ), .A1(n736), .Z(\c_prefetch_data[0][6] ));
Q_MX02 U809 ( .S(n103), .A0(\r_prefetch_data[0][5] ), .A1(n737), .Z(\c_prefetch_data[0][5] ));
Q_MX02 U810 ( .S(n103), .A0(\r_prefetch_data[0][4] ), .A1(n738), .Z(\c_prefetch_data[0][4] ));
Q_MX02 U811 ( .S(n103), .A0(\r_prefetch_data[0][3] ), .A1(n739), .Z(\c_prefetch_data[0][3] ));
Q_MX02 U812 ( .S(n103), .A0(\r_prefetch_data[0][2] ), .A1(n740), .Z(\c_prefetch_data[0][2] ));
Q_MX02 U813 ( .S(n103), .A0(\r_prefetch_data[0][1] ), .A1(n741), .Z(\c_prefetch_data[0][1] ));
Q_MX02 U814 ( .S(n103), .A0(\r_prefetch_data[0][0] ), .A1(n742), .Z(\c_prefetch_data[0][0] ));
Q_MX02 U815 ( .S(n104), .A0(\r_prefetch_data[1][83] ), .A1(n576), .Z(\c_prefetch_data[1][83] ));
Q_MX02 U816 ( .S(n104), .A0(\r_prefetch_data[1][82] ), .A1(n493), .Z(\c_prefetch_data[1][82] ));
Q_MX02 U817 ( .S(n104), .A0(\r_prefetch_data[1][81] ), .A1(n494), .Z(\c_prefetch_data[1][81] ));
Q_MX02 U818 ( .S(n104), .A0(\r_prefetch_data[1][80] ), .A1(n495), .Z(\c_prefetch_data[1][80] ));
Q_MX02 U819 ( .S(n104), .A0(\r_prefetch_data[1][79] ), .A1(n496), .Z(\c_prefetch_data[1][79] ));
Q_MX02 U820 ( .S(n104), .A0(\r_prefetch_data[1][78] ), .A1(n497), .Z(\c_prefetch_data[1][78] ));
Q_MX02 U821 ( .S(n104), .A0(\r_prefetch_data[1][77] ), .A1(n498), .Z(\c_prefetch_data[1][77] ));
Q_MX02 U822 ( .S(n104), .A0(\r_prefetch_data[1][76] ), .A1(n499), .Z(\c_prefetch_data[1][76] ));
Q_MX02 U823 ( .S(n104), .A0(\r_prefetch_data[1][75] ), .A1(n500), .Z(\c_prefetch_data[1][75] ));
Q_MX02 U824 ( .S(n104), .A0(\r_prefetch_data[1][74] ), .A1(n501), .Z(\c_prefetch_data[1][74] ));
Q_MX02 U825 ( .S(n104), .A0(\r_prefetch_data[1][73] ), .A1(n502), .Z(\c_prefetch_data[1][73] ));
Q_MX02 U826 ( .S(n104), .A0(\r_prefetch_data[1][72] ), .A1(n503), .Z(\c_prefetch_data[1][72] ));
Q_MX02 U827 ( .S(n104), .A0(\r_prefetch_data[1][71] ), .A1(n504), .Z(\c_prefetch_data[1][71] ));
Q_MX02 U828 ( .S(n104), .A0(\r_prefetch_data[1][70] ), .A1(n505), .Z(\c_prefetch_data[1][70] ));
Q_MX02 U829 ( .S(n104), .A0(\r_prefetch_data[1][69] ), .A1(n506), .Z(\c_prefetch_data[1][69] ));
Q_MX02 U830 ( .S(n104), .A0(\r_prefetch_data[1][68] ), .A1(n507), .Z(\c_prefetch_data[1][68] ));
Q_MX02 U831 ( .S(n104), .A0(\r_prefetch_data[1][67] ), .A1(n508), .Z(\c_prefetch_data[1][67] ));
Q_MX02 U832 ( .S(n104), .A0(\r_prefetch_data[1][66] ), .A1(n509), .Z(\c_prefetch_data[1][66] ));
Q_MX02 U833 ( .S(n104), .A0(\r_prefetch_data[1][65] ), .A1(n510), .Z(\c_prefetch_data[1][65] ));
Q_MX02 U834 ( .S(n104), .A0(\r_prefetch_data[1][64] ), .A1(n511), .Z(\c_prefetch_data[1][64] ));
Q_MX02 U835 ( .S(n104), .A0(\r_prefetch_data[1][63] ), .A1(n512), .Z(\c_prefetch_data[1][63] ));
Q_MX02 U836 ( .S(n104), .A0(\r_prefetch_data[1][62] ), .A1(n513), .Z(\c_prefetch_data[1][62] ));
Q_MX02 U837 ( .S(n104), .A0(\r_prefetch_data[1][61] ), .A1(n514), .Z(\c_prefetch_data[1][61] ));
Q_MX02 U838 ( .S(n104), .A0(\r_prefetch_data[1][60] ), .A1(n515), .Z(\c_prefetch_data[1][60] ));
Q_MX02 U839 ( .S(n104), .A0(\r_prefetch_data[1][59] ), .A1(n516), .Z(\c_prefetch_data[1][59] ));
Q_MX02 U840 ( .S(n104), .A0(\r_prefetch_data[1][58] ), .A1(n517), .Z(\c_prefetch_data[1][58] ));
Q_MX02 U841 ( .S(n104), .A0(\r_prefetch_data[1][57] ), .A1(n518), .Z(\c_prefetch_data[1][57] ));
Q_MX02 U842 ( .S(n104), .A0(\r_prefetch_data[1][56] ), .A1(n519), .Z(\c_prefetch_data[1][56] ));
Q_MX02 U843 ( .S(n104), .A0(\r_prefetch_data[1][55] ), .A1(n520), .Z(\c_prefetch_data[1][55] ));
Q_MX02 U844 ( .S(n104), .A0(\r_prefetch_data[1][54] ), .A1(n521), .Z(\c_prefetch_data[1][54] ));
Q_MX02 U845 ( .S(n104), .A0(\r_prefetch_data[1][53] ), .A1(n522), .Z(\c_prefetch_data[1][53] ));
Q_MX02 U846 ( .S(n104), .A0(\r_prefetch_data[1][52] ), .A1(n523), .Z(\c_prefetch_data[1][52] ));
Q_MX02 U847 ( .S(n104), .A0(\r_prefetch_data[1][51] ), .A1(n524), .Z(\c_prefetch_data[1][51] ));
Q_MX02 U848 ( .S(n104), .A0(\r_prefetch_data[1][50] ), .A1(n525), .Z(\c_prefetch_data[1][50] ));
Q_MX02 U849 ( .S(n104), .A0(\r_prefetch_data[1][49] ), .A1(n526), .Z(\c_prefetch_data[1][49] ));
Q_MX02 U850 ( .S(n104), .A0(\r_prefetch_data[1][48] ), .A1(n527), .Z(\c_prefetch_data[1][48] ));
Q_MX02 U851 ( .S(n104), .A0(\r_prefetch_data[1][47] ), .A1(n528), .Z(\c_prefetch_data[1][47] ));
Q_MX02 U852 ( .S(n104), .A0(\r_prefetch_data[1][46] ), .A1(n529), .Z(\c_prefetch_data[1][46] ));
Q_MX02 U853 ( .S(n104), .A0(\r_prefetch_data[1][45] ), .A1(n530), .Z(\c_prefetch_data[1][45] ));
Q_MX02 U854 ( .S(n104), .A0(\r_prefetch_data[1][44] ), .A1(n531), .Z(\c_prefetch_data[1][44] ));
Q_MX02 U855 ( .S(n104), .A0(\r_prefetch_data[1][43] ), .A1(n532), .Z(\c_prefetch_data[1][43] ));
Q_MX02 U856 ( .S(n104), .A0(\r_prefetch_data[1][42] ), .A1(n533), .Z(\c_prefetch_data[1][42] ));
Q_MX02 U857 ( .S(n104), .A0(\r_prefetch_data[1][41] ), .A1(n534), .Z(\c_prefetch_data[1][41] ));
Q_MX02 U858 ( .S(n104), .A0(\r_prefetch_data[1][40] ), .A1(n535), .Z(\c_prefetch_data[1][40] ));
Q_MX02 U859 ( .S(n104), .A0(\r_prefetch_data[1][39] ), .A1(n536), .Z(\c_prefetch_data[1][39] ));
Q_MX02 U860 ( .S(n104), .A0(\r_prefetch_data[1][38] ), .A1(n537), .Z(\c_prefetch_data[1][38] ));
Q_MX02 U861 ( .S(n104), .A0(\r_prefetch_data[1][37] ), .A1(n538), .Z(\c_prefetch_data[1][37] ));
Q_MX02 U862 ( .S(n104), .A0(\r_prefetch_data[1][36] ), .A1(n539), .Z(\c_prefetch_data[1][36] ));
Q_MX02 U863 ( .S(n104), .A0(\r_prefetch_data[1][35] ), .A1(n540), .Z(\c_prefetch_data[1][35] ));
Q_MX02 U864 ( .S(n104), .A0(\r_prefetch_data[1][34] ), .A1(n541), .Z(\c_prefetch_data[1][34] ));
Q_MX02 U865 ( .S(n104), .A0(\r_prefetch_data[1][33] ), .A1(n542), .Z(\c_prefetch_data[1][33] ));
Q_MX02 U866 ( .S(n104), .A0(\r_prefetch_data[1][32] ), .A1(n543), .Z(\c_prefetch_data[1][32] ));
Q_MX02 U867 ( .S(n104), .A0(\r_prefetch_data[1][31] ), .A1(n544), .Z(\c_prefetch_data[1][31] ));
Q_MX02 U868 ( .S(n104), .A0(\r_prefetch_data[1][30] ), .A1(n545), .Z(\c_prefetch_data[1][30] ));
Q_MX02 U869 ( .S(n104), .A0(\r_prefetch_data[1][29] ), .A1(n546), .Z(\c_prefetch_data[1][29] ));
Q_MX02 U870 ( .S(n104), .A0(\r_prefetch_data[1][28] ), .A1(n547), .Z(\c_prefetch_data[1][28] ));
Q_MX02 U871 ( .S(n104), .A0(\r_prefetch_data[1][27] ), .A1(n548), .Z(\c_prefetch_data[1][27] ));
Q_MX02 U872 ( .S(n104), .A0(\r_prefetch_data[1][26] ), .A1(n549), .Z(\c_prefetch_data[1][26] ));
Q_MX02 U873 ( .S(n104), .A0(\r_prefetch_data[1][25] ), .A1(n550), .Z(\c_prefetch_data[1][25] ));
Q_MX02 U874 ( .S(n104), .A0(\r_prefetch_data[1][24] ), .A1(n551), .Z(\c_prefetch_data[1][24] ));
Q_MX02 U875 ( .S(n104), .A0(\r_prefetch_data[1][23] ), .A1(n552), .Z(\c_prefetch_data[1][23] ));
Q_MX02 U876 ( .S(n104), .A0(\r_prefetch_data[1][22] ), .A1(n553), .Z(\c_prefetch_data[1][22] ));
Q_MX02 U877 ( .S(n104), .A0(\r_prefetch_data[1][21] ), .A1(n554), .Z(\c_prefetch_data[1][21] ));
Q_MX02 U878 ( .S(n104), .A0(\r_prefetch_data[1][20] ), .A1(n555), .Z(\c_prefetch_data[1][20] ));
Q_MX02 U879 ( .S(n104), .A0(\r_prefetch_data[1][19] ), .A1(n556), .Z(\c_prefetch_data[1][19] ));
Q_MX02 U880 ( .S(n104), .A0(\r_prefetch_data[1][18] ), .A1(n557), .Z(\c_prefetch_data[1][18] ));
Q_MX02 U881 ( .S(n104), .A0(\r_prefetch_data[1][17] ), .A1(n558), .Z(\c_prefetch_data[1][17] ));
Q_MX02 U882 ( .S(n104), .A0(\r_prefetch_data[1][16] ), .A1(n559), .Z(\c_prefetch_data[1][16] ));
Q_MX02 U883 ( .S(n104), .A0(\r_prefetch_data[1][15] ), .A1(n560), .Z(\c_prefetch_data[1][15] ));
Q_MX02 U884 ( .S(n104), .A0(\r_prefetch_data[1][14] ), .A1(n561), .Z(\c_prefetch_data[1][14] ));
Q_MX02 U885 ( .S(n104), .A0(\r_prefetch_data[1][13] ), .A1(n562), .Z(\c_prefetch_data[1][13] ));
Q_MX02 U886 ( .S(n104), .A0(\r_prefetch_data[1][12] ), .A1(n563), .Z(\c_prefetch_data[1][12] ));
Q_MX02 U887 ( .S(n104), .A0(\r_prefetch_data[1][11] ), .A1(n564), .Z(\c_prefetch_data[1][11] ));
Q_MX02 U888 ( .S(n104), .A0(\r_prefetch_data[1][10] ), .A1(n565), .Z(\c_prefetch_data[1][10] ));
Q_MX02 U889 ( .S(n104), .A0(\r_prefetch_data[1][9] ), .A1(n566), .Z(\c_prefetch_data[1][9] ));
Q_MX02 U890 ( .S(n104), .A0(\r_prefetch_data[1][8] ), .A1(n567), .Z(\c_prefetch_data[1][8] ));
Q_MX02 U891 ( .S(n104), .A0(\r_prefetch_data[1][7] ), .A1(n568), .Z(\c_prefetch_data[1][7] ));
Q_MX02 U892 ( .S(n104), .A0(\r_prefetch_data[1][6] ), .A1(n569), .Z(\c_prefetch_data[1][6] ));
Q_MX02 U893 ( .S(n104), .A0(\r_prefetch_data[1][5] ), .A1(n570), .Z(\c_prefetch_data[1][5] ));
Q_MX02 U894 ( .S(n104), .A0(\r_prefetch_data[1][4] ), .A1(n571), .Z(\c_prefetch_data[1][4] ));
Q_MX02 U895 ( .S(n104), .A0(\r_prefetch_data[1][3] ), .A1(n572), .Z(\c_prefetch_data[1][3] ));
Q_MX02 U896 ( .S(n104), .A0(\r_prefetch_data[1][2] ), .A1(n573), .Z(\c_prefetch_data[1][2] ));
Q_MX02 U897 ( .S(n104), .A0(\r_prefetch_data[1][1] ), .A1(n574), .Z(\c_prefetch_data[1][1] ));
Q_MX02 U898 ( .S(n104), .A0(\r_prefetch_data[1][0] ), .A1(n575), .Z(\c_prefetch_data[1][0] ));
Q_MX02 U899 ( .S(n105), .A0(\r_prefetch_data[2][83] ), .A1(n409), .Z(\c_prefetch_data[2][83] ));
Q_MX02 U900 ( .S(n105), .A0(\r_prefetch_data[2][82] ), .A1(n326), .Z(\c_prefetch_data[2][82] ));
Q_MX02 U901 ( .S(n105), .A0(\r_prefetch_data[2][81] ), .A1(n327), .Z(\c_prefetch_data[2][81] ));
Q_MX02 U902 ( .S(n105), .A0(\r_prefetch_data[2][80] ), .A1(n328), .Z(\c_prefetch_data[2][80] ));
Q_MX02 U903 ( .S(n105), .A0(\r_prefetch_data[2][79] ), .A1(n329), .Z(\c_prefetch_data[2][79] ));
Q_MX02 U904 ( .S(n105), .A0(\r_prefetch_data[2][78] ), .A1(n330), .Z(\c_prefetch_data[2][78] ));
Q_MX02 U905 ( .S(n105), .A0(\r_prefetch_data[2][77] ), .A1(n331), .Z(\c_prefetch_data[2][77] ));
Q_MX02 U906 ( .S(n105), .A0(\r_prefetch_data[2][76] ), .A1(n332), .Z(\c_prefetch_data[2][76] ));
Q_MX02 U907 ( .S(n105), .A0(\r_prefetch_data[2][75] ), .A1(n333), .Z(\c_prefetch_data[2][75] ));
Q_MX02 U908 ( .S(n105), .A0(\r_prefetch_data[2][74] ), .A1(n334), .Z(\c_prefetch_data[2][74] ));
Q_MX02 U909 ( .S(n105), .A0(\r_prefetch_data[2][73] ), .A1(n335), .Z(\c_prefetch_data[2][73] ));
Q_MX02 U910 ( .S(n105), .A0(\r_prefetch_data[2][72] ), .A1(n336), .Z(\c_prefetch_data[2][72] ));
Q_MX02 U911 ( .S(n105), .A0(\r_prefetch_data[2][71] ), .A1(n337), .Z(\c_prefetch_data[2][71] ));
Q_MX02 U912 ( .S(n105), .A0(\r_prefetch_data[2][70] ), .A1(n338), .Z(\c_prefetch_data[2][70] ));
Q_MX02 U913 ( .S(n105), .A0(\r_prefetch_data[2][69] ), .A1(n339), .Z(\c_prefetch_data[2][69] ));
Q_MX02 U914 ( .S(n105), .A0(\r_prefetch_data[2][68] ), .A1(n340), .Z(\c_prefetch_data[2][68] ));
Q_MX02 U915 ( .S(n105), .A0(\r_prefetch_data[2][67] ), .A1(n341), .Z(\c_prefetch_data[2][67] ));
Q_MX02 U916 ( .S(n105), .A0(\r_prefetch_data[2][66] ), .A1(n342), .Z(\c_prefetch_data[2][66] ));
Q_MX02 U917 ( .S(n105), .A0(\r_prefetch_data[2][65] ), .A1(n343), .Z(\c_prefetch_data[2][65] ));
Q_MX02 U918 ( .S(n105), .A0(\r_prefetch_data[2][64] ), .A1(n344), .Z(\c_prefetch_data[2][64] ));
Q_MX02 U919 ( .S(n105), .A0(\r_prefetch_data[2][63] ), .A1(n345), .Z(\c_prefetch_data[2][63] ));
Q_MX02 U920 ( .S(n105), .A0(\r_prefetch_data[2][62] ), .A1(n346), .Z(\c_prefetch_data[2][62] ));
Q_MX02 U921 ( .S(n105), .A0(\r_prefetch_data[2][61] ), .A1(n347), .Z(\c_prefetch_data[2][61] ));
Q_MX02 U922 ( .S(n105), .A0(\r_prefetch_data[2][60] ), .A1(n348), .Z(\c_prefetch_data[2][60] ));
Q_MX02 U923 ( .S(n105), .A0(\r_prefetch_data[2][59] ), .A1(n349), .Z(\c_prefetch_data[2][59] ));
Q_MX02 U924 ( .S(n105), .A0(\r_prefetch_data[2][58] ), .A1(n350), .Z(\c_prefetch_data[2][58] ));
Q_MX02 U925 ( .S(n105), .A0(\r_prefetch_data[2][57] ), .A1(n351), .Z(\c_prefetch_data[2][57] ));
Q_MX02 U926 ( .S(n105), .A0(\r_prefetch_data[2][56] ), .A1(n352), .Z(\c_prefetch_data[2][56] ));
Q_MX02 U927 ( .S(n105), .A0(\r_prefetch_data[2][55] ), .A1(n353), .Z(\c_prefetch_data[2][55] ));
Q_MX02 U928 ( .S(n105), .A0(\r_prefetch_data[2][54] ), .A1(n354), .Z(\c_prefetch_data[2][54] ));
Q_MX02 U929 ( .S(n105), .A0(\r_prefetch_data[2][53] ), .A1(n355), .Z(\c_prefetch_data[2][53] ));
Q_MX02 U930 ( .S(n105), .A0(\r_prefetch_data[2][52] ), .A1(n356), .Z(\c_prefetch_data[2][52] ));
Q_MX02 U931 ( .S(n105), .A0(\r_prefetch_data[2][51] ), .A1(n357), .Z(\c_prefetch_data[2][51] ));
Q_MX02 U932 ( .S(n105), .A0(\r_prefetch_data[2][50] ), .A1(n358), .Z(\c_prefetch_data[2][50] ));
Q_MX02 U933 ( .S(n105), .A0(\r_prefetch_data[2][49] ), .A1(n359), .Z(\c_prefetch_data[2][49] ));
Q_MX02 U934 ( .S(n105), .A0(\r_prefetch_data[2][48] ), .A1(n360), .Z(\c_prefetch_data[2][48] ));
Q_MX02 U935 ( .S(n105), .A0(\r_prefetch_data[2][47] ), .A1(n361), .Z(\c_prefetch_data[2][47] ));
Q_MX02 U936 ( .S(n105), .A0(\r_prefetch_data[2][46] ), .A1(n362), .Z(\c_prefetch_data[2][46] ));
Q_MX02 U937 ( .S(n105), .A0(\r_prefetch_data[2][45] ), .A1(n363), .Z(\c_prefetch_data[2][45] ));
Q_MX02 U938 ( .S(n105), .A0(\r_prefetch_data[2][44] ), .A1(n364), .Z(\c_prefetch_data[2][44] ));
Q_MX02 U939 ( .S(n105), .A0(\r_prefetch_data[2][43] ), .A1(n365), .Z(\c_prefetch_data[2][43] ));
Q_MX02 U940 ( .S(n105), .A0(\r_prefetch_data[2][42] ), .A1(n366), .Z(\c_prefetch_data[2][42] ));
Q_MX02 U941 ( .S(n105), .A0(\r_prefetch_data[2][41] ), .A1(n367), .Z(\c_prefetch_data[2][41] ));
Q_MX02 U942 ( .S(n105), .A0(\r_prefetch_data[2][40] ), .A1(n368), .Z(\c_prefetch_data[2][40] ));
Q_MX02 U943 ( .S(n105), .A0(\r_prefetch_data[2][39] ), .A1(n369), .Z(\c_prefetch_data[2][39] ));
Q_MX02 U944 ( .S(n105), .A0(\r_prefetch_data[2][38] ), .A1(n370), .Z(\c_prefetch_data[2][38] ));
Q_MX02 U945 ( .S(n105), .A0(\r_prefetch_data[2][37] ), .A1(n371), .Z(\c_prefetch_data[2][37] ));
Q_MX02 U946 ( .S(n105), .A0(\r_prefetch_data[2][36] ), .A1(n372), .Z(\c_prefetch_data[2][36] ));
Q_MX02 U947 ( .S(n105), .A0(\r_prefetch_data[2][35] ), .A1(n373), .Z(\c_prefetch_data[2][35] ));
Q_MX02 U948 ( .S(n105), .A0(\r_prefetch_data[2][34] ), .A1(n374), .Z(\c_prefetch_data[2][34] ));
Q_MX02 U949 ( .S(n105), .A0(\r_prefetch_data[2][33] ), .A1(n375), .Z(\c_prefetch_data[2][33] ));
Q_MX02 U950 ( .S(n105), .A0(\r_prefetch_data[2][32] ), .A1(n376), .Z(\c_prefetch_data[2][32] ));
Q_MX02 U951 ( .S(n105), .A0(\r_prefetch_data[2][31] ), .A1(n377), .Z(\c_prefetch_data[2][31] ));
Q_MX02 U952 ( .S(n105), .A0(\r_prefetch_data[2][30] ), .A1(n378), .Z(\c_prefetch_data[2][30] ));
Q_MX02 U953 ( .S(n105), .A0(\r_prefetch_data[2][29] ), .A1(n379), .Z(\c_prefetch_data[2][29] ));
Q_MX02 U954 ( .S(n105), .A0(\r_prefetch_data[2][28] ), .A1(n380), .Z(\c_prefetch_data[2][28] ));
Q_MX02 U955 ( .S(n105), .A0(\r_prefetch_data[2][27] ), .A1(n381), .Z(\c_prefetch_data[2][27] ));
Q_MX02 U956 ( .S(n105), .A0(\r_prefetch_data[2][26] ), .A1(n382), .Z(\c_prefetch_data[2][26] ));
Q_MX02 U957 ( .S(n105), .A0(\r_prefetch_data[2][25] ), .A1(n383), .Z(\c_prefetch_data[2][25] ));
Q_MX02 U958 ( .S(n105), .A0(\r_prefetch_data[2][24] ), .A1(n384), .Z(\c_prefetch_data[2][24] ));
Q_MX02 U959 ( .S(n105), .A0(\r_prefetch_data[2][23] ), .A1(n385), .Z(\c_prefetch_data[2][23] ));
Q_MX02 U960 ( .S(n105), .A0(\r_prefetch_data[2][22] ), .A1(n386), .Z(\c_prefetch_data[2][22] ));
Q_MX02 U961 ( .S(n105), .A0(\r_prefetch_data[2][21] ), .A1(n387), .Z(\c_prefetch_data[2][21] ));
Q_MX02 U962 ( .S(n105), .A0(\r_prefetch_data[2][20] ), .A1(n388), .Z(\c_prefetch_data[2][20] ));
Q_MX02 U963 ( .S(n105), .A0(\r_prefetch_data[2][19] ), .A1(n389), .Z(\c_prefetch_data[2][19] ));
Q_MX02 U964 ( .S(n105), .A0(\r_prefetch_data[2][18] ), .A1(n390), .Z(\c_prefetch_data[2][18] ));
Q_MX02 U965 ( .S(n105), .A0(\r_prefetch_data[2][17] ), .A1(n391), .Z(\c_prefetch_data[2][17] ));
Q_MX02 U966 ( .S(n105), .A0(\r_prefetch_data[2][16] ), .A1(n392), .Z(\c_prefetch_data[2][16] ));
Q_MX02 U967 ( .S(n105), .A0(\r_prefetch_data[2][15] ), .A1(n393), .Z(\c_prefetch_data[2][15] ));
Q_MX02 U968 ( .S(n105), .A0(\r_prefetch_data[2][14] ), .A1(n394), .Z(\c_prefetch_data[2][14] ));
Q_MX02 U969 ( .S(n105), .A0(\r_prefetch_data[2][13] ), .A1(n395), .Z(\c_prefetch_data[2][13] ));
Q_MX02 U970 ( .S(n105), .A0(\r_prefetch_data[2][12] ), .A1(n396), .Z(\c_prefetch_data[2][12] ));
Q_MX02 U971 ( .S(n105), .A0(\r_prefetch_data[2][11] ), .A1(n397), .Z(\c_prefetch_data[2][11] ));
Q_MX02 U972 ( .S(n105), .A0(\r_prefetch_data[2][10] ), .A1(n398), .Z(\c_prefetch_data[2][10] ));
Q_MX02 U973 ( .S(n105), .A0(\r_prefetch_data[2][9] ), .A1(n399), .Z(\c_prefetch_data[2][9] ));
Q_MX02 U974 ( .S(n105), .A0(\r_prefetch_data[2][8] ), .A1(n400), .Z(\c_prefetch_data[2][8] ));
Q_MX02 U975 ( .S(n105), .A0(\r_prefetch_data[2][7] ), .A1(n401), .Z(\c_prefetch_data[2][7] ));
Q_MX02 U976 ( .S(n105), .A0(\r_prefetch_data[2][6] ), .A1(n402), .Z(\c_prefetch_data[2][6] ));
Q_MX02 U977 ( .S(n105), .A0(\r_prefetch_data[2][5] ), .A1(n403), .Z(\c_prefetch_data[2][5] ));
Q_MX02 U978 ( .S(n105), .A0(\r_prefetch_data[2][4] ), .A1(n404), .Z(\c_prefetch_data[2][4] ));
Q_MX02 U979 ( .S(n105), .A0(\r_prefetch_data[2][3] ), .A1(n405), .Z(\c_prefetch_data[2][3] ));
Q_MX02 U980 ( .S(n105), .A0(\r_prefetch_data[2][2] ), .A1(n406), .Z(\c_prefetch_data[2][2] ));
Q_MX02 U981 ( .S(n105), .A0(\r_prefetch_data[2][1] ), .A1(n407), .Z(\c_prefetch_data[2][1] ));
Q_MX02 U982 ( .S(n105), .A0(\r_prefetch_data[2][0] ), .A1(n408), .Z(\c_prefetch_data[2][0] ));
Q_MX02 U983 ( .S(n139), .A0(n106), .A1(n325), .Z(c_prefetch_full));
Q_MX02 U984 ( .S(n106), .A0(n86), .A1(r_prefetch_full), .Z(n325));
Q_AN02 U985 ( .A0(prefetch_lden_mem[2]), .A1(mem_ecc_error), .Z(n409));
Q_AN02 U986 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[82]), .Z(n410));
Q_AN02 U987 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[81]), .Z(n411));
Q_AN02 U988 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[80]), .Z(n412));
Q_AN02 U989 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[79]), .Z(n413));
Q_AN02 U990 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[78]), .Z(n414));
Q_AN02 U991 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[77]), .Z(n415));
Q_AN02 U992 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[76]), .Z(n416));
Q_AN02 U993 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[75]), .Z(n417));
Q_AN02 U994 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[74]), .Z(n418));
Q_AN02 U995 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[73]), .Z(n419));
Q_AN02 U996 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[72]), .Z(n420));
Q_AN02 U997 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[71]), .Z(n421));
Q_AN02 U998 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[70]), .Z(n422));
Q_AN02 U999 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[69]), .Z(n423));
Q_AN02 U1000 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[68]), .Z(n424));
Q_AN02 U1001 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[67]), .Z(n425));
Q_AN02 U1002 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[66]), .Z(n426));
Q_AN02 U1003 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[65]), .Z(n427));
Q_AN02 U1004 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[64]), .Z(n428));
Q_AN02 U1005 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[63]), .Z(n429));
Q_AN02 U1006 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[62]), .Z(n430));
Q_AN02 U1007 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[61]), .Z(n431));
Q_AN02 U1008 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[60]), .Z(n432));
Q_AN02 U1009 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[59]), .Z(n433));
Q_AN02 U1010 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[58]), .Z(n434));
Q_AN02 U1011 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[57]), .Z(n435));
Q_AN02 U1012 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[56]), .Z(n436));
Q_AN02 U1013 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[55]), .Z(n437));
Q_AN02 U1014 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[54]), .Z(n438));
Q_AN02 U1015 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[53]), .Z(n439));
Q_AN02 U1016 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[52]), .Z(n440));
Q_AN02 U1017 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[51]), .Z(n441));
Q_AN02 U1018 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[50]), .Z(n442));
Q_AN02 U1019 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[49]), .Z(n443));
Q_AN02 U1020 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[48]), .Z(n444));
Q_AN02 U1021 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[47]), .Z(n445));
Q_AN02 U1022 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[46]), .Z(n446));
Q_AN02 U1023 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[45]), .Z(n447));
Q_AN02 U1024 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[44]), .Z(n448));
Q_AN02 U1025 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[43]), .Z(n449));
Q_AN02 U1026 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[42]), .Z(n450));
Q_AN02 U1027 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[41]), .Z(n451));
Q_AN02 U1028 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[40]), .Z(n452));
Q_AN02 U1029 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[39]), .Z(n453));
Q_AN02 U1030 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[38]), .Z(n454));
Q_AN02 U1031 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[37]), .Z(n455));
Q_AN02 U1032 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[36]), .Z(n456));
Q_AN02 U1033 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[35]), .Z(n457));
Q_AN02 U1034 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[34]), .Z(n458));
Q_AN02 U1035 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[33]), .Z(n459));
Q_AN02 U1036 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[32]), .Z(n460));
Q_AN02 U1037 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[31]), .Z(n461));
Q_AN02 U1038 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[30]), .Z(n462));
Q_AN02 U1039 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[29]), .Z(n463));
Q_AN02 U1040 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[28]), .Z(n464));
Q_AN02 U1041 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[27]), .Z(n465));
Q_AN02 U1042 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[26]), .Z(n466));
Q_AN02 U1043 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[25]), .Z(n467));
Q_AN02 U1044 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[24]), .Z(n468));
Q_AN02 U1045 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[23]), .Z(n469));
Q_AN02 U1046 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[22]), .Z(n470));
Q_AN02 U1047 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[21]), .Z(n471));
Q_AN02 U1048 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[20]), .Z(n472));
Q_AN02 U1049 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[19]), .Z(n473));
Q_AN02 U1050 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[18]), .Z(n474));
Q_AN02 U1051 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[17]), .Z(n475));
Q_AN02 U1052 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[16]), .Z(n476));
Q_AN02 U1053 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[15]), .Z(n477));
Q_AN02 U1054 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[14]), .Z(n478));
Q_AN02 U1055 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[13]), .Z(n479));
Q_AN02 U1056 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[12]), .Z(n480));
Q_AN02 U1057 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[11]), .Z(n481));
Q_AN02 U1058 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[10]), .Z(n482));
Q_AN02 U1059 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[9]), .Z(n483));
Q_AN02 U1060 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[8]), .Z(n484));
Q_AN02 U1061 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[7]), .Z(n485));
Q_AN02 U1062 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[6]), .Z(n486));
Q_AN02 U1063 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[5]), .Z(n487));
Q_AN02 U1064 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[4]), .Z(n488));
Q_AN02 U1065 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[3]), .Z(n489));
Q_AN02 U1066 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[2]), .Z(n490));
Q_AN02 U1067 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[1]), .Z(n491));
Q_AN02 U1068 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[0]), .Z(n492));
Q_AO21 U1069 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[82]), .B0(n410), .Z(n326));
Q_AO21 U1070 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[81]), .B0(n411), .Z(n327));
Q_AO21 U1071 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[80]), .B0(n412), .Z(n328));
Q_AO21 U1072 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[79]), .B0(n413), .Z(n329));
Q_AO21 U1073 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[78]), .B0(n414), .Z(n330));
Q_AO21 U1074 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[77]), .B0(n415), .Z(n331));
Q_AO21 U1075 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[76]), .B0(n416), .Z(n332));
Q_AO21 U1076 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[75]), .B0(n417), .Z(n333));
Q_AO21 U1077 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[74]), .B0(n418), .Z(n334));
Q_AO21 U1078 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[73]), .B0(n419), .Z(n335));
Q_AO21 U1079 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[72]), .B0(n420), .Z(n336));
Q_AO21 U1080 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[71]), .B0(n421), .Z(n337));
Q_AO21 U1081 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[70]), .B0(n422), .Z(n338));
Q_AO21 U1082 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[69]), .B0(n423), .Z(n339));
Q_AO21 U1083 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[68]), .B0(n424), .Z(n340));
Q_AO21 U1084 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[67]), .B0(n425), .Z(n341));
Q_AO21 U1085 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[66]), .B0(n426), .Z(n342));
Q_AO21 U1086 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[65]), .B0(n427), .Z(n343));
Q_AO21 U1087 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[64]), .B0(n428), .Z(n344));
Q_AO21 U1088 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[63]), .B0(n429), .Z(n345));
Q_AO21 U1089 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[62]), .B0(n430), .Z(n346));
Q_AO21 U1090 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[61]), .B0(n431), .Z(n347));
Q_AO21 U1091 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[60]), .B0(n432), .Z(n348));
Q_AO21 U1092 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[59]), .B0(n433), .Z(n349));
Q_AO21 U1093 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[58]), .B0(n434), .Z(n350));
Q_AO21 U1094 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[57]), .B0(n435), .Z(n351));
Q_AO21 U1095 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[56]), .B0(n436), .Z(n352));
Q_AO21 U1096 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[55]), .B0(n437), .Z(n353));
Q_AO21 U1097 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[54]), .B0(n438), .Z(n354));
Q_AO21 U1098 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[53]), .B0(n439), .Z(n355));
Q_AO21 U1099 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[52]), .B0(n440), .Z(n356));
Q_AO21 U1100 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[51]), .B0(n441), .Z(n357));
Q_AO21 U1101 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[50]), .B0(n442), .Z(n358));
Q_AO21 U1102 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[49]), .B0(n443), .Z(n359));
Q_AO21 U1103 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[48]), .B0(n444), .Z(n360));
Q_AO21 U1104 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[47]), .B0(n445), .Z(n361));
Q_AO21 U1105 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[46]), .B0(n446), .Z(n362));
Q_AO21 U1106 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[45]), .B0(n447), .Z(n363));
Q_AO21 U1107 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[44]), .B0(n448), .Z(n364));
Q_AO21 U1108 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[43]), .B0(n449), .Z(n365));
Q_AO21 U1109 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[42]), .B0(n450), .Z(n366));
Q_AO21 U1110 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[41]), .B0(n451), .Z(n367));
Q_AO21 U1111 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[40]), .B0(n452), .Z(n368));
Q_AO21 U1112 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[39]), .B0(n453), .Z(n369));
Q_AO21 U1113 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[38]), .B0(n454), .Z(n370));
Q_AO21 U1114 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[37]), .B0(n455), .Z(n371));
Q_AO21 U1115 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[36]), .B0(n456), .Z(n372));
Q_AO21 U1116 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[35]), .B0(n457), .Z(n373));
Q_AO21 U1117 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[34]), .B0(n458), .Z(n374));
Q_AO21 U1118 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[33]), .B0(n459), .Z(n375));
Q_AO21 U1119 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[32]), .B0(n460), .Z(n376));
Q_AO21 U1120 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[31]), .B0(n461), .Z(n377));
Q_AO21 U1121 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[30]), .B0(n462), .Z(n378));
Q_AO21 U1122 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[29]), .B0(n463), .Z(n379));
Q_AO21 U1123 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[28]), .B0(n464), .Z(n380));
Q_AO21 U1124 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[27]), .B0(n465), .Z(n381));
Q_AO21 U1125 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[26]), .B0(n466), .Z(n382));
Q_AO21 U1126 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[25]), .B0(n467), .Z(n383));
Q_AO21 U1127 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[24]), .B0(n468), .Z(n384));
Q_AO21 U1128 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[23]), .B0(n469), .Z(n385));
Q_AO21 U1129 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[22]), .B0(n470), .Z(n386));
Q_AO21 U1130 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[21]), .B0(n471), .Z(n387));
Q_AO21 U1131 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[20]), .B0(n472), .Z(n388));
Q_AO21 U1132 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[19]), .B0(n473), .Z(n389));
Q_AO21 U1133 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[18]), .B0(n474), .Z(n390));
Q_AO21 U1134 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[17]), .B0(n475), .Z(n391));
Q_AO21 U1135 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[16]), .B0(n476), .Z(n392));
Q_AO21 U1136 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[15]), .B0(n477), .Z(n393));
Q_AO21 U1137 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[14]), .B0(n478), .Z(n394));
Q_AO21 U1138 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[13]), .B0(n479), .Z(n395));
Q_AO21 U1139 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[12]), .B0(n480), .Z(n396));
Q_AO21 U1140 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[11]), .B0(n481), .Z(n397));
Q_AO21 U1141 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[10]), .B0(n482), .Z(n398));
Q_AO21 U1142 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[9]), .B0(n483), .Z(n399));
Q_AO21 U1143 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[8]), .B0(n484), .Z(n400));
Q_AO21 U1144 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[7]), .B0(n485), .Z(n401));
Q_AO21 U1145 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[6]), .B0(n486), .Z(n402));
Q_AO21 U1146 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[5]), .B0(n487), .Z(n403));
Q_AO21 U1147 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[4]), .B0(n488), .Z(n404));
Q_AO21 U1148 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[3]), .B0(n489), .Z(n405));
Q_AO21 U1149 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[2]), .B0(n490), .Z(n406));
Q_AO21 U1150 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[1]), .B0(n491), .Z(n407));
Q_AO21 U1151 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[0]), .B0(n492), .Z(n408));
Q_AN02 U1152 ( .A0(prefetch_lden_mem[1]), .A1(mem_ecc_error), .Z(n576));
Q_AN02 U1153 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[82]), .Z(n577));
Q_AN02 U1154 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[81]), .Z(n578));
Q_AN02 U1155 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[80]), .Z(n579));
Q_AN02 U1156 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[79]), .Z(n580));
Q_AN02 U1157 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[78]), .Z(n581));
Q_AN02 U1158 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[77]), .Z(n582));
Q_AN02 U1159 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[76]), .Z(n583));
Q_AN02 U1160 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[75]), .Z(n584));
Q_AN02 U1161 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[74]), .Z(n585));
Q_AN02 U1162 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[73]), .Z(n586));
Q_AN02 U1163 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[72]), .Z(n587));
Q_AN02 U1164 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[71]), .Z(n588));
Q_AN02 U1165 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[70]), .Z(n589));
Q_AN02 U1166 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[69]), .Z(n590));
Q_AN02 U1167 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[68]), .Z(n591));
Q_AN02 U1168 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[67]), .Z(n592));
Q_AN02 U1169 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[66]), .Z(n593));
Q_AN02 U1170 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[65]), .Z(n594));
Q_AN02 U1171 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[64]), .Z(n595));
Q_AN02 U1172 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[63]), .Z(n596));
Q_AN02 U1173 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[62]), .Z(n597));
Q_AN02 U1174 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[61]), .Z(n598));
Q_AN02 U1175 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[60]), .Z(n599));
Q_AN02 U1176 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[59]), .Z(n600));
Q_AN02 U1177 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[58]), .Z(n601));
Q_AN02 U1178 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[57]), .Z(n602));
Q_AN02 U1179 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[56]), .Z(n603));
Q_AN02 U1180 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[55]), .Z(n604));
Q_AN02 U1181 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[54]), .Z(n605));
Q_AN02 U1182 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[53]), .Z(n606));
Q_AN02 U1183 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[52]), .Z(n607));
Q_AN02 U1184 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[51]), .Z(n608));
Q_AN02 U1185 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[50]), .Z(n609));
Q_AN02 U1186 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[49]), .Z(n610));
Q_AN02 U1187 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[48]), .Z(n611));
Q_AN02 U1188 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[47]), .Z(n612));
Q_AN02 U1189 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[46]), .Z(n613));
Q_AN02 U1190 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[45]), .Z(n614));
Q_AN02 U1191 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[44]), .Z(n615));
Q_AN02 U1192 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[43]), .Z(n616));
Q_AN02 U1193 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[42]), .Z(n617));
Q_AN02 U1194 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[41]), .Z(n618));
Q_AN02 U1195 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[40]), .Z(n619));
Q_AN02 U1196 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[39]), .Z(n620));
Q_AN02 U1197 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[38]), .Z(n621));
Q_AN02 U1198 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[37]), .Z(n622));
Q_AN02 U1199 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[36]), .Z(n623));
Q_AN02 U1200 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[35]), .Z(n624));
Q_AN02 U1201 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[34]), .Z(n625));
Q_AN02 U1202 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[33]), .Z(n626));
Q_AN02 U1203 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[32]), .Z(n627));
Q_AN02 U1204 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[31]), .Z(n628));
Q_AN02 U1205 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[30]), .Z(n629));
Q_AN02 U1206 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[29]), .Z(n630));
Q_AN02 U1207 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[28]), .Z(n631));
Q_AN02 U1208 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[27]), .Z(n632));
Q_AN02 U1209 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[26]), .Z(n633));
Q_AN02 U1210 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[25]), .Z(n634));
Q_AN02 U1211 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[24]), .Z(n635));
Q_AN02 U1212 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[23]), .Z(n636));
Q_AN02 U1213 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[22]), .Z(n637));
Q_AN02 U1214 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[21]), .Z(n638));
Q_AN02 U1215 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[20]), .Z(n639));
Q_AN02 U1216 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[19]), .Z(n640));
Q_AN02 U1217 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[18]), .Z(n641));
Q_AN02 U1218 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[17]), .Z(n642));
Q_AN02 U1219 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[16]), .Z(n643));
Q_AN02 U1220 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[15]), .Z(n644));
Q_AN02 U1221 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[14]), .Z(n645));
Q_AN02 U1222 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[13]), .Z(n646));
Q_AN02 U1223 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[12]), .Z(n647));
Q_AN02 U1224 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[11]), .Z(n648));
Q_AN02 U1225 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[10]), .Z(n649));
Q_AN02 U1226 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[9]), .Z(n650));
Q_AN02 U1227 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[8]), .Z(n651));
Q_AN02 U1228 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[7]), .Z(n652));
Q_AN02 U1229 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[6]), .Z(n653));
Q_AN02 U1230 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[5]), .Z(n654));
Q_AN02 U1231 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[4]), .Z(n655));
Q_AN02 U1232 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[3]), .Z(n656));
Q_AN02 U1233 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[2]), .Z(n657));
Q_AN02 U1234 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[1]), .Z(n658));
Q_AN02 U1235 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[0]), .Z(n659));
Q_AO21 U1236 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[82]), .B0(n577), .Z(n493));
Q_AO21 U1237 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[81]), .B0(n578), .Z(n494));
Q_AO21 U1238 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[80]), .B0(n579), .Z(n495));
Q_AO21 U1239 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[79]), .B0(n580), .Z(n496));
Q_AO21 U1240 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[78]), .B0(n581), .Z(n497));
Q_AO21 U1241 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[77]), .B0(n582), .Z(n498));
Q_AO21 U1242 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[76]), .B0(n583), .Z(n499));
Q_AO21 U1243 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[75]), .B0(n584), .Z(n500));
Q_AO21 U1244 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[74]), .B0(n585), .Z(n501));
Q_AO21 U1245 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[73]), .B0(n586), .Z(n502));
Q_AO21 U1246 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[72]), .B0(n587), .Z(n503));
Q_AO21 U1247 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[71]), .B0(n588), .Z(n504));
Q_AO21 U1248 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[70]), .B0(n589), .Z(n505));
Q_AO21 U1249 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[69]), .B0(n590), .Z(n506));
Q_AO21 U1250 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[68]), .B0(n591), .Z(n507));
Q_AO21 U1251 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[67]), .B0(n592), .Z(n508));
Q_AO21 U1252 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[66]), .B0(n593), .Z(n509));
Q_AO21 U1253 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[65]), .B0(n594), .Z(n510));
Q_AO21 U1254 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[64]), .B0(n595), .Z(n511));
Q_AO21 U1255 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[63]), .B0(n596), .Z(n512));
Q_AO21 U1256 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[62]), .B0(n597), .Z(n513));
Q_AO21 U1257 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[61]), .B0(n598), .Z(n514));
Q_AO21 U1258 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[60]), .B0(n599), .Z(n515));
Q_AO21 U1259 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[59]), .B0(n600), .Z(n516));
Q_AO21 U1260 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[58]), .B0(n601), .Z(n517));
Q_AO21 U1261 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[57]), .B0(n602), .Z(n518));
Q_AO21 U1262 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[56]), .B0(n603), .Z(n519));
Q_AO21 U1263 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[55]), .B0(n604), .Z(n520));
Q_AO21 U1264 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[54]), .B0(n605), .Z(n521));
Q_AO21 U1265 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[53]), .B0(n606), .Z(n522));
Q_AO21 U1266 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[52]), .B0(n607), .Z(n523));
Q_AO21 U1267 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[51]), .B0(n608), .Z(n524));
Q_AO21 U1268 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[50]), .B0(n609), .Z(n525));
Q_AO21 U1269 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[49]), .B0(n610), .Z(n526));
Q_AO21 U1270 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[48]), .B0(n611), .Z(n527));
Q_AO21 U1271 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[47]), .B0(n612), .Z(n528));
Q_AO21 U1272 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[46]), .B0(n613), .Z(n529));
Q_AO21 U1273 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[45]), .B0(n614), .Z(n530));
Q_AO21 U1274 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[44]), .B0(n615), .Z(n531));
Q_AO21 U1275 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[43]), .B0(n616), .Z(n532));
Q_AO21 U1276 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[42]), .B0(n617), .Z(n533));
Q_AO21 U1277 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[41]), .B0(n618), .Z(n534));
Q_AO21 U1278 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[40]), .B0(n619), .Z(n535));
Q_AO21 U1279 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[39]), .B0(n620), .Z(n536));
Q_AO21 U1280 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[38]), .B0(n621), .Z(n537));
Q_AO21 U1281 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[37]), .B0(n622), .Z(n538));
Q_AO21 U1282 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[36]), .B0(n623), .Z(n539));
Q_AO21 U1283 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[35]), .B0(n624), .Z(n540));
Q_AO21 U1284 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[34]), .B0(n625), .Z(n541));
Q_AO21 U1285 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[33]), .B0(n626), .Z(n542));
Q_AO21 U1286 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[32]), .B0(n627), .Z(n543));
Q_AO21 U1287 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[31]), .B0(n628), .Z(n544));
Q_AO21 U1288 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[30]), .B0(n629), .Z(n545));
Q_AO21 U1289 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[29]), .B0(n630), .Z(n546));
Q_AO21 U1290 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[28]), .B0(n631), .Z(n547));
Q_AO21 U1291 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[27]), .B0(n632), .Z(n548));
Q_AO21 U1292 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[26]), .B0(n633), .Z(n549));
Q_AO21 U1293 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[25]), .B0(n634), .Z(n550));
Q_AO21 U1294 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[24]), .B0(n635), .Z(n551));
Q_AO21 U1295 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[23]), .B0(n636), .Z(n552));
Q_AO21 U1296 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[22]), .B0(n637), .Z(n553));
Q_AO21 U1297 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[21]), .B0(n638), .Z(n554));
Q_AO21 U1298 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[20]), .B0(n639), .Z(n555));
Q_AO21 U1299 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[19]), .B0(n640), .Z(n556));
Q_AO21 U1300 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[18]), .B0(n641), .Z(n557));
Q_AO21 U1301 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[17]), .B0(n642), .Z(n558));
Q_AO21 U1302 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[16]), .B0(n643), .Z(n559));
Q_AO21 U1303 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[15]), .B0(n644), .Z(n560));
Q_AO21 U1304 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[14]), .B0(n645), .Z(n561));
Q_AO21 U1305 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[13]), .B0(n646), .Z(n562));
Q_AO21 U1306 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[12]), .B0(n647), .Z(n563));
Q_AO21 U1307 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[11]), .B0(n648), .Z(n564));
Q_AO21 U1308 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[10]), .B0(n649), .Z(n565));
Q_AO21 U1309 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[9]), .B0(n650), .Z(n566));
Q_AO21 U1310 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[8]), .B0(n651), .Z(n567));
Q_AO21 U1311 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[7]), .B0(n652), .Z(n568));
Q_AO21 U1312 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[6]), .B0(n653), .Z(n569));
Q_AO21 U1313 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[5]), .B0(n654), .Z(n570));
Q_AO21 U1314 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[4]), .B0(n655), .Z(n571));
Q_AO21 U1315 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[3]), .B0(n656), .Z(n572));
Q_AO21 U1316 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[2]), .B0(n657), .Z(n573));
Q_AO21 U1317 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[1]), .B0(n658), .Z(n574));
Q_AO21 U1318 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[0]), .B0(n659), .Z(n575));
Q_AN02 U1319 ( .A0(prefetch_lden_mem[0]), .A1(mem_ecc_error), .Z(n743));
Q_AN02 U1320 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[82]), .Z(n744));
Q_AN02 U1321 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[81]), .Z(n745));
Q_AN02 U1322 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[80]), .Z(n746));
Q_AN02 U1323 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[79]), .Z(n747));
Q_AN02 U1324 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[78]), .Z(n748));
Q_AN02 U1325 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[77]), .Z(n749));
Q_AN02 U1326 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[76]), .Z(n750));
Q_AN02 U1327 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[75]), .Z(n751));
Q_AN02 U1328 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[74]), .Z(n752));
Q_AN02 U1329 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[73]), .Z(n753));
Q_AN02 U1330 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[72]), .Z(n754));
Q_AN02 U1331 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[71]), .Z(n755));
Q_AN02 U1332 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[70]), .Z(n756));
Q_AN02 U1333 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[69]), .Z(n757));
Q_AN02 U1334 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[68]), .Z(n758));
Q_AN02 U1335 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[67]), .Z(n759));
Q_AN02 U1336 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[66]), .Z(n760));
Q_AN02 U1337 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[65]), .Z(n761));
Q_AN02 U1338 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[64]), .Z(n762));
Q_AN02 U1339 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[63]), .Z(n763));
Q_AN02 U1340 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[62]), .Z(n764));
Q_AN02 U1341 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[61]), .Z(n765));
Q_AN02 U1342 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[60]), .Z(n766));
Q_AN02 U1343 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[59]), .Z(n767));
Q_AN02 U1344 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[58]), .Z(n768));
Q_AN02 U1345 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[57]), .Z(n769));
Q_AN02 U1346 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[56]), .Z(n770));
Q_AN02 U1347 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[55]), .Z(n771));
Q_AN02 U1348 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[54]), .Z(n772));
Q_AN02 U1349 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[53]), .Z(n773));
Q_AN02 U1350 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[52]), .Z(n774));
Q_AN02 U1351 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[51]), .Z(n775));
Q_AN02 U1352 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[50]), .Z(n776));
Q_AN02 U1353 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[49]), .Z(n777));
Q_AN02 U1354 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[48]), .Z(n778));
Q_AN02 U1355 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[47]), .Z(n779));
Q_AN02 U1356 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[46]), .Z(n780));
Q_AN02 U1357 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[45]), .Z(n781));
Q_AN02 U1358 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[44]), .Z(n782));
Q_AN02 U1359 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[43]), .Z(n783));
Q_AN02 U1360 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[42]), .Z(n784));
Q_AN02 U1361 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[41]), .Z(n785));
Q_AN02 U1362 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[40]), .Z(n786));
Q_AN02 U1363 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[39]), .Z(n787));
Q_AN02 U1364 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[38]), .Z(n788));
Q_AN02 U1365 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[37]), .Z(n789));
Q_AN02 U1366 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[36]), .Z(n790));
Q_AN02 U1367 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[35]), .Z(n791));
Q_AN02 U1368 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[34]), .Z(n792));
Q_AN02 U1369 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[33]), .Z(n793));
Q_AN02 U1370 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[32]), .Z(n794));
Q_AN02 U1371 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[31]), .Z(n795));
Q_AN02 U1372 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[30]), .Z(n796));
Q_AN02 U1373 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[29]), .Z(n797));
Q_AN02 U1374 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[28]), .Z(n798));
Q_AN02 U1375 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[27]), .Z(n799));
Q_AN02 U1376 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[26]), .Z(n800));
Q_AN02 U1377 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[25]), .Z(n801));
Q_AN02 U1378 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[24]), .Z(n802));
Q_AN02 U1379 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[23]), .Z(n803));
Q_AN02 U1380 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[22]), .Z(n804));
Q_AN02 U1381 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[21]), .Z(n805));
Q_AN02 U1382 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[20]), .Z(n806));
Q_AN02 U1383 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[19]), .Z(n807));
Q_AN02 U1384 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[18]), .Z(n808));
Q_AN02 U1385 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[17]), .Z(n809));
Q_AN02 U1386 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[16]), .Z(n810));
Q_AN02 U1387 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[15]), .Z(n811));
Q_AN02 U1388 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[14]), .Z(n812));
Q_AN02 U1389 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[13]), .Z(n813));
Q_AN02 U1390 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[12]), .Z(n814));
Q_AN02 U1391 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[11]), .Z(n815));
Q_AN02 U1392 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[10]), .Z(n816));
Q_AN02 U1393 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[9]), .Z(n817));
Q_AN02 U1394 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[8]), .Z(n818));
Q_AN02 U1395 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[7]), .Z(n819));
Q_AN02 U1396 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[6]), .Z(n820));
Q_AN02 U1397 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[5]), .Z(n821));
Q_AN02 U1398 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[4]), .Z(n822));
Q_AN02 U1399 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[3]), .Z(n823));
Q_AN02 U1400 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[2]), .Z(n824));
Q_AN02 U1401 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[1]), .Z(n825));
Q_AN02 U1402 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[0]), .Z(n826));
Q_AO21 U1403 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[82]), .B0(n744), .Z(n660));
Q_AO21 U1404 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[81]), .B0(n745), .Z(n661));
Q_AO21 U1405 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[80]), .B0(n746), .Z(n662));
Q_AO21 U1406 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[79]), .B0(n747), .Z(n663));
Q_AO21 U1407 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[78]), .B0(n748), .Z(n664));
Q_AO21 U1408 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[77]), .B0(n749), .Z(n665));
Q_AO21 U1409 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[76]), .B0(n750), .Z(n666));
Q_AO21 U1410 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[75]), .B0(n751), .Z(n667));
Q_AO21 U1411 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[74]), .B0(n752), .Z(n668));
Q_AO21 U1412 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[73]), .B0(n753), .Z(n669));
Q_AO21 U1413 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[72]), .B0(n754), .Z(n670));
Q_AO21 U1414 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[71]), .B0(n755), .Z(n671));
Q_AO21 U1415 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[70]), .B0(n756), .Z(n672));
Q_AO21 U1416 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[69]), .B0(n757), .Z(n673));
Q_AO21 U1417 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[68]), .B0(n758), .Z(n674));
Q_AO21 U1418 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[67]), .B0(n759), .Z(n675));
Q_AO21 U1419 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[66]), .B0(n760), .Z(n676));
Q_AO21 U1420 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[65]), .B0(n761), .Z(n677));
Q_AO21 U1421 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[64]), .B0(n762), .Z(n678));
Q_AO21 U1422 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[63]), .B0(n763), .Z(n679));
Q_AO21 U1423 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[62]), .B0(n764), .Z(n680));
Q_AO21 U1424 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[61]), .B0(n765), .Z(n681));
Q_AO21 U1425 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[60]), .B0(n766), .Z(n682));
Q_AO21 U1426 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[59]), .B0(n767), .Z(n683));
Q_AO21 U1427 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[58]), .B0(n768), .Z(n684));
Q_AO21 U1428 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[57]), .B0(n769), .Z(n685));
Q_AO21 U1429 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[56]), .B0(n770), .Z(n686));
Q_AO21 U1430 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[55]), .B0(n771), .Z(n687));
Q_AO21 U1431 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[54]), .B0(n772), .Z(n688));
Q_AO21 U1432 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[53]), .B0(n773), .Z(n689));
Q_AO21 U1433 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[52]), .B0(n774), .Z(n690));
Q_AO21 U1434 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[51]), .B0(n775), .Z(n691));
Q_AO21 U1435 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[50]), .B0(n776), .Z(n692));
Q_AO21 U1436 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[49]), .B0(n777), .Z(n693));
Q_AO21 U1437 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[48]), .B0(n778), .Z(n694));
Q_AO21 U1438 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[47]), .B0(n779), .Z(n695));
Q_AO21 U1439 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[46]), .B0(n780), .Z(n696));
Q_AO21 U1440 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[45]), .B0(n781), .Z(n697));
Q_AO21 U1441 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[44]), .B0(n782), .Z(n698));
Q_AO21 U1442 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[43]), .B0(n783), .Z(n699));
Q_AO21 U1443 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[42]), .B0(n784), .Z(n700));
Q_AO21 U1444 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[41]), .B0(n785), .Z(n701));
Q_AO21 U1445 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[40]), .B0(n786), .Z(n702));
Q_AO21 U1446 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[39]), .B0(n787), .Z(n703));
Q_AO21 U1447 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[38]), .B0(n788), .Z(n704));
Q_AO21 U1448 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[37]), .B0(n789), .Z(n705));
Q_AO21 U1449 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[36]), .B0(n790), .Z(n706));
Q_AO21 U1450 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[35]), .B0(n791), .Z(n707));
Q_AO21 U1451 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[34]), .B0(n792), .Z(n708));
Q_AO21 U1452 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[33]), .B0(n793), .Z(n709));
Q_AO21 U1453 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[32]), .B0(n794), .Z(n710));
Q_AO21 U1454 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[31]), .B0(n795), .Z(n711));
Q_AO21 U1455 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[30]), .B0(n796), .Z(n712));
Q_AO21 U1456 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[29]), .B0(n797), .Z(n713));
Q_AO21 U1457 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[28]), .B0(n798), .Z(n714));
Q_AO21 U1458 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[27]), .B0(n799), .Z(n715));
Q_AO21 U1459 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[26]), .B0(n800), .Z(n716));
Q_AO21 U1460 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[25]), .B0(n801), .Z(n717));
Q_AO21 U1461 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[24]), .B0(n802), .Z(n718));
Q_AO21 U1462 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[23]), .B0(n803), .Z(n719));
Q_AO21 U1463 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[22]), .B0(n804), .Z(n720));
Q_AO21 U1464 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[21]), .B0(n805), .Z(n721));
Q_AO21 U1465 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[20]), .B0(n806), .Z(n722));
Q_AO21 U1466 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[19]), .B0(n807), .Z(n723));
Q_AO21 U1467 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[18]), .B0(n808), .Z(n724));
Q_AO21 U1468 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[17]), .B0(n809), .Z(n725));
Q_AO21 U1469 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[16]), .B0(n810), .Z(n726));
Q_AO21 U1470 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[15]), .B0(n811), .Z(n727));
Q_AO21 U1471 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[14]), .B0(n812), .Z(n728));
Q_AO21 U1472 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[13]), .B0(n813), .Z(n729));
Q_AO21 U1473 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[12]), .B0(n814), .Z(n730));
Q_AO21 U1474 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[11]), .B0(n815), .Z(n731));
Q_AO21 U1475 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[10]), .B0(n816), .Z(n732));
Q_AO21 U1476 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[9]), .B0(n817), .Z(n733));
Q_AO21 U1477 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[8]), .B0(n818), .Z(n734));
Q_AO21 U1478 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[7]), .B0(n819), .Z(n735));
Q_AO21 U1479 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[6]), .B0(n820), .Z(n736));
Q_AO21 U1480 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[5]), .B0(n821), .Z(n737));
Q_AO21 U1481 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[4]), .B0(n822), .Z(n738));
Q_AO21 U1482 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[3]), .B0(n823), .Z(n739));
Q_AO21 U1483 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[2]), .B0(n824), .Z(n740));
Q_AO21 U1484 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[1]), .B0(n825), .Z(n741));
Q_AO21 U1485 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[0]), .B0(n826), .Z(n742));
Q_OR02 U1486 ( .A0(prefetch_lden_bypass[2]), .A1(prefetch_lden_mem[2]), .Z(n105));
Q_OR02 U1487 ( .A0(prefetch_lden_bypass[1]), .A1(prefetch_lden_mem[1]), .Z(n104));
Q_OR02 U1488 ( .A0(prefetch_lden_bypass[0]), .A1(prefetch_lden_mem[0]), .Z(n103));
Q_AN02 U1489 ( .A0(n109), .A1(\c_mem_prefetch_wptr_dly[0][2] ), .Z(prefetch_lden_bypass[2]));
Q_AN02 U1490 ( .A0(n109), .A1(\c_mem_prefetch_wptr_dly[0][1] ), .Z(prefetch_lden_bypass[1]));
Q_AN02 U1491 ( .A0(n109), .A1(\c_mem_prefetch_wptr_dly[0][0] ), .Z(prefetch_lden_bypass[0]));
Q_AN02 U1492 ( .A0(n149), .A1(n827), .Z(prefetch_lden_mem[2]));
Q_AN02 U1493 ( .A0(n149), .A1(n828), .Z(prefetch_lden_mem[1]));
Q_AN02 U1494 ( .A0(n149), .A1(n829), .Z(prefetch_lden_mem[0]));
Q_MX03 U1495 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(n829), .A1(n828), .A2(n827), .Z(n87));
Q_AN02 U1496 ( .A0(r_mem_ren_dly[2]), .A1(\r_mem_prefetch_wptr_dly[2][2] ), .Z(n827));
Q_AN02 U1497 ( .A0(r_mem_ren_dly[2]), .A1(\r_mem_prefetch_wptr_dly[2][1] ), .Z(n828));
Q_AN02 U1498 ( .A0(r_mem_ren_dly[2]), .A1(\r_mem_prefetch_wptr_dly[2][0] ), .Z(n829));
Q_AN02 U1499 ( .A0(n110), .A1(r_prefetch_full), .Z(n86));
Q_ND02 U1500 ( .A0(n831), .A1(n830), .Z(n89));
Q_AN03 U1501 ( .A0(r_mem_wptr[1]), .A1(r_mem_wptr[0]), .A2(n832), .Z(n830));
Q_AN03 U1502 ( .A0(n834), .A1(n835), .A2(r_mem_wptr[2]), .Z(n831));
Q_AN03 U1503 ( .A0(r_mem_wptr[7]), .A1(n833), .A2(r_mem_wptr[5]), .Z(n832));
Q_ND02 U1504 ( .A0(n837), .A1(n836), .Z(n90));
Q_AN03 U1505 ( .A0(r_mem_rptr[1]), .A1(r_mem_rptr[0]), .A2(n838), .Z(n836));
Q_AN03 U1506 ( .A0(n840), .A1(n841), .A2(r_mem_rptr[2]), .Z(n837));
Q_AN03 U1507 ( .A0(r_mem_rptr[7]), .A1(n839), .A2(r_mem_rptr[5]), .Z(n838));
Q_AN02 U1508 ( .A0(n842), .A1(r_prefetch_rptr[1]), .Z(n91));
Q_INV U1509 ( .A(_zy_sva_sf1hot_0), .Z(n844));
Q_AN02 U1510 ( .A0(rst_n), .A1(n844), .Z(n843));
ixc_assign_8 _zz_strnp_0 ( used_slots[7:0], r_used_slots[7:0]);
ixc_assign_8 _zz_strnp_1 ( free_slots[7:0], r_free_slots[7:0]);
ixc_assign_8 _zz_strnp_2 ( mem_waddr[7:0], r_mem_wptr[7:0]);
ixc_assign_8 _zz_strnp_3 ( mem_raddr[7:0], r_mem_rptr[7:0]);
ixc_assign_83 _zz_strnp_4 ( mem_wdata[82:0], wdata[82:0]);
ixc_assign _zz_strnp_5 ( empty, r_prefetch_empty);
ixc_assign _zz_strnp_6 ( full, r_mem_full);
ixc_assign _zz_strnp_7 ( _zy_simnet_mem_wen_0_w$, mem_wen);
ixc_assign_8 _zz_strnp_8 ( _zy_simnet_mem_waddr_1_w$[0:7], mem_waddr[7:0]);
ixc_assign_83 _zz_strnp_9 ( _zy_simnet_mem_wdata_2_w$[0:82], mem_wdata[82:0]);
ixc_assign _zz_strnp_10 ( _zy_simnet_mem_ren_3_w$, mem_ren);
ixc_assign_8 _zz_strnp_11 ( _zy_simnet_mem_raddr_4_w$[0:7], mem_raddr[7:0]);
ixc_assign _zz_strnp_12 ( _zy_simnet_empty_5_w$, empty);
ixc_assign _zz_strnp_13 ( _zy_simnet_full_6_w$, full);
ixc_assign_8 _zz_strnp_14 ( _zy_simnet_used_slots_7_w$[0:7], used_slots[7:0]);
ixc_assign_8 _zz_strnp_15 ( _zy_simnet_free_slots_8_w$[0:7], free_slots[7:0]);
ixc_assign _zz_strnp_16 ( _zy_simnet_rerr_9_w$, rerr);
ixc_assign_83 _zz_strnp_17 ( _zy_simnet_rdata_10_w$[0:82], rdata[82:0]);
ixc_assign _zz_strnp_18 ( _zy_simnet_underflow_11_w$, underflow);
ixc_assign _zz_strnp_19 ( _zy_simnet_overflow_12_w$, overflow);
Q_INV U1531 ( .A(rst_n), .Z(_zy_sva__asrtLbl279_1_reset_or));
Q_AO21 U1532 ( .A0(_zy_sva_b0[1]), .A1(_zy_sva_b0[2]), .B0(n851), .Z(n850));
Q_XOR2 U1533 ( .A0(_zy_sva_b0[1]), .A1(_zy_sva_b0[2]), .Z(n852));
Q_AN02 U1534 ( .A0(_zy_sva_b0[0]), .A1(n852), .Z(n851));
Q_XOR2 U1535 ( .A0(_zy_sva_b0[0]), .A1(n852), .Z(n849));
Q_INV U1536 ( .A(n850), .Z(n848));
Q_AN02 U1537 ( .A0(n848), .A1(n849), .Z(_zy_sva_sf1hot_0));
ixc_sample_logic_3_3 _zz_zy_sva_b0 ( _zy_sva_b0[2:0], { 
	\c_mem_prefetch_wptr_dly[0][2] , \c_mem_prefetch_wptr_dly[0][1] , 
	\c_mem_prefetch_wptr_dly[0][0] });
ixc_pio_call_0_0_0_0_1 _zzixc_tfport_1_0 ( _zyixc_port_1_0_ack, 
	_zyixc_port_1_0_s2hW, _zyixc_port_1_0_isf, _zyixc_port_1_0_req, n847, 
	_zyixc_port_1_0_osf, n846, n1);
wire [2:0] n855 = 3'b000;
Q_ASSERT _asrtLbl279 ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT( ), .FAIL_COUNT( ), .CHECK_COUNT( ), .KILL_SIGNAL( ), .SEVERITY(n855[0]));
// pragma CVASTRPROP INSTANCE "_asrtLbl279" HDL_ASSERT "$"
// pragma CVASTRPROP INSTANCE "_asrtLbl279" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/common/nx_library/nx_fifo_ctrl_ram_1r1w.v"
//pragma CVAINTPROP INSTANCE "_asrtLbl279" ASSERT_LINE 279
Q_AN02 U1541 ( .A0(r_free_slots[1]), .A1(r_free_slots[0]), .Z(n323));
Q_AN02 U1542 ( .A0(r_used_slots[1]), .A1(r_used_slots[0]), .Z(n310));
Q_XOR2 U1543 ( .A0(mem_ren), .A1(r_mem_rptr[0]), .Z(n213));
Q_XNR2 U1544 ( .A0(n133), .A1(n191), .Z(n189));
Q_XNR2 U1545 ( .A0(n114), .A1(n298), .Z(n166));
Q_XOR2 U1546 ( .A0(n147), .A1(n141), .Z(n112));
Q_INV U1547 ( .A(_zy_sva__asrtLbl279_1_1_fail[0]), .Z(n853));
Q_FDP4EP \_zy_sva__asrtLbl279_1_1_fail_REG[0] ( .CK(clk), .CE(n843), .R(n845), .D(n853), .Q(_zy_sva__asrtLbl279_1_1_fail[0]));
Q_INV U1549 ( .A(_zyixc_port_1_0_req), .Z(n854));
Q_FDP4EP _zyixc_port_1_0_req_REG  ( .CK(clk), .CE(n843), .R(n845), .D(n854), .Q(_zyixc_port_1_0_req));
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m1 "r_mem_prefetch_wptr_dly 1 2 0 2 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m2 "c_mem_prefetch_wptr_dly 1 2 0 2 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m3 "r_prefetch_data 1 83 0 2 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m4 "c_prefetch_data 1 83 0 2 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_NON_CMM "4"
// pragma CVASTRPROP MODULE HDLICE PROP_RANOFF TRUE
endmodule
