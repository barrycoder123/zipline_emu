architecture module of ixc_gfifo_bind_20_2 is

begin
end module;
