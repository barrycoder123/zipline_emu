
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
(* celldefine = 1 *) 
module nx_indirect_access_cntrl_v2_xcm125 ( clk, rst_n, wr_stb, reg_addr, 
	cmnd_op, cmnd_addr, cmnd_table_id, stat_code, stat_datawords, 
	stat_addr, stat_table_id, capability_lst, capability_type, enable, 
	.addr_limit( {\addr_limit[0][13] , \addr_limit[0][12] , 
	\addr_limit[0][11] , \addr_limit[0][10] , \addr_limit[0][9] , 
	\addr_limit[0][8] , \addr_limit[0][7] , \addr_limit[0][6] , 
	\addr_limit[0][5] , \addr_limit[0][4] , \addr_limit[0][3] , 
	\addr_limit[0][2] , \addr_limit[0][1] , \addr_limit[0][0] } ), 
	wr_dat, rd_dat, sw_cs, sw_ce, sw_we, sw_add, sw_wdat, sw_rdat, 
	sw_match, sw_aindex, grant, rsp, yield, reset);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
input clk;
input rst_n;
input wr_stb;
input [10:0] reg_addr;
input [3:0] cmnd_op;
input [13:0] cmnd_addr;
input [0:0] cmnd_table_id;
output [2:0] stat_code;
output [4:0] stat_datawords;
output [13:0] stat_addr;
output [0:0] stat_table_id;
output [15:0] capability_lst;
output [3:0] capability_type;
output enable;
input \addr_limit[0][13] ;
input \addr_limit[0][12] ;
input \addr_limit[0][11] ;
input \addr_limit[0][10] ;
input \addr_limit[0][9] ;
input \addr_limit[0][8] ;
input \addr_limit[0][7] ;
input \addr_limit[0][6] ;
input \addr_limit[0][5] ;
input \addr_limit[0][4] ;
input \addr_limit[0][3] ;
input \addr_limit[0][2] ;
input \addr_limit[0][1] ;
input \addr_limit[0][0] ;
input [37:0] wr_dat;
output [37:0] rd_dat;
output sw_cs;
output sw_ce;
output sw_we;
output [13:0] sw_add;
output [37:0] sw_wdat;
input [37:0] sw_rdat;
input sw_match;
input [12:0] sw_aindex;
input grant;
input rsp;
output yield;
output reset;
wire [0:2] _zy_simnet_stat_code_0_w$;
wire [0:4] _zy_simnet_stat_datawords_1_w$;
wire [0:13] _zy_simnet_stat_addr_2_w$;
wire _zy_simnet_stat_table_id_3_w$;
wire [0:15] _zy_simnet_capability_lst_4_w$;
wire [0:3] _zy_simnet_capability_type_5_w$;
wire _zy_simnet_enable_6_w$;
wire [0:37] _zy_simnet_rd_dat_7_w$;
wire _zy_simnet_sw_cs_8_w$;
wire _zy_simnet_sw_ce_9_w$;
wire _zy_simnet_sw_we_10_w$;
wire [0:13] _zy_simnet_sw_add_11_w$;
wire [0:37] _zy_simnet_sw_wdat_12_w$;
wire _zy_simnet_yield_13_w$;
wire _zy_simnet_reset_14_w$;
wire [3:0] cmnd;
wire init_r;
wire [0:0] inc_r;
wire init_inc_r;
wire sw_cs_r;
wire sw_ce_r;
wire rst_r;
wire rst_or_ini_r;
wire [13:0] rst_addr_r;
wire sw_we_r;
wire cmnd_rd_stb;
wire cmnd_wr_stb;
wire cmnd_ena_stb;
wire cmnd_dis_stb;
wire cmnd_rst_stb;
wire cmnd_ini_stb;
wire cmnd_inc_stb;
wire cmnd_sis_stb;
wire cmnd_tmo_stb;
wire cmnd_cmp_stb;
wire cmnd_issued;
wire ack_error;
wire unsupported_op;
wire [3:0] state_r;
wire [5:0] timer_r;
wire timeout;
wire sim_tmo_r;
wire [13:0] maxaddr;
wire badaddr;
wire igrant;
wire [2:0] stat;
supply0 n1;
supply1 n2;
Q_BUF U0 ( .A(n2), .Z(stat_datawords[0]));
Q_BUF U1 ( .A(n1), .Z(stat_datawords[1]));
Q_BUF U2 ( .A(n1), .Z(stat_datawords[2]));
Q_BUF U3 ( .A(n1), .Z(stat_datawords[3]));
Q_BUF U4 ( .A(n1), .Z(stat_datawords[4]));
Q_BUF U5 ( .A(n1), .Z(capability_type[0]));
Q_BUF U6 ( .A(n1), .Z(capability_type[1]));
Q_BUF U7 ( .A(n1), .Z(capability_type[2]));
Q_BUF U8 ( .A(n1), .Z(capability_type[3]));
Q_BUF U9 ( .A(n2), .Z(capability_lst[0]));
Q_BUF U10 ( .A(n2), .Z(capability_lst[1]));
Q_BUF U11 ( .A(n2), .Z(capability_lst[2]));
Q_BUF U12 ( .A(n2), .Z(capability_lst[3]));
Q_BUF U13 ( .A(n2), .Z(capability_lst[4]));
Q_BUF U14 ( .A(n2), .Z(capability_lst[5]));
Q_BUF U15 ( .A(n2), .Z(capability_lst[6]));
Q_BUF U16 ( .A(n1), .Z(capability_lst[7]));
Q_BUF U17 ( .A(n2), .Z(capability_lst[8]));
Q_BUF U18 ( .A(n1), .Z(capability_lst[9]));
Q_BUF U19 ( .A(n1), .Z(capability_lst[10]));
Q_BUF U20 ( .A(n1), .Z(capability_lst[11]));
Q_BUF U21 ( .A(n1), .Z(capability_lst[12]));
Q_BUF U22 ( .A(n1), .Z(capability_lst[13]));
Q_BUF U23 ( .A(n2), .Z(capability_lst[14]));
Q_BUF U24 ( .A(n2), .Z(capability_lst[15]));
Q_BUF U25 ( .A(n1), .Z(stat_table_id[0]));
ixc_assign_3 _zz_strnp_7 ( stat[2:0], stat_code[2:0]);
ixc_assign_4 _zz_strnp_1 ( cmnd[3:0], cmnd_op[3:0]);
ixc_assign \genblk1._zz_strnp_0 ( reset, rst_or_ini_r);
ixc_context_read_6 _zzixc_ctxrd_0 ( { stat_code[2], stat_code[1], 
	stat_code[0], stat[2], stat[1], stat[0]});
ixc_assign _zz_strnp_22 ( _zy_simnet_reset_14_w$, reset);
ixc_assign _zz_strnp_21 ( _zy_simnet_yield_13_w$, yield);
ixc_assign_38 _zz_strnp_20 ( _zy_simnet_sw_wdat_12_w$[0:37], sw_wdat[37:0]);
ixc_assign_14 _zz_strnp_19 ( _zy_simnet_sw_add_11_w$[0:13], sw_add[13:0]);
ixc_assign _zz_strnp_18 ( _zy_simnet_sw_we_10_w$, sw_we);
ixc_assign _zz_strnp_17 ( _zy_simnet_sw_ce_9_w$, sw_ce);
ixc_assign _zz_strnp_16 ( _zy_simnet_sw_cs_8_w$, sw_cs);
ixc_assign_38 _zz_strnp_15 ( _zy_simnet_rd_dat_7_w$[0:37], rd_dat[37:0]);
ixc_assign _zz_strnp_14 ( _zy_simnet_enable_6_w$, enable);
ixc_assign_4 _zz_strnp_13 ( _zy_simnet_capability_type_5_w$[0:3], { n1, n1, 
	n1, n1});
ixc_assign_16 _zz_strnp_12 ( _zy_simnet_capability_lst_4_w$[0:15], { n2, n2, 
	n1, n1, n1, n1, n1, n2, n1, n2, n2, n2, n2, n2, n2, n2});
ixc_assign _zz_strnp_11 ( _zy_simnet_stat_table_id_3_w$, n1);
ixc_assign_14 _zz_strnp_10 ( _zy_simnet_stat_addr_2_w$[0:13], stat_addr[13:0]);
ixc_assign_5 _zz_strnp_9 ( _zy_simnet_stat_datawords_1_w$[0:4], { n1, n1, n1, 
	n1, n2});
ixc_assign_3 _zz_strnp_8 ( _zy_simnet_stat_code_0_w$[0:2], stat_code[2:0]);
ixc_assign_14 _zz_strnp_6 ( stat_addr[13:0], maxaddr[13:0]);
Q_AN02 U46 ( .A0(n54), .A1(grant), .Z(igrant));
Q_OA21 U47 ( .A0(n53), .A1(n52), .B0(cmnd_issued), .Z(badaddr));
Q_AO21 U48 ( .A0(n17), .A1(n29), .B0(n16), .Z(n53));
Q_AO21 U49 ( .A0(n50), .A1(n42), .B0(n51), .Z(n52));
Q_AN03 U50 ( .A0(n50), .A1(n43), .A2(n49), .Z(n51));
Q_AN02 U51 ( .A0(n17), .A1(n30), .Z(n50));
Q_AO21 U52 ( .A0(n46), .A1(n48), .B0(n45), .Z(n49));
Q_AN02 U53 ( .A0(cmnd_addr[0]), .A1(n47), .Z(n48));
Q_INV U54 ( .A(maxaddr[0]), .Z(n47));
Q_OR02 U55 ( .A0(cmnd_addr[1]), .A1(n44), .Z(n46));
Q_AN02 U56 ( .A0(cmnd_addr[1]), .A1(n44), .Z(n45));
Q_INV U57 ( .A(maxaddr[1]), .Z(n44));
Q_OR03 U58 ( .A0(n39), .A1(n38), .A2(n41), .Z(n42));
Q_OA21 U59 ( .A0(cmnd_addr[2]), .A1(n35), .B0(n37), .Z(n43));
Q_AN03 U60 ( .A0(cmnd_addr[2]), .A1(n35), .A2(n37), .Z(n38));
Q_INV U61 ( .A(maxaddr[2]), .Z(n35));
Q_OA21 U62 ( .A0(cmnd_addr[3]), .A1(n34), .B0(n36), .Z(n37));
Q_AN03 U63 ( .A0(cmnd_addr[3]), .A1(n34), .A2(n36), .Z(n39));
Q_INV U64 ( .A(maxaddr[3]), .Z(n34));
Q_OA21 U65 ( .A0(cmnd_addr[4]), .A1(n33), .B0(n32), .Z(n36));
Q_AN03 U66 ( .A0(cmnd_addr[4]), .A1(n33), .A2(n32), .Z(n40));
Q_INV U67 ( .A(maxaddr[4]), .Z(n33));
Q_OR02 U68 ( .A0(cmnd_addr[5]), .A1(n31), .Z(n32));
Q_AO21 U69 ( .A0(cmnd_addr[5]), .A1(n31), .B0(n40), .Z(n41));
Q_INV U70 ( .A(maxaddr[5]), .Z(n31));
Q_OR03 U71 ( .A0(n26), .A1(n25), .A2(n28), .Z(n29));
Q_OA21 U72 ( .A0(cmnd_addr[6]), .A1(n22), .B0(n24), .Z(n30));
Q_AN03 U73 ( .A0(cmnd_addr[6]), .A1(n22), .A2(n24), .Z(n25));
Q_INV U74 ( .A(maxaddr[6]), .Z(n22));
Q_OA21 U75 ( .A0(cmnd_addr[7]), .A1(n21), .B0(n23), .Z(n24));
Q_AN03 U76 ( .A0(cmnd_addr[7]), .A1(n21), .A2(n23), .Z(n26));
Q_INV U77 ( .A(maxaddr[7]), .Z(n21));
Q_OA21 U78 ( .A0(cmnd_addr[8]), .A1(n20), .B0(n19), .Z(n23));
Q_AN03 U79 ( .A0(cmnd_addr[8]), .A1(n20), .A2(n19), .Z(n27));
Q_INV U80 ( .A(maxaddr[8]), .Z(n20));
Q_OR02 U81 ( .A0(cmnd_addr[9]), .A1(n18), .Z(n19));
Q_AO21 U82 ( .A0(cmnd_addr[9]), .A1(n18), .B0(n27), .Z(n28));
Q_INV U83 ( .A(maxaddr[9]), .Z(n18));
Q_OR03 U84 ( .A0(n13), .A1(n12), .A2(n15), .Z(n16));
Q_OA21 U85 ( .A0(cmnd_addr[10]), .A1(n9), .B0(n11), .Z(n17));
Q_AN03 U86 ( .A0(cmnd_addr[10]), .A1(n9), .A2(n11), .Z(n12));
Q_INV U87 ( .A(maxaddr[10]), .Z(n9));
Q_OA21 U88 ( .A0(cmnd_addr[11]), .A1(n8), .B0(n10), .Z(n11));
Q_AN03 U89 ( .A0(cmnd_addr[11]), .A1(n8), .A2(n10), .Z(n13));
Q_INV U90 ( .A(maxaddr[11]), .Z(n8));
Q_OA21 U91 ( .A0(cmnd_addr[12]), .A1(n7), .B0(n6), .Z(n10));
Q_AN03 U92 ( .A0(cmnd_addr[12]), .A1(n7), .A2(n6), .Z(n14));
Q_INV U93 ( .A(maxaddr[12]), .Z(n7));
Q_OR02 U94 ( .A0(cmnd_addr[13]), .A1(n5), .Z(n6));
Q_AO21 U95 ( .A0(cmnd_addr[13]), .A1(n5), .B0(n14), .Z(n15));
Q_INV U96 ( .A(maxaddr[13]), .Z(n5));
Q_AN02 U97 ( .A0(n3), .A1(n4), .Z(timeout));
Q_AN03 U98 ( .A0(timer_r[2]), .A1(timer_r[1]), .A2(timer_r[0]), .Z(n4));
Q_AN03 U99 ( .A0(timer_r[5]), .A1(timer_r[4]), .A2(timer_r[3]), .Z(n3));
ixc_assign _zz_strnp_5 ( yield, timer_r[5]);
ixc_assign _zz_strnp_4 ( sw_we, sw_we_r);
ixc_assign _zz_strnp_3 ( sw_ce, sw_ce_r);
ixc_assign _zz_strnp_2 ( sw_cs, sw_cs_r);
Q_MX02 U104 ( .S(rst_or_ini_r), .A0(cmnd_addr[0]), .A1(rst_addr_r[0]), .Z(sw_add[0]));
Q_MX02 U105 ( .S(rst_or_ini_r), .A0(cmnd_addr[1]), .A1(rst_addr_r[1]), .Z(sw_add[1]));
Q_MX02 U106 ( .S(rst_or_ini_r), .A0(cmnd_addr[2]), .A1(rst_addr_r[2]), .Z(sw_add[2]));
Q_MX02 U107 ( .S(rst_or_ini_r), .A0(cmnd_addr[3]), .A1(rst_addr_r[3]), .Z(sw_add[3]));
Q_MX02 U108 ( .S(rst_or_ini_r), .A0(cmnd_addr[4]), .A1(rst_addr_r[4]), .Z(sw_add[4]));
Q_MX02 U109 ( .S(rst_or_ini_r), .A0(cmnd_addr[5]), .A1(rst_addr_r[5]), .Z(sw_add[5]));
Q_MX02 U110 ( .S(rst_or_ini_r), .A0(cmnd_addr[6]), .A1(rst_addr_r[6]), .Z(sw_add[6]));
Q_MX02 U111 ( .S(rst_or_ini_r), .A0(cmnd_addr[7]), .A1(rst_addr_r[7]), .Z(sw_add[7]));
Q_MX02 U112 ( .S(rst_or_ini_r), .A0(cmnd_addr[8]), .A1(rst_addr_r[8]), .Z(sw_add[8]));
Q_MX02 U113 ( .S(rst_or_ini_r), .A0(cmnd_addr[9]), .A1(rst_addr_r[9]), .Z(sw_add[9]));
Q_MX02 U114 ( .S(rst_or_ini_r), .A0(cmnd_addr[10]), .A1(rst_addr_r[10]), .Z(sw_add[10]));
Q_MX02 U115 ( .S(rst_or_ini_r), .A0(cmnd_addr[11]), .A1(rst_addr_r[11]), .Z(sw_add[11]));
Q_MX02 U116 ( .S(rst_or_ini_r), .A0(cmnd_addr[12]), .A1(rst_addr_r[12]), .Z(sw_add[12]));
Q_MX02 U117 ( .S(rst_or_ini_r), .A0(cmnd_addr[13]), .A1(rst_addr_r[13]), .Z(sw_add[13]));
Q_AN02 U118 ( .A0(enable), .A1(\addr_limit[0][0] ), .Z(maxaddr[0]));
Q_AN02 U119 ( .A0(enable), .A1(\addr_limit[0][1] ), .Z(maxaddr[1]));
Q_AN02 U120 ( .A0(enable), .A1(\addr_limit[0][2] ), .Z(maxaddr[2]));
Q_AN02 U121 ( .A0(enable), .A1(\addr_limit[0][3] ), .Z(maxaddr[3]));
Q_AN02 U122 ( .A0(enable), .A1(\addr_limit[0][4] ), .Z(maxaddr[4]));
Q_AN02 U123 ( .A0(enable), .A1(\addr_limit[0][5] ), .Z(maxaddr[5]));
Q_AN02 U124 ( .A0(enable), .A1(\addr_limit[0][6] ), .Z(maxaddr[6]));
Q_AN02 U125 ( .A0(enable), .A1(\addr_limit[0][7] ), .Z(maxaddr[7]));
Q_AN02 U126 ( .A0(enable), .A1(\addr_limit[0][8] ), .Z(maxaddr[8]));
Q_AN02 U127 ( .A0(enable), .A1(\addr_limit[0][9] ), .Z(maxaddr[9]));
Q_AN02 U128 ( .A0(enable), .A1(\addr_limit[0][10] ), .Z(maxaddr[10]));
Q_AN02 U129 ( .A0(enable), .A1(\addr_limit[0][11] ), .Z(maxaddr[11]));
Q_AN02 U130 ( .A0(enable), .A1(\addr_limit[0][12] ), .Z(maxaddr[12]));
Q_AN02 U131 ( .A0(enable), .A1(\addr_limit[0][13] ), .Z(maxaddr[13]));
Q_INV U132 ( .A(reg_addr[3]), .Z(n55));
Q_INV U133 ( .A(reg_addr[4]), .Z(n56));
Q_INV U134 ( .A(reg_addr[5]), .Z(n57));
Q_INV U135 ( .A(reg_addr[7]), .Z(n58));
Q_INV U136 ( .A(reg_addr[8]), .Z(n59));
Q_OR03 U137 ( .A0(reg_addr[10]), .A1(reg_addr[9]), .A2(n59), .Z(n60));
Q_OR03 U138 ( .A0(n58), .A1(reg_addr[6]), .A2(n57), .Z(n61));
Q_OR03 U139 ( .A0(n56), .A1(n55), .A2(reg_addr[2]), .Z(n62));
Q_OR03 U140 ( .A0(reg_addr[1]), .A1(reg_addr[0]), .A2(n60), .Z(n63));
Q_NR03 U141 ( .A0(n61), .A1(n62), .A2(n63), .Z(n64));
Q_AN02 U142 ( .A0(wr_stb), .A1(n64), .Z(n87));
Q_INV U143 ( .A(n83), .Z(cmnd_issued));
Q_INV U144 ( .A(unsupported_op), .Z(n82));
Q_OA21 U145 ( .A0(n66), .A1(n67), .B0(n65), .Z(unsupported_op));
Q_AN02 U146 ( .A0(n65), .A1(n68), .Z(ack_error));
Q_AO21 U147 ( .A0(n70), .A1(n71), .B0(n69), .Z(n83));
Q_INV U148 ( .A(n87), .Z(n69));
Q_MX02 U149 ( .S(cmnd[3]), .A0(n74), .A1(n72), .Z(n70));
Q_INV U150 ( .A(cmnd_cmp_stb), .Z(n84));
Q_AN02 U151 ( .A0(n65), .A1(n75), .Z(cmnd_cmp_stb));
Q_AN02 U152 ( .A0(n65), .A1(n76), .Z(cmnd_tmo_stb));
Q_AN03 U153 ( .A0(n65), .A1(n71), .A2(n74), .Z(cmnd_sis_stb));
Q_AN02 U154 ( .A0(n87), .A1(cmnd[3]), .Z(n65));
Q_AN02 U155 ( .A0(n77), .A1(n68), .Z(cmnd_inc_stb));
Q_AN02 U156 ( .A0(n72), .A1(cmnd[0]), .Z(n68));
Q_AN02 U157 ( .A0(n77), .A1(n76), .Z(cmnd_ini_stb));
Q_AN02 U158 ( .A0(n72), .A1(n71), .Z(n76));
Q_AN02 U159 ( .A0(cmnd[2]), .A1(cmnd[1]), .Z(n72));
Q_INV U160 ( .A(cmnd_rst_stb), .Z(n85));
Q_AN02 U161 ( .A0(n67), .A1(n78), .Z(cmnd_rst_stb));
Q_AN02 U162 ( .A0(n77), .A1(cmnd[0]), .Z(n78));
Q_AN02 U163 ( .A0(n67), .A1(n79), .Z(cmnd_dis_stb));
Q_AN02 U164 ( .A0(n77), .A1(n71), .Z(n79));
Q_AN02 U165 ( .A0(cmnd[2]), .A1(n80), .Z(n67));
Q_AN02 U166 ( .A0(n66), .A1(n78), .Z(cmnd_ena_stb));
Q_INV U167 ( .A(cmnd_wr_stb), .Z(n86));
Q_AN02 U168 ( .A0(n66), .A1(n79), .Z(cmnd_wr_stb));
Q_INV U169 ( .A(cmnd[0]), .Z(n71));
Q_AN02 U170 ( .A0(n81), .A1(cmnd[1]), .Z(n66));
Q_AN02 U171 ( .A0(n77), .A1(n75), .Z(cmnd_rd_stb));
Q_AN02 U172 ( .A0(n74), .A1(cmnd[0]), .Z(n75));
Q_NR02 U173 ( .A0(cmnd[2]), .A1(cmnd[1]), .Z(n74));
Q_INV U174 ( .A(cmnd[1]), .Z(n80));
Q_INV U175 ( .A(cmnd[2]), .Z(n81));
Q_AN02 U176 ( .A0(n87), .A1(n73), .Z(n77));
Q_INV U177 ( .A(cmnd[3]), .Z(n73));
Q_OR02 U178 ( .A0(cmnd_ini_stb), .A1(cmnd_inc_stb), .Z(n436));
Q_XNR2 U179 ( .A0(rst_addr_r[0]), .A1(maxaddr[0]), .Z(n88));
Q_XNR2 U180 ( .A0(rst_addr_r[1]), .A1(maxaddr[1]), .Z(n89));
Q_XNR2 U181 ( .A0(rst_addr_r[2]), .A1(maxaddr[2]), .Z(n90));
Q_XNR2 U182 ( .A0(rst_addr_r[3]), .A1(maxaddr[3]), .Z(n91));
Q_XNR2 U183 ( .A0(rst_addr_r[4]), .A1(maxaddr[4]), .Z(n92));
Q_XNR2 U184 ( .A0(rst_addr_r[5]), .A1(maxaddr[5]), .Z(n93));
Q_XNR2 U185 ( .A0(rst_addr_r[6]), .A1(maxaddr[6]), .Z(n94));
Q_XNR2 U186 ( .A0(rst_addr_r[7]), .A1(maxaddr[7]), .Z(n95));
Q_XNR2 U187 ( .A0(rst_addr_r[8]), .A1(maxaddr[8]), .Z(n96));
Q_XNR2 U188 ( .A0(rst_addr_r[9]), .A1(maxaddr[9]), .Z(n97));
Q_XNR2 U189 ( .A0(rst_addr_r[10]), .A1(maxaddr[10]), .Z(n98));
Q_XNR2 U190 ( .A0(rst_addr_r[11]), .A1(maxaddr[11]), .Z(n99));
Q_XNR2 U191 ( .A0(rst_addr_r[12]), .A1(maxaddr[12]), .Z(n100));
Q_XNR2 U192 ( .A0(rst_addr_r[13]), .A1(maxaddr[13]), .Z(n101));
Q_AN03 U193 ( .A0(n101), .A1(n100), .A2(n99), .Z(n102));
Q_AN03 U194 ( .A0(n98), .A1(n97), .A2(n96), .Z(n103));
Q_AN03 U195 ( .A0(n95), .A1(n94), .A2(n93), .Z(n104));
Q_AN03 U196 ( .A0(n92), .A1(n91), .A2(n90), .Z(n105));
Q_AN03 U197 ( .A0(n89), .A1(n88), .A2(n102), .Z(n106));
Q_AN03 U198 ( .A0(n103), .A1(n104), .A2(n105), .Z(n107));
Q_AN02 U199 ( .A0(n106), .A1(n107), .Z(n437));
Q_XNR2 U200 ( .A0(rst_addr_r[0]), .A1(cmnd_addr[0]), .Z(n108));
Q_XNR2 U201 ( .A0(rst_addr_r[1]), .A1(cmnd_addr[1]), .Z(n109));
Q_XNR2 U202 ( .A0(rst_addr_r[2]), .A1(cmnd_addr[2]), .Z(n110));
Q_XNR2 U203 ( .A0(rst_addr_r[3]), .A1(cmnd_addr[3]), .Z(n111));
Q_XNR2 U204 ( .A0(rst_addr_r[4]), .A1(cmnd_addr[4]), .Z(n112));
Q_XNR2 U205 ( .A0(rst_addr_r[5]), .A1(cmnd_addr[5]), .Z(n113));
Q_XNR2 U206 ( .A0(rst_addr_r[6]), .A1(cmnd_addr[6]), .Z(n114));
Q_XNR2 U207 ( .A0(rst_addr_r[7]), .A1(cmnd_addr[7]), .Z(n115));
Q_XNR2 U208 ( .A0(rst_addr_r[8]), .A1(cmnd_addr[8]), .Z(n116));
Q_XNR2 U209 ( .A0(rst_addr_r[9]), .A1(cmnd_addr[9]), .Z(n117));
Q_XNR2 U210 ( .A0(rst_addr_r[10]), .A1(cmnd_addr[10]), .Z(n118));
Q_XNR2 U211 ( .A0(rst_addr_r[11]), .A1(cmnd_addr[11]), .Z(n119));
Q_XNR2 U212 ( .A0(rst_addr_r[12]), .A1(cmnd_addr[12]), .Z(n120));
Q_XNR2 U213 ( .A0(rst_addr_r[13]), .A1(cmnd_addr[13]), .Z(n121));
Q_AN03 U214 ( .A0(n121), .A1(n120), .A2(n119), .Z(n122));
Q_AN03 U215 ( .A0(n118), .A1(n117), .A2(n116), .Z(n123));
Q_AN03 U216 ( .A0(n115), .A1(n114), .A2(n113), .Z(n124));
Q_AN03 U217 ( .A0(n112), .A1(n111), .A2(n110), .Z(n125));
Q_AN03 U218 ( .A0(n109), .A1(n108), .A2(n122), .Z(n126));
Q_AN03 U219 ( .A0(n123), .A1(n124), .A2(n125), .Z(n127));
Q_AN02 U220 ( .A0(n126), .A1(n127), .Z(n438));
Q_AN02 U221 ( .A0(init_inc_r), .A1(igrant), .Z(n128));
Q_XOR2 U222 ( .A0(inc_r[0]), .A1(n128), .Z(n129));
Q_AD01HF U223 ( .A0(rst_addr_r[0]), .B0(igrant), .S(n130), .CO(n131));
Q_AD01HF U224 ( .A0(rst_addr_r[1]), .B0(n131), .S(n132), .CO(n133));
Q_AD01HF U225 ( .A0(rst_addr_r[2]), .B0(n133), .S(n134), .CO(n135));
Q_AD01HF U226 ( .A0(rst_addr_r[3]), .B0(n135), .S(n136), .CO(n137));
Q_AD01HF U227 ( .A0(rst_addr_r[4]), .B0(n137), .S(n138), .CO(n139));
Q_AD01HF U228 ( .A0(rst_addr_r[5]), .B0(n139), .S(n140), .CO(n141));
Q_AD01HF U229 ( .A0(rst_addr_r[6]), .B0(n141), .S(n142), .CO(n143));
Q_AD01HF U230 ( .A0(rst_addr_r[7]), .B0(n143), .S(n144), .CO(n145));
Q_AD01HF U231 ( .A0(rst_addr_r[8]), .B0(n145), .S(n146), .CO(n147));
Q_AD01HF U232 ( .A0(rst_addr_r[9]), .B0(n147), .S(n148), .CO(n149));
Q_AD01HF U233 ( .A0(rst_addr_r[10]), .B0(n149), .S(n150), .CO(n151));
Q_AD01HF U234 ( .A0(rst_addr_r[11]), .B0(n151), .S(n152), .CO(n153));
Q_AD01HF U235 ( .A0(rst_addr_r[12]), .B0(n153), .S(n154), .CO(n155));
Q_XOR2 U236 ( .A0(rst_addr_r[13]), .A1(n155), .Z(n156));
Q_AD01HF U237 ( .A0(timer_r[1]), .B0(timer_r[0]), .S(n158), .CO(n159));
Q_AD01HF U238 ( .A0(timer_r[2]), .B0(n159), .S(n160), .CO(n161));
Q_AD01HF U239 ( .A0(timer_r[3]), .B0(n161), .S(n162), .CO(n163));
Q_AD01HF U240 ( .A0(timer_r[4]), .B0(n163), .S(n164), .CO(n165));
Q_XOR2 U241 ( .A0(timer_r[5]), .A1(n165), .Z(n166));
Q_INV U242 ( .A(n167), .Z(n168));
Q_MX02 U243 ( .S(n359), .A0(n171), .A1(n169), .Z(n167));
Q_XOR2 U244 ( .A0(n414), .A1(n170), .Z(n169));
Q_AN02 U245 ( .A0(n413), .A1(n415), .Z(n170));
Q_OR02 U246 ( .A0(n414), .A1(n172), .Z(n171));
Q_INV U247 ( .A(n173), .Z(n174));
Q_MX02 U248 ( .S(n414), .A0(n175), .A1(n176), .Z(n173));
Q_ND02 U249 ( .A0(n292), .A1(n415), .Z(n176));
Q_AN02 U250 ( .A0(n359), .A1(n178), .Z(n177));
Q_MX02 U251 ( .S(n414), .A0(n179), .A1(n172), .Z(n178));
Q_NR02 U252 ( .A0(n292), .A1(n415), .Z(n179));
Q_OR02 U253 ( .A0(n413), .A1(n415), .Z(n172));
Q_NR03 U254 ( .A0(n416), .A1(n414), .A2(n181), .Z(n180));
Q_INV U255 ( .A(n175), .Z(n181));
Q_XOR2 U256 ( .A0(n292), .A1(n415), .Z(n175));
Q_AN02 U257 ( .A0(n416), .A1(n414), .Z(n182));
Q_AO21 U258 ( .A0(n182), .A1(state_r[3]), .B0(n180), .Z(n442));
Q_AO21 U259 ( .A0(n182), .A1(state_r[2]), .B0(n177), .Z(n441));
Q_AO21 U260 ( .A0(n182), .A1(state_r[1]), .B0(n174), .Z(n440));
Q_AO21 U261 ( .A0(n182), .A1(state_r[0]), .B0(n168), .Z(n439));
Q_AN02 U262 ( .A0(n417), .A1(n157), .Z(n183));
Q_AN02 U263 ( .A0(n417), .A1(n158), .Z(n184));
Q_AN02 U264 ( .A0(n417), .A1(n160), .Z(n185));
Q_AN02 U265 ( .A0(n417), .A1(n162), .Z(n186));
Q_AN02 U266 ( .A0(n417), .A1(n164), .Z(n187));
Q_AN02 U267 ( .A0(n417), .A1(n166), .Z(n188));
Q_AN02 U268 ( .A0(n419), .A1(cmnd_addr[0]), .Z(n189));
Q_MX02 U269 ( .S(n420), .A0(n189), .A1(n130), .Z(n190));
Q_AN02 U270 ( .A0(n419), .A1(cmnd_addr[1]), .Z(n191));
Q_MX02 U271 ( .S(n420), .A0(n191), .A1(n132), .Z(n192));
Q_AN02 U272 ( .A0(n419), .A1(cmnd_addr[2]), .Z(n193));
Q_MX02 U273 ( .S(n420), .A0(n193), .A1(n134), .Z(n194));
Q_AN02 U274 ( .A0(n419), .A1(cmnd_addr[3]), .Z(n195));
Q_MX02 U275 ( .S(n420), .A0(n195), .A1(n136), .Z(n196));
Q_AN02 U276 ( .A0(n419), .A1(cmnd_addr[4]), .Z(n197));
Q_MX02 U277 ( .S(n420), .A0(n197), .A1(n138), .Z(n198));
Q_AN02 U278 ( .A0(n419), .A1(cmnd_addr[5]), .Z(n199));
Q_MX02 U279 ( .S(n420), .A0(n199), .A1(n140), .Z(n200));
Q_AN02 U280 ( .A0(n419), .A1(cmnd_addr[6]), .Z(n201));
Q_MX02 U281 ( .S(n420), .A0(n201), .A1(n142), .Z(n202));
Q_AN02 U282 ( .A0(n419), .A1(cmnd_addr[7]), .Z(n203));
Q_MX02 U283 ( .S(n420), .A0(n203), .A1(n144), .Z(n204));
Q_AN02 U284 ( .A0(n419), .A1(cmnd_addr[8]), .Z(n205));
Q_MX02 U285 ( .S(n420), .A0(n205), .A1(n146), .Z(n206));
Q_AN02 U286 ( .A0(n419), .A1(cmnd_addr[9]), .Z(n207));
Q_MX02 U287 ( .S(n420), .A0(n207), .A1(n148), .Z(n208));
Q_AN02 U288 ( .A0(n419), .A1(cmnd_addr[10]), .Z(n209));
Q_MX02 U289 ( .S(n420), .A0(n209), .A1(n150), .Z(n210));
Q_AN02 U290 ( .A0(n419), .A1(cmnd_addr[11]), .Z(n211));
Q_MX02 U291 ( .S(n420), .A0(n211), .A1(n152), .Z(n212));
Q_AN02 U292 ( .A0(n419), .A1(cmnd_addr[12]), .Z(n213));
Q_MX02 U293 ( .S(n420), .A0(n213), .A1(n154), .Z(n214));
Q_AN02 U294 ( .A0(n419), .A1(cmnd_addr[13]), .Z(n215));
Q_MX02 U295 ( .S(n420), .A0(n215), .A1(n156), .Z(n216));
Q_AN02 U296 ( .A0(n425), .A1(n129), .Z(n217));
Q_MX03 U297 ( .S0(n427), .S1(n428), .A0(sw_aindex[0]), .A1(wr_dat[0]), .A2(sw_rdat[0]), .Z(n218));
Q_MX03 U298 ( .S0(n427), .S1(n428), .A0(sw_aindex[1]), .A1(wr_dat[1]), .A2(sw_rdat[1]), .Z(n219));
Q_MX03 U299 ( .S0(n427), .S1(n428), .A0(sw_aindex[2]), .A1(wr_dat[2]), .A2(sw_rdat[2]), .Z(n220));
Q_MX03 U300 ( .S0(n427), .S1(n428), .A0(sw_aindex[3]), .A1(wr_dat[3]), .A2(sw_rdat[3]), .Z(n221));
Q_MX03 U301 ( .S0(n427), .S1(n428), .A0(sw_aindex[4]), .A1(wr_dat[4]), .A2(sw_rdat[4]), .Z(n222));
Q_MX03 U302 ( .S0(n427), .S1(n428), .A0(sw_aindex[5]), .A1(wr_dat[5]), .A2(sw_rdat[5]), .Z(n223));
Q_MX03 U303 ( .S0(n427), .S1(n428), .A0(sw_aindex[6]), .A1(wr_dat[6]), .A2(sw_rdat[6]), .Z(n224));
Q_MX03 U304 ( .S0(n427), .S1(n428), .A0(sw_aindex[7]), .A1(wr_dat[7]), .A2(sw_rdat[7]), .Z(n225));
Q_MX03 U305 ( .S0(n427), .S1(n428), .A0(sw_aindex[8]), .A1(wr_dat[8]), .A2(sw_rdat[8]), .Z(n226));
Q_MX03 U306 ( .S0(n427), .S1(n428), .A0(sw_aindex[9]), .A1(wr_dat[9]), .A2(sw_rdat[9]), .Z(n227));
Q_MX03 U307 ( .S0(n427), .S1(n428), .A0(sw_aindex[10]), .A1(wr_dat[10]), .A2(sw_rdat[10]), .Z(n228));
Q_MX03 U308 ( .S0(n427), .S1(n428), .A0(sw_aindex[11]), .A1(wr_dat[11]), .A2(sw_rdat[11]), .Z(n229));
Q_MX03 U309 ( .S0(n427), .S1(n428), .A0(sw_aindex[12]), .A1(wr_dat[12]), .A2(sw_rdat[12]), .Z(n230));
Q_MX03 U310 ( .S0(n427), .S1(n428), .A0(sw_match), .A1(wr_dat[13]), .A2(sw_rdat[13]), .Z(n231));
Q_AN02 U311 ( .A0(n427), .A1(wr_dat[14]), .Z(n232));
Q_MX02 U312 ( .S(n428), .A0(n232), .A1(sw_rdat[14]), .Z(n233));
Q_AN02 U313 ( .A0(n427), .A1(wr_dat[15]), .Z(n234));
Q_MX02 U314 ( .S(n428), .A0(n234), .A1(sw_rdat[15]), .Z(n235));
Q_AN02 U315 ( .A0(n427), .A1(wr_dat[16]), .Z(n236));
Q_MX02 U316 ( .S(n428), .A0(n236), .A1(sw_rdat[16]), .Z(n237));
Q_AN02 U317 ( .A0(n427), .A1(wr_dat[17]), .Z(n238));
Q_MX02 U318 ( .S(n428), .A0(n238), .A1(sw_rdat[17]), .Z(n239));
Q_AN02 U319 ( .A0(n427), .A1(wr_dat[18]), .Z(n240));
Q_MX02 U320 ( .S(n428), .A0(n240), .A1(sw_rdat[18]), .Z(n241));
Q_AN02 U321 ( .A0(n427), .A1(wr_dat[19]), .Z(n242));
Q_MX02 U322 ( .S(n428), .A0(n242), .A1(sw_rdat[19]), .Z(n243));
Q_AN02 U323 ( .A0(n427), .A1(wr_dat[20]), .Z(n244));
Q_MX02 U324 ( .S(n428), .A0(n244), .A1(sw_rdat[20]), .Z(n245));
Q_AN02 U325 ( .A0(n427), .A1(wr_dat[21]), .Z(n246));
Q_MX02 U326 ( .S(n428), .A0(n246), .A1(sw_rdat[21]), .Z(n247));
Q_AN02 U327 ( .A0(n427), .A1(wr_dat[22]), .Z(n248));
Q_MX02 U328 ( .S(n428), .A0(n248), .A1(sw_rdat[22]), .Z(n249));
Q_AN02 U329 ( .A0(n427), .A1(wr_dat[23]), .Z(n250));
Q_MX02 U330 ( .S(n428), .A0(n250), .A1(sw_rdat[23]), .Z(n251));
Q_AN02 U331 ( .A0(n427), .A1(wr_dat[24]), .Z(n252));
Q_MX02 U332 ( .S(n428), .A0(n252), .A1(sw_rdat[24]), .Z(n253));
Q_AN02 U333 ( .A0(n427), .A1(wr_dat[25]), .Z(n254));
Q_MX02 U334 ( .S(n428), .A0(n254), .A1(sw_rdat[25]), .Z(n255));
Q_AN02 U335 ( .A0(n427), .A1(wr_dat[26]), .Z(n256));
Q_MX02 U336 ( .S(n428), .A0(n256), .A1(sw_rdat[26]), .Z(n257));
Q_AN02 U337 ( .A0(n427), .A1(wr_dat[27]), .Z(n258));
Q_MX02 U338 ( .S(n428), .A0(n258), .A1(sw_rdat[27]), .Z(n259));
Q_AN02 U339 ( .A0(n427), .A1(wr_dat[28]), .Z(n260));
Q_MX02 U340 ( .S(n428), .A0(n260), .A1(sw_rdat[28]), .Z(n261));
Q_AN02 U341 ( .A0(n427), .A1(wr_dat[29]), .Z(n262));
Q_MX02 U342 ( .S(n428), .A0(n262), .A1(sw_rdat[29]), .Z(n263));
Q_AN02 U343 ( .A0(n427), .A1(wr_dat[30]), .Z(n264));
Q_MX02 U344 ( .S(n428), .A0(n264), .A1(sw_rdat[30]), .Z(n265));
Q_AN02 U345 ( .A0(n427), .A1(wr_dat[31]), .Z(n266));
Q_MX02 U346 ( .S(n428), .A0(n266), .A1(sw_rdat[31]), .Z(n267));
Q_AN02 U347 ( .A0(n427), .A1(wr_dat[32]), .Z(n268));
Q_MX02 U348 ( .S(n428), .A0(n268), .A1(sw_rdat[32]), .Z(n269));
Q_AN02 U349 ( .A0(n427), .A1(wr_dat[33]), .Z(n270));
Q_MX02 U350 ( .S(n428), .A0(n270), .A1(sw_rdat[33]), .Z(n271));
Q_AN02 U351 ( .A0(n427), .A1(wr_dat[34]), .Z(n272));
Q_MX02 U352 ( .S(n428), .A0(n272), .A1(sw_rdat[34]), .Z(n273));
Q_AN02 U353 ( .A0(n427), .A1(wr_dat[35]), .Z(n274));
Q_MX02 U354 ( .S(n428), .A0(n274), .A1(sw_rdat[35]), .Z(n275));
Q_AN02 U355 ( .A0(n427), .A1(wr_dat[36]), .Z(n276));
Q_MX02 U356 ( .S(n428), .A0(n276), .A1(sw_rdat[36]), .Z(n277));
Q_AN02 U357 ( .A0(n427), .A1(wr_dat[37]), .Z(n278));
Q_MX02 U358 ( .S(n428), .A0(n278), .A1(sw_rdat[37]), .Z(n279));
Q_FDP1 \state_r_REG[3] ( .CK(clk), .R(rst_n), .D(n442), .Q(state_r[3]), .QN(n307));
Q_FDP1 \state_r_REG[2] ( .CK(clk), .R(rst_n), .D(n441), .Q(state_r[2]), .QN(n308));
Q_FDP1 \state_r_REG[1] ( .CK(clk), .R(rst_n), .D(n440), .Q(state_r[1]), .QN(n310));
Q_FDP1 \state_r_REG[0] ( .CK(clk), .R(rst_n), .D(n439), .Q(state_r[0]), .QN(n306));
Q_FDP1 \timer_r_REG[5] ( .CK(clk), .R(rst_n), .D(n188), .Q(timer_r[5]), .QN( ));
Q_FDP1 \timer_r_REG[4] ( .CK(clk), .R(rst_n), .D(n187), .Q(timer_r[4]), .QN( ));
Q_FDP1 \timer_r_REG[3] ( .CK(clk), .R(rst_n), .D(n186), .Q(timer_r[3]), .QN( ));
Q_FDP1 \timer_r_REG[2] ( .CK(clk), .R(rst_n), .D(n185), .Q(timer_r[2]), .QN( ));
Q_FDP1 \timer_r_REG[1] ( .CK(clk), .R(rst_n), .D(n184), .Q(timer_r[1]), .QN( ));
Q_FDP1 \timer_r_REG[0] ( .CK(clk), .R(rst_n), .D(n183), .Q(timer_r[0]), .QN(n157));
Q_ND02 U369 ( .A0(n281), .A1(n282), .Z(n280));
Q_ND02 U370 ( .A0(n283), .A1(n385), .Z(n282));
Q_OR02 U371 ( .A0(n284), .A1(n430), .Z(n283));
Q_INV U372 ( .A(n429), .Z(n284));
Q_ND02 U373 ( .A0(n281), .A1(n286), .Z(n285));
Q_ND02 U374 ( .A0(n429), .A1(n385), .Z(n286));
Q_OR03 U375 ( .A0(n429), .A1(n430), .A2(n385), .Z(n281));
Q_MX02 U376 ( .S(n385), .A0(n429), .A1(n430), .Z(n287));
Q_FDP2 \stat_code_REG[2] ( .CK(clk), .S(rst_n), .D(n288), .Q(stat_code[2]), .QN( ));
Q_MX02 U378 ( .S(n400), .A0(stat_code[2]), .A1(n287), .Z(n288));
Q_FDP2 \stat_code_REG[1] ( .CK(clk), .S(rst_n), .D(n289), .Q(stat_code[1]), .QN( ));
Q_MX02 U380 ( .S(n400), .A0(stat_code[1]), .A1(n285), .Z(n289));
Q_FDP2 \stat_code_REG[0] ( .CK(clk), .S(rst_n), .D(n290), .Q(stat_code[0]), .QN( ));
Q_MX02 U382 ( .S(n400), .A0(stat_code[0]), .A1(n280), .Z(n290));
Q_FDP2 init_r_REG  ( .CK(clk), .S(rst_n), .D(n291), .Q(init_r), .QN(enable));
Q_MX02 U384 ( .S(n432), .A0(init_r), .A1(n426), .Z(n291));
Q_FDP1 sw_cs_r_REG  ( .CK(clk), .R(rst_n), .D(n424), .Q(sw_cs_r), .QN( ));
Q_FDP1 sw_ce_r_REG  ( .CK(clk), .R(rst_n), .D(n423), .Q(sw_ce_r), .QN( ));
Q_FDP1 rst_r_REG  ( .CK(clk), .R(rst_n), .D(n422), .Q(rst_r), .QN(n443));
Q_FDP1 rst_or_ini_r_REG  ( .CK(clk), .R(rst_n), .D(n421), .Q(rst_or_ini_r), .QN( ));
Q_FDP1 sw_we_r_REG  ( .CK(clk), .R(rst_n), .D(n418), .Q(sw_we_r), .QN( ));
Q_INV U390 ( .A(n292), .Z(n413));
Q_OA21 U391 ( .A0(n294), .A1(n295), .B0(n293), .Z(n292));
Q_AN03 U392 ( .A0(state_r[0]), .A1(n299), .A2(n297), .Z(n298));
Q_OR03 U393 ( .A0(n301), .A1(n302), .A2(n296), .Z(n295));
Q_AO21 U394 ( .A0(n303), .A1(n304), .B0(n298), .Z(n300));
Q_AN02 U395 ( .A0(n305), .A1(n306), .Z(n304));
Q_NR02 U396 ( .A0(state_r[3]), .A1(state_r[2]), .Z(n305));
Q_MX02 U397 ( .S(state_r[1]), .A0(cmnd_ena_stb), .A1(n309), .Z(n303));
Q_AN02 U398 ( .A0(n312), .A1(n83), .Z(n311));
Q_AO21 U399 ( .A0(n313), .A1(n314), .B0(n300), .Z(n301));
Q_NR02 U400 ( .A0(cmnd_dis_stb), .A1(unsupported_op), .Z(n314));
Q_OA21 U401 ( .A0(n315), .A1(n316), .B0(n311), .Z(n302));
Q_AN03 U402 ( .A0(n318), .A1(state_r[3]), .A2(n309), .Z(n317));
Q_AN02 U403 ( .A0(ack_error), .A1(enable), .Z(n309));
Q_OR02 U404 ( .A0(n319), .A1(n317), .Z(n316));
Q_AN02 U405 ( .A0(n307), .A1(igrant), .Z(n320));
Q_OA21 U406 ( .A0(n321), .A1(n322), .B0(n320), .Z(n315));
Q_AN02 U407 ( .A0(n324), .A1(n437), .Z(n321));
Q_OA21 U408 ( .A0(state_r[0]), .A1(n438), .B0(n323), .Z(n322));
Q_AN02 U409 ( .A0(n328), .A1(n84), .Z(n326));
Q_AN03 U410 ( .A0(cmnd_rst_stb), .A1(n297), .A2(n326), .Z(n327));
Q_OR03 U411 ( .A0(n329), .A1(n327), .A2(n325), .Z(n294));
Q_AN02 U412 ( .A0(n330), .A1(n331), .Z(n329));
Q_NR02 U413 ( .A0(timeout), .A1(state_r[0]), .Z(n332));
Q_OA21 U414 ( .A0(n333), .A1(n296), .B0(n293), .Z(n414));
Q_OR02 U415 ( .A0(n334), .A1(n335), .Z(n333));
Q_AO21 U416 ( .A0(n338), .A1(n339), .B0(n336), .Z(n296));
Q_AN02 U417 ( .A0(n340), .A1(n83), .Z(n339));
Q_NR02 U418 ( .A0(timeout), .A1(state_r[3]), .Z(n340));
Q_OA21 U419 ( .A0(n341), .A1(n342), .B0(n337), .Z(n336));
Q_AN02 U420 ( .A0(n307), .A1(n343), .Z(n342));
Q_NR02 U421 ( .A0(state_r[0]), .A1(cmnd_ena_stb), .Z(n343));
Q_AN02 U422 ( .A0(n344), .A1(n345), .Z(n341));
Q_MX02 U423 ( .S(state_r[0]), .A0(n347), .A1(n346), .Z(n344));
Q_AO21 U424 ( .A0(n349), .A1(n324), .B0(n348), .Z(n338));
Q_OA21 U425 ( .A0(n350), .A1(n351), .B0(state_r[2]), .Z(n348));
Q_NR02 U426 ( .A0(n352), .A1(rsp), .Z(n351));
Q_INV U427 ( .A(rsp), .Z(n346));
Q_AO21 U428 ( .A0(n352), .A1(n347), .B0(n353), .Z(n350));
Q_NR02 U429 ( .A0(n354), .A1(n438), .Z(n353));
Q_ND02 U430 ( .A0(igrant), .A1(n437), .Z(n349));
Q_OA21 U431 ( .A0(n355), .A1(n356), .B0(n434), .Z(n415));
Q_AN02 U432 ( .A0(n357), .A1(n358), .Z(n355));
Q_INV U433 ( .A(n359), .Z(n416));
Q_OA21 U434 ( .A0(n360), .A1(n334), .B0(n293), .Z(n359));
Q_AN03 U435 ( .A0(n356), .A1(state_r[0]), .A2(n297), .Z(n335));
Q_INV U436 ( .A(n358), .Z(n356));
Q_AN02 U437 ( .A0(n86), .A1(cmnd_rd_stb), .Z(n299));
Q_AN03 U438 ( .A0(n297), .A1(n328), .A2(n357), .Z(n361));
Q_AO21 U439 ( .A0(cmnd_rst_stb), .A1(n84), .B0(cmnd_cmp_stb), .Z(n357));
Q_OR03 U440 ( .A0(n362), .A1(n361), .A2(n335), .Z(n360));
Q_AN02 U441 ( .A0(n363), .A1(n330), .Z(n362));
Q_AN03 U442 ( .A0(igrant), .A1(n83), .A2(n332), .Z(n330));
Q_AO21 U443 ( .A0(n364), .A1(n365), .B0(n325), .Z(n334));
Q_AN03 U444 ( .A0(n84), .A1(n436), .A2(n328), .Z(n365));
Q_AN02 U445 ( .A0(ack_error), .A1(init_r), .Z(n367));
Q_AO21 U446 ( .A0(n313), .A1(cmnd_dis_stb), .B0(n366), .Z(n325));
Q_AN03 U447 ( .A0(n328), .A1(n368), .A2(n364), .Z(n313));
Q_NR02 U448 ( .A0(cmnd_cmp_stb), .A1(n436), .Z(n368));
Q_AN02 U449 ( .A0(state_r[0]), .A1(n358), .Z(n328));
Q_NR02 U450 ( .A0(cmnd_wr_stb), .A1(cmnd_rd_stb), .Z(n358));
Q_AN02 U451 ( .A0(n85), .A1(n297), .Z(n364));
Q_OA21 U452 ( .A0(n369), .A1(n370), .B0(n367), .Z(n366));
Q_AN02 U453 ( .A0(n318), .A1(n345), .Z(n369));
Q_AN03 U454 ( .A0(n312), .A1(state_r[3]), .A2(n83), .Z(n345));
Q_INV U455 ( .A(n337), .Z(n318));
Q_AN02 U456 ( .A0(n347), .A1(n424), .Z(n417));
Q_INV U457 ( .A(igrant), .Z(n347));
Q_OA21 U458 ( .A0(n372), .A1(n373), .B0(n371), .Z(n418));
Q_AN02 U459 ( .A0(cmnd_sis_stb), .A1(n374), .Z(n419));
Q_INV U460 ( .A(n420), .Z(n374));
Q_OR02 U461 ( .A0(state_r[0]), .A1(state_r[1]), .Z(n354));
Q_ND02 U462 ( .A0(state_r[1]), .A1(state_r[0]), .Z(n352));
Q_OA21 U463 ( .A0(n372), .A1(n375), .B0(n371), .Z(n421));
Q_AN02 U464 ( .A0(n373), .A1(n376), .Z(n375));
Q_AN02 U465 ( .A0(n441), .A1(n377), .Z(n373));
Q_AN02 U466 ( .A0(n371), .A1(n372), .Z(n422));
Q_AN02 U467 ( .A0(n378), .A1(n439), .Z(n372));
Q_OR03 U468 ( .A0(n422), .A1(n379), .A2(n423), .Z(n424));
Q_AN02 U469 ( .A0(n442), .A1(n380), .Z(n423));
Q_AN03 U470 ( .A0(n371), .A1(n441), .A2(n381), .Z(n379));
Q_INV U471 ( .A(n382), .Z(n381));
Q_INV U472 ( .A(n383), .Z(n425));
Q_AN02 U473 ( .A0(n384), .A1(state_r[0]), .Z(n428));
Q_AN02 U474 ( .A0(n387), .A1(n388), .Z(n389));
Q_INV U475 ( .A(n390), .Z(n387));
Q_OR03 U476 ( .A0(n391), .A1(n389), .A2(n386), .Z(n385));
Q_AN03 U477 ( .A0(n393), .A1(n82), .A2(n392), .Z(n386));
Q_OR02 U478 ( .A0(n382), .A1(n394), .Z(n391));
Q_AN02 U479 ( .A0(n440), .A1(n439), .Z(n382));
Q_INV U480 ( .A(n395), .Z(n394));
Q_AN02 U481 ( .A0(n371), .A1(n396), .Z(n388));
Q_NR02 U482 ( .A0(n441), .A1(n439), .Z(n396));
Q_OA21 U483 ( .A0(n398), .A1(n377), .B0(n388), .Z(n429));
Q_AN02 U484 ( .A0(n82), .A1(n440), .Z(n390));
Q_OA21 U485 ( .A0(n393), .A1(badaddr), .B0(n390), .Z(n398));
Q_AN02 U486 ( .A0(timeout), .A1(n293), .Z(n393));
Q_NR02 U487 ( .A0(n442), .A1(n441), .Z(n395));
Q_OA21 U488 ( .A0(n399), .A1(n377), .B0(n395), .Z(n430));
Q_AN03 U489 ( .A0(n440), .A1(n376), .A2(unsupported_op), .Z(n399));
Q_ND02 U490 ( .A0(n370), .A1(n392), .Z(n400));
Q_AN02 U491 ( .A0(n378), .A1(n401), .Z(n392));
Q_NR02 U492 ( .A0(n442), .A1(n439), .Z(n401));
Q_AN02 U493 ( .A0(n397), .A1(n440), .Z(n378));
Q_AN02 U494 ( .A0(n402), .A1(n403), .Z(n370));
Q_NR02 U495 ( .A0(state_r[3]), .A1(state_r[0]), .Z(n402));
Q_OA21 U496 ( .A0(n427), .A1(n319), .B0(n293), .Z(n431));
Q_AN03 U497 ( .A0(state_r[0]), .A1(rsp), .A2(n363), .Z(n319));
Q_INV U498 ( .A(n426), .Z(n427));
Q_AN02 U499 ( .A0(n307), .A1(n337), .Z(n297));
Q_OR02 U500 ( .A0(n384), .A1(n331), .Z(n363));
Q_AN02 U501 ( .A0(state_r[3]), .A1(n337), .Z(n331));
Q_AN03 U502 ( .A0(state_r[2]), .A1(state_r[1]), .A2(n307), .Z(n384));
Q_AN03 U503 ( .A0(n426), .A1(n371), .A2(n380), .Z(n404));
Q_AN02 U504 ( .A0(n405), .A1(n376), .Z(n380));
Q_INV U505 ( .A(n439), .Z(n376));
Q_NR02 U506 ( .A0(n441), .A1(n440), .Z(n405));
Q_INV U507 ( .A(n440), .Z(n377));
Q_INV U508 ( .A(n441), .Z(n397));
Q_INV U509 ( .A(n442), .Z(n371));
Q_AO21 U510 ( .A0(n406), .A1(n407), .B0(n404), .Z(n432));
Q_AN02 U511 ( .A0(n306), .A1(cmnd_ena_stb), .Z(n407));
Q_OR02 U512 ( .A0(state_r[3]), .A1(state_r[1]), .Z(n408));
Q_OR03 U513 ( .A0(state_r[2]), .A1(state_r[0]), .A2(n408), .Z(n426));
Q_AN03 U514 ( .A0(n410), .A1(n310), .A2(n409), .Z(n433));
Q_AO21 U515 ( .A0(state_r[2]), .A1(n306), .B0(n383), .Z(n409));
Q_AN02 U516 ( .A0(n308), .A1(state_r[0]), .Z(n383));
Q_AN02 U517 ( .A0(n406), .A1(state_r[0]), .Z(n434));
Q_AN02 U518 ( .A0(n410), .A1(n337), .Z(n406));
Q_NR02 U519 ( .A0(state_r[2]), .A1(state_r[1]), .Z(n337));
Q_NR02 U520 ( .A0(badaddr), .A1(state_r[3]), .Z(n410));
Q_INV U521 ( .A(badaddr), .Z(n293));
Q_OR03 U522 ( .A0(cmnd_rst_stb), .A1(cmnd_sis_stb), .A2(n420), .Z(n435));
Q_OA21 U523 ( .A0(n324), .A1(n411), .B0(n410), .Z(n420));
Q_AN02 U524 ( .A0(n323), .A1(n306), .Z(n411));
Q_AN02 U525 ( .A0(state_r[2]), .A1(n310), .Z(n323));
Q_AN02 U526 ( .A0(n403), .A1(state_r[0]), .Z(n324));
Q_AN02 U527 ( .A0(n308), .A1(state_r[1]), .Z(n403));
Q_OR02 U528 ( .A0(cmnd_tmo_stb), .A1(timeout), .Z(n412));
Q_INV U529 ( .A(timeout), .Z(n312));
Q_AN02 U530 ( .A0(n443), .A1(wr_dat[0]), .Z(sw_wdat[0]));
Q_AN02 U531 ( .A0(n443), .A1(wr_dat[1]), .Z(sw_wdat[1]));
Q_AN02 U532 ( .A0(n443), .A1(wr_dat[2]), .Z(sw_wdat[2]));
Q_AN02 U533 ( .A0(n443), .A1(wr_dat[3]), .Z(sw_wdat[3]));
Q_AN02 U534 ( .A0(n443), .A1(wr_dat[4]), .Z(sw_wdat[4]));
Q_AN02 U535 ( .A0(n443), .A1(wr_dat[5]), .Z(sw_wdat[5]));
Q_AN02 U536 ( .A0(n443), .A1(wr_dat[6]), .Z(sw_wdat[6]));
Q_AN02 U537 ( .A0(n443), .A1(wr_dat[7]), .Z(sw_wdat[7]));
Q_AN02 U538 ( .A0(n443), .A1(wr_dat[8]), .Z(sw_wdat[8]));
Q_AN02 U539 ( .A0(n443), .A1(wr_dat[9]), .Z(sw_wdat[9]));
Q_AN02 U540 ( .A0(n443), .A1(wr_dat[10]), .Z(sw_wdat[10]));
Q_AN02 U541 ( .A0(n443), .A1(wr_dat[11]), .Z(sw_wdat[11]));
Q_AN02 U542 ( .A0(n443), .A1(wr_dat[12]), .Z(sw_wdat[12]));
Q_AN02 U543 ( .A0(n443), .A1(wr_dat[13]), .Z(sw_wdat[13]));
Q_AN02 U544 ( .A0(n443), .A1(wr_dat[14]), .Z(sw_wdat[14]));
Q_AN02 U545 ( .A0(n443), .A1(wr_dat[15]), .Z(sw_wdat[15]));
Q_AN02 U546 ( .A0(n443), .A1(wr_dat[16]), .Z(sw_wdat[16]));
Q_AN02 U547 ( .A0(n443), .A1(wr_dat[17]), .Z(sw_wdat[17]));
Q_AN02 U548 ( .A0(n443), .A1(wr_dat[18]), .Z(sw_wdat[18]));
Q_AN02 U549 ( .A0(n443), .A1(wr_dat[19]), .Z(sw_wdat[19]));
Q_AN02 U550 ( .A0(n443), .A1(wr_dat[20]), .Z(sw_wdat[20]));
Q_AN02 U551 ( .A0(n443), .A1(wr_dat[21]), .Z(sw_wdat[21]));
Q_AN02 U552 ( .A0(n443), .A1(wr_dat[22]), .Z(sw_wdat[22]));
Q_AN02 U553 ( .A0(n443), .A1(wr_dat[23]), .Z(sw_wdat[23]));
Q_AN02 U554 ( .A0(n443), .A1(wr_dat[24]), .Z(sw_wdat[24]));
Q_AN02 U555 ( .A0(n443), .A1(wr_dat[25]), .Z(sw_wdat[25]));
Q_AN02 U556 ( .A0(n443), .A1(wr_dat[26]), .Z(sw_wdat[26]));
Q_AN02 U557 ( .A0(n443), .A1(wr_dat[27]), .Z(sw_wdat[27]));
Q_AN02 U558 ( .A0(n443), .A1(wr_dat[28]), .Z(sw_wdat[28]));
Q_AN02 U559 ( .A0(n443), .A1(wr_dat[29]), .Z(sw_wdat[29]));
Q_AN02 U560 ( .A0(n443), .A1(wr_dat[30]), .Z(sw_wdat[30]));
Q_AN02 U561 ( .A0(n443), .A1(wr_dat[31]), .Z(sw_wdat[31]));
Q_AN02 U562 ( .A0(n443), .A1(wr_dat[32]), .Z(sw_wdat[32]));
Q_AN02 U563 ( .A0(n443), .A1(wr_dat[33]), .Z(sw_wdat[33]));
Q_AN02 U564 ( .A0(n443), .A1(wr_dat[34]), .Z(sw_wdat[34]));
Q_AN02 U565 ( .A0(n443), .A1(wr_dat[35]), .Z(sw_wdat[35]));
Q_AN02 U566 ( .A0(n443), .A1(wr_dat[36]), .Z(sw_wdat[36]));
Q_AN02 U567 ( .A0(n443), .A1(wr_dat[37]), .Z(sw_wdat[37]));
Q_FDP4EP sim_tmo_r_REG  ( .CK(clk), .CE(n412), .R(n444), .D(cmnd_tmo_stb), .Q(sim_tmo_r));
Q_INV U569 ( .A(rst_n), .Z(n444));
Q_INV U570 ( .A(sim_tmo_r), .Z(n54));
Q_FDP4EP \rst_addr_r_REG[0] ( .CK(clk), .CE(n435), .R(n444), .D(n190), .Q(rst_addr_r[0]));
Q_FDP4EP \rst_addr_r_REG[1] ( .CK(clk), .CE(n435), .R(n444), .D(n192), .Q(rst_addr_r[1]));
Q_FDP4EP \rst_addr_r_REG[2] ( .CK(clk), .CE(n435), .R(n444), .D(n194), .Q(rst_addr_r[2]));
Q_FDP4EP \rst_addr_r_REG[3] ( .CK(clk), .CE(n435), .R(n444), .D(n196), .Q(rst_addr_r[3]));
Q_FDP4EP \rst_addr_r_REG[4] ( .CK(clk), .CE(n435), .R(n444), .D(n198), .Q(rst_addr_r[4]));
Q_FDP4EP \rst_addr_r_REG[5] ( .CK(clk), .CE(n435), .R(n444), .D(n200), .Q(rst_addr_r[5]));
Q_FDP4EP \rst_addr_r_REG[6] ( .CK(clk), .CE(n435), .R(n444), .D(n202), .Q(rst_addr_r[6]));
Q_FDP4EP \rst_addr_r_REG[7] ( .CK(clk), .CE(n435), .R(n444), .D(n204), .Q(rst_addr_r[7]));
Q_FDP4EP \rst_addr_r_REG[8] ( .CK(clk), .CE(n435), .R(n444), .D(n206), .Q(rst_addr_r[8]));
Q_FDP4EP \rst_addr_r_REG[9] ( .CK(clk), .CE(n435), .R(n444), .D(n208), .Q(rst_addr_r[9]));
Q_FDP4EP \rst_addr_r_REG[10] ( .CK(clk), .CE(n435), .R(n444), .D(n210), .Q(rst_addr_r[10]));
Q_FDP4EP \rst_addr_r_REG[11] ( .CK(clk), .CE(n435), .R(n444), .D(n212), .Q(rst_addr_r[11]));
Q_FDP4EP \rst_addr_r_REG[12] ( .CK(clk), .CE(n435), .R(n444), .D(n214), .Q(rst_addr_r[12]));
Q_FDP4EP \rst_addr_r_REG[13] ( .CK(clk), .CE(n435), .R(n444), .D(n216), .Q(rst_addr_r[13]));
Q_FDP4EP \inc_r_REG[0] ( .CK(clk), .CE(n433), .R(n444), .D(n217), .Q(inc_r[0]));
Q_FDP4EP \rd_dat_REG[0] ( .CK(clk), .CE(n431), .R(n444), .D(n218), .Q(rd_dat[0]));
Q_FDP4EP \rd_dat_REG[1] ( .CK(clk), .CE(n431), .R(n444), .D(n219), .Q(rd_dat[1]));
Q_FDP4EP \rd_dat_REG[2] ( .CK(clk), .CE(n431), .R(n444), .D(n220), .Q(rd_dat[2]));
Q_FDP4EP \rd_dat_REG[3] ( .CK(clk), .CE(n431), .R(n444), .D(n221), .Q(rd_dat[3]));
Q_FDP4EP \rd_dat_REG[4] ( .CK(clk), .CE(n431), .R(n444), .D(n222), .Q(rd_dat[4]));
Q_FDP4EP \rd_dat_REG[5] ( .CK(clk), .CE(n431), .R(n444), .D(n223), .Q(rd_dat[5]));
Q_FDP4EP \rd_dat_REG[6] ( .CK(clk), .CE(n431), .R(n444), .D(n224), .Q(rd_dat[6]));
Q_FDP4EP \rd_dat_REG[7] ( .CK(clk), .CE(n431), .R(n444), .D(n225), .Q(rd_dat[7]));
Q_FDP4EP \rd_dat_REG[8] ( .CK(clk), .CE(n431), .R(n444), .D(n226), .Q(rd_dat[8]));
Q_FDP4EP \rd_dat_REG[9] ( .CK(clk), .CE(n431), .R(n444), .D(n227), .Q(rd_dat[9]));
Q_FDP4EP \rd_dat_REG[10] ( .CK(clk), .CE(n431), .R(n444), .D(n228), .Q(rd_dat[10]));
Q_FDP4EP \rd_dat_REG[11] ( .CK(clk), .CE(n431), .R(n444), .D(n229), .Q(rd_dat[11]));
Q_FDP4EP \rd_dat_REG[12] ( .CK(clk), .CE(n431), .R(n444), .D(n230), .Q(rd_dat[12]));
Q_FDP4EP \rd_dat_REG[13] ( .CK(clk), .CE(n431), .R(n444), .D(n231), .Q(rd_dat[13]));
Q_FDP4EP \rd_dat_REG[14] ( .CK(clk), .CE(n431), .R(n444), .D(n233), .Q(rd_dat[14]));
Q_FDP4EP \rd_dat_REG[15] ( .CK(clk), .CE(n431), .R(n444), .D(n235), .Q(rd_dat[15]));
Q_FDP4EP \rd_dat_REG[16] ( .CK(clk), .CE(n431), .R(n444), .D(n237), .Q(rd_dat[16]));
Q_FDP4EP \rd_dat_REG[17] ( .CK(clk), .CE(n431), .R(n444), .D(n239), .Q(rd_dat[17]));
Q_FDP4EP \rd_dat_REG[18] ( .CK(clk), .CE(n431), .R(n444), .D(n241), .Q(rd_dat[18]));
Q_FDP4EP \rd_dat_REG[19] ( .CK(clk), .CE(n431), .R(n444), .D(n243), .Q(rd_dat[19]));
Q_FDP4EP \rd_dat_REG[20] ( .CK(clk), .CE(n431), .R(n444), .D(n245), .Q(rd_dat[20]));
Q_FDP4EP \rd_dat_REG[21] ( .CK(clk), .CE(n431), .R(n444), .D(n247), .Q(rd_dat[21]));
Q_FDP4EP \rd_dat_REG[22] ( .CK(clk), .CE(n431), .R(n444), .D(n249), .Q(rd_dat[22]));
Q_FDP4EP \rd_dat_REG[23] ( .CK(clk), .CE(n431), .R(n444), .D(n251), .Q(rd_dat[23]));
Q_FDP4EP \rd_dat_REG[24] ( .CK(clk), .CE(n431), .R(n444), .D(n253), .Q(rd_dat[24]));
Q_FDP4EP \rd_dat_REG[25] ( .CK(clk), .CE(n431), .R(n444), .D(n255), .Q(rd_dat[25]));
Q_FDP4EP \rd_dat_REG[26] ( .CK(clk), .CE(n431), .R(n444), .D(n257), .Q(rd_dat[26]));
Q_FDP4EP \rd_dat_REG[27] ( .CK(clk), .CE(n431), .R(n444), .D(n259), .Q(rd_dat[27]));
Q_FDP4EP \rd_dat_REG[28] ( .CK(clk), .CE(n431), .R(n444), .D(n261), .Q(rd_dat[28]));
Q_FDP4EP \rd_dat_REG[29] ( .CK(clk), .CE(n431), .R(n444), .D(n263), .Q(rd_dat[29]));
Q_FDP4EP \rd_dat_REG[30] ( .CK(clk), .CE(n431), .R(n444), .D(n265), .Q(rd_dat[30]));
Q_FDP4EP \rd_dat_REG[31] ( .CK(clk), .CE(n431), .R(n444), .D(n267), .Q(rd_dat[31]));
Q_FDP4EP \rd_dat_REG[32] ( .CK(clk), .CE(n431), .R(n444), .D(n269), .Q(rd_dat[32]));
Q_FDP4EP \rd_dat_REG[33] ( .CK(clk), .CE(n431), .R(n444), .D(n271), .Q(rd_dat[33]));
Q_FDP4EP \rd_dat_REG[34] ( .CK(clk), .CE(n431), .R(n444), .D(n273), .Q(rd_dat[34]));
Q_FDP4EP \rd_dat_REG[35] ( .CK(clk), .CE(n431), .R(n444), .D(n275), .Q(rd_dat[35]));
Q_FDP4EP \rd_dat_REG[36] ( .CK(clk), .CE(n431), .R(n444), .D(n277), .Q(rd_dat[36]));
Q_FDP4EP \rd_dat_REG[37] ( .CK(clk), .CE(n431), .R(n444), .D(n279), .Q(rd_dat[37]));
Q_FDP4EP init_inc_r_REG  ( .CK(clk), .CE(n434), .R(n444), .D(n1), .Q(init_inc_r));
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "addr_limit (2,0) 1 13 0 0 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "1"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_1 "-1 genblk2  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_0 "-1 genblk1  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "genblk2"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "genblk1"
endmodule
