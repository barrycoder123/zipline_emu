architecture module of gfifo_conns is
  component gfifo_conns_0
  end component ;


begin
  gc0 : gfifo_conns_0
     ;
end module;
