
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module cr_kme_kim_drng_reader ( kimreader_parser_ack, kimreader_ckvreader_valid, 
	.kimreader_ckvreader_data( {\kimreader_ckvreader_data.sot [0], 
	\kimreader_ckvreader_data.eoi [0], \kimreader_ckvreader_data.eot [0], 
	\kimreader_ckvreader_data.id [3], \kimreader_ckvreader_data.id [2], 
	\kimreader_ckvreader_data.id [1], \kimreader_ckvreader_data.id [0], 
	\kimreader_ckvreader_data.tdata [63], 
	\kimreader_ckvreader_data.tdata [62], 
	\kimreader_ckvreader_data.tdata [61], 
	\kimreader_ckvreader_data.tdata [60], 
	\kimreader_ckvreader_data.tdata [59], 
	\kimreader_ckvreader_data.tdata [58], 
	\kimreader_ckvreader_data.tdata [57], 
	\kimreader_ckvreader_data.tdata [56], 
	\kimreader_ckvreader_data.tdata [55], 
	\kimreader_ckvreader_data.tdata [54], 
	\kimreader_ckvreader_data.tdata [53], 
	\kimreader_ckvreader_data.tdata [52], 
	\kimreader_ckvreader_data.tdata [51], 
	\kimreader_ckvreader_data.tdata [50], 
	\kimreader_ckvreader_data.tdata [49], 
	\kimreader_ckvreader_data.tdata [48], 
	\kimreader_ckvreader_data.tdata [47], 
	\kimreader_ckvreader_data.tdata [46], 
	\kimreader_ckvreader_data.tdata [45], 
	\kimreader_ckvreader_data.tdata [44], 
	\kimreader_ckvreader_data.tdata [43], 
	\kimreader_ckvreader_data.tdata [42], 
	\kimreader_ckvreader_data.tdata [41], 
	\kimreader_ckvreader_data.tdata [40], 
	\kimreader_ckvreader_data.tdata [39], 
	\kimreader_ckvreader_data.tdata [38], 
	\kimreader_ckvreader_data.tdata [37], 
	\kimreader_ckvreader_data.tdata [36], 
	\kimreader_ckvreader_data.tdata [35], 
	\kimreader_ckvreader_data.tdata [34], 
	\kimreader_ckvreader_data.tdata [33], 
	\kimreader_ckvreader_data.tdata [32], 
	\kimreader_ckvreader_data.tdata [31], 
	\kimreader_ckvreader_data.tdata [30], 
	\kimreader_ckvreader_data.tdata [29], 
	\kimreader_ckvreader_data.tdata [28], 
	\kimreader_ckvreader_data.tdata [27], 
	\kimreader_ckvreader_data.tdata [26], 
	\kimreader_ckvreader_data.tdata [25], 
	\kimreader_ckvreader_data.tdata [24], 
	\kimreader_ckvreader_data.tdata [23], 
	\kimreader_ckvreader_data.tdata [22], 
	\kimreader_ckvreader_data.tdata [21], 
	\kimreader_ckvreader_data.tdata [20], 
	\kimreader_ckvreader_data.tdata [19], 
	\kimreader_ckvreader_data.tdata [18], 
	\kimreader_ckvreader_data.tdata [17], 
	\kimreader_ckvreader_data.tdata [16], 
	\kimreader_ckvreader_data.tdata [15], 
	\kimreader_ckvreader_data.tdata [14], 
	\kimreader_ckvreader_data.tdata [13], 
	\kimreader_ckvreader_data.tdata [12], 
	\kimreader_ckvreader_data.tdata [11], 
	\kimreader_ckvreader_data.tdata [10], 
	\kimreader_ckvreader_data.tdata [9], 
	\kimreader_ckvreader_data.tdata [8], 
	\kimreader_ckvreader_data.tdata [7], 
	\kimreader_ckvreader_data.tdata [6], 
	\kimreader_ckvreader_data.tdata [5], 
	\kimreader_ckvreader_data.tdata [4], 
	\kimreader_ckvreader_data.tdata [3], 
	\kimreader_ckvreader_data.tdata [2], 
	\kimreader_ckvreader_data.tdata [1], 
	\kimreader_ckvreader_data.tdata [0]} ), drng_ack, kim_rd, kim_addr, 
	stat_req_with_expired_seed, stat_aux_key_type_0, stat_aux_key_type_1, 
	stat_aux_key_type_2, stat_aux_key_type_3, stat_aux_key_type_4, 
	stat_aux_key_type_5, stat_aux_key_type_6, stat_aux_key_type_7, 
	stat_aux_key_type_8, stat_aux_key_type_9, stat_aux_key_type_10, 
	stat_aux_key_type_11, stat_aux_key_type_12, stat_aux_key_type_13, 
	stat_aux_cmd_with_vf_pf_fail, clk, rst_n, parser_kimreader_valid, 
	.parser_kimreader_data( {\parser_kimreader_data.sot [0], 
	\parser_kimreader_data.eoi [0], \parser_kimreader_data.eot [0], 
	\parser_kimreader_data.id [3], \parser_kimreader_data.id [2], 
	\parser_kimreader_data.id [1], \parser_kimreader_data.id [0], 
	\parser_kimreader_data.tdata [63], \parser_kimreader_data.tdata [62], 
	\parser_kimreader_data.tdata [61], \parser_kimreader_data.tdata [60], 
	\parser_kimreader_data.tdata [59], \parser_kimreader_data.tdata [58], 
	\parser_kimreader_data.tdata [57], \parser_kimreader_data.tdata [56], 
	\parser_kimreader_data.tdata [55], \parser_kimreader_data.tdata [54], 
	\parser_kimreader_data.tdata [53], \parser_kimreader_data.tdata [52], 
	\parser_kimreader_data.tdata [51], \parser_kimreader_data.tdata [50], 
	\parser_kimreader_data.tdata [49], \parser_kimreader_data.tdata [48], 
	\parser_kimreader_data.tdata [47], \parser_kimreader_data.tdata [46], 
	\parser_kimreader_data.tdata [45], \parser_kimreader_data.tdata [44], 
	\parser_kimreader_data.tdata [43], \parser_kimreader_data.tdata [42], 
	\parser_kimreader_data.tdata [41], \parser_kimreader_data.tdata [40], 
	\parser_kimreader_data.tdata [39], \parser_kimreader_data.tdata [38], 
	\parser_kimreader_data.tdata [37], \parser_kimreader_data.tdata [36], 
	\parser_kimreader_data.tdata [35], \parser_kimreader_data.tdata [34], 
	\parser_kimreader_data.tdata [33], \parser_kimreader_data.tdata [32], 
	\parser_kimreader_data.tdata [31], \parser_kimreader_data.tdata [30], 
	\parser_kimreader_data.tdata [29], \parser_kimreader_data.tdata [28], 
	\parser_kimreader_data.tdata [27], \parser_kimreader_data.tdata [26], 
	\parser_kimreader_data.tdata [25], \parser_kimreader_data.tdata [24], 
	\parser_kimreader_data.tdata [23], \parser_kimreader_data.tdata [22], 
	\parser_kimreader_data.tdata [21], \parser_kimreader_data.tdata [20], 
	\parser_kimreader_data.tdata [19], \parser_kimreader_data.tdata [18], 
	\parser_kimreader_data.tdata [17], \parser_kimreader_data.tdata [16], 
	\parser_kimreader_data.tdata [15], \parser_kimreader_data.tdata [14], 
	\parser_kimreader_data.tdata [13], \parser_kimreader_data.tdata [12], 
	\parser_kimreader_data.tdata [11], \parser_kimreader_data.tdata [10], 
	\parser_kimreader_data.tdata [9], \parser_kimreader_data.tdata [8], 
	\parser_kimreader_data.tdata [7], \parser_kimreader_data.tdata [6], 
	\parser_kimreader_data.tdata [5], \parser_kimreader_data.tdata [4], 
	\parser_kimreader_data.tdata [3], \parser_kimreader_data.tdata [2], 
	\parser_kimreader_data.tdata [1], \parser_kimreader_data.tdata [0]} ), 
	ckvreader_kimreader_ack, drng_seed_expired, drng_health_fail, 
	drng_256_out, drng_valid, .kim_dout( {\kim_dout.valid [0], 
	\kim_dout.label_index [2], \kim_dout.label_index [1], 
	\kim_dout.label_index [0], \kim_dout.ckv_length [1], 
	\kim_dout.ckv_length [0], \kim_dout.ckv_pointer [14], 
	\kim_dout.ckv_pointer [13], \kim_dout.ckv_pointer [12], 
	\kim_dout.ckv_pointer [11], \kim_dout.ckv_pointer [10], 
	\kim_dout.ckv_pointer [9], \kim_dout.ckv_pointer [8], 
	\kim_dout.ckv_pointer [7], \kim_dout.ckv_pointer [6], 
	\kim_dout.ckv_pointer [5], \kim_dout.ckv_pointer [4], 
	\kim_dout.ckv_pointer [3], \kim_dout.ckv_pointer [2], 
	\kim_dout.ckv_pointer [1], \kim_dout.ckv_pointer [0], 
	\kim_dout.pf_num [3], \kim_dout.pf_num [2], \kim_dout.pf_num [1], 
	\kim_dout.pf_num [0], \kim_dout.vf_num [11], \kim_dout.vf_num [10], 
	\kim_dout.vf_num [9], \kim_dout.vf_num [8], \kim_dout.vf_num [7], 
	\kim_dout.vf_num [6], \kim_dout.vf_num [5], \kim_dout.vf_num [4], 
	\kim_dout.vf_num [3], \kim_dout.vf_num [2], \kim_dout.vf_num [1], 
	\kim_dout.vf_num [0], \kim_dout.vf_valid [0]} ), kim_mbe, 
	disable_unencrypted_keys);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output kimreader_parser_ack;
output kimreader_ckvreader_valid;
output [0:0] \kimreader_ckvreader_data.sot ;
output [0:0] \kimreader_ckvreader_data.eoi ;
output [0:0] \kimreader_ckvreader_data.eot ;
output [3:0] \kimreader_ckvreader_data.id ;
output [63:0] \kimreader_ckvreader_data.tdata ;
wire [70:0] kimreader_ckvreader_data;
output drng_ack;
output kim_rd;
output [13:0] kim_addr;
output stat_req_with_expired_seed;
output stat_aux_key_type_0;
output stat_aux_key_type_1;
output stat_aux_key_type_2;
output stat_aux_key_type_3;
output stat_aux_key_type_4;
output stat_aux_key_type_5;
output stat_aux_key_type_6;
output stat_aux_key_type_7;
output stat_aux_key_type_8;
output stat_aux_key_type_9;
output stat_aux_key_type_10;
output stat_aux_key_type_11;
output stat_aux_key_type_12;
output stat_aux_key_type_13;
output stat_aux_cmd_with_vf_pf_fail;
input clk;
input rst_n;
input parser_kimreader_valid;
input [0:0] \parser_kimreader_data.sot ;
input [0:0] \parser_kimreader_data.eoi ;
input [0:0] \parser_kimreader_data.eot ;
input [3:0] \parser_kimreader_data.id ;
input [63:0] \parser_kimreader_data.tdata ;
wire [70:0] parser_kimreader_data;
input ckvreader_kimreader_ack;
input drng_seed_expired;
input drng_health_fail;
input [127:0] drng_256_out;
input drng_valid;
input [0:0] \kim_dout.valid ;
input [2:0] \kim_dout.label_index ;
input [1:0] \kim_dout.ckv_length ;
input [14:0] \kim_dout.ckv_pointer ;
input [3:0] \kim_dout.pf_num ;
input [11:0] \kim_dout.vf_num ;
input [0:0] \kim_dout.vf_valid ;
wire [37:0] kim_dout;
input kim_mbe;
input disable_unencrypted_keys;
wire _zy_simnet_kimreader_parser_ack_0_w$;
wire _zy_simnet_kimreader_ckvreader_valid_1_w$;
wire [0:70] _zy_simnet_kimreader_ckvreader_data_2_w$;
wire _zy_simnet_drng_ack_3_w$;
wire _zy_simnet_kim_rd_4_w$;
wire [0:13] _zy_simnet_kim_addr_5_w$;
wire _zy_simnet_stat_req_with_expired_seed_6_w$;
wire _zy_simnet_stat_aux_key_type_0_7_w$;
wire _zy_simnet_stat_aux_key_type_1_8_w$;
wire _zy_simnet_stat_aux_key_type_2_9_w$;
wire _zy_simnet_stat_aux_key_type_3_10_w$;
wire _zy_simnet_stat_aux_key_type_4_11_w$;
wire _zy_simnet_stat_aux_key_type_5_12_w$;
wire _zy_simnet_stat_aux_key_type_6_13_w$;
wire _zy_simnet_stat_aux_key_type_7_14_w$;
wire _zy_simnet_stat_aux_key_type_8_15_w$;
wire _zy_simnet_stat_aux_key_type_9_16_w$;
wire _zy_simnet_stat_aux_key_type_10_17_w$;
wire _zy_simnet_stat_aux_key_type_11_18_w$;
wire _zy_simnet_stat_aux_key_type_12_19_w$;
wire _zy_simnet_stat_aux_key_type_13_20_w$;
wire _zy_simnet_stat_aux_cmd_with_vf_pf_fail_21_w$;
wire _zy_sva_disable_unenc_keys_1_reset_or;
wire _zy_sva_enable_unenc_keys_2_reset_or;
wire _zy_sva_disable_unenc_keys_3_reset_or;
wire _zy_sva_enable_unenc_keys_4_reset_or;
wire _zy_sva_disable_unenc_keys_5_reset_or;
wire _zy_sva_enable_unenc_keys_6_reset_or;
wire _zy_sva_disable_unenc_keys_7_reset_or;
wire _zy_sva_enable_unenc_keys_8_reset_or;
wire _zy_sva_disable_unenc_keys_9_reset_or;
wire _zy_sva_enable_unenc_keys_10_reset_or;
wire _zy_sva_b0_t;
wire _zy_sva_b1_t;
wire _zy_sva_b2_t;
wire _zy_sva_b3_t;
wire _zy_sva_b4_t;
wire _zy_sva_b5_t;
wire _zy_sva_b6_t;
wire _zy_sva_b7_t;
wire _zy_sva_b8_t;
wire _zy_sva_b9_t;
wire [2:0] cur_state;
wire [2:0] nxt_state;
wire [13:0] dek_ref_q;
wire [13:0] dak_ref_q;
wire dek_is_kdf_key_q;
wire dak_is_kdf_key_q;
wire [7:0] kim_errors_q;
wire [37:0] dek_kim_entry_q;
wire [37:0] dak_kim_entry_q;
wire dek_kim_mbe_q;
wire dak_kim_mbe_q;
wire kim_rd_q;
wire [63:0] tlv_word0;
wire [63:0] tlv_word8;
wire [63:0] tlv_word9;
wire [55:0] tlv_word42;
wire [31:0] aux_key_ctrl;
wire [5:0] aux_key_type;
`_2_ wire [0:0] _zy_sva_disable_unenc_keys_1_ccheck;
`_2_ wire [0:0] _zy_sva_disable_unenc_keys_1_cpass;
`_2_ wire _zy_sva_b0;
`_2_ wire [0:0] _zy_sva_enable_unenc_keys_2_ccheck;
`_2_ wire [0:0] _zy_sva_enable_unenc_keys_2_cpass;
`_2_ wire _zy_sva_b1;
`_2_ wire [0:0] _zy_sva_disable_unenc_keys_3_ccheck;
`_2_ wire [0:0] _zy_sva_disable_unenc_keys_3_cpass;
`_2_ wire _zy_sva_b2;
`_2_ wire [0:0] _zy_sva_enable_unenc_keys_4_ccheck;
`_2_ wire [0:0] _zy_sva_enable_unenc_keys_4_cpass;
`_2_ wire _zy_sva_b3;
`_2_ wire [0:0] _zy_sva_disable_unenc_keys_5_ccheck;
`_2_ wire [0:0] _zy_sva_disable_unenc_keys_5_cpass;
`_2_ wire _zy_sva_b4;
`_2_ wire [0:0] _zy_sva_enable_unenc_keys_6_ccheck;
`_2_ wire [0:0] _zy_sva_enable_unenc_keys_6_cpass;
`_2_ wire _zy_sva_b5;
`_2_ wire [0:0] _zy_sva_disable_unenc_keys_7_ccheck;
`_2_ wire [0:0] _zy_sva_disable_unenc_keys_7_cpass;
`_2_ wire _zy_sva_b6;
`_2_ wire [0:0] _zy_sva_enable_unenc_keys_8_ccheck;
`_2_ wire [0:0] _zy_sva_enable_unenc_keys_8_cpass;
`_2_ wire _zy_sva_b7;
`_2_ wire [0:0] _zy_sva_disable_unenc_keys_9_ccheck;
`_2_ wire [0:0] _zy_sva_disable_unenc_keys_9_cpass;
`_2_ wire _zy_sva_b8;
`_2_ wire [0:0] _zy_sva_enable_unenc_keys_10_ccheck;
`_2_ wire [0:0] _zy_sva_enable_unenc_keys_10_cpass;
`_2_ wire _zy_sva_b9;
wire _zyL438_tfiRv4;
wire _zyL444_tfiRv5;
wire _zyL468_tfiRv6;
wire _zyL473_tfiRv7;
supply0 n379;
supply1 n646;
wire [0:0] \dek_kim_entry_q.valid ;
wire [2:0] \dek_kim_entry_q.label_index ;
wire [1:0] \dek_kim_entry_q.ckv_length ;
wire [14:0] \dek_kim_entry_q.ckv_pointer ;
wire [3:0] \dek_kim_entry_q.pf_num ;
wire [11:0] \dek_kim_entry_q.vf_num ;
wire [0:0] \dek_kim_entry_q.vf_valid ;
wire [0:0] \dak_kim_entry_q.valid ;
wire [2:0] \dak_kim_entry_q.label_index ;
wire [1:0] \dak_kim_entry_q.ckv_length ;
wire [14:0] \dak_kim_entry_q.ckv_pointer ;
wire [3:0] \dak_kim_entry_q.pf_num ;
wire [11:0] \dak_kim_entry_q.vf_num ;
wire [0:0] \dak_kim_entry_q.vf_valid ;
wire [1:0] \tlv_word0.tlv_bip2 ;
wire [12:0] \tlv_word0.resv0 ;
wire [0:0] \tlv_word0.kdf_dek_iter ;
wire [0:0] \tlv_word0.keyless_algos ;
wire [0:0] \tlv_word0.needs_dek ;
wire [0:0] \tlv_word0.needs_dak ;
wire [5:0] \tlv_word0.key_type ;
wire [10:0] \tlv_word0.tlv_frame_num ;
wire [3:0] \tlv_word0.tlv_eng_id ;
wire [7:0] \tlv_word0.tlv_seq_num ;
wire [7:0] \tlv_word0.tlv_len ;
wire [7:0] \tlv_word0.tlv_type ;
wire [0:0] \tlv_word8.dek_kim_entry.valid ;
wire [2:0] \tlv_word8.dek_kim_entry.label_index ;
wire [1:0] \tlv_word8.dek_kim_entry.ckv_length ;
wire [14:0] \tlv_word8.dek_kim_entry.ckv_pointer ;
wire [3:0] \tlv_word8.dek_kim_entry.pf_num ;
wire [11:0] \tlv_word8.dek_kim_entry.vf_num ;
wire [0:0] \tlv_word8.dek_kim_entry.vf_valid ;
wire [5:0] \tlv_word8.unused ;
wire [0:0] \tlv_word8.missing_iv ;
wire [0:0] \tlv_word8.missing_guid ;
wire [0:0] \tlv_word8.validate_dek ;
wire [0:0] \tlv_word8.vf_valid ;
wire [3:0] \tlv_word8.pf_num ;
wire [11:0] \tlv_word8.vf_num ;
wire [0:0] \tlv_word9.dak_kim_entry.valid ;
wire [2:0] \tlv_word9.dak_kim_entry.label_index ;
wire [1:0] \tlv_word9.dak_kim_entry.ckv_length ;
wire [14:0] \tlv_word9.dak_kim_entry.ckv_pointer ;
wire [3:0] \tlv_word9.dak_kim_entry.pf_num ;
wire [11:0] \tlv_word9.dak_kim_entry.vf_num ;
wire [0:0] \tlv_word9.dak_kim_entry.vf_valid ;
wire [7:0] \tlv_word9.unused ;
wire [0:0] \tlv_word9.validate_dak ;
wire [0:0] \tlv_word9.vf_valid ;
wire [3:0] \tlv_word9.pf_num ;
wire [11:0] \tlv_word9.vf_num ;
wire [0:0] \tlv_word42.corrupt_crc32 ;
wire [46:0] \tlv_word42.unused ;
wire [7:0] \tlv_word42.error_code ;
wire [0:0] \aux_key_ctrl.dak_key_op ;
wire [13:0] \aux_key_ctrl.dak_key_ref ;
wire [1:0] \aux_key_ctrl.kdf_mode ;
wire [0:0] \aux_key_ctrl.dek_key_op ;
wire [13:0] \aux_key_ctrl.dek_key_ref ;
tran (kimreader_ckvreader_data[70], \kimreader_ckvreader_data.sot [0]);
tran (kimreader_ckvreader_data[69], \kimreader_ckvreader_data.eoi [0]);
tran (kimreader_ckvreader_data[68], \kimreader_ckvreader_data.eot [0]);
tran (kimreader_ckvreader_data[67], \kimreader_ckvreader_data.id [3]);
tran (kimreader_ckvreader_data[66], \kimreader_ckvreader_data.id [2]);
tran (kimreader_ckvreader_data[65], \kimreader_ckvreader_data.id [1]);
tran (kimreader_ckvreader_data[64], \kimreader_ckvreader_data.id [0]);
tran (kimreader_ckvreader_data[63], \kimreader_ckvreader_data.tdata [63]);
tran (kimreader_ckvreader_data[62], \kimreader_ckvreader_data.tdata [62]);
tran (kimreader_ckvreader_data[61], \kimreader_ckvreader_data.tdata [61]);
tran (kimreader_ckvreader_data[60], \kimreader_ckvreader_data.tdata [60]);
tran (kimreader_ckvreader_data[59], \kimreader_ckvreader_data.tdata [59]);
tran (kimreader_ckvreader_data[58], \kimreader_ckvreader_data.tdata [58]);
tran (kimreader_ckvreader_data[57], \kimreader_ckvreader_data.tdata [57]);
tran (kimreader_ckvreader_data[56], \kimreader_ckvreader_data.tdata [56]);
tran (kimreader_ckvreader_data[55], \kimreader_ckvreader_data.tdata [55]);
tran (kimreader_ckvreader_data[54], \kimreader_ckvreader_data.tdata [54]);
tran (kimreader_ckvreader_data[53], \kimreader_ckvreader_data.tdata [53]);
tran (kimreader_ckvreader_data[52], \kimreader_ckvreader_data.tdata [52]);
tran (kimreader_ckvreader_data[51], \kimreader_ckvreader_data.tdata [51]);
tran (kimreader_ckvreader_data[50], \kimreader_ckvreader_data.tdata [50]);
tran (kimreader_ckvreader_data[49], \kimreader_ckvreader_data.tdata [49]);
tran (kimreader_ckvreader_data[48], \kimreader_ckvreader_data.tdata [48]);
tran (kimreader_ckvreader_data[47], \kimreader_ckvreader_data.tdata [47]);
tran (kimreader_ckvreader_data[46], \kimreader_ckvreader_data.tdata [46]);
tran (kimreader_ckvreader_data[45], \kimreader_ckvreader_data.tdata [45]);
tran (kimreader_ckvreader_data[44], \kimreader_ckvreader_data.tdata [44]);
tran (kimreader_ckvreader_data[43], \kimreader_ckvreader_data.tdata [43]);
tran (kimreader_ckvreader_data[42], \kimreader_ckvreader_data.tdata [42]);
tran (kimreader_ckvreader_data[41], \kimreader_ckvreader_data.tdata [41]);
tran (kimreader_ckvreader_data[40], \kimreader_ckvreader_data.tdata [40]);
tran (kimreader_ckvreader_data[39], \kimreader_ckvreader_data.tdata [39]);
tran (kimreader_ckvreader_data[38], \kimreader_ckvreader_data.tdata [38]);
tran (kimreader_ckvreader_data[37], \kimreader_ckvreader_data.tdata [37]);
tran (kimreader_ckvreader_data[36], \kimreader_ckvreader_data.tdata [36]);
tran (kimreader_ckvreader_data[35], \kimreader_ckvreader_data.tdata [35]);
tran (kimreader_ckvreader_data[34], \kimreader_ckvreader_data.tdata [34]);
tran (kimreader_ckvreader_data[33], \kimreader_ckvreader_data.tdata [33]);
tran (kimreader_ckvreader_data[32], \kimreader_ckvreader_data.tdata [32]);
tran (kimreader_ckvreader_data[31], \kimreader_ckvreader_data.tdata [31]);
tran (kimreader_ckvreader_data[30], \kimreader_ckvreader_data.tdata [30]);
tran (kimreader_ckvreader_data[29], \kimreader_ckvreader_data.tdata [29]);
tran (kimreader_ckvreader_data[28], \kimreader_ckvreader_data.tdata [28]);
tran (kimreader_ckvreader_data[27], \kimreader_ckvreader_data.tdata [27]);
tran (kimreader_ckvreader_data[26], \kimreader_ckvreader_data.tdata [26]);
tran (kimreader_ckvreader_data[25], \kimreader_ckvreader_data.tdata [25]);
tran (kimreader_ckvreader_data[24], \kimreader_ckvreader_data.tdata [24]);
tran (kimreader_ckvreader_data[23], \kimreader_ckvreader_data.tdata [23]);
tran (kimreader_ckvreader_data[22], \kimreader_ckvreader_data.tdata [22]);
tran (kimreader_ckvreader_data[21], \kimreader_ckvreader_data.tdata [21]);
tran (kimreader_ckvreader_data[20], \kimreader_ckvreader_data.tdata [20]);
tran (kimreader_ckvreader_data[19], \kimreader_ckvreader_data.tdata [19]);
tran (kimreader_ckvreader_data[18], \kimreader_ckvreader_data.tdata [18]);
tran (kimreader_ckvreader_data[17], \kimreader_ckvreader_data.tdata [17]);
tran (kimreader_ckvreader_data[16], \kimreader_ckvreader_data.tdata [16]);
tran (kimreader_ckvreader_data[15], \kimreader_ckvreader_data.tdata [15]);
tran (kimreader_ckvreader_data[14], \kimreader_ckvreader_data.tdata [14]);
tran (kimreader_ckvreader_data[13], \kimreader_ckvreader_data.tdata [13]);
tran (kimreader_ckvreader_data[12], \kimreader_ckvreader_data.tdata [12]);
tran (kimreader_ckvreader_data[11], \kimreader_ckvreader_data.tdata [11]);
tran (kimreader_ckvreader_data[10], \kimreader_ckvreader_data.tdata [10]);
tran (kimreader_ckvreader_data[9], \kimreader_ckvreader_data.tdata [9]);
tran (kimreader_ckvreader_data[8], \kimreader_ckvreader_data.tdata [8]);
tran (kimreader_ckvreader_data[7], \kimreader_ckvreader_data.tdata [7]);
tran (kimreader_ckvreader_data[6], \kimreader_ckvreader_data.tdata [6]);
tran (kimreader_ckvreader_data[5], \kimreader_ckvreader_data.tdata [5]);
tran (kimreader_ckvreader_data[4], \kimreader_ckvreader_data.tdata [4]);
tran (kimreader_ckvreader_data[3], \kimreader_ckvreader_data.tdata [3]);
tran (kimreader_ckvreader_data[2], \kimreader_ckvreader_data.tdata [2]);
tran (kimreader_ckvreader_data[1], \kimreader_ckvreader_data.tdata [1]);
tran (kimreader_ckvreader_data[0], \kimreader_ckvreader_data.tdata [0]);
tran (parser_kimreader_data[70], \parser_kimreader_data.sot [0]);
tran (parser_kimreader_data[69], \parser_kimreader_data.eoi [0]);
tran (parser_kimreader_data[68], \parser_kimreader_data.eot [0]);
tran (parser_kimreader_data[67], \parser_kimreader_data.id [3]);
tran (parser_kimreader_data[66], \parser_kimreader_data.id [2]);
tran (parser_kimreader_data[65], \parser_kimreader_data.id [1]);
tran (parser_kimreader_data[64], \parser_kimreader_data.id [0]);
tran (parser_kimreader_data[63], \parser_kimreader_data.tdata [63]);
tran (parser_kimreader_data[62], \parser_kimreader_data.tdata [62]);
tran (parser_kimreader_data[61], \parser_kimreader_data.tdata [61]);
tran (parser_kimreader_data[60], \parser_kimreader_data.tdata [60]);
tran (parser_kimreader_data[59], \parser_kimreader_data.tdata [59]);
tran (parser_kimreader_data[58], \parser_kimreader_data.tdata [58]);
tran (parser_kimreader_data[57], \parser_kimreader_data.tdata [57]);
tran (parser_kimreader_data[56], \parser_kimreader_data.tdata [56]);
tran (parser_kimreader_data[55], \parser_kimreader_data.tdata [55]);
tran (parser_kimreader_data[54], \parser_kimreader_data.tdata [54]);
tran (parser_kimreader_data[53], \parser_kimreader_data.tdata [53]);
tran (parser_kimreader_data[52], \parser_kimreader_data.tdata [52]);
tran (parser_kimreader_data[51], \parser_kimreader_data.tdata [51]);
tran (parser_kimreader_data[50], \parser_kimreader_data.tdata [50]);
tran (parser_kimreader_data[49], \parser_kimreader_data.tdata [49]);
tran (parser_kimreader_data[48], \parser_kimreader_data.tdata [48]);
tran (parser_kimreader_data[47], \parser_kimreader_data.tdata [47]);
tran (parser_kimreader_data[46], \parser_kimreader_data.tdata [46]);
tran (parser_kimreader_data[45], \parser_kimreader_data.tdata [45]);
tran (parser_kimreader_data[44], \parser_kimreader_data.tdata [44]);
tran (parser_kimreader_data[43], \parser_kimreader_data.tdata [43]);
tran (parser_kimreader_data[42], \parser_kimreader_data.tdata [42]);
tran (parser_kimreader_data[41], \parser_kimreader_data.tdata [41]);
tran (parser_kimreader_data[40], \parser_kimreader_data.tdata [40]);
tran (parser_kimreader_data[39], \parser_kimreader_data.tdata [39]);
tran (parser_kimreader_data[38], \parser_kimreader_data.tdata [38]);
tran (parser_kimreader_data[37], \parser_kimreader_data.tdata [37]);
tran (parser_kimreader_data[36], \parser_kimreader_data.tdata [36]);
tran (parser_kimreader_data[35], \parser_kimreader_data.tdata [35]);
tran (parser_kimreader_data[34], \parser_kimreader_data.tdata [34]);
tran (parser_kimreader_data[33], \parser_kimreader_data.tdata [33]);
tran (parser_kimreader_data[32], \parser_kimreader_data.tdata [32]);
tran (parser_kimreader_data[31], \parser_kimreader_data.tdata [31]);
tran (parser_kimreader_data[30], \parser_kimreader_data.tdata [30]);
tran (parser_kimreader_data[29], \parser_kimreader_data.tdata [29]);
tran (parser_kimreader_data[28], \parser_kimreader_data.tdata [28]);
tran (parser_kimreader_data[27], \parser_kimreader_data.tdata [27]);
tran (parser_kimreader_data[26], \parser_kimreader_data.tdata [26]);
tran (parser_kimreader_data[25], \parser_kimreader_data.tdata [25]);
tran (parser_kimreader_data[24], \parser_kimreader_data.tdata [24]);
tran (parser_kimreader_data[23], \parser_kimreader_data.tdata [23]);
tran (parser_kimreader_data[22], \parser_kimreader_data.tdata [22]);
tran (parser_kimreader_data[21], \parser_kimreader_data.tdata [21]);
tran (parser_kimreader_data[20], \parser_kimreader_data.tdata [20]);
tran (parser_kimreader_data[19], \parser_kimreader_data.tdata [19]);
tran (parser_kimreader_data[18], \parser_kimreader_data.tdata [18]);
tran (parser_kimreader_data[17], \parser_kimreader_data.tdata [17]);
tran (parser_kimreader_data[16], \parser_kimreader_data.tdata [16]);
tran (parser_kimreader_data[15], \parser_kimreader_data.tdata [15]);
tran (parser_kimreader_data[14], \parser_kimreader_data.tdata [14]);
tran (parser_kimreader_data[13], \parser_kimreader_data.tdata [13]);
tran (parser_kimreader_data[12], \parser_kimreader_data.tdata [12]);
tran (parser_kimreader_data[11], \parser_kimreader_data.tdata [11]);
tran (parser_kimreader_data[10], \parser_kimreader_data.tdata [10]);
tran (parser_kimreader_data[9], \parser_kimreader_data.tdata [9]);
tran (parser_kimreader_data[8], \parser_kimreader_data.tdata [8]);
tran (parser_kimreader_data[7], \parser_kimreader_data.tdata [7]);
tran (parser_kimreader_data[6], \parser_kimreader_data.tdata [6]);
tran (parser_kimreader_data[5], \parser_kimreader_data.tdata [5]);
tran (parser_kimreader_data[4], \parser_kimreader_data.tdata [4]);
tran (parser_kimreader_data[3], \parser_kimreader_data.tdata [3]);
tran (parser_kimreader_data[2], \parser_kimreader_data.tdata [2]);
tran (parser_kimreader_data[1], \parser_kimreader_data.tdata [1]);
tran (parser_kimreader_data[0], \parser_kimreader_data.tdata [0]);
tran (kim_dout[37], \kim_dout.valid [0]);
tran (kim_dout[36], \kim_dout.label_index [2]);
tran (kim_dout[35], \kim_dout.label_index [1]);
tran (kim_dout[34], \kim_dout.label_index [0]);
tran (kim_dout[33], \kim_dout.ckv_length [1]);
tran (kim_dout[32], \kim_dout.ckv_length [0]);
tran (kim_dout[31], \kim_dout.ckv_pointer [14]);
tran (kim_dout[30], \kim_dout.ckv_pointer [13]);
tran (kim_dout[29], \kim_dout.ckv_pointer [12]);
tran (kim_dout[28], \kim_dout.ckv_pointer [11]);
tran (kim_dout[27], \kim_dout.ckv_pointer [10]);
tran (kim_dout[26], \kim_dout.ckv_pointer [9]);
tran (kim_dout[25], \kim_dout.ckv_pointer [8]);
tran (kim_dout[24], \kim_dout.ckv_pointer [7]);
tran (kim_dout[23], \kim_dout.ckv_pointer [6]);
tran (kim_dout[22], \kim_dout.ckv_pointer [5]);
tran (kim_dout[21], \kim_dout.ckv_pointer [4]);
tran (kim_dout[20], \kim_dout.ckv_pointer [3]);
tran (kim_dout[19], \kim_dout.ckv_pointer [2]);
tran (kim_dout[18], \kim_dout.ckv_pointer [1]);
tran (kim_dout[17], \kim_dout.ckv_pointer [0]);
tran (kim_dout[16], \kim_dout.pf_num [3]);
tran (kim_dout[15], \kim_dout.pf_num [2]);
tran (kim_dout[14], \kim_dout.pf_num [1]);
tran (kim_dout[13], \kim_dout.pf_num [0]);
tran (kim_dout[12], \kim_dout.vf_num [11]);
tran (kim_dout[11], \kim_dout.vf_num [10]);
tran (kim_dout[10], \kim_dout.vf_num [9]);
tran (kim_dout[9], \kim_dout.vf_num [8]);
tran (kim_dout[8], \kim_dout.vf_num [7]);
tran (kim_dout[7], \kim_dout.vf_num [6]);
tran (kim_dout[6], \kim_dout.vf_num [5]);
tran (kim_dout[5], \kim_dout.vf_num [4]);
tran (kim_dout[4], \kim_dout.vf_num [3]);
tran (kim_dout[3], \kim_dout.vf_num [2]);
tran (kim_dout[2], \kim_dout.vf_num [1]);
tran (kim_dout[1], \kim_dout.vf_num [0]);
tran (kim_dout[0], \kim_dout.vf_valid [0]);
tran (tlv_word0[0], \tlv_word0.tlv_type [0]);
tran (aux_key_ctrl[0], \aux_key_ctrl.dek_key_ref [0]);
tran (tlv_word0[1], \tlv_word0.tlv_type [1]);
tran (aux_key_ctrl[1], \aux_key_ctrl.dek_key_ref [1]);
tran (tlv_word0[2], \tlv_word0.tlv_type [2]);
tran (aux_key_ctrl[2], \aux_key_ctrl.dek_key_ref [2]);
tran (tlv_word0[3], \tlv_word0.tlv_type [3]);
tran (aux_key_ctrl[3], \aux_key_ctrl.dek_key_ref [3]);
tran (tlv_word0[4], \tlv_word0.tlv_type [4]);
tran (aux_key_ctrl[4], \aux_key_ctrl.dek_key_ref [4]);
tran (tlv_word0[5], \tlv_word0.tlv_type [5]);
tran (aux_key_ctrl[5], \aux_key_ctrl.dek_key_ref [5]);
tran (tlv_word0[6], \tlv_word0.tlv_type [6]);
tran (aux_key_ctrl[6], \aux_key_ctrl.dek_key_ref [6]);
tran (tlv_word0[7], \tlv_word0.tlv_type [7]);
tran (aux_key_ctrl[7], \aux_key_ctrl.dek_key_ref [7]);
tran (tlv_word0[8], \tlv_word0.tlv_len [0]);
tran (tlv_word42[8], \tlv_word42.unused [0]);
tran (aux_key_ctrl[8], \aux_key_ctrl.dek_key_ref [8]);
tran (tlv_word0[9], \tlv_word0.tlv_len [1]);
tran (tlv_word42[9], \tlv_word42.unused [1]);
tran (aux_key_ctrl[9], \aux_key_ctrl.dek_key_ref [9]);
tran (tlv_word0[10], \tlv_word0.tlv_len [2]);
tran (tlv_word42[10], \tlv_word42.unused [2]);
tran (aux_key_ctrl[10], \aux_key_ctrl.dek_key_ref [10]);
tran (tlv_word0[11], \tlv_word0.tlv_len [3]);
tran (tlv_word42[11], \tlv_word42.unused [3]);
tran (aux_key_ctrl[11], \aux_key_ctrl.dek_key_ref [11]);
tran (tlv_word0[12], \tlv_word0.tlv_len [4]);
tran (tlv_word42[12], \tlv_word42.unused [4]);
tran (aux_key_ctrl[12], \aux_key_ctrl.dek_key_ref [12]);
tran (tlv_word0[13], \tlv_word0.tlv_len [5]);
tran (tlv_word42[13], \tlv_word42.unused [5]);
tran (aux_key_ctrl[13], \aux_key_ctrl.dek_key_ref [13]);
tran (tlv_word0[14], \tlv_word0.tlv_len [6]);
tran (tlv_word42[14], \tlv_word42.unused [6]);
tran (aux_key_ctrl[14], \aux_key_ctrl.dek_key_op [0]);
tran (tlv_word0[15], \tlv_word0.tlv_len [7]);
tran (tlv_word42[15], \tlv_word42.unused [7]);
tran (aux_key_ctrl[15], \aux_key_ctrl.kdf_mode [0]);
tran (tlv_word0[16], \tlv_word0.tlv_seq_num [0]);
tran (tlv_word42[16], \tlv_word42.unused [8]);
tran (aux_key_ctrl[16], \aux_key_ctrl.kdf_mode [1]);
tran (tlv_word0[17], \tlv_word0.tlv_seq_num [1]);
tran (tlv_word42[17], \tlv_word42.unused [9]);
tran (aux_key_ctrl[17], \aux_key_ctrl.dak_key_ref [0]);
tran (tlv_word0[18], \tlv_word0.tlv_seq_num [2]);
tran (tlv_word42[18], \tlv_word42.unused [10]);
tran (aux_key_ctrl[18], \aux_key_ctrl.dak_key_ref [1]);
tran (tlv_word0[19], \tlv_word0.tlv_seq_num [3]);
tran (tlv_word42[19], \tlv_word42.unused [11]);
tran (aux_key_ctrl[19], \aux_key_ctrl.dak_key_ref [2]);
tran (tlv_word0[20], \tlv_word0.tlv_seq_num [4]);
tran (tlv_word42[20], \tlv_word42.unused [12]);
tran (aux_key_ctrl[20], \aux_key_ctrl.dak_key_ref [3]);
tran (tlv_word0[21], \tlv_word0.tlv_seq_num [5]);
tran (tlv_word42[21], \tlv_word42.unused [13]);
tran (aux_key_ctrl[21], \aux_key_ctrl.dak_key_ref [4]);
tran (tlv_word0[22], \tlv_word0.tlv_seq_num [6]);
tran (tlv_word42[22], \tlv_word42.unused [14]);
tran (aux_key_ctrl[22], \aux_key_ctrl.dak_key_ref [5]);
tran (tlv_word0[23], \tlv_word0.tlv_seq_num [7]);
tran (tlv_word42[23], \tlv_word42.unused [15]);
tran (aux_key_ctrl[23], \aux_key_ctrl.dak_key_ref [6]);
tran (tlv_word0[24], \tlv_word0.tlv_eng_id [0]);
tran (tlv_word42[24], \tlv_word42.unused [16]);
tran (aux_key_ctrl[24], \aux_key_ctrl.dak_key_ref [7]);
tran (tlv_word0[25], \tlv_word0.tlv_eng_id [1]);
tran (tlv_word42[25], \tlv_word42.unused [17]);
tran (aux_key_ctrl[25], \aux_key_ctrl.dak_key_ref [8]);
tran (tlv_word0[26], \tlv_word0.tlv_eng_id [2]);
tran (tlv_word42[26], \tlv_word42.unused [18]);
tran (aux_key_ctrl[26], \aux_key_ctrl.dak_key_ref [9]);
tran (tlv_word0[27], \tlv_word0.tlv_eng_id [3]);
tran (tlv_word42[27], \tlv_word42.unused [19]);
tran (aux_key_ctrl[27], \aux_key_ctrl.dak_key_ref [10]);
tran (tlv_word0[28], \tlv_word0.tlv_frame_num [0]);
tran (tlv_word42[28], \tlv_word42.unused [20]);
tran (aux_key_ctrl[28], \aux_key_ctrl.dak_key_ref [11]);
tran (tlv_word0[29], \tlv_word0.tlv_frame_num [1]);
tran (tlv_word42[29], \tlv_word42.unused [21]);
tran (aux_key_ctrl[29], \aux_key_ctrl.dak_key_ref [12]);
tran (tlv_word0[30], \tlv_word0.tlv_frame_num [2]);
tran (tlv_word42[30], \tlv_word42.unused [22]);
tran (aux_key_ctrl[30], \aux_key_ctrl.dak_key_ref [13]);
tran (tlv_word0[31], \tlv_word0.tlv_frame_num [3]);
tran (tlv_word42[31], \tlv_word42.unused [23]);
tran (aux_key_ctrl[31], \aux_key_ctrl.dak_key_op [0]);
tran (tlv_word42[0], \tlv_word42.error_code [0]);
tran (tlv_word42[1], \tlv_word42.error_code [1]);
tran (tlv_word42[2], \tlv_word42.error_code [2]);
tran (tlv_word42[3], \tlv_word42.error_code [3]);
tran (tlv_word42[4], \tlv_word42.error_code [4]);
tran (tlv_word42[5], \tlv_word42.error_code [5]);
tran (tlv_word42[6], \tlv_word42.error_code [6]);
tran (tlv_word42[7], \tlv_word42.error_code [7]);
tran (tlv_word0[32], \tlv_word0.tlv_frame_num [4]);
tran (tlv_word42[32], \tlv_word42.unused [24]);
tran (tlv_word0[33], \tlv_word0.tlv_frame_num [5]);
tran (tlv_word42[33], \tlv_word42.unused [25]);
tran (tlv_word0[34], \tlv_word0.tlv_frame_num [6]);
tran (tlv_word42[34], \tlv_word42.unused [26]);
tran (tlv_word0[35], \tlv_word0.tlv_frame_num [7]);
tran (tlv_word42[35], \tlv_word42.unused [27]);
tran (tlv_word0[36], \tlv_word0.tlv_frame_num [8]);
tran (tlv_word42[36], \tlv_word42.unused [28]);
tran (tlv_word0[37], \tlv_word0.tlv_frame_num [9]);
tran (tlv_word42[37], \tlv_word42.unused [29]);
tran (tlv_word0[38], \tlv_word0.tlv_frame_num [10]);
tran (tlv_word42[38], \tlv_word42.unused [30]);
tran (tlv_word0[39], \tlv_word0.key_type [0]);
tran (tlv_word42[39], \tlv_word42.unused [31]);
tran (tlv_word0[40], \tlv_word0.key_type [1]);
tran (tlv_word42[40], \tlv_word42.unused [32]);
tran (tlv_word0[41], \tlv_word0.key_type [2]);
tran (tlv_word42[41], \tlv_word42.unused [33]);
tran (tlv_word0[42], \tlv_word0.key_type [3]);
tran (tlv_word42[42], \tlv_word42.unused [34]);
tran (tlv_word0[43], \tlv_word0.key_type [4]);
tran (tlv_word42[43], \tlv_word42.unused [35]);
tran (tlv_word0[44], \tlv_word0.key_type [5]);
tran (tlv_word42[44], \tlv_word42.unused [36]);
tran (tlv_word0[45], \tlv_word0.needs_dak [0]);
tran (tlv_word42[45], \tlv_word42.unused [37]);
tran (tlv_word0[46], \tlv_word0.needs_dek [0]);
tran (tlv_word42[46], \tlv_word42.unused [38]);
tran (tlv_word0[47], \tlv_word0.keyless_algos [0]);
tran (tlv_word42[47], \tlv_word42.unused [39]);
tran (tlv_word0[48], \tlv_word0.kdf_dek_iter [0]);
tran (tlv_word42[48], \tlv_word42.unused [40]);
tran (tlv_word0[49], \tlv_word0.resv0 [0]);
tran (tlv_word42[49], \tlv_word42.unused [41]);
tran (tlv_word0[50], \tlv_word0.resv0 [1]);
tran (tlv_word42[50], \tlv_word42.unused [42]);
tran (tlv_word0[51], \tlv_word0.resv0 [2]);
tran (tlv_word42[51], \tlv_word42.unused [43]);
tran (tlv_word0[52], \tlv_word0.resv0 [3]);
tran (tlv_word42[52], \tlv_word42.unused [44]);
tran (tlv_word0[53], \tlv_word0.resv0 [4]);
tran (tlv_word42[53], \tlv_word42.unused [45]);
tran (tlv_word0[54], \tlv_word0.resv0 [5]);
tran (tlv_word42[54], \tlv_word42.unused [46]);
tran (tlv_word0[55], \tlv_word0.resv0 [6]);
tran (tlv_word42[55], \tlv_word42.corrupt_crc32 [0]);
tran (tlv_word9[17], \tlv_word9.validate_dak [0]);
tran (tlv_word9[18], \tlv_word9.unused [0]);
tran (tlv_word9[19], \tlv_word9.unused [1]);
tran (tlv_word8[0], \tlv_word8.vf_num [0]);
tran (tlv_word8[1], \tlv_word8.vf_num [1]);
tran (tlv_word8[2], \tlv_word8.vf_num [2]);
tran (tlv_word8[3], \tlv_word8.vf_num [3]);
tran (tlv_word8[4], \tlv_word8.vf_num [4]);
tran (tlv_word8[5], \tlv_word8.vf_num [5]);
tran (tlv_word8[6], \tlv_word8.vf_num [6]);
tran (tlv_word8[7], \tlv_word8.vf_num [7]);
tran (tlv_word8[8], \tlv_word8.vf_num [8]);
tran (tlv_word8[9], \tlv_word8.vf_num [9]);
tran (tlv_word8[10], \tlv_word8.vf_num [10]);
tran (tlv_word8[11], \tlv_word8.vf_num [11]);
tran (tlv_word8[12], \tlv_word8.pf_num [0]);
tran (tlv_word8[13], \tlv_word8.pf_num [1]);
tran (tlv_word8[14], \tlv_word8.pf_num [2]);
tran (tlv_word8[15], \tlv_word8.pf_num [3]);
tran (tlv_word8[16], \tlv_word8.vf_valid [0]);
tran (tlv_word8[20], \tlv_word8.unused [0]);
tran (tlv_word8[21], \tlv_word8.unused [1]);
tran (tlv_word8[22], \tlv_word8.unused [2]);
tran (tlv_word8[23], \tlv_word8.unused [3]);
tran (tlv_word8[24], \tlv_word8.unused [4]);
tran (tlv_word8[25], \tlv_word8.unused [5]);
tran (tlv_word0[56], \tlv_word0.resv0 [7]);
tran (tlv_word0[57], \tlv_word0.resv0 [8]);
tran (tlv_word0[58], \tlv_word0.resv0 [9]);
tran (tlv_word0[59], \tlv_word0.resv0 [10]);
tran (tlv_word0[60], \tlv_word0.resv0 [11]);
tran (tlv_word0[61], \tlv_word0.resv0 [12]);
tran (tlv_word0[62], \tlv_word0.tlv_bip2 [0]);
tran (tlv_word0[63], \tlv_word0.tlv_bip2 [1]);
tran (tlv_word8[63], \tlv_word8.dek_kim_entry.valid [0]);
tran (tlv_word8[62], \tlv_word8.dek_kim_entry.label_index [2]);
tran (tlv_word8[61], \tlv_word8.dek_kim_entry.label_index [1]);
tran (tlv_word8[60], \tlv_word8.dek_kim_entry.label_index [0]);
tran (tlv_word8[59], \tlv_word8.dek_kim_entry.ckv_length [1]);
tran (tlv_word8[58], \tlv_word8.dek_kim_entry.ckv_length [0]);
tran (tlv_word8[57], \tlv_word8.dek_kim_entry.ckv_pointer [14]);
tran (tlv_word8[56], \tlv_word8.dek_kim_entry.ckv_pointer [13]);
tran (tlv_word8[55], \tlv_word8.dek_kim_entry.ckv_pointer [12]);
tran (tlv_word8[54], \tlv_word8.dek_kim_entry.ckv_pointer [11]);
tran (tlv_word8[53], \tlv_word8.dek_kim_entry.ckv_pointer [10]);
tran (tlv_word8[52], \tlv_word8.dek_kim_entry.ckv_pointer [9]);
tran (tlv_word8[51], \tlv_word8.dek_kim_entry.ckv_pointer [8]);
tran (tlv_word8[50], \tlv_word8.dek_kim_entry.ckv_pointer [7]);
tran (tlv_word8[49], \tlv_word8.dek_kim_entry.ckv_pointer [6]);
tran (tlv_word8[48], \tlv_word8.dek_kim_entry.ckv_pointer [5]);
tran (tlv_word8[47], \tlv_word8.dek_kim_entry.ckv_pointer [4]);
tran (tlv_word8[46], \tlv_word8.dek_kim_entry.ckv_pointer [3]);
tran (tlv_word8[45], \tlv_word8.dek_kim_entry.ckv_pointer [2]);
tran (tlv_word8[44], \tlv_word8.dek_kim_entry.ckv_pointer [1]);
tran (tlv_word8[43], \tlv_word8.dek_kim_entry.ckv_pointer [0]);
tran (tlv_word8[42], \tlv_word8.dek_kim_entry.pf_num [3]);
tran (tlv_word8[41], \tlv_word8.dek_kim_entry.pf_num [2]);
tran (tlv_word8[40], \tlv_word8.dek_kim_entry.pf_num [1]);
tran (tlv_word8[39], \tlv_word8.dek_kim_entry.pf_num [0]);
tran (tlv_word8[38], \tlv_word8.dek_kim_entry.vf_num [11]);
tran (tlv_word8[37], \tlv_word8.dek_kim_entry.vf_num [10]);
tran (tlv_word8[36], \tlv_word8.dek_kim_entry.vf_num [9]);
tran (tlv_word8[35], \tlv_word8.dek_kim_entry.vf_num [8]);
tran (tlv_word8[34], \tlv_word8.dek_kim_entry.vf_num [7]);
tran (tlv_word8[33], \tlv_word8.dek_kim_entry.vf_num [6]);
tran (tlv_word8[32], \tlv_word8.dek_kim_entry.vf_num [5]);
tran (tlv_word8[31], \tlv_word8.dek_kim_entry.vf_num [4]);
tran (tlv_word8[30], \tlv_word8.dek_kim_entry.vf_num [3]);
tran (tlv_word8[29], \tlv_word8.dek_kim_entry.vf_num [2]);
tran (tlv_word8[28], \tlv_word8.dek_kim_entry.vf_num [1]);
tran (tlv_word8[27], \tlv_word8.dek_kim_entry.vf_num [0]);
tran (tlv_word8[26], \tlv_word8.dek_kim_entry.vf_valid [0]);
tran (tlv_word9[25], \tlv_word9.unused [7]);
tran (tlv_word9[24], \tlv_word9.unused [6]);
tran (tlv_word9[23], \tlv_word9.unused [5]);
tran (tlv_word9[22], \tlv_word9.unused [4]);
tran (tlv_word9[21], \tlv_word9.unused [3]);
tran (tlv_word9[20], \tlv_word9.unused [2]);
tran (tlv_word9[16], \tlv_word9.vf_valid [0]);
tran (tlv_word9[15], \tlv_word9.pf_num [3]);
tran (tlv_word9[14], \tlv_word9.pf_num [2]);
tran (tlv_word9[13], \tlv_word9.pf_num [1]);
tran (tlv_word9[12], \tlv_word9.pf_num [0]);
tran (tlv_word9[11], \tlv_word9.vf_num [11]);
tran (tlv_word9[10], \tlv_word9.vf_num [10]);
tran (tlv_word9[9], \tlv_word9.vf_num [9]);
tran (tlv_word9[8], \tlv_word9.vf_num [8]);
tran (tlv_word9[7], \tlv_word9.vf_num [7]);
tran (tlv_word9[6], \tlv_word9.vf_num [6]);
tran (tlv_word9[5], \tlv_word9.vf_num [5]);
tran (tlv_word9[4], \tlv_word9.vf_num [4]);
tran (tlv_word9[3], \tlv_word9.vf_num [3]);
tran (tlv_word9[2], \tlv_word9.vf_num [2]);
tran (tlv_word9[1], \tlv_word9.vf_num [1]);
tran (tlv_word9[0], \tlv_word9.vf_num [0]);
tran (tlv_word9[63], \tlv_word9.dak_kim_entry.valid [0]);
tran (tlv_word9[62], \tlv_word9.dak_kim_entry.label_index [2]);
tran (tlv_word9[61], \tlv_word9.dak_kim_entry.label_index [1]);
tran (tlv_word9[60], \tlv_word9.dak_kim_entry.label_index [0]);
tran (tlv_word9[59], \tlv_word9.dak_kim_entry.ckv_length [1]);
tran (tlv_word9[58], \tlv_word9.dak_kim_entry.ckv_length [0]);
tran (tlv_word9[57], \tlv_word9.dak_kim_entry.ckv_pointer [14]);
tran (tlv_word9[56], \tlv_word9.dak_kim_entry.ckv_pointer [13]);
tran (tlv_word9[55], \tlv_word9.dak_kim_entry.ckv_pointer [12]);
tran (tlv_word9[54], \tlv_word9.dak_kim_entry.ckv_pointer [11]);
tran (tlv_word9[53], \tlv_word9.dak_kim_entry.ckv_pointer [10]);
tran (tlv_word9[52], \tlv_word9.dak_kim_entry.ckv_pointer [9]);
tran (tlv_word9[51], \tlv_word9.dak_kim_entry.ckv_pointer [8]);
tran (tlv_word9[50], \tlv_word9.dak_kim_entry.ckv_pointer [7]);
tran (tlv_word9[49], \tlv_word9.dak_kim_entry.ckv_pointer [6]);
tran (tlv_word9[48], \tlv_word9.dak_kim_entry.ckv_pointer [5]);
tran (tlv_word9[47], \tlv_word9.dak_kim_entry.ckv_pointer [4]);
tran (tlv_word9[46], \tlv_word9.dak_kim_entry.ckv_pointer [3]);
tran (tlv_word9[45], \tlv_word9.dak_kim_entry.ckv_pointer [2]);
tran (tlv_word9[44], \tlv_word9.dak_kim_entry.ckv_pointer [1]);
tran (tlv_word9[43], \tlv_word9.dak_kim_entry.ckv_pointer [0]);
tran (tlv_word9[42], \tlv_word9.dak_kim_entry.pf_num [3]);
tran (tlv_word9[41], \tlv_word9.dak_kim_entry.pf_num [2]);
tran (tlv_word9[40], \tlv_word9.dak_kim_entry.pf_num [1]);
tran (tlv_word9[39], \tlv_word9.dak_kim_entry.pf_num [0]);
tran (tlv_word9[38], \tlv_word9.dak_kim_entry.vf_num [11]);
tran (tlv_word9[37], \tlv_word9.dak_kim_entry.vf_num [10]);
tran (tlv_word9[36], \tlv_word9.dak_kim_entry.vf_num [9]);
tran (tlv_word9[35], \tlv_word9.dak_kim_entry.vf_num [8]);
tran (tlv_word9[34], \tlv_word9.dak_kim_entry.vf_num [7]);
tran (tlv_word9[33], \tlv_word9.dak_kim_entry.vf_num [6]);
tran (tlv_word9[32], \tlv_word9.dak_kim_entry.vf_num [5]);
tran (tlv_word9[31], \tlv_word9.dak_kim_entry.vf_num [4]);
tran (tlv_word9[30], \tlv_word9.dak_kim_entry.vf_num [3]);
tran (tlv_word9[29], \tlv_word9.dak_kim_entry.vf_num [2]);
tran (tlv_word9[28], \tlv_word9.dak_kim_entry.vf_num [1]);
tran (tlv_word9[27], \tlv_word9.dak_kim_entry.vf_num [0]);
tran (tlv_word9[26], \tlv_word9.dak_kim_entry.vf_valid [0]);
tran (tlv_word8[19], \tlv_word8.missing_iv [0]);
tran (tlv_word8[18], \tlv_word8.missing_guid [0]);
tran (tlv_word8[17], \tlv_word8.validate_dek [0]);
tran (dek_kim_entry_q[37], \dek_kim_entry_q.valid [0]);
tran (dek_kim_entry_q[36], \dek_kim_entry_q.label_index [2]);
tran (dek_kim_entry_q[35], \dek_kim_entry_q.label_index [1]);
tran (dek_kim_entry_q[34], \dek_kim_entry_q.label_index [0]);
tran (dek_kim_entry_q[33], \dek_kim_entry_q.ckv_length [1]);
tran (dek_kim_entry_q[32], \dek_kim_entry_q.ckv_length [0]);
tran (dek_kim_entry_q[31], \dek_kim_entry_q.ckv_pointer [14]);
tran (dek_kim_entry_q[30], \dek_kim_entry_q.ckv_pointer [13]);
tran (dek_kim_entry_q[29], \dek_kim_entry_q.ckv_pointer [12]);
tran (dek_kim_entry_q[28], \dek_kim_entry_q.ckv_pointer [11]);
tran (dek_kim_entry_q[27], \dek_kim_entry_q.ckv_pointer [10]);
tran (dek_kim_entry_q[26], \dek_kim_entry_q.ckv_pointer [9]);
tran (dek_kim_entry_q[25], \dek_kim_entry_q.ckv_pointer [8]);
tran (dek_kim_entry_q[24], \dek_kim_entry_q.ckv_pointer [7]);
tran (dek_kim_entry_q[23], \dek_kim_entry_q.ckv_pointer [6]);
tran (dek_kim_entry_q[22], \dek_kim_entry_q.ckv_pointer [5]);
tran (dek_kim_entry_q[21], \dek_kim_entry_q.ckv_pointer [4]);
tran (dek_kim_entry_q[20], \dek_kim_entry_q.ckv_pointer [3]);
tran (dek_kim_entry_q[19], \dek_kim_entry_q.ckv_pointer [2]);
tran (dek_kim_entry_q[18], \dek_kim_entry_q.ckv_pointer [1]);
tran (dek_kim_entry_q[17], \dek_kim_entry_q.ckv_pointer [0]);
tran (dek_kim_entry_q[16], \dek_kim_entry_q.pf_num [3]);
tran (dek_kim_entry_q[15], \dek_kim_entry_q.pf_num [2]);
tran (dek_kim_entry_q[14], \dek_kim_entry_q.pf_num [1]);
tran (dek_kim_entry_q[13], \dek_kim_entry_q.pf_num [0]);
tran (dek_kim_entry_q[12], \dek_kim_entry_q.vf_num [11]);
tran (dek_kim_entry_q[11], \dek_kim_entry_q.vf_num [10]);
tran (dek_kim_entry_q[10], \dek_kim_entry_q.vf_num [9]);
tran (dek_kim_entry_q[9], \dek_kim_entry_q.vf_num [8]);
tran (dek_kim_entry_q[8], \dek_kim_entry_q.vf_num [7]);
tran (dek_kim_entry_q[7], \dek_kim_entry_q.vf_num [6]);
tran (dek_kim_entry_q[6], \dek_kim_entry_q.vf_num [5]);
tran (dek_kim_entry_q[5], \dek_kim_entry_q.vf_num [4]);
tran (dek_kim_entry_q[4], \dek_kim_entry_q.vf_num [3]);
tran (dek_kim_entry_q[3], \dek_kim_entry_q.vf_num [2]);
tran (dek_kim_entry_q[2], \dek_kim_entry_q.vf_num [1]);
tran (dek_kim_entry_q[1], \dek_kim_entry_q.vf_num [0]);
tran (dek_kim_entry_q[0], \dek_kim_entry_q.vf_valid [0]);
tran (dak_kim_entry_q[37], \dak_kim_entry_q.valid [0]);
tran (dak_kim_entry_q[36], \dak_kim_entry_q.label_index [2]);
tran (dak_kim_entry_q[35], \dak_kim_entry_q.label_index [1]);
tran (dak_kim_entry_q[34], \dak_kim_entry_q.label_index [0]);
tran (dak_kim_entry_q[33], \dak_kim_entry_q.ckv_length [1]);
tran (dak_kim_entry_q[32], \dak_kim_entry_q.ckv_length [0]);
tran (dak_kim_entry_q[31], \dak_kim_entry_q.ckv_pointer [14]);
tran (dak_kim_entry_q[30], \dak_kim_entry_q.ckv_pointer [13]);
tran (dak_kim_entry_q[29], \dak_kim_entry_q.ckv_pointer [12]);
tran (dak_kim_entry_q[28], \dak_kim_entry_q.ckv_pointer [11]);
tran (dak_kim_entry_q[27], \dak_kim_entry_q.ckv_pointer [10]);
tran (dak_kim_entry_q[26], \dak_kim_entry_q.ckv_pointer [9]);
tran (dak_kim_entry_q[25], \dak_kim_entry_q.ckv_pointer [8]);
tran (dak_kim_entry_q[24], \dak_kim_entry_q.ckv_pointer [7]);
tran (dak_kim_entry_q[23], \dak_kim_entry_q.ckv_pointer [6]);
tran (dak_kim_entry_q[22], \dak_kim_entry_q.ckv_pointer [5]);
tran (dak_kim_entry_q[21], \dak_kim_entry_q.ckv_pointer [4]);
tran (dak_kim_entry_q[20], \dak_kim_entry_q.ckv_pointer [3]);
tran (dak_kim_entry_q[19], \dak_kim_entry_q.ckv_pointer [2]);
tran (dak_kim_entry_q[18], \dak_kim_entry_q.ckv_pointer [1]);
tran (dak_kim_entry_q[17], \dak_kim_entry_q.ckv_pointer [0]);
tran (dak_kim_entry_q[16], \dak_kim_entry_q.pf_num [3]);
tran (dak_kim_entry_q[15], \dak_kim_entry_q.pf_num [2]);
tran (dak_kim_entry_q[14], \dak_kim_entry_q.pf_num [1]);
tran (dak_kim_entry_q[13], \dak_kim_entry_q.pf_num [0]);
tran (dak_kim_entry_q[12], \dak_kim_entry_q.vf_num [11]);
tran (dak_kim_entry_q[11], \dak_kim_entry_q.vf_num [10]);
tran (dak_kim_entry_q[10], \dak_kim_entry_q.vf_num [9]);
tran (dak_kim_entry_q[9], \dak_kim_entry_q.vf_num [8]);
tran (dak_kim_entry_q[8], \dak_kim_entry_q.vf_num [7]);
tran (dak_kim_entry_q[7], \dak_kim_entry_q.vf_num [6]);
tran (dak_kim_entry_q[6], \dak_kim_entry_q.vf_num [5]);
tran (dak_kim_entry_q[5], \dak_kim_entry_q.vf_num [4]);
tran (dak_kim_entry_q[4], \dak_kim_entry_q.vf_num [3]);
tran (dak_kim_entry_q[3], \dak_kim_entry_q.vf_num [2]);
tran (dak_kim_entry_q[2], \dak_kim_entry_q.vf_num [1]);
tran (dak_kim_entry_q[1], \dak_kim_entry_q.vf_num [0]);
tran (dak_kim_entry_q[0], \dak_kim_entry_q.vf_valid [0]);
Q_BUF U0 ( .A(_zy_sva_disable_unenc_keys_3_reset_or), .Z(_zy_sva_enable_unenc_keys_2_reset_or));
Q_BUF U1 ( .A(_zy_sva_enable_unenc_keys_4_reset_or), .Z(_zy_sva_disable_unenc_keys_3_reset_or));
Q_BUF U2 ( .A(_zy_sva_disable_unenc_keys_5_reset_or), .Z(_zy_sva_enable_unenc_keys_4_reset_or));
Q_BUF U3 ( .A(_zy_sva_enable_unenc_keys_6_reset_or), .Z(_zy_sva_disable_unenc_keys_5_reset_or));
Q_BUF U4 ( .A(_zy_sva_disable_unenc_keys_7_reset_or), .Z(_zy_sva_enable_unenc_keys_6_reset_or));
Q_BUF U5 ( .A(_zy_sva_enable_unenc_keys_8_reset_or), .Z(_zy_sva_disable_unenc_keys_7_reset_or));
Q_BUF U6 ( .A(_zy_sva_disable_unenc_keys_9_reset_or), .Z(_zy_sva_enable_unenc_keys_8_reset_or));
Q_BUF U7 ( .A(_zy_sva_enable_unenc_keys_10_reset_or), .Z(_zy_sva_disable_unenc_keys_9_reset_or));
Q_BUF U8 ( .A(_zy_sva_disable_unenc_keys_1_reset_or), .Z(_zy_sva_enable_unenc_keys_10_reset_or));
Q_ASSIGN U9 ( .B(parser_kimreader_data[0]), .A(tlv_word0[0]));
Q_ASSIGN U10 ( .B(parser_kimreader_data[0]), .A(aux_key_ctrl[0]));
Q_ASSIGN U11 ( .B(parser_kimreader_data[1]), .A(tlv_word0[1]));
Q_ASSIGN U12 ( .B(parser_kimreader_data[1]), .A(aux_key_ctrl[1]));
Q_ASSIGN U13 ( .B(parser_kimreader_data[2]), .A(tlv_word0[2]));
Q_ASSIGN U14 ( .B(parser_kimreader_data[2]), .A(aux_key_ctrl[2]));
Q_ASSIGN U15 ( .B(parser_kimreader_data[3]), .A(tlv_word0[3]));
Q_ASSIGN U16 ( .B(parser_kimreader_data[3]), .A(aux_key_ctrl[3]));
Q_ASSIGN U17 ( .B(parser_kimreader_data[4]), .A(tlv_word0[4]));
Q_ASSIGN U18 ( .B(parser_kimreader_data[4]), .A(aux_key_ctrl[4]));
Q_ASSIGN U19 ( .B(parser_kimreader_data[5]), .A(tlv_word0[5]));
Q_ASSIGN U20 ( .B(parser_kimreader_data[5]), .A(aux_key_ctrl[5]));
Q_ASSIGN U21 ( .B(parser_kimreader_data[6]), .A(tlv_word0[6]));
Q_ASSIGN U22 ( .B(parser_kimreader_data[6]), .A(aux_key_ctrl[6]));
Q_ASSIGN U23 ( .B(parser_kimreader_data[7]), .A(tlv_word0[7]));
Q_ASSIGN U24 ( .B(parser_kimreader_data[7]), .A(aux_key_ctrl[7]));
Q_ASSIGN U25 ( .B(parser_kimreader_data[8]), .A(tlv_word0[8]));
Q_ASSIGN U26 ( .B(parser_kimreader_data[8]), .A(tlv_word42[8]));
Q_ASSIGN U27 ( .B(parser_kimreader_data[8]), .A(aux_key_ctrl[8]));
Q_ASSIGN U28 ( .B(parser_kimreader_data[9]), .A(tlv_word0[9]));
Q_ASSIGN U29 ( .B(parser_kimreader_data[9]), .A(tlv_word42[9]));
Q_ASSIGN U30 ( .B(parser_kimreader_data[9]), .A(aux_key_ctrl[9]));
Q_ASSIGN U31 ( .B(parser_kimreader_data[10]), .A(tlv_word0[10]));
Q_ASSIGN U32 ( .B(parser_kimreader_data[10]), .A(tlv_word42[10]));
Q_ASSIGN U33 ( .B(parser_kimreader_data[10]), .A(aux_key_ctrl[10]));
Q_ASSIGN U34 ( .B(parser_kimreader_data[11]), .A(tlv_word0[11]));
Q_ASSIGN U35 ( .B(parser_kimreader_data[11]), .A(tlv_word42[11]));
Q_ASSIGN U36 ( .B(parser_kimreader_data[11]), .A(aux_key_ctrl[11]));
Q_ASSIGN U37 ( .B(parser_kimreader_data[12]), .A(tlv_word0[12]));
Q_ASSIGN U38 ( .B(parser_kimreader_data[12]), .A(tlv_word42[12]));
Q_ASSIGN U39 ( .B(parser_kimreader_data[12]), .A(aux_key_ctrl[12]));
Q_ASSIGN U40 ( .B(parser_kimreader_data[13]), .A(tlv_word0[13]));
Q_ASSIGN U41 ( .B(parser_kimreader_data[13]), .A(tlv_word42[13]));
Q_ASSIGN U42 ( .B(parser_kimreader_data[13]), .A(aux_key_ctrl[13]));
Q_ASSIGN U43 ( .B(parser_kimreader_data[14]), .A(tlv_word0[14]));
Q_ASSIGN U44 ( .B(parser_kimreader_data[14]), .A(tlv_word42[14]));
Q_ASSIGN U45 ( .B(parser_kimreader_data[14]), .A(aux_key_ctrl[14]));
Q_ASSIGN U46 ( .B(parser_kimreader_data[15]), .A(tlv_word0[15]));
Q_ASSIGN U47 ( .B(parser_kimreader_data[15]), .A(tlv_word42[15]));
Q_ASSIGN U48 ( .B(parser_kimreader_data[15]), .A(aux_key_ctrl[15]));
Q_ASSIGN U49 ( .B(parser_kimreader_data[16]), .A(tlv_word0[16]));
Q_ASSIGN U50 ( .B(parser_kimreader_data[16]), .A(tlv_word42[16]));
Q_ASSIGN U51 ( .B(parser_kimreader_data[16]), .A(aux_key_ctrl[16]));
Q_ASSIGN U52 ( .B(parser_kimreader_data[17]), .A(tlv_word0[17]));
Q_ASSIGN U53 ( .B(parser_kimreader_data[17]), .A(tlv_word42[17]));
Q_ASSIGN U54 ( .B(parser_kimreader_data[17]), .A(aux_key_ctrl[17]));
Q_ASSIGN U55 ( .B(parser_kimreader_data[18]), .A(tlv_word0[18]));
Q_ASSIGN U56 ( .B(parser_kimreader_data[18]), .A(tlv_word42[18]));
Q_ASSIGN U57 ( .B(parser_kimreader_data[18]), .A(aux_key_ctrl[18]));
Q_ASSIGN U58 ( .B(parser_kimreader_data[19]), .A(tlv_word0[19]));
Q_ASSIGN U59 ( .B(parser_kimreader_data[19]), .A(tlv_word42[19]));
Q_ASSIGN U60 ( .B(parser_kimreader_data[19]), .A(aux_key_ctrl[19]));
Q_ASSIGN U61 ( .B(parser_kimreader_data[20]), .A(tlv_word0[20]));
Q_ASSIGN U62 ( .B(parser_kimreader_data[20]), .A(tlv_word42[20]));
Q_ASSIGN U63 ( .B(parser_kimreader_data[20]), .A(aux_key_ctrl[20]));
Q_ASSIGN U64 ( .B(parser_kimreader_data[21]), .A(tlv_word0[21]));
Q_ASSIGN U65 ( .B(parser_kimreader_data[21]), .A(tlv_word42[21]));
Q_ASSIGN U66 ( .B(parser_kimreader_data[21]), .A(aux_key_ctrl[21]));
Q_ASSIGN U67 ( .B(parser_kimreader_data[22]), .A(tlv_word0[22]));
Q_ASSIGN U68 ( .B(parser_kimreader_data[22]), .A(tlv_word42[22]));
Q_ASSIGN U69 ( .B(parser_kimreader_data[22]), .A(aux_key_ctrl[22]));
Q_ASSIGN U70 ( .B(parser_kimreader_data[23]), .A(tlv_word0[23]));
Q_ASSIGN U71 ( .B(parser_kimreader_data[23]), .A(tlv_word42[23]));
Q_ASSIGN U72 ( .B(parser_kimreader_data[23]), .A(aux_key_ctrl[23]));
Q_ASSIGN U73 ( .B(parser_kimreader_data[24]), .A(tlv_word0[24]));
Q_ASSIGN U74 ( .B(parser_kimreader_data[24]), .A(tlv_word42[24]));
Q_ASSIGN U75 ( .B(parser_kimreader_data[24]), .A(aux_key_ctrl[24]));
Q_ASSIGN U76 ( .B(parser_kimreader_data[25]), .A(tlv_word0[25]));
Q_ASSIGN U77 ( .B(parser_kimreader_data[25]), .A(tlv_word42[25]));
Q_ASSIGN U78 ( .B(parser_kimreader_data[25]), .A(aux_key_ctrl[25]));
Q_ASSIGN U79 ( .B(parser_kimreader_data[26]), .A(tlv_word0[26]));
Q_ASSIGN U80 ( .B(parser_kimreader_data[26]), .A(tlv_word42[26]));
Q_ASSIGN U81 ( .B(parser_kimreader_data[26]), .A(aux_key_ctrl[26]));
Q_ASSIGN U82 ( .B(parser_kimreader_data[27]), .A(tlv_word0[27]));
Q_ASSIGN U83 ( .B(parser_kimreader_data[27]), .A(tlv_word42[27]));
Q_ASSIGN U84 ( .B(parser_kimreader_data[27]), .A(aux_key_ctrl[27]));
Q_ASSIGN U85 ( .B(parser_kimreader_data[28]), .A(tlv_word0[28]));
Q_ASSIGN U86 ( .B(parser_kimreader_data[28]), .A(tlv_word42[28]));
Q_ASSIGN U87 ( .B(parser_kimreader_data[28]), .A(aux_key_ctrl[28]));
Q_ASSIGN U88 ( .B(parser_kimreader_data[29]), .A(tlv_word0[29]));
Q_ASSIGN U89 ( .B(parser_kimreader_data[29]), .A(tlv_word42[29]));
Q_ASSIGN U90 ( .B(parser_kimreader_data[29]), .A(aux_key_ctrl[29]));
Q_ASSIGN U91 ( .B(parser_kimreader_data[30]), .A(tlv_word0[30]));
Q_ASSIGN U92 ( .B(parser_kimreader_data[30]), .A(tlv_word42[30]));
Q_ASSIGN U93 ( .B(parser_kimreader_data[30]), .A(aux_key_ctrl[30]));
Q_ASSIGN U94 ( .B(parser_kimreader_data[31]), .A(tlv_word0[31]));
Q_ASSIGN U95 ( .B(parser_kimreader_data[31]), .A(tlv_word42[31]));
Q_ASSIGN U96 ( .B(parser_kimreader_data[31]), .A(aux_key_ctrl[31]));
Q_BUF U97 ( .A(kim_errors_q[0]), .Z(tlv_word42[0]));
Q_BUF U98 ( .A(kim_errors_q[1]), .Z(tlv_word42[1]));
Q_BUF U99 ( .A(kim_errors_q[2]), .Z(tlv_word42[2]));
Q_BUF U100 ( .A(kim_errors_q[3]), .Z(tlv_word42[3]));
Q_BUF U101 ( .A(kim_errors_q[4]), .Z(tlv_word42[4]));
Q_BUF U102 ( .A(kim_errors_q[5]), .Z(tlv_word42[5]));
Q_BUF U103 ( .A(kim_errors_q[6]), .Z(tlv_word42[6]));
Q_BUF U104 ( .A(kim_errors_q[7]), .Z(tlv_word42[7]));
Q_ASSIGN U105 ( .B(parser_kimreader_data[32]), .A(tlv_word0[32]));
Q_ASSIGN U106 ( .B(parser_kimreader_data[32]), .A(tlv_word42[32]));
Q_ASSIGN U107 ( .B(parser_kimreader_data[33]), .A(tlv_word0[33]));
Q_ASSIGN U108 ( .B(parser_kimreader_data[33]), .A(tlv_word42[33]));
Q_ASSIGN U109 ( .B(parser_kimreader_data[34]), .A(tlv_word0[34]));
Q_ASSIGN U110 ( .B(parser_kimreader_data[34]), .A(tlv_word42[34]));
Q_ASSIGN U111 ( .B(parser_kimreader_data[35]), .A(tlv_word0[35]));
Q_ASSIGN U112 ( .B(parser_kimreader_data[35]), .A(tlv_word42[35]));
Q_ASSIGN U113 ( .B(parser_kimreader_data[36]), .A(tlv_word0[36]));
Q_ASSIGN U114 ( .B(parser_kimreader_data[36]), .A(tlv_word42[36]));
Q_ASSIGN U115 ( .B(parser_kimreader_data[37]), .A(tlv_word0[37]));
Q_ASSIGN U116 ( .B(parser_kimreader_data[37]), .A(tlv_word42[37]));
Q_ASSIGN U117 ( .B(parser_kimreader_data[38]), .A(tlv_word0[38]));
Q_ASSIGN U118 ( .B(parser_kimreader_data[38]), .A(tlv_word42[38]));
Q_ASSIGN U119 ( .B(parser_kimreader_data[39]), .A(tlv_word0[39]));
Q_ASSIGN U120 ( .B(parser_kimreader_data[39]), .A(tlv_word42[39]));
Q_ASSIGN U121 ( .B(parser_kimreader_data[40]), .A(tlv_word0[40]));
Q_ASSIGN U122 ( .B(parser_kimreader_data[40]), .A(tlv_word42[40]));
Q_ASSIGN U123 ( .B(parser_kimreader_data[41]), .A(tlv_word0[41]));
Q_ASSIGN U124 ( .B(parser_kimreader_data[41]), .A(tlv_word42[41]));
Q_ASSIGN U125 ( .B(parser_kimreader_data[42]), .A(tlv_word0[42]));
Q_ASSIGN U126 ( .B(parser_kimreader_data[42]), .A(tlv_word42[42]));
Q_ASSIGN U127 ( .B(parser_kimreader_data[43]), .A(tlv_word0[43]));
Q_ASSIGN U128 ( .B(parser_kimreader_data[43]), .A(tlv_word42[43]));
Q_ASSIGN U129 ( .B(parser_kimreader_data[44]), .A(tlv_word0[44]));
Q_ASSIGN U130 ( .B(parser_kimreader_data[44]), .A(tlv_word42[44]));
Q_ASSIGN U131 ( .B(parser_kimreader_data[45]), .A(tlv_word0[45]));
Q_ASSIGN U132 ( .B(parser_kimreader_data[45]), .A(tlv_word42[45]));
Q_ASSIGN U133 ( .B(parser_kimreader_data[46]), .A(tlv_word0[46]));
Q_ASSIGN U134 ( .B(parser_kimreader_data[46]), .A(tlv_word42[46]));
Q_ASSIGN U135 ( .B(parser_kimreader_data[47]), .A(tlv_word0[47]));
Q_ASSIGN U136 ( .B(parser_kimreader_data[47]), .A(tlv_word42[47]));
Q_ASSIGN U137 ( .B(parser_kimreader_data[48]), .A(tlv_word0[48]));
Q_ASSIGN U138 ( .B(parser_kimreader_data[48]), .A(tlv_word42[48]));
Q_ASSIGN U139 ( .B(parser_kimreader_data[49]), .A(tlv_word0[49]));
Q_ASSIGN U140 ( .B(parser_kimreader_data[49]), .A(tlv_word42[49]));
Q_ASSIGN U141 ( .B(parser_kimreader_data[50]), .A(tlv_word0[50]));
Q_ASSIGN U142 ( .B(parser_kimreader_data[50]), .A(tlv_word42[50]));
Q_ASSIGN U143 ( .B(parser_kimreader_data[51]), .A(tlv_word0[51]));
Q_ASSIGN U144 ( .B(parser_kimreader_data[51]), .A(tlv_word42[51]));
Q_ASSIGN U145 ( .B(parser_kimreader_data[52]), .A(tlv_word0[52]));
Q_ASSIGN U146 ( .B(parser_kimreader_data[52]), .A(tlv_word42[52]));
Q_ASSIGN U147 ( .B(parser_kimreader_data[53]), .A(tlv_word0[53]));
Q_ASSIGN U148 ( .B(parser_kimreader_data[53]), .A(tlv_word42[53]));
Q_ASSIGN U149 ( .B(parser_kimreader_data[54]), .A(tlv_word0[54]));
Q_ASSIGN U150 ( .B(parser_kimreader_data[54]), .A(tlv_word42[54]));
Q_ASSIGN U151 ( .B(parser_kimreader_data[55]), .A(tlv_word0[55]));
Q_ASSIGN U152 ( .B(parser_kimreader_data[55]), .A(tlv_word42[55]));
Q_BUF U153 ( .A(tlv_word8[17]), .Z(tlv_word9[17]));
Q_BUF U154 ( .A(tlv_word8[18]), .Z(tlv_word9[18]));
Q_BUF U155 ( .A(tlv_word8[19]), .Z(tlv_word9[19]));
Q_BUF U156 ( .A(tlv_word9[0]), .Z(tlv_word8[0]));
Q_BUF U157 ( .A(tlv_word9[1]), .Z(tlv_word8[1]));
Q_BUF U158 ( .A(tlv_word9[2]), .Z(tlv_word8[2]));
Q_BUF U159 ( .A(tlv_word9[3]), .Z(tlv_word8[3]));
Q_BUF U160 ( .A(tlv_word9[4]), .Z(tlv_word8[4]));
Q_BUF U161 ( .A(tlv_word9[5]), .Z(tlv_word8[5]));
Q_BUF U162 ( .A(tlv_word9[6]), .Z(tlv_word8[6]));
Q_BUF U163 ( .A(tlv_word9[7]), .Z(tlv_word8[7]));
Q_BUF U164 ( .A(tlv_word9[8]), .Z(tlv_word8[8]));
Q_BUF U165 ( .A(tlv_word9[9]), .Z(tlv_word8[9]));
Q_BUF U166 ( .A(tlv_word9[10]), .Z(tlv_word8[10]));
Q_BUF U167 ( .A(tlv_word9[11]), .Z(tlv_word8[11]));
Q_BUF U168 ( .A(tlv_word9[12]), .Z(tlv_word8[12]));
Q_BUF U169 ( .A(tlv_word9[13]), .Z(tlv_word8[13]));
Q_BUF U170 ( .A(tlv_word9[14]), .Z(tlv_word8[14]));
Q_BUF U171 ( .A(tlv_word9[15]), .Z(tlv_word8[15]));
Q_BUF U172 ( .A(tlv_word9[16]), .Z(tlv_word8[16]));
Q_BUF U173 ( .A(tlv_word9[20]), .Z(tlv_word8[20]));
Q_BUF U174 ( .A(tlv_word9[21]), .Z(tlv_word8[21]));
Q_BUF U175 ( .A(tlv_word9[22]), .Z(tlv_word8[22]));
Q_BUF U176 ( .A(tlv_word9[23]), .Z(tlv_word8[23]));
Q_BUF U177 ( .A(tlv_word9[24]), .Z(tlv_word8[24]));
Q_BUF U178 ( .A(tlv_word9[25]), .Z(tlv_word8[25]));
Q_ASSIGN U179 ( .B(parser_kimreader_data[56]), .A(tlv_word0[56]));
Q_ASSIGN U180 ( .B(parser_kimreader_data[57]), .A(tlv_word0[57]));
Q_ASSIGN U181 ( .B(parser_kimreader_data[58]), .A(tlv_word0[58]));
Q_ASSIGN U182 ( .B(parser_kimreader_data[59]), .A(tlv_word0[59]));
Q_ASSIGN U183 ( .B(parser_kimreader_data[60]), .A(tlv_word0[60]));
Q_ASSIGN U184 ( .B(parser_kimreader_data[61]), .A(tlv_word0[61]));
Q_ASSIGN U185 ( .B(parser_kimreader_data[62]), .A(tlv_word0[62]));
Q_ASSIGN U186 ( .B(parser_kimreader_data[63]), .A(tlv_word0[63]));
Q_OR02 U187 ( .A0(n373), .A1(n374), .Z(n1));
wire [2:0] n651 = 3'b000;
Q_ASSERT \key_type_enc_dek_6_.enable_unenc_keys  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_enable_unenc_keys_10_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_enable_unenc_keys_10_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n651[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_6_.enable_unenc_keys " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_6_.enable_unenc_keys " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kim_drng_reader.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_6_.enable_unenc_keys " ASSERT_LINE 596
wire [2:0] n652 = 3'b000;
Q_ASSERT \key_type_enc_dek_6_.disable_unenc_keys  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_disable_unenc_keys_9_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_disable_unenc_keys_9_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n652[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_6_.disable_unenc_keys " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_6_.disable_unenc_keys " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kim_drng_reader.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_6_.disable_unenc_keys " ASSERT_LINE 591
wire [2:0] n653 = 3'b000;
Q_ASSERT \key_type_enc_dek_5_.enable_unenc_keys  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_enable_unenc_keys_8_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_enable_unenc_keys_8_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n653[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_5_.enable_unenc_keys " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_5_.enable_unenc_keys " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kim_drng_reader.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_5_.enable_unenc_keys " ASSERT_LINE 596
wire [2:0] n654 = 3'b000;
Q_ASSERT \key_type_enc_dek_5_.disable_unenc_keys  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_disable_unenc_keys_7_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_disable_unenc_keys_7_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n654[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_5_.disable_unenc_keys " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_5_.disable_unenc_keys " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kim_drng_reader.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_5_.disable_unenc_keys " ASSERT_LINE 591
wire [2:0] n655 = 3'b000;
Q_ASSERT \key_type_enc_dek_4_.enable_unenc_keys  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_enable_unenc_keys_6_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_enable_unenc_keys_6_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n655[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_4_.enable_unenc_keys " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_4_.enable_unenc_keys " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kim_drng_reader.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_4_.enable_unenc_keys " ASSERT_LINE 596
wire [2:0] n656 = 3'b000;
Q_ASSERT \key_type_enc_dek_4_.disable_unenc_keys  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_disable_unenc_keys_5_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_disable_unenc_keys_5_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n656[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_4_.disable_unenc_keys " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_4_.disable_unenc_keys " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kim_drng_reader.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_4_.disable_unenc_keys " ASSERT_LINE 591
wire [2:0] n657 = 3'b000;
Q_ASSERT \key_type_enc_dek_3_.enable_unenc_keys  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_enable_unenc_keys_4_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_enable_unenc_keys_4_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n657[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_3_.enable_unenc_keys " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_3_.enable_unenc_keys " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kim_drng_reader.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_3_.enable_unenc_keys " ASSERT_LINE 596
wire [2:0] n658 = 3'b000;
Q_ASSERT \key_type_enc_dek_3_.disable_unenc_keys  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_disable_unenc_keys_3_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_disable_unenc_keys_3_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n658[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_3_.disable_unenc_keys " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_3_.disable_unenc_keys " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kim_drng_reader.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_3_.disable_unenc_keys " ASSERT_LINE 591
wire [2:0] n659 = 3'b000;
Q_ASSERT \key_type_enc_dek_2_.enable_unenc_keys  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_enable_unenc_keys_2_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_enable_unenc_keys_2_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n659[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_2_.enable_unenc_keys " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_2_.enable_unenc_keys " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kim_drng_reader.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_2_.enable_unenc_keys " ASSERT_LINE 596
wire [2:0] n660 = 3'b000;
Q_ASSERT \key_type_enc_dek_2_.disable_unenc_keys  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_disable_unenc_keys_1_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_disable_unenc_keys_1_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n660[0]));
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_2_.disable_unenc_keys " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\key_type_enc_dek_2_.disable_unenc_keys " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kim_drng_reader.v"
//pragma CVAINTPROP INSTANCE "\key_type_enc_dek_2_.disable_unenc_keys " ASSERT_LINE 591
ixc_sample_logic_1_3 _zz_zy_sva_b9 ( _zy_sva_b9, _zy_sva_b9_t);
ixc_sample_logic_1_3 _zz_zy_sva_b8 ( _zy_sva_b8, _zy_sva_b8_t);
ixc_sample_logic_1_3 _zz_zy_sva_b7 ( _zy_sva_b7, _zy_sva_b7_t);
ixc_sample_logic_1_3 _zz_zy_sva_b6 ( _zy_sva_b6, _zy_sva_b6_t);
ixc_sample_logic_1_3 _zz_zy_sva_b5 ( _zy_sva_b5, _zy_sva_b5_t);
ixc_sample_logic_1_3 _zz_zy_sva_b4 ( _zy_sva_b4, _zy_sva_b4_t);
ixc_sample_logic_1_3 _zz_zy_sva_b3 ( _zy_sva_b3, _zy_sva_b3_t);
ixc_sample_logic_1_3 _zz_zy_sva_b2 ( _zy_sva_b2, _zy_sva_b2_t);
ixc_sample_logic_1_3 _zz_zy_sva_b1 ( _zy_sva_b1, _zy_sva_b1_t);
ixc_sample_logic_1_3 _zz_zy_sva_b0 ( _zy_sva_b0, _zy_sva_b0_t);
Q_NR03 U208 ( .A0(n3), .A1(disable_unencrypted_keys), .A2(n22), .Z(_zy_sva_b9_t));
Q_AN03 U209 ( .A0(n4), .A1(disable_unencrypted_keys), .A2(n23), .Z(_zy_sva_b8_t));
Q_INV U210 ( .A(n22), .Z(n23));
Q_OR02 U211 ( .A0(n6), .A1(n21), .Z(n22));
Q_OR03 U212 ( .A0(n14), .A1(n5), .A2(parser_kimreader_data[39]), .Z(n21));
Q_NR03 U213 ( .A0(n3), .A1(disable_unencrypted_keys), .A2(n19), .Z(_zy_sva_b7_t));
Q_AN03 U214 ( .A0(n4), .A1(disable_unencrypted_keys), .A2(n20), .Z(_zy_sva_b6_t));
Q_INV U215 ( .A(n19), .Z(n20));
Q_OR02 U216 ( .A0(n6), .A1(n18), .Z(n19));
Q_OR03 U217 ( .A0(n14), .A1(parser_kimreader_data[40]), .A2(n10), .Z(n18));
Q_NR03 U218 ( .A0(n3), .A1(disable_unencrypted_keys), .A2(n16), .Z(_zy_sva_b5_t));
Q_AN03 U219 ( .A0(n4), .A1(disable_unencrypted_keys), .A2(n17), .Z(_zy_sva_b4_t));
Q_INV U220 ( .A(n16), .Z(n17));
Q_OR02 U221 ( .A0(n6), .A1(n15), .Z(n16));
Q_OR03 U222 ( .A0(n14), .A1(parser_kimreader_data[40]), .A2(parser_kimreader_data[39]), .Z(n15));
Q_INV U223 ( .A(parser_kimreader_data[41]), .Z(n14));
Q_NR03 U224 ( .A0(n3), .A1(disable_unencrypted_keys), .A2(n12), .Z(_zy_sva_b3_t));
Q_AN03 U225 ( .A0(n4), .A1(disable_unencrypted_keys), .A2(n13), .Z(_zy_sva_b2_t));
Q_INV U226 ( .A(n12), .Z(n13));
Q_OR02 U227 ( .A0(n6), .A1(n11), .Z(n12));
Q_OR03 U228 ( .A0(parser_kimreader_data[41]), .A1(n5), .A2(n10), .Z(n11));
Q_INV U229 ( .A(parser_kimreader_data[39]), .Z(n10));
Q_NR03 U230 ( .A0(n3), .A1(disable_unencrypted_keys), .A2(n8), .Z(_zy_sva_b1_t));
Q_AN03 U231 ( .A0(n4), .A1(disable_unencrypted_keys), .A2(n9), .Z(_zy_sva_b0_t));
Q_INV U232 ( .A(n8), .Z(n9));
Q_OR02 U233 ( .A0(n6), .A1(n7), .Z(n8));
Q_OR03 U234 ( .A0(parser_kimreader_data[41]), .A1(n5), .A2(parser_kimreader_data[39]), .Z(n7));
Q_OR03 U235 ( .A0(parser_kimreader_data[44]), .A1(parser_kimreader_data[43]), .A2(parser_kimreader_data[42]), .Z(n6));
Q_INV U236 ( .A(parser_kimreader_data[40]), .Z(n5));
Q_INV U237 ( .A(n3), .Z(n4));
Q_OR02 U238 ( .A0(parser_kimreader_data[64]), .A1(n2), .Z(n3));
Q_OR03 U239 ( .A0(parser_kimreader_data[67]), .A1(parser_kimreader_data[66]), .A2(parser_kimreader_data[65]), .Z(n2));
Q_INV U240 ( .A(rst_n), .Z(_zy_sva_disable_unenc_keys_1_reset_or));
ixc_assign _zz_strnp_21 ( _zy_simnet_stat_aux_cmd_with_vf_pf_fail_21_w$, 
	stat_aux_cmd_with_vf_pf_fail);
ixc_assign _zz_strnp_20 ( _zy_simnet_stat_aux_key_type_13_20_w$, 
	stat_aux_key_type_13);
ixc_assign _zz_strnp_19 ( _zy_simnet_stat_aux_key_type_12_19_w$, 
	stat_aux_key_type_12);
ixc_assign _zz_strnp_18 ( _zy_simnet_stat_aux_key_type_11_18_w$, 
	stat_aux_key_type_11);
ixc_assign _zz_strnp_17 ( _zy_simnet_stat_aux_key_type_10_17_w$, 
	stat_aux_key_type_10);
ixc_assign _zz_strnp_16 ( _zy_simnet_stat_aux_key_type_9_16_w$, 
	stat_aux_key_type_9);
ixc_assign _zz_strnp_15 ( _zy_simnet_stat_aux_key_type_8_15_w$, 
	stat_aux_key_type_8);
ixc_assign _zz_strnp_14 ( _zy_simnet_stat_aux_key_type_7_14_w$, 
	stat_aux_key_type_7);
ixc_assign _zz_strnp_13 ( _zy_simnet_stat_aux_key_type_6_13_w$, 
	stat_aux_key_type_6);
ixc_assign _zz_strnp_12 ( _zy_simnet_stat_aux_key_type_5_12_w$, 
	stat_aux_key_type_5);
ixc_assign _zz_strnp_11 ( _zy_simnet_stat_aux_key_type_4_11_w$, 
	stat_aux_key_type_4);
ixc_assign _zz_strnp_10 ( _zy_simnet_stat_aux_key_type_3_10_w$, 
	stat_aux_key_type_3);
ixc_assign _zz_strnp_9 ( _zy_simnet_stat_aux_key_type_2_9_w$, 
	stat_aux_key_type_2);
ixc_assign _zz_strnp_8 ( _zy_simnet_stat_aux_key_type_1_8_w$, 
	stat_aux_key_type_1);
ixc_assign _zz_strnp_7 ( _zy_simnet_stat_aux_key_type_0_7_w$, 
	stat_aux_key_type_0);
ixc_assign _zz_strnp_6 ( _zy_simnet_stat_req_with_expired_seed_6_w$, 
	stat_req_with_expired_seed);
ixc_assign_14 _zz_strnp_5 ( _zy_simnet_kim_addr_5_w$[0:13], kim_addr[13:0]);
ixc_assign _zz_strnp_4 ( _zy_simnet_kim_rd_4_w$, kim_rd);
ixc_assign _zz_strnp_3 ( _zy_simnet_drng_ack_3_w$, drng_ack);
ixc_assign_71 _zz_strnp_2 ( _zy_simnet_kimreader_ckvreader_data_2_w$[0:70], 
	kimreader_ckvreader_data[70:0]);
ixc_assign _zz_strnp_1 ( _zy_simnet_kimreader_ckvreader_valid_1_w$, 
	kimreader_ckvreader_valid);
ixc_assign _zz_strnp_0 ( _zy_simnet_kimreader_parser_ack_0_w$, 
	kimreader_parser_ack);
Q_AN02 U263 ( .A0(rst_n), .A1(_zy_sva_b0), .Z(n24));
Q_AN02 U264 ( .A0(rst_n), .A1(_zy_sva_b1), .Z(n25));
Q_AN02 U265 ( .A0(rst_n), .A1(_zy_sva_b2), .Z(n26));
Q_AN02 U266 ( .A0(rst_n), .A1(_zy_sva_b3), .Z(n27));
Q_AN02 U267 ( .A0(rst_n), .A1(_zy_sva_b4), .Z(n28));
Q_AN02 U268 ( .A0(rst_n), .A1(_zy_sva_b5), .Z(n29));
Q_AN02 U269 ( .A0(rst_n), .A1(_zy_sva_b6), .Z(n30));
Q_AN02 U270 ( .A0(rst_n), .A1(_zy_sva_b7), .Z(n31));
Q_AN02 U271 ( .A0(rst_n), .A1(_zy_sva_b8), .Z(n32));
Q_AN02 U272 ( .A0(rst_n), .A1(_zy_sva_b9), .Z(n33));
Q_FDP1 kim_rd_q_REG  ( .CK(clk), .R(rst_n), .D(kim_rd), .Q(kim_rd_q), .QN(n642));
Q_FDP1 \cur_state_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_state[0]), .Q(cur_state[0]), .QN(n51));
Q_FDP1 \cur_state_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_state[1]), .Q(cur_state[1]), .QN(n46));
Q_FDP1 \cur_state_REG[2] ( .CK(clk), .R(rst_n), .D(nxt_state[2]), .Q(cur_state[2]), .QN(n53));
Q_INV U277 ( .A(parser_kimreader_data[65]), .Z(n34));
Q_OR03 U278 ( .A0(parser_kimreader_data[67]), .A1(parser_kimreader_data[66]), .A2(n34), .Z(n35));
Q_NR02 U279 ( .A0(parser_kimreader_data[64]), .A1(n35), .Z(n36));
Q_AN02 U280 ( .A0(n36), .A1(parser_kimreader_data[69]), .Z(n70));
Q_INV U281 ( .A(parser_kimreader_data[64]), .Z(n37));
Q_NR02 U282 ( .A0(n37), .A1(n2), .Z(n38));
Q_OR02 U283 ( .A0(parser_kimreader_data[14]), .A1(parser_kimreader_data[31]), .Z(n39));
Q_AN03 U284 ( .A0(n38), .A1(n39), .A2(parser_kimreader_data[15]), .Z(n71));
Q_AN03 U285 ( .A0(kimreader_ckvreader_valid), .A1(kimreader_ckvreader_data[69]), .A2(ckvreader_kimreader_ack), .Z(n72));
Q_XNR2 U286 ( .A0(n67), .A1(n40), .Z(nxt_state[0]));
Q_AN02 U287 ( .A0(n68), .A1(n69), .Z(n40));
Q_INV U288 ( .A(n69), .Z(nxt_state[1]));
Q_INV U289 ( .A(n41), .Z(nxt_state[2]));
Q_MX02 U290 ( .S(n67), .A0(n42), .A1(n43), .Z(n41));
Q_NR02 U291 ( .A0(n68), .A1(n69), .Z(n42));
Q_OR02 U292 ( .A0(n56), .A1(n69), .Z(n43));
Q_MX02 U293 ( .S(cur_state[2]), .A0(n44), .A1(n52), .Z(n67));
Q_MX02 U294 ( .S(cur_state[1]), .A0(n45), .A1(n50), .Z(n44));
Q_OR03 U295 ( .A0(cur_state[0]), .A1(n48), .A2(n47), .Z(n45));
Q_INV U296 ( .A(kimreader_parser_ack), .Z(n48));
Q_OR02 U297 ( .A0(n70), .A1(n49), .Z(n47));
Q_INV U298 ( .A(n71), .Z(n49));
Q_MX02 U299 ( .S(cur_state[0]), .A0(n348), .A1(n72), .Z(n50));
Q_MX02 U300 ( .S(cur_state[1]), .A0(n54), .A1(n55), .Z(n52));
Q_INV U301 ( .A(n56), .Z(n68));
Q_MX02 U302 ( .S(cur_state[2]), .A0(n57), .A1(n61), .Z(n56));
Q_OR03 U303 ( .A0(n58), .A1(n59), .A2(cur_state[1]), .Z(n57));
Q_NR02 U304 ( .A0(n60), .A1(cur_state[0]), .Z(n59));
Q_OA21 U305 ( .A0(n70), .A1(n71), .B0(kimreader_parser_ack), .Z(n60));
Q_AN02 U306 ( .A0(kim_rd), .A1(cur_state[0]), .Z(n58));
Q_MX02 U307 ( .S(cur_state[1]), .A0(n62), .A1(n54), .Z(n61));
Q_INV U308 ( .A(n55), .Z(n62));
Q_XNR2 U309 ( .A0(cur_state[0]), .A1(ckvreader_kimreader_ack), .Z(n55));
Q_MX02 U310 ( .S(cur_state[2]), .A0(n63), .A1(n66), .Z(n69));
Q_MX02 U311 ( .S(cur_state[1]), .A0(n64), .A1(n65), .Z(n63));
Q_INV U312 ( .A(n58), .Z(n64));
Q_AN02 U313 ( .A0(cur_state[0]), .A1(n72), .Z(n65));
Q_XNR2 U314 ( .A0(cur_state[1]), .A1(n54), .Z(n66));
Q_AN02 U315 ( .A0(cur_state[0]), .A1(ckvreader_kimreader_ack), .Z(n54));
Q_AN03 U316 ( .A0(parser_kimreader_data[67]), .A1(parser_kimreader_data[66]), .A2(parser_kimreader_data[65]), .Z(n73));
Q_AN02 U317 ( .A0(parser_kimreader_data[64]), .A1(n73), .Z(n378));
Q_INV U318 ( .A(parser_kimreader_data[66]), .Z(n74));
Q_OR03 U319 ( .A0(parser_kimreader_data[67]), .A1(n74), .A2(parser_kimreader_data[65]), .Z(n75));
Q_NR02 U320 ( .A0(parser_kimreader_data[64]), .A1(n75), .Z(n76));
Q_AN02 U321 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[0]), .Z(n77));
Q_AN02 U322 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[1]), .Z(n78));
Q_AN02 U323 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[2]), .Z(n79));
Q_AN02 U324 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[3]), .Z(n80));
Q_AN02 U325 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[4]), .Z(n81));
Q_AN02 U326 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[5]), .Z(n82));
Q_AN02 U327 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[6]), .Z(n83));
Q_AN02 U328 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[7]), .Z(n84));
Q_AN02 U329 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[8]), .Z(n85));
Q_AN02 U330 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[9]), .Z(n86));
Q_AN02 U331 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[10]), .Z(n87));
Q_AN02 U332 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[11]), .Z(n88));
Q_AN02 U333 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[12]), .Z(n89));
Q_AN02 U334 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[13]), .Z(n90));
Q_AN02 U335 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[14]), .Z(n91));
Q_AN02 U336 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[15]), .Z(n92));
Q_AN02 U337 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[16]), .Z(n93));
Q_AN02 U338 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[17]), .Z(n94));
Q_AN02 U339 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[18]), .Z(n95));
Q_AN02 U340 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[19]), .Z(n96));
Q_AN02 U341 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[20]), .Z(n97));
Q_AN02 U342 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[21]), .Z(n98));
Q_AN02 U343 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[22]), .Z(n99));
Q_AN02 U344 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[23]), .Z(n100));
Q_AN02 U345 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[24]), .Z(n101));
Q_AN02 U346 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[25]), .Z(n102));
Q_AN02 U347 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[26]), .Z(n103));
Q_AN02 U348 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[27]), .Z(n104));
Q_AN02 U349 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[28]), .Z(n105));
Q_AN02 U350 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[29]), .Z(n106));
Q_AN02 U351 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[30]), .Z(n107));
Q_AN02 U352 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[31]), .Z(n108));
Q_AN02 U353 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[32]), .Z(n109));
Q_AN02 U354 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[33]), .Z(n110));
Q_AN02 U355 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[34]), .Z(n111));
Q_AN02 U356 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[35]), .Z(n112));
Q_AN02 U357 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[36]), .Z(n113));
Q_AN02 U358 ( .A0(parser_kimreader_data[17]), .A1(dek_kim_entry_q[37]), .Z(n114));
Q_AN02 U359 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[0]), .Z(n115));
Q_AN02 U360 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[1]), .Z(n116));
Q_AN02 U361 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[2]), .Z(n117));
Q_AN02 U362 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[3]), .Z(n118));
Q_AN02 U363 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[4]), .Z(n119));
Q_AN02 U364 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[5]), .Z(n120));
Q_AN02 U365 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[6]), .Z(n121));
Q_AN02 U366 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[7]), .Z(n122));
Q_AN02 U367 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[8]), .Z(n123));
Q_AN02 U368 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[9]), .Z(n124));
Q_AN02 U369 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[10]), .Z(n125));
Q_AN02 U370 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[11]), .Z(n126));
Q_AN02 U371 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[12]), .Z(n127));
Q_AN02 U372 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[13]), .Z(n128));
Q_AN02 U373 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[14]), .Z(n129));
Q_AN02 U374 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[15]), .Z(n130));
Q_AN02 U375 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[16]), .Z(n131));
Q_AN02 U376 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[17]), .Z(n132));
Q_AN02 U377 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[18]), .Z(n133));
Q_AN02 U378 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[19]), .Z(n134));
Q_AN02 U379 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[20]), .Z(n135));
Q_AN02 U380 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[21]), .Z(n136));
Q_AN02 U381 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[22]), .Z(n137));
Q_AN02 U382 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[23]), .Z(n138));
Q_AN02 U383 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[24]), .Z(n139));
Q_AN02 U384 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[25]), .Z(n140));
Q_AN02 U385 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[26]), .Z(n141));
Q_AN02 U386 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[27]), .Z(n142));
Q_AN02 U387 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[28]), .Z(n143));
Q_AN02 U388 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[29]), .Z(n144));
Q_AN02 U389 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[30]), .Z(n145));
Q_AN02 U390 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[31]), .Z(n146));
Q_AN02 U391 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[32]), .Z(n147));
Q_AN02 U392 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[33]), .Z(n148));
Q_AN02 U393 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[34]), .Z(n149));
Q_AN02 U394 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[35]), .Z(n150));
Q_AN02 U395 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[36]), .Z(n151));
Q_AN02 U396 ( .A0(parser_kimreader_data[17]), .A1(dak_kim_entry_q[37]), .Z(n152));
Q_AN02 U397 ( .A0(n342), .A1(n77), .Z(tlv_word8[26]));
Q_AN02 U398 ( .A0(n342), .A1(n78), .Z(tlv_word8[27]));
Q_AN02 U399 ( .A0(n342), .A1(n79), .Z(tlv_word8[28]));
Q_AN02 U400 ( .A0(n342), .A1(n80), .Z(tlv_word8[29]));
Q_AN02 U401 ( .A0(n342), .A1(n81), .Z(tlv_word8[30]));
Q_AN02 U402 ( .A0(n342), .A1(n82), .Z(tlv_word8[31]));
Q_AN02 U403 ( .A0(n342), .A1(n83), .Z(tlv_word8[32]));
Q_AN02 U404 ( .A0(n342), .A1(n84), .Z(tlv_word8[33]));
Q_AN02 U405 ( .A0(n342), .A1(n85), .Z(tlv_word8[34]));
Q_AN02 U406 ( .A0(n342), .A1(n86), .Z(tlv_word8[35]));
Q_AN02 U407 ( .A0(n342), .A1(n87), .Z(tlv_word8[36]));
Q_AN02 U408 ( .A0(n342), .A1(n88), .Z(tlv_word8[37]));
Q_AN02 U409 ( .A0(n342), .A1(n89), .Z(tlv_word8[38]));
Q_AN02 U410 ( .A0(n342), .A1(n90), .Z(tlv_word8[39]));
Q_AN02 U411 ( .A0(n342), .A1(n91), .Z(tlv_word8[40]));
Q_AN02 U412 ( .A0(n342), .A1(n92), .Z(tlv_word8[41]));
Q_AN02 U413 ( .A0(n342), .A1(n93), .Z(tlv_word8[42]));
Q_AN02 U414 ( .A0(n342), .A1(n94), .Z(tlv_word8[43]));
Q_AN02 U415 ( .A0(n342), .A1(n95), .Z(tlv_word8[44]));
Q_AN02 U416 ( .A0(n342), .A1(n96), .Z(tlv_word8[45]));
Q_AN02 U417 ( .A0(n342), .A1(n97), .Z(tlv_word8[46]));
Q_AN02 U418 ( .A0(n342), .A1(n98), .Z(tlv_word8[47]));
Q_AN02 U419 ( .A0(n342), .A1(n99), .Z(tlv_word8[48]));
Q_AN02 U420 ( .A0(n342), .A1(n100), .Z(tlv_word8[49]));
Q_AN02 U421 ( .A0(n342), .A1(n101), .Z(tlv_word8[50]));
Q_AN02 U422 ( .A0(n342), .A1(n102), .Z(tlv_word8[51]));
Q_AN02 U423 ( .A0(n342), .A1(n103), .Z(tlv_word8[52]));
Q_AN02 U424 ( .A0(n342), .A1(n104), .Z(tlv_word8[53]));
Q_AN02 U425 ( .A0(n342), .A1(n105), .Z(tlv_word8[54]));
Q_AN02 U426 ( .A0(n342), .A1(n106), .Z(tlv_word8[55]));
Q_AN02 U427 ( .A0(n342), .A1(n107), .Z(tlv_word8[56]));
Q_AN02 U428 ( .A0(n342), .A1(n108), .Z(tlv_word8[57]));
Q_AN02 U429 ( .A0(n342), .A1(n109), .Z(tlv_word8[58]));
Q_AN02 U430 ( .A0(n342), .A1(n110), .Z(tlv_word8[59]));
Q_AN02 U431 ( .A0(n342), .A1(n111), .Z(tlv_word8[60]));
Q_AN02 U432 ( .A0(n342), .A1(n112), .Z(tlv_word8[61]));
Q_AN02 U433 ( .A0(n342), .A1(n113), .Z(tlv_word8[62]));
Q_AN02 U434 ( .A0(n342), .A1(n114), .Z(tlv_word8[63]));
Q_AN02 U435 ( .A0(n342), .A1(parser_kimreader_data[0]), .Z(tlv_word9[0]));
Q_AN02 U436 ( .A0(n342), .A1(parser_kimreader_data[1]), .Z(tlv_word9[1]));
Q_AN02 U437 ( .A0(n342), .A1(parser_kimreader_data[2]), .Z(tlv_word9[2]));
Q_AN02 U438 ( .A0(n342), .A1(parser_kimreader_data[3]), .Z(tlv_word9[3]));
Q_AN02 U439 ( .A0(n342), .A1(parser_kimreader_data[4]), .Z(tlv_word9[4]));
Q_AN02 U440 ( .A0(n342), .A1(parser_kimreader_data[5]), .Z(tlv_word9[5]));
Q_AN02 U441 ( .A0(n342), .A1(parser_kimreader_data[6]), .Z(tlv_word9[6]));
Q_AN02 U442 ( .A0(n342), .A1(parser_kimreader_data[7]), .Z(tlv_word9[7]));
Q_AN02 U443 ( .A0(n342), .A1(parser_kimreader_data[8]), .Z(tlv_word9[8]));
Q_AN02 U444 ( .A0(n342), .A1(parser_kimreader_data[9]), .Z(tlv_word9[9]));
Q_AN02 U445 ( .A0(n342), .A1(parser_kimreader_data[10]), .Z(tlv_word9[10]));
Q_AN02 U446 ( .A0(n342), .A1(parser_kimreader_data[11]), .Z(tlv_word9[11]));
Q_AN02 U447 ( .A0(n342), .A1(parser_kimreader_data[12]), .Z(tlv_word9[12]));
Q_AN02 U448 ( .A0(n342), .A1(parser_kimreader_data[13]), .Z(tlv_word9[13]));
Q_AN02 U449 ( .A0(n342), .A1(parser_kimreader_data[14]), .Z(tlv_word9[14]));
Q_AN02 U450 ( .A0(n342), .A1(parser_kimreader_data[15]), .Z(tlv_word9[15]));
Q_AN02 U451 ( .A0(n342), .A1(parser_kimreader_data[16]), .Z(tlv_word9[16]));
Q_AN02 U452 ( .A0(n342), .A1(parser_kimreader_data[20]), .Z(tlv_word9[20]));
Q_AN02 U453 ( .A0(n342), .A1(parser_kimreader_data[21]), .Z(tlv_word9[21]));
Q_AN02 U454 ( .A0(n342), .A1(parser_kimreader_data[22]), .Z(tlv_word9[22]));
Q_AN02 U455 ( .A0(n342), .A1(parser_kimreader_data[23]), .Z(tlv_word9[23]));
Q_AN02 U456 ( .A0(n342), .A1(parser_kimreader_data[24]), .Z(tlv_word9[24]));
Q_AN02 U457 ( .A0(n342), .A1(parser_kimreader_data[25]), .Z(tlv_word9[25]));
Q_AN02 U458 ( .A0(n342), .A1(n115), .Z(tlv_word9[26]));
Q_AN02 U459 ( .A0(n342), .A1(n116), .Z(tlv_word9[27]));
Q_AN02 U460 ( .A0(n342), .A1(n117), .Z(tlv_word9[28]));
Q_AN02 U461 ( .A0(n342), .A1(n118), .Z(tlv_word9[29]));
Q_AN02 U462 ( .A0(n342), .A1(n119), .Z(tlv_word9[30]));
Q_AN02 U463 ( .A0(n342), .A1(n120), .Z(tlv_word9[31]));
Q_AN02 U464 ( .A0(n342), .A1(n121), .Z(tlv_word9[32]));
Q_AN02 U465 ( .A0(n342), .A1(n122), .Z(tlv_word9[33]));
Q_AN02 U466 ( .A0(n342), .A1(n123), .Z(tlv_word9[34]));
Q_AN02 U467 ( .A0(n342), .A1(n124), .Z(tlv_word9[35]));
Q_AN02 U468 ( .A0(n342), .A1(n125), .Z(tlv_word9[36]));
Q_AN02 U469 ( .A0(n342), .A1(n126), .Z(tlv_word9[37]));
Q_AN02 U470 ( .A0(n342), .A1(n127), .Z(tlv_word9[38]));
Q_AN02 U471 ( .A0(n342), .A1(n128), .Z(tlv_word9[39]));
Q_AN02 U472 ( .A0(n342), .A1(n129), .Z(tlv_word9[40]));
Q_AN02 U473 ( .A0(n342), .A1(n130), .Z(tlv_word9[41]));
Q_AN02 U474 ( .A0(n342), .A1(n131), .Z(tlv_word9[42]));
Q_AN02 U475 ( .A0(n342), .A1(n132), .Z(tlv_word9[43]));
Q_AN02 U476 ( .A0(n342), .A1(n133), .Z(tlv_word9[44]));
Q_AN02 U477 ( .A0(n342), .A1(n134), .Z(tlv_word9[45]));
Q_AN02 U478 ( .A0(n342), .A1(n135), .Z(tlv_word9[46]));
Q_AN02 U479 ( .A0(n342), .A1(n136), .Z(tlv_word9[47]));
Q_AN02 U480 ( .A0(n342), .A1(n137), .Z(tlv_word9[48]));
Q_AN02 U481 ( .A0(n342), .A1(n138), .Z(tlv_word9[49]));
Q_AN02 U482 ( .A0(n342), .A1(n139), .Z(tlv_word9[50]));
Q_AN02 U483 ( .A0(n342), .A1(n140), .Z(tlv_word9[51]));
Q_AN02 U484 ( .A0(n342), .A1(n141), .Z(tlv_word9[52]));
Q_AN02 U485 ( .A0(n342), .A1(n142), .Z(tlv_word9[53]));
Q_AN02 U486 ( .A0(n342), .A1(n143), .Z(tlv_word9[54]));
Q_AN02 U487 ( .A0(n342), .A1(n144), .Z(tlv_word9[55]));
Q_AN02 U488 ( .A0(n342), .A1(n145), .Z(tlv_word9[56]));
Q_AN02 U489 ( .A0(n342), .A1(n146), .Z(tlv_word9[57]));
Q_AN02 U490 ( .A0(n342), .A1(n147), .Z(tlv_word9[58]));
Q_AN02 U491 ( .A0(n342), .A1(n148), .Z(tlv_word9[59]));
Q_AN02 U492 ( .A0(n342), .A1(n149), .Z(tlv_word9[60]));
Q_AN02 U493 ( .A0(n342), .A1(n150), .Z(tlv_word9[61]));
Q_AN02 U494 ( .A0(n342), .A1(n151), .Z(tlv_word9[62]));
Q_AN02 U495 ( .A0(n342), .A1(n152), .Z(tlv_word9[63]));
Q_AN02 U496 ( .A0(n342), .A1(parser_kimreader_data[17]), .Z(tlv_word8[17]));
Q_AN02 U497 ( .A0(n342), .A1(parser_kimreader_data[18]), .Z(tlv_word8[18]));
Q_AN02 U498 ( .A0(n342), .A1(parser_kimreader_data[19]), .Z(tlv_word8[19]));
Q_AN02 U499 ( .A0(n345), .A1(dek_ref_q[0]), .Z(n153));
Q_MX02 U500 ( .S(n346), .A0(n153), .A1(dak_ref_q[0]), .Z(kim_addr[0]));
Q_AN02 U501 ( .A0(n345), .A1(dek_ref_q[1]), .Z(n154));
Q_MX02 U502 ( .S(n346), .A0(n154), .A1(dak_ref_q[1]), .Z(kim_addr[1]));
Q_AN02 U503 ( .A0(n345), .A1(dek_ref_q[2]), .Z(n155));
Q_MX02 U504 ( .S(n346), .A0(n155), .A1(dak_ref_q[2]), .Z(kim_addr[2]));
Q_AN02 U505 ( .A0(n345), .A1(dek_ref_q[3]), .Z(n156));
Q_MX02 U506 ( .S(n346), .A0(n156), .A1(dak_ref_q[3]), .Z(kim_addr[3]));
Q_AN02 U507 ( .A0(n345), .A1(dek_ref_q[4]), .Z(n157));
Q_MX02 U508 ( .S(n346), .A0(n157), .A1(dak_ref_q[4]), .Z(kim_addr[4]));
Q_AN02 U509 ( .A0(n345), .A1(dek_ref_q[5]), .Z(n158));
Q_MX02 U510 ( .S(n346), .A0(n158), .A1(dak_ref_q[5]), .Z(kim_addr[5]));
Q_AN02 U511 ( .A0(n345), .A1(dek_ref_q[6]), .Z(n159));
Q_MX02 U512 ( .S(n346), .A0(n159), .A1(dak_ref_q[6]), .Z(kim_addr[6]));
Q_AN02 U513 ( .A0(n345), .A1(dek_ref_q[7]), .Z(n160));
Q_MX02 U514 ( .S(n346), .A0(n160), .A1(dak_ref_q[7]), .Z(kim_addr[7]));
Q_AN02 U515 ( .A0(n345), .A1(dek_ref_q[8]), .Z(n161));
Q_MX02 U516 ( .S(n346), .A0(n161), .A1(dak_ref_q[8]), .Z(kim_addr[8]));
Q_AN02 U517 ( .A0(n345), .A1(dek_ref_q[9]), .Z(n162));
Q_MX02 U518 ( .S(n346), .A0(n162), .A1(dak_ref_q[9]), .Z(kim_addr[9]));
Q_AN02 U519 ( .A0(n345), .A1(dek_ref_q[10]), .Z(n163));
Q_MX02 U520 ( .S(n346), .A0(n163), .A1(dak_ref_q[10]), .Z(kim_addr[10]));
Q_AN02 U521 ( .A0(n345), .A1(dek_ref_q[11]), .Z(n164));
Q_MX02 U522 ( .S(n346), .A0(n164), .A1(dak_ref_q[11]), .Z(kim_addr[11]));
Q_AN02 U523 ( .A0(n345), .A1(dek_ref_q[12]), .Z(n165));
Q_MX02 U524 ( .S(n346), .A0(n165), .A1(dak_ref_q[12]), .Z(kim_addr[12]));
Q_AN02 U525 ( .A0(n345), .A1(dek_ref_q[13]), .Z(n166));
Q_MX02 U526 ( .S(n346), .A0(n166), .A1(dak_ref_q[13]), .Z(kim_addr[13]));
Q_MX03 U527 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[0]), .A1(drng_256_out[0]), .A2(drng_256_out[64]), .Z(n167));
Q_MX02 U528 ( .S(n373), .A0(parser_kimreader_data[0]), .A1(tlv_word42[0]), .Z(n168));
Q_AN02 U529 ( .A0(n373), .A1(parser_kimreader_data[0]), .Z(n169));
Q_MX03 U530 ( .S0(n374), .S1(n375), .A0(n169), .A1(n168), .A2(n167), .Z(kimreader_ckvreader_data[0]));
Q_MX03 U531 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[1]), .A1(drng_256_out[1]), .A2(drng_256_out[65]), .Z(n170));
Q_MX02 U532 ( .S(n373), .A0(parser_kimreader_data[1]), .A1(tlv_word42[1]), .Z(n171));
Q_AN02 U533 ( .A0(n373), .A1(parser_kimreader_data[1]), .Z(n172));
Q_MX03 U534 ( .S0(n374), .S1(n375), .A0(n172), .A1(n171), .A2(n170), .Z(kimreader_ckvreader_data[1]));
Q_MX03 U535 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[2]), .A1(drng_256_out[2]), .A2(drng_256_out[66]), .Z(n173));
Q_MX02 U536 ( .S(n373), .A0(parser_kimreader_data[2]), .A1(tlv_word42[2]), .Z(n174));
Q_AN02 U537 ( .A0(n373), .A1(parser_kimreader_data[2]), .Z(n175));
Q_MX03 U538 ( .S0(n374), .S1(n375), .A0(n175), .A1(n174), .A2(n173), .Z(kimreader_ckvreader_data[2]));
Q_MX03 U539 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[3]), .A1(drng_256_out[3]), .A2(drng_256_out[67]), .Z(n176));
Q_MX02 U540 ( .S(n373), .A0(parser_kimreader_data[3]), .A1(tlv_word42[3]), .Z(n177));
Q_AN02 U541 ( .A0(n373), .A1(parser_kimreader_data[3]), .Z(n178));
Q_MX03 U542 ( .S0(n374), .S1(n375), .A0(n178), .A1(n177), .A2(n176), .Z(kimreader_ckvreader_data[3]));
Q_MX03 U543 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[4]), .A1(drng_256_out[4]), .A2(drng_256_out[68]), .Z(n179));
Q_MX02 U544 ( .S(n373), .A0(parser_kimreader_data[4]), .A1(tlv_word42[4]), .Z(n180));
Q_AN02 U545 ( .A0(n373), .A1(parser_kimreader_data[4]), .Z(n181));
Q_MX03 U546 ( .S0(n374), .S1(n375), .A0(n181), .A1(n180), .A2(n179), .Z(kimreader_ckvreader_data[4]));
Q_MX03 U547 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[5]), .A1(drng_256_out[5]), .A2(drng_256_out[69]), .Z(n182));
Q_MX02 U548 ( .S(n373), .A0(parser_kimreader_data[5]), .A1(tlv_word42[5]), .Z(n183));
Q_AN02 U549 ( .A0(n373), .A1(parser_kimreader_data[5]), .Z(n184));
Q_MX03 U550 ( .S0(n374), .S1(n375), .A0(n184), .A1(n183), .A2(n182), .Z(kimreader_ckvreader_data[5]));
Q_MX03 U551 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[6]), .A1(drng_256_out[6]), .A2(drng_256_out[70]), .Z(n185));
Q_MX02 U552 ( .S(n373), .A0(parser_kimreader_data[6]), .A1(tlv_word42[6]), .Z(n186));
Q_AN02 U553 ( .A0(n373), .A1(parser_kimreader_data[6]), .Z(n187));
Q_MX03 U554 ( .S0(n374), .S1(n375), .A0(n187), .A1(n186), .A2(n185), .Z(kimreader_ckvreader_data[6]));
Q_MX03 U555 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[7]), .A1(drng_256_out[7]), .A2(drng_256_out[71]), .Z(n188));
Q_MX02 U556 ( .S(n373), .A0(parser_kimreader_data[7]), .A1(tlv_word42[7]), .Z(n189));
Q_AN02 U557 ( .A0(n373), .A1(parser_kimreader_data[7]), .Z(n190));
Q_MX03 U558 ( .S0(n374), .S1(n375), .A0(n190), .A1(n189), .A2(n188), .Z(kimreader_ckvreader_data[7]));
Q_MX03 U559 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[8]), .A1(drng_256_out[8]), .A2(drng_256_out[72]), .Z(n191));
Q_AN02 U560 ( .A0(n1), .A1(parser_kimreader_data[8]), .Z(n192));
Q_MX02 U561 ( .S(n375), .A0(n192), .A1(n191), .Z(kimreader_ckvreader_data[8]));
Q_MX03 U562 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[9]), .A1(drng_256_out[9]), .A2(drng_256_out[73]), .Z(n193));
Q_AN02 U563 ( .A0(n1), .A1(parser_kimreader_data[9]), .Z(n194));
Q_MX02 U564 ( .S(n375), .A0(n194), .A1(n193), .Z(kimreader_ckvreader_data[9]));
Q_MX03 U565 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[10]), .A1(drng_256_out[10]), .A2(drng_256_out[74]), .Z(n195));
Q_AN02 U566 ( .A0(n1), .A1(parser_kimreader_data[10]), .Z(n196));
Q_MX02 U567 ( .S(n375), .A0(n196), .A1(n195), .Z(kimreader_ckvreader_data[10]));
Q_MX03 U568 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[11]), .A1(drng_256_out[11]), .A2(drng_256_out[75]), .Z(n197));
Q_AN02 U569 ( .A0(n1), .A1(parser_kimreader_data[11]), .Z(n198));
Q_MX02 U570 ( .S(n375), .A0(n198), .A1(n197), .Z(kimreader_ckvreader_data[11]));
Q_MX03 U571 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[12]), .A1(drng_256_out[12]), .A2(drng_256_out[76]), .Z(n199));
Q_AN02 U572 ( .A0(n1), .A1(parser_kimreader_data[12]), .Z(n200));
Q_MX02 U573 ( .S(n375), .A0(n200), .A1(n199), .Z(kimreader_ckvreader_data[12]));
Q_MX03 U574 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[13]), .A1(drng_256_out[13]), .A2(drng_256_out[77]), .Z(n201));
Q_AN02 U575 ( .A0(n1), .A1(parser_kimreader_data[13]), .Z(n202));
Q_MX02 U576 ( .S(n375), .A0(n202), .A1(n201), .Z(kimreader_ckvreader_data[13]));
Q_MX03 U577 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[14]), .A1(drng_256_out[14]), .A2(drng_256_out[78]), .Z(n203));
Q_AN02 U578 ( .A0(n1), .A1(parser_kimreader_data[14]), .Z(n204));
Q_MX02 U579 ( .S(n375), .A0(n204), .A1(n203), .Z(kimreader_ckvreader_data[14]));
Q_MX03 U580 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[15]), .A1(drng_256_out[15]), .A2(drng_256_out[79]), .Z(n205));
Q_AN02 U581 ( .A0(n1), .A1(parser_kimreader_data[15]), .Z(n206));
Q_MX02 U582 ( .S(n375), .A0(n206), .A1(n205), .Z(kimreader_ckvreader_data[15]));
Q_MX03 U583 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[16]), .A1(drng_256_out[16]), .A2(drng_256_out[80]), .Z(n207));
Q_AN02 U584 ( .A0(n1), .A1(parser_kimreader_data[16]), .Z(n208));
Q_MX02 U585 ( .S(n375), .A0(n208), .A1(n207), .Z(kimreader_ckvreader_data[16]));
Q_MX03 U586 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[17]), .A1(drng_256_out[17]), .A2(drng_256_out[81]), .Z(n209));
Q_AN02 U587 ( .A0(n1), .A1(parser_kimreader_data[17]), .Z(n210));
Q_MX02 U588 ( .S(n375), .A0(n210), .A1(n209), .Z(kimreader_ckvreader_data[17]));
Q_MX03 U589 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[18]), .A1(drng_256_out[18]), .A2(drng_256_out[82]), .Z(n211));
Q_AN02 U590 ( .A0(n1), .A1(parser_kimreader_data[18]), .Z(n212));
Q_MX02 U591 ( .S(n375), .A0(n212), .A1(n211), .Z(kimreader_ckvreader_data[18]));
Q_MX03 U592 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[19]), .A1(drng_256_out[19]), .A2(drng_256_out[83]), .Z(n213));
Q_AN02 U593 ( .A0(n1), .A1(parser_kimreader_data[19]), .Z(n214));
Q_MX02 U594 ( .S(n375), .A0(n214), .A1(n213), .Z(kimreader_ckvreader_data[19]));
Q_MX03 U595 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[20]), .A1(drng_256_out[20]), .A2(drng_256_out[84]), .Z(n215));
Q_AN02 U596 ( .A0(n1), .A1(parser_kimreader_data[20]), .Z(n216));
Q_MX02 U597 ( .S(n375), .A0(n216), .A1(n215), .Z(kimreader_ckvreader_data[20]));
Q_MX03 U598 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[21]), .A1(drng_256_out[21]), .A2(drng_256_out[85]), .Z(n217));
Q_AN02 U599 ( .A0(n1), .A1(parser_kimreader_data[21]), .Z(n218));
Q_MX02 U600 ( .S(n375), .A0(n218), .A1(n217), .Z(kimreader_ckvreader_data[21]));
Q_MX03 U601 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[22]), .A1(drng_256_out[22]), .A2(drng_256_out[86]), .Z(n219));
Q_AN02 U602 ( .A0(n1), .A1(parser_kimreader_data[22]), .Z(n220));
Q_MX02 U603 ( .S(n375), .A0(n220), .A1(n219), .Z(kimreader_ckvreader_data[22]));
Q_MX03 U604 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[23]), .A1(drng_256_out[23]), .A2(drng_256_out[87]), .Z(n221));
Q_AN02 U605 ( .A0(n1), .A1(parser_kimreader_data[23]), .Z(n222));
Q_MX02 U606 ( .S(n375), .A0(n222), .A1(n221), .Z(kimreader_ckvreader_data[23]));
Q_MX03 U607 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[24]), .A1(drng_256_out[24]), .A2(drng_256_out[88]), .Z(n223));
Q_AN02 U608 ( .A0(n1), .A1(parser_kimreader_data[24]), .Z(n224));
Q_MX02 U609 ( .S(n375), .A0(n224), .A1(n223), .Z(kimreader_ckvreader_data[24]));
Q_MX03 U610 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[25]), .A1(drng_256_out[25]), .A2(drng_256_out[89]), .Z(n225));
Q_AN02 U611 ( .A0(n1), .A1(parser_kimreader_data[25]), .Z(n226));
Q_MX02 U612 ( .S(n375), .A0(n226), .A1(n225), .Z(kimreader_ckvreader_data[25]));
Q_MX03 U613 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[26]), .A1(drng_256_out[26]), .A2(drng_256_out[90]), .Z(n227));
Q_MX02 U614 ( .S(n373), .A0(n77), .A1(parser_kimreader_data[26]), .Z(n228));
Q_AN02 U615 ( .A0(n373), .A1(n115), .Z(n229));
Q_MX03 U616 ( .S0(n374), .S1(n375), .A0(n229), .A1(n228), .A2(n227), .Z(kimreader_ckvreader_data[26]));
Q_MX03 U617 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[27]), .A1(drng_256_out[27]), .A2(drng_256_out[91]), .Z(n230));
Q_MX02 U618 ( .S(n373), .A0(n78), .A1(parser_kimreader_data[27]), .Z(n231));
Q_AN02 U619 ( .A0(n373), .A1(n116), .Z(n232));
Q_MX03 U620 ( .S0(n374), .S1(n375), .A0(n232), .A1(n231), .A2(n230), .Z(kimreader_ckvreader_data[27]));
Q_MX03 U621 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[28]), .A1(drng_256_out[28]), .A2(drng_256_out[92]), .Z(n233));
Q_MX02 U622 ( .S(n373), .A0(n79), .A1(parser_kimreader_data[28]), .Z(n234));
Q_AN02 U623 ( .A0(n373), .A1(n117), .Z(n235));
Q_MX03 U624 ( .S0(n374), .S1(n375), .A0(n235), .A1(n234), .A2(n233), .Z(kimreader_ckvreader_data[28]));
Q_MX03 U625 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[29]), .A1(drng_256_out[29]), .A2(drng_256_out[93]), .Z(n236));
Q_MX02 U626 ( .S(n373), .A0(n80), .A1(parser_kimreader_data[29]), .Z(n237));
Q_AN02 U627 ( .A0(n373), .A1(n118), .Z(n238));
Q_MX03 U628 ( .S0(n374), .S1(n375), .A0(n238), .A1(n237), .A2(n236), .Z(kimreader_ckvreader_data[29]));
Q_MX03 U629 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[30]), .A1(drng_256_out[30]), .A2(drng_256_out[94]), .Z(n239));
Q_MX02 U630 ( .S(n373), .A0(n81), .A1(parser_kimreader_data[30]), .Z(n240));
Q_AN02 U631 ( .A0(n373), .A1(n119), .Z(n241));
Q_MX03 U632 ( .S0(n374), .S1(n375), .A0(n241), .A1(n240), .A2(n239), .Z(kimreader_ckvreader_data[30]));
Q_MX03 U633 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[31]), .A1(drng_256_out[31]), .A2(drng_256_out[95]), .Z(n242));
Q_MX02 U634 ( .S(n373), .A0(n82), .A1(parser_kimreader_data[31]), .Z(n243));
Q_AN02 U635 ( .A0(n373), .A1(n120), .Z(n244));
Q_MX03 U636 ( .S0(n374), .S1(n375), .A0(n244), .A1(n243), .A2(n242), .Z(kimreader_ckvreader_data[31]));
Q_MX03 U637 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[32]), .A1(drng_256_out[32]), .A2(drng_256_out[96]), .Z(n245));
Q_MX02 U638 ( .S(n373), .A0(n83), .A1(parser_kimreader_data[32]), .Z(n246));
Q_AN02 U639 ( .A0(n373), .A1(n121), .Z(n247));
Q_MX03 U640 ( .S0(n374), .S1(n375), .A0(n247), .A1(n246), .A2(n245), .Z(kimreader_ckvreader_data[32]));
Q_MX03 U641 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[33]), .A1(drng_256_out[33]), .A2(drng_256_out[97]), .Z(n248));
Q_MX02 U642 ( .S(n373), .A0(n84), .A1(parser_kimreader_data[33]), .Z(n249));
Q_AN02 U643 ( .A0(n373), .A1(n122), .Z(n250));
Q_MX03 U644 ( .S0(n374), .S1(n375), .A0(n250), .A1(n249), .A2(n248), .Z(kimreader_ckvreader_data[33]));
Q_MX03 U645 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[34]), .A1(drng_256_out[34]), .A2(drng_256_out[98]), .Z(n251));
Q_MX02 U646 ( .S(n373), .A0(n85), .A1(parser_kimreader_data[34]), .Z(n252));
Q_AN02 U647 ( .A0(n373), .A1(n123), .Z(n253));
Q_MX03 U648 ( .S0(n374), .S1(n375), .A0(n253), .A1(n252), .A2(n251), .Z(kimreader_ckvreader_data[34]));
Q_MX03 U649 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[35]), .A1(drng_256_out[35]), .A2(drng_256_out[99]), .Z(n254));
Q_MX02 U650 ( .S(n373), .A0(n86), .A1(parser_kimreader_data[35]), .Z(n255));
Q_AN02 U651 ( .A0(n373), .A1(n124), .Z(n256));
Q_MX03 U652 ( .S0(n374), .S1(n375), .A0(n256), .A1(n255), .A2(n254), .Z(kimreader_ckvreader_data[35]));
Q_MX03 U653 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[36]), .A1(drng_256_out[36]), .A2(drng_256_out[100]), .Z(n257));
Q_MX02 U654 ( .S(n373), .A0(n87), .A1(parser_kimreader_data[36]), .Z(n258));
Q_AN02 U655 ( .A0(n373), .A1(n125), .Z(n259));
Q_MX03 U656 ( .S0(n374), .S1(n375), .A0(n259), .A1(n258), .A2(n257), .Z(kimreader_ckvreader_data[36]));
Q_MX03 U657 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[37]), .A1(drng_256_out[37]), .A2(drng_256_out[101]), .Z(n260));
Q_MX02 U658 ( .S(n373), .A0(n88), .A1(parser_kimreader_data[37]), .Z(n261));
Q_AN02 U659 ( .A0(n373), .A1(n126), .Z(n262));
Q_MX03 U660 ( .S0(n374), .S1(n375), .A0(n262), .A1(n261), .A2(n260), .Z(kimreader_ckvreader_data[37]));
Q_MX03 U661 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[38]), .A1(drng_256_out[38]), .A2(drng_256_out[102]), .Z(n263));
Q_MX02 U662 ( .S(n373), .A0(n89), .A1(parser_kimreader_data[38]), .Z(n264));
Q_AN02 U663 ( .A0(n373), .A1(n127), .Z(n265));
Q_MX03 U664 ( .S0(n374), .S1(n375), .A0(n265), .A1(n264), .A2(n263), .Z(kimreader_ckvreader_data[38]));
Q_MX03 U665 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[39]), .A1(drng_256_out[39]), .A2(drng_256_out[103]), .Z(n266));
Q_MX02 U666 ( .S(n373), .A0(n90), .A1(parser_kimreader_data[39]), .Z(n267));
Q_AN02 U667 ( .A0(n373), .A1(n128), .Z(n268));
Q_MX03 U668 ( .S0(n374), .S1(n375), .A0(n268), .A1(n267), .A2(n266), .Z(kimreader_ckvreader_data[39]));
Q_MX03 U669 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[40]), .A1(drng_256_out[40]), .A2(drng_256_out[104]), .Z(n269));
Q_MX02 U670 ( .S(n373), .A0(n91), .A1(parser_kimreader_data[40]), .Z(n270));
Q_AN02 U671 ( .A0(n373), .A1(n129), .Z(n271));
Q_MX03 U672 ( .S0(n374), .S1(n375), .A0(n271), .A1(n270), .A2(n269), .Z(kimreader_ckvreader_data[40]));
Q_MX03 U673 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[41]), .A1(drng_256_out[41]), .A2(drng_256_out[105]), .Z(n272));
Q_MX02 U674 ( .S(n373), .A0(n92), .A1(parser_kimreader_data[41]), .Z(n273));
Q_AN02 U675 ( .A0(n373), .A1(n130), .Z(n274));
Q_MX03 U676 ( .S0(n374), .S1(n375), .A0(n274), .A1(n273), .A2(n272), .Z(kimreader_ckvreader_data[41]));
Q_MX03 U677 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[42]), .A1(drng_256_out[42]), .A2(drng_256_out[106]), .Z(n275));
Q_MX02 U678 ( .S(n373), .A0(n93), .A1(parser_kimreader_data[42]), .Z(n276));
Q_AN02 U679 ( .A0(n373), .A1(n131), .Z(n277));
Q_MX03 U680 ( .S0(n374), .S1(n375), .A0(n277), .A1(n276), .A2(n275), .Z(kimreader_ckvreader_data[42]));
Q_MX03 U681 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[43]), .A1(drng_256_out[43]), .A2(drng_256_out[107]), .Z(n278));
Q_MX02 U682 ( .S(n373), .A0(n94), .A1(parser_kimreader_data[43]), .Z(n279));
Q_AN02 U683 ( .A0(n373), .A1(n132), .Z(n280));
Q_MX03 U684 ( .S0(n374), .S1(n375), .A0(n280), .A1(n279), .A2(n278), .Z(kimreader_ckvreader_data[43]));
Q_MX03 U685 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[44]), .A1(drng_256_out[44]), .A2(drng_256_out[108]), .Z(n281));
Q_MX02 U686 ( .S(n373), .A0(n95), .A1(parser_kimreader_data[44]), .Z(n282));
Q_AN02 U687 ( .A0(n373), .A1(n133), .Z(n283));
Q_MX03 U688 ( .S0(n374), .S1(n375), .A0(n283), .A1(n282), .A2(n281), .Z(kimreader_ckvreader_data[44]));
Q_MX03 U689 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[45]), .A1(drng_256_out[45]), .A2(drng_256_out[109]), .Z(n284));
Q_MX02 U690 ( .S(n373), .A0(n96), .A1(parser_kimreader_data[45]), .Z(n285));
Q_AN02 U691 ( .A0(n373), .A1(n134), .Z(n286));
Q_MX03 U692 ( .S0(n374), .S1(n375), .A0(n286), .A1(n285), .A2(n284), .Z(kimreader_ckvreader_data[45]));
Q_MX03 U693 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[46]), .A1(drng_256_out[46]), .A2(drng_256_out[110]), .Z(n287));
Q_MX02 U694 ( .S(n373), .A0(n97), .A1(parser_kimreader_data[46]), .Z(n288));
Q_AN02 U695 ( .A0(n373), .A1(n135), .Z(n289));
Q_MX03 U696 ( .S0(n374), .S1(n375), .A0(n289), .A1(n288), .A2(n287), .Z(kimreader_ckvreader_data[46]));
Q_MX03 U697 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[47]), .A1(drng_256_out[47]), .A2(drng_256_out[111]), .Z(n290));
Q_MX02 U698 ( .S(n373), .A0(n98), .A1(parser_kimreader_data[47]), .Z(n291));
Q_AN02 U699 ( .A0(n373), .A1(n136), .Z(n292));
Q_MX03 U700 ( .S0(n374), .S1(n375), .A0(n292), .A1(n291), .A2(n290), .Z(kimreader_ckvreader_data[47]));
Q_MX03 U701 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[48]), .A1(drng_256_out[48]), .A2(drng_256_out[112]), .Z(n293));
Q_MX02 U702 ( .S(n373), .A0(n99), .A1(parser_kimreader_data[48]), .Z(n294));
Q_AN02 U703 ( .A0(n373), .A1(n137), .Z(n295));
Q_MX03 U704 ( .S0(n374), .S1(n375), .A0(n295), .A1(n294), .A2(n293), .Z(kimreader_ckvreader_data[48]));
Q_MX03 U705 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[49]), .A1(drng_256_out[49]), .A2(drng_256_out[113]), .Z(n296));
Q_MX02 U706 ( .S(n373), .A0(n100), .A1(parser_kimreader_data[49]), .Z(n297));
Q_AN02 U707 ( .A0(n373), .A1(n138), .Z(n298));
Q_MX03 U708 ( .S0(n374), .S1(n375), .A0(n298), .A1(n297), .A2(n296), .Z(kimreader_ckvreader_data[49]));
Q_MX03 U709 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[50]), .A1(drng_256_out[50]), .A2(drng_256_out[114]), .Z(n299));
Q_MX02 U710 ( .S(n373), .A0(n101), .A1(parser_kimreader_data[50]), .Z(n300));
Q_AN02 U711 ( .A0(n373), .A1(n139), .Z(n301));
Q_MX03 U712 ( .S0(n374), .S1(n375), .A0(n301), .A1(n300), .A2(n299), .Z(kimreader_ckvreader_data[50]));
Q_MX03 U713 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[51]), .A1(drng_256_out[51]), .A2(drng_256_out[115]), .Z(n302));
Q_MX02 U714 ( .S(n373), .A0(n102), .A1(parser_kimreader_data[51]), .Z(n303));
Q_AN02 U715 ( .A0(n373), .A1(n140), .Z(n304));
Q_MX03 U716 ( .S0(n374), .S1(n375), .A0(n304), .A1(n303), .A2(n302), .Z(kimreader_ckvreader_data[51]));
Q_MX03 U717 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[52]), .A1(drng_256_out[52]), .A2(drng_256_out[116]), .Z(n305));
Q_MX02 U718 ( .S(n373), .A0(n103), .A1(parser_kimreader_data[52]), .Z(n306));
Q_AN02 U719 ( .A0(n373), .A1(n141), .Z(n307));
Q_MX03 U720 ( .S0(n374), .S1(n375), .A0(n307), .A1(n306), .A2(n305), .Z(kimreader_ckvreader_data[52]));
Q_MX03 U721 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[53]), .A1(drng_256_out[53]), .A2(drng_256_out[117]), .Z(n308));
Q_MX02 U722 ( .S(n373), .A0(n104), .A1(parser_kimreader_data[53]), .Z(n309));
Q_AN02 U723 ( .A0(n373), .A1(n142), .Z(n310));
Q_MX03 U724 ( .S0(n374), .S1(n375), .A0(n310), .A1(n309), .A2(n308), .Z(kimreader_ckvreader_data[53]));
Q_MX03 U725 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[54]), .A1(drng_256_out[54]), .A2(drng_256_out[118]), .Z(n311));
Q_MX02 U726 ( .S(n373), .A0(n105), .A1(parser_kimreader_data[54]), .Z(n312));
Q_AN02 U727 ( .A0(n373), .A1(n143), .Z(n313));
Q_MX03 U728 ( .S0(n374), .S1(n375), .A0(n313), .A1(n312), .A2(n311), .Z(kimreader_ckvreader_data[54]));
Q_MX03 U729 ( .S0(n373), .S1(n374), .A0(parser_kimreader_data[55]), .A1(drng_256_out[55]), .A2(drng_256_out[119]), .Z(n314));
Q_MX02 U730 ( .S(n373), .A0(n106), .A1(parser_kimreader_data[55]), .Z(n315));
Q_AN02 U731 ( .A0(n373), .A1(n144), .Z(n316));
Q_MX03 U732 ( .S0(n374), .S1(n375), .A0(n316), .A1(n315), .A2(n314), .Z(kimreader_ckvreader_data[55]));
Q_MX03 U733 ( .S0(n373), .S1(n374), .A0(tlv_word0[56]), .A1(drng_256_out[56]), .A2(drng_256_out[120]), .Z(n317));
Q_INV U734 ( .A(n373), .Z(n318));
Q_AN02 U735 ( .A0(n318), .A1(n107), .Z(n319));
Q_AN02 U736 ( .A0(n373), .A1(n145), .Z(n320));
Q_MX03 U737 ( .S0(n374), .S1(n375), .A0(n320), .A1(n319), .A2(n317), .Z(kimreader_ckvreader_data[56]));
Q_MX03 U738 ( .S0(n373), .S1(n374), .A0(tlv_word0[57]), .A1(drng_256_out[57]), .A2(drng_256_out[121]), .Z(n321));
Q_AN02 U739 ( .A0(n318), .A1(n108), .Z(n322));
Q_AN02 U740 ( .A0(n373), .A1(n146), .Z(n323));
Q_MX03 U741 ( .S0(n374), .S1(n375), .A0(n323), .A1(n322), .A2(n321), .Z(kimreader_ckvreader_data[57]));
Q_MX03 U742 ( .S0(n373), .S1(n374), .A0(tlv_word0[58]), .A1(drng_256_out[58]), .A2(drng_256_out[122]), .Z(n324));
Q_AN02 U743 ( .A0(n318), .A1(n109), .Z(n325));
Q_AN02 U744 ( .A0(n373), .A1(n147), .Z(n326));
Q_MX03 U745 ( .S0(n374), .S1(n375), .A0(n326), .A1(n325), .A2(n324), .Z(kimreader_ckvreader_data[58]));
Q_MX03 U746 ( .S0(n373), .S1(n374), .A0(tlv_word0[59]), .A1(drng_256_out[59]), .A2(drng_256_out[123]), .Z(n327));
Q_AN02 U747 ( .A0(n318), .A1(n110), .Z(n328));
Q_AN02 U748 ( .A0(n373), .A1(n148), .Z(n329));
Q_MX03 U749 ( .S0(n374), .S1(n375), .A0(n329), .A1(n328), .A2(n327), .Z(kimreader_ckvreader_data[59]));
Q_MX03 U750 ( .S0(n373), .S1(n374), .A0(tlv_word0[60]), .A1(drng_256_out[60]), .A2(drng_256_out[124]), .Z(n330));
Q_AN02 U751 ( .A0(n318), .A1(n111), .Z(n331));
Q_AN02 U752 ( .A0(n373), .A1(n149), .Z(n332));
Q_MX03 U753 ( .S0(n374), .S1(n375), .A0(n332), .A1(n331), .A2(n330), .Z(kimreader_ckvreader_data[60]));
Q_MX03 U754 ( .S0(n373), .S1(n374), .A0(tlv_word0[61]), .A1(drng_256_out[61]), .A2(drng_256_out[125]), .Z(n333));
Q_AN02 U755 ( .A0(n318), .A1(n112), .Z(n334));
Q_AN02 U756 ( .A0(n373), .A1(n150), .Z(n335));
Q_MX03 U757 ( .S0(n374), .S1(n375), .A0(n335), .A1(n334), .A2(n333), .Z(kimreader_ckvreader_data[61]));
Q_MX03 U758 ( .S0(n373), .S1(n374), .A0(tlv_word0[62]), .A1(drng_256_out[62]), .A2(drng_256_out[126]), .Z(n336));
Q_AN02 U759 ( .A0(n318), .A1(n113), .Z(n337));
Q_AN02 U760 ( .A0(n373), .A1(n151), .Z(n338));
Q_MX03 U761 ( .S0(n374), .S1(n375), .A0(n338), .A1(n337), .A2(n336), .Z(kimreader_ckvreader_data[62]));
Q_MX03 U762 ( .S0(n373), .S1(n374), .A0(tlv_word0[63]), .A1(drng_256_out[63]), .A2(drng_256_out[127]), .Z(n339));
Q_AN02 U763 ( .A0(n318), .A1(n114), .Z(n340));
Q_AN02 U764 ( .A0(n373), .A1(n152), .Z(n341));
Q_MX03 U765 ( .S0(n374), .S1(n375), .A0(n341), .A1(n340), .A2(n339), .Z(kimreader_ckvreader_data[63]));
Q_AN02 U766 ( .A0(n376), .A1(parser_kimreader_data[64]), .Z(kimreader_ckvreader_data[64]));
Q_AN02 U767 ( .A0(n376), .A1(parser_kimreader_data[65]), .Z(kimreader_ckvreader_data[65]));
Q_AN02 U768 ( .A0(n376), .A1(parser_kimreader_data[66]), .Z(kimreader_ckvreader_data[66]));
Q_AN02 U769 ( .A0(n376), .A1(parser_kimreader_data[67]), .Z(kimreader_ckvreader_data[67]));
Q_AN02 U770 ( .A0(n376), .A1(parser_kimreader_data[68]), .Z(kimreader_ckvreader_data[68]));
Q_AN02 U771 ( .A0(n376), .A1(parser_kimreader_data[69]), .Z(kimreader_ckvreader_data[69]));
Q_AN02 U772 ( .A0(n376), .A1(parser_kimreader_data[70]), .Z(kimreader_ckvreader_data[70]));
Q_MX02 U773 ( .S(n369), .A0(n377), .A1(parser_kimreader_valid), .Z(kimreader_ckvreader_valid));
Q_AN02 U774 ( .A0(n376), .A1(ckvreader_kimreader_ack), .Z(kimreader_parser_ack));
Q_NR02 U775 ( .A0(cur_state[2]), .A1(n343), .Z(n342));
Q_INV U776 ( .A(n344), .Z(n343));
Q_AN02 U777 ( .A0(cur_state[0]), .A1(cur_state[1]), .Z(n344));
Q_NR03 U778 ( .A0(n51), .A1(cur_state[1]), .A2(cur_state[2]), .Z(n345));
Q_NR02 U779 ( .A0(cur_state[2]), .A1(n347), .Z(n346));
Q_OR02 U780 ( .A0(cur_state[0]), .A1(n46), .Z(n347));
Q_INV U781 ( .A(n348), .Z(kim_rd));
Q_OR02 U782 ( .A0(cur_state[2]), .A1(n349), .Z(n348));
Q_XOR2 U783 ( .A0(cur_state[0]), .A1(n46), .Z(n349));
Q_AN03 U784 ( .A0(cur_state[2]), .A1(n350), .A2(ckvreader_kimreader_ack), .Z(drng_ack));
Q_MX02 U785 ( .S(cur_state[2]), .A0(n351), .A1(n350), .Z(n373));
Q_MX02 U786 ( .S(cur_state[0]), .A0(n352), .A1(n354), .Z(n351));
Q_INV U787 ( .A(n353), .Z(n352));
Q_AN02 U788 ( .A0(parser_kimreader_data[69]), .A1(n355), .Z(n354));
Q_AN02 U789 ( .A0(cur_state[0]), .A1(n356), .Z(n350));
Q_INV U790 ( .A(n357), .Z(n374));
Q_MX02 U791 ( .S(cur_state[2]), .A0(n358), .A1(n362), .Z(n357));
Q_MX02 U792 ( .S(cur_state[0]), .A0(n353), .A1(n360), .Z(n358));
Q_OR02 U793 ( .A0(n359), .A1(cur_state[1]), .Z(n353));
Q_INV U794 ( .A(n378), .Z(n359));
Q_OR02 U795 ( .A0(parser_kimreader_data[69]), .A1(n361), .Z(n360));
Q_INV U796 ( .A(n355), .Z(n361));
Q_OR02 U797 ( .A0(cur_state[0]), .A1(n363), .Z(n362));
Q_INV U798 ( .A(n356), .Z(n363));
Q_AN02 U799 ( .A0(parser_kimreader_valid), .A1(drng_valid), .Z(n356));
Q_OR02 U800 ( .A0(n364), .A1(n365), .Z(n375));
Q_NR02 U801 ( .A0(n366), .A1(cur_state[2]), .Z(n365));
Q_OR03 U802 ( .A0(n378), .A1(cur_state[1]), .A2(cur_state[0]), .Z(n366));
Q_AN02 U803 ( .A0(n367), .A1(cur_state[2]), .Z(n364));
Q_AO21 U804 ( .A0(n368), .A1(n53), .B0(n364), .Z(n377));
Q_AN02 U805 ( .A0(cur_state[0]), .A1(n355), .Z(n368));
Q_NR02 U806 ( .A0(cur_state[2]), .A1(n370), .Z(n369));
Q_OR02 U807 ( .A0(cur_state[0]), .A1(cur_state[1]), .Z(n370));
Q_MX02 U808 ( .S(cur_state[2]), .A0(n371), .A1(n367), .Z(n376));
Q_OR02 U809 ( .A0(n368), .A1(n372), .Z(n371));
Q_INV U810 ( .A(n370), .Z(n372));
Q_AN02 U811 ( .A0(cur_state[1]), .A1(n76), .Z(n355));
Q_OA21 U812 ( .A0(drng_valid), .A1(drng_seed_expired), .B0(parser_kimreader_valid), .Z(n367));
Q_FDP1 stat_req_with_expired_seed_REG  ( .CK(clk), .R(rst_n), .D(n379), .Q(stat_req_with_expired_seed), .QN( ));
Q_INV U814 ( .A(parser_kimreader_data[67]), .Z(n380));
Q_AN03 U815 ( .A0(parser_kimreader_data[64]), .A1(n648), .A2(parser_kimreader_data[69]), .Z(n594));
Q_OR03 U816 ( .A0(n383), .A1(tlv_word42[6]), .A2(tlv_word42[5]), .Z(n384));
Q_OR03 U817 ( .A0(tlv_word42[4]), .A1(tlv_word42[3]), .A2(n382), .Z(n385));
Q_OR03 U818 ( .A0(tlv_word42[1]), .A1(n381), .A2(n384), .Z(n386));
Q_OR02 U819 ( .A0(n385), .A1(n386), .Z(n387));
Q_OR03 U820 ( .A0(tlv_word42[4]), .A1(tlv_word42[3]), .A2(tlv_word42[2]), .Z(n389));
Q_OR03 U821 ( .A0(n388), .A1(n381), .A2(n384), .Z(n390));
Q_OR02 U822 ( .A0(n389), .A1(n390), .Z(n391));
Q_AN03 U823 ( .A0(n380), .A1(parser_kimreader_data[66]), .A2(parser_kimreader_data[65]), .Z(n392));
Q_AN03 U824 ( .A0(n37), .A1(n392), .A2(n393), .Z(n571));
Q_OR02 U825 ( .A0(dek_kim_mbe_q), .A1(dak_kim_mbe_q), .Z(n393));
Q_OR03 U826 ( .A0(aux_key_type[5]), .A1(aux_key_type[4]), .A2(aux_key_type[3]), .Z(n394));
Q_OR03 U827 ( .A0(aux_key_type[2]), .A1(aux_key_type[1]), .A2(aux_key_type[0]), .Z(n395));
Q_OA21 U828 ( .A0(n394), .A1(n395), .B0(n76), .Z(n591));
Q_XNR2 U829 ( .A0(tlv_word8[0]), .A1(tlv_word8[27]), .Z(n396));
Q_XNR2 U830 ( .A0(tlv_word8[1]), .A1(tlv_word8[28]), .Z(n397));
Q_XNR2 U831 ( .A0(tlv_word8[2]), .A1(tlv_word8[29]), .Z(n398));
Q_XNR2 U832 ( .A0(tlv_word8[3]), .A1(tlv_word8[30]), .Z(n399));
Q_XNR2 U833 ( .A0(tlv_word8[4]), .A1(tlv_word8[31]), .Z(n400));
Q_XNR2 U834 ( .A0(tlv_word8[5]), .A1(tlv_word8[32]), .Z(n401));
Q_XNR2 U835 ( .A0(tlv_word8[6]), .A1(tlv_word8[33]), .Z(n402));
Q_XNR2 U836 ( .A0(tlv_word8[7]), .A1(tlv_word8[34]), .Z(n403));
Q_XNR2 U837 ( .A0(tlv_word8[8]), .A1(tlv_word8[35]), .Z(n404));
Q_XNR2 U838 ( .A0(tlv_word8[9]), .A1(tlv_word8[36]), .Z(n405));
Q_XNR2 U839 ( .A0(tlv_word8[10]), .A1(tlv_word8[37]), .Z(n406));
Q_XNR2 U840 ( .A0(tlv_word8[11]), .A1(tlv_word8[38]), .Z(n407));
Q_AN03 U841 ( .A0(n407), .A1(n406), .A2(n405), .Z(n408));
Q_AN03 U842 ( .A0(n404), .A1(n403), .A2(n402), .Z(n409));
Q_AN03 U843 ( .A0(n401), .A1(n400), .A2(n399), .Z(n410));
Q_AN03 U844 ( .A0(n398), .A1(n397), .A2(n396), .Z(n411));
Q_AN03 U845 ( .A0(n408), .A1(n409), .A2(n410), .Z(n412));
Q_ND02 U846 ( .A0(n411), .A1(n412), .Z(n413));
Q_AN02 U847 ( .A0(tlv_word8[16]), .A1(n413), .Z(n592));
Q_XNR2 U848 ( .A0(tlv_word8[16]), .A1(tlv_word8[26]), .Z(n414));
Q_INV U849 ( .A(n414), .Z(n595));
Q_XNR2 U850 ( .A0(tlv_word8[12]), .A1(tlv_word8[39]), .Z(n415));
Q_INV U851 ( .A(n415), .Z(n596));
Q_XNR2 U852 ( .A0(tlv_word8[0]), .A1(tlv_word9[27]), .Z(n416));
Q_XNR2 U853 ( .A0(tlv_word8[1]), .A1(tlv_word9[28]), .Z(n417));
Q_XNR2 U854 ( .A0(tlv_word8[2]), .A1(tlv_word9[29]), .Z(n418));
Q_XNR2 U855 ( .A0(tlv_word8[3]), .A1(tlv_word9[30]), .Z(n419));
Q_XNR2 U856 ( .A0(tlv_word8[4]), .A1(tlv_word9[31]), .Z(n420));
Q_XNR2 U857 ( .A0(tlv_word8[5]), .A1(tlv_word9[32]), .Z(n421));
Q_XNR2 U858 ( .A0(tlv_word8[6]), .A1(tlv_word9[33]), .Z(n422));
Q_XNR2 U859 ( .A0(tlv_word8[7]), .A1(tlv_word9[34]), .Z(n423));
Q_XNR2 U860 ( .A0(tlv_word8[8]), .A1(tlv_word9[35]), .Z(n424));
Q_XNR2 U861 ( .A0(tlv_word8[9]), .A1(tlv_word9[36]), .Z(n425));
Q_XNR2 U862 ( .A0(tlv_word8[10]), .A1(tlv_word9[37]), .Z(n426));
Q_XNR2 U863 ( .A0(tlv_word8[11]), .A1(tlv_word9[38]), .Z(n427));
Q_AN03 U864 ( .A0(n427), .A1(n426), .A2(n425), .Z(n428));
Q_AN03 U865 ( .A0(n424), .A1(n423), .A2(n422), .Z(n429));
Q_AN03 U866 ( .A0(n421), .A1(n420), .A2(n419), .Z(n430));
Q_AN03 U867 ( .A0(n418), .A1(n417), .A2(n416), .Z(n431));
Q_AN03 U868 ( .A0(n428), .A1(n429), .A2(n430), .Z(n432));
Q_ND02 U869 ( .A0(n431), .A1(n432), .Z(n433));
Q_AN02 U870 ( .A0(tlv_word8[16]), .A1(n433), .Z(n593));
Q_XNR2 U871 ( .A0(tlv_word8[16]), .A1(tlv_word9[26]), .Z(n434));
Q_INV U872 ( .A(n434), .Z(n597));
Q_XNR2 U873 ( .A0(tlv_word8[12]), .A1(tlv_word9[39]), .Z(n435));
Q_INV U874 ( .A(n435), .Z(n598));
Q_AO21 U875 ( .A0(n469), .A1(n437), .B0(n571), .Z(n436));
Q_OR02 U876 ( .A0(n569), .A1(n570), .Z(n437));
Q_XOR2 U877 ( .A0(n469), .A1(n442), .Z(n439));
Q_NR02 U878 ( .A0(n571), .A1(n441), .Z(n440));
Q_MX02 U879 ( .S(n469), .A0(n443), .A1(n438), .Z(n441));
Q_INV U880 ( .A(n442), .Z(n438));
Q_XOR2 U881 ( .A0(n453), .A1(n570), .Z(n442));
Q_ND02 U882 ( .A0(n453), .A1(n570), .Z(n443));
Q_MX02 U883 ( .S(n469), .A0(n445), .A1(n453), .Z(n444));
Q_AN02 U884 ( .A0(n569), .A1(n570), .Z(n445));
Q_OR03 U885 ( .A0(n453), .A1(n570), .A2(n469), .Z(n446));
Q_FDP1 stat_aux_key_type_0_REG  ( .CK(clk), .R(rst_n), .D(n586), .Q(stat_aux_key_type_0), .QN( ));
Q_FDP1 stat_aux_key_type_1_REG  ( .CK(clk), .R(rst_n), .D(n585), .Q(stat_aux_key_type_1), .QN( ));
Q_FDP1 stat_aux_key_type_2_REG  ( .CK(clk), .R(rst_n), .D(n584), .Q(stat_aux_key_type_2), .QN( ));
Q_FDP1 stat_aux_key_type_3_REG  ( .CK(clk), .R(rst_n), .D(n583), .Q(stat_aux_key_type_3), .QN( ));
Q_FDP1 stat_aux_key_type_4_REG  ( .CK(clk), .R(rst_n), .D(n582), .Q(stat_aux_key_type_4), .QN( ));
Q_FDP1 stat_aux_key_type_5_REG  ( .CK(clk), .R(rst_n), .D(n581), .Q(stat_aux_key_type_5), .QN( ));
Q_FDP1 stat_aux_key_type_6_REG  ( .CK(clk), .R(rst_n), .D(n580), .Q(stat_aux_key_type_6), .QN( ));
Q_FDP1 stat_aux_key_type_7_REG  ( .CK(clk), .R(rst_n), .D(n579), .Q(stat_aux_key_type_7), .QN( ));
Q_FDP1 stat_aux_key_type_8_REG  ( .CK(clk), .R(rst_n), .D(n578), .Q(stat_aux_key_type_8), .QN( ));
Q_FDP1 stat_aux_key_type_9_REG  ( .CK(clk), .R(rst_n), .D(n577), .Q(stat_aux_key_type_9), .QN( ));
Q_FDP1 stat_aux_key_type_10_REG  ( .CK(clk), .R(rst_n), .D(n576), .Q(stat_aux_key_type_10), .QN( ));
Q_FDP1 stat_aux_key_type_11_REG  ( .CK(clk), .R(rst_n), .D(n575), .Q(stat_aux_key_type_11), .QN( ));
Q_FDP1 stat_aux_key_type_12_REG  ( .CK(clk), .R(rst_n), .D(n574), .Q(stat_aux_key_type_12), .QN( ));
Q_FDP1 stat_aux_key_type_13_REG  ( .CK(clk), .R(rst_n), .D(n573), .Q(stat_aux_key_type_13), .QN( ));
Q_FDP1 stat_aux_cmd_with_vf_pf_fail_REG  ( .CK(clk), .R(rst_n), .D(n572), .Q(stat_aux_cmd_with_vf_pf_fail), .QN( ));
Q_AN02 U901 ( .A0(rst_n), .A1(n589), .Z(n447));
Q_AN02 U902 ( .A0(rst_n), .A1(n590), .Z(n448));
Q_INV U903 ( .A(n451), .Z(n567));
Q_INV U904 ( .A(n452), .Z(n568));
Q_INV U905 ( .A(n453), .Z(n569));
Q_AO21 U906 ( .A0(n455), .A1(n456), .B0(n454), .Z(n453));
Q_AN02 U907 ( .A0(n457), .A1(n458), .Z(n456));
Q_AO21 U908 ( .A0(n460), .A1(n461), .B0(n459), .Z(n454));
Q_AN03 U909 ( .A0(n463), .A1(n458), .A2(n462), .Z(n461));
Q_AO21 U910 ( .A0(n463), .A1(n464), .B0(n571), .Z(n459));
Q_NR02 U911 ( .A0(tlv_word8[63]), .A1(n571), .Z(n464));
Q_INV U912 ( .A(tlv_word9[63]), .Z(n466));
Q_AO21 U913 ( .A0(n467), .A1(n468), .B0(n466), .Z(n455));
Q_AN03 U914 ( .A0(tlv_word9[63]), .A1(n458), .A2(n457), .Z(n471));
Q_OR02 U915 ( .A0(n472), .A1(n571), .Z(n470));
Q_AO21 U916 ( .A0(n473), .A1(n474), .B0(n470), .Z(n469));
Q_AN03 U917 ( .A0(tlv_word8[63]), .A1(n458), .A2(n463), .Z(n474));
Q_OA21 U918 ( .A0(n475), .A1(n476), .B0(n471), .Z(n472));
Q_NR02 U919 ( .A0(n477), .A1(n476), .Z(n475));
Q_OR03 U920 ( .A0(n593), .A1(n598), .A2(n597), .Z(n476));
Q_INV U921 ( .A(n477), .Z(n467));
Q_OA21 U922 ( .A0(n478), .A1(n479), .B0(n458), .Z(n570));
Q_AN03 U923 ( .A0(n463), .A1(tlv_word8[63]), .A2(n473), .Z(n480));
Q_AO21 U924 ( .A0(n463), .A1(n465), .B0(n481), .Z(n484));
Q_INV U925 ( .A(tlv_word8[63]), .Z(n465));
Q_AN03 U926 ( .A0(n483), .A1(tlv_word9[17]), .A2(n482), .Z(n463));
Q_AN03 U927 ( .A0(n486), .A1(n487), .A2(disable_unencrypted_keys), .Z(n485));
Q_AN02 U928 ( .A0(n488), .A1(parser_kimreader_data[41]), .Z(n487));
Q_AN03 U929 ( .A0(n490), .A1(n489), .A2(n485), .Z(n479));
Q_ND02 U930 ( .A0(parser_kimreader_data[40]), .A1(parser_kimreader_data[39]), .Z(n489));
Q_AN03 U931 ( .A0(n492), .A1(n493), .A2(n490), .Z(n491));
Q_AN02 U932 ( .A0(parser_kimreader_data[40]), .A1(disable_unencrypted_keys), .Z(n493));
Q_AO21 U933 ( .A0(n495), .A1(n496), .B0(n494), .Z(n490));
Q_OR03 U934 ( .A0(n497), .A1(n498), .A2(n491), .Z(n478));
Q_AN03 U935 ( .A0(n500), .A1(n496), .A2(n495), .Z(n499));
Q_OR02 U936 ( .A0(n484), .A1(n499), .Z(n497));
Q_AN02 U937 ( .A0(n494), .A1(n500), .Z(n498));
Q_AN03 U938 ( .A0(n501), .A1(n502), .A2(n492), .Z(n500));
Q_INV U939 ( .A(parser_kimreader_data[47]), .Z(n502));
Q_NR02 U940 ( .A0(parser_kimreader_data[40]), .A1(parser_kimreader_data[39]), .Z(n501));
Q_AN02 U941 ( .A0(n486), .A1(n503), .Z(n492));
Q_NR02 U942 ( .A0(parser_kimreader_data[42]), .A1(parser_kimreader_data[41]), .Z(n503));
Q_INV U943 ( .A(parser_kimreader_data[42]), .Z(n488));
Q_NR02 U944 ( .A0(parser_kimreader_data[44]), .A1(parser_kimreader_data[43]), .Z(n486));
Q_AO21 U945 ( .A0(n504), .A1(n483), .B0(n480), .Z(n481));
Q_AO21 U946 ( .A0(n506), .A1(parser_kimreader_data[69]), .B0(n505), .Z(n494));
Q_INV U947 ( .A(n482), .Z(n504));
Q_OR02 U948 ( .A0(n507), .A1(n508), .Z(n473));
Q_NR02 U949 ( .A0(n509), .A1(n508), .Z(n507));
Q_OR03 U950 ( .A0(n592), .A1(n596), .A2(n595), .Z(n508));
Q_INV U951 ( .A(n509), .Z(n460));
Q_AN02 U952 ( .A0(n510), .A1(n511), .Z(n572));
Q_AN02 U953 ( .A0(kimreader_parser_ack), .A1(n594), .Z(n510));
Q_ND02 U954 ( .A0(n391), .A1(n387), .Z(n511));
Q_AN02 U955 ( .A0(n512), .A1(n513), .Z(n573));
Q_AN02 U956 ( .A0(n514), .A1(n510), .Z(n513));
Q_AN02 U957 ( .A0(n512), .A1(n515), .Z(n574));
Q_AN02 U958 ( .A0(n516), .A1(n510), .Z(n515));
Q_AN02 U959 ( .A0(n517), .A1(n518), .Z(n512));
Q_AN02 U960 ( .A0(n519), .A1(n520), .Z(n575));
Q_AN02 U961 ( .A0(n521), .A1(n510), .Z(n520));
Q_AN02 U962 ( .A0(n519), .A1(n522), .Z(n576));
Q_AN02 U963 ( .A0(n519), .A1(n513), .Z(n577));
Q_AN02 U964 ( .A0(n519), .A1(n515), .Z(n578));
Q_AN03 U965 ( .A0(aux_key_type[3]), .A1(n523), .A2(n517), .Z(n519));
Q_AN02 U966 ( .A0(n524), .A1(n520), .Z(n579));
Q_AN02 U967 ( .A0(n524), .A1(n522), .Z(n580));
Q_AN02 U968 ( .A0(n524), .A1(n513), .Z(n581));
Q_AN02 U969 ( .A0(n524), .A1(n515), .Z(n582));
Q_AN02 U970 ( .A0(n517), .A1(n525), .Z(n524));
Q_AN02 U971 ( .A0(n526), .A1(n520), .Z(n583));
Q_AN02 U972 ( .A0(n526), .A1(n522), .Z(n584));
Q_AN03 U973 ( .A0(aux_key_type[1]), .A1(n527), .A2(n510), .Z(n522));
Q_AN02 U974 ( .A0(n526), .A1(n513), .Z(n585));
Q_INV U975 ( .A(n528), .Z(n514));
Q_AN02 U976 ( .A0(n526), .A1(n515), .Z(n586));
Q_AN02 U977 ( .A0(n517), .A1(n529), .Z(n526));
Q_NR02 U978 ( .A0(aux_key_type[3]), .A1(aux_key_type[2]), .Z(n529));
Q_AN02 U979 ( .A0(kimreader_parser_ack), .A1(n38), .Z(n587));
Q_AN03 U980 ( .A0(n534), .A1(n458), .A2(n506), .Z(n533));
Q_AN02 U981 ( .A0(n3), .A1(parser_kimreader_data[69]), .Z(n534));
Q_AO21 U982 ( .A0(n477), .A1(n468), .B0(n535), .Z(n506));
Q_AN03 U983 ( .A0(tlv_word9[63]), .A1(n435), .A2(n536), .Z(n468));
Q_AN02 U984 ( .A0(n537), .A1(n434), .Z(n536));
Q_INV U985 ( .A(n593), .Z(n537));
Q_INV U986 ( .A(tlv_word9[17]), .Z(n535));
Q_AN02 U987 ( .A0(n452), .A1(n539), .Z(n538));
Q_AO21 U988 ( .A0(n540), .A1(n541), .B0(n538), .Z(n477));
Q_AN02 U989 ( .A0(n542), .A1(tlv_word9[42]), .Z(n541));
Q_INV U990 ( .A(n543), .Z(n542));
Q_OR02 U991 ( .A0(n543), .A1(n544), .Z(n452));
Q_ND02 U992 ( .A0(n517), .A1(aux_key_type[3]), .Z(n543));
Q_INV U993 ( .A(n540), .Z(n544));
Q_INV U994 ( .A(n545), .Z(n516));
Q_AO21 U995 ( .A0(n545), .A1(n523), .B0(n546), .Z(n540));
Q_OR02 U996 ( .A0(aux_key_type[0]), .A1(aux_key_type[1]), .Z(n545));
Q_OR03 U997 ( .A0(n48), .A1(n533), .A2(n532), .Z(n531));
Q_AN02 U998 ( .A0(n3), .A1(n458), .Z(n547));
Q_INV U999 ( .A(n571), .Z(n458));
Q_OA21 U1000 ( .A0(n505), .A1(n548), .B0(n547), .Z(n532));
Q_AN03 U1001 ( .A0(n496), .A1(n482), .A2(n495), .Z(n548));
Q_INV U1002 ( .A(n591), .Z(n505));
Q_AO21 U1003 ( .A0(n509), .A1(n462), .B0(n535), .Z(n495));
Q_AN02 U1004 ( .A0(n414), .A1(n415), .Z(n549));
Q_AN03 U1005 ( .A0(tlv_word8[63]), .A1(n550), .A2(n549), .Z(n462));
Q_INV U1006 ( .A(n592), .Z(n550));
Q_AN02 U1007 ( .A0(tlv_word8[42]), .A1(n517), .Z(n552));
Q_NR02 U1008 ( .A0(aux_key_type[5]), .A1(aux_key_type[4]), .Z(n517));
Q_AO21 U1009 ( .A0(n451), .A1(n553), .B0(n551), .Z(n509));
Q_OA21 U1010 ( .A0(n554), .A1(n555), .B0(n552), .Z(n551));
Q_AN02 U1011 ( .A0(n525), .A1(n521), .Z(n554));
Q_AN02 U1012 ( .A0(aux_key_type[1]), .A1(aux_key_type[0]), .Z(n521));
Q_AN02 U1013 ( .A0(n530), .A1(aux_key_type[2]), .Z(n525));
Q_OA21 U1014 ( .A0(n556), .A1(n546), .B0(aux_key_type[3]), .Z(n555));
Q_AN02 U1015 ( .A0(aux_key_type[2]), .A1(n557), .Z(n546));
Q_AN02 U1016 ( .A0(n528), .A1(n523), .Z(n556));
Q_OR02 U1017 ( .A0(n527), .A1(aux_key_type[1]), .Z(n528));
Q_AO21 U1018 ( .A0(n518), .A1(aux_key_type[1]), .B0(aux_key_type[5]), .Z(n559));
Q_AN02 U1019 ( .A0(aux_key_type[3]), .A1(aux_key_type[2]), .Z(n518));
Q_OR03 U1020 ( .A0(n560), .A1(n559), .A2(n558), .Z(n451));
Q_AO21 U1021 ( .A0(n561), .A1(n557), .B0(aux_key_type[4]), .Z(n558));
Q_AN02 U1022 ( .A0(n562), .A1(n530), .Z(n560));
Q_AO21 U1023 ( .A0(n523), .A1(aux_key_type[0]), .B0(n530), .Z(n561));
Q_ND02 U1024 ( .A0(aux_key_type[2]), .A1(aux_key_type[0]), .Z(n562));
Q_AN02 U1025 ( .A0(kimreader_parser_ack), .A1(n4), .Z(n588));
Q_AN02 U1026 ( .A0(kimreader_parser_ack), .A1(n483), .Z(n563));
Q_AN03 U1027 ( .A0(n482), .A1(n564), .A2(n563), .Z(n589));
Q_AN02 U1028 ( .A0(tlv_word9[17]), .A1(tlv_word8[42]), .Z(n564));
Q_AN03 U1029 ( .A0(n482), .A1(n565), .A2(n563), .Z(n590));
Q_AN02 U1030 ( .A0(tlv_word9[17]), .A1(n553), .Z(n565));
Q_INV U1031 ( .A(tlv_word8[42]), .Z(n553));
Q_NR02 U1032 ( .A0(tlv_word9[18]), .A1(tlv_word9[19]), .Z(n482));
Q_AN02 U1033 ( .A0(n591), .A1(n496), .Z(n483));
Q_INV U1034 ( .A(parser_kimreader_data[69]), .Z(n496));
Q_AN03 U1035 ( .A0(n566), .A1(tlv_word9[42]), .A2(rst_n), .Z(n449));
Q_AN03 U1036 ( .A0(n566), .A1(n539), .A2(rst_n), .Z(n450));
Q_INV U1037 ( .A(tlv_word9[42]), .Z(n539));
Q_AN02 U1038 ( .A0(kimreader_parser_ack), .A1(n457), .Z(n566));
Q_AN03 U1039 ( .A0(parser_kimreader_data[69]), .A1(tlv_word9[17]), .A2(n591), .Z(n457));
Q_AN03 U1040 ( .A0(kimreader_ckvreader_data[67]), .A1(kimreader_ckvreader_data[66]), .A2(kimreader_ckvreader_data[65]), .Z(n599));
Q_AN02 U1041 ( .A0(kimreader_ckvreader_data[64]), .A1(n599), .Z(n600));
Q_AN03 U1042 ( .A0(kimreader_ckvreader_valid), .A1(n600), .A2(ckvreader_kimreader_ack), .Z(n645));
Q_AN02 U1043 ( .A0(kim_rd_q), .A1(kim_mbe), .Z(n601));
Q_AN02 U1044 ( .A0(kim_rd_q), .A1(kim_dout[0]), .Z(n602));
Q_AN02 U1045 ( .A0(kim_rd_q), .A1(kim_dout[1]), .Z(n603));
Q_AN02 U1046 ( .A0(kim_rd_q), .A1(kim_dout[2]), .Z(n604));
Q_AN02 U1047 ( .A0(kim_rd_q), .A1(kim_dout[3]), .Z(n605));
Q_AN02 U1048 ( .A0(kim_rd_q), .A1(kim_dout[4]), .Z(n606));
Q_AN02 U1049 ( .A0(kim_rd_q), .A1(kim_dout[5]), .Z(n607));
Q_AN02 U1050 ( .A0(kim_rd_q), .A1(kim_dout[6]), .Z(n608));
Q_AN02 U1051 ( .A0(kim_rd_q), .A1(kim_dout[7]), .Z(n609));
Q_AN02 U1052 ( .A0(kim_rd_q), .A1(kim_dout[8]), .Z(n610));
Q_AN02 U1053 ( .A0(kim_rd_q), .A1(kim_dout[9]), .Z(n611));
Q_AN02 U1054 ( .A0(kim_rd_q), .A1(kim_dout[10]), .Z(n612));
Q_AN02 U1055 ( .A0(kim_rd_q), .A1(kim_dout[11]), .Z(n613));
Q_AN02 U1056 ( .A0(kim_rd_q), .A1(kim_dout[12]), .Z(n614));
Q_AN02 U1057 ( .A0(kim_rd_q), .A1(kim_dout[13]), .Z(n615));
Q_AN02 U1058 ( .A0(kim_rd_q), .A1(kim_dout[14]), .Z(n616));
Q_AN02 U1059 ( .A0(kim_rd_q), .A1(kim_dout[15]), .Z(n617));
Q_AN02 U1060 ( .A0(kim_rd_q), .A1(kim_dout[16]), .Z(n618));
Q_AN02 U1061 ( .A0(kim_rd_q), .A1(kim_dout[17]), .Z(n619));
Q_AN02 U1062 ( .A0(kim_rd_q), .A1(kim_dout[18]), .Z(n620));
Q_AN02 U1063 ( .A0(kim_rd_q), .A1(kim_dout[19]), .Z(n621));
Q_AN02 U1064 ( .A0(kim_rd_q), .A1(kim_dout[20]), .Z(n622));
Q_AN02 U1065 ( .A0(kim_rd_q), .A1(kim_dout[21]), .Z(n623));
Q_AN02 U1066 ( .A0(kim_rd_q), .A1(kim_dout[22]), .Z(n624));
Q_AN02 U1067 ( .A0(kim_rd_q), .A1(kim_dout[23]), .Z(n625));
Q_AN02 U1068 ( .A0(kim_rd_q), .A1(kim_dout[24]), .Z(n626));
Q_AN02 U1069 ( .A0(kim_rd_q), .A1(kim_dout[25]), .Z(n627));
Q_AN02 U1070 ( .A0(kim_rd_q), .A1(kim_dout[26]), .Z(n628));
Q_AN02 U1071 ( .A0(kim_rd_q), .A1(kim_dout[27]), .Z(n629));
Q_AN02 U1072 ( .A0(kim_rd_q), .A1(kim_dout[28]), .Z(n630));
Q_AN02 U1073 ( .A0(kim_rd_q), .A1(kim_dout[29]), .Z(n631));
Q_AN02 U1074 ( .A0(kim_rd_q), .A1(kim_dout[30]), .Z(n632));
Q_AN02 U1075 ( .A0(kim_rd_q), .A1(kim_dout[31]), .Z(n633));
Q_AN02 U1076 ( .A0(kim_rd_q), .A1(kim_dout[32]), .Z(n634));
Q_AN02 U1077 ( .A0(kim_rd_q), .A1(kim_dout[33]), .Z(n635));
Q_AN02 U1078 ( .A0(kim_rd_q), .A1(kim_dout[34]), .Z(n636));
Q_AN02 U1079 ( .A0(kim_rd_q), .A1(kim_dout[35]), .Z(n637));
Q_AN02 U1080 ( .A0(kim_rd_q), .A1(kim_dout[36]), .Z(n638));
Q_AN02 U1081 ( .A0(kim_rd_q), .A1(kim_dout[37]), .Z(n639));
Q_AO21 U1082 ( .A0(n641), .A1(n647), .B0(n640), .Z(n643));
Q_AO21 U1083 ( .A0(n641), .A1(n344), .B0(n640), .Z(n644));
Q_AN02 U1084 ( .A0(kim_rd_q), .A1(n53), .Z(n641));
Q_AN02 U1085 ( .A0(n642), .A1(n645), .Z(n640));
Q_INV U1086 ( .A(n347), .Z(n647));
Q_INV U1087 ( .A(n75), .Z(n648));
Q_FDP4EP dak_kim_mbe_q_REG  ( .CK(clk), .CE(n644), .R(n649), .D(n601), .Q(dak_kim_mbe_q));
Q_INV U1089 ( .A(rst_n), .Z(n649));
Q_FDP4EP dek_kim_mbe_q_REG  ( .CK(clk), .CE(n643), .R(n649), .D(n601), .Q(dek_kim_mbe_q));
Q_FDP4EP \dak_kim_entry_q_REG[0] ( .CK(clk), .CE(n644), .R(n649), .D(n602), .Q(dak_kim_entry_q[0]));
Q_FDP4EP \dak_kim_entry_q_REG[1] ( .CK(clk), .CE(n644), .R(n649), .D(n603), .Q(dak_kim_entry_q[1]));
Q_FDP4EP \dak_kim_entry_q_REG[2] ( .CK(clk), .CE(n644), .R(n649), .D(n604), .Q(dak_kim_entry_q[2]));
Q_FDP4EP \dak_kim_entry_q_REG[3] ( .CK(clk), .CE(n644), .R(n649), .D(n605), .Q(dak_kim_entry_q[3]));
Q_FDP4EP \dak_kim_entry_q_REG[4] ( .CK(clk), .CE(n644), .R(n649), .D(n606), .Q(dak_kim_entry_q[4]));
Q_FDP4EP \dak_kim_entry_q_REG[5] ( .CK(clk), .CE(n644), .R(n649), .D(n607), .Q(dak_kim_entry_q[5]));
Q_FDP4EP \dak_kim_entry_q_REG[6] ( .CK(clk), .CE(n644), .R(n649), .D(n608), .Q(dak_kim_entry_q[6]));
Q_FDP4EP \dak_kim_entry_q_REG[7] ( .CK(clk), .CE(n644), .R(n649), .D(n609), .Q(dak_kim_entry_q[7]));
Q_FDP4EP \dak_kim_entry_q_REG[8] ( .CK(clk), .CE(n644), .R(n649), .D(n610), .Q(dak_kim_entry_q[8]));
Q_FDP4EP \dak_kim_entry_q_REG[9] ( .CK(clk), .CE(n644), .R(n649), .D(n611), .Q(dak_kim_entry_q[9]));
Q_FDP4EP \dak_kim_entry_q_REG[10] ( .CK(clk), .CE(n644), .R(n649), .D(n612), .Q(dak_kim_entry_q[10]));
Q_FDP4EP \dak_kim_entry_q_REG[11] ( .CK(clk), .CE(n644), .R(n649), .D(n613), .Q(dak_kim_entry_q[11]));
Q_FDP4EP \dak_kim_entry_q_REG[12] ( .CK(clk), .CE(n644), .R(n649), .D(n614), .Q(dak_kim_entry_q[12]));
Q_FDP4EP \dak_kim_entry_q_REG[13] ( .CK(clk), .CE(n644), .R(n649), .D(n615), .Q(dak_kim_entry_q[13]));
Q_FDP4EP \dak_kim_entry_q_REG[14] ( .CK(clk), .CE(n644), .R(n649), .D(n616), .Q(dak_kim_entry_q[14]));
Q_FDP4EP \dak_kim_entry_q_REG[15] ( .CK(clk), .CE(n644), .R(n649), .D(n617), .Q(dak_kim_entry_q[15]));
Q_FDP4EP \dak_kim_entry_q_REG[16] ( .CK(clk), .CE(n644), .R(n649), .D(n618), .Q(dak_kim_entry_q[16]));
Q_FDP4EP \dak_kim_entry_q_REG[17] ( .CK(clk), .CE(n644), .R(n649), .D(n619), .Q(dak_kim_entry_q[17]));
Q_FDP4EP \dak_kim_entry_q_REG[18] ( .CK(clk), .CE(n644), .R(n649), .D(n620), .Q(dak_kim_entry_q[18]));
Q_FDP4EP \dak_kim_entry_q_REG[19] ( .CK(clk), .CE(n644), .R(n649), .D(n621), .Q(dak_kim_entry_q[19]));
Q_FDP4EP \dak_kim_entry_q_REG[20] ( .CK(clk), .CE(n644), .R(n649), .D(n622), .Q(dak_kim_entry_q[20]));
Q_FDP4EP \dak_kim_entry_q_REG[21] ( .CK(clk), .CE(n644), .R(n649), .D(n623), .Q(dak_kim_entry_q[21]));
Q_FDP4EP \dak_kim_entry_q_REG[22] ( .CK(clk), .CE(n644), .R(n649), .D(n624), .Q(dak_kim_entry_q[22]));
Q_FDP4EP \dak_kim_entry_q_REG[23] ( .CK(clk), .CE(n644), .R(n649), .D(n625), .Q(dak_kim_entry_q[23]));
Q_FDP4EP \dak_kim_entry_q_REG[24] ( .CK(clk), .CE(n644), .R(n649), .D(n626), .Q(dak_kim_entry_q[24]));
Q_FDP4EP \dak_kim_entry_q_REG[25] ( .CK(clk), .CE(n644), .R(n649), .D(n627), .Q(dak_kim_entry_q[25]));
Q_FDP4EP \dak_kim_entry_q_REG[26] ( .CK(clk), .CE(n644), .R(n649), .D(n628), .Q(dak_kim_entry_q[26]));
Q_FDP4EP \dak_kim_entry_q_REG[27] ( .CK(clk), .CE(n644), .R(n649), .D(n629), .Q(dak_kim_entry_q[27]));
Q_FDP4EP \dak_kim_entry_q_REG[28] ( .CK(clk), .CE(n644), .R(n649), .D(n630), .Q(dak_kim_entry_q[28]));
Q_FDP4EP \dak_kim_entry_q_REG[29] ( .CK(clk), .CE(n644), .R(n649), .D(n631), .Q(dak_kim_entry_q[29]));
Q_FDP4EP \dak_kim_entry_q_REG[30] ( .CK(clk), .CE(n644), .R(n649), .D(n632), .Q(dak_kim_entry_q[30]));
Q_FDP4EP \dak_kim_entry_q_REG[31] ( .CK(clk), .CE(n644), .R(n649), .D(n633), .Q(dak_kim_entry_q[31]));
Q_FDP4EP \dak_kim_entry_q_REG[32] ( .CK(clk), .CE(n644), .R(n649), .D(n634), .Q(dak_kim_entry_q[32]));
Q_FDP4EP \dak_kim_entry_q_REG[33] ( .CK(clk), .CE(n644), .R(n649), .D(n635), .Q(dak_kim_entry_q[33]));
Q_FDP4EP \dak_kim_entry_q_REG[34] ( .CK(clk), .CE(n644), .R(n649), .D(n636), .Q(dak_kim_entry_q[34]));
Q_FDP4EP \dak_kim_entry_q_REG[35] ( .CK(clk), .CE(n644), .R(n649), .D(n637), .Q(dak_kim_entry_q[35]));
Q_FDP4EP \dak_kim_entry_q_REG[36] ( .CK(clk), .CE(n644), .R(n649), .D(n638), .Q(dak_kim_entry_q[36]));
Q_FDP4EP \dak_kim_entry_q_REG[37] ( .CK(clk), .CE(n644), .R(n649), .D(n639), .Q(dak_kim_entry_q[37]));
Q_FDP4EP \dek_kim_entry_q_REG[0] ( .CK(clk), .CE(n643), .R(n649), .D(n602), .Q(dek_kim_entry_q[0]));
Q_FDP4EP \dek_kim_entry_q_REG[1] ( .CK(clk), .CE(n643), .R(n649), .D(n603), .Q(dek_kim_entry_q[1]));
Q_FDP4EP \dek_kim_entry_q_REG[2] ( .CK(clk), .CE(n643), .R(n649), .D(n604), .Q(dek_kim_entry_q[2]));
Q_FDP4EP \dek_kim_entry_q_REG[3] ( .CK(clk), .CE(n643), .R(n649), .D(n605), .Q(dek_kim_entry_q[3]));
Q_FDP4EP \dek_kim_entry_q_REG[4] ( .CK(clk), .CE(n643), .R(n649), .D(n606), .Q(dek_kim_entry_q[4]));
Q_FDP4EP \dek_kim_entry_q_REG[5] ( .CK(clk), .CE(n643), .R(n649), .D(n607), .Q(dek_kim_entry_q[5]));
Q_FDP4EP \dek_kim_entry_q_REG[6] ( .CK(clk), .CE(n643), .R(n649), .D(n608), .Q(dek_kim_entry_q[6]));
Q_FDP4EP \dek_kim_entry_q_REG[7] ( .CK(clk), .CE(n643), .R(n649), .D(n609), .Q(dek_kim_entry_q[7]));
Q_FDP4EP \dek_kim_entry_q_REG[8] ( .CK(clk), .CE(n643), .R(n649), .D(n610), .Q(dek_kim_entry_q[8]));
Q_FDP4EP \dek_kim_entry_q_REG[9] ( .CK(clk), .CE(n643), .R(n649), .D(n611), .Q(dek_kim_entry_q[9]));
Q_FDP4EP \dek_kim_entry_q_REG[10] ( .CK(clk), .CE(n643), .R(n649), .D(n612), .Q(dek_kim_entry_q[10]));
Q_FDP4EP \dek_kim_entry_q_REG[11] ( .CK(clk), .CE(n643), .R(n649), .D(n613), .Q(dek_kim_entry_q[11]));
Q_FDP4EP \dek_kim_entry_q_REG[12] ( .CK(clk), .CE(n643), .R(n649), .D(n614), .Q(dek_kim_entry_q[12]));
Q_FDP4EP \dek_kim_entry_q_REG[13] ( .CK(clk), .CE(n643), .R(n649), .D(n615), .Q(dek_kim_entry_q[13]));
Q_FDP4EP \dek_kim_entry_q_REG[14] ( .CK(clk), .CE(n643), .R(n649), .D(n616), .Q(dek_kim_entry_q[14]));
Q_FDP4EP \dek_kim_entry_q_REG[15] ( .CK(clk), .CE(n643), .R(n649), .D(n617), .Q(dek_kim_entry_q[15]));
Q_FDP4EP \dek_kim_entry_q_REG[16] ( .CK(clk), .CE(n643), .R(n649), .D(n618), .Q(dek_kim_entry_q[16]));
Q_FDP4EP \dek_kim_entry_q_REG[17] ( .CK(clk), .CE(n643), .R(n649), .D(n619), .Q(dek_kim_entry_q[17]));
Q_FDP4EP \dek_kim_entry_q_REG[18] ( .CK(clk), .CE(n643), .R(n649), .D(n620), .Q(dek_kim_entry_q[18]));
Q_FDP4EP \dek_kim_entry_q_REG[19] ( .CK(clk), .CE(n643), .R(n649), .D(n621), .Q(dek_kim_entry_q[19]));
Q_FDP4EP \dek_kim_entry_q_REG[20] ( .CK(clk), .CE(n643), .R(n649), .D(n622), .Q(dek_kim_entry_q[20]));
Q_FDP4EP \dek_kim_entry_q_REG[21] ( .CK(clk), .CE(n643), .R(n649), .D(n623), .Q(dek_kim_entry_q[21]));
Q_FDP4EP \dek_kim_entry_q_REG[22] ( .CK(clk), .CE(n643), .R(n649), .D(n624), .Q(dek_kim_entry_q[22]));
Q_FDP4EP \dek_kim_entry_q_REG[23] ( .CK(clk), .CE(n643), .R(n649), .D(n625), .Q(dek_kim_entry_q[23]));
Q_FDP4EP \dek_kim_entry_q_REG[24] ( .CK(clk), .CE(n643), .R(n649), .D(n626), .Q(dek_kim_entry_q[24]));
Q_FDP4EP \dek_kim_entry_q_REG[25] ( .CK(clk), .CE(n643), .R(n649), .D(n627), .Q(dek_kim_entry_q[25]));
Q_FDP4EP \dek_kim_entry_q_REG[26] ( .CK(clk), .CE(n643), .R(n649), .D(n628), .Q(dek_kim_entry_q[26]));
Q_FDP4EP \dek_kim_entry_q_REG[27] ( .CK(clk), .CE(n643), .R(n649), .D(n629), .Q(dek_kim_entry_q[27]));
Q_FDP4EP \dek_kim_entry_q_REG[28] ( .CK(clk), .CE(n643), .R(n649), .D(n630), .Q(dek_kim_entry_q[28]));
Q_FDP4EP \dek_kim_entry_q_REG[29] ( .CK(clk), .CE(n643), .R(n649), .D(n631), .Q(dek_kim_entry_q[29]));
Q_FDP4EP \dek_kim_entry_q_REG[30] ( .CK(clk), .CE(n643), .R(n649), .D(n632), .Q(dek_kim_entry_q[30]));
Q_FDP4EP \dek_kim_entry_q_REG[31] ( .CK(clk), .CE(n643), .R(n649), .D(n633), .Q(dek_kim_entry_q[31]));
Q_FDP4EP \dek_kim_entry_q_REG[32] ( .CK(clk), .CE(n643), .R(n649), .D(n634), .Q(dek_kim_entry_q[32]));
Q_FDP4EP \dek_kim_entry_q_REG[33] ( .CK(clk), .CE(n643), .R(n649), .D(n635), .Q(dek_kim_entry_q[33]));
Q_FDP4EP \dek_kim_entry_q_REG[34] ( .CK(clk), .CE(n643), .R(n649), .D(n636), .Q(dek_kim_entry_q[34]));
Q_FDP4EP \dek_kim_entry_q_REG[35] ( .CK(clk), .CE(n643), .R(n649), .D(n637), .Q(dek_kim_entry_q[35]));
Q_FDP4EP \dek_kim_entry_q_REG[36] ( .CK(clk), .CE(n643), .R(n649), .D(n638), .Q(dek_kim_entry_q[36]));
Q_FDP4EP \dek_kim_entry_q_REG[37] ( .CK(clk), .CE(n643), .R(n649), .D(n639), .Q(dek_kim_entry_q[37]));
Q_FDP4EP _zyL473_tfiRv7_REG  ( .CK(clk), .CE(n450), .R(n379), .D(n568), .Q(_zyL473_tfiRv7));
Q_FDP4EP _zyL468_tfiRv6_REG  ( .CK(clk), .CE(n449), .R(n379), .D(n568), .Q(_zyL468_tfiRv6));
Q_FDP4EP _zyL444_tfiRv5_REG  ( .CK(clk), .CE(n448), .R(n379), .D(n567), .Q(_zyL444_tfiRv5));
Q_FDP4EP _zyL438_tfiRv4_REG  ( .CK(clk), .CE(n447), .R(n379), .D(n567), .Q(_zyL438_tfiRv4));
Q_INV U1171 ( .A(n531), .Z(n650));
Q_FDP4EP \kim_errors_q_REG[0] ( .CK(clk), .CE(n650), .R(n649), .D(n436), .Q(kim_errors_q[0]));
Q_INV U1173 ( .A(tlv_word42[0]), .Z(n381));
Q_FDP4EP \kim_errors_q_REG[1] ( .CK(clk), .CE(n650), .R(n649), .D(n439), .Q(kim_errors_q[1]));
Q_INV U1175 ( .A(tlv_word42[1]), .Z(n388));
Q_FDP4EP \kim_errors_q_REG[2] ( .CK(clk), .CE(n650), .R(n649), .D(n440), .Q(kim_errors_q[2]));
Q_INV U1177 ( .A(tlv_word42[2]), .Z(n382));
Q_FDP4EP \kim_errors_q_REG[3] ( .CK(clk), .CE(n650), .R(n649), .D(n444), .Q(kim_errors_q[3]));
Q_FDP4EP \kim_errors_q_REG[4] ( .CK(clk), .CE(n650), .R(n649), .D(n379), .Q(kim_errors_q[4]));
Q_FDP4EP \kim_errors_q_REG[5] ( .CK(clk), .CE(n650), .R(n649), .D(n379), .Q(kim_errors_q[5]));
Q_FDP4EP \kim_errors_q_REG[6] ( .CK(clk), .CE(n650), .R(n649), .D(n379), .Q(kim_errors_q[6]));
Q_FDP4EP \kim_errors_q_REG[7] ( .CK(clk), .CE(n650), .R(n649), .D(n446), .Q(kim_errors_q[7]));
Q_INV U1183 ( .A(tlv_word42[7]), .Z(n383));
Q_FDP4EP dak_is_kdf_key_q_REG  ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[31]), .Q(dak_is_kdf_key_q));
Q_FDP4EP dek_is_kdf_key_q_REG  ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[14]), .Q(dek_is_kdf_key_q));
Q_FDP4EP \aux_key_type_REG[0] ( .CK(clk), .CE(n588), .R(n649), .D(parser_kimreader_data[39]), .Q(aux_key_type[0]));
Q_INV U1187 ( .A(aux_key_type[0]), .Z(n527));
Q_FDP4EP \aux_key_type_REG[1] ( .CK(clk), .CE(n588), .R(n649), .D(parser_kimreader_data[40]), .Q(aux_key_type[1]));
Q_INV U1189 ( .A(aux_key_type[1]), .Z(n557));
Q_FDP4EP \aux_key_type_REG[2] ( .CK(clk), .CE(n588), .R(n649), .D(parser_kimreader_data[41]), .Q(aux_key_type[2]));
Q_INV U1191 ( .A(aux_key_type[2]), .Z(n523));
Q_FDP4EP \aux_key_type_REG[3] ( .CK(clk), .CE(n588), .R(n649), .D(parser_kimreader_data[42]), .Q(aux_key_type[3]));
Q_INV U1193 ( .A(aux_key_type[3]), .Z(n530));
Q_FDP4EP \aux_key_type_REG[4] ( .CK(clk), .CE(n588), .R(n649), .D(parser_kimreader_data[43]), .Q(aux_key_type[4]));
Q_FDP4EP \aux_key_type_REG[5] ( .CK(clk), .CE(n588), .R(n649), .D(parser_kimreader_data[44]), .Q(aux_key_type[5]));
Q_FDP4EP \dak_ref_q_REG[0] ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[17]), .Q(dak_ref_q[0]));
Q_FDP4EP \dak_ref_q_REG[1] ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[18]), .Q(dak_ref_q[1]));
Q_FDP4EP \dak_ref_q_REG[2] ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[19]), .Q(dak_ref_q[2]));
Q_FDP4EP \dak_ref_q_REG[3] ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[20]), .Q(dak_ref_q[3]));
Q_FDP4EP \dak_ref_q_REG[4] ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[21]), .Q(dak_ref_q[4]));
Q_FDP4EP \dak_ref_q_REG[5] ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[22]), .Q(dak_ref_q[5]));
Q_FDP4EP \dak_ref_q_REG[6] ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[23]), .Q(dak_ref_q[6]));
Q_FDP4EP \dak_ref_q_REG[7] ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[24]), .Q(dak_ref_q[7]));
Q_FDP4EP \dak_ref_q_REG[8] ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[25]), .Q(dak_ref_q[8]));
Q_FDP4EP \dak_ref_q_REG[9] ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[26]), .Q(dak_ref_q[9]));
Q_FDP4EP \dak_ref_q_REG[10] ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[27]), .Q(dak_ref_q[10]));
Q_FDP4EP \dak_ref_q_REG[11] ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[28]), .Q(dak_ref_q[11]));
Q_FDP4EP \dak_ref_q_REG[12] ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[29]), .Q(dak_ref_q[12]));
Q_FDP4EP \dak_ref_q_REG[13] ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[30]), .Q(dak_ref_q[13]));
Q_FDP4EP \dek_ref_q_REG[0] ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[0]), .Q(dek_ref_q[0]));
Q_FDP4EP \dek_ref_q_REG[1] ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[1]), .Q(dek_ref_q[1]));
Q_FDP4EP \dek_ref_q_REG[2] ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[2]), .Q(dek_ref_q[2]));
Q_FDP4EP \dek_ref_q_REG[3] ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[3]), .Q(dek_ref_q[3]));
Q_FDP4EP \dek_ref_q_REG[4] ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[4]), .Q(dek_ref_q[4]));
Q_FDP4EP \dek_ref_q_REG[5] ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[5]), .Q(dek_ref_q[5]));
Q_FDP4EP \dek_ref_q_REG[6] ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[6]), .Q(dek_ref_q[6]));
Q_FDP4EP \dek_ref_q_REG[7] ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[7]), .Q(dek_ref_q[7]));
Q_FDP4EP \dek_ref_q_REG[8] ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[8]), .Q(dek_ref_q[8]));
Q_FDP4EP \dek_ref_q_REG[9] ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[9]), .Q(dek_ref_q[9]));
Q_FDP4EP \dek_ref_q_REG[10] ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[10]), .Q(dek_ref_q[10]));
Q_FDP4EP \dek_ref_q_REG[11] ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[11]), .Q(dek_ref_q[11]));
Q_FDP4EP \dek_ref_q_REG[12] ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[12]), .Q(dek_ref_q[12]));
Q_FDP4EP \dek_ref_q_REG[13] ( .CK(clk), .CE(n587), .R(n649), .D(parser_kimreader_data[13]), .Q(dek_ref_q[13]));
Q_FDP4EP \_zy_sva_enable_unenc_keys_10_cpass_REG[0] ( .CK(clk), .CE(n33), .R(n379), .D(n646), .Q(_zy_sva_enable_unenc_keys_10_cpass[0]));
Q_FDP4EP \_zy_sva_enable_unenc_keys_10_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n379), .D(n646), .Q(_zy_sva_enable_unenc_keys_10_ccheck[0]));
Q_FDP4EP \_zy_sva_disable_unenc_keys_9_cpass_REG[0] ( .CK(clk), .CE(n32), .R(n379), .D(n646), .Q(_zy_sva_disable_unenc_keys_9_cpass[0]));
Q_FDP4EP \_zy_sva_disable_unenc_keys_9_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n379), .D(n646), .Q(_zy_sva_disable_unenc_keys_9_ccheck[0]));
Q_FDP4EP \_zy_sva_enable_unenc_keys_8_cpass_REG[0] ( .CK(clk), .CE(n31), .R(n379), .D(n646), .Q(_zy_sva_enable_unenc_keys_8_cpass[0]));
Q_FDP4EP \_zy_sva_enable_unenc_keys_8_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n379), .D(n646), .Q(_zy_sva_enable_unenc_keys_8_ccheck[0]));
Q_FDP4EP \_zy_sva_disable_unenc_keys_7_cpass_REG[0] ( .CK(clk), .CE(n30), .R(n379), .D(n646), .Q(_zy_sva_disable_unenc_keys_7_cpass[0]));
Q_FDP4EP \_zy_sva_disable_unenc_keys_7_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n379), .D(n646), .Q(_zy_sva_disable_unenc_keys_7_ccheck[0]));
Q_FDP4EP \_zy_sva_enable_unenc_keys_6_cpass_REG[0] ( .CK(clk), .CE(n29), .R(n379), .D(n646), .Q(_zy_sva_enable_unenc_keys_6_cpass[0]));
Q_FDP4EP \_zy_sva_enable_unenc_keys_6_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n379), .D(n646), .Q(_zy_sva_enable_unenc_keys_6_ccheck[0]));
Q_FDP4EP \_zy_sva_disable_unenc_keys_5_cpass_REG[0] ( .CK(clk), .CE(n28), .R(n379), .D(n646), .Q(_zy_sva_disable_unenc_keys_5_cpass[0]));
Q_FDP4EP \_zy_sva_disable_unenc_keys_5_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n379), .D(n646), .Q(_zy_sva_disable_unenc_keys_5_ccheck[0]));
Q_FDP4EP \_zy_sva_enable_unenc_keys_4_cpass_REG[0] ( .CK(clk), .CE(n27), .R(n379), .D(n646), .Q(_zy_sva_enable_unenc_keys_4_cpass[0]));
Q_FDP4EP \_zy_sva_enable_unenc_keys_4_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n379), .D(n646), .Q(_zy_sva_enable_unenc_keys_4_ccheck[0]));
Q_FDP4EP \_zy_sva_disable_unenc_keys_3_cpass_REG[0] ( .CK(clk), .CE(n26), .R(n379), .D(n646), .Q(_zy_sva_disable_unenc_keys_3_cpass[0]));
Q_FDP4EP \_zy_sva_disable_unenc_keys_3_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n379), .D(n646), .Q(_zy_sva_disable_unenc_keys_3_ccheck[0]));
Q_FDP4EP \_zy_sva_enable_unenc_keys_2_cpass_REG[0] ( .CK(clk), .CE(n25), .R(n379), .D(n646), .Q(_zy_sva_enable_unenc_keys_2_cpass[0]));
Q_FDP4EP \_zy_sva_enable_unenc_keys_2_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n379), .D(n646), .Q(_zy_sva_enable_unenc_keys_2_ccheck[0]));
Q_FDP4EP \_zy_sva_disable_unenc_keys_1_cpass_REG[0] ( .CK(clk), .CE(n24), .R(n379), .D(n646), .Q(_zy_sva_disable_unenc_keys_1_cpass[0]));
Q_FDP4EP \_zy_sva_disable_unenc_keys_1_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n379), .D(n646), .Q(_zy_sva_disable_unenc_keys_1_ccheck[0]));
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "\kimreader_ckvreader_data.sot  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m2 "\kimreader_ckvreader_data.eoi  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m3 "\kimreader_ckvreader_data.eot  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m4 "\kimreader_ckvreader_data.id  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m5 "\kimreader_ckvreader_data.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m6 "\parser_kimreader_data.sot  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m7 "\parser_kimreader_data.eoi  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m8 "\parser_kimreader_data.eot  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m9 "\parser_kimreader_data.id  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m10 "\parser_kimreader_data.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m11 "\kim_dout.valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m12 "\kim_dout.label_index  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m13 "\kim_dout.ckv_length  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m14 "\kim_dout.ckv_pointer  (1,0) 1 14 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m15 "\kim_dout.pf_num  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m16 "\kim_dout.vf_num  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m17 "\kim_dout.vf_valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m18 "\dek_kim_entry_q.valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m19 "\dek_kim_entry_q.label_index  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m20 "\dek_kim_entry_q.ckv_length  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m21 "\dek_kim_entry_q.ckv_pointer  (1,0) 1 14 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m22 "\dek_kim_entry_q.pf_num  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m23 "\dek_kim_entry_q.vf_num  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m24 "\dek_kim_entry_q.vf_valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m25 "\dak_kim_entry_q.valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m26 "\dak_kim_entry_q.label_index  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m27 "\dak_kim_entry_q.ckv_length  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m28 "\dak_kim_entry_q.ckv_pointer  (1,0) 1 14 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m29 "\dak_kim_entry_q.pf_num  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m30 "\dak_kim_entry_q.vf_num  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m31 "\dak_kim_entry_q.vf_valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m32 "\tlv_word0.tlv_bip2  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m33 "\tlv_word0.resv0  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m34 "\tlv_word0.kdf_dek_iter  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m35 "\tlv_word0.keyless_algos  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m36 "\tlv_word0.needs_dek  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m37 "\tlv_word0.needs_dak  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m38 "\tlv_word0.key_type  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m39 "\tlv_word0.tlv_frame_num  (1,0) 1 10 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m40 "\tlv_word0.tlv_eng_id  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m41 "\tlv_word0.tlv_seq_num  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m42 "\tlv_word0.tlv_len  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m43 "\tlv_word0.tlv_type  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m44 "\tlv_word8.dek_kim_entry.valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m45 "\tlv_word8.dek_kim_entry.label_index  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m46 "\tlv_word8.dek_kim_entry.ckv_length  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m47 "\tlv_word8.dek_kim_entry.ckv_pointer  (1,0) 1 14 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m48 "\tlv_word8.dek_kim_entry.pf_num  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m49 "\tlv_word8.dek_kim_entry.vf_num  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m50 "\tlv_word8.dek_kim_entry.vf_valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m51 "\tlv_word8.unused  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m52 "\tlv_word8.missing_iv  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m53 "\tlv_word8.missing_guid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m54 "\tlv_word8.validate_dek  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m55 "\tlv_word8.vf_valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m56 "\tlv_word8.pf_num  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m57 "\tlv_word8.vf_num  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m58 "\tlv_word9.dak_kim_entry.valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m59 "\tlv_word9.dak_kim_entry.label_index  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m60 "\tlv_word9.dak_kim_entry.ckv_length  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m61 "\tlv_word9.dak_kim_entry.ckv_pointer  (1,0) 1 14 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m62 "\tlv_word9.dak_kim_entry.pf_num  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m63 "\tlv_word9.dak_kim_entry.vf_num  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m64 "\tlv_word9.dak_kim_entry.vf_valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m65 "\tlv_word9.unused  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m66 "\tlv_word9.validate_dak  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m67 "\tlv_word9.vf_valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m68 "\tlv_word9.pf_num  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m69 "\tlv_word9.vf_num  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m70 "\tlv_word42.corrupt_crc32  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m71 "\tlv_word42.unused  (1,0) 1 46 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m72 "\tlv_word42.error_code  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m73 "\aux_key_ctrl.dak_key_op  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m74 "\aux_key_ctrl.dak_key_ref  (1,0) 1 13 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m75 "\aux_key_ctrl.kdf_mode  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m76 "\aux_key_ctrl.dek_key_op  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m77 "\aux_key_ctrl.dek_key_ref  (1,0) 1 13 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "77"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r1 "kimreader_ckvreader_data 5 \kimreader_ckvreader_data.sot  \kimreader_ckvreader_data.eoi  \kimreader_ckvreader_data.eot  \kimreader_ckvreader_data.id  \kimreader_ckvreader_data.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r2 "parser_kimreader_data 5 \parser_kimreader_data.sot  \parser_kimreader_data.eoi  \parser_kimreader_data.eot  \parser_kimreader_data.id  \parser_kimreader_data.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r3 "kim_dout 7 \kim_dout.valid  \kim_dout.label_index  \kim_dout.ckv_length  \kim_dout.ckv_pointer  \kim_dout.pf_num  \kim_dout.vf_num  \kim_dout.vf_valid "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r4 "dek_kim_entry_q 7 \dek_kim_entry_q.valid  \dek_kim_entry_q.label_index  \dek_kim_entry_q.ckv_length  \dek_kim_entry_q.ckv_pointer  \dek_kim_entry_q.pf_num  \dek_kim_entry_q.vf_num  \dek_kim_entry_q.vf_valid "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r5 "dak_kim_entry_q 7 \dak_kim_entry_q.valid  \dak_kim_entry_q.label_index  \dak_kim_entry_q.ckv_length  \dak_kim_entry_q.ckv_pointer  \dak_kim_entry_q.pf_num  \dak_kim_entry_q.vf_num  \dak_kim_entry_q.vf_valid "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r6 "tlv_word0 12 \tlv_word0.tlv_bip2  \tlv_word0.resv0  \tlv_word0.kdf_dek_iter  \tlv_word0.keyless_algos  \tlv_word0.needs_dek  \tlv_word0.needs_dak  \tlv_word0.key_type  \tlv_word0.tlv_frame_num  \tlv_word0.tlv_eng_id  \tlv_word0.tlv_seq_num  \tlv_word0.tlv_len  \tlv_word0.tlv_type "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r7 "tlv_word8 8 \tlv_word8.dek_kim_entry  { \tlv_word8.dek_kim_entry.valid  \tlv_word8.dek_kim_entry.label_index  \tlv_word8.dek_kim_entry.ckv_length  \tlv_word8.dek_kim_entry.ckv_pointer  \tlv_word8.dek_kim_entry.pf_num  \tlv_word8.dek_kim_entry.vf_num  \tlv_word8.dek_kim_entry.vf_valid  } \tlv_word8.unused  \tlv_word8.missing_iv  \tlv_word8.missing_guid  \tlv_word8.validate_dek  \tlv_word8.vf_valid  \tlv_word8.pf_num  \tlv_word8.vf_num "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r8 "tlv_word9 6 \tlv_word9.dak_kim_entry  { \tlv_word9.dak_kim_entry.valid  \tlv_word9.dak_kim_entry.label_index  \tlv_word9.dak_kim_entry.ckv_length  \tlv_word9.dak_kim_entry.ckv_pointer  \tlv_word9.dak_kim_entry.pf_num  \tlv_word9.dak_kim_entry.vf_num  \tlv_word9.dak_kim_entry.vf_valid  } \tlv_word9.unused  \tlv_word9.validate_dak  \tlv_word9.vf_valid  \tlv_word9.pf_num  \tlv_word9.vf_num "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r9 "tlv_word42 3 \tlv_word42.corrupt_crc32  \tlv_word42.unused  \tlv_word42.error_code "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r10 "aux_key_ctrl 5 \aux_key_ctrl.dak_key_op  \aux_key_ctrl.dak_key_ref  \aux_key_ctrl.kdf_mode  \aux_key_ctrl.dek_key_op  \aux_key_ctrl.dek_key_ref "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_NUM "10"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_0 "-1 key_type_enc_dek 2 6 "
// pragma CVASTRPROP MODULE HDLICE PROP_RANOFF TRUE
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type_enc_dek[6]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type_enc_dek[5]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type_enc_dek[4]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type_enc_dek[3]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type_enc_dek[2]"
endmodule
