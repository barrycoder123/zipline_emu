
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module ixc_assign_611 ( L, R);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output [610:0] L;
input [610:0] R;
Q_ASSIGN U0 ( .B(R[0]), .A(L[0]));
Q_ASSIGN U1 ( .B(R[1]), .A(L[1]));
Q_ASSIGN U2 ( .B(R[2]), .A(L[2]));
Q_ASSIGN U3 ( .B(R[3]), .A(L[3]));
Q_ASSIGN U4 ( .B(R[4]), .A(L[4]));
Q_ASSIGN U5 ( .B(R[5]), .A(L[5]));
Q_ASSIGN U6 ( .B(R[6]), .A(L[6]));
Q_ASSIGN U7 ( .B(R[7]), .A(L[7]));
Q_ASSIGN U8 ( .B(R[8]), .A(L[8]));
Q_ASSIGN U9 ( .B(R[9]), .A(L[9]));
Q_ASSIGN U10 ( .B(R[10]), .A(L[10]));
Q_ASSIGN U11 ( .B(R[11]), .A(L[11]));
Q_ASSIGN U12 ( .B(R[12]), .A(L[12]));
Q_ASSIGN U13 ( .B(R[13]), .A(L[13]));
Q_ASSIGN U14 ( .B(R[14]), .A(L[14]));
Q_ASSIGN U15 ( .B(R[15]), .A(L[15]));
Q_ASSIGN U16 ( .B(R[16]), .A(L[16]));
Q_ASSIGN U17 ( .B(R[17]), .A(L[17]));
Q_ASSIGN U18 ( .B(R[18]), .A(L[18]));
Q_ASSIGN U19 ( .B(R[19]), .A(L[19]));
Q_ASSIGN U20 ( .B(R[20]), .A(L[20]));
Q_ASSIGN U21 ( .B(R[21]), .A(L[21]));
Q_ASSIGN U22 ( .B(R[22]), .A(L[22]));
Q_ASSIGN U23 ( .B(R[23]), .A(L[23]));
Q_ASSIGN U24 ( .B(R[24]), .A(L[24]));
Q_ASSIGN U25 ( .B(R[25]), .A(L[25]));
Q_ASSIGN U26 ( .B(R[26]), .A(L[26]));
Q_ASSIGN U27 ( .B(R[27]), .A(L[27]));
Q_ASSIGN U28 ( .B(R[28]), .A(L[28]));
Q_ASSIGN U29 ( .B(R[29]), .A(L[29]));
Q_ASSIGN U30 ( .B(R[30]), .A(L[30]));
Q_ASSIGN U31 ( .B(R[31]), .A(L[31]));
Q_ASSIGN U32 ( .B(R[32]), .A(L[32]));
Q_ASSIGN U33 ( .B(R[33]), .A(L[33]));
Q_ASSIGN U34 ( .B(R[34]), .A(L[34]));
Q_ASSIGN U35 ( .B(R[35]), .A(L[35]));
Q_ASSIGN U36 ( .B(R[36]), .A(L[36]));
Q_ASSIGN U37 ( .B(R[37]), .A(L[37]));
Q_ASSIGN U38 ( .B(R[38]), .A(L[38]));
Q_ASSIGN U39 ( .B(R[39]), .A(L[39]));
Q_ASSIGN U40 ( .B(R[40]), .A(L[40]));
Q_ASSIGN U41 ( .B(R[41]), .A(L[41]));
Q_ASSIGN U42 ( .B(R[42]), .A(L[42]));
Q_ASSIGN U43 ( .B(R[43]), .A(L[43]));
Q_ASSIGN U44 ( .B(R[44]), .A(L[44]));
Q_ASSIGN U45 ( .B(R[45]), .A(L[45]));
Q_ASSIGN U46 ( .B(R[46]), .A(L[46]));
Q_ASSIGN U47 ( .B(R[47]), .A(L[47]));
Q_ASSIGN U48 ( .B(R[48]), .A(L[48]));
Q_ASSIGN U49 ( .B(R[49]), .A(L[49]));
Q_ASSIGN U50 ( .B(R[50]), .A(L[50]));
Q_ASSIGN U51 ( .B(R[51]), .A(L[51]));
Q_ASSIGN U52 ( .B(R[52]), .A(L[52]));
Q_ASSIGN U53 ( .B(R[53]), .A(L[53]));
Q_ASSIGN U54 ( .B(R[54]), .A(L[54]));
Q_ASSIGN U55 ( .B(R[55]), .A(L[55]));
Q_ASSIGN U56 ( .B(R[56]), .A(L[56]));
Q_ASSIGN U57 ( .B(R[57]), .A(L[57]));
Q_ASSIGN U58 ( .B(R[58]), .A(L[58]));
Q_ASSIGN U59 ( .B(R[59]), .A(L[59]));
Q_ASSIGN U60 ( .B(R[60]), .A(L[60]));
Q_ASSIGN U61 ( .B(R[61]), .A(L[61]));
Q_ASSIGN U62 ( .B(R[62]), .A(L[62]));
Q_ASSIGN U63 ( .B(R[63]), .A(L[63]));
Q_ASSIGN U64 ( .B(R[64]), .A(L[64]));
Q_ASSIGN U65 ( .B(R[65]), .A(L[65]));
Q_ASSIGN U66 ( .B(R[66]), .A(L[66]));
Q_ASSIGN U67 ( .B(R[67]), .A(L[67]));
Q_ASSIGN U68 ( .B(R[68]), .A(L[68]));
Q_ASSIGN U69 ( .B(R[69]), .A(L[69]));
Q_ASSIGN U70 ( .B(R[70]), .A(L[70]));
Q_ASSIGN U71 ( .B(R[71]), .A(L[71]));
Q_ASSIGN U72 ( .B(R[72]), .A(L[72]));
Q_ASSIGN U73 ( .B(R[73]), .A(L[73]));
Q_ASSIGN U74 ( .B(R[74]), .A(L[74]));
Q_ASSIGN U75 ( .B(R[75]), .A(L[75]));
Q_ASSIGN U76 ( .B(R[76]), .A(L[76]));
Q_ASSIGN U77 ( .B(R[77]), .A(L[77]));
Q_ASSIGN U78 ( .B(R[78]), .A(L[78]));
Q_ASSIGN U79 ( .B(R[79]), .A(L[79]));
Q_ASSIGN U80 ( .B(R[80]), .A(L[80]));
Q_ASSIGN U81 ( .B(R[81]), .A(L[81]));
Q_ASSIGN U82 ( .B(R[82]), .A(L[82]));
Q_ASSIGN U83 ( .B(R[83]), .A(L[83]));
Q_ASSIGN U84 ( .B(R[84]), .A(L[84]));
Q_ASSIGN U85 ( .B(R[85]), .A(L[85]));
Q_ASSIGN U86 ( .B(R[86]), .A(L[86]));
Q_ASSIGN U87 ( .B(R[87]), .A(L[87]));
Q_ASSIGN U88 ( .B(R[88]), .A(L[88]));
Q_ASSIGN U89 ( .B(R[89]), .A(L[89]));
Q_ASSIGN U90 ( .B(R[90]), .A(L[90]));
Q_ASSIGN U91 ( .B(R[91]), .A(L[91]));
Q_ASSIGN U92 ( .B(R[92]), .A(L[92]));
Q_ASSIGN U93 ( .B(R[93]), .A(L[93]));
Q_ASSIGN U94 ( .B(R[94]), .A(L[94]));
Q_ASSIGN U95 ( .B(R[95]), .A(L[95]));
Q_ASSIGN U96 ( .B(R[96]), .A(L[96]));
Q_ASSIGN U97 ( .B(R[97]), .A(L[97]));
Q_ASSIGN U98 ( .B(R[98]), .A(L[98]));
Q_ASSIGN U99 ( .B(R[99]), .A(L[99]));
Q_ASSIGN U100 ( .B(R[100]), .A(L[100]));
Q_ASSIGN U101 ( .B(R[101]), .A(L[101]));
Q_ASSIGN U102 ( .B(R[102]), .A(L[102]));
Q_ASSIGN U103 ( .B(R[103]), .A(L[103]));
Q_ASSIGN U104 ( .B(R[104]), .A(L[104]));
Q_ASSIGN U105 ( .B(R[105]), .A(L[105]));
Q_ASSIGN U106 ( .B(R[106]), .A(L[106]));
Q_ASSIGN U107 ( .B(R[107]), .A(L[107]));
Q_ASSIGN U108 ( .B(R[108]), .A(L[108]));
Q_ASSIGN U109 ( .B(R[109]), .A(L[109]));
Q_ASSIGN U110 ( .B(R[110]), .A(L[110]));
Q_ASSIGN U111 ( .B(R[111]), .A(L[111]));
Q_ASSIGN U112 ( .B(R[112]), .A(L[112]));
Q_ASSIGN U113 ( .B(R[113]), .A(L[113]));
Q_ASSIGN U114 ( .B(R[114]), .A(L[114]));
Q_ASSIGN U115 ( .B(R[115]), .A(L[115]));
Q_ASSIGN U116 ( .B(R[116]), .A(L[116]));
Q_ASSIGN U117 ( .B(R[117]), .A(L[117]));
Q_ASSIGN U118 ( .B(R[118]), .A(L[118]));
Q_ASSIGN U119 ( .B(R[119]), .A(L[119]));
Q_ASSIGN U120 ( .B(R[120]), .A(L[120]));
Q_ASSIGN U121 ( .B(R[121]), .A(L[121]));
Q_ASSIGN U122 ( .B(R[122]), .A(L[122]));
Q_ASSIGN U123 ( .B(R[123]), .A(L[123]));
Q_ASSIGN U124 ( .B(R[124]), .A(L[124]));
Q_ASSIGN U125 ( .B(R[125]), .A(L[125]));
Q_ASSIGN U126 ( .B(R[126]), .A(L[126]));
Q_ASSIGN U127 ( .B(R[127]), .A(L[127]));
Q_ASSIGN U128 ( .B(R[128]), .A(L[128]));
Q_ASSIGN U129 ( .B(R[129]), .A(L[129]));
Q_ASSIGN U130 ( .B(R[130]), .A(L[130]));
Q_ASSIGN U131 ( .B(R[131]), .A(L[131]));
Q_ASSIGN U132 ( .B(R[132]), .A(L[132]));
Q_ASSIGN U133 ( .B(R[133]), .A(L[133]));
Q_ASSIGN U134 ( .B(R[134]), .A(L[134]));
Q_ASSIGN U135 ( .B(R[135]), .A(L[135]));
Q_ASSIGN U136 ( .B(R[136]), .A(L[136]));
Q_ASSIGN U137 ( .B(R[137]), .A(L[137]));
Q_ASSIGN U138 ( .B(R[138]), .A(L[138]));
Q_ASSIGN U139 ( .B(R[139]), .A(L[139]));
Q_ASSIGN U140 ( .B(R[140]), .A(L[140]));
Q_ASSIGN U141 ( .B(R[141]), .A(L[141]));
Q_ASSIGN U142 ( .B(R[142]), .A(L[142]));
Q_ASSIGN U143 ( .B(R[143]), .A(L[143]));
Q_ASSIGN U144 ( .B(R[144]), .A(L[144]));
Q_ASSIGN U145 ( .B(R[145]), .A(L[145]));
Q_ASSIGN U146 ( .B(R[146]), .A(L[146]));
Q_ASSIGN U147 ( .B(R[147]), .A(L[147]));
Q_ASSIGN U148 ( .B(R[148]), .A(L[148]));
Q_ASSIGN U149 ( .B(R[149]), .A(L[149]));
Q_ASSIGN U150 ( .B(R[150]), .A(L[150]));
Q_ASSIGN U151 ( .B(R[151]), .A(L[151]));
Q_ASSIGN U152 ( .B(R[152]), .A(L[152]));
Q_ASSIGN U153 ( .B(R[153]), .A(L[153]));
Q_ASSIGN U154 ( .B(R[154]), .A(L[154]));
Q_ASSIGN U155 ( .B(R[155]), .A(L[155]));
Q_ASSIGN U156 ( .B(R[156]), .A(L[156]));
Q_ASSIGN U157 ( .B(R[157]), .A(L[157]));
Q_ASSIGN U158 ( .B(R[158]), .A(L[158]));
Q_ASSIGN U159 ( .B(R[159]), .A(L[159]));
Q_ASSIGN U160 ( .B(R[160]), .A(L[160]));
Q_ASSIGN U161 ( .B(R[161]), .A(L[161]));
Q_ASSIGN U162 ( .B(R[162]), .A(L[162]));
Q_ASSIGN U163 ( .B(R[163]), .A(L[163]));
Q_ASSIGN U164 ( .B(R[164]), .A(L[164]));
Q_ASSIGN U165 ( .B(R[165]), .A(L[165]));
Q_ASSIGN U166 ( .B(R[166]), .A(L[166]));
Q_ASSIGN U167 ( .B(R[167]), .A(L[167]));
Q_ASSIGN U168 ( .B(R[168]), .A(L[168]));
Q_ASSIGN U169 ( .B(R[169]), .A(L[169]));
Q_ASSIGN U170 ( .B(R[170]), .A(L[170]));
Q_ASSIGN U171 ( .B(R[171]), .A(L[171]));
Q_ASSIGN U172 ( .B(R[172]), .A(L[172]));
Q_ASSIGN U173 ( .B(R[173]), .A(L[173]));
Q_ASSIGN U174 ( .B(R[174]), .A(L[174]));
Q_ASSIGN U175 ( .B(R[175]), .A(L[175]));
Q_ASSIGN U176 ( .B(R[176]), .A(L[176]));
Q_ASSIGN U177 ( .B(R[177]), .A(L[177]));
Q_ASSIGN U178 ( .B(R[178]), .A(L[178]));
Q_ASSIGN U179 ( .B(R[179]), .A(L[179]));
Q_ASSIGN U180 ( .B(R[180]), .A(L[180]));
Q_ASSIGN U181 ( .B(R[181]), .A(L[181]));
Q_ASSIGN U182 ( .B(R[182]), .A(L[182]));
Q_ASSIGN U183 ( .B(R[183]), .A(L[183]));
Q_ASSIGN U184 ( .B(R[184]), .A(L[184]));
Q_ASSIGN U185 ( .B(R[185]), .A(L[185]));
Q_ASSIGN U186 ( .B(R[186]), .A(L[186]));
Q_ASSIGN U187 ( .B(R[187]), .A(L[187]));
Q_ASSIGN U188 ( .B(R[188]), .A(L[188]));
Q_ASSIGN U189 ( .B(R[189]), .A(L[189]));
Q_ASSIGN U190 ( .B(R[190]), .A(L[190]));
Q_ASSIGN U191 ( .B(R[191]), .A(L[191]));
Q_ASSIGN U192 ( .B(R[192]), .A(L[192]));
Q_ASSIGN U193 ( .B(R[193]), .A(L[193]));
Q_ASSIGN U194 ( .B(R[194]), .A(L[194]));
Q_ASSIGN U195 ( .B(R[195]), .A(L[195]));
Q_ASSIGN U196 ( .B(R[196]), .A(L[196]));
Q_ASSIGN U197 ( .B(R[197]), .A(L[197]));
Q_ASSIGN U198 ( .B(R[198]), .A(L[198]));
Q_ASSIGN U199 ( .B(R[199]), .A(L[199]));
Q_ASSIGN U200 ( .B(R[200]), .A(L[200]));
Q_ASSIGN U201 ( .B(R[201]), .A(L[201]));
Q_ASSIGN U202 ( .B(R[202]), .A(L[202]));
Q_ASSIGN U203 ( .B(R[203]), .A(L[203]));
Q_ASSIGN U204 ( .B(R[204]), .A(L[204]));
Q_ASSIGN U205 ( .B(R[205]), .A(L[205]));
Q_ASSIGN U206 ( .B(R[206]), .A(L[206]));
Q_ASSIGN U207 ( .B(R[207]), .A(L[207]));
Q_ASSIGN U208 ( .B(R[208]), .A(L[208]));
Q_ASSIGN U209 ( .B(R[209]), .A(L[209]));
Q_ASSIGN U210 ( .B(R[210]), .A(L[210]));
Q_ASSIGN U211 ( .B(R[211]), .A(L[211]));
Q_ASSIGN U212 ( .B(R[212]), .A(L[212]));
Q_ASSIGN U213 ( .B(R[213]), .A(L[213]));
Q_ASSIGN U214 ( .B(R[214]), .A(L[214]));
Q_ASSIGN U215 ( .B(R[215]), .A(L[215]));
Q_ASSIGN U216 ( .B(R[216]), .A(L[216]));
Q_ASSIGN U217 ( .B(R[217]), .A(L[217]));
Q_ASSIGN U218 ( .B(R[218]), .A(L[218]));
Q_ASSIGN U219 ( .B(R[219]), .A(L[219]));
Q_ASSIGN U220 ( .B(R[220]), .A(L[220]));
Q_ASSIGN U221 ( .B(R[221]), .A(L[221]));
Q_ASSIGN U222 ( .B(R[222]), .A(L[222]));
Q_ASSIGN U223 ( .B(R[223]), .A(L[223]));
Q_ASSIGN U224 ( .B(R[224]), .A(L[224]));
Q_ASSIGN U225 ( .B(R[225]), .A(L[225]));
Q_ASSIGN U226 ( .B(R[226]), .A(L[226]));
Q_ASSIGN U227 ( .B(R[227]), .A(L[227]));
Q_ASSIGN U228 ( .B(R[228]), .A(L[228]));
Q_ASSIGN U229 ( .B(R[229]), .A(L[229]));
Q_ASSIGN U230 ( .B(R[230]), .A(L[230]));
Q_ASSIGN U231 ( .B(R[231]), .A(L[231]));
Q_ASSIGN U232 ( .B(R[232]), .A(L[232]));
Q_ASSIGN U233 ( .B(R[233]), .A(L[233]));
Q_ASSIGN U234 ( .B(R[234]), .A(L[234]));
Q_ASSIGN U235 ( .B(R[235]), .A(L[235]));
Q_ASSIGN U236 ( .B(R[236]), .A(L[236]));
Q_ASSIGN U237 ( .B(R[237]), .A(L[237]));
Q_ASSIGN U238 ( .B(R[238]), .A(L[238]));
Q_ASSIGN U239 ( .B(R[239]), .A(L[239]));
Q_ASSIGN U240 ( .B(R[240]), .A(L[240]));
Q_ASSIGN U241 ( .B(R[241]), .A(L[241]));
Q_ASSIGN U242 ( .B(R[242]), .A(L[242]));
Q_ASSIGN U243 ( .B(R[243]), .A(L[243]));
Q_ASSIGN U244 ( .B(R[244]), .A(L[244]));
Q_ASSIGN U245 ( .B(R[245]), .A(L[245]));
Q_ASSIGN U246 ( .B(R[246]), .A(L[246]));
Q_ASSIGN U247 ( .B(R[247]), .A(L[247]));
Q_ASSIGN U248 ( .B(R[248]), .A(L[248]));
Q_ASSIGN U249 ( .B(R[249]), .A(L[249]));
Q_ASSIGN U250 ( .B(R[250]), .A(L[250]));
Q_ASSIGN U251 ( .B(R[251]), .A(L[251]));
Q_ASSIGN U252 ( .B(R[252]), .A(L[252]));
Q_ASSIGN U253 ( .B(R[253]), .A(L[253]));
Q_ASSIGN U254 ( .B(R[254]), .A(L[254]));
Q_ASSIGN U255 ( .B(R[255]), .A(L[255]));
Q_ASSIGN U256 ( .B(R[256]), .A(L[256]));
Q_ASSIGN U257 ( .B(R[257]), .A(L[257]));
Q_ASSIGN U258 ( .B(R[258]), .A(L[258]));
Q_ASSIGN U259 ( .B(R[259]), .A(L[259]));
Q_ASSIGN U260 ( .B(R[260]), .A(L[260]));
Q_ASSIGN U261 ( .B(R[261]), .A(L[261]));
Q_ASSIGN U262 ( .B(R[262]), .A(L[262]));
Q_ASSIGN U263 ( .B(R[263]), .A(L[263]));
Q_ASSIGN U264 ( .B(R[264]), .A(L[264]));
Q_ASSIGN U265 ( .B(R[265]), .A(L[265]));
Q_ASSIGN U266 ( .B(R[266]), .A(L[266]));
Q_ASSIGN U267 ( .B(R[267]), .A(L[267]));
Q_ASSIGN U268 ( .B(R[268]), .A(L[268]));
Q_ASSIGN U269 ( .B(R[269]), .A(L[269]));
Q_ASSIGN U270 ( .B(R[270]), .A(L[270]));
Q_ASSIGN U271 ( .B(R[271]), .A(L[271]));
Q_ASSIGN U272 ( .B(R[272]), .A(L[272]));
Q_ASSIGN U273 ( .B(R[273]), .A(L[273]));
Q_ASSIGN U274 ( .B(R[274]), .A(L[274]));
Q_ASSIGN U275 ( .B(R[275]), .A(L[275]));
Q_ASSIGN U276 ( .B(R[276]), .A(L[276]));
Q_ASSIGN U277 ( .B(R[277]), .A(L[277]));
Q_ASSIGN U278 ( .B(R[278]), .A(L[278]));
Q_ASSIGN U279 ( .B(R[279]), .A(L[279]));
Q_ASSIGN U280 ( .B(R[280]), .A(L[280]));
Q_ASSIGN U281 ( .B(R[281]), .A(L[281]));
Q_ASSIGN U282 ( .B(R[282]), .A(L[282]));
Q_ASSIGN U283 ( .B(R[283]), .A(L[283]));
Q_ASSIGN U284 ( .B(R[284]), .A(L[284]));
Q_ASSIGN U285 ( .B(R[285]), .A(L[285]));
Q_ASSIGN U286 ( .B(R[286]), .A(L[286]));
Q_ASSIGN U287 ( .B(R[287]), .A(L[287]));
Q_ASSIGN U288 ( .B(R[288]), .A(L[288]));
Q_ASSIGN U289 ( .B(R[289]), .A(L[289]));
Q_ASSIGN U290 ( .B(R[290]), .A(L[290]));
Q_ASSIGN U291 ( .B(R[291]), .A(L[291]));
Q_ASSIGN U292 ( .B(R[292]), .A(L[292]));
Q_ASSIGN U293 ( .B(R[293]), .A(L[293]));
Q_ASSIGN U294 ( .B(R[294]), .A(L[294]));
Q_ASSIGN U295 ( .B(R[295]), .A(L[295]));
Q_ASSIGN U296 ( .B(R[296]), .A(L[296]));
Q_ASSIGN U297 ( .B(R[297]), .A(L[297]));
Q_ASSIGN U298 ( .B(R[298]), .A(L[298]));
Q_ASSIGN U299 ( .B(R[299]), .A(L[299]));
Q_ASSIGN U300 ( .B(R[300]), .A(L[300]));
Q_ASSIGN U301 ( .B(R[301]), .A(L[301]));
Q_ASSIGN U302 ( .B(R[302]), .A(L[302]));
Q_ASSIGN U303 ( .B(R[303]), .A(L[303]));
Q_ASSIGN U304 ( .B(R[304]), .A(L[304]));
Q_ASSIGN U305 ( .B(R[305]), .A(L[305]));
Q_ASSIGN U306 ( .B(R[306]), .A(L[306]));
Q_ASSIGN U307 ( .B(R[307]), .A(L[307]));
Q_ASSIGN U308 ( .B(R[308]), .A(L[308]));
Q_ASSIGN U309 ( .B(R[309]), .A(L[309]));
Q_ASSIGN U310 ( .B(R[310]), .A(L[310]));
Q_ASSIGN U311 ( .B(R[311]), .A(L[311]));
Q_ASSIGN U312 ( .B(R[312]), .A(L[312]));
Q_ASSIGN U313 ( .B(R[313]), .A(L[313]));
Q_ASSIGN U314 ( .B(R[314]), .A(L[314]));
Q_ASSIGN U315 ( .B(R[315]), .A(L[315]));
Q_ASSIGN U316 ( .B(R[316]), .A(L[316]));
Q_ASSIGN U317 ( .B(R[317]), .A(L[317]));
Q_ASSIGN U318 ( .B(R[318]), .A(L[318]));
Q_ASSIGN U319 ( .B(R[319]), .A(L[319]));
Q_ASSIGN U320 ( .B(R[320]), .A(L[320]));
Q_ASSIGN U321 ( .B(R[321]), .A(L[321]));
Q_ASSIGN U322 ( .B(R[322]), .A(L[322]));
Q_ASSIGN U323 ( .B(R[323]), .A(L[323]));
Q_ASSIGN U324 ( .B(R[324]), .A(L[324]));
Q_ASSIGN U325 ( .B(R[325]), .A(L[325]));
Q_ASSIGN U326 ( .B(R[326]), .A(L[326]));
Q_ASSIGN U327 ( .B(R[327]), .A(L[327]));
Q_ASSIGN U328 ( .B(R[328]), .A(L[328]));
Q_ASSIGN U329 ( .B(R[329]), .A(L[329]));
Q_ASSIGN U330 ( .B(R[330]), .A(L[330]));
Q_ASSIGN U331 ( .B(R[331]), .A(L[331]));
Q_ASSIGN U332 ( .B(R[332]), .A(L[332]));
Q_ASSIGN U333 ( .B(R[333]), .A(L[333]));
Q_ASSIGN U334 ( .B(R[334]), .A(L[334]));
Q_ASSIGN U335 ( .B(R[335]), .A(L[335]));
Q_ASSIGN U336 ( .B(R[336]), .A(L[336]));
Q_ASSIGN U337 ( .B(R[337]), .A(L[337]));
Q_ASSIGN U338 ( .B(R[338]), .A(L[338]));
Q_ASSIGN U339 ( .B(R[339]), .A(L[339]));
Q_ASSIGN U340 ( .B(R[340]), .A(L[340]));
Q_ASSIGN U341 ( .B(R[341]), .A(L[341]));
Q_ASSIGN U342 ( .B(R[342]), .A(L[342]));
Q_ASSIGN U343 ( .B(R[343]), .A(L[343]));
Q_ASSIGN U344 ( .B(R[344]), .A(L[344]));
Q_ASSIGN U345 ( .B(R[345]), .A(L[345]));
Q_ASSIGN U346 ( .B(R[346]), .A(L[346]));
Q_ASSIGN U347 ( .B(R[347]), .A(L[347]));
Q_ASSIGN U348 ( .B(R[348]), .A(L[348]));
Q_ASSIGN U349 ( .B(R[349]), .A(L[349]));
Q_ASSIGN U350 ( .B(R[350]), .A(L[350]));
Q_ASSIGN U351 ( .B(R[351]), .A(L[351]));
Q_ASSIGN U352 ( .B(R[352]), .A(L[352]));
Q_ASSIGN U353 ( .B(R[353]), .A(L[353]));
Q_ASSIGN U354 ( .B(R[354]), .A(L[354]));
Q_ASSIGN U355 ( .B(R[355]), .A(L[355]));
Q_ASSIGN U356 ( .B(R[356]), .A(L[356]));
Q_ASSIGN U357 ( .B(R[357]), .A(L[357]));
Q_ASSIGN U358 ( .B(R[358]), .A(L[358]));
Q_ASSIGN U359 ( .B(R[359]), .A(L[359]));
Q_ASSIGN U360 ( .B(R[360]), .A(L[360]));
Q_ASSIGN U361 ( .B(R[361]), .A(L[361]));
Q_ASSIGN U362 ( .B(R[362]), .A(L[362]));
Q_ASSIGN U363 ( .B(R[363]), .A(L[363]));
Q_ASSIGN U364 ( .B(R[364]), .A(L[364]));
Q_ASSIGN U365 ( .B(R[365]), .A(L[365]));
Q_ASSIGN U366 ( .B(R[366]), .A(L[366]));
Q_ASSIGN U367 ( .B(R[367]), .A(L[367]));
Q_ASSIGN U368 ( .B(R[368]), .A(L[368]));
Q_ASSIGN U369 ( .B(R[369]), .A(L[369]));
Q_ASSIGN U370 ( .B(R[370]), .A(L[370]));
Q_ASSIGN U371 ( .B(R[371]), .A(L[371]));
Q_ASSIGN U372 ( .B(R[372]), .A(L[372]));
Q_ASSIGN U373 ( .B(R[373]), .A(L[373]));
Q_ASSIGN U374 ( .B(R[374]), .A(L[374]));
Q_ASSIGN U375 ( .B(R[375]), .A(L[375]));
Q_ASSIGN U376 ( .B(R[376]), .A(L[376]));
Q_ASSIGN U377 ( .B(R[377]), .A(L[377]));
Q_ASSIGN U378 ( .B(R[378]), .A(L[378]));
Q_ASSIGN U379 ( .B(R[379]), .A(L[379]));
Q_ASSIGN U380 ( .B(R[380]), .A(L[380]));
Q_ASSIGN U381 ( .B(R[381]), .A(L[381]));
Q_ASSIGN U382 ( .B(R[382]), .A(L[382]));
Q_ASSIGN U383 ( .B(R[383]), .A(L[383]));
Q_ASSIGN U384 ( .B(R[384]), .A(L[384]));
Q_ASSIGN U385 ( .B(R[385]), .A(L[385]));
Q_ASSIGN U386 ( .B(R[386]), .A(L[386]));
Q_ASSIGN U387 ( .B(R[387]), .A(L[387]));
Q_ASSIGN U388 ( .B(R[388]), .A(L[388]));
Q_ASSIGN U389 ( .B(R[389]), .A(L[389]));
Q_ASSIGN U390 ( .B(R[390]), .A(L[390]));
Q_ASSIGN U391 ( .B(R[391]), .A(L[391]));
Q_ASSIGN U392 ( .B(R[392]), .A(L[392]));
Q_ASSIGN U393 ( .B(R[393]), .A(L[393]));
Q_ASSIGN U394 ( .B(R[394]), .A(L[394]));
Q_ASSIGN U395 ( .B(R[395]), .A(L[395]));
Q_ASSIGN U396 ( .B(R[396]), .A(L[396]));
Q_ASSIGN U397 ( .B(R[397]), .A(L[397]));
Q_ASSIGN U398 ( .B(R[398]), .A(L[398]));
Q_ASSIGN U399 ( .B(R[399]), .A(L[399]));
Q_ASSIGN U400 ( .B(R[400]), .A(L[400]));
Q_ASSIGN U401 ( .B(R[401]), .A(L[401]));
Q_ASSIGN U402 ( .B(R[402]), .A(L[402]));
Q_ASSIGN U403 ( .B(R[403]), .A(L[403]));
Q_ASSIGN U404 ( .B(R[404]), .A(L[404]));
Q_ASSIGN U405 ( .B(R[405]), .A(L[405]));
Q_ASSIGN U406 ( .B(R[406]), .A(L[406]));
Q_ASSIGN U407 ( .B(R[407]), .A(L[407]));
Q_ASSIGN U408 ( .B(R[408]), .A(L[408]));
Q_ASSIGN U409 ( .B(R[409]), .A(L[409]));
Q_ASSIGN U410 ( .B(R[410]), .A(L[410]));
Q_ASSIGN U411 ( .B(R[411]), .A(L[411]));
Q_ASSIGN U412 ( .B(R[412]), .A(L[412]));
Q_ASSIGN U413 ( .B(R[413]), .A(L[413]));
Q_ASSIGN U414 ( .B(R[414]), .A(L[414]));
Q_ASSIGN U415 ( .B(R[415]), .A(L[415]));
Q_ASSIGN U416 ( .B(R[416]), .A(L[416]));
Q_ASSIGN U417 ( .B(R[417]), .A(L[417]));
Q_ASSIGN U418 ( .B(R[418]), .A(L[418]));
Q_ASSIGN U419 ( .B(R[419]), .A(L[419]));
Q_ASSIGN U420 ( .B(R[420]), .A(L[420]));
Q_ASSIGN U421 ( .B(R[421]), .A(L[421]));
Q_ASSIGN U422 ( .B(R[422]), .A(L[422]));
Q_ASSIGN U423 ( .B(R[423]), .A(L[423]));
Q_ASSIGN U424 ( .B(R[424]), .A(L[424]));
Q_ASSIGN U425 ( .B(R[425]), .A(L[425]));
Q_ASSIGN U426 ( .B(R[426]), .A(L[426]));
Q_ASSIGN U427 ( .B(R[427]), .A(L[427]));
Q_ASSIGN U428 ( .B(R[428]), .A(L[428]));
Q_ASSIGN U429 ( .B(R[429]), .A(L[429]));
Q_ASSIGN U430 ( .B(R[430]), .A(L[430]));
Q_ASSIGN U431 ( .B(R[431]), .A(L[431]));
Q_ASSIGN U432 ( .B(R[432]), .A(L[432]));
Q_ASSIGN U433 ( .B(R[433]), .A(L[433]));
Q_ASSIGN U434 ( .B(R[434]), .A(L[434]));
Q_ASSIGN U435 ( .B(R[435]), .A(L[435]));
Q_ASSIGN U436 ( .B(R[436]), .A(L[436]));
Q_ASSIGN U437 ( .B(R[437]), .A(L[437]));
Q_ASSIGN U438 ( .B(R[438]), .A(L[438]));
Q_ASSIGN U439 ( .B(R[439]), .A(L[439]));
Q_ASSIGN U440 ( .B(R[440]), .A(L[440]));
Q_ASSIGN U441 ( .B(R[441]), .A(L[441]));
Q_ASSIGN U442 ( .B(R[442]), .A(L[442]));
Q_ASSIGN U443 ( .B(R[443]), .A(L[443]));
Q_ASSIGN U444 ( .B(R[444]), .A(L[444]));
Q_ASSIGN U445 ( .B(R[445]), .A(L[445]));
Q_ASSIGN U446 ( .B(R[446]), .A(L[446]));
Q_ASSIGN U447 ( .B(R[447]), .A(L[447]));
Q_ASSIGN U448 ( .B(R[448]), .A(L[448]));
Q_ASSIGN U449 ( .B(R[449]), .A(L[449]));
Q_ASSIGN U450 ( .B(R[450]), .A(L[450]));
Q_ASSIGN U451 ( .B(R[451]), .A(L[451]));
Q_ASSIGN U452 ( .B(R[452]), .A(L[452]));
Q_ASSIGN U453 ( .B(R[453]), .A(L[453]));
Q_ASSIGN U454 ( .B(R[454]), .A(L[454]));
Q_ASSIGN U455 ( .B(R[455]), .A(L[455]));
Q_ASSIGN U456 ( .B(R[456]), .A(L[456]));
Q_ASSIGN U457 ( .B(R[457]), .A(L[457]));
Q_ASSIGN U458 ( .B(R[458]), .A(L[458]));
Q_ASSIGN U459 ( .B(R[459]), .A(L[459]));
Q_ASSIGN U460 ( .B(R[460]), .A(L[460]));
Q_ASSIGN U461 ( .B(R[461]), .A(L[461]));
Q_ASSIGN U462 ( .B(R[462]), .A(L[462]));
Q_ASSIGN U463 ( .B(R[463]), .A(L[463]));
Q_ASSIGN U464 ( .B(R[464]), .A(L[464]));
Q_ASSIGN U465 ( .B(R[465]), .A(L[465]));
Q_ASSIGN U466 ( .B(R[466]), .A(L[466]));
Q_ASSIGN U467 ( .B(R[467]), .A(L[467]));
Q_ASSIGN U468 ( .B(R[468]), .A(L[468]));
Q_ASSIGN U469 ( .B(R[469]), .A(L[469]));
Q_ASSIGN U470 ( .B(R[470]), .A(L[470]));
Q_ASSIGN U471 ( .B(R[471]), .A(L[471]));
Q_ASSIGN U472 ( .B(R[472]), .A(L[472]));
Q_ASSIGN U473 ( .B(R[473]), .A(L[473]));
Q_ASSIGN U474 ( .B(R[474]), .A(L[474]));
Q_ASSIGN U475 ( .B(R[475]), .A(L[475]));
Q_ASSIGN U476 ( .B(R[476]), .A(L[476]));
Q_ASSIGN U477 ( .B(R[477]), .A(L[477]));
Q_ASSIGN U478 ( .B(R[478]), .A(L[478]));
Q_ASSIGN U479 ( .B(R[479]), .A(L[479]));
Q_ASSIGN U480 ( .B(R[480]), .A(L[480]));
Q_ASSIGN U481 ( .B(R[481]), .A(L[481]));
Q_ASSIGN U482 ( .B(R[482]), .A(L[482]));
Q_ASSIGN U483 ( .B(R[483]), .A(L[483]));
Q_ASSIGN U484 ( .B(R[484]), .A(L[484]));
Q_ASSIGN U485 ( .B(R[485]), .A(L[485]));
Q_ASSIGN U486 ( .B(R[486]), .A(L[486]));
Q_ASSIGN U487 ( .B(R[487]), .A(L[487]));
Q_ASSIGN U488 ( .B(R[488]), .A(L[488]));
Q_ASSIGN U489 ( .B(R[489]), .A(L[489]));
Q_ASSIGN U490 ( .B(R[490]), .A(L[490]));
Q_ASSIGN U491 ( .B(R[491]), .A(L[491]));
Q_ASSIGN U492 ( .B(R[492]), .A(L[492]));
Q_ASSIGN U493 ( .B(R[493]), .A(L[493]));
Q_ASSIGN U494 ( .B(R[494]), .A(L[494]));
Q_ASSIGN U495 ( .B(R[495]), .A(L[495]));
Q_ASSIGN U496 ( .B(R[496]), .A(L[496]));
Q_ASSIGN U497 ( .B(R[497]), .A(L[497]));
Q_ASSIGN U498 ( .B(R[498]), .A(L[498]));
Q_ASSIGN U499 ( .B(R[499]), .A(L[499]));
Q_ASSIGN U500 ( .B(R[500]), .A(L[500]));
Q_ASSIGN U501 ( .B(R[501]), .A(L[501]));
Q_ASSIGN U502 ( .B(R[502]), .A(L[502]));
Q_ASSIGN U503 ( .B(R[503]), .A(L[503]));
Q_ASSIGN U504 ( .B(R[504]), .A(L[504]));
Q_ASSIGN U505 ( .B(R[505]), .A(L[505]));
Q_ASSIGN U506 ( .B(R[506]), .A(L[506]));
Q_ASSIGN U507 ( .B(R[507]), .A(L[507]));
Q_ASSIGN U508 ( .B(R[508]), .A(L[508]));
Q_ASSIGN U509 ( .B(R[509]), .A(L[509]));
Q_ASSIGN U510 ( .B(R[510]), .A(L[510]));
Q_ASSIGN U511 ( .B(R[511]), .A(L[511]));
Q_ASSIGN U512 ( .B(R[512]), .A(L[512]));
Q_ASSIGN U513 ( .B(R[513]), .A(L[513]));
Q_ASSIGN U514 ( .B(R[514]), .A(L[514]));
Q_ASSIGN U515 ( .B(R[515]), .A(L[515]));
Q_ASSIGN U516 ( .B(R[516]), .A(L[516]));
Q_ASSIGN U517 ( .B(R[517]), .A(L[517]));
Q_ASSIGN U518 ( .B(R[518]), .A(L[518]));
Q_ASSIGN U519 ( .B(R[519]), .A(L[519]));
Q_ASSIGN U520 ( .B(R[520]), .A(L[520]));
Q_ASSIGN U521 ( .B(R[521]), .A(L[521]));
Q_ASSIGN U522 ( .B(R[522]), .A(L[522]));
Q_ASSIGN U523 ( .B(R[523]), .A(L[523]));
Q_ASSIGN U524 ( .B(R[524]), .A(L[524]));
Q_ASSIGN U525 ( .B(R[525]), .A(L[525]));
Q_ASSIGN U526 ( .B(R[526]), .A(L[526]));
Q_ASSIGN U527 ( .B(R[527]), .A(L[527]));
Q_ASSIGN U528 ( .B(R[528]), .A(L[528]));
Q_ASSIGN U529 ( .B(R[529]), .A(L[529]));
Q_ASSIGN U530 ( .B(R[530]), .A(L[530]));
Q_ASSIGN U531 ( .B(R[531]), .A(L[531]));
Q_ASSIGN U532 ( .B(R[532]), .A(L[532]));
Q_ASSIGN U533 ( .B(R[533]), .A(L[533]));
Q_ASSIGN U534 ( .B(R[534]), .A(L[534]));
Q_ASSIGN U535 ( .B(R[535]), .A(L[535]));
Q_ASSIGN U536 ( .B(R[536]), .A(L[536]));
Q_ASSIGN U537 ( .B(R[537]), .A(L[537]));
Q_ASSIGN U538 ( .B(R[538]), .A(L[538]));
Q_ASSIGN U539 ( .B(R[539]), .A(L[539]));
Q_ASSIGN U540 ( .B(R[540]), .A(L[540]));
Q_ASSIGN U541 ( .B(R[541]), .A(L[541]));
Q_ASSIGN U542 ( .B(R[542]), .A(L[542]));
Q_ASSIGN U543 ( .B(R[543]), .A(L[543]));
Q_ASSIGN U544 ( .B(R[544]), .A(L[544]));
Q_ASSIGN U545 ( .B(R[545]), .A(L[545]));
Q_ASSIGN U546 ( .B(R[546]), .A(L[546]));
Q_ASSIGN U547 ( .B(R[547]), .A(L[547]));
Q_ASSIGN U548 ( .B(R[548]), .A(L[548]));
Q_ASSIGN U549 ( .B(R[549]), .A(L[549]));
Q_ASSIGN U550 ( .B(R[550]), .A(L[550]));
Q_ASSIGN U551 ( .B(R[551]), .A(L[551]));
Q_ASSIGN U552 ( .B(R[552]), .A(L[552]));
Q_ASSIGN U553 ( .B(R[553]), .A(L[553]));
Q_ASSIGN U554 ( .B(R[554]), .A(L[554]));
Q_ASSIGN U555 ( .B(R[555]), .A(L[555]));
Q_ASSIGN U556 ( .B(R[556]), .A(L[556]));
Q_ASSIGN U557 ( .B(R[557]), .A(L[557]));
Q_ASSIGN U558 ( .B(R[558]), .A(L[558]));
Q_ASSIGN U559 ( .B(R[559]), .A(L[559]));
Q_ASSIGN U560 ( .B(R[560]), .A(L[560]));
Q_ASSIGN U561 ( .B(R[561]), .A(L[561]));
Q_ASSIGN U562 ( .B(R[562]), .A(L[562]));
Q_ASSIGN U563 ( .B(R[563]), .A(L[563]));
Q_ASSIGN U564 ( .B(R[564]), .A(L[564]));
Q_ASSIGN U565 ( .B(R[565]), .A(L[565]));
Q_ASSIGN U566 ( .B(R[566]), .A(L[566]));
Q_ASSIGN U567 ( .B(R[567]), .A(L[567]));
Q_ASSIGN U568 ( .B(R[568]), .A(L[568]));
Q_ASSIGN U569 ( .B(R[569]), .A(L[569]));
Q_ASSIGN U570 ( .B(R[570]), .A(L[570]));
Q_ASSIGN U571 ( .B(R[571]), .A(L[571]));
Q_ASSIGN U572 ( .B(R[572]), .A(L[572]));
Q_ASSIGN U573 ( .B(R[573]), .A(L[573]));
Q_ASSIGN U574 ( .B(R[574]), .A(L[574]));
Q_ASSIGN U575 ( .B(R[575]), .A(L[575]));
Q_ASSIGN U576 ( .B(R[576]), .A(L[576]));
Q_ASSIGN U577 ( .B(R[577]), .A(L[577]));
Q_ASSIGN U578 ( .B(R[578]), .A(L[578]));
Q_ASSIGN U579 ( .B(R[579]), .A(L[579]));
Q_ASSIGN U580 ( .B(R[580]), .A(L[580]));
Q_ASSIGN U581 ( .B(R[581]), .A(L[581]));
Q_ASSIGN U582 ( .B(R[582]), .A(L[582]));
Q_ASSIGN U583 ( .B(R[583]), .A(L[583]));
Q_ASSIGN U584 ( .B(R[584]), .A(L[584]));
Q_ASSIGN U585 ( .B(R[585]), .A(L[585]));
Q_ASSIGN U586 ( .B(R[586]), .A(L[586]));
Q_ASSIGN U587 ( .B(R[587]), .A(L[587]));
Q_ASSIGN U588 ( .B(R[588]), .A(L[588]));
Q_ASSIGN U589 ( .B(R[589]), .A(L[589]));
Q_ASSIGN U590 ( .B(R[590]), .A(L[590]));
Q_ASSIGN U591 ( .B(R[591]), .A(L[591]));
Q_ASSIGN U592 ( .B(R[592]), .A(L[592]));
Q_ASSIGN U593 ( .B(R[593]), .A(L[593]));
Q_ASSIGN U594 ( .B(R[594]), .A(L[594]));
Q_ASSIGN U595 ( .B(R[595]), .A(L[595]));
Q_ASSIGN U596 ( .B(R[596]), .A(L[596]));
Q_ASSIGN U597 ( .B(R[597]), .A(L[597]));
Q_ASSIGN U598 ( .B(R[598]), .A(L[598]));
Q_ASSIGN U599 ( .B(R[599]), .A(L[599]));
Q_ASSIGN U600 ( .B(R[600]), .A(L[600]));
Q_ASSIGN U601 ( .B(R[601]), .A(L[601]));
Q_ASSIGN U602 ( .B(R[602]), .A(L[602]));
Q_ASSIGN U603 ( .B(R[603]), .A(L[603]));
Q_ASSIGN U604 ( .B(R[604]), .A(L[604]));
Q_ASSIGN U605 ( .B(R[605]), .A(L[605]));
Q_ASSIGN U606 ( .B(R[606]), .A(L[606]));
Q_ASSIGN U607 ( .B(R[607]), .A(L[607]));
Q_ASSIGN U608 ( .B(R[608]), .A(L[608]));
Q_ASSIGN U609 ( .B(R[609]), .A(L[609]));
Q_ASSIGN U610 ( .B(R[610]), .A(L[610]));
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE "ixc_assign"
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE_LIB "IXCOM_TEMP_LIBRARY"
endmodule
