architecture module of tb_top is
  component kme_tb
  end component ;


begin
  kme_tb_dut : kme_tb
     ;
end module;
