ARCHITECTURE module OF ixc_assign_29 IS

BEGIN

  PROCESS --:o53
  (*)
  BEGIN
    L <= R ;
  END PROCESS ;
END module;