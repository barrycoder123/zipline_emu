
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
(* celldefine = 1 *) 
module nx_fifo_ctrl_ram_1r1w_xcm16 ( mem_wen, mem_waddr, mem_wdata, mem_ren, 
	mem_raddr, empty, full, used_slots, free_slots, rerr, rdata, 
	underflow, overflow, clk, rst_n, mem_rdata, mem_ecc_error, wen, 
	wdata, ren, clear);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output mem_wen;
output [10:0] mem_waddr;
output [70:0] mem_wdata;
output mem_ren;
output [10:0] mem_raddr;
output empty;
output full;
output [11:0] used_slots;
output [11:0] free_slots;
output rerr;
output [70:0] rdata;
output underflow;
output overflow;
input clk;
input rst_n;
input [70:0] mem_rdata;
input mem_ecc_error;
input wen;
input [70:0] wdata;
input ren;
input clear;
wire _zy_simnet_mem_wen_0_w$;
wire [0:10] _zy_simnet_mem_waddr_1_w$;
wire [0:70] _zy_simnet_mem_wdata_2_w$;
wire _zy_simnet_mem_ren_3_w$;
wire [0:10] _zy_simnet_mem_raddr_4_w$;
wire _zy_simnet_empty_5_w$;
wire _zy_simnet_full_6_w$;
wire [0:11] _zy_simnet_used_slots_7_w$;
wire [0:11] _zy_simnet_free_slots_8_w$;
wire _zy_simnet_rerr_9_w$;
wire [0:70] _zy_simnet_rdata_10_w$;
wire _zy_simnet_underflow_11_w$;
wire _zy_simnet_overflow_12_w$;
wire _zy_sva__asrtLbl279_1_reset_or;
wire _zy_sva_sf1hot_0;
wire _zyixc_port_1_0_s2hW;
wire [11:0] r_used_slots;
wire [11:0] c_used_slots;
wire [11:0] r_free_slots;
wire [11:0] c_free_slots;
wire [2:0] r_mem_ren_dly;
wire [2:0] c_mem_ren_dly;
wire [10:0] r_mem_wptr;
wire [10:0] c_mem_wptr;
wire [10:0] r_mem_rptr;
wire [10:0] c_mem_rptr;
wire r_mem_empty;
wire c_mem_empty;
wire r_mem_full;
wire c_mem_full;
wire [2:0] r_prefetch_wptr;
wire [2:0] c_prefetch_wptr;
wire [1:0] r_prefetch_rptr;
wire [1:0] c_prefetch_rptr;
wire [1:0] r_prefetch_depth;
wire [1:0] c_prefetch_depth;
wire r_prefetch_empty;
wire c_prefetch_empty;
wire r_prefetch_full;
wire c_prefetch_full;
wire prefetch_wen;
wire [2:0] prefetch_lden_bypass;
wire [2:0] prefetch_lden_mem;
`_2_ wire [2:0] _zy_sva_b0;
`_2_ wire [0:0] _zy_sva__asrtLbl279_1_1_fail;
`_2_ wire _zyixc_port_1_0_req;
`_2_ wire _zyixc_port_1_0_ack;
`_2_ wire _zyixc_port_1_0_isf;
`_2_ wire _zyixc_port_1_0_osf;
supply0 n838;
supply0 n839;
supply0 n840;
Q_BUF U0 ( .A(r_prefetch_wptr[2]), .Z(\c_mem_prefetch_wptr_dly[0][2] ));
Q_BUF U1 ( .A(r_prefetch_wptr[1]), .Z(\c_mem_prefetch_wptr_dly[0][1] ));
Q_BUF U2 ( .A(r_prefetch_wptr[0]), .Z(\c_mem_prefetch_wptr_dly[0][0] ));
Q_BUF U3 ( .A(\r_mem_prefetch_wptr_dly[0][0] ), .Z(\c_mem_prefetch_wptr_dly[1][0] ));
Q_BUF U4 ( .A(\r_mem_prefetch_wptr_dly[0][1] ), .Z(\c_mem_prefetch_wptr_dly[1][1] ));
Q_BUF U5 ( .A(\r_mem_prefetch_wptr_dly[0][2] ), .Z(\c_mem_prefetch_wptr_dly[1][2] ));
Q_BUF U6 ( .A(\r_mem_prefetch_wptr_dly[1][0] ), .Z(\c_mem_prefetch_wptr_dly[2][0] ));
Q_BUF U7 ( .A(\r_mem_prefetch_wptr_dly[1][1] ), .Z(\c_mem_prefetch_wptr_dly[2][1] ));
Q_BUF U8 ( .A(\r_mem_prefetch_wptr_dly[1][2] ), .Z(\c_mem_prefetch_wptr_dly[2][2] ));
Q_BUF U9 ( .A(n838), .Z(n1));
Q_MX03 U10 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][71] ), .A1(\r_prefetch_data[1][71] ), .A2(\r_prefetch_data[2][71] ), .Z(n2));
Q_MX03 U11 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][70] ), .A1(\r_prefetch_data[1][70] ), .A2(\r_prefetch_data[2][70] ), .Z(n3));
Q_MX03 U12 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][69] ), .A1(\r_prefetch_data[1][69] ), .A2(\r_prefetch_data[2][69] ), .Z(n4));
Q_MX03 U13 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][68] ), .A1(\r_prefetch_data[1][68] ), .A2(\r_prefetch_data[2][68] ), .Z(n5));
Q_MX03 U14 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][67] ), .A1(\r_prefetch_data[1][67] ), .A2(\r_prefetch_data[2][67] ), .Z(n6));
Q_MX03 U15 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][66] ), .A1(\r_prefetch_data[1][66] ), .A2(\r_prefetch_data[2][66] ), .Z(n7));
Q_MX03 U16 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][65] ), .A1(\r_prefetch_data[1][65] ), .A2(\r_prefetch_data[2][65] ), .Z(n8));
Q_MX03 U17 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][64] ), .A1(\r_prefetch_data[1][64] ), .A2(\r_prefetch_data[2][64] ), .Z(n9));
Q_MX03 U18 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][63] ), .A1(\r_prefetch_data[1][63] ), .A2(\r_prefetch_data[2][63] ), .Z(n10));
Q_MX03 U19 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][62] ), .A1(\r_prefetch_data[1][62] ), .A2(\r_prefetch_data[2][62] ), .Z(n11));
Q_MX03 U20 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][61] ), .A1(\r_prefetch_data[1][61] ), .A2(\r_prefetch_data[2][61] ), .Z(n12));
Q_MX03 U21 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][60] ), .A1(\r_prefetch_data[1][60] ), .A2(\r_prefetch_data[2][60] ), .Z(n13));
Q_MX03 U22 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][59] ), .A1(\r_prefetch_data[1][59] ), .A2(\r_prefetch_data[2][59] ), .Z(n14));
Q_MX03 U23 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][58] ), .A1(\r_prefetch_data[1][58] ), .A2(\r_prefetch_data[2][58] ), .Z(n15));
Q_MX03 U24 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][57] ), .A1(\r_prefetch_data[1][57] ), .A2(\r_prefetch_data[2][57] ), .Z(n16));
Q_MX03 U25 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][56] ), .A1(\r_prefetch_data[1][56] ), .A2(\r_prefetch_data[2][56] ), .Z(n17));
Q_MX03 U26 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][55] ), .A1(\r_prefetch_data[1][55] ), .A2(\r_prefetch_data[2][55] ), .Z(n18));
Q_MX03 U27 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][54] ), .A1(\r_prefetch_data[1][54] ), .A2(\r_prefetch_data[2][54] ), .Z(n19));
Q_MX03 U28 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][53] ), .A1(\r_prefetch_data[1][53] ), .A2(\r_prefetch_data[2][53] ), .Z(n20));
Q_MX03 U29 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][52] ), .A1(\r_prefetch_data[1][52] ), .A2(\r_prefetch_data[2][52] ), .Z(n21));
Q_MX03 U30 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][51] ), .A1(\r_prefetch_data[1][51] ), .A2(\r_prefetch_data[2][51] ), .Z(n22));
Q_MX03 U31 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][50] ), .A1(\r_prefetch_data[1][50] ), .A2(\r_prefetch_data[2][50] ), .Z(n23));
Q_MX03 U32 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][49] ), .A1(\r_prefetch_data[1][49] ), .A2(\r_prefetch_data[2][49] ), .Z(n24));
Q_MX03 U33 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][48] ), .A1(\r_prefetch_data[1][48] ), .A2(\r_prefetch_data[2][48] ), .Z(n25));
Q_MX03 U34 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][47] ), .A1(\r_prefetch_data[1][47] ), .A2(\r_prefetch_data[2][47] ), .Z(n26));
Q_MX03 U35 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][46] ), .A1(\r_prefetch_data[1][46] ), .A2(\r_prefetch_data[2][46] ), .Z(n27));
Q_MX03 U36 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][45] ), .A1(\r_prefetch_data[1][45] ), .A2(\r_prefetch_data[2][45] ), .Z(n28));
Q_MX03 U37 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][44] ), .A1(\r_prefetch_data[1][44] ), .A2(\r_prefetch_data[2][44] ), .Z(n29));
Q_MX03 U38 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][43] ), .A1(\r_prefetch_data[1][43] ), .A2(\r_prefetch_data[2][43] ), .Z(n30));
Q_MX03 U39 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][42] ), .A1(\r_prefetch_data[1][42] ), .A2(\r_prefetch_data[2][42] ), .Z(n31));
Q_MX03 U40 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][41] ), .A1(\r_prefetch_data[1][41] ), .A2(\r_prefetch_data[2][41] ), .Z(n32));
Q_MX03 U41 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][40] ), .A1(\r_prefetch_data[1][40] ), .A2(\r_prefetch_data[2][40] ), .Z(n33));
Q_MX03 U42 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][39] ), .A1(\r_prefetch_data[1][39] ), .A2(\r_prefetch_data[2][39] ), .Z(n34));
Q_MX03 U43 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][38] ), .A1(\r_prefetch_data[1][38] ), .A2(\r_prefetch_data[2][38] ), .Z(n35));
Q_MX03 U44 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][37] ), .A1(\r_prefetch_data[1][37] ), .A2(\r_prefetch_data[2][37] ), .Z(n36));
Q_MX03 U45 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][36] ), .A1(\r_prefetch_data[1][36] ), .A2(\r_prefetch_data[2][36] ), .Z(n37));
Q_MX03 U46 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][35] ), .A1(\r_prefetch_data[1][35] ), .A2(\r_prefetch_data[2][35] ), .Z(n38));
Q_MX03 U47 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][34] ), .A1(\r_prefetch_data[1][34] ), .A2(\r_prefetch_data[2][34] ), .Z(n39));
Q_MX03 U48 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][33] ), .A1(\r_prefetch_data[1][33] ), .A2(\r_prefetch_data[2][33] ), .Z(n40));
Q_MX03 U49 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][32] ), .A1(\r_prefetch_data[1][32] ), .A2(\r_prefetch_data[2][32] ), .Z(n41));
Q_MX03 U50 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][31] ), .A1(\r_prefetch_data[1][31] ), .A2(\r_prefetch_data[2][31] ), .Z(n42));
Q_MX03 U51 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][30] ), .A1(\r_prefetch_data[1][30] ), .A2(\r_prefetch_data[2][30] ), .Z(n43));
Q_MX03 U52 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][29] ), .A1(\r_prefetch_data[1][29] ), .A2(\r_prefetch_data[2][29] ), .Z(n44));
Q_MX03 U53 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][28] ), .A1(\r_prefetch_data[1][28] ), .A2(\r_prefetch_data[2][28] ), .Z(n45));
Q_MX03 U54 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][27] ), .A1(\r_prefetch_data[1][27] ), .A2(\r_prefetch_data[2][27] ), .Z(n46));
Q_MX03 U55 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][26] ), .A1(\r_prefetch_data[1][26] ), .A2(\r_prefetch_data[2][26] ), .Z(n47));
Q_MX03 U56 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][25] ), .A1(\r_prefetch_data[1][25] ), .A2(\r_prefetch_data[2][25] ), .Z(n48));
Q_MX03 U57 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][24] ), .A1(\r_prefetch_data[1][24] ), .A2(\r_prefetch_data[2][24] ), .Z(n49));
Q_MX03 U58 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][23] ), .A1(\r_prefetch_data[1][23] ), .A2(\r_prefetch_data[2][23] ), .Z(n50));
Q_MX03 U59 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][22] ), .A1(\r_prefetch_data[1][22] ), .A2(\r_prefetch_data[2][22] ), .Z(n51));
Q_MX03 U60 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][21] ), .A1(\r_prefetch_data[1][21] ), .A2(\r_prefetch_data[2][21] ), .Z(n52));
Q_MX03 U61 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][20] ), .A1(\r_prefetch_data[1][20] ), .A2(\r_prefetch_data[2][20] ), .Z(n53));
Q_MX03 U62 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][19] ), .A1(\r_prefetch_data[1][19] ), .A2(\r_prefetch_data[2][19] ), .Z(n54));
Q_MX03 U63 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][18] ), .A1(\r_prefetch_data[1][18] ), .A2(\r_prefetch_data[2][18] ), .Z(n55));
Q_MX03 U64 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][17] ), .A1(\r_prefetch_data[1][17] ), .A2(\r_prefetch_data[2][17] ), .Z(n56));
Q_MX03 U65 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][16] ), .A1(\r_prefetch_data[1][16] ), .A2(\r_prefetch_data[2][16] ), .Z(n57));
Q_MX03 U66 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][15] ), .A1(\r_prefetch_data[1][15] ), .A2(\r_prefetch_data[2][15] ), .Z(n58));
Q_MX03 U67 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][14] ), .A1(\r_prefetch_data[1][14] ), .A2(\r_prefetch_data[2][14] ), .Z(n59));
Q_MX03 U68 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][13] ), .A1(\r_prefetch_data[1][13] ), .A2(\r_prefetch_data[2][13] ), .Z(n60));
Q_MX03 U69 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][12] ), .A1(\r_prefetch_data[1][12] ), .A2(\r_prefetch_data[2][12] ), .Z(n61));
Q_MX03 U70 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][11] ), .A1(\r_prefetch_data[1][11] ), .A2(\r_prefetch_data[2][11] ), .Z(n62));
Q_MX03 U71 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][10] ), .A1(\r_prefetch_data[1][10] ), .A2(\r_prefetch_data[2][10] ), .Z(n63));
Q_MX03 U72 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][9] ), .A1(\r_prefetch_data[1][9] ), .A2(\r_prefetch_data[2][9] ), .Z(n64));
Q_MX03 U73 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][8] ), .A1(\r_prefetch_data[1][8] ), .A2(\r_prefetch_data[2][8] ), .Z(n65));
Q_MX03 U74 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][7] ), .A1(\r_prefetch_data[1][7] ), .A2(\r_prefetch_data[2][7] ), .Z(n66));
Q_MX03 U75 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][6] ), .A1(\r_prefetch_data[1][6] ), .A2(\r_prefetch_data[2][6] ), .Z(n67));
Q_MX03 U76 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][5] ), .A1(\r_prefetch_data[1][5] ), .A2(\r_prefetch_data[2][5] ), .Z(n68));
Q_MX03 U77 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][4] ), .A1(\r_prefetch_data[1][4] ), .A2(\r_prefetch_data[2][4] ), .Z(n69));
Q_MX03 U78 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][3] ), .A1(\r_prefetch_data[1][3] ), .A2(\r_prefetch_data[2][3] ), .Z(n70));
Q_MX03 U79 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][2] ), .A1(\r_prefetch_data[1][2] ), .A2(\r_prefetch_data[2][2] ), .Z(n71));
Q_MX03 U80 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][1] ), .A1(\r_prefetch_data[1][1] ), .A2(\r_prefetch_data[2][1] ), .Z(n72));
Q_MX03 U81 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(\r_prefetch_data[0][0] ), .A1(\r_prefetch_data[1][0] ), .A2(\r_prefetch_data[2][0] ), .Z(n73));
Q_FDP0 \r_mem_prefetch_wptr_dly_REG[2][2] ( .CK(clk), .D(\c_mem_prefetch_wptr_dly[2][2] ), .Q(\r_mem_prefetch_wptr_dly[2][2] ), .QN( ));
Q_FDP0 \r_mem_prefetch_wptr_dly_REG[2][1] ( .CK(clk), .D(\c_mem_prefetch_wptr_dly[2][1] ), .Q(\r_mem_prefetch_wptr_dly[2][1] ), .QN( ));
Q_FDP0 \r_mem_prefetch_wptr_dly_REG[2][0] ( .CK(clk), .D(\c_mem_prefetch_wptr_dly[2][0] ), .Q(\r_mem_prefetch_wptr_dly[2][0] ), .QN( ));
Q_FDP0 \r_mem_prefetch_wptr_dly_REG[1][2] ( .CK(clk), .D(\c_mem_prefetch_wptr_dly[1][2] ), .Q(\r_mem_prefetch_wptr_dly[1][2] ), .QN( ));
Q_FDP0 \r_mem_prefetch_wptr_dly_REG[1][1] ( .CK(clk), .D(\c_mem_prefetch_wptr_dly[1][1] ), .Q(\r_mem_prefetch_wptr_dly[1][1] ), .QN( ));
Q_FDP0 \r_mem_prefetch_wptr_dly_REG[1][0] ( .CK(clk), .D(\c_mem_prefetch_wptr_dly[1][0] ), .Q(\r_mem_prefetch_wptr_dly[1][0] ), .QN( ));
Q_FDP0 \r_mem_prefetch_wptr_dly_REG[0][2] ( .CK(clk), .D(\c_mem_prefetch_wptr_dly[0][2] ), .Q(\r_mem_prefetch_wptr_dly[0][2] ), .QN( ));
Q_FDP0 \r_mem_prefetch_wptr_dly_REG[0][1] ( .CK(clk), .D(\c_mem_prefetch_wptr_dly[0][1] ), .Q(\r_mem_prefetch_wptr_dly[0][1] ), .QN( ));
Q_FDP0 \r_mem_prefetch_wptr_dly_REG[0][0] ( .CK(clk), .D(\c_mem_prefetch_wptr_dly[0][0] ), .Q(\r_mem_prefetch_wptr_dly[0][0] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][71] ( .CK(clk), .D(\c_prefetch_data[2][71] ), .Q(\r_prefetch_data[2][71] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][70] ( .CK(clk), .D(\c_prefetch_data[2][70] ), .Q(\r_prefetch_data[2][70] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][69] ( .CK(clk), .D(\c_prefetch_data[2][69] ), .Q(\r_prefetch_data[2][69] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][68] ( .CK(clk), .D(\c_prefetch_data[2][68] ), .Q(\r_prefetch_data[2][68] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][67] ( .CK(clk), .D(\c_prefetch_data[2][67] ), .Q(\r_prefetch_data[2][67] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][66] ( .CK(clk), .D(\c_prefetch_data[2][66] ), .Q(\r_prefetch_data[2][66] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][65] ( .CK(clk), .D(\c_prefetch_data[2][65] ), .Q(\r_prefetch_data[2][65] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][64] ( .CK(clk), .D(\c_prefetch_data[2][64] ), .Q(\r_prefetch_data[2][64] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][63] ( .CK(clk), .D(\c_prefetch_data[2][63] ), .Q(\r_prefetch_data[2][63] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][62] ( .CK(clk), .D(\c_prefetch_data[2][62] ), .Q(\r_prefetch_data[2][62] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][61] ( .CK(clk), .D(\c_prefetch_data[2][61] ), .Q(\r_prefetch_data[2][61] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][60] ( .CK(clk), .D(\c_prefetch_data[2][60] ), .Q(\r_prefetch_data[2][60] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][59] ( .CK(clk), .D(\c_prefetch_data[2][59] ), .Q(\r_prefetch_data[2][59] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][58] ( .CK(clk), .D(\c_prefetch_data[2][58] ), .Q(\r_prefetch_data[2][58] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][57] ( .CK(clk), .D(\c_prefetch_data[2][57] ), .Q(\r_prefetch_data[2][57] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][56] ( .CK(clk), .D(\c_prefetch_data[2][56] ), .Q(\r_prefetch_data[2][56] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][55] ( .CK(clk), .D(\c_prefetch_data[2][55] ), .Q(\r_prefetch_data[2][55] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][54] ( .CK(clk), .D(\c_prefetch_data[2][54] ), .Q(\r_prefetch_data[2][54] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][53] ( .CK(clk), .D(\c_prefetch_data[2][53] ), .Q(\r_prefetch_data[2][53] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][52] ( .CK(clk), .D(\c_prefetch_data[2][52] ), .Q(\r_prefetch_data[2][52] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][51] ( .CK(clk), .D(\c_prefetch_data[2][51] ), .Q(\r_prefetch_data[2][51] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][50] ( .CK(clk), .D(\c_prefetch_data[2][50] ), .Q(\r_prefetch_data[2][50] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][49] ( .CK(clk), .D(\c_prefetch_data[2][49] ), .Q(\r_prefetch_data[2][49] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][48] ( .CK(clk), .D(\c_prefetch_data[2][48] ), .Q(\r_prefetch_data[2][48] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][47] ( .CK(clk), .D(\c_prefetch_data[2][47] ), .Q(\r_prefetch_data[2][47] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][46] ( .CK(clk), .D(\c_prefetch_data[2][46] ), .Q(\r_prefetch_data[2][46] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][45] ( .CK(clk), .D(\c_prefetch_data[2][45] ), .Q(\r_prefetch_data[2][45] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][44] ( .CK(clk), .D(\c_prefetch_data[2][44] ), .Q(\r_prefetch_data[2][44] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][43] ( .CK(clk), .D(\c_prefetch_data[2][43] ), .Q(\r_prefetch_data[2][43] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][42] ( .CK(clk), .D(\c_prefetch_data[2][42] ), .Q(\r_prefetch_data[2][42] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][41] ( .CK(clk), .D(\c_prefetch_data[2][41] ), .Q(\r_prefetch_data[2][41] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][40] ( .CK(clk), .D(\c_prefetch_data[2][40] ), .Q(\r_prefetch_data[2][40] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][39] ( .CK(clk), .D(\c_prefetch_data[2][39] ), .Q(\r_prefetch_data[2][39] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][38] ( .CK(clk), .D(\c_prefetch_data[2][38] ), .Q(\r_prefetch_data[2][38] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][37] ( .CK(clk), .D(\c_prefetch_data[2][37] ), .Q(\r_prefetch_data[2][37] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][36] ( .CK(clk), .D(\c_prefetch_data[2][36] ), .Q(\r_prefetch_data[2][36] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][35] ( .CK(clk), .D(\c_prefetch_data[2][35] ), .Q(\r_prefetch_data[2][35] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][34] ( .CK(clk), .D(\c_prefetch_data[2][34] ), .Q(\r_prefetch_data[2][34] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][33] ( .CK(clk), .D(\c_prefetch_data[2][33] ), .Q(\r_prefetch_data[2][33] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][32] ( .CK(clk), .D(\c_prefetch_data[2][32] ), .Q(\r_prefetch_data[2][32] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][31] ( .CK(clk), .D(\c_prefetch_data[2][31] ), .Q(\r_prefetch_data[2][31] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][30] ( .CK(clk), .D(\c_prefetch_data[2][30] ), .Q(\r_prefetch_data[2][30] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][29] ( .CK(clk), .D(\c_prefetch_data[2][29] ), .Q(\r_prefetch_data[2][29] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][28] ( .CK(clk), .D(\c_prefetch_data[2][28] ), .Q(\r_prefetch_data[2][28] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][27] ( .CK(clk), .D(\c_prefetch_data[2][27] ), .Q(\r_prefetch_data[2][27] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][26] ( .CK(clk), .D(\c_prefetch_data[2][26] ), .Q(\r_prefetch_data[2][26] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][25] ( .CK(clk), .D(\c_prefetch_data[2][25] ), .Q(\r_prefetch_data[2][25] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][24] ( .CK(clk), .D(\c_prefetch_data[2][24] ), .Q(\r_prefetch_data[2][24] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][23] ( .CK(clk), .D(\c_prefetch_data[2][23] ), .Q(\r_prefetch_data[2][23] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][22] ( .CK(clk), .D(\c_prefetch_data[2][22] ), .Q(\r_prefetch_data[2][22] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][21] ( .CK(clk), .D(\c_prefetch_data[2][21] ), .Q(\r_prefetch_data[2][21] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][20] ( .CK(clk), .D(\c_prefetch_data[2][20] ), .Q(\r_prefetch_data[2][20] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][19] ( .CK(clk), .D(\c_prefetch_data[2][19] ), .Q(\r_prefetch_data[2][19] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][18] ( .CK(clk), .D(\c_prefetch_data[2][18] ), .Q(\r_prefetch_data[2][18] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][17] ( .CK(clk), .D(\c_prefetch_data[2][17] ), .Q(\r_prefetch_data[2][17] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][16] ( .CK(clk), .D(\c_prefetch_data[2][16] ), .Q(\r_prefetch_data[2][16] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][15] ( .CK(clk), .D(\c_prefetch_data[2][15] ), .Q(\r_prefetch_data[2][15] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][14] ( .CK(clk), .D(\c_prefetch_data[2][14] ), .Q(\r_prefetch_data[2][14] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][13] ( .CK(clk), .D(\c_prefetch_data[2][13] ), .Q(\r_prefetch_data[2][13] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][12] ( .CK(clk), .D(\c_prefetch_data[2][12] ), .Q(\r_prefetch_data[2][12] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][11] ( .CK(clk), .D(\c_prefetch_data[2][11] ), .Q(\r_prefetch_data[2][11] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][10] ( .CK(clk), .D(\c_prefetch_data[2][10] ), .Q(\r_prefetch_data[2][10] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][9] ( .CK(clk), .D(\c_prefetch_data[2][9] ), .Q(\r_prefetch_data[2][9] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][8] ( .CK(clk), .D(\c_prefetch_data[2][8] ), .Q(\r_prefetch_data[2][8] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][7] ( .CK(clk), .D(\c_prefetch_data[2][7] ), .Q(\r_prefetch_data[2][7] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][6] ( .CK(clk), .D(\c_prefetch_data[2][6] ), .Q(\r_prefetch_data[2][6] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][5] ( .CK(clk), .D(\c_prefetch_data[2][5] ), .Q(\r_prefetch_data[2][5] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][4] ( .CK(clk), .D(\c_prefetch_data[2][4] ), .Q(\r_prefetch_data[2][4] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][3] ( .CK(clk), .D(\c_prefetch_data[2][3] ), .Q(\r_prefetch_data[2][3] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][2] ( .CK(clk), .D(\c_prefetch_data[2][2] ), .Q(\r_prefetch_data[2][2] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][1] ( .CK(clk), .D(\c_prefetch_data[2][1] ), .Q(\r_prefetch_data[2][1] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[2][0] ( .CK(clk), .D(\c_prefetch_data[2][0] ), .Q(\r_prefetch_data[2][0] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][71] ( .CK(clk), .D(\c_prefetch_data[1][71] ), .Q(\r_prefetch_data[1][71] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][70] ( .CK(clk), .D(\c_prefetch_data[1][70] ), .Q(\r_prefetch_data[1][70] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][69] ( .CK(clk), .D(\c_prefetch_data[1][69] ), .Q(\r_prefetch_data[1][69] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][68] ( .CK(clk), .D(\c_prefetch_data[1][68] ), .Q(\r_prefetch_data[1][68] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][67] ( .CK(clk), .D(\c_prefetch_data[1][67] ), .Q(\r_prefetch_data[1][67] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][66] ( .CK(clk), .D(\c_prefetch_data[1][66] ), .Q(\r_prefetch_data[1][66] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][65] ( .CK(clk), .D(\c_prefetch_data[1][65] ), .Q(\r_prefetch_data[1][65] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][64] ( .CK(clk), .D(\c_prefetch_data[1][64] ), .Q(\r_prefetch_data[1][64] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][63] ( .CK(clk), .D(\c_prefetch_data[1][63] ), .Q(\r_prefetch_data[1][63] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][62] ( .CK(clk), .D(\c_prefetch_data[1][62] ), .Q(\r_prefetch_data[1][62] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][61] ( .CK(clk), .D(\c_prefetch_data[1][61] ), .Q(\r_prefetch_data[1][61] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][60] ( .CK(clk), .D(\c_prefetch_data[1][60] ), .Q(\r_prefetch_data[1][60] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][59] ( .CK(clk), .D(\c_prefetch_data[1][59] ), .Q(\r_prefetch_data[1][59] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][58] ( .CK(clk), .D(\c_prefetch_data[1][58] ), .Q(\r_prefetch_data[1][58] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][57] ( .CK(clk), .D(\c_prefetch_data[1][57] ), .Q(\r_prefetch_data[1][57] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][56] ( .CK(clk), .D(\c_prefetch_data[1][56] ), .Q(\r_prefetch_data[1][56] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][55] ( .CK(clk), .D(\c_prefetch_data[1][55] ), .Q(\r_prefetch_data[1][55] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][54] ( .CK(clk), .D(\c_prefetch_data[1][54] ), .Q(\r_prefetch_data[1][54] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][53] ( .CK(clk), .D(\c_prefetch_data[1][53] ), .Q(\r_prefetch_data[1][53] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][52] ( .CK(clk), .D(\c_prefetch_data[1][52] ), .Q(\r_prefetch_data[1][52] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][51] ( .CK(clk), .D(\c_prefetch_data[1][51] ), .Q(\r_prefetch_data[1][51] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][50] ( .CK(clk), .D(\c_prefetch_data[1][50] ), .Q(\r_prefetch_data[1][50] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][49] ( .CK(clk), .D(\c_prefetch_data[1][49] ), .Q(\r_prefetch_data[1][49] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][48] ( .CK(clk), .D(\c_prefetch_data[1][48] ), .Q(\r_prefetch_data[1][48] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][47] ( .CK(clk), .D(\c_prefetch_data[1][47] ), .Q(\r_prefetch_data[1][47] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][46] ( .CK(clk), .D(\c_prefetch_data[1][46] ), .Q(\r_prefetch_data[1][46] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][45] ( .CK(clk), .D(\c_prefetch_data[1][45] ), .Q(\r_prefetch_data[1][45] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][44] ( .CK(clk), .D(\c_prefetch_data[1][44] ), .Q(\r_prefetch_data[1][44] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][43] ( .CK(clk), .D(\c_prefetch_data[1][43] ), .Q(\r_prefetch_data[1][43] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][42] ( .CK(clk), .D(\c_prefetch_data[1][42] ), .Q(\r_prefetch_data[1][42] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][41] ( .CK(clk), .D(\c_prefetch_data[1][41] ), .Q(\r_prefetch_data[1][41] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][40] ( .CK(clk), .D(\c_prefetch_data[1][40] ), .Q(\r_prefetch_data[1][40] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][39] ( .CK(clk), .D(\c_prefetch_data[1][39] ), .Q(\r_prefetch_data[1][39] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][38] ( .CK(clk), .D(\c_prefetch_data[1][38] ), .Q(\r_prefetch_data[1][38] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][37] ( .CK(clk), .D(\c_prefetch_data[1][37] ), .Q(\r_prefetch_data[1][37] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][36] ( .CK(clk), .D(\c_prefetch_data[1][36] ), .Q(\r_prefetch_data[1][36] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][35] ( .CK(clk), .D(\c_prefetch_data[1][35] ), .Q(\r_prefetch_data[1][35] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][34] ( .CK(clk), .D(\c_prefetch_data[1][34] ), .Q(\r_prefetch_data[1][34] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][33] ( .CK(clk), .D(\c_prefetch_data[1][33] ), .Q(\r_prefetch_data[1][33] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][32] ( .CK(clk), .D(\c_prefetch_data[1][32] ), .Q(\r_prefetch_data[1][32] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][31] ( .CK(clk), .D(\c_prefetch_data[1][31] ), .Q(\r_prefetch_data[1][31] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][30] ( .CK(clk), .D(\c_prefetch_data[1][30] ), .Q(\r_prefetch_data[1][30] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][29] ( .CK(clk), .D(\c_prefetch_data[1][29] ), .Q(\r_prefetch_data[1][29] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][28] ( .CK(clk), .D(\c_prefetch_data[1][28] ), .Q(\r_prefetch_data[1][28] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][27] ( .CK(clk), .D(\c_prefetch_data[1][27] ), .Q(\r_prefetch_data[1][27] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][26] ( .CK(clk), .D(\c_prefetch_data[1][26] ), .Q(\r_prefetch_data[1][26] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][25] ( .CK(clk), .D(\c_prefetch_data[1][25] ), .Q(\r_prefetch_data[1][25] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][24] ( .CK(clk), .D(\c_prefetch_data[1][24] ), .Q(\r_prefetch_data[1][24] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][23] ( .CK(clk), .D(\c_prefetch_data[1][23] ), .Q(\r_prefetch_data[1][23] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][22] ( .CK(clk), .D(\c_prefetch_data[1][22] ), .Q(\r_prefetch_data[1][22] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][21] ( .CK(clk), .D(\c_prefetch_data[1][21] ), .Q(\r_prefetch_data[1][21] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][20] ( .CK(clk), .D(\c_prefetch_data[1][20] ), .Q(\r_prefetch_data[1][20] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][19] ( .CK(clk), .D(\c_prefetch_data[1][19] ), .Q(\r_prefetch_data[1][19] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][18] ( .CK(clk), .D(\c_prefetch_data[1][18] ), .Q(\r_prefetch_data[1][18] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][17] ( .CK(clk), .D(\c_prefetch_data[1][17] ), .Q(\r_prefetch_data[1][17] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][16] ( .CK(clk), .D(\c_prefetch_data[1][16] ), .Q(\r_prefetch_data[1][16] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][15] ( .CK(clk), .D(\c_prefetch_data[1][15] ), .Q(\r_prefetch_data[1][15] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][14] ( .CK(clk), .D(\c_prefetch_data[1][14] ), .Q(\r_prefetch_data[1][14] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][13] ( .CK(clk), .D(\c_prefetch_data[1][13] ), .Q(\r_prefetch_data[1][13] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][12] ( .CK(clk), .D(\c_prefetch_data[1][12] ), .Q(\r_prefetch_data[1][12] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][11] ( .CK(clk), .D(\c_prefetch_data[1][11] ), .Q(\r_prefetch_data[1][11] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][10] ( .CK(clk), .D(\c_prefetch_data[1][10] ), .Q(\r_prefetch_data[1][10] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][9] ( .CK(clk), .D(\c_prefetch_data[1][9] ), .Q(\r_prefetch_data[1][9] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][8] ( .CK(clk), .D(\c_prefetch_data[1][8] ), .Q(\r_prefetch_data[1][8] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][7] ( .CK(clk), .D(\c_prefetch_data[1][7] ), .Q(\r_prefetch_data[1][7] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][6] ( .CK(clk), .D(\c_prefetch_data[1][6] ), .Q(\r_prefetch_data[1][6] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][5] ( .CK(clk), .D(\c_prefetch_data[1][5] ), .Q(\r_prefetch_data[1][5] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][4] ( .CK(clk), .D(\c_prefetch_data[1][4] ), .Q(\r_prefetch_data[1][4] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][3] ( .CK(clk), .D(\c_prefetch_data[1][3] ), .Q(\r_prefetch_data[1][3] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][2] ( .CK(clk), .D(\c_prefetch_data[1][2] ), .Q(\r_prefetch_data[1][2] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][1] ( .CK(clk), .D(\c_prefetch_data[1][1] ), .Q(\r_prefetch_data[1][1] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[1][0] ( .CK(clk), .D(\c_prefetch_data[1][0] ), .Q(\r_prefetch_data[1][0] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][71] ( .CK(clk), .D(\c_prefetch_data[0][71] ), .Q(\r_prefetch_data[0][71] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][70] ( .CK(clk), .D(\c_prefetch_data[0][70] ), .Q(\r_prefetch_data[0][70] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][69] ( .CK(clk), .D(\c_prefetch_data[0][69] ), .Q(\r_prefetch_data[0][69] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][68] ( .CK(clk), .D(\c_prefetch_data[0][68] ), .Q(\r_prefetch_data[0][68] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][67] ( .CK(clk), .D(\c_prefetch_data[0][67] ), .Q(\r_prefetch_data[0][67] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][66] ( .CK(clk), .D(\c_prefetch_data[0][66] ), .Q(\r_prefetch_data[0][66] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][65] ( .CK(clk), .D(\c_prefetch_data[0][65] ), .Q(\r_prefetch_data[0][65] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][64] ( .CK(clk), .D(\c_prefetch_data[0][64] ), .Q(\r_prefetch_data[0][64] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][63] ( .CK(clk), .D(\c_prefetch_data[0][63] ), .Q(\r_prefetch_data[0][63] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][62] ( .CK(clk), .D(\c_prefetch_data[0][62] ), .Q(\r_prefetch_data[0][62] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][61] ( .CK(clk), .D(\c_prefetch_data[0][61] ), .Q(\r_prefetch_data[0][61] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][60] ( .CK(clk), .D(\c_prefetch_data[0][60] ), .Q(\r_prefetch_data[0][60] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][59] ( .CK(clk), .D(\c_prefetch_data[0][59] ), .Q(\r_prefetch_data[0][59] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][58] ( .CK(clk), .D(\c_prefetch_data[0][58] ), .Q(\r_prefetch_data[0][58] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][57] ( .CK(clk), .D(\c_prefetch_data[0][57] ), .Q(\r_prefetch_data[0][57] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][56] ( .CK(clk), .D(\c_prefetch_data[0][56] ), .Q(\r_prefetch_data[0][56] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][55] ( .CK(clk), .D(\c_prefetch_data[0][55] ), .Q(\r_prefetch_data[0][55] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][54] ( .CK(clk), .D(\c_prefetch_data[0][54] ), .Q(\r_prefetch_data[0][54] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][53] ( .CK(clk), .D(\c_prefetch_data[0][53] ), .Q(\r_prefetch_data[0][53] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][52] ( .CK(clk), .D(\c_prefetch_data[0][52] ), .Q(\r_prefetch_data[0][52] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][51] ( .CK(clk), .D(\c_prefetch_data[0][51] ), .Q(\r_prefetch_data[0][51] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][50] ( .CK(clk), .D(\c_prefetch_data[0][50] ), .Q(\r_prefetch_data[0][50] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][49] ( .CK(clk), .D(\c_prefetch_data[0][49] ), .Q(\r_prefetch_data[0][49] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][48] ( .CK(clk), .D(\c_prefetch_data[0][48] ), .Q(\r_prefetch_data[0][48] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][47] ( .CK(clk), .D(\c_prefetch_data[0][47] ), .Q(\r_prefetch_data[0][47] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][46] ( .CK(clk), .D(\c_prefetch_data[0][46] ), .Q(\r_prefetch_data[0][46] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][45] ( .CK(clk), .D(\c_prefetch_data[0][45] ), .Q(\r_prefetch_data[0][45] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][44] ( .CK(clk), .D(\c_prefetch_data[0][44] ), .Q(\r_prefetch_data[0][44] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][43] ( .CK(clk), .D(\c_prefetch_data[0][43] ), .Q(\r_prefetch_data[0][43] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][42] ( .CK(clk), .D(\c_prefetch_data[0][42] ), .Q(\r_prefetch_data[0][42] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][41] ( .CK(clk), .D(\c_prefetch_data[0][41] ), .Q(\r_prefetch_data[0][41] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][40] ( .CK(clk), .D(\c_prefetch_data[0][40] ), .Q(\r_prefetch_data[0][40] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][39] ( .CK(clk), .D(\c_prefetch_data[0][39] ), .Q(\r_prefetch_data[0][39] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][38] ( .CK(clk), .D(\c_prefetch_data[0][38] ), .Q(\r_prefetch_data[0][38] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][37] ( .CK(clk), .D(\c_prefetch_data[0][37] ), .Q(\r_prefetch_data[0][37] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][36] ( .CK(clk), .D(\c_prefetch_data[0][36] ), .Q(\r_prefetch_data[0][36] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][35] ( .CK(clk), .D(\c_prefetch_data[0][35] ), .Q(\r_prefetch_data[0][35] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][34] ( .CK(clk), .D(\c_prefetch_data[0][34] ), .Q(\r_prefetch_data[0][34] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][33] ( .CK(clk), .D(\c_prefetch_data[0][33] ), .Q(\r_prefetch_data[0][33] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][32] ( .CK(clk), .D(\c_prefetch_data[0][32] ), .Q(\r_prefetch_data[0][32] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][31] ( .CK(clk), .D(\c_prefetch_data[0][31] ), .Q(\r_prefetch_data[0][31] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][30] ( .CK(clk), .D(\c_prefetch_data[0][30] ), .Q(\r_prefetch_data[0][30] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][29] ( .CK(clk), .D(\c_prefetch_data[0][29] ), .Q(\r_prefetch_data[0][29] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][28] ( .CK(clk), .D(\c_prefetch_data[0][28] ), .Q(\r_prefetch_data[0][28] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][27] ( .CK(clk), .D(\c_prefetch_data[0][27] ), .Q(\r_prefetch_data[0][27] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][26] ( .CK(clk), .D(\c_prefetch_data[0][26] ), .Q(\r_prefetch_data[0][26] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][25] ( .CK(clk), .D(\c_prefetch_data[0][25] ), .Q(\r_prefetch_data[0][25] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][24] ( .CK(clk), .D(\c_prefetch_data[0][24] ), .Q(\r_prefetch_data[0][24] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][23] ( .CK(clk), .D(\c_prefetch_data[0][23] ), .Q(\r_prefetch_data[0][23] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][22] ( .CK(clk), .D(\c_prefetch_data[0][22] ), .Q(\r_prefetch_data[0][22] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][21] ( .CK(clk), .D(\c_prefetch_data[0][21] ), .Q(\r_prefetch_data[0][21] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][20] ( .CK(clk), .D(\c_prefetch_data[0][20] ), .Q(\r_prefetch_data[0][20] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][19] ( .CK(clk), .D(\c_prefetch_data[0][19] ), .Q(\r_prefetch_data[0][19] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][18] ( .CK(clk), .D(\c_prefetch_data[0][18] ), .Q(\r_prefetch_data[0][18] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][17] ( .CK(clk), .D(\c_prefetch_data[0][17] ), .Q(\r_prefetch_data[0][17] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][16] ( .CK(clk), .D(\c_prefetch_data[0][16] ), .Q(\r_prefetch_data[0][16] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][15] ( .CK(clk), .D(\c_prefetch_data[0][15] ), .Q(\r_prefetch_data[0][15] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][14] ( .CK(clk), .D(\c_prefetch_data[0][14] ), .Q(\r_prefetch_data[0][14] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][13] ( .CK(clk), .D(\c_prefetch_data[0][13] ), .Q(\r_prefetch_data[0][13] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][12] ( .CK(clk), .D(\c_prefetch_data[0][12] ), .Q(\r_prefetch_data[0][12] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][11] ( .CK(clk), .D(\c_prefetch_data[0][11] ), .Q(\r_prefetch_data[0][11] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][10] ( .CK(clk), .D(\c_prefetch_data[0][10] ), .Q(\r_prefetch_data[0][10] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][9] ( .CK(clk), .D(\c_prefetch_data[0][9] ), .Q(\r_prefetch_data[0][9] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][8] ( .CK(clk), .D(\c_prefetch_data[0][8] ), .Q(\r_prefetch_data[0][8] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][7] ( .CK(clk), .D(\c_prefetch_data[0][7] ), .Q(\r_prefetch_data[0][7] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][6] ( .CK(clk), .D(\c_prefetch_data[0][6] ), .Q(\r_prefetch_data[0][6] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][5] ( .CK(clk), .D(\c_prefetch_data[0][5] ), .Q(\r_prefetch_data[0][5] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][4] ( .CK(clk), .D(\c_prefetch_data[0][4] ), .Q(\r_prefetch_data[0][4] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][3] ( .CK(clk), .D(\c_prefetch_data[0][3] ), .Q(\r_prefetch_data[0][3] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][2] ( .CK(clk), .D(\c_prefetch_data[0][2] ), .Q(\r_prefetch_data[0][2] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][1] ( .CK(clk), .D(\c_prefetch_data[0][1] ), .Q(\r_prefetch_data[0][1] ), .QN( ));
Q_FDP0 \r_prefetch_data_REG[0][0] ( .CK(clk), .D(\c_prefetch_data[0][0] ), .Q(\r_prefetch_data[0][0] ), .QN( ));
Q_FDP1 \r_mem_ren_dly_REG[2] ( .CK(clk), .R(rst_n), .D(c_mem_ren_dly[2]), .Q(r_mem_ren_dly[2]), .QN( ));
Q_FDP1 \r_mem_ren_dly_REG[1] ( .CK(clk), .R(rst_n), .D(c_mem_ren_dly[1]), .Q(r_mem_ren_dly[1]), .QN( ));
Q_FDP1 \r_mem_ren_dly_REG[0] ( .CK(clk), .R(rst_n), .D(c_mem_ren_dly[0]), .Q(r_mem_ren_dly[0]), .QN( ));
Q_FDP2 r_mem_empty_REG  ( .CK(clk), .S(rst_n), .D(c_mem_empty), .Q(r_mem_empty), .QN( ));
Q_FDP1 r_mem_full_REG  ( .CK(clk), .R(rst_n), .D(c_mem_full), .Q(r_mem_full), .QN(n118));
Q_FDP1 \r_mem_wptr_REG[10] ( .CK(clk), .R(rst_n), .D(c_mem_wptr[10]), .Q(r_mem_wptr[10]), .QN( ));
Q_FDP1 \r_mem_wptr_REG[9] ( .CK(clk), .R(rst_n), .D(c_mem_wptr[9]), .Q(r_mem_wptr[9]), .QN( ));
Q_FDP1 \r_mem_wptr_REG[8] ( .CK(clk), .R(rst_n), .D(c_mem_wptr[8]), .Q(r_mem_wptr[8]), .QN( ));
Q_FDP1 \r_mem_wptr_REG[7] ( .CK(clk), .R(rst_n), .D(c_mem_wptr[7]), .Q(r_mem_wptr[7]), .QN( ));
Q_FDP1 \r_mem_wptr_REG[6] ( .CK(clk), .R(rst_n), .D(c_mem_wptr[6]), .Q(r_mem_wptr[6]), .QN( ));
Q_FDP1 \r_mem_wptr_REG[5] ( .CK(clk), .R(rst_n), .D(c_mem_wptr[5]), .Q(r_mem_wptr[5]), .QN( ));
Q_FDP1 \r_mem_wptr_REG[4] ( .CK(clk), .R(rst_n), .D(c_mem_wptr[4]), .Q(r_mem_wptr[4]), .QN( ));
Q_FDP1 \r_mem_wptr_REG[3] ( .CK(clk), .R(rst_n), .D(c_mem_wptr[3]), .Q(r_mem_wptr[3]), .QN( ));
Q_FDP1 \r_mem_wptr_REG[2] ( .CK(clk), .R(rst_n), .D(c_mem_wptr[2]), .Q(r_mem_wptr[2]), .QN( ));
Q_FDP1 \r_mem_wptr_REG[1] ( .CK(clk), .R(rst_n), .D(c_mem_wptr[1]), .Q(r_mem_wptr[1]), .QN( ));
Q_FDP1 \r_mem_wptr_REG[0] ( .CK(clk), .R(rst_n), .D(c_mem_wptr[0]), .Q(r_mem_wptr[0]), .QN(n308));
Q_FDP1 \r_mem_rptr_REG[10] ( .CK(clk), .R(rst_n), .D(c_mem_rptr[10]), .Q(r_mem_rptr[10]), .QN( ));
Q_FDP1 \r_mem_rptr_REG[9] ( .CK(clk), .R(rst_n), .D(c_mem_rptr[9]), .Q(r_mem_rptr[9]), .QN( ));
Q_FDP1 \r_mem_rptr_REG[8] ( .CK(clk), .R(rst_n), .D(c_mem_rptr[8]), .Q(r_mem_rptr[8]), .QN( ));
Q_FDP1 \r_mem_rptr_REG[7] ( .CK(clk), .R(rst_n), .D(c_mem_rptr[7]), .Q(r_mem_rptr[7]), .QN( ));
Q_FDP1 \r_mem_rptr_REG[6] ( .CK(clk), .R(rst_n), .D(c_mem_rptr[6]), .Q(r_mem_rptr[6]), .QN( ));
Q_FDP1 \r_mem_rptr_REG[5] ( .CK(clk), .R(rst_n), .D(c_mem_rptr[5]), .Q(r_mem_rptr[5]), .QN( ));
Q_FDP1 \r_mem_rptr_REG[4] ( .CK(clk), .R(rst_n), .D(c_mem_rptr[4]), .Q(r_mem_rptr[4]), .QN( ));
Q_FDP1 \r_mem_rptr_REG[3] ( .CK(clk), .R(rst_n), .D(c_mem_rptr[3]), .Q(r_mem_rptr[3]), .QN( ));
Q_FDP1 \r_mem_rptr_REG[2] ( .CK(clk), .R(rst_n), .D(c_mem_rptr[2]), .Q(r_mem_rptr[2]), .QN( ));
Q_FDP1 \r_mem_rptr_REG[1] ( .CK(clk), .R(rst_n), .D(c_mem_rptr[1]), .Q(r_mem_rptr[1]), .QN( ));
Q_FDP1 \r_mem_rptr_REG[0] ( .CK(clk), .R(rst_n), .D(c_mem_rptr[0]), .Q(r_mem_rptr[0]), .QN( ));
Q_FDP2 r_prefetch_empty_REG  ( .CK(clk), .S(rst_n), .D(c_prefetch_empty), .Q(r_prefetch_empty), .QN( ));
Q_FDP1 r_prefetch_full_REG  ( .CK(clk), .R(rst_n), .D(c_prefetch_full), .Q(r_prefetch_full), .QN( ));
Q_FDP1 \r_prefetch_wptr_REG[2] ( .CK(clk), .R(rst_n), .D(c_prefetch_wptr[2]), .Q(r_prefetch_wptr[2]), .QN( ));
Q_FDP1 \r_prefetch_wptr_REG[1] ( .CK(clk), .R(rst_n), .D(c_prefetch_wptr[1]), .Q(r_prefetch_wptr[1]), .QN( ));
Q_FDP2 \r_prefetch_wptr_REG[0] ( .CK(clk), .S(rst_n), .D(c_prefetch_wptr[0]), .Q(r_prefetch_wptr[0]), .QN( ));
Q_FDP1 \r_prefetch_rptr_REG[1] ( .CK(clk), .R(rst_n), .D(c_prefetch_rptr[1]), .Q(r_prefetch_rptr[1]), .QN( ));
Q_FDP1 \r_prefetch_rptr_REG[0] ( .CK(clk), .R(rst_n), .D(c_prefetch_rptr[0]), .Q(r_prefetch_rptr[0]), .QN(n835));
Q_FDP1 \r_prefetch_depth_REG[1] ( .CK(clk), .R(rst_n), .D(c_prefetch_depth[1]), .Q(r_prefetch_depth[1]), .QN(n195));
Q_FDP1 \r_prefetch_depth_REG[0] ( .CK(clk), .R(rst_n), .D(c_prefetch_depth[0]), .Q(r_prefetch_depth[0]), .QN(n196));
Q_FDP1 \r_used_slots_REG[11] ( .CK(clk), .R(rst_n), .D(c_used_slots[11]), .Q(r_used_slots[11]), .QN( ));
Q_FDP1 \r_used_slots_REG[10] ( .CK(clk), .R(rst_n), .D(c_used_slots[10]), .Q(r_used_slots[10]), .QN( ));
Q_FDP1 \r_used_slots_REG[9] ( .CK(clk), .R(rst_n), .D(c_used_slots[9]), .Q(r_used_slots[9]), .QN( ));
Q_FDP1 \r_used_slots_REG[8] ( .CK(clk), .R(rst_n), .D(c_used_slots[8]), .Q(r_used_slots[8]), .QN( ));
Q_FDP1 \r_used_slots_REG[7] ( .CK(clk), .R(rst_n), .D(c_used_slots[7]), .Q(r_used_slots[7]), .QN( ));
Q_FDP1 \r_used_slots_REG[6] ( .CK(clk), .R(rst_n), .D(c_used_slots[6]), .Q(r_used_slots[6]), .QN( ));
Q_FDP1 \r_used_slots_REG[5] ( .CK(clk), .R(rst_n), .D(c_used_slots[5]), .Q(r_used_slots[5]), .QN( ));
Q_FDP1 \r_used_slots_REG[4] ( .CK(clk), .R(rst_n), .D(c_used_slots[4]), .Q(r_used_slots[4]), .QN( ));
Q_FDP1 \r_used_slots_REG[3] ( .CK(clk), .R(rst_n), .D(c_used_slots[3]), .Q(r_used_slots[3]), .QN( ));
Q_FDP1 \r_used_slots_REG[2] ( .CK(clk), .R(rst_n), .D(c_used_slots[2]), .Q(r_used_slots[2]), .QN( ));
Q_FDP1 \r_used_slots_REG[1] ( .CK(clk), .R(rst_n), .D(c_used_slots[1]), .Q(r_used_slots[1]), .QN( ));
Q_FDP1 \r_used_slots_REG[0] ( .CK(clk), .R(rst_n), .D(c_used_slots[0]), .Q(r_used_slots[0]), .QN(n370));
Q_FDP2 \r_free_slots_REG[11] ( .CK(clk), .S(rst_n), .D(c_free_slots[11]), .Q(r_free_slots[11]), .QN( ));
Q_FDP1 \r_free_slots_REG[10] ( .CK(clk), .R(rst_n), .D(c_free_slots[10]), .Q(r_free_slots[10]), .QN( ));
Q_FDP1 \r_free_slots_REG[9] ( .CK(clk), .R(rst_n), .D(c_free_slots[9]), .Q(r_free_slots[9]), .QN( ));
Q_FDP1 \r_free_slots_REG[8] ( .CK(clk), .R(rst_n), .D(c_free_slots[8]), .Q(r_free_slots[8]), .QN( ));
Q_FDP1 \r_free_slots_REG[7] ( .CK(clk), .R(rst_n), .D(c_free_slots[7]), .Q(r_free_slots[7]), .QN( ));
Q_FDP1 \r_free_slots_REG[6] ( .CK(clk), .R(rst_n), .D(c_free_slots[6]), .Q(r_free_slots[6]), .QN( ));
Q_FDP1 \r_free_slots_REG[5] ( .CK(clk), .R(rst_n), .D(c_free_slots[5]), .Q(r_free_slots[5]), .QN( ));
Q_FDP1 \r_free_slots_REG[4] ( .CK(clk), .R(rst_n), .D(c_free_slots[4]), .Q(r_free_slots[4]), .QN( ));
Q_FDP1 \r_free_slots_REG[3] ( .CK(clk), .R(rst_n), .D(c_free_slots[3]), .Q(r_free_slots[3]), .QN( ));
Q_FDP1 \r_free_slots_REG[2] ( .CK(clk), .R(rst_n), .D(c_free_slots[2]), .Q(r_free_slots[2]), .QN( ));
Q_FDP2 \r_free_slots_REG[1] ( .CK(clk), .S(rst_n), .D(c_free_slots[1]), .Q(r_free_slots[1]), .QN( ));
Q_FDP2 \r_free_slots_REG[0] ( .CK(clk), .S(rst_n), .D(c_free_slots[0]), .Q(r_free_slots[0]), .QN(n391));
Q_NR02 U367 ( .A0(r_mem_full), .A1(n80), .Z(n117));
Q_AN02 U368 ( .A0(wen), .A1(n117), .Z(mem_wen));
Q_AN02 U369 ( .A0(ren), .A1(empty), .Z(underflow));
Q_AN02 U370 ( .A0(wen), .A1(r_mem_full), .Z(overflow));
Q_INV U371 ( .A(wen), .Z(n106));
Q_OR02 U372 ( .A0(n106), .A1(r_mem_full), .Z(n114));
Q_INV U373 ( .A(ren), .Z(n99));
Q_OR02 U374 ( .A0(n99), .A1(empty), .Z(n121));
Q_INV U375 ( .A(n121), .Z(n135));
Q_INV U376 ( .A(clear), .Z(n96));
Q_AN02 U377 ( .A0(n96), .A1(n100), .Z(n81));
Q_NR02 U378 ( .A0(r_mem_full), .A1(clear), .Z(n101));
Q_AN03 U379 ( .A0(n121), .A1(wen), .A2(n101), .Z(n102));
Q_NR02 U380 ( .A0(n102), .A1(clear), .Z(n103));
Q_AN02 U381 ( .A0(n114), .A1(n96), .Z(n104));
Q_AO21 U382 ( .A0(n135), .A1(n104), .B0(clear), .Z(n105));
Q_INV U383 ( .A(n105), .Z(n82));
Q_AN02 U384 ( .A0(n77), .A1(n106), .Z(n107));
Q_AO21 U385 ( .A0(mem_ren), .A1(n107), .B0(n110), .Z(n83));
Q_OR02 U386 ( .A0(clear), .A1(n108), .Z(n110));
Q_INV U387 ( .A(n117), .Z(n109));
Q_AN03 U388 ( .A0(mem_ren), .A1(n77), .A2(n109), .Z(n108));
Q_AN03 U389 ( .A0(wen), .A1(n96), .A2(n117), .Z(n97));
Q_NR02 U390 ( .A0(n97), .A1(n83), .Z(n111));
Q_INV U391 ( .A(n75), .Z(n112));
Q_OR02 U392 ( .A0(n80), .A1(n112), .Z(n113));
Q_OA21 U393 ( .A0(n114), .A1(n113), .B0(n115), .Z(n84));
Q_INV U394 ( .A(mem_ren), .Z(n127));
Q_NR02 U395 ( .A0(mem_ren), .A1(clear), .Z(n115));
Q_AN02 U396 ( .A0(n75), .A1(n96), .Z(n116));
Q_AN03 U397 ( .A0(n117), .A1(n116), .A2(wen), .Z(n85));
Q_AN03 U398 ( .A0(n118), .A1(n80), .A2(wen), .Z(n98));
Q_OR02 U399 ( .A0(mem_ren), .A1(n98), .Z(prefetch_wen));
Q_AN02 U400 ( .A0(n96), .A1(prefetch_wen), .Z(n86));
Q_OR02 U401 ( .A0(n86), .A1(clear), .Z(n119));
Q_INV U402 ( .A(n119), .Z(n87));
Q_NR02 U403 ( .A0(n79), .A1(clear), .Z(n120));
Q_AN02 U404 ( .A0(n135), .A1(n120), .Z(n88));
Q_AN02 U405 ( .A0(n96), .A1(n121), .Z(n89));
Q_INV U406 ( .A(n98), .Z(n129));
Q_OA21 U407 ( .A0(n99), .A1(empty), .B0(prefetch_wen), .Z(n134));
Q_NR02 U408 ( .A0(n121), .A1(mem_ren), .Z(n122));
Q_AN02 U409 ( .A0(n129), .A1(n122), .Z(n123));
Q_OA21 U410 ( .A0(n123), .A1(n134), .B0(n96), .Z(n90));
Q_AN02 U411 ( .A0(n134), .A1(n96), .Z(n124));
Q_NR02 U412 ( .A0(n124), .A1(clear), .Z(n125));
Q_AN03 U413 ( .A0(n195), .A1(n126), .A2(n135), .Z(n128));
Q_AN02 U414 ( .A0(r_prefetch_depth[0]), .A1(n127), .Z(n126));
Q_AO21 U415 ( .A0(n129), .A1(n128), .B0(clear), .Z(n91));
Q_NR02 U416 ( .A0(n86), .A1(n91), .Z(n130));
Q_AN02 U417 ( .A0(r_prefetch_depth[1]), .A1(n196), .Z(n133));
Q_AN03 U418 ( .A0(n133), .A1(n96), .A2(n134), .Z(n131));
Q_NR02 U419 ( .A0(n131), .A1(clear), .Z(n132));
Q_AN02 U420 ( .A0(n134), .A1(n133), .Z(n137));
Q_AN02 U421 ( .A0(prefetch_wen), .A1(n135), .Z(n136));
Q_OA21 U422 ( .A0(n137), .A1(n136), .B0(n96), .Z(n95));
Q_NR02 U423 ( .A0(n97), .A1(clear), .Z(n138));
Q_ND02 U424 ( .A0(ren), .A1(n74), .Z(n139));
Q_AN02 U425 ( .A0(n96), .A1(r_mem_ren_dly[1]), .Z(c_mem_ren_dly[2]));
Q_AN02 U426 ( .A0(n96), .A1(r_mem_ren_dly[0]), .Z(c_mem_ren_dly[1]));
Q_AN02 U427 ( .A0(n96), .A1(mem_ren), .Z(c_mem_ren_dly[0]));
Q_MX02 U428 ( .S(n74), .A0(n2), .A1(mem_ecc_error), .Z(rerr));
Q_MX02 U429 ( .S(n74), .A0(n3), .A1(mem_rdata[70]), .Z(rdata[70]));
Q_MX02 U430 ( .S(n74), .A0(n4), .A1(mem_rdata[69]), .Z(rdata[69]));
Q_MX02 U431 ( .S(n74), .A0(n5), .A1(mem_rdata[68]), .Z(rdata[68]));
Q_MX02 U432 ( .S(n74), .A0(n6), .A1(mem_rdata[67]), .Z(rdata[67]));
Q_MX02 U433 ( .S(n74), .A0(n7), .A1(mem_rdata[66]), .Z(rdata[66]));
Q_MX02 U434 ( .S(n74), .A0(n8), .A1(mem_rdata[65]), .Z(rdata[65]));
Q_MX02 U435 ( .S(n74), .A0(n9), .A1(mem_rdata[64]), .Z(rdata[64]));
Q_MX02 U436 ( .S(n74), .A0(n10), .A1(mem_rdata[63]), .Z(rdata[63]));
Q_MX02 U437 ( .S(n74), .A0(n11), .A1(mem_rdata[62]), .Z(rdata[62]));
Q_MX02 U438 ( .S(n74), .A0(n12), .A1(mem_rdata[61]), .Z(rdata[61]));
Q_MX02 U439 ( .S(n74), .A0(n13), .A1(mem_rdata[60]), .Z(rdata[60]));
Q_MX02 U440 ( .S(n74), .A0(n14), .A1(mem_rdata[59]), .Z(rdata[59]));
Q_MX02 U441 ( .S(n74), .A0(n15), .A1(mem_rdata[58]), .Z(rdata[58]));
Q_MX02 U442 ( .S(n74), .A0(n16), .A1(mem_rdata[57]), .Z(rdata[57]));
Q_MX02 U443 ( .S(n74), .A0(n17), .A1(mem_rdata[56]), .Z(rdata[56]));
Q_MX02 U444 ( .S(n74), .A0(n18), .A1(mem_rdata[55]), .Z(rdata[55]));
Q_MX02 U445 ( .S(n74), .A0(n19), .A1(mem_rdata[54]), .Z(rdata[54]));
Q_MX02 U446 ( .S(n74), .A0(n20), .A1(mem_rdata[53]), .Z(rdata[53]));
Q_MX02 U447 ( .S(n74), .A0(n21), .A1(mem_rdata[52]), .Z(rdata[52]));
Q_MX02 U448 ( .S(n74), .A0(n22), .A1(mem_rdata[51]), .Z(rdata[51]));
Q_MX02 U449 ( .S(n74), .A0(n23), .A1(mem_rdata[50]), .Z(rdata[50]));
Q_MX02 U450 ( .S(n74), .A0(n24), .A1(mem_rdata[49]), .Z(rdata[49]));
Q_MX02 U451 ( .S(n74), .A0(n25), .A1(mem_rdata[48]), .Z(rdata[48]));
Q_MX02 U452 ( .S(n74), .A0(n26), .A1(mem_rdata[47]), .Z(rdata[47]));
Q_MX02 U453 ( .S(n74), .A0(n27), .A1(mem_rdata[46]), .Z(rdata[46]));
Q_MX02 U454 ( .S(n74), .A0(n28), .A1(mem_rdata[45]), .Z(rdata[45]));
Q_MX02 U455 ( .S(n74), .A0(n29), .A1(mem_rdata[44]), .Z(rdata[44]));
Q_MX02 U456 ( .S(n74), .A0(n30), .A1(mem_rdata[43]), .Z(rdata[43]));
Q_MX02 U457 ( .S(n74), .A0(n31), .A1(mem_rdata[42]), .Z(rdata[42]));
Q_MX02 U458 ( .S(n74), .A0(n32), .A1(mem_rdata[41]), .Z(rdata[41]));
Q_MX02 U459 ( .S(n74), .A0(n33), .A1(mem_rdata[40]), .Z(rdata[40]));
Q_MX02 U460 ( .S(n74), .A0(n34), .A1(mem_rdata[39]), .Z(rdata[39]));
Q_MX02 U461 ( .S(n74), .A0(n35), .A1(mem_rdata[38]), .Z(rdata[38]));
Q_MX02 U462 ( .S(n74), .A0(n36), .A1(mem_rdata[37]), .Z(rdata[37]));
Q_MX02 U463 ( .S(n74), .A0(n37), .A1(mem_rdata[36]), .Z(rdata[36]));
Q_MX02 U464 ( .S(n74), .A0(n38), .A1(mem_rdata[35]), .Z(rdata[35]));
Q_MX02 U465 ( .S(n74), .A0(n39), .A1(mem_rdata[34]), .Z(rdata[34]));
Q_MX02 U466 ( .S(n74), .A0(n40), .A1(mem_rdata[33]), .Z(rdata[33]));
Q_MX02 U467 ( .S(n74), .A0(n41), .A1(mem_rdata[32]), .Z(rdata[32]));
Q_MX02 U468 ( .S(n74), .A0(n42), .A1(mem_rdata[31]), .Z(rdata[31]));
Q_MX02 U469 ( .S(n74), .A0(n43), .A1(mem_rdata[30]), .Z(rdata[30]));
Q_MX02 U470 ( .S(n74), .A0(n44), .A1(mem_rdata[29]), .Z(rdata[29]));
Q_MX02 U471 ( .S(n74), .A0(n45), .A1(mem_rdata[28]), .Z(rdata[28]));
Q_MX02 U472 ( .S(n74), .A0(n46), .A1(mem_rdata[27]), .Z(rdata[27]));
Q_MX02 U473 ( .S(n74), .A0(n47), .A1(mem_rdata[26]), .Z(rdata[26]));
Q_MX02 U474 ( .S(n74), .A0(n48), .A1(mem_rdata[25]), .Z(rdata[25]));
Q_MX02 U475 ( .S(n74), .A0(n49), .A1(mem_rdata[24]), .Z(rdata[24]));
Q_MX02 U476 ( .S(n74), .A0(n50), .A1(mem_rdata[23]), .Z(rdata[23]));
Q_MX02 U477 ( .S(n74), .A0(n51), .A1(mem_rdata[22]), .Z(rdata[22]));
Q_MX02 U478 ( .S(n74), .A0(n52), .A1(mem_rdata[21]), .Z(rdata[21]));
Q_MX02 U479 ( .S(n74), .A0(n53), .A1(mem_rdata[20]), .Z(rdata[20]));
Q_MX02 U480 ( .S(n74), .A0(n54), .A1(mem_rdata[19]), .Z(rdata[19]));
Q_MX02 U481 ( .S(n74), .A0(n55), .A1(mem_rdata[18]), .Z(rdata[18]));
Q_MX02 U482 ( .S(n74), .A0(n56), .A1(mem_rdata[17]), .Z(rdata[17]));
Q_MX02 U483 ( .S(n74), .A0(n57), .A1(mem_rdata[16]), .Z(rdata[16]));
Q_MX02 U484 ( .S(n74), .A0(n58), .A1(mem_rdata[15]), .Z(rdata[15]));
Q_MX02 U485 ( .S(n74), .A0(n59), .A1(mem_rdata[14]), .Z(rdata[14]));
Q_MX02 U486 ( .S(n74), .A0(n60), .A1(mem_rdata[13]), .Z(rdata[13]));
Q_MX02 U487 ( .S(n74), .A0(n61), .A1(mem_rdata[12]), .Z(rdata[12]));
Q_MX02 U488 ( .S(n74), .A0(n62), .A1(mem_rdata[11]), .Z(rdata[11]));
Q_MX02 U489 ( .S(n74), .A0(n63), .A1(mem_rdata[10]), .Z(rdata[10]));
Q_MX02 U490 ( .S(n74), .A0(n64), .A1(mem_rdata[9]), .Z(rdata[9]));
Q_MX02 U491 ( .S(n74), .A0(n65), .A1(mem_rdata[8]), .Z(rdata[8]));
Q_MX02 U492 ( .S(n74), .A0(n66), .A1(mem_rdata[7]), .Z(rdata[7]));
Q_MX02 U493 ( .S(n74), .A0(n67), .A1(mem_rdata[6]), .Z(rdata[6]));
Q_MX02 U494 ( .S(n74), .A0(n68), .A1(mem_rdata[5]), .Z(rdata[5]));
Q_MX02 U495 ( .S(n74), .A0(n69), .A1(mem_rdata[4]), .Z(rdata[4]));
Q_MX02 U496 ( .S(n74), .A0(n70), .A1(mem_rdata[3]), .Z(rdata[3]));
Q_MX02 U497 ( .S(n74), .A0(n71), .A1(mem_rdata[2]), .Z(rdata[2]));
Q_MX02 U498 ( .S(n74), .A0(n72), .A1(mem_rdata[1]), .Z(rdata[1]));
Q_MX02 U499 ( .S(n74), .A0(n73), .A1(mem_rdata[0]), .Z(rdata[0]));
Q_MX02 U500 ( .S(n81), .A0(n140), .A1(n141), .Z(c_used_slots[11]));
Q_AN02 U501 ( .A0(n103), .A1(r_used_slots[11]), .Z(n140));
Q_MX02 U502 ( .S(n103), .A0(n350), .A1(n329), .Z(n141));
Q_MX02 U503 ( .S(n81), .A0(n142), .A1(n143), .Z(c_used_slots[10]));
Q_AN02 U504 ( .A0(n103), .A1(r_used_slots[10]), .Z(n142));
Q_MX02 U505 ( .S(n103), .A0(n352), .A1(n331), .Z(n143));
Q_MX02 U506 ( .S(n81), .A0(n144), .A1(n145), .Z(c_used_slots[9]));
Q_AN02 U507 ( .A0(n103), .A1(r_used_slots[9]), .Z(n144));
Q_MX02 U508 ( .S(n103), .A0(n354), .A1(n333), .Z(n145));
Q_MX02 U509 ( .S(n81), .A0(n146), .A1(n147), .Z(c_used_slots[8]));
Q_AN02 U510 ( .A0(n103), .A1(r_used_slots[8]), .Z(n146));
Q_MX02 U511 ( .S(n103), .A0(n356), .A1(n335), .Z(n147));
Q_MX02 U512 ( .S(n81), .A0(n148), .A1(n149), .Z(c_used_slots[7]));
Q_AN02 U513 ( .A0(n103), .A1(r_used_slots[7]), .Z(n148));
Q_MX02 U514 ( .S(n103), .A0(n358), .A1(n337), .Z(n149));
Q_MX02 U515 ( .S(n81), .A0(n150), .A1(n151), .Z(c_used_slots[6]));
Q_AN02 U516 ( .A0(n103), .A1(r_used_slots[6]), .Z(n150));
Q_MX02 U517 ( .S(n103), .A0(n360), .A1(n339), .Z(n151));
Q_MX02 U518 ( .S(n81), .A0(n152), .A1(n153), .Z(c_used_slots[5]));
Q_AN02 U519 ( .A0(n103), .A1(r_used_slots[5]), .Z(n152));
Q_MX02 U520 ( .S(n103), .A0(n362), .A1(n341), .Z(n153));
Q_MX02 U521 ( .S(n81), .A0(n154), .A1(n155), .Z(c_used_slots[4]));
Q_AN02 U522 ( .A0(n103), .A1(r_used_slots[4]), .Z(n154));
Q_MX02 U523 ( .S(n103), .A0(n364), .A1(n343), .Z(n155));
Q_MX02 U524 ( .S(n81), .A0(n156), .A1(n157), .Z(c_used_slots[3]));
Q_AN02 U525 ( .A0(n103), .A1(r_used_slots[3]), .Z(n156));
Q_MX02 U526 ( .S(n103), .A0(n366), .A1(n345), .Z(n157));
Q_MX02 U527 ( .S(n81), .A0(n158), .A1(n159), .Z(c_used_slots[2]));
Q_AN02 U528 ( .A0(n103), .A1(r_used_slots[2]), .Z(n158));
Q_MX02 U529 ( .S(n103), .A0(n368), .A1(n347), .Z(n159));
Q_MX02 U530 ( .S(n81), .A0(n160), .A1(n161), .Z(c_used_slots[1]));
Q_AN02 U531 ( .A0(n103), .A1(r_used_slots[1]), .Z(n160));
Q_MX02 U532 ( .S(n81), .A0(n162), .A1(n370), .Z(c_used_slots[0]));
Q_AN02 U533 ( .A0(n103), .A1(r_used_slots[0]), .Z(n162));
Q_MX02 U534 ( .S(n81), .A0(n163), .A1(n164), .Z(c_free_slots[11]));
Q_OR02 U535 ( .A0(n105), .A1(r_free_slots[11]), .Z(n163));
Q_MX02 U536 ( .S(n105), .A0(n309), .A1(n371), .Z(n164));
Q_MX02 U537 ( .S(n81), .A0(n165), .A1(n166), .Z(c_free_slots[10]));
Q_AN02 U538 ( .A0(n82), .A1(r_free_slots[10]), .Z(n165));
Q_MX02 U539 ( .S(n105), .A0(n311), .A1(n373), .Z(n166));
Q_MX02 U540 ( .S(n81), .A0(n167), .A1(n168), .Z(c_free_slots[9]));
Q_AN02 U541 ( .A0(n82), .A1(r_free_slots[9]), .Z(n167));
Q_MX02 U542 ( .S(n105), .A0(n313), .A1(n375), .Z(n168));
Q_MX02 U543 ( .S(n81), .A0(n169), .A1(n170), .Z(c_free_slots[8]));
Q_AN02 U544 ( .A0(n82), .A1(r_free_slots[8]), .Z(n169));
Q_MX02 U545 ( .S(n105), .A0(n315), .A1(n377), .Z(n170));
Q_MX02 U546 ( .S(n81), .A0(n171), .A1(n172), .Z(c_free_slots[7]));
Q_AN02 U547 ( .A0(n82), .A1(r_free_slots[7]), .Z(n171));
Q_MX02 U548 ( .S(n105), .A0(n317), .A1(n379), .Z(n172));
Q_MX02 U549 ( .S(n81), .A0(n173), .A1(n174), .Z(c_free_slots[6]));
Q_AN02 U550 ( .A0(n82), .A1(r_free_slots[6]), .Z(n173));
Q_MX02 U551 ( .S(n105), .A0(n319), .A1(n381), .Z(n174));
Q_MX02 U552 ( .S(n81), .A0(n175), .A1(n176), .Z(c_free_slots[5]));
Q_AN02 U553 ( .A0(n82), .A1(r_free_slots[5]), .Z(n175));
Q_MX02 U554 ( .S(n105), .A0(n321), .A1(n383), .Z(n176));
Q_MX02 U555 ( .S(n81), .A0(n177), .A1(n178), .Z(c_free_slots[4]));
Q_AN02 U556 ( .A0(n82), .A1(r_free_slots[4]), .Z(n177));
Q_MX02 U557 ( .S(n105), .A0(n323), .A1(n385), .Z(n178));
Q_MX02 U558 ( .S(n81), .A0(n179), .A1(n180), .Z(c_free_slots[3]));
Q_AN02 U559 ( .A0(n82), .A1(r_free_slots[3]), .Z(n179));
Q_MX02 U560 ( .S(n105), .A0(n325), .A1(n387), .Z(n180));
Q_MX02 U561 ( .S(n81), .A0(n181), .A1(n182), .Z(c_free_slots[2]));
Q_AN02 U562 ( .A0(n82), .A1(r_free_slots[2]), .Z(n181));
Q_MX02 U563 ( .S(n105), .A0(n327), .A1(n389), .Z(n182));
Q_MX02 U564 ( .S(n81), .A0(n183), .A1(n184), .Z(c_free_slots[1]));
Q_OR02 U565 ( .A0(n105), .A1(r_free_slots[1]), .Z(n183));
Q_MX02 U566 ( .S(n81), .A0(n185), .A1(n391), .Z(c_free_slots[0]));
Q_OR02 U567 ( .A0(n105), .A1(r_free_slots[0]), .Z(n185));
Q_MX02 U568 ( .S(n111), .A0(n83), .A1(r_mem_empty), .Z(c_mem_empty));
Q_MX02 U569 ( .S(n84), .A0(n85), .A1(r_mem_full), .Z(c_mem_full));
Q_MX02 U570 ( .S(n86), .A0(n186), .A1(\c_mem_prefetch_wptr_dly[0][1] ), .Z(c_prefetch_wptr[2]));
Q_AN02 U571 ( .A0(n87), .A1(\c_mem_prefetch_wptr_dly[0][2] ), .Z(n186));
Q_MX02 U572 ( .S(n86), .A0(n187), .A1(\c_mem_prefetch_wptr_dly[0][0] ), .Z(c_prefetch_wptr[1]));
Q_AN02 U573 ( .A0(n87), .A1(\c_mem_prefetch_wptr_dly[0][1] ), .Z(n187));
Q_MX02 U574 ( .S(n86), .A0(n188), .A1(\c_mem_prefetch_wptr_dly[0][2] ), .Z(c_prefetch_wptr[0]));
Q_OR02 U575 ( .A0(n119), .A1(\c_mem_prefetch_wptr_dly[0][0] ), .Z(n188));
Q_MX02 U576 ( .S(n88), .A0(n189), .A1(n197), .Z(c_prefetch_rptr[1]));
Q_AN02 U577 ( .A0(n89), .A1(r_prefetch_rptr[1]), .Z(n189));
Q_MX02 U578 ( .S(n88), .A0(n190), .A1(n835), .Z(c_prefetch_rptr[0]));
Q_AN02 U579 ( .A0(n89), .A1(r_prefetch_rptr[0]), .Z(n190));
Q_MX02 U580 ( .S(n90), .A0(n191), .A1(n192), .Z(c_prefetch_depth[1]));
Q_AN02 U581 ( .A0(n125), .A1(r_prefetch_depth[1]), .Z(n191));
Q_MX02 U582 ( .S(n90), .A0(n193), .A1(n196), .Z(c_prefetch_depth[0]));
Q_AN02 U583 ( .A0(n125), .A1(r_prefetch_depth[0]), .Z(n193));
Q_MX02 U584 ( .S(n130), .A0(n91), .A1(r_prefetch_empty), .Z(c_prefetch_empty));
Q_XOR2 U585 ( .A0(r_prefetch_depth[0]), .A1(n195), .Z(n194));
Q_XOR2 U586 ( .A0(r_prefetch_rptr[1]), .A1(r_prefetch_rptr[0]), .Z(n197));
Q_AN02 U587 ( .A0(n96), .A1(n213), .Z(c_mem_rptr[10]));
Q_AN02 U588 ( .A0(n96), .A1(n214), .Z(c_mem_rptr[9]));
Q_AN02 U589 ( .A0(n96), .A1(n215), .Z(c_mem_rptr[8]));
Q_AN02 U590 ( .A0(n96), .A1(n216), .Z(c_mem_rptr[7]));
Q_AN02 U591 ( .A0(n96), .A1(n217), .Z(c_mem_rptr[6]));
Q_AN02 U592 ( .A0(n96), .A1(n218), .Z(c_mem_rptr[5]));
Q_AN02 U593 ( .A0(n96), .A1(n219), .Z(c_mem_rptr[4]));
Q_AN02 U594 ( .A0(n96), .A1(n220), .Z(c_mem_rptr[3]));
Q_AN02 U595 ( .A0(n96), .A1(n221), .Z(c_mem_rptr[2]));
Q_AN02 U596 ( .A0(n96), .A1(n222), .Z(c_mem_rptr[1]));
Q_AN02 U597 ( .A0(n96), .A1(n223), .Z(c_mem_rptr[0]));
Q_AN03 U598 ( .A0(n200), .A1(n199), .A2(n198), .Z(n75));
Q_AN03 U599 ( .A0(n203), .A1(n202), .A2(n201), .Z(n198));
Q_AN03 U600 ( .A0(n206), .A1(n205), .A2(n204), .Z(n199));
Q_AN03 U601 ( .A0(n209), .A1(n208), .A2(n207), .Z(n200));
Q_AN03 U602 ( .A0(n212), .A1(n211), .A2(n210), .Z(n201));
Q_XNR2 U603 ( .A0(n279), .A1(n213), .Z(n202));
Q_XNR2 U604 ( .A0(n280), .A1(n214), .Z(n203));
Q_XNR2 U605 ( .A0(n281), .A1(n215), .Z(n204));
Q_XNR2 U606 ( .A0(n282), .A1(n216), .Z(n205));
Q_XNR2 U607 ( .A0(n283), .A1(n217), .Z(n206));
Q_XNR2 U608 ( .A0(n284), .A1(n218), .Z(n207));
Q_XNR2 U609 ( .A0(n285), .A1(n219), .Z(n208));
Q_XNR2 U610 ( .A0(n286), .A1(n220), .Z(n209));
Q_XNR2 U611 ( .A0(n287), .A1(n221), .Z(n210));
Q_XNR2 U612 ( .A0(n288), .A1(n222), .Z(n211));
Q_XNR2 U613 ( .A0(n308), .A1(n223), .Z(n212));
Q_MX02 U614 ( .S(mem_ren), .A0(r_mem_rptr[10]), .A1(n239), .Z(n213));
Q_MX02 U615 ( .S(mem_ren), .A0(r_mem_rptr[9]), .A1(n240), .Z(n214));
Q_MX02 U616 ( .S(mem_ren), .A0(r_mem_rptr[8]), .A1(n241), .Z(n215));
Q_MX02 U617 ( .S(mem_ren), .A0(r_mem_rptr[7]), .A1(n242), .Z(n216));
Q_MX02 U618 ( .S(mem_ren), .A0(r_mem_rptr[6]), .A1(n243), .Z(n217));
Q_MX02 U619 ( .S(mem_ren), .A0(r_mem_rptr[5]), .A1(n244), .Z(n218));
Q_MX02 U620 ( .S(mem_ren), .A0(r_mem_rptr[4]), .A1(n245), .Z(n219));
Q_MX02 U621 ( .S(mem_ren), .A0(r_mem_rptr[3]), .A1(n246), .Z(n220));
Q_MX02 U622 ( .S(mem_ren), .A0(r_mem_rptr[2]), .A1(n247), .Z(n221));
Q_MX02 U623 ( .S(mem_ren), .A0(r_mem_rptr[1]), .A1(n248), .Z(n222));
Q_AN03 U624 ( .A0(n226), .A1(n225), .A2(n224), .Z(n77));
Q_AN03 U625 ( .A0(n229), .A1(n228), .A2(n227), .Z(n224));
Q_AN03 U626 ( .A0(n232), .A1(n231), .A2(n230), .Z(n225));
Q_AN03 U627 ( .A0(n235), .A1(n234), .A2(n233), .Z(n226));
Q_AN03 U628 ( .A0(n238), .A1(n237), .A2(n236), .Z(n227));
Q_XNR2 U629 ( .A0(n239), .A1(r_mem_wptr[10]), .Z(n228));
Q_XNR2 U630 ( .A0(n240), .A1(r_mem_wptr[9]), .Z(n229));
Q_XNR2 U631 ( .A0(n241), .A1(r_mem_wptr[8]), .Z(n230));
Q_XNR2 U632 ( .A0(n242), .A1(r_mem_wptr[7]), .Z(n231));
Q_XNR2 U633 ( .A0(n243), .A1(r_mem_wptr[6]), .Z(n232));
Q_XNR2 U634 ( .A0(n244), .A1(r_mem_wptr[5]), .Z(n233));
Q_XNR2 U635 ( .A0(n245), .A1(r_mem_wptr[4]), .Z(n234));
Q_XNR2 U636 ( .A0(n246), .A1(r_mem_wptr[3]), .Z(n235));
Q_XNR2 U637 ( .A0(n247), .A1(r_mem_wptr[2]), .Z(n236));
Q_XNR2 U638 ( .A0(n248), .A1(r_mem_wptr[1]), .Z(n237));
Q_XOR2 U639 ( .A0(r_mem_rptr[0]), .A1(r_mem_wptr[0]), .Z(n238));
Q_AN02 U640 ( .A0(n78), .A1(n249), .Z(n239));
Q_AN02 U641 ( .A0(n78), .A1(n251), .Z(n240));
Q_AN02 U642 ( .A0(n78), .A1(n253), .Z(n241));
Q_AN02 U643 ( .A0(n78), .A1(n255), .Z(n242));
Q_AN02 U644 ( .A0(n78), .A1(n257), .Z(n243));
Q_AN02 U645 ( .A0(n78), .A1(n259), .Z(n244));
Q_AN02 U646 ( .A0(n78), .A1(n261), .Z(n245));
Q_AN02 U647 ( .A0(n78), .A1(n263), .Z(n246));
Q_AN02 U648 ( .A0(n78), .A1(n265), .Z(n247));
Q_AN02 U649 ( .A0(n78), .A1(n267), .Z(n248));
Q_XOR2 U650 ( .A0(r_mem_rptr[10]), .A1(n250), .Z(n249));
Q_AD01HF U651 ( .A0(r_mem_rptr[9]), .B0(n252), .S(n251), .CO(n250));
Q_AD01HF U652 ( .A0(r_mem_rptr[8]), .B0(n254), .S(n253), .CO(n252));
Q_AD01HF U653 ( .A0(r_mem_rptr[7]), .B0(n256), .S(n255), .CO(n254));
Q_AD01HF U654 ( .A0(r_mem_rptr[6]), .B0(n258), .S(n257), .CO(n256));
Q_AD01HF U655 ( .A0(r_mem_rptr[5]), .B0(n260), .S(n259), .CO(n258));
Q_AD01HF U656 ( .A0(r_mem_rptr[4]), .B0(n262), .S(n261), .CO(n260));
Q_AD01HF U657 ( .A0(r_mem_rptr[3]), .B0(n264), .S(n263), .CO(n262));
Q_AD01HF U658 ( .A0(r_mem_rptr[2]), .B0(n266), .S(n265), .CO(n264));
Q_AD01HF U659 ( .A0(r_mem_rptr[1]), .B0(r_mem_rptr[0]), .S(n267), .CO(n266));
Q_MX02 U660 ( .S(n97), .A0(n268), .A1(n279), .Z(c_mem_wptr[10]));
Q_AN02 U661 ( .A0(n138), .A1(r_mem_wptr[10]), .Z(n268));
Q_MX02 U662 ( .S(n97), .A0(n269), .A1(n280), .Z(c_mem_wptr[9]));
Q_AN02 U663 ( .A0(n138), .A1(r_mem_wptr[9]), .Z(n269));
Q_MX02 U664 ( .S(n97), .A0(n270), .A1(n281), .Z(c_mem_wptr[8]));
Q_AN02 U665 ( .A0(n138), .A1(r_mem_wptr[8]), .Z(n270));
Q_MX02 U666 ( .S(n97), .A0(n271), .A1(n282), .Z(c_mem_wptr[7]));
Q_AN02 U667 ( .A0(n138), .A1(r_mem_wptr[7]), .Z(n271));
Q_MX02 U668 ( .S(n97), .A0(n272), .A1(n283), .Z(c_mem_wptr[6]));
Q_AN02 U669 ( .A0(n138), .A1(r_mem_wptr[6]), .Z(n272));
Q_MX02 U670 ( .S(n97), .A0(n273), .A1(n284), .Z(c_mem_wptr[5]));
Q_AN02 U671 ( .A0(n138), .A1(r_mem_wptr[5]), .Z(n273));
Q_MX02 U672 ( .S(n97), .A0(n274), .A1(n285), .Z(c_mem_wptr[4]));
Q_AN02 U673 ( .A0(n138), .A1(r_mem_wptr[4]), .Z(n274));
Q_MX02 U674 ( .S(n97), .A0(n275), .A1(n286), .Z(c_mem_wptr[3]));
Q_AN02 U675 ( .A0(n138), .A1(r_mem_wptr[3]), .Z(n275));
Q_MX02 U676 ( .S(n97), .A0(n276), .A1(n287), .Z(c_mem_wptr[2]));
Q_AN02 U677 ( .A0(n138), .A1(r_mem_wptr[2]), .Z(n276));
Q_MX02 U678 ( .S(n97), .A0(n277), .A1(n288), .Z(c_mem_wptr[1]));
Q_AN02 U679 ( .A0(n138), .A1(r_mem_wptr[1]), .Z(n277));
Q_MX02 U680 ( .S(n97), .A0(n278), .A1(n308), .Z(c_mem_wptr[0]));
Q_AN02 U681 ( .A0(n138), .A1(r_mem_wptr[0]), .Z(n278));
Q_AN02 U682 ( .A0(n76), .A1(n289), .Z(n279));
Q_AN02 U683 ( .A0(n76), .A1(n291), .Z(n280));
Q_AN02 U684 ( .A0(n76), .A1(n293), .Z(n281));
Q_AN02 U685 ( .A0(n76), .A1(n295), .Z(n282));
Q_AN02 U686 ( .A0(n76), .A1(n297), .Z(n283));
Q_AN02 U687 ( .A0(n76), .A1(n299), .Z(n284));
Q_AN02 U688 ( .A0(n76), .A1(n301), .Z(n285));
Q_AN02 U689 ( .A0(n76), .A1(n303), .Z(n286));
Q_AN02 U690 ( .A0(n76), .A1(n305), .Z(n287));
Q_AN02 U691 ( .A0(n76), .A1(n307), .Z(n288));
Q_XOR2 U692 ( .A0(r_mem_wptr[10]), .A1(n290), .Z(n289));
Q_AD01HF U693 ( .A0(r_mem_wptr[9]), .B0(n292), .S(n291), .CO(n290));
Q_AD01HF U694 ( .A0(r_mem_wptr[8]), .B0(n294), .S(n293), .CO(n292));
Q_AD01HF U695 ( .A0(r_mem_wptr[7]), .B0(n296), .S(n295), .CO(n294));
Q_AD01HF U696 ( .A0(r_mem_wptr[6]), .B0(n298), .S(n297), .CO(n296));
Q_AD01HF U697 ( .A0(r_mem_wptr[5]), .B0(n300), .S(n299), .CO(n298));
Q_AD01HF U698 ( .A0(r_mem_wptr[4]), .B0(n302), .S(n301), .CO(n300));
Q_AD01HF U699 ( .A0(r_mem_wptr[3]), .B0(n304), .S(n303), .CO(n302));
Q_AD01HF U700 ( .A0(r_mem_wptr[2]), .B0(n306), .S(n305), .CO(n304));
Q_AD01HF U701 ( .A0(r_mem_wptr[1]), .B0(r_mem_wptr[0]), .S(n307), .CO(n306));
Q_XNR2 U702 ( .A0(r_free_slots[11]), .A1(n310), .Z(n309));
Q_OR02 U703 ( .A0(r_free_slots[10]), .A1(n312), .Z(n310));
Q_XNR2 U704 ( .A0(r_free_slots[10]), .A1(n312), .Z(n311));
Q_OR02 U705 ( .A0(r_free_slots[9]), .A1(n314), .Z(n312));
Q_XNR2 U706 ( .A0(r_free_slots[9]), .A1(n314), .Z(n313));
Q_OR02 U707 ( .A0(r_free_slots[8]), .A1(n316), .Z(n314));
Q_XNR2 U708 ( .A0(r_free_slots[8]), .A1(n316), .Z(n315));
Q_OR02 U709 ( .A0(r_free_slots[7]), .A1(n318), .Z(n316));
Q_XNR2 U710 ( .A0(r_free_slots[7]), .A1(n318), .Z(n317));
Q_OR02 U711 ( .A0(r_free_slots[6]), .A1(n320), .Z(n318));
Q_XNR2 U712 ( .A0(r_free_slots[6]), .A1(n320), .Z(n319));
Q_OR02 U713 ( .A0(r_free_slots[5]), .A1(n322), .Z(n320));
Q_XNR2 U714 ( .A0(r_free_slots[5]), .A1(n322), .Z(n321));
Q_OR02 U715 ( .A0(r_free_slots[4]), .A1(n324), .Z(n322));
Q_XNR2 U716 ( .A0(r_free_slots[4]), .A1(n324), .Z(n323));
Q_OR02 U717 ( .A0(r_free_slots[3]), .A1(n326), .Z(n324));
Q_XNR2 U718 ( .A0(r_free_slots[3]), .A1(n326), .Z(n325));
Q_OR02 U719 ( .A0(r_free_slots[2]), .A1(n328), .Z(n326));
Q_XNR2 U720 ( .A0(r_free_slots[2]), .A1(n328), .Z(n327));
Q_OR02 U721 ( .A0(r_free_slots[1]), .A1(r_free_slots[0]), .Z(n328));
Q_XNR3 U722 ( .A0(r_free_slots[1]), .A1(r_free_slots[0]), .A2(n105), .Z(n184));
Q_XNR2 U723 ( .A0(r_used_slots[11]), .A1(n330), .Z(n329));
Q_OR02 U724 ( .A0(r_used_slots[10]), .A1(n332), .Z(n330));
Q_XNR2 U725 ( .A0(r_used_slots[10]), .A1(n332), .Z(n331));
Q_OR02 U726 ( .A0(r_used_slots[9]), .A1(n334), .Z(n332));
Q_XNR2 U727 ( .A0(r_used_slots[9]), .A1(n334), .Z(n333));
Q_OR02 U728 ( .A0(r_used_slots[8]), .A1(n336), .Z(n334));
Q_XNR2 U729 ( .A0(r_used_slots[8]), .A1(n336), .Z(n335));
Q_OR02 U730 ( .A0(r_used_slots[7]), .A1(n338), .Z(n336));
Q_XNR2 U731 ( .A0(r_used_slots[7]), .A1(n338), .Z(n337));
Q_OR02 U732 ( .A0(r_used_slots[6]), .A1(n340), .Z(n338));
Q_XNR2 U733 ( .A0(r_used_slots[6]), .A1(n340), .Z(n339));
Q_OR02 U734 ( .A0(r_used_slots[5]), .A1(n342), .Z(n340));
Q_XNR2 U735 ( .A0(r_used_slots[5]), .A1(n342), .Z(n341));
Q_OR02 U736 ( .A0(r_used_slots[4]), .A1(n344), .Z(n342));
Q_XNR2 U737 ( .A0(r_used_slots[4]), .A1(n344), .Z(n343));
Q_OR02 U738 ( .A0(r_used_slots[3]), .A1(n346), .Z(n344));
Q_XNR2 U739 ( .A0(r_used_slots[3]), .A1(n346), .Z(n345));
Q_OR02 U740 ( .A0(r_used_slots[2]), .A1(n348), .Z(n346));
Q_XNR2 U741 ( .A0(r_used_slots[2]), .A1(n348), .Z(n347));
Q_OR02 U742 ( .A0(r_used_slots[1]), .A1(r_used_slots[0]), .Z(n348));
Q_XNR2 U743 ( .A0(r_used_slots[1]), .A1(r_used_slots[0]), .Z(n349));
Q_XOR2 U744 ( .A0(r_used_slots[11]), .A1(n351), .Z(n350));
Q_AD01HF U745 ( .A0(r_used_slots[10]), .B0(n353), .S(n352), .CO(n351));
Q_AD01HF U746 ( .A0(r_used_slots[9]), .B0(n355), .S(n354), .CO(n353));
Q_AD01HF U747 ( .A0(r_used_slots[8]), .B0(n357), .S(n356), .CO(n355));
Q_AD01HF U748 ( .A0(r_used_slots[7]), .B0(n359), .S(n358), .CO(n357));
Q_AD01HF U749 ( .A0(r_used_slots[6]), .B0(n361), .S(n360), .CO(n359));
Q_AD01HF U750 ( .A0(r_used_slots[5]), .B0(n363), .S(n362), .CO(n361));
Q_AD01HF U751 ( .A0(r_used_slots[4]), .B0(n365), .S(n364), .CO(n363));
Q_AD01HF U752 ( .A0(r_used_slots[3]), .B0(n367), .S(n366), .CO(n365));
Q_AD01HF U753 ( .A0(r_used_slots[2]), .B0(n369), .S(n368), .CO(n367));
Q_XOR2 U754 ( .A0(r_free_slots[11]), .A1(n372), .Z(n371));
Q_AD01HF U755 ( .A0(r_free_slots[10]), .B0(n374), .S(n373), .CO(n372));
Q_AD01HF U756 ( .A0(r_free_slots[9]), .B0(n376), .S(n375), .CO(n374));
Q_AD01HF U757 ( .A0(r_free_slots[8]), .B0(n378), .S(n377), .CO(n376));
Q_AD01HF U758 ( .A0(r_free_slots[7]), .B0(n380), .S(n379), .CO(n378));
Q_AD01HF U759 ( .A0(r_free_slots[6]), .B0(n382), .S(n381), .CO(n380));
Q_AD01HF U760 ( .A0(r_free_slots[5]), .B0(n384), .S(n383), .CO(n382));
Q_AD01HF U761 ( .A0(r_free_slots[4]), .B0(n386), .S(n385), .CO(n384));
Q_AD01HF U762 ( .A0(r_free_slots[3]), .B0(n388), .S(n387), .CO(n386));
Q_AD01HF U763 ( .A0(r_free_slots[2]), .B0(n390), .S(n389), .CO(n388));
Q_MX02 U764 ( .S(n92), .A0(\r_prefetch_data[0][71] ), .A1(n750), .Z(\c_prefetch_data[0][71] ));
Q_MX02 U765 ( .S(n92), .A0(\r_prefetch_data[0][70] ), .A1(n679), .Z(\c_prefetch_data[0][70] ));
Q_MX02 U766 ( .S(n92), .A0(\r_prefetch_data[0][69] ), .A1(n680), .Z(\c_prefetch_data[0][69] ));
Q_MX02 U767 ( .S(n92), .A0(\r_prefetch_data[0][68] ), .A1(n681), .Z(\c_prefetch_data[0][68] ));
Q_MX02 U768 ( .S(n92), .A0(\r_prefetch_data[0][67] ), .A1(n682), .Z(\c_prefetch_data[0][67] ));
Q_MX02 U769 ( .S(n92), .A0(\r_prefetch_data[0][66] ), .A1(n683), .Z(\c_prefetch_data[0][66] ));
Q_MX02 U770 ( .S(n92), .A0(\r_prefetch_data[0][65] ), .A1(n684), .Z(\c_prefetch_data[0][65] ));
Q_MX02 U771 ( .S(n92), .A0(\r_prefetch_data[0][64] ), .A1(n685), .Z(\c_prefetch_data[0][64] ));
Q_MX02 U772 ( .S(n92), .A0(\r_prefetch_data[0][63] ), .A1(n686), .Z(\c_prefetch_data[0][63] ));
Q_MX02 U773 ( .S(n92), .A0(\r_prefetch_data[0][62] ), .A1(n687), .Z(\c_prefetch_data[0][62] ));
Q_MX02 U774 ( .S(n92), .A0(\r_prefetch_data[0][61] ), .A1(n688), .Z(\c_prefetch_data[0][61] ));
Q_MX02 U775 ( .S(n92), .A0(\r_prefetch_data[0][60] ), .A1(n689), .Z(\c_prefetch_data[0][60] ));
Q_MX02 U776 ( .S(n92), .A0(\r_prefetch_data[0][59] ), .A1(n690), .Z(\c_prefetch_data[0][59] ));
Q_MX02 U777 ( .S(n92), .A0(\r_prefetch_data[0][58] ), .A1(n691), .Z(\c_prefetch_data[0][58] ));
Q_MX02 U778 ( .S(n92), .A0(\r_prefetch_data[0][57] ), .A1(n692), .Z(\c_prefetch_data[0][57] ));
Q_MX02 U779 ( .S(n92), .A0(\r_prefetch_data[0][56] ), .A1(n693), .Z(\c_prefetch_data[0][56] ));
Q_MX02 U780 ( .S(n92), .A0(\r_prefetch_data[0][55] ), .A1(n694), .Z(\c_prefetch_data[0][55] ));
Q_MX02 U781 ( .S(n92), .A0(\r_prefetch_data[0][54] ), .A1(n695), .Z(\c_prefetch_data[0][54] ));
Q_MX02 U782 ( .S(n92), .A0(\r_prefetch_data[0][53] ), .A1(n696), .Z(\c_prefetch_data[0][53] ));
Q_MX02 U783 ( .S(n92), .A0(\r_prefetch_data[0][52] ), .A1(n697), .Z(\c_prefetch_data[0][52] ));
Q_MX02 U784 ( .S(n92), .A0(\r_prefetch_data[0][51] ), .A1(n698), .Z(\c_prefetch_data[0][51] ));
Q_MX02 U785 ( .S(n92), .A0(\r_prefetch_data[0][50] ), .A1(n699), .Z(\c_prefetch_data[0][50] ));
Q_MX02 U786 ( .S(n92), .A0(\r_prefetch_data[0][49] ), .A1(n700), .Z(\c_prefetch_data[0][49] ));
Q_MX02 U787 ( .S(n92), .A0(\r_prefetch_data[0][48] ), .A1(n701), .Z(\c_prefetch_data[0][48] ));
Q_MX02 U788 ( .S(n92), .A0(\r_prefetch_data[0][47] ), .A1(n702), .Z(\c_prefetch_data[0][47] ));
Q_MX02 U789 ( .S(n92), .A0(\r_prefetch_data[0][46] ), .A1(n703), .Z(\c_prefetch_data[0][46] ));
Q_MX02 U790 ( .S(n92), .A0(\r_prefetch_data[0][45] ), .A1(n704), .Z(\c_prefetch_data[0][45] ));
Q_MX02 U791 ( .S(n92), .A0(\r_prefetch_data[0][44] ), .A1(n705), .Z(\c_prefetch_data[0][44] ));
Q_MX02 U792 ( .S(n92), .A0(\r_prefetch_data[0][43] ), .A1(n706), .Z(\c_prefetch_data[0][43] ));
Q_MX02 U793 ( .S(n92), .A0(\r_prefetch_data[0][42] ), .A1(n707), .Z(\c_prefetch_data[0][42] ));
Q_MX02 U794 ( .S(n92), .A0(\r_prefetch_data[0][41] ), .A1(n708), .Z(\c_prefetch_data[0][41] ));
Q_MX02 U795 ( .S(n92), .A0(\r_prefetch_data[0][40] ), .A1(n709), .Z(\c_prefetch_data[0][40] ));
Q_MX02 U796 ( .S(n92), .A0(\r_prefetch_data[0][39] ), .A1(n710), .Z(\c_prefetch_data[0][39] ));
Q_MX02 U797 ( .S(n92), .A0(\r_prefetch_data[0][38] ), .A1(n711), .Z(\c_prefetch_data[0][38] ));
Q_MX02 U798 ( .S(n92), .A0(\r_prefetch_data[0][37] ), .A1(n712), .Z(\c_prefetch_data[0][37] ));
Q_MX02 U799 ( .S(n92), .A0(\r_prefetch_data[0][36] ), .A1(n713), .Z(\c_prefetch_data[0][36] ));
Q_MX02 U800 ( .S(n92), .A0(\r_prefetch_data[0][35] ), .A1(n714), .Z(\c_prefetch_data[0][35] ));
Q_MX02 U801 ( .S(n92), .A0(\r_prefetch_data[0][34] ), .A1(n715), .Z(\c_prefetch_data[0][34] ));
Q_MX02 U802 ( .S(n92), .A0(\r_prefetch_data[0][33] ), .A1(n716), .Z(\c_prefetch_data[0][33] ));
Q_MX02 U803 ( .S(n92), .A0(\r_prefetch_data[0][32] ), .A1(n717), .Z(\c_prefetch_data[0][32] ));
Q_MX02 U804 ( .S(n92), .A0(\r_prefetch_data[0][31] ), .A1(n718), .Z(\c_prefetch_data[0][31] ));
Q_MX02 U805 ( .S(n92), .A0(\r_prefetch_data[0][30] ), .A1(n719), .Z(\c_prefetch_data[0][30] ));
Q_MX02 U806 ( .S(n92), .A0(\r_prefetch_data[0][29] ), .A1(n720), .Z(\c_prefetch_data[0][29] ));
Q_MX02 U807 ( .S(n92), .A0(\r_prefetch_data[0][28] ), .A1(n721), .Z(\c_prefetch_data[0][28] ));
Q_MX02 U808 ( .S(n92), .A0(\r_prefetch_data[0][27] ), .A1(n722), .Z(\c_prefetch_data[0][27] ));
Q_MX02 U809 ( .S(n92), .A0(\r_prefetch_data[0][26] ), .A1(n723), .Z(\c_prefetch_data[0][26] ));
Q_MX02 U810 ( .S(n92), .A0(\r_prefetch_data[0][25] ), .A1(n724), .Z(\c_prefetch_data[0][25] ));
Q_MX02 U811 ( .S(n92), .A0(\r_prefetch_data[0][24] ), .A1(n725), .Z(\c_prefetch_data[0][24] ));
Q_MX02 U812 ( .S(n92), .A0(\r_prefetch_data[0][23] ), .A1(n726), .Z(\c_prefetch_data[0][23] ));
Q_MX02 U813 ( .S(n92), .A0(\r_prefetch_data[0][22] ), .A1(n727), .Z(\c_prefetch_data[0][22] ));
Q_MX02 U814 ( .S(n92), .A0(\r_prefetch_data[0][21] ), .A1(n728), .Z(\c_prefetch_data[0][21] ));
Q_MX02 U815 ( .S(n92), .A0(\r_prefetch_data[0][20] ), .A1(n729), .Z(\c_prefetch_data[0][20] ));
Q_MX02 U816 ( .S(n92), .A0(\r_prefetch_data[0][19] ), .A1(n730), .Z(\c_prefetch_data[0][19] ));
Q_MX02 U817 ( .S(n92), .A0(\r_prefetch_data[0][18] ), .A1(n731), .Z(\c_prefetch_data[0][18] ));
Q_MX02 U818 ( .S(n92), .A0(\r_prefetch_data[0][17] ), .A1(n732), .Z(\c_prefetch_data[0][17] ));
Q_MX02 U819 ( .S(n92), .A0(\r_prefetch_data[0][16] ), .A1(n733), .Z(\c_prefetch_data[0][16] ));
Q_MX02 U820 ( .S(n92), .A0(\r_prefetch_data[0][15] ), .A1(n734), .Z(\c_prefetch_data[0][15] ));
Q_MX02 U821 ( .S(n92), .A0(\r_prefetch_data[0][14] ), .A1(n735), .Z(\c_prefetch_data[0][14] ));
Q_MX02 U822 ( .S(n92), .A0(\r_prefetch_data[0][13] ), .A1(n736), .Z(\c_prefetch_data[0][13] ));
Q_MX02 U823 ( .S(n92), .A0(\r_prefetch_data[0][12] ), .A1(n737), .Z(\c_prefetch_data[0][12] ));
Q_MX02 U824 ( .S(n92), .A0(\r_prefetch_data[0][11] ), .A1(n738), .Z(\c_prefetch_data[0][11] ));
Q_MX02 U825 ( .S(n92), .A0(\r_prefetch_data[0][10] ), .A1(n739), .Z(\c_prefetch_data[0][10] ));
Q_MX02 U826 ( .S(n92), .A0(\r_prefetch_data[0][9] ), .A1(n740), .Z(\c_prefetch_data[0][9] ));
Q_MX02 U827 ( .S(n92), .A0(\r_prefetch_data[0][8] ), .A1(n741), .Z(\c_prefetch_data[0][8] ));
Q_MX02 U828 ( .S(n92), .A0(\r_prefetch_data[0][7] ), .A1(n742), .Z(\c_prefetch_data[0][7] ));
Q_MX02 U829 ( .S(n92), .A0(\r_prefetch_data[0][6] ), .A1(n743), .Z(\c_prefetch_data[0][6] ));
Q_MX02 U830 ( .S(n92), .A0(\r_prefetch_data[0][5] ), .A1(n744), .Z(\c_prefetch_data[0][5] ));
Q_MX02 U831 ( .S(n92), .A0(\r_prefetch_data[0][4] ), .A1(n745), .Z(\c_prefetch_data[0][4] ));
Q_MX02 U832 ( .S(n92), .A0(\r_prefetch_data[0][3] ), .A1(n746), .Z(\c_prefetch_data[0][3] ));
Q_MX02 U833 ( .S(n92), .A0(\r_prefetch_data[0][2] ), .A1(n747), .Z(\c_prefetch_data[0][2] ));
Q_MX02 U834 ( .S(n92), .A0(\r_prefetch_data[0][1] ), .A1(n748), .Z(\c_prefetch_data[0][1] ));
Q_MX02 U835 ( .S(n92), .A0(\r_prefetch_data[0][0] ), .A1(n749), .Z(\c_prefetch_data[0][0] ));
Q_MX02 U836 ( .S(n93), .A0(\r_prefetch_data[1][71] ), .A1(n607), .Z(\c_prefetch_data[1][71] ));
Q_MX02 U837 ( .S(n93), .A0(\r_prefetch_data[1][70] ), .A1(n536), .Z(\c_prefetch_data[1][70] ));
Q_MX02 U838 ( .S(n93), .A0(\r_prefetch_data[1][69] ), .A1(n537), .Z(\c_prefetch_data[1][69] ));
Q_MX02 U839 ( .S(n93), .A0(\r_prefetch_data[1][68] ), .A1(n538), .Z(\c_prefetch_data[1][68] ));
Q_MX02 U840 ( .S(n93), .A0(\r_prefetch_data[1][67] ), .A1(n539), .Z(\c_prefetch_data[1][67] ));
Q_MX02 U841 ( .S(n93), .A0(\r_prefetch_data[1][66] ), .A1(n540), .Z(\c_prefetch_data[1][66] ));
Q_MX02 U842 ( .S(n93), .A0(\r_prefetch_data[1][65] ), .A1(n541), .Z(\c_prefetch_data[1][65] ));
Q_MX02 U843 ( .S(n93), .A0(\r_prefetch_data[1][64] ), .A1(n542), .Z(\c_prefetch_data[1][64] ));
Q_MX02 U844 ( .S(n93), .A0(\r_prefetch_data[1][63] ), .A1(n543), .Z(\c_prefetch_data[1][63] ));
Q_MX02 U845 ( .S(n93), .A0(\r_prefetch_data[1][62] ), .A1(n544), .Z(\c_prefetch_data[1][62] ));
Q_MX02 U846 ( .S(n93), .A0(\r_prefetch_data[1][61] ), .A1(n545), .Z(\c_prefetch_data[1][61] ));
Q_MX02 U847 ( .S(n93), .A0(\r_prefetch_data[1][60] ), .A1(n546), .Z(\c_prefetch_data[1][60] ));
Q_MX02 U848 ( .S(n93), .A0(\r_prefetch_data[1][59] ), .A1(n547), .Z(\c_prefetch_data[1][59] ));
Q_MX02 U849 ( .S(n93), .A0(\r_prefetch_data[1][58] ), .A1(n548), .Z(\c_prefetch_data[1][58] ));
Q_MX02 U850 ( .S(n93), .A0(\r_prefetch_data[1][57] ), .A1(n549), .Z(\c_prefetch_data[1][57] ));
Q_MX02 U851 ( .S(n93), .A0(\r_prefetch_data[1][56] ), .A1(n550), .Z(\c_prefetch_data[1][56] ));
Q_MX02 U852 ( .S(n93), .A0(\r_prefetch_data[1][55] ), .A1(n551), .Z(\c_prefetch_data[1][55] ));
Q_MX02 U853 ( .S(n93), .A0(\r_prefetch_data[1][54] ), .A1(n552), .Z(\c_prefetch_data[1][54] ));
Q_MX02 U854 ( .S(n93), .A0(\r_prefetch_data[1][53] ), .A1(n553), .Z(\c_prefetch_data[1][53] ));
Q_MX02 U855 ( .S(n93), .A0(\r_prefetch_data[1][52] ), .A1(n554), .Z(\c_prefetch_data[1][52] ));
Q_MX02 U856 ( .S(n93), .A0(\r_prefetch_data[1][51] ), .A1(n555), .Z(\c_prefetch_data[1][51] ));
Q_MX02 U857 ( .S(n93), .A0(\r_prefetch_data[1][50] ), .A1(n556), .Z(\c_prefetch_data[1][50] ));
Q_MX02 U858 ( .S(n93), .A0(\r_prefetch_data[1][49] ), .A1(n557), .Z(\c_prefetch_data[1][49] ));
Q_MX02 U859 ( .S(n93), .A0(\r_prefetch_data[1][48] ), .A1(n558), .Z(\c_prefetch_data[1][48] ));
Q_MX02 U860 ( .S(n93), .A0(\r_prefetch_data[1][47] ), .A1(n559), .Z(\c_prefetch_data[1][47] ));
Q_MX02 U861 ( .S(n93), .A0(\r_prefetch_data[1][46] ), .A1(n560), .Z(\c_prefetch_data[1][46] ));
Q_MX02 U862 ( .S(n93), .A0(\r_prefetch_data[1][45] ), .A1(n561), .Z(\c_prefetch_data[1][45] ));
Q_MX02 U863 ( .S(n93), .A0(\r_prefetch_data[1][44] ), .A1(n562), .Z(\c_prefetch_data[1][44] ));
Q_MX02 U864 ( .S(n93), .A0(\r_prefetch_data[1][43] ), .A1(n563), .Z(\c_prefetch_data[1][43] ));
Q_MX02 U865 ( .S(n93), .A0(\r_prefetch_data[1][42] ), .A1(n564), .Z(\c_prefetch_data[1][42] ));
Q_MX02 U866 ( .S(n93), .A0(\r_prefetch_data[1][41] ), .A1(n565), .Z(\c_prefetch_data[1][41] ));
Q_MX02 U867 ( .S(n93), .A0(\r_prefetch_data[1][40] ), .A1(n566), .Z(\c_prefetch_data[1][40] ));
Q_MX02 U868 ( .S(n93), .A0(\r_prefetch_data[1][39] ), .A1(n567), .Z(\c_prefetch_data[1][39] ));
Q_MX02 U869 ( .S(n93), .A0(\r_prefetch_data[1][38] ), .A1(n568), .Z(\c_prefetch_data[1][38] ));
Q_MX02 U870 ( .S(n93), .A0(\r_prefetch_data[1][37] ), .A1(n569), .Z(\c_prefetch_data[1][37] ));
Q_MX02 U871 ( .S(n93), .A0(\r_prefetch_data[1][36] ), .A1(n570), .Z(\c_prefetch_data[1][36] ));
Q_MX02 U872 ( .S(n93), .A0(\r_prefetch_data[1][35] ), .A1(n571), .Z(\c_prefetch_data[1][35] ));
Q_MX02 U873 ( .S(n93), .A0(\r_prefetch_data[1][34] ), .A1(n572), .Z(\c_prefetch_data[1][34] ));
Q_MX02 U874 ( .S(n93), .A0(\r_prefetch_data[1][33] ), .A1(n573), .Z(\c_prefetch_data[1][33] ));
Q_MX02 U875 ( .S(n93), .A0(\r_prefetch_data[1][32] ), .A1(n574), .Z(\c_prefetch_data[1][32] ));
Q_MX02 U876 ( .S(n93), .A0(\r_prefetch_data[1][31] ), .A1(n575), .Z(\c_prefetch_data[1][31] ));
Q_MX02 U877 ( .S(n93), .A0(\r_prefetch_data[1][30] ), .A1(n576), .Z(\c_prefetch_data[1][30] ));
Q_MX02 U878 ( .S(n93), .A0(\r_prefetch_data[1][29] ), .A1(n577), .Z(\c_prefetch_data[1][29] ));
Q_MX02 U879 ( .S(n93), .A0(\r_prefetch_data[1][28] ), .A1(n578), .Z(\c_prefetch_data[1][28] ));
Q_MX02 U880 ( .S(n93), .A0(\r_prefetch_data[1][27] ), .A1(n579), .Z(\c_prefetch_data[1][27] ));
Q_MX02 U881 ( .S(n93), .A0(\r_prefetch_data[1][26] ), .A1(n580), .Z(\c_prefetch_data[1][26] ));
Q_MX02 U882 ( .S(n93), .A0(\r_prefetch_data[1][25] ), .A1(n581), .Z(\c_prefetch_data[1][25] ));
Q_MX02 U883 ( .S(n93), .A0(\r_prefetch_data[1][24] ), .A1(n582), .Z(\c_prefetch_data[1][24] ));
Q_MX02 U884 ( .S(n93), .A0(\r_prefetch_data[1][23] ), .A1(n583), .Z(\c_prefetch_data[1][23] ));
Q_MX02 U885 ( .S(n93), .A0(\r_prefetch_data[1][22] ), .A1(n584), .Z(\c_prefetch_data[1][22] ));
Q_MX02 U886 ( .S(n93), .A0(\r_prefetch_data[1][21] ), .A1(n585), .Z(\c_prefetch_data[1][21] ));
Q_MX02 U887 ( .S(n93), .A0(\r_prefetch_data[1][20] ), .A1(n586), .Z(\c_prefetch_data[1][20] ));
Q_MX02 U888 ( .S(n93), .A0(\r_prefetch_data[1][19] ), .A1(n587), .Z(\c_prefetch_data[1][19] ));
Q_MX02 U889 ( .S(n93), .A0(\r_prefetch_data[1][18] ), .A1(n588), .Z(\c_prefetch_data[1][18] ));
Q_MX02 U890 ( .S(n93), .A0(\r_prefetch_data[1][17] ), .A1(n589), .Z(\c_prefetch_data[1][17] ));
Q_MX02 U891 ( .S(n93), .A0(\r_prefetch_data[1][16] ), .A1(n590), .Z(\c_prefetch_data[1][16] ));
Q_MX02 U892 ( .S(n93), .A0(\r_prefetch_data[1][15] ), .A1(n591), .Z(\c_prefetch_data[1][15] ));
Q_MX02 U893 ( .S(n93), .A0(\r_prefetch_data[1][14] ), .A1(n592), .Z(\c_prefetch_data[1][14] ));
Q_MX02 U894 ( .S(n93), .A0(\r_prefetch_data[1][13] ), .A1(n593), .Z(\c_prefetch_data[1][13] ));
Q_MX02 U895 ( .S(n93), .A0(\r_prefetch_data[1][12] ), .A1(n594), .Z(\c_prefetch_data[1][12] ));
Q_MX02 U896 ( .S(n93), .A0(\r_prefetch_data[1][11] ), .A1(n595), .Z(\c_prefetch_data[1][11] ));
Q_MX02 U897 ( .S(n93), .A0(\r_prefetch_data[1][10] ), .A1(n596), .Z(\c_prefetch_data[1][10] ));
Q_MX02 U898 ( .S(n93), .A0(\r_prefetch_data[1][9] ), .A1(n597), .Z(\c_prefetch_data[1][9] ));
Q_MX02 U899 ( .S(n93), .A0(\r_prefetch_data[1][8] ), .A1(n598), .Z(\c_prefetch_data[1][8] ));
Q_MX02 U900 ( .S(n93), .A0(\r_prefetch_data[1][7] ), .A1(n599), .Z(\c_prefetch_data[1][7] ));
Q_MX02 U901 ( .S(n93), .A0(\r_prefetch_data[1][6] ), .A1(n600), .Z(\c_prefetch_data[1][6] ));
Q_MX02 U902 ( .S(n93), .A0(\r_prefetch_data[1][5] ), .A1(n601), .Z(\c_prefetch_data[1][5] ));
Q_MX02 U903 ( .S(n93), .A0(\r_prefetch_data[1][4] ), .A1(n602), .Z(\c_prefetch_data[1][4] ));
Q_MX02 U904 ( .S(n93), .A0(\r_prefetch_data[1][3] ), .A1(n603), .Z(\c_prefetch_data[1][3] ));
Q_MX02 U905 ( .S(n93), .A0(\r_prefetch_data[1][2] ), .A1(n604), .Z(\c_prefetch_data[1][2] ));
Q_MX02 U906 ( .S(n93), .A0(\r_prefetch_data[1][1] ), .A1(n605), .Z(\c_prefetch_data[1][1] ));
Q_MX02 U907 ( .S(n93), .A0(\r_prefetch_data[1][0] ), .A1(n606), .Z(\c_prefetch_data[1][0] ));
Q_MX02 U908 ( .S(n94), .A0(\r_prefetch_data[2][71] ), .A1(n464), .Z(\c_prefetch_data[2][71] ));
Q_MX02 U909 ( .S(n94), .A0(\r_prefetch_data[2][70] ), .A1(n393), .Z(\c_prefetch_data[2][70] ));
Q_MX02 U910 ( .S(n94), .A0(\r_prefetch_data[2][69] ), .A1(n394), .Z(\c_prefetch_data[2][69] ));
Q_MX02 U911 ( .S(n94), .A0(\r_prefetch_data[2][68] ), .A1(n395), .Z(\c_prefetch_data[2][68] ));
Q_MX02 U912 ( .S(n94), .A0(\r_prefetch_data[2][67] ), .A1(n396), .Z(\c_prefetch_data[2][67] ));
Q_MX02 U913 ( .S(n94), .A0(\r_prefetch_data[2][66] ), .A1(n397), .Z(\c_prefetch_data[2][66] ));
Q_MX02 U914 ( .S(n94), .A0(\r_prefetch_data[2][65] ), .A1(n398), .Z(\c_prefetch_data[2][65] ));
Q_MX02 U915 ( .S(n94), .A0(\r_prefetch_data[2][64] ), .A1(n399), .Z(\c_prefetch_data[2][64] ));
Q_MX02 U916 ( .S(n94), .A0(\r_prefetch_data[2][63] ), .A1(n400), .Z(\c_prefetch_data[2][63] ));
Q_MX02 U917 ( .S(n94), .A0(\r_prefetch_data[2][62] ), .A1(n401), .Z(\c_prefetch_data[2][62] ));
Q_MX02 U918 ( .S(n94), .A0(\r_prefetch_data[2][61] ), .A1(n402), .Z(\c_prefetch_data[2][61] ));
Q_MX02 U919 ( .S(n94), .A0(\r_prefetch_data[2][60] ), .A1(n403), .Z(\c_prefetch_data[2][60] ));
Q_MX02 U920 ( .S(n94), .A0(\r_prefetch_data[2][59] ), .A1(n404), .Z(\c_prefetch_data[2][59] ));
Q_MX02 U921 ( .S(n94), .A0(\r_prefetch_data[2][58] ), .A1(n405), .Z(\c_prefetch_data[2][58] ));
Q_MX02 U922 ( .S(n94), .A0(\r_prefetch_data[2][57] ), .A1(n406), .Z(\c_prefetch_data[2][57] ));
Q_MX02 U923 ( .S(n94), .A0(\r_prefetch_data[2][56] ), .A1(n407), .Z(\c_prefetch_data[2][56] ));
Q_MX02 U924 ( .S(n94), .A0(\r_prefetch_data[2][55] ), .A1(n408), .Z(\c_prefetch_data[2][55] ));
Q_MX02 U925 ( .S(n94), .A0(\r_prefetch_data[2][54] ), .A1(n409), .Z(\c_prefetch_data[2][54] ));
Q_MX02 U926 ( .S(n94), .A0(\r_prefetch_data[2][53] ), .A1(n410), .Z(\c_prefetch_data[2][53] ));
Q_MX02 U927 ( .S(n94), .A0(\r_prefetch_data[2][52] ), .A1(n411), .Z(\c_prefetch_data[2][52] ));
Q_MX02 U928 ( .S(n94), .A0(\r_prefetch_data[2][51] ), .A1(n412), .Z(\c_prefetch_data[2][51] ));
Q_MX02 U929 ( .S(n94), .A0(\r_prefetch_data[2][50] ), .A1(n413), .Z(\c_prefetch_data[2][50] ));
Q_MX02 U930 ( .S(n94), .A0(\r_prefetch_data[2][49] ), .A1(n414), .Z(\c_prefetch_data[2][49] ));
Q_MX02 U931 ( .S(n94), .A0(\r_prefetch_data[2][48] ), .A1(n415), .Z(\c_prefetch_data[2][48] ));
Q_MX02 U932 ( .S(n94), .A0(\r_prefetch_data[2][47] ), .A1(n416), .Z(\c_prefetch_data[2][47] ));
Q_MX02 U933 ( .S(n94), .A0(\r_prefetch_data[2][46] ), .A1(n417), .Z(\c_prefetch_data[2][46] ));
Q_MX02 U934 ( .S(n94), .A0(\r_prefetch_data[2][45] ), .A1(n418), .Z(\c_prefetch_data[2][45] ));
Q_MX02 U935 ( .S(n94), .A0(\r_prefetch_data[2][44] ), .A1(n419), .Z(\c_prefetch_data[2][44] ));
Q_MX02 U936 ( .S(n94), .A0(\r_prefetch_data[2][43] ), .A1(n420), .Z(\c_prefetch_data[2][43] ));
Q_MX02 U937 ( .S(n94), .A0(\r_prefetch_data[2][42] ), .A1(n421), .Z(\c_prefetch_data[2][42] ));
Q_MX02 U938 ( .S(n94), .A0(\r_prefetch_data[2][41] ), .A1(n422), .Z(\c_prefetch_data[2][41] ));
Q_MX02 U939 ( .S(n94), .A0(\r_prefetch_data[2][40] ), .A1(n423), .Z(\c_prefetch_data[2][40] ));
Q_MX02 U940 ( .S(n94), .A0(\r_prefetch_data[2][39] ), .A1(n424), .Z(\c_prefetch_data[2][39] ));
Q_MX02 U941 ( .S(n94), .A0(\r_prefetch_data[2][38] ), .A1(n425), .Z(\c_prefetch_data[2][38] ));
Q_MX02 U942 ( .S(n94), .A0(\r_prefetch_data[2][37] ), .A1(n426), .Z(\c_prefetch_data[2][37] ));
Q_MX02 U943 ( .S(n94), .A0(\r_prefetch_data[2][36] ), .A1(n427), .Z(\c_prefetch_data[2][36] ));
Q_MX02 U944 ( .S(n94), .A0(\r_prefetch_data[2][35] ), .A1(n428), .Z(\c_prefetch_data[2][35] ));
Q_MX02 U945 ( .S(n94), .A0(\r_prefetch_data[2][34] ), .A1(n429), .Z(\c_prefetch_data[2][34] ));
Q_MX02 U946 ( .S(n94), .A0(\r_prefetch_data[2][33] ), .A1(n430), .Z(\c_prefetch_data[2][33] ));
Q_MX02 U947 ( .S(n94), .A0(\r_prefetch_data[2][32] ), .A1(n431), .Z(\c_prefetch_data[2][32] ));
Q_MX02 U948 ( .S(n94), .A0(\r_prefetch_data[2][31] ), .A1(n432), .Z(\c_prefetch_data[2][31] ));
Q_MX02 U949 ( .S(n94), .A0(\r_prefetch_data[2][30] ), .A1(n433), .Z(\c_prefetch_data[2][30] ));
Q_MX02 U950 ( .S(n94), .A0(\r_prefetch_data[2][29] ), .A1(n434), .Z(\c_prefetch_data[2][29] ));
Q_MX02 U951 ( .S(n94), .A0(\r_prefetch_data[2][28] ), .A1(n435), .Z(\c_prefetch_data[2][28] ));
Q_MX02 U952 ( .S(n94), .A0(\r_prefetch_data[2][27] ), .A1(n436), .Z(\c_prefetch_data[2][27] ));
Q_MX02 U953 ( .S(n94), .A0(\r_prefetch_data[2][26] ), .A1(n437), .Z(\c_prefetch_data[2][26] ));
Q_MX02 U954 ( .S(n94), .A0(\r_prefetch_data[2][25] ), .A1(n438), .Z(\c_prefetch_data[2][25] ));
Q_MX02 U955 ( .S(n94), .A0(\r_prefetch_data[2][24] ), .A1(n439), .Z(\c_prefetch_data[2][24] ));
Q_MX02 U956 ( .S(n94), .A0(\r_prefetch_data[2][23] ), .A1(n440), .Z(\c_prefetch_data[2][23] ));
Q_MX02 U957 ( .S(n94), .A0(\r_prefetch_data[2][22] ), .A1(n441), .Z(\c_prefetch_data[2][22] ));
Q_MX02 U958 ( .S(n94), .A0(\r_prefetch_data[2][21] ), .A1(n442), .Z(\c_prefetch_data[2][21] ));
Q_MX02 U959 ( .S(n94), .A0(\r_prefetch_data[2][20] ), .A1(n443), .Z(\c_prefetch_data[2][20] ));
Q_MX02 U960 ( .S(n94), .A0(\r_prefetch_data[2][19] ), .A1(n444), .Z(\c_prefetch_data[2][19] ));
Q_MX02 U961 ( .S(n94), .A0(\r_prefetch_data[2][18] ), .A1(n445), .Z(\c_prefetch_data[2][18] ));
Q_MX02 U962 ( .S(n94), .A0(\r_prefetch_data[2][17] ), .A1(n446), .Z(\c_prefetch_data[2][17] ));
Q_MX02 U963 ( .S(n94), .A0(\r_prefetch_data[2][16] ), .A1(n447), .Z(\c_prefetch_data[2][16] ));
Q_MX02 U964 ( .S(n94), .A0(\r_prefetch_data[2][15] ), .A1(n448), .Z(\c_prefetch_data[2][15] ));
Q_MX02 U965 ( .S(n94), .A0(\r_prefetch_data[2][14] ), .A1(n449), .Z(\c_prefetch_data[2][14] ));
Q_MX02 U966 ( .S(n94), .A0(\r_prefetch_data[2][13] ), .A1(n450), .Z(\c_prefetch_data[2][13] ));
Q_MX02 U967 ( .S(n94), .A0(\r_prefetch_data[2][12] ), .A1(n451), .Z(\c_prefetch_data[2][12] ));
Q_MX02 U968 ( .S(n94), .A0(\r_prefetch_data[2][11] ), .A1(n452), .Z(\c_prefetch_data[2][11] ));
Q_MX02 U969 ( .S(n94), .A0(\r_prefetch_data[2][10] ), .A1(n453), .Z(\c_prefetch_data[2][10] ));
Q_MX02 U970 ( .S(n94), .A0(\r_prefetch_data[2][9] ), .A1(n454), .Z(\c_prefetch_data[2][9] ));
Q_MX02 U971 ( .S(n94), .A0(\r_prefetch_data[2][8] ), .A1(n455), .Z(\c_prefetch_data[2][8] ));
Q_MX02 U972 ( .S(n94), .A0(\r_prefetch_data[2][7] ), .A1(n456), .Z(\c_prefetch_data[2][7] ));
Q_MX02 U973 ( .S(n94), .A0(\r_prefetch_data[2][6] ), .A1(n457), .Z(\c_prefetch_data[2][6] ));
Q_MX02 U974 ( .S(n94), .A0(\r_prefetch_data[2][5] ), .A1(n458), .Z(\c_prefetch_data[2][5] ));
Q_MX02 U975 ( .S(n94), .A0(\r_prefetch_data[2][4] ), .A1(n459), .Z(\c_prefetch_data[2][4] ));
Q_MX02 U976 ( .S(n94), .A0(\r_prefetch_data[2][3] ), .A1(n460), .Z(\c_prefetch_data[2][3] ));
Q_MX02 U977 ( .S(n94), .A0(\r_prefetch_data[2][2] ), .A1(n461), .Z(\c_prefetch_data[2][2] ));
Q_MX02 U978 ( .S(n94), .A0(\r_prefetch_data[2][1] ), .A1(n462), .Z(\c_prefetch_data[2][1] ));
Q_MX02 U979 ( .S(n94), .A0(\r_prefetch_data[2][0] ), .A1(n463), .Z(\c_prefetch_data[2][0] ));
Q_MX02 U980 ( .S(n132), .A0(n95), .A1(n392), .Z(c_prefetch_full));
Q_MX02 U981 ( .S(n95), .A0(n826), .A1(r_prefetch_full), .Z(n392));
Q_AN02 U982 ( .A0(prefetch_lden_mem[2]), .A1(mem_ecc_error), .Z(n464));
Q_AN02 U983 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[70]), .Z(n465));
Q_AN02 U984 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[69]), .Z(n466));
Q_AN02 U985 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[68]), .Z(n467));
Q_AN02 U986 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[67]), .Z(n468));
Q_AN02 U987 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[66]), .Z(n469));
Q_AN02 U988 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[65]), .Z(n470));
Q_AN02 U989 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[64]), .Z(n471));
Q_AN02 U990 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[63]), .Z(n472));
Q_AN02 U991 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[62]), .Z(n473));
Q_AN02 U992 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[61]), .Z(n474));
Q_AN02 U993 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[60]), .Z(n475));
Q_AN02 U994 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[59]), .Z(n476));
Q_AN02 U995 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[58]), .Z(n477));
Q_AN02 U996 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[57]), .Z(n478));
Q_AN02 U997 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[56]), .Z(n479));
Q_AN02 U998 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[55]), .Z(n480));
Q_AN02 U999 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[54]), .Z(n481));
Q_AN02 U1000 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[53]), .Z(n482));
Q_AN02 U1001 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[52]), .Z(n483));
Q_AN02 U1002 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[51]), .Z(n484));
Q_AN02 U1003 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[50]), .Z(n485));
Q_AN02 U1004 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[49]), .Z(n486));
Q_AN02 U1005 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[48]), .Z(n487));
Q_AN02 U1006 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[47]), .Z(n488));
Q_AN02 U1007 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[46]), .Z(n489));
Q_AN02 U1008 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[45]), .Z(n490));
Q_AN02 U1009 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[44]), .Z(n491));
Q_AN02 U1010 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[43]), .Z(n492));
Q_AN02 U1011 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[42]), .Z(n493));
Q_AN02 U1012 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[41]), .Z(n494));
Q_AN02 U1013 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[40]), .Z(n495));
Q_AN02 U1014 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[39]), .Z(n496));
Q_AN02 U1015 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[38]), .Z(n497));
Q_AN02 U1016 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[37]), .Z(n498));
Q_AN02 U1017 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[36]), .Z(n499));
Q_AN02 U1018 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[35]), .Z(n500));
Q_AN02 U1019 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[34]), .Z(n501));
Q_AN02 U1020 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[33]), .Z(n502));
Q_AN02 U1021 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[32]), .Z(n503));
Q_AN02 U1022 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[31]), .Z(n504));
Q_AN02 U1023 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[30]), .Z(n505));
Q_AN02 U1024 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[29]), .Z(n506));
Q_AN02 U1025 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[28]), .Z(n507));
Q_AN02 U1026 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[27]), .Z(n508));
Q_AN02 U1027 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[26]), .Z(n509));
Q_AN02 U1028 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[25]), .Z(n510));
Q_AN02 U1029 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[24]), .Z(n511));
Q_AN02 U1030 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[23]), .Z(n512));
Q_AN02 U1031 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[22]), .Z(n513));
Q_AN02 U1032 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[21]), .Z(n514));
Q_AN02 U1033 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[20]), .Z(n515));
Q_AN02 U1034 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[19]), .Z(n516));
Q_AN02 U1035 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[18]), .Z(n517));
Q_AN02 U1036 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[17]), .Z(n518));
Q_AN02 U1037 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[16]), .Z(n519));
Q_AN02 U1038 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[15]), .Z(n520));
Q_AN02 U1039 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[14]), .Z(n521));
Q_AN02 U1040 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[13]), .Z(n522));
Q_AN02 U1041 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[12]), .Z(n523));
Q_AN02 U1042 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[11]), .Z(n524));
Q_AN02 U1043 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[10]), .Z(n525));
Q_AN02 U1044 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[9]), .Z(n526));
Q_AN02 U1045 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[8]), .Z(n527));
Q_AN02 U1046 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[7]), .Z(n528));
Q_AN02 U1047 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[6]), .Z(n529));
Q_AN02 U1048 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[5]), .Z(n530));
Q_AN02 U1049 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[4]), .Z(n531));
Q_AN02 U1050 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[3]), .Z(n532));
Q_AN02 U1051 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[2]), .Z(n533));
Q_AN02 U1052 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[1]), .Z(n534));
Q_AN02 U1053 ( .A0(prefetch_lden_mem[2]), .A1(mem_rdata[0]), .Z(n535));
Q_AO21 U1054 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[70]), .B0(n465), .Z(n393));
Q_AO21 U1055 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[69]), .B0(n466), .Z(n394));
Q_AO21 U1056 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[68]), .B0(n467), .Z(n395));
Q_AO21 U1057 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[67]), .B0(n468), .Z(n396));
Q_AO21 U1058 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[66]), .B0(n469), .Z(n397));
Q_AO21 U1059 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[65]), .B0(n470), .Z(n398));
Q_AO21 U1060 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[64]), .B0(n471), .Z(n399));
Q_AO21 U1061 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[63]), .B0(n472), .Z(n400));
Q_AO21 U1062 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[62]), .B0(n473), .Z(n401));
Q_AO21 U1063 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[61]), .B0(n474), .Z(n402));
Q_AO21 U1064 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[60]), .B0(n475), .Z(n403));
Q_AO21 U1065 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[59]), .B0(n476), .Z(n404));
Q_AO21 U1066 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[58]), .B0(n477), .Z(n405));
Q_AO21 U1067 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[57]), .B0(n478), .Z(n406));
Q_AO21 U1068 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[56]), .B0(n479), .Z(n407));
Q_AO21 U1069 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[55]), .B0(n480), .Z(n408));
Q_AO21 U1070 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[54]), .B0(n481), .Z(n409));
Q_AO21 U1071 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[53]), .B0(n482), .Z(n410));
Q_AO21 U1072 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[52]), .B0(n483), .Z(n411));
Q_AO21 U1073 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[51]), .B0(n484), .Z(n412));
Q_AO21 U1074 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[50]), .B0(n485), .Z(n413));
Q_AO21 U1075 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[49]), .B0(n486), .Z(n414));
Q_AO21 U1076 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[48]), .B0(n487), .Z(n415));
Q_AO21 U1077 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[47]), .B0(n488), .Z(n416));
Q_AO21 U1078 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[46]), .B0(n489), .Z(n417));
Q_AO21 U1079 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[45]), .B0(n490), .Z(n418));
Q_AO21 U1080 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[44]), .B0(n491), .Z(n419));
Q_AO21 U1081 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[43]), .B0(n492), .Z(n420));
Q_AO21 U1082 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[42]), .B0(n493), .Z(n421));
Q_AO21 U1083 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[41]), .B0(n494), .Z(n422));
Q_AO21 U1084 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[40]), .B0(n495), .Z(n423));
Q_AO21 U1085 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[39]), .B0(n496), .Z(n424));
Q_AO21 U1086 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[38]), .B0(n497), .Z(n425));
Q_AO21 U1087 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[37]), .B0(n498), .Z(n426));
Q_AO21 U1088 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[36]), .B0(n499), .Z(n427));
Q_AO21 U1089 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[35]), .B0(n500), .Z(n428));
Q_AO21 U1090 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[34]), .B0(n501), .Z(n429));
Q_AO21 U1091 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[33]), .B0(n502), .Z(n430));
Q_AO21 U1092 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[32]), .B0(n503), .Z(n431));
Q_AO21 U1093 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[31]), .B0(n504), .Z(n432));
Q_AO21 U1094 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[30]), .B0(n505), .Z(n433));
Q_AO21 U1095 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[29]), .B0(n506), .Z(n434));
Q_AO21 U1096 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[28]), .B0(n507), .Z(n435));
Q_AO21 U1097 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[27]), .B0(n508), .Z(n436));
Q_AO21 U1098 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[26]), .B0(n509), .Z(n437));
Q_AO21 U1099 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[25]), .B0(n510), .Z(n438));
Q_AO21 U1100 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[24]), .B0(n511), .Z(n439));
Q_AO21 U1101 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[23]), .B0(n512), .Z(n440));
Q_AO21 U1102 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[22]), .B0(n513), .Z(n441));
Q_AO21 U1103 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[21]), .B0(n514), .Z(n442));
Q_AO21 U1104 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[20]), .B0(n515), .Z(n443));
Q_AO21 U1105 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[19]), .B0(n516), .Z(n444));
Q_AO21 U1106 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[18]), .B0(n517), .Z(n445));
Q_AO21 U1107 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[17]), .B0(n518), .Z(n446));
Q_AO21 U1108 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[16]), .B0(n519), .Z(n447));
Q_AO21 U1109 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[15]), .B0(n520), .Z(n448));
Q_AO21 U1110 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[14]), .B0(n521), .Z(n449));
Q_AO21 U1111 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[13]), .B0(n522), .Z(n450));
Q_AO21 U1112 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[12]), .B0(n523), .Z(n451));
Q_AO21 U1113 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[11]), .B0(n524), .Z(n452));
Q_AO21 U1114 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[10]), .B0(n525), .Z(n453));
Q_AO21 U1115 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[9]), .B0(n526), .Z(n454));
Q_AO21 U1116 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[8]), .B0(n527), .Z(n455));
Q_AO21 U1117 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[7]), .B0(n528), .Z(n456));
Q_AO21 U1118 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[6]), .B0(n529), .Z(n457));
Q_AO21 U1119 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[5]), .B0(n530), .Z(n458));
Q_AO21 U1120 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[4]), .B0(n531), .Z(n459));
Q_AO21 U1121 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[3]), .B0(n532), .Z(n460));
Q_AO21 U1122 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[2]), .B0(n533), .Z(n461));
Q_AO21 U1123 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[1]), .B0(n534), .Z(n462));
Q_AO21 U1124 ( .A0(prefetch_lden_bypass[2]), .A1(wdata[0]), .B0(n535), .Z(n463));
Q_AN02 U1125 ( .A0(prefetch_lden_mem[1]), .A1(mem_ecc_error), .Z(n607));
Q_AN02 U1126 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[70]), .Z(n608));
Q_AN02 U1127 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[69]), .Z(n609));
Q_AN02 U1128 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[68]), .Z(n610));
Q_AN02 U1129 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[67]), .Z(n611));
Q_AN02 U1130 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[66]), .Z(n612));
Q_AN02 U1131 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[65]), .Z(n613));
Q_AN02 U1132 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[64]), .Z(n614));
Q_AN02 U1133 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[63]), .Z(n615));
Q_AN02 U1134 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[62]), .Z(n616));
Q_AN02 U1135 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[61]), .Z(n617));
Q_AN02 U1136 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[60]), .Z(n618));
Q_AN02 U1137 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[59]), .Z(n619));
Q_AN02 U1138 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[58]), .Z(n620));
Q_AN02 U1139 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[57]), .Z(n621));
Q_AN02 U1140 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[56]), .Z(n622));
Q_AN02 U1141 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[55]), .Z(n623));
Q_AN02 U1142 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[54]), .Z(n624));
Q_AN02 U1143 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[53]), .Z(n625));
Q_AN02 U1144 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[52]), .Z(n626));
Q_AN02 U1145 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[51]), .Z(n627));
Q_AN02 U1146 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[50]), .Z(n628));
Q_AN02 U1147 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[49]), .Z(n629));
Q_AN02 U1148 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[48]), .Z(n630));
Q_AN02 U1149 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[47]), .Z(n631));
Q_AN02 U1150 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[46]), .Z(n632));
Q_AN02 U1151 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[45]), .Z(n633));
Q_AN02 U1152 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[44]), .Z(n634));
Q_AN02 U1153 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[43]), .Z(n635));
Q_AN02 U1154 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[42]), .Z(n636));
Q_AN02 U1155 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[41]), .Z(n637));
Q_AN02 U1156 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[40]), .Z(n638));
Q_AN02 U1157 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[39]), .Z(n639));
Q_AN02 U1158 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[38]), .Z(n640));
Q_AN02 U1159 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[37]), .Z(n641));
Q_AN02 U1160 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[36]), .Z(n642));
Q_AN02 U1161 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[35]), .Z(n643));
Q_AN02 U1162 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[34]), .Z(n644));
Q_AN02 U1163 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[33]), .Z(n645));
Q_AN02 U1164 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[32]), .Z(n646));
Q_AN02 U1165 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[31]), .Z(n647));
Q_AN02 U1166 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[30]), .Z(n648));
Q_AN02 U1167 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[29]), .Z(n649));
Q_AN02 U1168 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[28]), .Z(n650));
Q_AN02 U1169 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[27]), .Z(n651));
Q_AN02 U1170 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[26]), .Z(n652));
Q_AN02 U1171 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[25]), .Z(n653));
Q_AN02 U1172 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[24]), .Z(n654));
Q_AN02 U1173 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[23]), .Z(n655));
Q_AN02 U1174 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[22]), .Z(n656));
Q_AN02 U1175 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[21]), .Z(n657));
Q_AN02 U1176 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[20]), .Z(n658));
Q_AN02 U1177 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[19]), .Z(n659));
Q_AN02 U1178 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[18]), .Z(n660));
Q_AN02 U1179 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[17]), .Z(n661));
Q_AN02 U1180 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[16]), .Z(n662));
Q_AN02 U1181 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[15]), .Z(n663));
Q_AN02 U1182 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[14]), .Z(n664));
Q_AN02 U1183 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[13]), .Z(n665));
Q_AN02 U1184 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[12]), .Z(n666));
Q_AN02 U1185 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[11]), .Z(n667));
Q_AN02 U1186 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[10]), .Z(n668));
Q_AN02 U1187 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[9]), .Z(n669));
Q_AN02 U1188 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[8]), .Z(n670));
Q_AN02 U1189 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[7]), .Z(n671));
Q_AN02 U1190 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[6]), .Z(n672));
Q_AN02 U1191 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[5]), .Z(n673));
Q_AN02 U1192 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[4]), .Z(n674));
Q_AN02 U1193 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[3]), .Z(n675));
Q_AN02 U1194 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[2]), .Z(n676));
Q_AN02 U1195 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[1]), .Z(n677));
Q_AN02 U1196 ( .A0(prefetch_lden_mem[1]), .A1(mem_rdata[0]), .Z(n678));
Q_AO21 U1197 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[70]), .B0(n608), .Z(n536));
Q_AO21 U1198 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[69]), .B0(n609), .Z(n537));
Q_AO21 U1199 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[68]), .B0(n610), .Z(n538));
Q_AO21 U1200 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[67]), .B0(n611), .Z(n539));
Q_AO21 U1201 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[66]), .B0(n612), .Z(n540));
Q_AO21 U1202 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[65]), .B0(n613), .Z(n541));
Q_AO21 U1203 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[64]), .B0(n614), .Z(n542));
Q_AO21 U1204 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[63]), .B0(n615), .Z(n543));
Q_AO21 U1205 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[62]), .B0(n616), .Z(n544));
Q_AO21 U1206 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[61]), .B0(n617), .Z(n545));
Q_AO21 U1207 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[60]), .B0(n618), .Z(n546));
Q_AO21 U1208 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[59]), .B0(n619), .Z(n547));
Q_AO21 U1209 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[58]), .B0(n620), .Z(n548));
Q_AO21 U1210 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[57]), .B0(n621), .Z(n549));
Q_AO21 U1211 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[56]), .B0(n622), .Z(n550));
Q_AO21 U1212 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[55]), .B0(n623), .Z(n551));
Q_AO21 U1213 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[54]), .B0(n624), .Z(n552));
Q_AO21 U1214 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[53]), .B0(n625), .Z(n553));
Q_AO21 U1215 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[52]), .B0(n626), .Z(n554));
Q_AO21 U1216 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[51]), .B0(n627), .Z(n555));
Q_AO21 U1217 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[50]), .B0(n628), .Z(n556));
Q_AO21 U1218 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[49]), .B0(n629), .Z(n557));
Q_AO21 U1219 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[48]), .B0(n630), .Z(n558));
Q_AO21 U1220 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[47]), .B0(n631), .Z(n559));
Q_AO21 U1221 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[46]), .B0(n632), .Z(n560));
Q_AO21 U1222 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[45]), .B0(n633), .Z(n561));
Q_AO21 U1223 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[44]), .B0(n634), .Z(n562));
Q_AO21 U1224 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[43]), .B0(n635), .Z(n563));
Q_AO21 U1225 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[42]), .B0(n636), .Z(n564));
Q_AO21 U1226 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[41]), .B0(n637), .Z(n565));
Q_AO21 U1227 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[40]), .B0(n638), .Z(n566));
Q_AO21 U1228 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[39]), .B0(n639), .Z(n567));
Q_AO21 U1229 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[38]), .B0(n640), .Z(n568));
Q_AO21 U1230 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[37]), .B0(n641), .Z(n569));
Q_AO21 U1231 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[36]), .B0(n642), .Z(n570));
Q_AO21 U1232 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[35]), .B0(n643), .Z(n571));
Q_AO21 U1233 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[34]), .B0(n644), .Z(n572));
Q_AO21 U1234 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[33]), .B0(n645), .Z(n573));
Q_AO21 U1235 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[32]), .B0(n646), .Z(n574));
Q_AO21 U1236 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[31]), .B0(n647), .Z(n575));
Q_AO21 U1237 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[30]), .B0(n648), .Z(n576));
Q_AO21 U1238 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[29]), .B0(n649), .Z(n577));
Q_AO21 U1239 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[28]), .B0(n650), .Z(n578));
Q_AO21 U1240 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[27]), .B0(n651), .Z(n579));
Q_AO21 U1241 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[26]), .B0(n652), .Z(n580));
Q_AO21 U1242 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[25]), .B0(n653), .Z(n581));
Q_AO21 U1243 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[24]), .B0(n654), .Z(n582));
Q_AO21 U1244 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[23]), .B0(n655), .Z(n583));
Q_AO21 U1245 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[22]), .B0(n656), .Z(n584));
Q_AO21 U1246 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[21]), .B0(n657), .Z(n585));
Q_AO21 U1247 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[20]), .B0(n658), .Z(n586));
Q_AO21 U1248 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[19]), .B0(n659), .Z(n587));
Q_AO21 U1249 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[18]), .B0(n660), .Z(n588));
Q_AO21 U1250 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[17]), .B0(n661), .Z(n589));
Q_AO21 U1251 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[16]), .B0(n662), .Z(n590));
Q_AO21 U1252 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[15]), .B0(n663), .Z(n591));
Q_AO21 U1253 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[14]), .B0(n664), .Z(n592));
Q_AO21 U1254 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[13]), .B0(n665), .Z(n593));
Q_AO21 U1255 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[12]), .B0(n666), .Z(n594));
Q_AO21 U1256 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[11]), .B0(n667), .Z(n595));
Q_AO21 U1257 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[10]), .B0(n668), .Z(n596));
Q_AO21 U1258 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[9]), .B0(n669), .Z(n597));
Q_AO21 U1259 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[8]), .B0(n670), .Z(n598));
Q_AO21 U1260 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[7]), .B0(n671), .Z(n599));
Q_AO21 U1261 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[6]), .B0(n672), .Z(n600));
Q_AO21 U1262 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[5]), .B0(n673), .Z(n601));
Q_AO21 U1263 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[4]), .B0(n674), .Z(n602));
Q_AO21 U1264 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[3]), .B0(n675), .Z(n603));
Q_AO21 U1265 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[2]), .B0(n676), .Z(n604));
Q_AO21 U1266 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[1]), .B0(n677), .Z(n605));
Q_AO21 U1267 ( .A0(prefetch_lden_bypass[1]), .A1(wdata[0]), .B0(n678), .Z(n606));
Q_AN02 U1268 ( .A0(prefetch_lden_mem[0]), .A1(mem_ecc_error), .Z(n750));
Q_AN02 U1269 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[70]), .Z(n751));
Q_AN02 U1270 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[69]), .Z(n752));
Q_AN02 U1271 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[68]), .Z(n753));
Q_AN02 U1272 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[67]), .Z(n754));
Q_AN02 U1273 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[66]), .Z(n755));
Q_AN02 U1274 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[65]), .Z(n756));
Q_AN02 U1275 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[64]), .Z(n757));
Q_AN02 U1276 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[63]), .Z(n758));
Q_AN02 U1277 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[62]), .Z(n759));
Q_AN02 U1278 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[61]), .Z(n760));
Q_AN02 U1279 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[60]), .Z(n761));
Q_AN02 U1280 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[59]), .Z(n762));
Q_AN02 U1281 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[58]), .Z(n763));
Q_AN02 U1282 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[57]), .Z(n764));
Q_AN02 U1283 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[56]), .Z(n765));
Q_AN02 U1284 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[55]), .Z(n766));
Q_AN02 U1285 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[54]), .Z(n767));
Q_AN02 U1286 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[53]), .Z(n768));
Q_AN02 U1287 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[52]), .Z(n769));
Q_AN02 U1288 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[51]), .Z(n770));
Q_AN02 U1289 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[50]), .Z(n771));
Q_AN02 U1290 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[49]), .Z(n772));
Q_AN02 U1291 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[48]), .Z(n773));
Q_AN02 U1292 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[47]), .Z(n774));
Q_AN02 U1293 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[46]), .Z(n775));
Q_AN02 U1294 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[45]), .Z(n776));
Q_AN02 U1295 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[44]), .Z(n777));
Q_AN02 U1296 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[43]), .Z(n778));
Q_AN02 U1297 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[42]), .Z(n779));
Q_AN02 U1298 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[41]), .Z(n780));
Q_AN02 U1299 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[40]), .Z(n781));
Q_AN02 U1300 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[39]), .Z(n782));
Q_AN02 U1301 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[38]), .Z(n783));
Q_AN02 U1302 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[37]), .Z(n784));
Q_AN02 U1303 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[36]), .Z(n785));
Q_AN02 U1304 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[35]), .Z(n786));
Q_AN02 U1305 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[34]), .Z(n787));
Q_AN02 U1306 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[33]), .Z(n788));
Q_AN02 U1307 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[32]), .Z(n789));
Q_AN02 U1308 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[31]), .Z(n790));
Q_AN02 U1309 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[30]), .Z(n791));
Q_AN02 U1310 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[29]), .Z(n792));
Q_AN02 U1311 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[28]), .Z(n793));
Q_AN02 U1312 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[27]), .Z(n794));
Q_AN02 U1313 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[26]), .Z(n795));
Q_AN02 U1314 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[25]), .Z(n796));
Q_AN02 U1315 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[24]), .Z(n797));
Q_AN02 U1316 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[23]), .Z(n798));
Q_AN02 U1317 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[22]), .Z(n799));
Q_AN02 U1318 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[21]), .Z(n800));
Q_AN02 U1319 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[20]), .Z(n801));
Q_AN02 U1320 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[19]), .Z(n802));
Q_AN02 U1321 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[18]), .Z(n803));
Q_AN02 U1322 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[17]), .Z(n804));
Q_AN02 U1323 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[16]), .Z(n805));
Q_AN02 U1324 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[15]), .Z(n806));
Q_AN02 U1325 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[14]), .Z(n807));
Q_AN02 U1326 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[13]), .Z(n808));
Q_AN02 U1327 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[12]), .Z(n809));
Q_AN02 U1328 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[11]), .Z(n810));
Q_AN02 U1329 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[10]), .Z(n811));
Q_AN02 U1330 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[9]), .Z(n812));
Q_AN02 U1331 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[8]), .Z(n813));
Q_AN02 U1332 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[7]), .Z(n814));
Q_AN02 U1333 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[6]), .Z(n815));
Q_AN02 U1334 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[5]), .Z(n816));
Q_AN02 U1335 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[4]), .Z(n817));
Q_AN02 U1336 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[3]), .Z(n818));
Q_AN02 U1337 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[2]), .Z(n819));
Q_AN02 U1338 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[1]), .Z(n820));
Q_AN02 U1339 ( .A0(prefetch_lden_mem[0]), .A1(mem_rdata[0]), .Z(n821));
Q_AO21 U1340 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[70]), .B0(n751), .Z(n679));
Q_AO21 U1341 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[69]), .B0(n752), .Z(n680));
Q_AO21 U1342 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[68]), .B0(n753), .Z(n681));
Q_AO21 U1343 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[67]), .B0(n754), .Z(n682));
Q_AO21 U1344 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[66]), .B0(n755), .Z(n683));
Q_AO21 U1345 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[65]), .B0(n756), .Z(n684));
Q_AO21 U1346 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[64]), .B0(n757), .Z(n685));
Q_AO21 U1347 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[63]), .B0(n758), .Z(n686));
Q_AO21 U1348 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[62]), .B0(n759), .Z(n687));
Q_AO21 U1349 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[61]), .B0(n760), .Z(n688));
Q_AO21 U1350 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[60]), .B0(n761), .Z(n689));
Q_AO21 U1351 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[59]), .B0(n762), .Z(n690));
Q_AO21 U1352 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[58]), .B0(n763), .Z(n691));
Q_AO21 U1353 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[57]), .B0(n764), .Z(n692));
Q_AO21 U1354 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[56]), .B0(n765), .Z(n693));
Q_AO21 U1355 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[55]), .B0(n766), .Z(n694));
Q_AO21 U1356 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[54]), .B0(n767), .Z(n695));
Q_AO21 U1357 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[53]), .B0(n768), .Z(n696));
Q_AO21 U1358 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[52]), .B0(n769), .Z(n697));
Q_AO21 U1359 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[51]), .B0(n770), .Z(n698));
Q_AO21 U1360 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[50]), .B0(n771), .Z(n699));
Q_AO21 U1361 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[49]), .B0(n772), .Z(n700));
Q_AO21 U1362 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[48]), .B0(n773), .Z(n701));
Q_AO21 U1363 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[47]), .B0(n774), .Z(n702));
Q_AO21 U1364 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[46]), .B0(n775), .Z(n703));
Q_AO21 U1365 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[45]), .B0(n776), .Z(n704));
Q_AO21 U1366 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[44]), .B0(n777), .Z(n705));
Q_AO21 U1367 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[43]), .B0(n778), .Z(n706));
Q_AO21 U1368 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[42]), .B0(n779), .Z(n707));
Q_AO21 U1369 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[41]), .B0(n780), .Z(n708));
Q_AO21 U1370 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[40]), .B0(n781), .Z(n709));
Q_AO21 U1371 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[39]), .B0(n782), .Z(n710));
Q_AO21 U1372 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[38]), .B0(n783), .Z(n711));
Q_AO21 U1373 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[37]), .B0(n784), .Z(n712));
Q_AO21 U1374 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[36]), .B0(n785), .Z(n713));
Q_AO21 U1375 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[35]), .B0(n786), .Z(n714));
Q_AO21 U1376 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[34]), .B0(n787), .Z(n715));
Q_AO21 U1377 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[33]), .B0(n788), .Z(n716));
Q_AO21 U1378 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[32]), .B0(n789), .Z(n717));
Q_AO21 U1379 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[31]), .B0(n790), .Z(n718));
Q_AO21 U1380 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[30]), .B0(n791), .Z(n719));
Q_AO21 U1381 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[29]), .B0(n792), .Z(n720));
Q_AO21 U1382 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[28]), .B0(n793), .Z(n721));
Q_AO21 U1383 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[27]), .B0(n794), .Z(n722));
Q_AO21 U1384 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[26]), .B0(n795), .Z(n723));
Q_AO21 U1385 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[25]), .B0(n796), .Z(n724));
Q_AO21 U1386 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[24]), .B0(n797), .Z(n725));
Q_AO21 U1387 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[23]), .B0(n798), .Z(n726));
Q_AO21 U1388 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[22]), .B0(n799), .Z(n727));
Q_AO21 U1389 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[21]), .B0(n800), .Z(n728));
Q_AO21 U1390 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[20]), .B0(n801), .Z(n729));
Q_AO21 U1391 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[19]), .B0(n802), .Z(n730));
Q_AO21 U1392 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[18]), .B0(n803), .Z(n731));
Q_AO21 U1393 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[17]), .B0(n804), .Z(n732));
Q_AO21 U1394 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[16]), .B0(n805), .Z(n733));
Q_AO21 U1395 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[15]), .B0(n806), .Z(n734));
Q_AO21 U1396 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[14]), .B0(n807), .Z(n735));
Q_AO21 U1397 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[13]), .B0(n808), .Z(n736));
Q_AO21 U1398 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[12]), .B0(n809), .Z(n737));
Q_AO21 U1399 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[11]), .B0(n810), .Z(n738));
Q_AO21 U1400 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[10]), .B0(n811), .Z(n739));
Q_AO21 U1401 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[9]), .B0(n812), .Z(n740));
Q_AO21 U1402 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[8]), .B0(n813), .Z(n741));
Q_AO21 U1403 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[7]), .B0(n814), .Z(n742));
Q_AO21 U1404 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[6]), .B0(n815), .Z(n743));
Q_AO21 U1405 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[5]), .B0(n816), .Z(n744));
Q_AO21 U1406 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[4]), .B0(n817), .Z(n745));
Q_AO21 U1407 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[3]), .B0(n818), .Z(n746));
Q_AO21 U1408 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[2]), .B0(n819), .Z(n747));
Q_AO21 U1409 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[1]), .B0(n820), .Z(n748));
Q_AO21 U1410 ( .A0(prefetch_lden_bypass[0]), .A1(wdata[0]), .B0(n821), .Z(n749));
Q_OR02 U1411 ( .A0(prefetch_lden_bypass[2]), .A1(prefetch_lden_mem[2]), .Z(n94));
Q_OR02 U1412 ( .A0(prefetch_lden_bypass[1]), .A1(prefetch_lden_mem[1]), .Z(n93));
Q_OR02 U1413 ( .A0(prefetch_lden_bypass[0]), .A1(prefetch_lden_mem[0]), .Z(n92));
Q_AN02 U1414 ( .A0(n98), .A1(\c_mem_prefetch_wptr_dly[0][2] ), .Z(prefetch_lden_bypass[2]));
Q_AN02 U1415 ( .A0(n98), .A1(\c_mem_prefetch_wptr_dly[0][1] ), .Z(prefetch_lden_bypass[1]));
Q_AN02 U1416 ( .A0(n98), .A1(\c_mem_prefetch_wptr_dly[0][0] ), .Z(prefetch_lden_bypass[0]));
Q_AN02 U1417 ( .A0(n139), .A1(n822), .Z(prefetch_lden_mem[2]));
Q_AN02 U1418 ( .A0(n139), .A1(n823), .Z(prefetch_lden_mem[1]));
Q_AN02 U1419 ( .A0(n139), .A1(n824), .Z(prefetch_lden_mem[0]));
Q_MX03 U1420 ( .S0(r_prefetch_rptr[0]), .S1(r_prefetch_rptr[1]), .A0(n824), .A1(n823), .A2(n822), .Z(n74));
Q_AN02 U1421 ( .A0(r_mem_ren_dly[2]), .A1(\r_mem_prefetch_wptr_dly[2][2] ), .Z(n822));
Q_AN02 U1422 ( .A0(r_mem_ren_dly[2]), .A1(\r_mem_prefetch_wptr_dly[2][1] ), .Z(n823));
Q_AN02 U1423 ( .A0(r_mem_ren_dly[2]), .A1(\r_mem_prefetch_wptr_dly[2][0] ), .Z(n824));
Q_AN02 U1424 ( .A0(r_mem_empty), .A1(n825), .Z(n80));
Q_NR02 U1425 ( .A0(n826), .A1(r_mem_empty), .Z(mem_ren));
Q_INV U1426 ( .A(n826), .Z(n825));
Q_AN02 U1427 ( .A0(n99), .A1(r_prefetch_full), .Z(n826));
Q_ND03 U1428 ( .A0(n829), .A1(n828), .A2(n827), .Z(n76));
Q_AN03 U1429 ( .A0(r_mem_wptr[1]), .A1(r_mem_wptr[0]), .A2(n830), .Z(n827));
Q_AN03 U1430 ( .A0(r_mem_wptr[4]), .A1(r_mem_wptr[3]), .A2(r_mem_wptr[2]), .Z(n828));
Q_AN03 U1431 ( .A0(r_mem_wptr[7]), .A1(r_mem_wptr[6]), .A2(r_mem_wptr[5]), .Z(n829));
Q_AN03 U1432 ( .A0(r_mem_wptr[10]), .A1(r_mem_wptr[9]), .A2(r_mem_wptr[8]), .Z(n830));
Q_ND03 U1433 ( .A0(n833), .A1(n832), .A2(n831), .Z(n78));
Q_AN03 U1434 ( .A0(r_mem_rptr[1]), .A1(r_mem_rptr[0]), .A2(n834), .Z(n831));
Q_AN03 U1435 ( .A0(r_mem_rptr[4]), .A1(r_mem_rptr[3]), .A2(r_mem_rptr[2]), .Z(n832));
Q_AN03 U1436 ( .A0(r_mem_rptr[7]), .A1(r_mem_rptr[6]), .A2(r_mem_rptr[5]), .Z(n833));
Q_AN03 U1437 ( .A0(r_mem_rptr[10]), .A1(r_mem_rptr[9]), .A2(r_mem_rptr[8]), .Z(n834));
Q_AN02 U1438 ( .A0(n835), .A1(r_prefetch_rptr[1]), .Z(n79));
Q_INV U1439 ( .A(_zy_sva_sf1hot_0), .Z(n837));
Q_AN02 U1440 ( .A0(rst_n), .A1(n837), .Z(n836));
ixc_assign_12 _zz_strnp_0 ( used_slots[11:0], r_used_slots[11:0]);
ixc_assign_12 _zz_strnp_1 ( free_slots[11:0], r_free_slots[11:0]);
ixc_assign_11 _zz_strnp_2 ( mem_waddr[10:0], r_mem_wptr[10:0]);
ixc_assign_11 _zz_strnp_3 ( mem_raddr[10:0], r_mem_rptr[10:0]);
ixc_assign_71 _zz_strnp_4 ( mem_wdata[70:0], wdata[70:0]);
ixc_assign _zz_strnp_5 ( empty, r_prefetch_empty);
ixc_assign _zz_strnp_6 ( full, r_mem_full);
ixc_assign _zz_strnp_7 ( _zy_simnet_mem_wen_0_w$, mem_wen);
ixc_assign_11 _zz_strnp_8 ( _zy_simnet_mem_waddr_1_w$[0:10], mem_waddr[10:0]);
ixc_assign_71 _zz_strnp_9 ( _zy_simnet_mem_wdata_2_w$[0:70], mem_wdata[70:0]);
ixc_assign _zz_strnp_10 ( _zy_simnet_mem_ren_3_w$, mem_ren);
ixc_assign_11 _zz_strnp_11 ( _zy_simnet_mem_raddr_4_w$[0:10], mem_raddr[10:0]);
ixc_assign _zz_strnp_12 ( _zy_simnet_empty_5_w$, empty);
ixc_assign _zz_strnp_13 ( _zy_simnet_full_6_w$, full);
ixc_assign_12 _zz_strnp_14 ( _zy_simnet_used_slots_7_w$[0:11], 
	used_slots[11:0]);
ixc_assign_12 _zz_strnp_15 ( _zy_simnet_free_slots_8_w$[0:11], 
	free_slots[11:0]);
ixc_assign _zz_strnp_16 ( _zy_simnet_rerr_9_w$, rerr);
ixc_assign_71 _zz_strnp_17 ( _zy_simnet_rdata_10_w$[0:70], rdata[70:0]);
ixc_assign _zz_strnp_18 ( _zy_simnet_underflow_11_w$, underflow);
ixc_assign _zz_strnp_19 ( _zy_simnet_overflow_12_w$, overflow);
Q_INV U1461 ( .A(rst_n), .Z(_zy_sva__asrtLbl279_1_reset_or));
Q_AO21 U1462 ( .A0(_zy_sva_b0[1]), .A1(_zy_sva_b0[2]), .B0(n844), .Z(n843));
Q_XOR2 U1463 ( .A0(_zy_sva_b0[1]), .A1(_zy_sva_b0[2]), .Z(n845));
Q_AN02 U1464 ( .A0(_zy_sva_b0[0]), .A1(n845), .Z(n844));
Q_XOR2 U1465 ( .A0(_zy_sva_b0[0]), .A1(n845), .Z(n842));
Q_INV U1466 ( .A(n843), .Z(n841));
Q_AN02 U1467 ( .A0(n841), .A1(n842), .Z(_zy_sva_sf1hot_0));
ixc_sample_logic_3_3 _zz_zy_sva_b0 ( _zy_sva_b0[2:0], { 
	\c_mem_prefetch_wptr_dly[0][2] , \c_mem_prefetch_wptr_dly[0][1] , 
	\c_mem_prefetch_wptr_dly[0][0] });
ixc_pio_call_0_0_0_0_1 _zzixc_tfport_1_0 ( _zyixc_port_1_0_ack, 
	_zyixc_port_1_0_s2hW, _zyixc_port_1_0_isf, _zyixc_port_1_0_req, n840, 
	_zyixc_port_1_0_osf, n839, n1);
wire [2:0] n848 = 3'b000;
Q_ASSERT _asrtLbl279 ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT( ), .FAIL_COUNT( ), .CHECK_COUNT( ), .KILL_SIGNAL( ), .SEVERITY(n848[0]));
// pragma CVASTRPROP INSTANCE "_asrtLbl279" HDL_ASSERT "$"
// pragma CVASTRPROP INSTANCE "_asrtLbl279" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/common/nx_library/nx_fifo_ctrl_ram_1r1w.v"
//pragma CVAINTPROP INSTANCE "_asrtLbl279" ASSERT_LINE 279
Q_AN02 U1471 ( .A0(r_free_slots[1]), .A1(r_free_slots[0]), .Z(n390));
Q_AN02 U1472 ( .A0(r_used_slots[1]), .A1(r_used_slots[0]), .Z(n369));
Q_XOR2 U1473 ( .A0(mem_ren), .A1(r_mem_rptr[0]), .Z(n223));
Q_XNR2 U1474 ( .A0(n125), .A1(n194), .Z(n192));
Q_XNR2 U1475 ( .A0(n103), .A1(n349), .Z(n161));
Q_XOR2 U1476 ( .A0(n114), .A1(n121), .Z(n100));
Q_INV U1477 ( .A(_zy_sva__asrtLbl279_1_1_fail[0]), .Z(n846));
Q_FDP4EP \_zy_sva__asrtLbl279_1_1_fail_REG[0] ( .CK(clk), .CE(n836), .R(n838), .D(n846), .Q(_zy_sva__asrtLbl279_1_1_fail[0]));
Q_INV U1479 ( .A(_zyixc_port_1_0_req), .Z(n847));
Q_FDP4EP _zyixc_port_1_0_req_REG  ( .CK(clk), .CE(n836), .R(n838), .D(n847), .Q(_zyixc_port_1_0_req));
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m1 "r_mem_prefetch_wptr_dly 1 2 0 2 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m2 "c_mem_prefetch_wptr_dly 1 2 0 2 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m3 "r_prefetch_data 1 71 0 2 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m4 "c_prefetch_data 1 71 0 2 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_NON_CMM "4"
// pragma CVASTRPROP MODULE HDLICE PROP_RANOFF TRUE
endmodule
