
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
(* celldefine = 1 *) 
module nx_roreg_indirect_access_xcm131 ( stat_code, stat_datawords, stat_addr, 
	capability_lst, capability_type, rd_dat, clk, rst_n, addr, cmnd_op, 
	cmnd_addr, wr_stb, wr_dat, .mem_a( {\mem_a[0][63] , \mem_a[0][62] , 
	\mem_a[0][61] , \mem_a[0][60] , \mem_a[0][59] , \mem_a[0][58] , 
	\mem_a[0][57] , \mem_a[0][56] , \mem_a[0][55] , \mem_a[0][54] , 
	\mem_a[0][53] , \mem_a[0][52] , \mem_a[0][51] , \mem_a[0][50] , 
	\mem_a[0][49] , \mem_a[0][48] , \mem_a[0][47] , \mem_a[0][46] , 
	\mem_a[0][45] , \mem_a[0][44] , \mem_a[0][43] , \mem_a[0][42] , 
	\mem_a[0][41] , \mem_a[0][40] , \mem_a[0][39] , \mem_a[0][38] , 
	\mem_a[0][37] , \mem_a[0][36] , \mem_a[0][35] , \mem_a[0][34] , 
	\mem_a[0][33] , \mem_a[0][32] , \mem_a[0][31] , \mem_a[0][30] , 
	\mem_a[0][29] , \mem_a[0][28] , \mem_a[0][27] , \mem_a[0][26] , 
	\mem_a[0][25] , \mem_a[0][24] , \mem_a[0][23] , \mem_a[0][22] , 
	\mem_a[0][21] , \mem_a[0][20] , \mem_a[0][19] , \mem_a[0][18] , 
	\mem_a[0][17] , \mem_a[0][16] , \mem_a[0][15] , \mem_a[0][14] , 
	\mem_a[0][13] , \mem_a[0][12] , \mem_a[0][11] , \mem_a[0][10] , 
	\mem_a[0][9] , \mem_a[0][8] , \mem_a[0][7] , \mem_a[0][6] , 
	\mem_a[0][5] , \mem_a[0][4] , \mem_a[0][3] , \mem_a[0][2] , 
	\mem_a[0][1] , \mem_a[0][0] , \mem_a[1][63] , \mem_a[1][62] , 
	\mem_a[1][61] , \mem_a[1][60] , \mem_a[1][59] , \mem_a[1][58] , 
	\mem_a[1][57] , \mem_a[1][56] , \mem_a[1][55] , \mem_a[1][54] , 
	\mem_a[1][53] , \mem_a[1][52] , \mem_a[1][51] , \mem_a[1][50] , 
	\mem_a[1][49] , \mem_a[1][48] , \mem_a[1][47] , \mem_a[1][46] , 
	\mem_a[1][45] , \mem_a[1][44] , \mem_a[1][43] , \mem_a[1][42] , 
	\mem_a[1][41] , \mem_a[1][40] , \mem_a[1][39] , \mem_a[1][38] , 
	\mem_a[1][37] , \mem_a[1][36] , \mem_a[1][35] , \mem_a[1][34] , 
	\mem_a[1][33] , \mem_a[1][32] , \mem_a[1][31] , \mem_a[1][30] , 
	\mem_a[1][29] , \mem_a[1][28] , \mem_a[1][27] , \mem_a[1][26] , 
	\mem_a[1][25] , \mem_a[1][24] , \mem_a[1][23] , \mem_a[1][22] , 
	\mem_a[1][21] , \mem_a[1][20] , \mem_a[1][19] , \mem_a[1][18] , 
	\mem_a[1][17] , \mem_a[1][16] , \mem_a[1][15] , \mem_a[1][14] , 
	\mem_a[1][13] , \mem_a[1][12] , \mem_a[1][11] , \mem_a[1][10] , 
	\mem_a[1][9] , \mem_a[1][8] , \mem_a[1][7] , \mem_a[1][6] , 
	\mem_a[1][5] , \mem_a[1][4] , \mem_a[1][3] , \mem_a[1][2] , 
	\mem_a[1][1] , \mem_a[1][0] , \mem_a[2][63] , \mem_a[2][62] , 
	\mem_a[2][61] , \mem_a[2][60] , \mem_a[2][59] , \mem_a[2][58] , 
	\mem_a[2][57] , \mem_a[2][56] , \mem_a[2][55] , \mem_a[2][54] , 
	\mem_a[2][53] , \mem_a[2][52] , \mem_a[2][51] , \mem_a[2][50] , 
	\mem_a[2][49] , \mem_a[2][48] , \mem_a[2][47] , \mem_a[2][46] , 
	\mem_a[2][45] , \mem_a[2][44] , \mem_a[2][43] , \mem_a[2][42] , 
	\mem_a[2][41] , \mem_a[2][40] , \mem_a[2][39] , \mem_a[2][38] , 
	\mem_a[2][37] , \mem_a[2][36] , \mem_a[2][35] , \mem_a[2][34] , 
	\mem_a[2][33] , \mem_a[2][32] , \mem_a[2][31] , \mem_a[2][30] , 
	\mem_a[2][29] , \mem_a[2][28] , \mem_a[2][27] , \mem_a[2][26] , 
	\mem_a[2][25] , \mem_a[2][24] , \mem_a[2][23] , \mem_a[2][22] , 
	\mem_a[2][21] , \mem_a[2][20] , \mem_a[2][19] , \mem_a[2][18] , 
	\mem_a[2][17] , \mem_a[2][16] , \mem_a[2][15] , \mem_a[2][14] , 
	\mem_a[2][13] , \mem_a[2][12] , \mem_a[2][11] , \mem_a[2][10] , 
	\mem_a[2][9] , \mem_a[2][8] , \mem_a[2][7] , \mem_a[2][6] , 
	\mem_a[2][5] , \mem_a[2][4] , \mem_a[2][3] , \mem_a[2][2] , 
	\mem_a[2][1] , \mem_a[2][0] , \mem_a[3][63] , \mem_a[3][62] , 
	\mem_a[3][61] , \mem_a[3][60] , \mem_a[3][59] , \mem_a[3][58] , 
	\mem_a[3][57] , \mem_a[3][56] , \mem_a[3][55] , \mem_a[3][54] , 
	\mem_a[3][53] , \mem_a[3][52] , \mem_a[3][51] , \mem_a[3][50] , 
	\mem_a[3][49] , \mem_a[3][48] , \mem_a[3][47] , \mem_a[3][46] , 
	\mem_a[3][45] , \mem_a[3][44] , \mem_a[3][43] , \mem_a[3][42] , 
	\mem_a[3][41] , \mem_a[3][40] , \mem_a[3][39] , \mem_a[3][38] , 
	\mem_a[3][37] , \mem_a[3][36] , \mem_a[3][35] , \mem_a[3][34] , 
	\mem_a[3][33] , \mem_a[3][32] , \mem_a[3][31] , \mem_a[3][30] , 
	\mem_a[3][29] , \mem_a[3][28] , \mem_a[3][27] , \mem_a[3][26] , 
	\mem_a[3][25] , \mem_a[3][24] , \mem_a[3][23] , \mem_a[3][22] , 
	\mem_a[3][21] , \mem_a[3][20] , \mem_a[3][19] , \mem_a[3][18] , 
	\mem_a[3][17] , \mem_a[3][16] , \mem_a[3][15] , \mem_a[3][14] , 
	\mem_a[3][13] , \mem_a[3][12] , \mem_a[3][11] , \mem_a[3][10] , 
	\mem_a[3][9] , \mem_a[3][8] , \mem_a[3][7] , \mem_a[3][6] , 
	\mem_a[3][5] , \mem_a[3][4] , \mem_a[3][3] , \mem_a[3][2] , 
	\mem_a[3][1] , \mem_a[3][0] , \mem_a[4][63] , \mem_a[4][62] , 
	\mem_a[4][61] , \mem_a[4][60] , \mem_a[4][59] , \mem_a[4][58] , 
	\mem_a[4][57] , \mem_a[4][56] , \mem_a[4][55] , \mem_a[4][54] , 
	\mem_a[4][53] , \mem_a[4][52] , \mem_a[4][51] , \mem_a[4][50] , 
	\mem_a[4][49] , \mem_a[4][48] , \mem_a[4][47] , \mem_a[4][46] , 
	\mem_a[4][45] , \mem_a[4][44] , \mem_a[4][43] , \mem_a[4][42] , 
	\mem_a[4][41] , \mem_a[4][40] , \mem_a[4][39] , \mem_a[4][38] , 
	\mem_a[4][37] , \mem_a[4][36] , \mem_a[4][35] , \mem_a[4][34] , 
	\mem_a[4][33] , \mem_a[4][32] , \mem_a[4][31] , \mem_a[4][30] , 
	\mem_a[4][29] , \mem_a[4][28] , \mem_a[4][27] , \mem_a[4][26] , 
	\mem_a[4][25] , \mem_a[4][24] , \mem_a[4][23] , \mem_a[4][22] , 
	\mem_a[4][21] , \mem_a[4][20] , \mem_a[4][19] , \mem_a[4][18] , 
	\mem_a[4][17] , \mem_a[4][16] , \mem_a[4][15] , \mem_a[4][14] , 
	\mem_a[4][13] , \mem_a[4][12] , \mem_a[4][11] , \mem_a[4][10] , 
	\mem_a[4][9] , \mem_a[4][8] , \mem_a[4][7] , \mem_a[4][6] , 
	\mem_a[4][5] , \mem_a[4][4] , \mem_a[4][3] , \mem_a[4][2] , 
	\mem_a[4][1] , \mem_a[4][0] , \mem_a[5][63] , \mem_a[5][62] , 
	\mem_a[5][61] , \mem_a[5][60] , \mem_a[5][59] , \mem_a[5][58] , 
	\mem_a[5][57] , \mem_a[5][56] , \mem_a[5][55] , \mem_a[5][54] , 
	\mem_a[5][53] , \mem_a[5][52] , \mem_a[5][51] , \mem_a[5][50] , 
	\mem_a[5][49] , \mem_a[5][48] , \mem_a[5][47] , \mem_a[5][46] , 
	\mem_a[5][45] , \mem_a[5][44] , \mem_a[5][43] , \mem_a[5][42] , 
	\mem_a[5][41] , \mem_a[5][40] , \mem_a[5][39] , \mem_a[5][38] , 
	\mem_a[5][37] , \mem_a[5][36] , \mem_a[5][35] , \mem_a[5][34] , 
	\mem_a[5][33] , \mem_a[5][32] , \mem_a[5][31] , \mem_a[5][30] , 
	\mem_a[5][29] , \mem_a[5][28] , \mem_a[5][27] , \mem_a[5][26] , 
	\mem_a[5][25] , \mem_a[5][24] , \mem_a[5][23] , \mem_a[5][22] , 
	\mem_a[5][21] , \mem_a[5][20] , \mem_a[5][19] , \mem_a[5][18] , 
	\mem_a[5][17] , \mem_a[5][16] , \mem_a[5][15] , \mem_a[5][14] , 
	\mem_a[5][13] , \mem_a[5][12] , \mem_a[5][11] , \mem_a[5][10] , 
	\mem_a[5][9] , \mem_a[5][8] , \mem_a[5][7] , \mem_a[5][6] , 
	\mem_a[5][5] , \mem_a[5][4] , \mem_a[5][3] , \mem_a[5][2] , 
	\mem_a[5][1] , \mem_a[5][0] , \mem_a[6][63] , \mem_a[6][62] , 
	\mem_a[6][61] , \mem_a[6][60] , \mem_a[6][59] , \mem_a[6][58] , 
	\mem_a[6][57] , \mem_a[6][56] , \mem_a[6][55] , \mem_a[6][54] , 
	\mem_a[6][53] , \mem_a[6][52] , \mem_a[6][51] , \mem_a[6][50] , 
	\mem_a[6][49] , \mem_a[6][48] , \mem_a[6][47] , \mem_a[6][46] , 
	\mem_a[6][45] , \mem_a[6][44] , \mem_a[6][43] , \mem_a[6][42] , 
	\mem_a[6][41] , \mem_a[6][40] , \mem_a[6][39] , \mem_a[6][38] , 
	\mem_a[6][37] , \mem_a[6][36] , \mem_a[6][35] , \mem_a[6][34] , 
	\mem_a[6][33] , \mem_a[6][32] , \mem_a[6][31] , \mem_a[6][30] , 
	\mem_a[6][29] , \mem_a[6][28] , \mem_a[6][27] , \mem_a[6][26] , 
	\mem_a[6][25] , \mem_a[6][24] , \mem_a[6][23] , \mem_a[6][22] , 
	\mem_a[6][21] , \mem_a[6][20] , \mem_a[6][19] , \mem_a[6][18] , 
	\mem_a[6][17] , \mem_a[6][16] , \mem_a[6][15] , \mem_a[6][14] , 
	\mem_a[6][13] , \mem_a[6][12] , \mem_a[6][11] , \mem_a[6][10] , 
	\mem_a[6][9] , \mem_a[6][8] , \mem_a[6][7] , \mem_a[6][6] , 
	\mem_a[6][5] , \mem_a[6][4] , \mem_a[6][3] , \mem_a[6][2] , 
	\mem_a[6][1] , \mem_a[6][0] , \mem_a[7][63] , \mem_a[7][62] , 
	\mem_a[7][61] , \mem_a[7][60] , \mem_a[7][59] , \mem_a[7][58] , 
	\mem_a[7][57] , \mem_a[7][56] , \mem_a[7][55] , \mem_a[7][54] , 
	\mem_a[7][53] , \mem_a[7][52] , \mem_a[7][51] , \mem_a[7][50] , 
	\mem_a[7][49] , \mem_a[7][48] , \mem_a[7][47] , \mem_a[7][46] , 
	\mem_a[7][45] , \mem_a[7][44] , \mem_a[7][43] , \mem_a[7][42] , 
	\mem_a[7][41] , \mem_a[7][40] , \mem_a[7][39] , \mem_a[7][38] , 
	\mem_a[7][37] , \mem_a[7][36] , \mem_a[7][35] , \mem_a[7][34] , 
	\mem_a[7][33] , \mem_a[7][32] , \mem_a[7][31] , \mem_a[7][30] , 
	\mem_a[7][29] , \mem_a[7][28] , \mem_a[7][27] , \mem_a[7][26] , 
	\mem_a[7][25] , \mem_a[7][24] , \mem_a[7][23] , \mem_a[7][22] , 
	\mem_a[7][21] , \mem_a[7][20] , \mem_a[7][19] , \mem_a[7][18] , 
	\mem_a[7][17] , \mem_a[7][16] , \mem_a[7][15] , \mem_a[7][14] , 
	\mem_a[7][13] , \mem_a[7][12] , \mem_a[7][11] , \mem_a[7][10] , 
	\mem_a[7][9] , \mem_a[7][8] , \mem_a[7][7] , \mem_a[7][6] , 
	\mem_a[7][5] , \mem_a[7][4] , \mem_a[7][3] , \mem_a[7][2] , 
	\mem_a[7][1] , \mem_a[7][0] , \mem_a[8][63] , \mem_a[8][62] , 
	\mem_a[8][61] , \mem_a[8][60] , \mem_a[8][59] , \mem_a[8][58] , 
	\mem_a[8][57] , \mem_a[8][56] , \mem_a[8][55] , \mem_a[8][54] , 
	\mem_a[8][53] , \mem_a[8][52] , \mem_a[8][51] , \mem_a[8][50] , 
	\mem_a[8][49] , \mem_a[8][48] , \mem_a[8][47] , \mem_a[8][46] , 
	\mem_a[8][45] , \mem_a[8][44] , \mem_a[8][43] , \mem_a[8][42] , 
	\mem_a[8][41] , \mem_a[8][40] , \mem_a[8][39] , \mem_a[8][38] , 
	\mem_a[8][37] , \mem_a[8][36] , \mem_a[8][35] , \mem_a[8][34] , 
	\mem_a[8][33] , \mem_a[8][32] , \mem_a[8][31] , \mem_a[8][30] , 
	\mem_a[8][29] , \mem_a[8][28] , \mem_a[8][27] , \mem_a[8][26] , 
	\mem_a[8][25] , \mem_a[8][24] , \mem_a[8][23] , \mem_a[8][22] , 
	\mem_a[8][21] , \mem_a[8][20] , \mem_a[8][19] , \mem_a[8][18] , 
	\mem_a[8][17] , \mem_a[8][16] , \mem_a[8][15] , \mem_a[8][14] , 
	\mem_a[8][13] , \mem_a[8][12] , \mem_a[8][11] , \mem_a[8][10] , 
	\mem_a[8][9] , \mem_a[8][8] , \mem_a[8][7] , \mem_a[8][6] , 
	\mem_a[8][5] , \mem_a[8][4] , \mem_a[8][3] , \mem_a[8][2] , 
	\mem_a[8][1] , \mem_a[8][0] , \mem_a[9][63] , \mem_a[9][62] , 
	\mem_a[9][61] , \mem_a[9][60] , \mem_a[9][59] , \mem_a[9][58] , 
	\mem_a[9][57] , \mem_a[9][56] , \mem_a[9][55] , \mem_a[9][54] , 
	\mem_a[9][53] , \mem_a[9][52] , \mem_a[9][51] , \mem_a[9][50] , 
	\mem_a[9][49] , \mem_a[9][48] , \mem_a[9][47] , \mem_a[9][46] , 
	\mem_a[9][45] , \mem_a[9][44] , \mem_a[9][43] , \mem_a[9][42] , 
	\mem_a[9][41] , \mem_a[9][40] , \mem_a[9][39] , \mem_a[9][38] , 
	\mem_a[9][37] , \mem_a[9][36] , \mem_a[9][35] , \mem_a[9][34] , 
	\mem_a[9][33] , \mem_a[9][32] , \mem_a[9][31] , \mem_a[9][30] , 
	\mem_a[9][29] , \mem_a[9][28] , \mem_a[9][27] , \mem_a[9][26] , 
	\mem_a[9][25] , \mem_a[9][24] , \mem_a[9][23] , \mem_a[9][22] , 
	\mem_a[9][21] , \mem_a[9][20] , \mem_a[9][19] , \mem_a[9][18] , 
	\mem_a[9][17] , \mem_a[9][16] , \mem_a[9][15] , \mem_a[9][14] , 
	\mem_a[9][13] , \mem_a[9][12] , \mem_a[9][11] , \mem_a[9][10] , 
	\mem_a[9][9] , \mem_a[9][8] , \mem_a[9][7] , \mem_a[9][6] , 
	\mem_a[9][5] , \mem_a[9][4] , \mem_a[9][3] , \mem_a[9][2] , 
	\mem_a[9][1] , \mem_a[9][0] , \mem_a[10][63] , \mem_a[10][62] , 
	\mem_a[10][61] , \mem_a[10][60] , \mem_a[10][59] , \mem_a[10][58] , 
	\mem_a[10][57] , \mem_a[10][56] , \mem_a[10][55] , \mem_a[10][54] , 
	\mem_a[10][53] , \mem_a[10][52] , \mem_a[10][51] , \mem_a[10][50] , 
	\mem_a[10][49] , \mem_a[10][48] , \mem_a[10][47] , \mem_a[10][46] , 
	\mem_a[10][45] , \mem_a[10][44] , \mem_a[10][43] , \mem_a[10][42] , 
	\mem_a[10][41] , \mem_a[10][40] , \mem_a[10][39] , \mem_a[10][38] , 
	\mem_a[10][37] , \mem_a[10][36] , \mem_a[10][35] , \mem_a[10][34] , 
	\mem_a[10][33] , \mem_a[10][32] , \mem_a[10][31] , \mem_a[10][30] , 
	\mem_a[10][29] , \mem_a[10][28] , \mem_a[10][27] , \mem_a[10][26] , 
	\mem_a[10][25] , \mem_a[10][24] , \mem_a[10][23] , \mem_a[10][22] , 
	\mem_a[10][21] , \mem_a[10][20] , \mem_a[10][19] , \mem_a[10][18] , 
	\mem_a[10][17] , \mem_a[10][16] , \mem_a[10][15] , \mem_a[10][14] , 
	\mem_a[10][13] , \mem_a[10][12] , \mem_a[10][11] , \mem_a[10][10] , 
	\mem_a[10][9] , \mem_a[10][8] , \mem_a[10][7] , \mem_a[10][6] , 
	\mem_a[10][5] , \mem_a[10][4] , \mem_a[10][3] , \mem_a[10][2] , 
	\mem_a[10][1] , \mem_a[10][0] , \mem_a[11][63] , \mem_a[11][62] , 
	\mem_a[11][61] , \mem_a[11][60] , \mem_a[11][59] , \mem_a[11][58] , 
	\mem_a[11][57] , \mem_a[11][56] , \mem_a[11][55] , \mem_a[11][54] , 
	\mem_a[11][53] , \mem_a[11][52] , \mem_a[11][51] , \mem_a[11][50] , 
	\mem_a[11][49] , \mem_a[11][48] , \mem_a[11][47] , \mem_a[11][46] , 
	\mem_a[11][45] , \mem_a[11][44] , \mem_a[11][43] , \mem_a[11][42] , 
	\mem_a[11][41] , \mem_a[11][40] , \mem_a[11][39] , \mem_a[11][38] , 
	\mem_a[11][37] , \mem_a[11][36] , \mem_a[11][35] , \mem_a[11][34] , 
	\mem_a[11][33] , \mem_a[11][32] , \mem_a[11][31] , \mem_a[11][30] , 
	\mem_a[11][29] , \mem_a[11][28] , \mem_a[11][27] , \mem_a[11][26] , 
	\mem_a[11][25] , \mem_a[11][24] , \mem_a[11][23] , \mem_a[11][22] , 
	\mem_a[11][21] , \mem_a[11][20] , \mem_a[11][19] , \mem_a[11][18] , 
	\mem_a[11][17] , \mem_a[11][16] , \mem_a[11][15] , \mem_a[11][14] , 
	\mem_a[11][13] , \mem_a[11][12] , \mem_a[11][11] , \mem_a[11][10] , 
	\mem_a[11][9] , \mem_a[11][8] , \mem_a[11][7] , \mem_a[11][6] , 
	\mem_a[11][5] , \mem_a[11][4] , \mem_a[11][3] , \mem_a[11][2] , 
	\mem_a[11][1] , \mem_a[11][0] , \mem_a[12][63] , \mem_a[12][62] , 
	\mem_a[12][61] , \mem_a[12][60] , \mem_a[12][59] , \mem_a[12][58] , 
	\mem_a[12][57] , \mem_a[12][56] , \mem_a[12][55] , \mem_a[12][54] , 
	\mem_a[12][53] , \mem_a[12][52] , \mem_a[12][51] , \mem_a[12][50] , 
	\mem_a[12][49] , \mem_a[12][48] , \mem_a[12][47] , \mem_a[12][46] , 
	\mem_a[12][45] , \mem_a[12][44] , \mem_a[12][43] , \mem_a[12][42] , 
	\mem_a[12][41] , \mem_a[12][40] , \mem_a[12][39] , \mem_a[12][38] , 
	\mem_a[12][37] , \mem_a[12][36] , \mem_a[12][35] , \mem_a[12][34] , 
	\mem_a[12][33] , \mem_a[12][32] , \mem_a[12][31] , \mem_a[12][30] , 
	\mem_a[12][29] , \mem_a[12][28] , \mem_a[12][27] , \mem_a[12][26] , 
	\mem_a[12][25] , \mem_a[12][24] , \mem_a[12][23] , \mem_a[12][22] , 
	\mem_a[12][21] , \mem_a[12][20] , \mem_a[12][19] , \mem_a[12][18] , 
	\mem_a[12][17] , \mem_a[12][16] , \mem_a[12][15] , \mem_a[12][14] , 
	\mem_a[12][13] , \mem_a[12][12] , \mem_a[12][11] , \mem_a[12][10] , 
	\mem_a[12][9] , \mem_a[12][8] , \mem_a[12][7] , \mem_a[12][6] , 
	\mem_a[12][5] , \mem_a[12][4] , \mem_a[12][3] , \mem_a[12][2] , 
	\mem_a[12][1] , \mem_a[12][0] , \mem_a[13][63] , \mem_a[13][62] , 
	\mem_a[13][61] , \mem_a[13][60] , \mem_a[13][59] , \mem_a[13][58] , 
	\mem_a[13][57] , \mem_a[13][56] , \mem_a[13][55] , \mem_a[13][54] , 
	\mem_a[13][53] , \mem_a[13][52] , \mem_a[13][51] , \mem_a[13][50] , 
	\mem_a[13][49] , \mem_a[13][48] , \mem_a[13][47] , \mem_a[13][46] , 
	\mem_a[13][45] , \mem_a[13][44] , \mem_a[13][43] , \mem_a[13][42] , 
	\mem_a[13][41] , \mem_a[13][40] , \mem_a[13][39] , \mem_a[13][38] , 
	\mem_a[13][37] , \mem_a[13][36] , \mem_a[13][35] , \mem_a[13][34] , 
	\mem_a[13][33] , \mem_a[13][32] , \mem_a[13][31] , \mem_a[13][30] , 
	\mem_a[13][29] , \mem_a[13][28] , \mem_a[13][27] , \mem_a[13][26] , 
	\mem_a[13][25] , \mem_a[13][24] , \mem_a[13][23] , \mem_a[13][22] , 
	\mem_a[13][21] , \mem_a[13][20] , \mem_a[13][19] , \mem_a[13][18] , 
	\mem_a[13][17] , \mem_a[13][16] , \mem_a[13][15] , \mem_a[13][14] , 
	\mem_a[13][13] , \mem_a[13][12] , \mem_a[13][11] , \mem_a[13][10] , 
	\mem_a[13][9] , \mem_a[13][8] , \mem_a[13][7] , \mem_a[13][6] , 
	\mem_a[13][5] , \mem_a[13][4] , \mem_a[13][3] , \mem_a[13][2] , 
	\mem_a[13][1] , \mem_a[13][0] , \mem_a[14][63] , \mem_a[14][62] , 
	\mem_a[14][61] , \mem_a[14][60] , \mem_a[14][59] , \mem_a[14][58] , 
	\mem_a[14][57] , \mem_a[14][56] , \mem_a[14][55] , \mem_a[14][54] , 
	\mem_a[14][53] , \mem_a[14][52] , \mem_a[14][51] , \mem_a[14][50] , 
	\mem_a[14][49] , \mem_a[14][48] , \mem_a[14][47] , \mem_a[14][46] , 
	\mem_a[14][45] , \mem_a[14][44] , \mem_a[14][43] , \mem_a[14][42] , 
	\mem_a[14][41] , \mem_a[14][40] , \mem_a[14][39] , \mem_a[14][38] , 
	\mem_a[14][37] , \mem_a[14][36] , \mem_a[14][35] , \mem_a[14][34] , 
	\mem_a[14][33] , \mem_a[14][32] , \mem_a[14][31] , \mem_a[14][30] , 
	\mem_a[14][29] , \mem_a[14][28] , \mem_a[14][27] , \mem_a[14][26] , 
	\mem_a[14][25] , \mem_a[14][24] , \mem_a[14][23] , \mem_a[14][22] , 
	\mem_a[14][21] , \mem_a[14][20] , \mem_a[14][19] , \mem_a[14][18] , 
	\mem_a[14][17] , \mem_a[14][16] , \mem_a[14][15] , \mem_a[14][14] , 
	\mem_a[14][13] , \mem_a[14][12] , \mem_a[14][11] , \mem_a[14][10] , 
	\mem_a[14][9] , \mem_a[14][8] , \mem_a[14][7] , \mem_a[14][6] , 
	\mem_a[14][5] , \mem_a[14][4] , \mem_a[14][3] , \mem_a[14][2] , 
	\mem_a[14][1] , \mem_a[14][0] , \mem_a[15][63] , \mem_a[15][62] , 
	\mem_a[15][61] , \mem_a[15][60] , \mem_a[15][59] , \mem_a[15][58] , 
	\mem_a[15][57] , \mem_a[15][56] , \mem_a[15][55] , \mem_a[15][54] , 
	\mem_a[15][53] , \mem_a[15][52] , \mem_a[15][51] , \mem_a[15][50] , 
	\mem_a[15][49] , \mem_a[15][48] , \mem_a[15][47] , \mem_a[15][46] , 
	\mem_a[15][45] , \mem_a[15][44] , \mem_a[15][43] , \mem_a[15][42] , 
	\mem_a[15][41] , \mem_a[15][40] , \mem_a[15][39] , \mem_a[15][38] , 
	\mem_a[15][37] , \mem_a[15][36] , \mem_a[15][35] , \mem_a[15][34] , 
	\mem_a[15][33] , \mem_a[15][32] , \mem_a[15][31] , \mem_a[15][30] , 
	\mem_a[15][29] , \mem_a[15][28] , \mem_a[15][27] , \mem_a[15][26] , 
	\mem_a[15][25] , \mem_a[15][24] , \mem_a[15][23] , \mem_a[15][22] , 
	\mem_a[15][21] , \mem_a[15][20] , \mem_a[15][19] , \mem_a[15][18] , 
	\mem_a[15][17] , \mem_a[15][16] , \mem_a[15][15] , \mem_a[15][14] , 
	\mem_a[15][13] , \mem_a[15][12] , \mem_a[15][11] , \mem_a[15][10] , 
	\mem_a[15][9] , \mem_a[15][8] , \mem_a[15][7] , \mem_a[15][6] , 
	\mem_a[15][5] , \mem_a[15][4] , \mem_a[15][3] , \mem_a[15][2] , 
	\mem_a[15][1] , \mem_a[15][0] , \mem_a[16][63] , \mem_a[16][62] , 
	\mem_a[16][61] , \mem_a[16][60] , \mem_a[16][59] , \mem_a[16][58] , 
	\mem_a[16][57] , \mem_a[16][56] , \mem_a[16][55] , \mem_a[16][54] , 
	\mem_a[16][53] , \mem_a[16][52] , \mem_a[16][51] , \mem_a[16][50] , 
	\mem_a[16][49] , \mem_a[16][48] , \mem_a[16][47] , \mem_a[16][46] , 
	\mem_a[16][45] , \mem_a[16][44] , \mem_a[16][43] , \mem_a[16][42] , 
	\mem_a[16][41] , \mem_a[16][40] , \mem_a[16][39] , \mem_a[16][38] , 
	\mem_a[16][37] , \mem_a[16][36] , \mem_a[16][35] , \mem_a[16][34] , 
	\mem_a[16][33] , \mem_a[16][32] , \mem_a[16][31] , \mem_a[16][30] , 
	\mem_a[16][29] , \mem_a[16][28] , \mem_a[16][27] , \mem_a[16][26] , 
	\mem_a[16][25] , \mem_a[16][24] , \mem_a[16][23] , \mem_a[16][22] , 
	\mem_a[16][21] , \mem_a[16][20] , \mem_a[16][19] , \mem_a[16][18] , 
	\mem_a[16][17] , \mem_a[16][16] , \mem_a[16][15] , \mem_a[16][14] , 
	\mem_a[16][13] , \mem_a[16][12] , \mem_a[16][11] , \mem_a[16][10] , 
	\mem_a[16][9] , \mem_a[16][8] , \mem_a[16][7] , \mem_a[16][6] , 
	\mem_a[16][5] , \mem_a[16][4] , \mem_a[16][3] , \mem_a[16][2] , 
	\mem_a[16][1] , \mem_a[16][0] , \mem_a[17][63] , \mem_a[17][62] , 
	\mem_a[17][61] , \mem_a[17][60] , \mem_a[17][59] , \mem_a[17][58] , 
	\mem_a[17][57] , \mem_a[17][56] , \mem_a[17][55] , \mem_a[17][54] , 
	\mem_a[17][53] , \mem_a[17][52] , \mem_a[17][51] , \mem_a[17][50] , 
	\mem_a[17][49] , \mem_a[17][48] , \mem_a[17][47] , \mem_a[17][46] , 
	\mem_a[17][45] , \mem_a[17][44] , \mem_a[17][43] , \mem_a[17][42] , 
	\mem_a[17][41] , \mem_a[17][40] , \mem_a[17][39] , \mem_a[17][38] , 
	\mem_a[17][37] , \mem_a[17][36] , \mem_a[17][35] , \mem_a[17][34] , 
	\mem_a[17][33] , \mem_a[17][32] , \mem_a[17][31] , \mem_a[17][30] , 
	\mem_a[17][29] , \mem_a[17][28] , \mem_a[17][27] , \mem_a[17][26] , 
	\mem_a[17][25] , \mem_a[17][24] , \mem_a[17][23] , \mem_a[17][22] , 
	\mem_a[17][21] , \mem_a[17][20] , \mem_a[17][19] , \mem_a[17][18] , 
	\mem_a[17][17] , \mem_a[17][16] , \mem_a[17][15] , \mem_a[17][14] , 
	\mem_a[17][13] , \mem_a[17][12] , \mem_a[17][11] , \mem_a[17][10] , 
	\mem_a[17][9] , \mem_a[17][8] , \mem_a[17][7] , \mem_a[17][6] , 
	\mem_a[17][5] , \mem_a[17][4] , \mem_a[17][3] , \mem_a[17][2] , 
	\mem_a[17][1] , \mem_a[17][0] , \mem_a[18][63] , \mem_a[18][62] , 
	\mem_a[18][61] , \mem_a[18][60] , \mem_a[18][59] , \mem_a[18][58] , 
	\mem_a[18][57] , \mem_a[18][56] , \mem_a[18][55] , \mem_a[18][54] , 
	\mem_a[18][53] , \mem_a[18][52] , \mem_a[18][51] , \mem_a[18][50] , 
	\mem_a[18][49] , \mem_a[18][48] , \mem_a[18][47] , \mem_a[18][46] , 
	\mem_a[18][45] , \mem_a[18][44] , \mem_a[18][43] , \mem_a[18][42] , 
	\mem_a[18][41] , \mem_a[18][40] , \mem_a[18][39] , \mem_a[18][38] , 
	\mem_a[18][37] , \mem_a[18][36] , \mem_a[18][35] , \mem_a[18][34] , 
	\mem_a[18][33] , \mem_a[18][32] , \mem_a[18][31] , \mem_a[18][30] , 
	\mem_a[18][29] , \mem_a[18][28] , \mem_a[18][27] , \mem_a[18][26] , 
	\mem_a[18][25] , \mem_a[18][24] , \mem_a[18][23] , \mem_a[18][22] , 
	\mem_a[18][21] , \mem_a[18][20] , \mem_a[18][19] , \mem_a[18][18] , 
	\mem_a[18][17] , \mem_a[18][16] , \mem_a[18][15] , \mem_a[18][14] , 
	\mem_a[18][13] , \mem_a[18][12] , \mem_a[18][11] , \mem_a[18][10] , 
	\mem_a[18][9] , \mem_a[18][8] , \mem_a[18][7] , \mem_a[18][6] , 
	\mem_a[18][5] , \mem_a[18][4] , \mem_a[18][3] , \mem_a[18][2] , 
	\mem_a[18][1] , \mem_a[18][0] , \mem_a[19][63] , \mem_a[19][62] , 
	\mem_a[19][61] , \mem_a[19][60] , \mem_a[19][59] , \mem_a[19][58] , 
	\mem_a[19][57] , \mem_a[19][56] , \mem_a[19][55] , \mem_a[19][54] , 
	\mem_a[19][53] , \mem_a[19][52] , \mem_a[19][51] , \mem_a[19][50] , 
	\mem_a[19][49] , \mem_a[19][48] , \mem_a[19][47] , \mem_a[19][46] , 
	\mem_a[19][45] , \mem_a[19][44] , \mem_a[19][43] , \mem_a[19][42] , 
	\mem_a[19][41] , \mem_a[19][40] , \mem_a[19][39] , \mem_a[19][38] , 
	\mem_a[19][37] , \mem_a[19][36] , \mem_a[19][35] , \mem_a[19][34] , 
	\mem_a[19][33] , \mem_a[19][32] , \mem_a[19][31] , \mem_a[19][30] , 
	\mem_a[19][29] , \mem_a[19][28] , \mem_a[19][27] , \mem_a[19][26] , 
	\mem_a[19][25] , \mem_a[19][24] , \mem_a[19][23] , \mem_a[19][22] , 
	\mem_a[19][21] , \mem_a[19][20] , \mem_a[19][19] , \mem_a[19][18] , 
	\mem_a[19][17] , \mem_a[19][16] , \mem_a[19][15] , \mem_a[19][14] , 
	\mem_a[19][13] , \mem_a[19][12] , \mem_a[19][11] , \mem_a[19][10] , 
	\mem_a[19][9] , \mem_a[19][8] , \mem_a[19][7] , \mem_a[19][6] , 
	\mem_a[19][5] , \mem_a[19][4] , \mem_a[19][3] , \mem_a[19][2] , 
	\mem_a[19][1] , \mem_a[19][0] , \mem_a[20][63] , \mem_a[20][62] , 
	\mem_a[20][61] , \mem_a[20][60] , \mem_a[20][59] , \mem_a[20][58] , 
	\mem_a[20][57] , \mem_a[20][56] , \mem_a[20][55] , \mem_a[20][54] , 
	\mem_a[20][53] , \mem_a[20][52] , \mem_a[20][51] , \mem_a[20][50] , 
	\mem_a[20][49] , \mem_a[20][48] , \mem_a[20][47] , \mem_a[20][46] , 
	\mem_a[20][45] , \mem_a[20][44] , \mem_a[20][43] , \mem_a[20][42] , 
	\mem_a[20][41] , \mem_a[20][40] , \mem_a[20][39] , \mem_a[20][38] , 
	\mem_a[20][37] , \mem_a[20][36] , \mem_a[20][35] , \mem_a[20][34] , 
	\mem_a[20][33] , \mem_a[20][32] , \mem_a[20][31] , \mem_a[20][30] , 
	\mem_a[20][29] , \mem_a[20][28] , \mem_a[20][27] , \mem_a[20][26] , 
	\mem_a[20][25] , \mem_a[20][24] , \mem_a[20][23] , \mem_a[20][22] , 
	\mem_a[20][21] , \mem_a[20][20] , \mem_a[20][19] , \mem_a[20][18] , 
	\mem_a[20][17] , \mem_a[20][16] , \mem_a[20][15] , \mem_a[20][14] , 
	\mem_a[20][13] , \mem_a[20][12] , \mem_a[20][11] , \mem_a[20][10] , 
	\mem_a[20][9] , \mem_a[20][8] , \mem_a[20][7] , \mem_a[20][6] , 
	\mem_a[20][5] , \mem_a[20][4] , \mem_a[20][3] , \mem_a[20][2] , 
	\mem_a[20][1] , \mem_a[20][0] , \mem_a[21][63] , \mem_a[21][62] , 
	\mem_a[21][61] , \mem_a[21][60] , \mem_a[21][59] , \mem_a[21][58] , 
	\mem_a[21][57] , \mem_a[21][56] , \mem_a[21][55] , \mem_a[21][54] , 
	\mem_a[21][53] , \mem_a[21][52] , \mem_a[21][51] , \mem_a[21][50] , 
	\mem_a[21][49] , \mem_a[21][48] , \mem_a[21][47] , \mem_a[21][46] , 
	\mem_a[21][45] , \mem_a[21][44] , \mem_a[21][43] , \mem_a[21][42] , 
	\mem_a[21][41] , \mem_a[21][40] , \mem_a[21][39] , \mem_a[21][38] , 
	\mem_a[21][37] , \mem_a[21][36] , \mem_a[21][35] , \mem_a[21][34] , 
	\mem_a[21][33] , \mem_a[21][32] , \mem_a[21][31] , \mem_a[21][30] , 
	\mem_a[21][29] , \mem_a[21][28] , \mem_a[21][27] , \mem_a[21][26] , 
	\mem_a[21][25] , \mem_a[21][24] , \mem_a[21][23] , \mem_a[21][22] , 
	\mem_a[21][21] , \mem_a[21][20] , \mem_a[21][19] , \mem_a[21][18] , 
	\mem_a[21][17] , \mem_a[21][16] , \mem_a[21][15] , \mem_a[21][14] , 
	\mem_a[21][13] , \mem_a[21][12] , \mem_a[21][11] , \mem_a[21][10] , 
	\mem_a[21][9] , \mem_a[21][8] , \mem_a[21][7] , \mem_a[21][6] , 
	\mem_a[21][5] , \mem_a[21][4] , \mem_a[21][3] , \mem_a[21][2] , 
	\mem_a[21][1] , \mem_a[21][0] , \mem_a[22][63] , \mem_a[22][62] , 
	\mem_a[22][61] , \mem_a[22][60] , \mem_a[22][59] , \mem_a[22][58] , 
	\mem_a[22][57] , \mem_a[22][56] , \mem_a[22][55] , \mem_a[22][54] , 
	\mem_a[22][53] , \mem_a[22][52] , \mem_a[22][51] , \mem_a[22][50] , 
	\mem_a[22][49] , \mem_a[22][48] , \mem_a[22][47] , \mem_a[22][46] , 
	\mem_a[22][45] , \mem_a[22][44] , \mem_a[22][43] , \mem_a[22][42] , 
	\mem_a[22][41] , \mem_a[22][40] , \mem_a[22][39] , \mem_a[22][38] , 
	\mem_a[22][37] , \mem_a[22][36] , \mem_a[22][35] , \mem_a[22][34] , 
	\mem_a[22][33] , \mem_a[22][32] , \mem_a[22][31] , \mem_a[22][30] , 
	\mem_a[22][29] , \mem_a[22][28] , \mem_a[22][27] , \mem_a[22][26] , 
	\mem_a[22][25] , \mem_a[22][24] , \mem_a[22][23] , \mem_a[22][22] , 
	\mem_a[22][21] , \mem_a[22][20] , \mem_a[22][19] , \mem_a[22][18] , 
	\mem_a[22][17] , \mem_a[22][16] , \mem_a[22][15] , \mem_a[22][14] , 
	\mem_a[22][13] , \mem_a[22][12] , \mem_a[22][11] , \mem_a[22][10] , 
	\mem_a[22][9] , \mem_a[22][8] , \mem_a[22][7] , \mem_a[22][6] , 
	\mem_a[22][5] , \mem_a[22][4] , \mem_a[22][3] , \mem_a[22][2] , 
	\mem_a[22][1] , \mem_a[22][0] , \mem_a[23][63] , \mem_a[23][62] , 
	\mem_a[23][61] , \mem_a[23][60] , \mem_a[23][59] , \mem_a[23][58] , 
	\mem_a[23][57] , \mem_a[23][56] , \mem_a[23][55] , \mem_a[23][54] , 
	\mem_a[23][53] , \mem_a[23][52] , \mem_a[23][51] , \mem_a[23][50] , 
	\mem_a[23][49] , \mem_a[23][48] , \mem_a[23][47] , \mem_a[23][46] , 
	\mem_a[23][45] , \mem_a[23][44] , \mem_a[23][43] , \mem_a[23][42] , 
	\mem_a[23][41] , \mem_a[23][40] , \mem_a[23][39] , \mem_a[23][38] , 
	\mem_a[23][37] , \mem_a[23][36] , \mem_a[23][35] , \mem_a[23][34] , 
	\mem_a[23][33] , \mem_a[23][32] , \mem_a[23][31] , \mem_a[23][30] , 
	\mem_a[23][29] , \mem_a[23][28] , \mem_a[23][27] , \mem_a[23][26] , 
	\mem_a[23][25] , \mem_a[23][24] , \mem_a[23][23] , \mem_a[23][22] , 
	\mem_a[23][21] , \mem_a[23][20] , \mem_a[23][19] , \mem_a[23][18] , 
	\mem_a[23][17] , \mem_a[23][16] , \mem_a[23][15] , \mem_a[23][14] , 
	\mem_a[23][13] , \mem_a[23][12] , \mem_a[23][11] , \mem_a[23][10] , 
	\mem_a[23][9] , \mem_a[23][8] , \mem_a[23][7] , \mem_a[23][6] , 
	\mem_a[23][5] , \mem_a[23][4] , \mem_a[23][3] , \mem_a[23][2] , 
	\mem_a[23][1] , \mem_a[23][0] , \mem_a[24][63] , \mem_a[24][62] , 
	\mem_a[24][61] , \mem_a[24][60] , \mem_a[24][59] , \mem_a[24][58] , 
	\mem_a[24][57] , \mem_a[24][56] , \mem_a[24][55] , \mem_a[24][54] , 
	\mem_a[24][53] , \mem_a[24][52] , \mem_a[24][51] , \mem_a[24][50] , 
	\mem_a[24][49] , \mem_a[24][48] , \mem_a[24][47] , \mem_a[24][46] , 
	\mem_a[24][45] , \mem_a[24][44] , \mem_a[24][43] , \mem_a[24][42] , 
	\mem_a[24][41] , \mem_a[24][40] , \mem_a[24][39] , \mem_a[24][38] , 
	\mem_a[24][37] , \mem_a[24][36] , \mem_a[24][35] , \mem_a[24][34] , 
	\mem_a[24][33] , \mem_a[24][32] , \mem_a[24][31] , \mem_a[24][30] , 
	\mem_a[24][29] , \mem_a[24][28] , \mem_a[24][27] , \mem_a[24][26] , 
	\mem_a[24][25] , \mem_a[24][24] , \mem_a[24][23] , \mem_a[24][22] , 
	\mem_a[24][21] , \mem_a[24][20] , \mem_a[24][19] , \mem_a[24][18] , 
	\mem_a[24][17] , \mem_a[24][16] , \mem_a[24][15] , \mem_a[24][14] , 
	\mem_a[24][13] , \mem_a[24][12] , \mem_a[24][11] , \mem_a[24][10] , 
	\mem_a[24][9] , \mem_a[24][8] , \mem_a[24][7] , \mem_a[24][6] , 
	\mem_a[24][5] , \mem_a[24][4] , \mem_a[24][3] , \mem_a[24][2] , 
	\mem_a[24][1] , \mem_a[24][0] , \mem_a[25][63] , \mem_a[25][62] , 
	\mem_a[25][61] , \mem_a[25][60] , \mem_a[25][59] , \mem_a[25][58] , 
	\mem_a[25][57] , \mem_a[25][56] , \mem_a[25][55] , \mem_a[25][54] , 
	\mem_a[25][53] , \mem_a[25][52] , \mem_a[25][51] , \mem_a[25][50] , 
	\mem_a[25][49] , \mem_a[25][48] , \mem_a[25][47] , \mem_a[25][46] , 
	\mem_a[25][45] , \mem_a[25][44] , \mem_a[25][43] , \mem_a[25][42] , 
	\mem_a[25][41] , \mem_a[25][40] , \mem_a[25][39] , \mem_a[25][38] , 
	\mem_a[25][37] , \mem_a[25][36] , \mem_a[25][35] , \mem_a[25][34] , 
	\mem_a[25][33] , \mem_a[25][32] , \mem_a[25][31] , \mem_a[25][30] , 
	\mem_a[25][29] , \mem_a[25][28] , \mem_a[25][27] , \mem_a[25][26] , 
	\mem_a[25][25] , \mem_a[25][24] , \mem_a[25][23] , \mem_a[25][22] , 
	\mem_a[25][21] , \mem_a[25][20] , \mem_a[25][19] , \mem_a[25][18] , 
	\mem_a[25][17] , \mem_a[25][16] , \mem_a[25][15] , \mem_a[25][14] , 
	\mem_a[25][13] , \mem_a[25][12] , \mem_a[25][11] , \mem_a[25][10] , 
	\mem_a[25][9] , \mem_a[25][8] , \mem_a[25][7] , \mem_a[25][6] , 
	\mem_a[25][5] , \mem_a[25][4] , \mem_a[25][3] , \mem_a[25][2] , 
	\mem_a[25][1] , \mem_a[25][0] , \mem_a[26][63] , \mem_a[26][62] , 
	\mem_a[26][61] , \mem_a[26][60] , \mem_a[26][59] , \mem_a[26][58] , 
	\mem_a[26][57] , \mem_a[26][56] , \mem_a[26][55] , \mem_a[26][54] , 
	\mem_a[26][53] , \mem_a[26][52] , \mem_a[26][51] , \mem_a[26][50] , 
	\mem_a[26][49] , \mem_a[26][48] , \mem_a[26][47] , \mem_a[26][46] , 
	\mem_a[26][45] , \mem_a[26][44] , \mem_a[26][43] , \mem_a[26][42] , 
	\mem_a[26][41] , \mem_a[26][40] , \mem_a[26][39] , \mem_a[26][38] , 
	\mem_a[26][37] , \mem_a[26][36] , \mem_a[26][35] , \mem_a[26][34] , 
	\mem_a[26][33] , \mem_a[26][32] , \mem_a[26][31] , \mem_a[26][30] , 
	\mem_a[26][29] , \mem_a[26][28] , \mem_a[26][27] , \mem_a[26][26] , 
	\mem_a[26][25] , \mem_a[26][24] , \mem_a[26][23] , \mem_a[26][22] , 
	\mem_a[26][21] , \mem_a[26][20] , \mem_a[26][19] , \mem_a[26][18] , 
	\mem_a[26][17] , \mem_a[26][16] , \mem_a[26][15] , \mem_a[26][14] , 
	\mem_a[26][13] , \mem_a[26][12] , \mem_a[26][11] , \mem_a[26][10] , 
	\mem_a[26][9] , \mem_a[26][8] , \mem_a[26][7] , \mem_a[26][6] , 
	\mem_a[26][5] , \mem_a[26][4] , \mem_a[26][3] , \mem_a[26][2] , 
	\mem_a[26][1] , \mem_a[26][0] , \mem_a[27][63] , \mem_a[27][62] , 
	\mem_a[27][61] , \mem_a[27][60] , \mem_a[27][59] , \mem_a[27][58] , 
	\mem_a[27][57] , \mem_a[27][56] , \mem_a[27][55] , \mem_a[27][54] , 
	\mem_a[27][53] , \mem_a[27][52] , \mem_a[27][51] , \mem_a[27][50] , 
	\mem_a[27][49] , \mem_a[27][48] , \mem_a[27][47] , \mem_a[27][46] , 
	\mem_a[27][45] , \mem_a[27][44] , \mem_a[27][43] , \mem_a[27][42] , 
	\mem_a[27][41] , \mem_a[27][40] , \mem_a[27][39] , \mem_a[27][38] , 
	\mem_a[27][37] , \mem_a[27][36] , \mem_a[27][35] , \mem_a[27][34] , 
	\mem_a[27][33] , \mem_a[27][32] , \mem_a[27][31] , \mem_a[27][30] , 
	\mem_a[27][29] , \mem_a[27][28] , \mem_a[27][27] , \mem_a[27][26] , 
	\mem_a[27][25] , \mem_a[27][24] , \mem_a[27][23] , \mem_a[27][22] , 
	\mem_a[27][21] , \mem_a[27][20] , \mem_a[27][19] , \mem_a[27][18] , 
	\mem_a[27][17] , \mem_a[27][16] , \mem_a[27][15] , \mem_a[27][14] , 
	\mem_a[27][13] , \mem_a[27][12] , \mem_a[27][11] , \mem_a[27][10] , 
	\mem_a[27][9] , \mem_a[27][8] , \mem_a[27][7] , \mem_a[27][6] , 
	\mem_a[27][5] , \mem_a[27][4] , \mem_a[27][3] , \mem_a[27][2] , 
	\mem_a[27][1] , \mem_a[27][0] , \mem_a[28][63] , \mem_a[28][62] , 
	\mem_a[28][61] , \mem_a[28][60] , \mem_a[28][59] , \mem_a[28][58] , 
	\mem_a[28][57] , \mem_a[28][56] , \mem_a[28][55] , \mem_a[28][54] , 
	\mem_a[28][53] , \mem_a[28][52] , \mem_a[28][51] , \mem_a[28][50] , 
	\mem_a[28][49] , \mem_a[28][48] , \mem_a[28][47] , \mem_a[28][46] , 
	\mem_a[28][45] , \mem_a[28][44] , \mem_a[28][43] , \mem_a[28][42] , 
	\mem_a[28][41] , \mem_a[28][40] , \mem_a[28][39] , \mem_a[28][38] , 
	\mem_a[28][37] , \mem_a[28][36] , \mem_a[28][35] , \mem_a[28][34] , 
	\mem_a[28][33] , \mem_a[28][32] , \mem_a[28][31] , \mem_a[28][30] , 
	\mem_a[28][29] , \mem_a[28][28] , \mem_a[28][27] , \mem_a[28][26] , 
	\mem_a[28][25] , \mem_a[28][24] , \mem_a[28][23] , \mem_a[28][22] , 
	\mem_a[28][21] , \mem_a[28][20] , \mem_a[28][19] , \mem_a[28][18] , 
	\mem_a[28][17] , \mem_a[28][16] , \mem_a[28][15] , \mem_a[28][14] , 
	\mem_a[28][13] , \mem_a[28][12] , \mem_a[28][11] , \mem_a[28][10] , 
	\mem_a[28][9] , \mem_a[28][8] , \mem_a[28][7] , \mem_a[28][6] , 
	\mem_a[28][5] , \mem_a[28][4] , \mem_a[28][3] , \mem_a[28][2] , 
	\mem_a[28][1] , \mem_a[28][0] , \mem_a[29][63] , \mem_a[29][62] , 
	\mem_a[29][61] , \mem_a[29][60] , \mem_a[29][59] , \mem_a[29][58] , 
	\mem_a[29][57] , \mem_a[29][56] , \mem_a[29][55] , \mem_a[29][54] , 
	\mem_a[29][53] , \mem_a[29][52] , \mem_a[29][51] , \mem_a[29][50] , 
	\mem_a[29][49] , \mem_a[29][48] , \mem_a[29][47] , \mem_a[29][46] , 
	\mem_a[29][45] , \mem_a[29][44] , \mem_a[29][43] , \mem_a[29][42] , 
	\mem_a[29][41] , \mem_a[29][40] , \mem_a[29][39] , \mem_a[29][38] , 
	\mem_a[29][37] , \mem_a[29][36] , \mem_a[29][35] , \mem_a[29][34] , 
	\mem_a[29][33] , \mem_a[29][32] , \mem_a[29][31] , \mem_a[29][30] , 
	\mem_a[29][29] , \mem_a[29][28] , \mem_a[29][27] , \mem_a[29][26] , 
	\mem_a[29][25] , \mem_a[29][24] , \mem_a[29][23] , \mem_a[29][22] , 
	\mem_a[29][21] , \mem_a[29][20] , \mem_a[29][19] , \mem_a[29][18] , 
	\mem_a[29][17] , \mem_a[29][16] , \mem_a[29][15] , \mem_a[29][14] , 
	\mem_a[29][13] , \mem_a[29][12] , \mem_a[29][11] , \mem_a[29][10] , 
	\mem_a[29][9] , \mem_a[29][8] , \mem_a[29][7] , \mem_a[29][6] , 
	\mem_a[29][5] , \mem_a[29][4] , \mem_a[29][3] , \mem_a[29][2] , 
	\mem_a[29][1] , \mem_a[29][0] , \mem_a[30][63] , \mem_a[30][62] , 
	\mem_a[30][61] , \mem_a[30][60] , \mem_a[30][59] , \mem_a[30][58] , 
	\mem_a[30][57] , \mem_a[30][56] , \mem_a[30][55] , \mem_a[30][54] , 
	\mem_a[30][53] , \mem_a[30][52] , \mem_a[30][51] , \mem_a[30][50] , 
	\mem_a[30][49] , \mem_a[30][48] , \mem_a[30][47] , \mem_a[30][46] , 
	\mem_a[30][45] , \mem_a[30][44] , \mem_a[30][43] , \mem_a[30][42] , 
	\mem_a[30][41] , \mem_a[30][40] , \mem_a[30][39] , \mem_a[30][38] , 
	\mem_a[30][37] , \mem_a[30][36] , \mem_a[30][35] , \mem_a[30][34] , 
	\mem_a[30][33] , \mem_a[30][32] , \mem_a[30][31] , \mem_a[30][30] , 
	\mem_a[30][29] , \mem_a[30][28] , \mem_a[30][27] , \mem_a[30][26] , 
	\mem_a[30][25] , \mem_a[30][24] , \mem_a[30][23] , \mem_a[30][22] , 
	\mem_a[30][21] , \mem_a[30][20] , \mem_a[30][19] , \mem_a[30][18] , 
	\mem_a[30][17] , \mem_a[30][16] , \mem_a[30][15] , \mem_a[30][14] , 
	\mem_a[30][13] , \mem_a[30][12] , \mem_a[30][11] , \mem_a[30][10] , 
	\mem_a[30][9] , \mem_a[30][8] , \mem_a[30][7] , \mem_a[30][6] , 
	\mem_a[30][5] , \mem_a[30][4] , \mem_a[30][3] , \mem_a[30][2] , 
	\mem_a[30][1] , \mem_a[30][0] , \mem_a[31][63] , \mem_a[31][62] , 
	\mem_a[31][61] , \mem_a[31][60] , \mem_a[31][59] , \mem_a[31][58] , 
	\mem_a[31][57] , \mem_a[31][56] , \mem_a[31][55] , \mem_a[31][54] , 
	\mem_a[31][53] , \mem_a[31][52] , \mem_a[31][51] , \mem_a[31][50] , 
	\mem_a[31][49] , \mem_a[31][48] , \mem_a[31][47] , \mem_a[31][46] , 
	\mem_a[31][45] , \mem_a[31][44] , \mem_a[31][43] , \mem_a[31][42] , 
	\mem_a[31][41] , \mem_a[31][40] , \mem_a[31][39] , \mem_a[31][38] , 
	\mem_a[31][37] , \mem_a[31][36] , \mem_a[31][35] , \mem_a[31][34] , 
	\mem_a[31][33] , \mem_a[31][32] , \mem_a[31][31] , \mem_a[31][30] , 
	\mem_a[31][29] , \mem_a[31][28] , \mem_a[31][27] , \mem_a[31][26] , 
	\mem_a[31][25] , \mem_a[31][24] , \mem_a[31][23] , \mem_a[31][22] , 
	\mem_a[31][21] , \mem_a[31][20] , \mem_a[31][19] , \mem_a[31][18] , 
	\mem_a[31][17] , \mem_a[31][16] , \mem_a[31][15] , \mem_a[31][14] , 
	\mem_a[31][13] , \mem_a[31][12] , \mem_a[31][11] , \mem_a[31][10] , 
	\mem_a[31][9] , \mem_a[31][8] , \mem_a[31][7] , \mem_a[31][6] , 
	\mem_a[31][5] , \mem_a[31][4] , \mem_a[31][3] , \mem_a[31][2] , 
	\mem_a[31][1] , \mem_a[31][0] } ));
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output [2:0] stat_code;
output [4:0] stat_datawords;
output [4:0] stat_addr;
output [15:0] capability_lst;
output [3:0] capability_type;
output [63:0] rd_dat;
input clk;
input rst_n;
input [10:0] addr;
input [3:0] cmnd_op;
input [4:0] cmnd_addr;
input wr_stb;
input [63:0] wr_dat;
input \mem_a[0][63] ;
input \mem_a[0][62] ;
input \mem_a[0][61] ;
input \mem_a[0][60] ;
input \mem_a[0][59] ;
input \mem_a[0][58] ;
input \mem_a[0][57] ;
input \mem_a[0][56] ;
input \mem_a[0][55] ;
input \mem_a[0][54] ;
input \mem_a[0][53] ;
input \mem_a[0][52] ;
input \mem_a[0][51] ;
input \mem_a[0][50] ;
input \mem_a[0][49] ;
input \mem_a[0][48] ;
input \mem_a[0][47] ;
input \mem_a[0][46] ;
input \mem_a[0][45] ;
input \mem_a[0][44] ;
input \mem_a[0][43] ;
input \mem_a[0][42] ;
input \mem_a[0][41] ;
input \mem_a[0][40] ;
input \mem_a[0][39] ;
input \mem_a[0][38] ;
input \mem_a[0][37] ;
input \mem_a[0][36] ;
input \mem_a[0][35] ;
input \mem_a[0][34] ;
input \mem_a[0][33] ;
input \mem_a[0][32] ;
input \mem_a[0][31] ;
input \mem_a[0][30] ;
input \mem_a[0][29] ;
input \mem_a[0][28] ;
input \mem_a[0][27] ;
input \mem_a[0][26] ;
input \mem_a[0][25] ;
input \mem_a[0][24] ;
input \mem_a[0][23] ;
input \mem_a[0][22] ;
input \mem_a[0][21] ;
input \mem_a[0][20] ;
input \mem_a[0][19] ;
input \mem_a[0][18] ;
input \mem_a[0][17] ;
input \mem_a[0][16] ;
input \mem_a[0][15] ;
input \mem_a[0][14] ;
input \mem_a[0][13] ;
input \mem_a[0][12] ;
input \mem_a[0][11] ;
input \mem_a[0][10] ;
input \mem_a[0][9] ;
input \mem_a[0][8] ;
input \mem_a[0][7] ;
input \mem_a[0][6] ;
input \mem_a[0][5] ;
input \mem_a[0][4] ;
input \mem_a[0][3] ;
input \mem_a[0][2] ;
input \mem_a[0][1] ;
input \mem_a[0][0] ;
input \mem_a[1][63] ;
input \mem_a[1][62] ;
input \mem_a[1][61] ;
input \mem_a[1][60] ;
input \mem_a[1][59] ;
input \mem_a[1][58] ;
input \mem_a[1][57] ;
input \mem_a[1][56] ;
input \mem_a[1][55] ;
input \mem_a[1][54] ;
input \mem_a[1][53] ;
input \mem_a[1][52] ;
input \mem_a[1][51] ;
input \mem_a[1][50] ;
input \mem_a[1][49] ;
input \mem_a[1][48] ;
input \mem_a[1][47] ;
input \mem_a[1][46] ;
input \mem_a[1][45] ;
input \mem_a[1][44] ;
input \mem_a[1][43] ;
input \mem_a[1][42] ;
input \mem_a[1][41] ;
input \mem_a[1][40] ;
input \mem_a[1][39] ;
input \mem_a[1][38] ;
input \mem_a[1][37] ;
input \mem_a[1][36] ;
input \mem_a[1][35] ;
input \mem_a[1][34] ;
input \mem_a[1][33] ;
input \mem_a[1][32] ;
input \mem_a[1][31] ;
input \mem_a[1][30] ;
input \mem_a[1][29] ;
input \mem_a[1][28] ;
input \mem_a[1][27] ;
input \mem_a[1][26] ;
input \mem_a[1][25] ;
input \mem_a[1][24] ;
input \mem_a[1][23] ;
input \mem_a[1][22] ;
input \mem_a[1][21] ;
input \mem_a[1][20] ;
input \mem_a[1][19] ;
input \mem_a[1][18] ;
input \mem_a[1][17] ;
input \mem_a[1][16] ;
input \mem_a[1][15] ;
input \mem_a[1][14] ;
input \mem_a[1][13] ;
input \mem_a[1][12] ;
input \mem_a[1][11] ;
input \mem_a[1][10] ;
input \mem_a[1][9] ;
input \mem_a[1][8] ;
input \mem_a[1][7] ;
input \mem_a[1][6] ;
input \mem_a[1][5] ;
input \mem_a[1][4] ;
input \mem_a[1][3] ;
input \mem_a[1][2] ;
input \mem_a[1][1] ;
input \mem_a[1][0] ;
input \mem_a[2][63] ;
input \mem_a[2][62] ;
input \mem_a[2][61] ;
input \mem_a[2][60] ;
input \mem_a[2][59] ;
input \mem_a[2][58] ;
input \mem_a[2][57] ;
input \mem_a[2][56] ;
input \mem_a[2][55] ;
input \mem_a[2][54] ;
input \mem_a[2][53] ;
input \mem_a[2][52] ;
input \mem_a[2][51] ;
input \mem_a[2][50] ;
input \mem_a[2][49] ;
input \mem_a[2][48] ;
input \mem_a[2][47] ;
input \mem_a[2][46] ;
input \mem_a[2][45] ;
input \mem_a[2][44] ;
input \mem_a[2][43] ;
input \mem_a[2][42] ;
input \mem_a[2][41] ;
input \mem_a[2][40] ;
input \mem_a[2][39] ;
input \mem_a[2][38] ;
input \mem_a[2][37] ;
input \mem_a[2][36] ;
input \mem_a[2][35] ;
input \mem_a[2][34] ;
input \mem_a[2][33] ;
input \mem_a[2][32] ;
input \mem_a[2][31] ;
input \mem_a[2][30] ;
input \mem_a[2][29] ;
input \mem_a[2][28] ;
input \mem_a[2][27] ;
input \mem_a[2][26] ;
input \mem_a[2][25] ;
input \mem_a[2][24] ;
input \mem_a[2][23] ;
input \mem_a[2][22] ;
input \mem_a[2][21] ;
input \mem_a[2][20] ;
input \mem_a[2][19] ;
input \mem_a[2][18] ;
input \mem_a[2][17] ;
input \mem_a[2][16] ;
input \mem_a[2][15] ;
input \mem_a[2][14] ;
input \mem_a[2][13] ;
input \mem_a[2][12] ;
input \mem_a[2][11] ;
input \mem_a[2][10] ;
input \mem_a[2][9] ;
input \mem_a[2][8] ;
input \mem_a[2][7] ;
input \mem_a[2][6] ;
input \mem_a[2][5] ;
input \mem_a[2][4] ;
input \mem_a[2][3] ;
input \mem_a[2][2] ;
input \mem_a[2][1] ;
input \mem_a[2][0] ;
input \mem_a[3][63] ;
input \mem_a[3][62] ;
input \mem_a[3][61] ;
input \mem_a[3][60] ;
input \mem_a[3][59] ;
input \mem_a[3][58] ;
input \mem_a[3][57] ;
input \mem_a[3][56] ;
input \mem_a[3][55] ;
input \mem_a[3][54] ;
input \mem_a[3][53] ;
input \mem_a[3][52] ;
input \mem_a[3][51] ;
input \mem_a[3][50] ;
input \mem_a[3][49] ;
input \mem_a[3][48] ;
input \mem_a[3][47] ;
input \mem_a[3][46] ;
input \mem_a[3][45] ;
input \mem_a[3][44] ;
input \mem_a[3][43] ;
input \mem_a[3][42] ;
input \mem_a[3][41] ;
input \mem_a[3][40] ;
input \mem_a[3][39] ;
input \mem_a[3][38] ;
input \mem_a[3][37] ;
input \mem_a[3][36] ;
input \mem_a[3][35] ;
input \mem_a[3][34] ;
input \mem_a[3][33] ;
input \mem_a[3][32] ;
input \mem_a[3][31] ;
input \mem_a[3][30] ;
input \mem_a[3][29] ;
input \mem_a[3][28] ;
input \mem_a[3][27] ;
input \mem_a[3][26] ;
input \mem_a[3][25] ;
input \mem_a[3][24] ;
input \mem_a[3][23] ;
input \mem_a[3][22] ;
input \mem_a[3][21] ;
input \mem_a[3][20] ;
input \mem_a[3][19] ;
input \mem_a[3][18] ;
input \mem_a[3][17] ;
input \mem_a[3][16] ;
input \mem_a[3][15] ;
input \mem_a[3][14] ;
input \mem_a[3][13] ;
input \mem_a[3][12] ;
input \mem_a[3][11] ;
input \mem_a[3][10] ;
input \mem_a[3][9] ;
input \mem_a[3][8] ;
input \mem_a[3][7] ;
input \mem_a[3][6] ;
input \mem_a[3][5] ;
input \mem_a[3][4] ;
input \mem_a[3][3] ;
input \mem_a[3][2] ;
input \mem_a[3][1] ;
input \mem_a[3][0] ;
input \mem_a[4][63] ;
input \mem_a[4][62] ;
input \mem_a[4][61] ;
input \mem_a[4][60] ;
input \mem_a[4][59] ;
input \mem_a[4][58] ;
input \mem_a[4][57] ;
input \mem_a[4][56] ;
input \mem_a[4][55] ;
input \mem_a[4][54] ;
input \mem_a[4][53] ;
input \mem_a[4][52] ;
input \mem_a[4][51] ;
input \mem_a[4][50] ;
input \mem_a[4][49] ;
input \mem_a[4][48] ;
input \mem_a[4][47] ;
input \mem_a[4][46] ;
input \mem_a[4][45] ;
input \mem_a[4][44] ;
input \mem_a[4][43] ;
input \mem_a[4][42] ;
input \mem_a[4][41] ;
input \mem_a[4][40] ;
input \mem_a[4][39] ;
input \mem_a[4][38] ;
input \mem_a[4][37] ;
input \mem_a[4][36] ;
input \mem_a[4][35] ;
input \mem_a[4][34] ;
input \mem_a[4][33] ;
input \mem_a[4][32] ;
input \mem_a[4][31] ;
input \mem_a[4][30] ;
input \mem_a[4][29] ;
input \mem_a[4][28] ;
input \mem_a[4][27] ;
input \mem_a[4][26] ;
input \mem_a[4][25] ;
input \mem_a[4][24] ;
input \mem_a[4][23] ;
input \mem_a[4][22] ;
input \mem_a[4][21] ;
input \mem_a[4][20] ;
input \mem_a[4][19] ;
input \mem_a[4][18] ;
input \mem_a[4][17] ;
input \mem_a[4][16] ;
input \mem_a[4][15] ;
input \mem_a[4][14] ;
input \mem_a[4][13] ;
input \mem_a[4][12] ;
input \mem_a[4][11] ;
input \mem_a[4][10] ;
input \mem_a[4][9] ;
input \mem_a[4][8] ;
input \mem_a[4][7] ;
input \mem_a[4][6] ;
input \mem_a[4][5] ;
input \mem_a[4][4] ;
input \mem_a[4][3] ;
input \mem_a[4][2] ;
input \mem_a[4][1] ;
input \mem_a[4][0] ;
input \mem_a[5][63] ;
input \mem_a[5][62] ;
input \mem_a[5][61] ;
input \mem_a[5][60] ;
input \mem_a[5][59] ;
input \mem_a[5][58] ;
input \mem_a[5][57] ;
input \mem_a[5][56] ;
input \mem_a[5][55] ;
input \mem_a[5][54] ;
input \mem_a[5][53] ;
input \mem_a[5][52] ;
input \mem_a[5][51] ;
input \mem_a[5][50] ;
input \mem_a[5][49] ;
input \mem_a[5][48] ;
input \mem_a[5][47] ;
input \mem_a[5][46] ;
input \mem_a[5][45] ;
input \mem_a[5][44] ;
input \mem_a[5][43] ;
input \mem_a[5][42] ;
input \mem_a[5][41] ;
input \mem_a[5][40] ;
input \mem_a[5][39] ;
input \mem_a[5][38] ;
input \mem_a[5][37] ;
input \mem_a[5][36] ;
input \mem_a[5][35] ;
input \mem_a[5][34] ;
input \mem_a[5][33] ;
input \mem_a[5][32] ;
input \mem_a[5][31] ;
input \mem_a[5][30] ;
input \mem_a[5][29] ;
input \mem_a[5][28] ;
input \mem_a[5][27] ;
input \mem_a[5][26] ;
input \mem_a[5][25] ;
input \mem_a[5][24] ;
input \mem_a[5][23] ;
input \mem_a[5][22] ;
input \mem_a[5][21] ;
input \mem_a[5][20] ;
input \mem_a[5][19] ;
input \mem_a[5][18] ;
input \mem_a[5][17] ;
input \mem_a[5][16] ;
input \mem_a[5][15] ;
input \mem_a[5][14] ;
input \mem_a[5][13] ;
input \mem_a[5][12] ;
input \mem_a[5][11] ;
input \mem_a[5][10] ;
input \mem_a[5][9] ;
input \mem_a[5][8] ;
input \mem_a[5][7] ;
input \mem_a[5][6] ;
input \mem_a[5][5] ;
input \mem_a[5][4] ;
input \mem_a[5][3] ;
input \mem_a[5][2] ;
input \mem_a[5][1] ;
input \mem_a[5][0] ;
input \mem_a[6][63] ;
input \mem_a[6][62] ;
input \mem_a[6][61] ;
input \mem_a[6][60] ;
input \mem_a[6][59] ;
input \mem_a[6][58] ;
input \mem_a[6][57] ;
input \mem_a[6][56] ;
input \mem_a[6][55] ;
input \mem_a[6][54] ;
input \mem_a[6][53] ;
input \mem_a[6][52] ;
input \mem_a[6][51] ;
input \mem_a[6][50] ;
input \mem_a[6][49] ;
input \mem_a[6][48] ;
input \mem_a[6][47] ;
input \mem_a[6][46] ;
input \mem_a[6][45] ;
input \mem_a[6][44] ;
input \mem_a[6][43] ;
input \mem_a[6][42] ;
input \mem_a[6][41] ;
input \mem_a[6][40] ;
input \mem_a[6][39] ;
input \mem_a[6][38] ;
input \mem_a[6][37] ;
input \mem_a[6][36] ;
input \mem_a[6][35] ;
input \mem_a[6][34] ;
input \mem_a[6][33] ;
input \mem_a[6][32] ;
input \mem_a[6][31] ;
input \mem_a[6][30] ;
input \mem_a[6][29] ;
input \mem_a[6][28] ;
input \mem_a[6][27] ;
input \mem_a[6][26] ;
input \mem_a[6][25] ;
input \mem_a[6][24] ;
input \mem_a[6][23] ;
input \mem_a[6][22] ;
input \mem_a[6][21] ;
input \mem_a[6][20] ;
input \mem_a[6][19] ;
input \mem_a[6][18] ;
input \mem_a[6][17] ;
input \mem_a[6][16] ;
input \mem_a[6][15] ;
input \mem_a[6][14] ;
input \mem_a[6][13] ;
input \mem_a[6][12] ;
input \mem_a[6][11] ;
input \mem_a[6][10] ;
input \mem_a[6][9] ;
input \mem_a[6][8] ;
input \mem_a[6][7] ;
input \mem_a[6][6] ;
input \mem_a[6][5] ;
input \mem_a[6][4] ;
input \mem_a[6][3] ;
input \mem_a[6][2] ;
input \mem_a[6][1] ;
input \mem_a[6][0] ;
input \mem_a[7][63] ;
input \mem_a[7][62] ;
input \mem_a[7][61] ;
input \mem_a[7][60] ;
input \mem_a[7][59] ;
input \mem_a[7][58] ;
input \mem_a[7][57] ;
input \mem_a[7][56] ;
input \mem_a[7][55] ;
input \mem_a[7][54] ;
input \mem_a[7][53] ;
input \mem_a[7][52] ;
input \mem_a[7][51] ;
input \mem_a[7][50] ;
input \mem_a[7][49] ;
input \mem_a[7][48] ;
input \mem_a[7][47] ;
input \mem_a[7][46] ;
input \mem_a[7][45] ;
input \mem_a[7][44] ;
input \mem_a[7][43] ;
input \mem_a[7][42] ;
input \mem_a[7][41] ;
input \mem_a[7][40] ;
input \mem_a[7][39] ;
input \mem_a[7][38] ;
input \mem_a[7][37] ;
input \mem_a[7][36] ;
input \mem_a[7][35] ;
input \mem_a[7][34] ;
input \mem_a[7][33] ;
input \mem_a[7][32] ;
input \mem_a[7][31] ;
input \mem_a[7][30] ;
input \mem_a[7][29] ;
input \mem_a[7][28] ;
input \mem_a[7][27] ;
input \mem_a[7][26] ;
input \mem_a[7][25] ;
input \mem_a[7][24] ;
input \mem_a[7][23] ;
input \mem_a[7][22] ;
input \mem_a[7][21] ;
input \mem_a[7][20] ;
input \mem_a[7][19] ;
input \mem_a[7][18] ;
input \mem_a[7][17] ;
input \mem_a[7][16] ;
input \mem_a[7][15] ;
input \mem_a[7][14] ;
input \mem_a[7][13] ;
input \mem_a[7][12] ;
input \mem_a[7][11] ;
input \mem_a[7][10] ;
input \mem_a[7][9] ;
input \mem_a[7][8] ;
input \mem_a[7][7] ;
input \mem_a[7][6] ;
input \mem_a[7][5] ;
input \mem_a[7][4] ;
input \mem_a[7][3] ;
input \mem_a[7][2] ;
input \mem_a[7][1] ;
input \mem_a[7][0] ;
input \mem_a[8][63] ;
input \mem_a[8][62] ;
input \mem_a[8][61] ;
input \mem_a[8][60] ;
input \mem_a[8][59] ;
input \mem_a[8][58] ;
input \mem_a[8][57] ;
input \mem_a[8][56] ;
input \mem_a[8][55] ;
input \mem_a[8][54] ;
input \mem_a[8][53] ;
input \mem_a[8][52] ;
input \mem_a[8][51] ;
input \mem_a[8][50] ;
input \mem_a[8][49] ;
input \mem_a[8][48] ;
input \mem_a[8][47] ;
input \mem_a[8][46] ;
input \mem_a[8][45] ;
input \mem_a[8][44] ;
input \mem_a[8][43] ;
input \mem_a[8][42] ;
input \mem_a[8][41] ;
input \mem_a[8][40] ;
input \mem_a[8][39] ;
input \mem_a[8][38] ;
input \mem_a[8][37] ;
input \mem_a[8][36] ;
input \mem_a[8][35] ;
input \mem_a[8][34] ;
input \mem_a[8][33] ;
input \mem_a[8][32] ;
input \mem_a[8][31] ;
input \mem_a[8][30] ;
input \mem_a[8][29] ;
input \mem_a[8][28] ;
input \mem_a[8][27] ;
input \mem_a[8][26] ;
input \mem_a[8][25] ;
input \mem_a[8][24] ;
input \mem_a[8][23] ;
input \mem_a[8][22] ;
input \mem_a[8][21] ;
input \mem_a[8][20] ;
input \mem_a[8][19] ;
input \mem_a[8][18] ;
input \mem_a[8][17] ;
input \mem_a[8][16] ;
input \mem_a[8][15] ;
input \mem_a[8][14] ;
input \mem_a[8][13] ;
input \mem_a[8][12] ;
input \mem_a[8][11] ;
input \mem_a[8][10] ;
input \mem_a[8][9] ;
input \mem_a[8][8] ;
input \mem_a[8][7] ;
input \mem_a[8][6] ;
input \mem_a[8][5] ;
input \mem_a[8][4] ;
input \mem_a[8][3] ;
input \mem_a[8][2] ;
input \mem_a[8][1] ;
input \mem_a[8][0] ;
input \mem_a[9][63] ;
input \mem_a[9][62] ;
input \mem_a[9][61] ;
input \mem_a[9][60] ;
input \mem_a[9][59] ;
input \mem_a[9][58] ;
input \mem_a[9][57] ;
input \mem_a[9][56] ;
input \mem_a[9][55] ;
input \mem_a[9][54] ;
input \mem_a[9][53] ;
input \mem_a[9][52] ;
input \mem_a[9][51] ;
input \mem_a[9][50] ;
input \mem_a[9][49] ;
input \mem_a[9][48] ;
input \mem_a[9][47] ;
input \mem_a[9][46] ;
input \mem_a[9][45] ;
input \mem_a[9][44] ;
input \mem_a[9][43] ;
input \mem_a[9][42] ;
input \mem_a[9][41] ;
input \mem_a[9][40] ;
input \mem_a[9][39] ;
input \mem_a[9][38] ;
input \mem_a[9][37] ;
input \mem_a[9][36] ;
input \mem_a[9][35] ;
input \mem_a[9][34] ;
input \mem_a[9][33] ;
input \mem_a[9][32] ;
input \mem_a[9][31] ;
input \mem_a[9][30] ;
input \mem_a[9][29] ;
input \mem_a[9][28] ;
input \mem_a[9][27] ;
input \mem_a[9][26] ;
input \mem_a[9][25] ;
input \mem_a[9][24] ;
input \mem_a[9][23] ;
input \mem_a[9][22] ;
input \mem_a[9][21] ;
input \mem_a[9][20] ;
input \mem_a[9][19] ;
input \mem_a[9][18] ;
input \mem_a[9][17] ;
input \mem_a[9][16] ;
input \mem_a[9][15] ;
input \mem_a[9][14] ;
input \mem_a[9][13] ;
input \mem_a[9][12] ;
input \mem_a[9][11] ;
input \mem_a[9][10] ;
input \mem_a[9][9] ;
input \mem_a[9][8] ;
input \mem_a[9][7] ;
input \mem_a[9][6] ;
input \mem_a[9][5] ;
input \mem_a[9][4] ;
input \mem_a[9][3] ;
input \mem_a[9][2] ;
input \mem_a[9][1] ;
input \mem_a[9][0] ;
input \mem_a[10][63] ;
input \mem_a[10][62] ;
input \mem_a[10][61] ;
input \mem_a[10][60] ;
input \mem_a[10][59] ;
input \mem_a[10][58] ;
input \mem_a[10][57] ;
input \mem_a[10][56] ;
input \mem_a[10][55] ;
input \mem_a[10][54] ;
input \mem_a[10][53] ;
input \mem_a[10][52] ;
input \mem_a[10][51] ;
input \mem_a[10][50] ;
input \mem_a[10][49] ;
input \mem_a[10][48] ;
input \mem_a[10][47] ;
input \mem_a[10][46] ;
input \mem_a[10][45] ;
input \mem_a[10][44] ;
input \mem_a[10][43] ;
input \mem_a[10][42] ;
input \mem_a[10][41] ;
input \mem_a[10][40] ;
input \mem_a[10][39] ;
input \mem_a[10][38] ;
input \mem_a[10][37] ;
input \mem_a[10][36] ;
input \mem_a[10][35] ;
input \mem_a[10][34] ;
input \mem_a[10][33] ;
input \mem_a[10][32] ;
input \mem_a[10][31] ;
input \mem_a[10][30] ;
input \mem_a[10][29] ;
input \mem_a[10][28] ;
input \mem_a[10][27] ;
input \mem_a[10][26] ;
input \mem_a[10][25] ;
input \mem_a[10][24] ;
input \mem_a[10][23] ;
input \mem_a[10][22] ;
input \mem_a[10][21] ;
input \mem_a[10][20] ;
input \mem_a[10][19] ;
input \mem_a[10][18] ;
input \mem_a[10][17] ;
input \mem_a[10][16] ;
input \mem_a[10][15] ;
input \mem_a[10][14] ;
input \mem_a[10][13] ;
input \mem_a[10][12] ;
input \mem_a[10][11] ;
input \mem_a[10][10] ;
input \mem_a[10][9] ;
input \mem_a[10][8] ;
input \mem_a[10][7] ;
input \mem_a[10][6] ;
input \mem_a[10][5] ;
input \mem_a[10][4] ;
input \mem_a[10][3] ;
input \mem_a[10][2] ;
input \mem_a[10][1] ;
input \mem_a[10][0] ;
input \mem_a[11][63] ;
input \mem_a[11][62] ;
input \mem_a[11][61] ;
input \mem_a[11][60] ;
input \mem_a[11][59] ;
input \mem_a[11][58] ;
input \mem_a[11][57] ;
input \mem_a[11][56] ;
input \mem_a[11][55] ;
input \mem_a[11][54] ;
input \mem_a[11][53] ;
input \mem_a[11][52] ;
input \mem_a[11][51] ;
input \mem_a[11][50] ;
input \mem_a[11][49] ;
input \mem_a[11][48] ;
input \mem_a[11][47] ;
input \mem_a[11][46] ;
input \mem_a[11][45] ;
input \mem_a[11][44] ;
input \mem_a[11][43] ;
input \mem_a[11][42] ;
input \mem_a[11][41] ;
input \mem_a[11][40] ;
input \mem_a[11][39] ;
input \mem_a[11][38] ;
input \mem_a[11][37] ;
input \mem_a[11][36] ;
input \mem_a[11][35] ;
input \mem_a[11][34] ;
input \mem_a[11][33] ;
input \mem_a[11][32] ;
input \mem_a[11][31] ;
input \mem_a[11][30] ;
input \mem_a[11][29] ;
input \mem_a[11][28] ;
input \mem_a[11][27] ;
input \mem_a[11][26] ;
input \mem_a[11][25] ;
input \mem_a[11][24] ;
input \mem_a[11][23] ;
input \mem_a[11][22] ;
input \mem_a[11][21] ;
input \mem_a[11][20] ;
input \mem_a[11][19] ;
input \mem_a[11][18] ;
input \mem_a[11][17] ;
input \mem_a[11][16] ;
input \mem_a[11][15] ;
input \mem_a[11][14] ;
input \mem_a[11][13] ;
input \mem_a[11][12] ;
input \mem_a[11][11] ;
input \mem_a[11][10] ;
input \mem_a[11][9] ;
input \mem_a[11][8] ;
input \mem_a[11][7] ;
input \mem_a[11][6] ;
input \mem_a[11][5] ;
input \mem_a[11][4] ;
input \mem_a[11][3] ;
input \mem_a[11][2] ;
input \mem_a[11][1] ;
input \mem_a[11][0] ;
input \mem_a[12][63] ;
input \mem_a[12][62] ;
input \mem_a[12][61] ;
input \mem_a[12][60] ;
input \mem_a[12][59] ;
input \mem_a[12][58] ;
input \mem_a[12][57] ;
input \mem_a[12][56] ;
input \mem_a[12][55] ;
input \mem_a[12][54] ;
input \mem_a[12][53] ;
input \mem_a[12][52] ;
input \mem_a[12][51] ;
input \mem_a[12][50] ;
input \mem_a[12][49] ;
input \mem_a[12][48] ;
input \mem_a[12][47] ;
input \mem_a[12][46] ;
input \mem_a[12][45] ;
input \mem_a[12][44] ;
input \mem_a[12][43] ;
input \mem_a[12][42] ;
input \mem_a[12][41] ;
input \mem_a[12][40] ;
input \mem_a[12][39] ;
input \mem_a[12][38] ;
input \mem_a[12][37] ;
input \mem_a[12][36] ;
input \mem_a[12][35] ;
input \mem_a[12][34] ;
input \mem_a[12][33] ;
input \mem_a[12][32] ;
input \mem_a[12][31] ;
input \mem_a[12][30] ;
input \mem_a[12][29] ;
input \mem_a[12][28] ;
input \mem_a[12][27] ;
input \mem_a[12][26] ;
input \mem_a[12][25] ;
input \mem_a[12][24] ;
input \mem_a[12][23] ;
input \mem_a[12][22] ;
input \mem_a[12][21] ;
input \mem_a[12][20] ;
input \mem_a[12][19] ;
input \mem_a[12][18] ;
input \mem_a[12][17] ;
input \mem_a[12][16] ;
input \mem_a[12][15] ;
input \mem_a[12][14] ;
input \mem_a[12][13] ;
input \mem_a[12][12] ;
input \mem_a[12][11] ;
input \mem_a[12][10] ;
input \mem_a[12][9] ;
input \mem_a[12][8] ;
input \mem_a[12][7] ;
input \mem_a[12][6] ;
input \mem_a[12][5] ;
input \mem_a[12][4] ;
input \mem_a[12][3] ;
input \mem_a[12][2] ;
input \mem_a[12][1] ;
input \mem_a[12][0] ;
input \mem_a[13][63] ;
input \mem_a[13][62] ;
input \mem_a[13][61] ;
input \mem_a[13][60] ;
input \mem_a[13][59] ;
input \mem_a[13][58] ;
input \mem_a[13][57] ;
input \mem_a[13][56] ;
input \mem_a[13][55] ;
input \mem_a[13][54] ;
input \mem_a[13][53] ;
input \mem_a[13][52] ;
input \mem_a[13][51] ;
input \mem_a[13][50] ;
input \mem_a[13][49] ;
input \mem_a[13][48] ;
input \mem_a[13][47] ;
input \mem_a[13][46] ;
input \mem_a[13][45] ;
input \mem_a[13][44] ;
input \mem_a[13][43] ;
input \mem_a[13][42] ;
input \mem_a[13][41] ;
input \mem_a[13][40] ;
input \mem_a[13][39] ;
input \mem_a[13][38] ;
input \mem_a[13][37] ;
input \mem_a[13][36] ;
input \mem_a[13][35] ;
input \mem_a[13][34] ;
input \mem_a[13][33] ;
input \mem_a[13][32] ;
input \mem_a[13][31] ;
input \mem_a[13][30] ;
input \mem_a[13][29] ;
input \mem_a[13][28] ;
input \mem_a[13][27] ;
input \mem_a[13][26] ;
input \mem_a[13][25] ;
input \mem_a[13][24] ;
input \mem_a[13][23] ;
input \mem_a[13][22] ;
input \mem_a[13][21] ;
input \mem_a[13][20] ;
input \mem_a[13][19] ;
input \mem_a[13][18] ;
input \mem_a[13][17] ;
input \mem_a[13][16] ;
input \mem_a[13][15] ;
input \mem_a[13][14] ;
input \mem_a[13][13] ;
input \mem_a[13][12] ;
input \mem_a[13][11] ;
input \mem_a[13][10] ;
input \mem_a[13][9] ;
input \mem_a[13][8] ;
input \mem_a[13][7] ;
input \mem_a[13][6] ;
input \mem_a[13][5] ;
input \mem_a[13][4] ;
input \mem_a[13][3] ;
input \mem_a[13][2] ;
input \mem_a[13][1] ;
input \mem_a[13][0] ;
input \mem_a[14][63] ;
input \mem_a[14][62] ;
input \mem_a[14][61] ;
input \mem_a[14][60] ;
input \mem_a[14][59] ;
input \mem_a[14][58] ;
input \mem_a[14][57] ;
input \mem_a[14][56] ;
input \mem_a[14][55] ;
input \mem_a[14][54] ;
input \mem_a[14][53] ;
input \mem_a[14][52] ;
input \mem_a[14][51] ;
input \mem_a[14][50] ;
input \mem_a[14][49] ;
input \mem_a[14][48] ;
input \mem_a[14][47] ;
input \mem_a[14][46] ;
input \mem_a[14][45] ;
input \mem_a[14][44] ;
input \mem_a[14][43] ;
input \mem_a[14][42] ;
input \mem_a[14][41] ;
input \mem_a[14][40] ;
input \mem_a[14][39] ;
input \mem_a[14][38] ;
input \mem_a[14][37] ;
input \mem_a[14][36] ;
input \mem_a[14][35] ;
input \mem_a[14][34] ;
input \mem_a[14][33] ;
input \mem_a[14][32] ;
input \mem_a[14][31] ;
input \mem_a[14][30] ;
input \mem_a[14][29] ;
input \mem_a[14][28] ;
input \mem_a[14][27] ;
input \mem_a[14][26] ;
input \mem_a[14][25] ;
input \mem_a[14][24] ;
input \mem_a[14][23] ;
input \mem_a[14][22] ;
input \mem_a[14][21] ;
input \mem_a[14][20] ;
input \mem_a[14][19] ;
input \mem_a[14][18] ;
input \mem_a[14][17] ;
input \mem_a[14][16] ;
input \mem_a[14][15] ;
input \mem_a[14][14] ;
input \mem_a[14][13] ;
input \mem_a[14][12] ;
input \mem_a[14][11] ;
input \mem_a[14][10] ;
input \mem_a[14][9] ;
input \mem_a[14][8] ;
input \mem_a[14][7] ;
input \mem_a[14][6] ;
input \mem_a[14][5] ;
input \mem_a[14][4] ;
input \mem_a[14][3] ;
input \mem_a[14][2] ;
input \mem_a[14][1] ;
input \mem_a[14][0] ;
input \mem_a[15][63] ;
input \mem_a[15][62] ;
input \mem_a[15][61] ;
input \mem_a[15][60] ;
input \mem_a[15][59] ;
input \mem_a[15][58] ;
input \mem_a[15][57] ;
input \mem_a[15][56] ;
input \mem_a[15][55] ;
input \mem_a[15][54] ;
input \mem_a[15][53] ;
input \mem_a[15][52] ;
input \mem_a[15][51] ;
input \mem_a[15][50] ;
input \mem_a[15][49] ;
input \mem_a[15][48] ;
input \mem_a[15][47] ;
input \mem_a[15][46] ;
input \mem_a[15][45] ;
input \mem_a[15][44] ;
input \mem_a[15][43] ;
input \mem_a[15][42] ;
input \mem_a[15][41] ;
input \mem_a[15][40] ;
input \mem_a[15][39] ;
input \mem_a[15][38] ;
input \mem_a[15][37] ;
input \mem_a[15][36] ;
input \mem_a[15][35] ;
input \mem_a[15][34] ;
input \mem_a[15][33] ;
input \mem_a[15][32] ;
input \mem_a[15][31] ;
input \mem_a[15][30] ;
input \mem_a[15][29] ;
input \mem_a[15][28] ;
input \mem_a[15][27] ;
input \mem_a[15][26] ;
input \mem_a[15][25] ;
input \mem_a[15][24] ;
input \mem_a[15][23] ;
input \mem_a[15][22] ;
input \mem_a[15][21] ;
input \mem_a[15][20] ;
input \mem_a[15][19] ;
input \mem_a[15][18] ;
input \mem_a[15][17] ;
input \mem_a[15][16] ;
input \mem_a[15][15] ;
input \mem_a[15][14] ;
input \mem_a[15][13] ;
input \mem_a[15][12] ;
input \mem_a[15][11] ;
input \mem_a[15][10] ;
input \mem_a[15][9] ;
input \mem_a[15][8] ;
input \mem_a[15][7] ;
input \mem_a[15][6] ;
input \mem_a[15][5] ;
input \mem_a[15][4] ;
input \mem_a[15][3] ;
input \mem_a[15][2] ;
input \mem_a[15][1] ;
input \mem_a[15][0] ;
input \mem_a[16][63] ;
input \mem_a[16][62] ;
input \mem_a[16][61] ;
input \mem_a[16][60] ;
input \mem_a[16][59] ;
input \mem_a[16][58] ;
input \mem_a[16][57] ;
input \mem_a[16][56] ;
input \mem_a[16][55] ;
input \mem_a[16][54] ;
input \mem_a[16][53] ;
input \mem_a[16][52] ;
input \mem_a[16][51] ;
input \mem_a[16][50] ;
input \mem_a[16][49] ;
input \mem_a[16][48] ;
input \mem_a[16][47] ;
input \mem_a[16][46] ;
input \mem_a[16][45] ;
input \mem_a[16][44] ;
input \mem_a[16][43] ;
input \mem_a[16][42] ;
input \mem_a[16][41] ;
input \mem_a[16][40] ;
input \mem_a[16][39] ;
input \mem_a[16][38] ;
input \mem_a[16][37] ;
input \mem_a[16][36] ;
input \mem_a[16][35] ;
input \mem_a[16][34] ;
input \mem_a[16][33] ;
input \mem_a[16][32] ;
input \mem_a[16][31] ;
input \mem_a[16][30] ;
input \mem_a[16][29] ;
input \mem_a[16][28] ;
input \mem_a[16][27] ;
input \mem_a[16][26] ;
input \mem_a[16][25] ;
input \mem_a[16][24] ;
input \mem_a[16][23] ;
input \mem_a[16][22] ;
input \mem_a[16][21] ;
input \mem_a[16][20] ;
input \mem_a[16][19] ;
input \mem_a[16][18] ;
input \mem_a[16][17] ;
input \mem_a[16][16] ;
input \mem_a[16][15] ;
input \mem_a[16][14] ;
input \mem_a[16][13] ;
input \mem_a[16][12] ;
input \mem_a[16][11] ;
input \mem_a[16][10] ;
input \mem_a[16][9] ;
input \mem_a[16][8] ;
input \mem_a[16][7] ;
input \mem_a[16][6] ;
input \mem_a[16][5] ;
input \mem_a[16][4] ;
input \mem_a[16][3] ;
input \mem_a[16][2] ;
input \mem_a[16][1] ;
input \mem_a[16][0] ;
input \mem_a[17][63] ;
input \mem_a[17][62] ;
input \mem_a[17][61] ;
input \mem_a[17][60] ;
input \mem_a[17][59] ;
input \mem_a[17][58] ;
input \mem_a[17][57] ;
input \mem_a[17][56] ;
input \mem_a[17][55] ;
input \mem_a[17][54] ;
input \mem_a[17][53] ;
input \mem_a[17][52] ;
input \mem_a[17][51] ;
input \mem_a[17][50] ;
input \mem_a[17][49] ;
input \mem_a[17][48] ;
input \mem_a[17][47] ;
input \mem_a[17][46] ;
input \mem_a[17][45] ;
input \mem_a[17][44] ;
input \mem_a[17][43] ;
input \mem_a[17][42] ;
input \mem_a[17][41] ;
input \mem_a[17][40] ;
input \mem_a[17][39] ;
input \mem_a[17][38] ;
input \mem_a[17][37] ;
input \mem_a[17][36] ;
input \mem_a[17][35] ;
input \mem_a[17][34] ;
input \mem_a[17][33] ;
input \mem_a[17][32] ;
input \mem_a[17][31] ;
input \mem_a[17][30] ;
input \mem_a[17][29] ;
input \mem_a[17][28] ;
input \mem_a[17][27] ;
input \mem_a[17][26] ;
input \mem_a[17][25] ;
input \mem_a[17][24] ;
input \mem_a[17][23] ;
input \mem_a[17][22] ;
input \mem_a[17][21] ;
input \mem_a[17][20] ;
input \mem_a[17][19] ;
input \mem_a[17][18] ;
input \mem_a[17][17] ;
input \mem_a[17][16] ;
input \mem_a[17][15] ;
input \mem_a[17][14] ;
input \mem_a[17][13] ;
input \mem_a[17][12] ;
input \mem_a[17][11] ;
input \mem_a[17][10] ;
input \mem_a[17][9] ;
input \mem_a[17][8] ;
input \mem_a[17][7] ;
input \mem_a[17][6] ;
input \mem_a[17][5] ;
input \mem_a[17][4] ;
input \mem_a[17][3] ;
input \mem_a[17][2] ;
input \mem_a[17][1] ;
input \mem_a[17][0] ;
input \mem_a[18][63] ;
input \mem_a[18][62] ;
input \mem_a[18][61] ;
input \mem_a[18][60] ;
input \mem_a[18][59] ;
input \mem_a[18][58] ;
input \mem_a[18][57] ;
input \mem_a[18][56] ;
input \mem_a[18][55] ;
input \mem_a[18][54] ;
input \mem_a[18][53] ;
input \mem_a[18][52] ;
input \mem_a[18][51] ;
input \mem_a[18][50] ;
input \mem_a[18][49] ;
input \mem_a[18][48] ;
input \mem_a[18][47] ;
input \mem_a[18][46] ;
input \mem_a[18][45] ;
input \mem_a[18][44] ;
input \mem_a[18][43] ;
input \mem_a[18][42] ;
input \mem_a[18][41] ;
input \mem_a[18][40] ;
input \mem_a[18][39] ;
input \mem_a[18][38] ;
input \mem_a[18][37] ;
input \mem_a[18][36] ;
input \mem_a[18][35] ;
input \mem_a[18][34] ;
input \mem_a[18][33] ;
input \mem_a[18][32] ;
input \mem_a[18][31] ;
input \mem_a[18][30] ;
input \mem_a[18][29] ;
input \mem_a[18][28] ;
input \mem_a[18][27] ;
input \mem_a[18][26] ;
input \mem_a[18][25] ;
input \mem_a[18][24] ;
input \mem_a[18][23] ;
input \mem_a[18][22] ;
input \mem_a[18][21] ;
input \mem_a[18][20] ;
input \mem_a[18][19] ;
input \mem_a[18][18] ;
input \mem_a[18][17] ;
input \mem_a[18][16] ;
input \mem_a[18][15] ;
input \mem_a[18][14] ;
input \mem_a[18][13] ;
input \mem_a[18][12] ;
input \mem_a[18][11] ;
input \mem_a[18][10] ;
input \mem_a[18][9] ;
input \mem_a[18][8] ;
input \mem_a[18][7] ;
input \mem_a[18][6] ;
input \mem_a[18][5] ;
input \mem_a[18][4] ;
input \mem_a[18][3] ;
input \mem_a[18][2] ;
input \mem_a[18][1] ;
input \mem_a[18][0] ;
input \mem_a[19][63] ;
input \mem_a[19][62] ;
input \mem_a[19][61] ;
input \mem_a[19][60] ;
input \mem_a[19][59] ;
input \mem_a[19][58] ;
input \mem_a[19][57] ;
input \mem_a[19][56] ;
input \mem_a[19][55] ;
input \mem_a[19][54] ;
input \mem_a[19][53] ;
input \mem_a[19][52] ;
input \mem_a[19][51] ;
input \mem_a[19][50] ;
input \mem_a[19][49] ;
input \mem_a[19][48] ;
input \mem_a[19][47] ;
input \mem_a[19][46] ;
input \mem_a[19][45] ;
input \mem_a[19][44] ;
input \mem_a[19][43] ;
input \mem_a[19][42] ;
input \mem_a[19][41] ;
input \mem_a[19][40] ;
input \mem_a[19][39] ;
input \mem_a[19][38] ;
input \mem_a[19][37] ;
input \mem_a[19][36] ;
input \mem_a[19][35] ;
input \mem_a[19][34] ;
input \mem_a[19][33] ;
input \mem_a[19][32] ;
input \mem_a[19][31] ;
input \mem_a[19][30] ;
input \mem_a[19][29] ;
input \mem_a[19][28] ;
input \mem_a[19][27] ;
input \mem_a[19][26] ;
input \mem_a[19][25] ;
input \mem_a[19][24] ;
input \mem_a[19][23] ;
input \mem_a[19][22] ;
input \mem_a[19][21] ;
input \mem_a[19][20] ;
input \mem_a[19][19] ;
input \mem_a[19][18] ;
input \mem_a[19][17] ;
input \mem_a[19][16] ;
input \mem_a[19][15] ;
input \mem_a[19][14] ;
input \mem_a[19][13] ;
input \mem_a[19][12] ;
input \mem_a[19][11] ;
input \mem_a[19][10] ;
input \mem_a[19][9] ;
input \mem_a[19][8] ;
input \mem_a[19][7] ;
input \mem_a[19][6] ;
input \mem_a[19][5] ;
input \mem_a[19][4] ;
input \mem_a[19][3] ;
input \mem_a[19][2] ;
input \mem_a[19][1] ;
input \mem_a[19][0] ;
input \mem_a[20][63] ;
input \mem_a[20][62] ;
input \mem_a[20][61] ;
input \mem_a[20][60] ;
input \mem_a[20][59] ;
input \mem_a[20][58] ;
input \mem_a[20][57] ;
input \mem_a[20][56] ;
input \mem_a[20][55] ;
input \mem_a[20][54] ;
input \mem_a[20][53] ;
input \mem_a[20][52] ;
input \mem_a[20][51] ;
input \mem_a[20][50] ;
input \mem_a[20][49] ;
input \mem_a[20][48] ;
input \mem_a[20][47] ;
input \mem_a[20][46] ;
input \mem_a[20][45] ;
input \mem_a[20][44] ;
input \mem_a[20][43] ;
input \mem_a[20][42] ;
input \mem_a[20][41] ;
input \mem_a[20][40] ;
input \mem_a[20][39] ;
input \mem_a[20][38] ;
input \mem_a[20][37] ;
input \mem_a[20][36] ;
input \mem_a[20][35] ;
input \mem_a[20][34] ;
input \mem_a[20][33] ;
input \mem_a[20][32] ;
input \mem_a[20][31] ;
input \mem_a[20][30] ;
input \mem_a[20][29] ;
input \mem_a[20][28] ;
input \mem_a[20][27] ;
input \mem_a[20][26] ;
input \mem_a[20][25] ;
input \mem_a[20][24] ;
input \mem_a[20][23] ;
input \mem_a[20][22] ;
input \mem_a[20][21] ;
input \mem_a[20][20] ;
input \mem_a[20][19] ;
input \mem_a[20][18] ;
input \mem_a[20][17] ;
input \mem_a[20][16] ;
input \mem_a[20][15] ;
input \mem_a[20][14] ;
input \mem_a[20][13] ;
input \mem_a[20][12] ;
input \mem_a[20][11] ;
input \mem_a[20][10] ;
input \mem_a[20][9] ;
input \mem_a[20][8] ;
input \mem_a[20][7] ;
input \mem_a[20][6] ;
input \mem_a[20][5] ;
input \mem_a[20][4] ;
input \mem_a[20][3] ;
input \mem_a[20][2] ;
input \mem_a[20][1] ;
input \mem_a[20][0] ;
input \mem_a[21][63] ;
input \mem_a[21][62] ;
input \mem_a[21][61] ;
input \mem_a[21][60] ;
input \mem_a[21][59] ;
input \mem_a[21][58] ;
input \mem_a[21][57] ;
input \mem_a[21][56] ;
input \mem_a[21][55] ;
input \mem_a[21][54] ;
input \mem_a[21][53] ;
input \mem_a[21][52] ;
input \mem_a[21][51] ;
input \mem_a[21][50] ;
input \mem_a[21][49] ;
input \mem_a[21][48] ;
input \mem_a[21][47] ;
input \mem_a[21][46] ;
input \mem_a[21][45] ;
input \mem_a[21][44] ;
input \mem_a[21][43] ;
input \mem_a[21][42] ;
input \mem_a[21][41] ;
input \mem_a[21][40] ;
input \mem_a[21][39] ;
input \mem_a[21][38] ;
input \mem_a[21][37] ;
input \mem_a[21][36] ;
input \mem_a[21][35] ;
input \mem_a[21][34] ;
input \mem_a[21][33] ;
input \mem_a[21][32] ;
input \mem_a[21][31] ;
input \mem_a[21][30] ;
input \mem_a[21][29] ;
input \mem_a[21][28] ;
input \mem_a[21][27] ;
input \mem_a[21][26] ;
input \mem_a[21][25] ;
input \mem_a[21][24] ;
input \mem_a[21][23] ;
input \mem_a[21][22] ;
input \mem_a[21][21] ;
input \mem_a[21][20] ;
input \mem_a[21][19] ;
input \mem_a[21][18] ;
input \mem_a[21][17] ;
input \mem_a[21][16] ;
input \mem_a[21][15] ;
input \mem_a[21][14] ;
input \mem_a[21][13] ;
input \mem_a[21][12] ;
input \mem_a[21][11] ;
input \mem_a[21][10] ;
input \mem_a[21][9] ;
input \mem_a[21][8] ;
input \mem_a[21][7] ;
input \mem_a[21][6] ;
input \mem_a[21][5] ;
input \mem_a[21][4] ;
input \mem_a[21][3] ;
input \mem_a[21][2] ;
input \mem_a[21][1] ;
input \mem_a[21][0] ;
input \mem_a[22][63] ;
input \mem_a[22][62] ;
input \mem_a[22][61] ;
input \mem_a[22][60] ;
input \mem_a[22][59] ;
input \mem_a[22][58] ;
input \mem_a[22][57] ;
input \mem_a[22][56] ;
input \mem_a[22][55] ;
input \mem_a[22][54] ;
input \mem_a[22][53] ;
input \mem_a[22][52] ;
input \mem_a[22][51] ;
input \mem_a[22][50] ;
input \mem_a[22][49] ;
input \mem_a[22][48] ;
input \mem_a[22][47] ;
input \mem_a[22][46] ;
input \mem_a[22][45] ;
input \mem_a[22][44] ;
input \mem_a[22][43] ;
input \mem_a[22][42] ;
input \mem_a[22][41] ;
input \mem_a[22][40] ;
input \mem_a[22][39] ;
input \mem_a[22][38] ;
input \mem_a[22][37] ;
input \mem_a[22][36] ;
input \mem_a[22][35] ;
input \mem_a[22][34] ;
input \mem_a[22][33] ;
input \mem_a[22][32] ;
input \mem_a[22][31] ;
input \mem_a[22][30] ;
input \mem_a[22][29] ;
input \mem_a[22][28] ;
input \mem_a[22][27] ;
input \mem_a[22][26] ;
input \mem_a[22][25] ;
input \mem_a[22][24] ;
input \mem_a[22][23] ;
input \mem_a[22][22] ;
input \mem_a[22][21] ;
input \mem_a[22][20] ;
input \mem_a[22][19] ;
input \mem_a[22][18] ;
input \mem_a[22][17] ;
input \mem_a[22][16] ;
input \mem_a[22][15] ;
input \mem_a[22][14] ;
input \mem_a[22][13] ;
input \mem_a[22][12] ;
input \mem_a[22][11] ;
input \mem_a[22][10] ;
input \mem_a[22][9] ;
input \mem_a[22][8] ;
input \mem_a[22][7] ;
input \mem_a[22][6] ;
input \mem_a[22][5] ;
input \mem_a[22][4] ;
input \mem_a[22][3] ;
input \mem_a[22][2] ;
input \mem_a[22][1] ;
input \mem_a[22][0] ;
input \mem_a[23][63] ;
input \mem_a[23][62] ;
input \mem_a[23][61] ;
input \mem_a[23][60] ;
input \mem_a[23][59] ;
input \mem_a[23][58] ;
input \mem_a[23][57] ;
input \mem_a[23][56] ;
input \mem_a[23][55] ;
input \mem_a[23][54] ;
input \mem_a[23][53] ;
input \mem_a[23][52] ;
input \mem_a[23][51] ;
input \mem_a[23][50] ;
input \mem_a[23][49] ;
input \mem_a[23][48] ;
input \mem_a[23][47] ;
input \mem_a[23][46] ;
input \mem_a[23][45] ;
input \mem_a[23][44] ;
input \mem_a[23][43] ;
input \mem_a[23][42] ;
input \mem_a[23][41] ;
input \mem_a[23][40] ;
input \mem_a[23][39] ;
input \mem_a[23][38] ;
input \mem_a[23][37] ;
input \mem_a[23][36] ;
input \mem_a[23][35] ;
input \mem_a[23][34] ;
input \mem_a[23][33] ;
input \mem_a[23][32] ;
input \mem_a[23][31] ;
input \mem_a[23][30] ;
input \mem_a[23][29] ;
input \mem_a[23][28] ;
input \mem_a[23][27] ;
input \mem_a[23][26] ;
input \mem_a[23][25] ;
input \mem_a[23][24] ;
input \mem_a[23][23] ;
input \mem_a[23][22] ;
input \mem_a[23][21] ;
input \mem_a[23][20] ;
input \mem_a[23][19] ;
input \mem_a[23][18] ;
input \mem_a[23][17] ;
input \mem_a[23][16] ;
input \mem_a[23][15] ;
input \mem_a[23][14] ;
input \mem_a[23][13] ;
input \mem_a[23][12] ;
input \mem_a[23][11] ;
input \mem_a[23][10] ;
input \mem_a[23][9] ;
input \mem_a[23][8] ;
input \mem_a[23][7] ;
input \mem_a[23][6] ;
input \mem_a[23][5] ;
input \mem_a[23][4] ;
input \mem_a[23][3] ;
input \mem_a[23][2] ;
input \mem_a[23][1] ;
input \mem_a[23][0] ;
input \mem_a[24][63] ;
input \mem_a[24][62] ;
input \mem_a[24][61] ;
input \mem_a[24][60] ;
input \mem_a[24][59] ;
input \mem_a[24][58] ;
input \mem_a[24][57] ;
input \mem_a[24][56] ;
input \mem_a[24][55] ;
input \mem_a[24][54] ;
input \mem_a[24][53] ;
input \mem_a[24][52] ;
input \mem_a[24][51] ;
input \mem_a[24][50] ;
input \mem_a[24][49] ;
input \mem_a[24][48] ;
input \mem_a[24][47] ;
input \mem_a[24][46] ;
input \mem_a[24][45] ;
input \mem_a[24][44] ;
input \mem_a[24][43] ;
input \mem_a[24][42] ;
input \mem_a[24][41] ;
input \mem_a[24][40] ;
input \mem_a[24][39] ;
input \mem_a[24][38] ;
input \mem_a[24][37] ;
input \mem_a[24][36] ;
input \mem_a[24][35] ;
input \mem_a[24][34] ;
input \mem_a[24][33] ;
input \mem_a[24][32] ;
input \mem_a[24][31] ;
input \mem_a[24][30] ;
input \mem_a[24][29] ;
input \mem_a[24][28] ;
input \mem_a[24][27] ;
input \mem_a[24][26] ;
input \mem_a[24][25] ;
input \mem_a[24][24] ;
input \mem_a[24][23] ;
input \mem_a[24][22] ;
input \mem_a[24][21] ;
input \mem_a[24][20] ;
input \mem_a[24][19] ;
input \mem_a[24][18] ;
input \mem_a[24][17] ;
input \mem_a[24][16] ;
input \mem_a[24][15] ;
input \mem_a[24][14] ;
input \mem_a[24][13] ;
input \mem_a[24][12] ;
input \mem_a[24][11] ;
input \mem_a[24][10] ;
input \mem_a[24][9] ;
input \mem_a[24][8] ;
input \mem_a[24][7] ;
input \mem_a[24][6] ;
input \mem_a[24][5] ;
input \mem_a[24][4] ;
input \mem_a[24][3] ;
input \mem_a[24][2] ;
input \mem_a[24][1] ;
input \mem_a[24][0] ;
input \mem_a[25][63] ;
input \mem_a[25][62] ;
input \mem_a[25][61] ;
input \mem_a[25][60] ;
input \mem_a[25][59] ;
input \mem_a[25][58] ;
input \mem_a[25][57] ;
input \mem_a[25][56] ;
input \mem_a[25][55] ;
input \mem_a[25][54] ;
input \mem_a[25][53] ;
input \mem_a[25][52] ;
input \mem_a[25][51] ;
input \mem_a[25][50] ;
input \mem_a[25][49] ;
input \mem_a[25][48] ;
input \mem_a[25][47] ;
input \mem_a[25][46] ;
input \mem_a[25][45] ;
input \mem_a[25][44] ;
input \mem_a[25][43] ;
input \mem_a[25][42] ;
input \mem_a[25][41] ;
input \mem_a[25][40] ;
input \mem_a[25][39] ;
input \mem_a[25][38] ;
input \mem_a[25][37] ;
input \mem_a[25][36] ;
input \mem_a[25][35] ;
input \mem_a[25][34] ;
input \mem_a[25][33] ;
input \mem_a[25][32] ;
input \mem_a[25][31] ;
input \mem_a[25][30] ;
input \mem_a[25][29] ;
input \mem_a[25][28] ;
input \mem_a[25][27] ;
input \mem_a[25][26] ;
input \mem_a[25][25] ;
input \mem_a[25][24] ;
input \mem_a[25][23] ;
input \mem_a[25][22] ;
input \mem_a[25][21] ;
input \mem_a[25][20] ;
input \mem_a[25][19] ;
input \mem_a[25][18] ;
input \mem_a[25][17] ;
input \mem_a[25][16] ;
input \mem_a[25][15] ;
input \mem_a[25][14] ;
input \mem_a[25][13] ;
input \mem_a[25][12] ;
input \mem_a[25][11] ;
input \mem_a[25][10] ;
input \mem_a[25][9] ;
input \mem_a[25][8] ;
input \mem_a[25][7] ;
input \mem_a[25][6] ;
input \mem_a[25][5] ;
input \mem_a[25][4] ;
input \mem_a[25][3] ;
input \mem_a[25][2] ;
input \mem_a[25][1] ;
input \mem_a[25][0] ;
input \mem_a[26][63] ;
input \mem_a[26][62] ;
input \mem_a[26][61] ;
input \mem_a[26][60] ;
input \mem_a[26][59] ;
input \mem_a[26][58] ;
input \mem_a[26][57] ;
input \mem_a[26][56] ;
input \mem_a[26][55] ;
input \mem_a[26][54] ;
input \mem_a[26][53] ;
input \mem_a[26][52] ;
input \mem_a[26][51] ;
input \mem_a[26][50] ;
input \mem_a[26][49] ;
input \mem_a[26][48] ;
input \mem_a[26][47] ;
input \mem_a[26][46] ;
input \mem_a[26][45] ;
input \mem_a[26][44] ;
input \mem_a[26][43] ;
input \mem_a[26][42] ;
input \mem_a[26][41] ;
input \mem_a[26][40] ;
input \mem_a[26][39] ;
input \mem_a[26][38] ;
input \mem_a[26][37] ;
input \mem_a[26][36] ;
input \mem_a[26][35] ;
input \mem_a[26][34] ;
input \mem_a[26][33] ;
input \mem_a[26][32] ;
input \mem_a[26][31] ;
input \mem_a[26][30] ;
input \mem_a[26][29] ;
input \mem_a[26][28] ;
input \mem_a[26][27] ;
input \mem_a[26][26] ;
input \mem_a[26][25] ;
input \mem_a[26][24] ;
input \mem_a[26][23] ;
input \mem_a[26][22] ;
input \mem_a[26][21] ;
input \mem_a[26][20] ;
input \mem_a[26][19] ;
input \mem_a[26][18] ;
input \mem_a[26][17] ;
input \mem_a[26][16] ;
input \mem_a[26][15] ;
input \mem_a[26][14] ;
input \mem_a[26][13] ;
input \mem_a[26][12] ;
input \mem_a[26][11] ;
input \mem_a[26][10] ;
input \mem_a[26][9] ;
input \mem_a[26][8] ;
input \mem_a[26][7] ;
input \mem_a[26][6] ;
input \mem_a[26][5] ;
input \mem_a[26][4] ;
input \mem_a[26][3] ;
input \mem_a[26][2] ;
input \mem_a[26][1] ;
input \mem_a[26][0] ;
input \mem_a[27][63] ;
input \mem_a[27][62] ;
input \mem_a[27][61] ;
input \mem_a[27][60] ;
input \mem_a[27][59] ;
input \mem_a[27][58] ;
input \mem_a[27][57] ;
input \mem_a[27][56] ;
input \mem_a[27][55] ;
input \mem_a[27][54] ;
input \mem_a[27][53] ;
input \mem_a[27][52] ;
input \mem_a[27][51] ;
input \mem_a[27][50] ;
input \mem_a[27][49] ;
input \mem_a[27][48] ;
input \mem_a[27][47] ;
input \mem_a[27][46] ;
input \mem_a[27][45] ;
input \mem_a[27][44] ;
input \mem_a[27][43] ;
input \mem_a[27][42] ;
input \mem_a[27][41] ;
input \mem_a[27][40] ;
input \mem_a[27][39] ;
input \mem_a[27][38] ;
input \mem_a[27][37] ;
input \mem_a[27][36] ;
input \mem_a[27][35] ;
input \mem_a[27][34] ;
input \mem_a[27][33] ;
input \mem_a[27][32] ;
input \mem_a[27][31] ;
input \mem_a[27][30] ;
input \mem_a[27][29] ;
input \mem_a[27][28] ;
input \mem_a[27][27] ;
input \mem_a[27][26] ;
input \mem_a[27][25] ;
input \mem_a[27][24] ;
input \mem_a[27][23] ;
input \mem_a[27][22] ;
input \mem_a[27][21] ;
input \mem_a[27][20] ;
input \mem_a[27][19] ;
input \mem_a[27][18] ;
input \mem_a[27][17] ;
input \mem_a[27][16] ;
input \mem_a[27][15] ;
input \mem_a[27][14] ;
input \mem_a[27][13] ;
input \mem_a[27][12] ;
input \mem_a[27][11] ;
input \mem_a[27][10] ;
input \mem_a[27][9] ;
input \mem_a[27][8] ;
input \mem_a[27][7] ;
input \mem_a[27][6] ;
input \mem_a[27][5] ;
input \mem_a[27][4] ;
input \mem_a[27][3] ;
input \mem_a[27][2] ;
input \mem_a[27][1] ;
input \mem_a[27][0] ;
input \mem_a[28][63] ;
input \mem_a[28][62] ;
input \mem_a[28][61] ;
input \mem_a[28][60] ;
input \mem_a[28][59] ;
input \mem_a[28][58] ;
input \mem_a[28][57] ;
input \mem_a[28][56] ;
input \mem_a[28][55] ;
input \mem_a[28][54] ;
input \mem_a[28][53] ;
input \mem_a[28][52] ;
input \mem_a[28][51] ;
input \mem_a[28][50] ;
input \mem_a[28][49] ;
input \mem_a[28][48] ;
input \mem_a[28][47] ;
input \mem_a[28][46] ;
input \mem_a[28][45] ;
input \mem_a[28][44] ;
input \mem_a[28][43] ;
input \mem_a[28][42] ;
input \mem_a[28][41] ;
input \mem_a[28][40] ;
input \mem_a[28][39] ;
input \mem_a[28][38] ;
input \mem_a[28][37] ;
input \mem_a[28][36] ;
input \mem_a[28][35] ;
input \mem_a[28][34] ;
input \mem_a[28][33] ;
input \mem_a[28][32] ;
input \mem_a[28][31] ;
input \mem_a[28][30] ;
input \mem_a[28][29] ;
input \mem_a[28][28] ;
input \mem_a[28][27] ;
input \mem_a[28][26] ;
input \mem_a[28][25] ;
input \mem_a[28][24] ;
input \mem_a[28][23] ;
input \mem_a[28][22] ;
input \mem_a[28][21] ;
input \mem_a[28][20] ;
input \mem_a[28][19] ;
input \mem_a[28][18] ;
input \mem_a[28][17] ;
input \mem_a[28][16] ;
input \mem_a[28][15] ;
input \mem_a[28][14] ;
input \mem_a[28][13] ;
input \mem_a[28][12] ;
input \mem_a[28][11] ;
input \mem_a[28][10] ;
input \mem_a[28][9] ;
input \mem_a[28][8] ;
input \mem_a[28][7] ;
input \mem_a[28][6] ;
input \mem_a[28][5] ;
input \mem_a[28][4] ;
input \mem_a[28][3] ;
input \mem_a[28][2] ;
input \mem_a[28][1] ;
input \mem_a[28][0] ;
input \mem_a[29][63] ;
input \mem_a[29][62] ;
input \mem_a[29][61] ;
input \mem_a[29][60] ;
input \mem_a[29][59] ;
input \mem_a[29][58] ;
input \mem_a[29][57] ;
input \mem_a[29][56] ;
input \mem_a[29][55] ;
input \mem_a[29][54] ;
input \mem_a[29][53] ;
input \mem_a[29][52] ;
input \mem_a[29][51] ;
input \mem_a[29][50] ;
input \mem_a[29][49] ;
input \mem_a[29][48] ;
input \mem_a[29][47] ;
input \mem_a[29][46] ;
input \mem_a[29][45] ;
input \mem_a[29][44] ;
input \mem_a[29][43] ;
input \mem_a[29][42] ;
input \mem_a[29][41] ;
input \mem_a[29][40] ;
input \mem_a[29][39] ;
input \mem_a[29][38] ;
input \mem_a[29][37] ;
input \mem_a[29][36] ;
input \mem_a[29][35] ;
input \mem_a[29][34] ;
input \mem_a[29][33] ;
input \mem_a[29][32] ;
input \mem_a[29][31] ;
input \mem_a[29][30] ;
input \mem_a[29][29] ;
input \mem_a[29][28] ;
input \mem_a[29][27] ;
input \mem_a[29][26] ;
input \mem_a[29][25] ;
input \mem_a[29][24] ;
input \mem_a[29][23] ;
input \mem_a[29][22] ;
input \mem_a[29][21] ;
input \mem_a[29][20] ;
input \mem_a[29][19] ;
input \mem_a[29][18] ;
input \mem_a[29][17] ;
input \mem_a[29][16] ;
input \mem_a[29][15] ;
input \mem_a[29][14] ;
input \mem_a[29][13] ;
input \mem_a[29][12] ;
input \mem_a[29][11] ;
input \mem_a[29][10] ;
input \mem_a[29][9] ;
input \mem_a[29][8] ;
input \mem_a[29][7] ;
input \mem_a[29][6] ;
input \mem_a[29][5] ;
input \mem_a[29][4] ;
input \mem_a[29][3] ;
input \mem_a[29][2] ;
input \mem_a[29][1] ;
input \mem_a[29][0] ;
input \mem_a[30][63] ;
input \mem_a[30][62] ;
input \mem_a[30][61] ;
input \mem_a[30][60] ;
input \mem_a[30][59] ;
input \mem_a[30][58] ;
input \mem_a[30][57] ;
input \mem_a[30][56] ;
input \mem_a[30][55] ;
input \mem_a[30][54] ;
input \mem_a[30][53] ;
input \mem_a[30][52] ;
input \mem_a[30][51] ;
input \mem_a[30][50] ;
input \mem_a[30][49] ;
input \mem_a[30][48] ;
input \mem_a[30][47] ;
input \mem_a[30][46] ;
input \mem_a[30][45] ;
input \mem_a[30][44] ;
input \mem_a[30][43] ;
input \mem_a[30][42] ;
input \mem_a[30][41] ;
input \mem_a[30][40] ;
input \mem_a[30][39] ;
input \mem_a[30][38] ;
input \mem_a[30][37] ;
input \mem_a[30][36] ;
input \mem_a[30][35] ;
input \mem_a[30][34] ;
input \mem_a[30][33] ;
input \mem_a[30][32] ;
input \mem_a[30][31] ;
input \mem_a[30][30] ;
input \mem_a[30][29] ;
input \mem_a[30][28] ;
input \mem_a[30][27] ;
input \mem_a[30][26] ;
input \mem_a[30][25] ;
input \mem_a[30][24] ;
input \mem_a[30][23] ;
input \mem_a[30][22] ;
input \mem_a[30][21] ;
input \mem_a[30][20] ;
input \mem_a[30][19] ;
input \mem_a[30][18] ;
input \mem_a[30][17] ;
input \mem_a[30][16] ;
input \mem_a[30][15] ;
input \mem_a[30][14] ;
input \mem_a[30][13] ;
input \mem_a[30][12] ;
input \mem_a[30][11] ;
input \mem_a[30][10] ;
input \mem_a[30][9] ;
input \mem_a[30][8] ;
input \mem_a[30][7] ;
input \mem_a[30][6] ;
input \mem_a[30][5] ;
input \mem_a[30][4] ;
input \mem_a[30][3] ;
input \mem_a[30][2] ;
input \mem_a[30][1] ;
input \mem_a[30][0] ;
input \mem_a[31][63] ;
input \mem_a[31][62] ;
input \mem_a[31][61] ;
input \mem_a[31][60] ;
input \mem_a[31][59] ;
input \mem_a[31][58] ;
input \mem_a[31][57] ;
input \mem_a[31][56] ;
input \mem_a[31][55] ;
input \mem_a[31][54] ;
input \mem_a[31][53] ;
input \mem_a[31][52] ;
input \mem_a[31][51] ;
input \mem_a[31][50] ;
input \mem_a[31][49] ;
input \mem_a[31][48] ;
input \mem_a[31][47] ;
input \mem_a[31][46] ;
input \mem_a[31][45] ;
input \mem_a[31][44] ;
input \mem_a[31][43] ;
input \mem_a[31][42] ;
input \mem_a[31][41] ;
input \mem_a[31][40] ;
input \mem_a[31][39] ;
input \mem_a[31][38] ;
input \mem_a[31][37] ;
input \mem_a[31][36] ;
input \mem_a[31][35] ;
input \mem_a[31][34] ;
input \mem_a[31][33] ;
input \mem_a[31][32] ;
input \mem_a[31][31] ;
input \mem_a[31][30] ;
input \mem_a[31][29] ;
input \mem_a[31][28] ;
input \mem_a[31][27] ;
input \mem_a[31][26] ;
input \mem_a[31][25] ;
input \mem_a[31][24] ;
input \mem_a[31][23] ;
input \mem_a[31][22] ;
input \mem_a[31][21] ;
input \mem_a[31][20] ;
input \mem_a[31][19] ;
input \mem_a[31][18] ;
input \mem_a[31][17] ;
input \mem_a[31][16] ;
input \mem_a[31][15] ;
input \mem_a[31][14] ;
input \mem_a[31][13] ;
input \mem_a[31][12] ;
input \mem_a[31][11] ;
input \mem_a[31][10] ;
input \mem_a[31][9] ;
input \mem_a[31][8] ;
input \mem_a[31][7] ;
input \mem_a[31][6] ;
input \mem_a[31][5] ;
input \mem_a[31][4] ;
input \mem_a[31][3] ;
input \mem_a[31][2] ;
input \mem_a[31][1] ;
input \mem_a[31][0] ;
wire [0:2] _zy_simnet_stat_code_0_w$;
wire [0:4] _zy_simnet_stat_datawords_1_w$;
wire [0:4] _zy_simnet_stat_addr_2_w$;
wire [0:15] _zy_simnet_capability_lst_3_w$;
wire [0:3] _zy_simnet_capability_type_4_w$;
wire [0:63] _zy_simnet_rd_dat_5_w$;
wire _zy_simnet_cio_6;
wire [0:2] _zy_simnet_stat_code_7_w$;
wire [0:4] _zy_simnet_stat_datawords_8_w$;
wire [0:4] _zy_simnet_stat_addr_9_w$;
wire _zy_simnet_dio_10;
wire [0:15] _zy_simnet_capability_lst_11_w$;
wire [0:3] _zy_simnet_capability_type_12_w$;
wire _zy_simnet_dio_13;
wire [0:4] _zy_simnet_addr_limit_14_w$;
wire [0:63] _zy_simnet_cio_15;
wire [0:63] _zy_simnet_rd_dat_16_w$;
wire _zy_simnet_sw_cs_17_w$;
wire _zy_simnet_dio_18;
wire _zy_simnet_sw_we_19_w$;
wire [0:4] _zy_simnet_sw_add_20_w$;
wire [0:63] _zy_simnet_sw_wdat_21_w$;
wire [0:63] _zy_simnet_sw_rdat_22_w$;
wire _zy_simnet_cio_23;
wire [0:3] _zy_simnet_cio_24;
wire _zy_simnet_cio_25;
wire _zy_simnet_dio_26;
wire _zy_simnet_reset_27_w$;
wire reset;
wire [4:0] sw_add;
wire sw_cs;
wire [63:0] sw_wdat;
wire [63:0] sw_rdat;
wire sw_we;
wire [4:0] addr_limit;
wire [63:0] _svmls_var_L189_0;
wire [31:0] _svmls_mah_L0_0;
wire [31:0] _svmls_dummy_ret;
supply0 n1;
supply1 n2;
Q_BUF U0 ( .A(n2), .Z(_zy_simnet_cio_25));
Q_BUF U1 ( .A(n1), .Z(_zy_simnet_cio_24[3]));
Q_BUF U2 ( .A(n1), .Z(_zy_simnet_cio_24[2]));
Q_BUF U3 ( .A(n1), .Z(_zy_simnet_cio_24[1]));
Q_BUF U4 ( .A(n1), .Z(_zy_simnet_cio_24[0]));
Q_BUF U5 ( .A(n1), .Z(_zy_simnet_cio_23));
Q_BUF U6 ( .A(n1), .Z(_zy_simnet_cio_15[63]));
Q_BUF U7 ( .A(n1), .Z(_zy_simnet_cio_15[62]));
Q_BUF U8 ( .A(n1), .Z(_zy_simnet_cio_15[61]));
Q_BUF U9 ( .A(n1), .Z(_zy_simnet_cio_15[60]));
Q_BUF U10 ( .A(n1), .Z(_zy_simnet_cio_15[59]));
Q_BUF U11 ( .A(n1), .Z(_zy_simnet_cio_15[58]));
Q_BUF U12 ( .A(n1), .Z(_zy_simnet_cio_15[57]));
Q_BUF U13 ( .A(n1), .Z(_zy_simnet_cio_15[56]));
Q_BUF U14 ( .A(n1), .Z(_zy_simnet_cio_15[55]));
Q_BUF U15 ( .A(n1), .Z(_zy_simnet_cio_15[54]));
Q_BUF U16 ( .A(n1), .Z(_zy_simnet_cio_15[53]));
Q_BUF U17 ( .A(n1), .Z(_zy_simnet_cio_15[52]));
Q_BUF U18 ( .A(n1), .Z(_zy_simnet_cio_15[51]));
Q_BUF U19 ( .A(n1), .Z(_zy_simnet_cio_15[50]));
Q_BUF U20 ( .A(n1), .Z(_zy_simnet_cio_15[49]));
Q_BUF U21 ( .A(n1), .Z(_zy_simnet_cio_15[48]));
Q_BUF U22 ( .A(n1), .Z(_zy_simnet_cio_15[47]));
Q_BUF U23 ( .A(n1), .Z(_zy_simnet_cio_15[46]));
Q_BUF U24 ( .A(n1), .Z(_zy_simnet_cio_15[45]));
Q_BUF U25 ( .A(n1), .Z(_zy_simnet_cio_15[44]));
Q_BUF U26 ( .A(n1), .Z(_zy_simnet_cio_15[43]));
Q_BUF U27 ( .A(n1), .Z(_zy_simnet_cio_15[42]));
Q_BUF U28 ( .A(n1), .Z(_zy_simnet_cio_15[41]));
Q_BUF U29 ( .A(n1), .Z(_zy_simnet_cio_15[40]));
Q_BUF U30 ( .A(n1), .Z(_zy_simnet_cio_15[39]));
Q_BUF U31 ( .A(n1), .Z(_zy_simnet_cio_15[38]));
Q_BUF U32 ( .A(n1), .Z(_zy_simnet_cio_15[37]));
Q_BUF U33 ( .A(n1), .Z(_zy_simnet_cio_15[36]));
Q_BUF U34 ( .A(n1), .Z(_zy_simnet_cio_15[35]));
Q_BUF U35 ( .A(n1), .Z(_zy_simnet_cio_15[34]));
Q_BUF U36 ( .A(n1), .Z(_zy_simnet_cio_15[33]));
Q_BUF U37 ( .A(n1), .Z(_zy_simnet_cio_15[32]));
Q_BUF U38 ( .A(n1), .Z(_zy_simnet_cio_15[31]));
Q_BUF U39 ( .A(n1), .Z(_zy_simnet_cio_15[30]));
Q_BUF U40 ( .A(n1), .Z(_zy_simnet_cio_15[29]));
Q_BUF U41 ( .A(n1), .Z(_zy_simnet_cio_15[28]));
Q_BUF U42 ( .A(n1), .Z(_zy_simnet_cio_15[27]));
Q_BUF U43 ( .A(n1), .Z(_zy_simnet_cio_15[26]));
Q_BUF U44 ( .A(n1), .Z(_zy_simnet_cio_15[25]));
Q_BUF U45 ( .A(n1), .Z(_zy_simnet_cio_15[24]));
Q_BUF U46 ( .A(n1), .Z(_zy_simnet_cio_15[23]));
Q_BUF U47 ( .A(n1), .Z(_zy_simnet_cio_15[22]));
Q_BUF U48 ( .A(n1), .Z(_zy_simnet_cio_15[21]));
Q_BUF U49 ( .A(n1), .Z(_zy_simnet_cio_15[20]));
Q_BUF U50 ( .A(n1), .Z(_zy_simnet_cio_15[19]));
Q_BUF U51 ( .A(n1), .Z(_zy_simnet_cio_15[18]));
Q_BUF U52 ( .A(n1), .Z(_zy_simnet_cio_15[17]));
Q_BUF U53 ( .A(n1), .Z(_zy_simnet_cio_15[16]));
Q_BUF U54 ( .A(n1), .Z(_zy_simnet_cio_15[15]));
Q_BUF U55 ( .A(n1), .Z(_zy_simnet_cio_15[14]));
Q_BUF U56 ( .A(n1), .Z(_zy_simnet_cio_15[13]));
Q_BUF U57 ( .A(n1), .Z(_zy_simnet_cio_15[12]));
Q_BUF U58 ( .A(n1), .Z(_zy_simnet_cio_15[11]));
Q_BUF U59 ( .A(n1), .Z(_zy_simnet_cio_15[10]));
Q_BUF U60 ( .A(n1), .Z(_zy_simnet_cio_15[9]));
Q_BUF U61 ( .A(n1), .Z(_zy_simnet_cio_15[8]));
Q_BUF U62 ( .A(n1), .Z(_zy_simnet_cio_15[7]));
Q_BUF U63 ( .A(n1), .Z(_zy_simnet_cio_15[6]));
Q_BUF U64 ( .A(n1), .Z(_zy_simnet_cio_15[5]));
Q_BUF U65 ( .A(n1), .Z(_zy_simnet_cio_15[4]));
Q_BUF U66 ( .A(n1), .Z(_zy_simnet_cio_15[3]));
Q_BUF U67 ( .A(n1), .Z(_zy_simnet_cio_15[2]));
Q_BUF U68 ( .A(n1), .Z(_zy_simnet_cio_15[1]));
Q_BUF U69 ( .A(n1), .Z(_zy_simnet_cio_15[0]));
Q_BUF U70 ( .A(n1), .Z(_zy_simnet_cio_6));
Q_BUF U71 ( .A(n2), .Z(addr_limit[0]));
Q_BUF U72 ( .A(n2), .Z(addr_limit[1]));
Q_BUF U73 ( .A(n2), .Z(addr_limit[2]));
Q_BUF U74 ( .A(n2), .Z(addr_limit[3]));
Q_BUF U75 ( .A(n2), .Z(addr_limit[4]));
nx_indirect_access_cntrl_xcm113 u_cntrl ( .clk( clk), .rst_n( rst_n), 
	.wr_stb( wr_stb), .reg_addr( addr[10:0]), .cmnd_op( cmnd_op[3:0]), 
	.cmnd_addr( cmnd_addr[4:0]), .cmnd_table_id( _zy_simnet_cio_6), 
	.stat_code( _zy_simnet_stat_code_7_w$[0:2]), .stat_datawords( 
	_zy_simnet_stat_datawords_8_w$[0:4]), .stat_addr( 
	_zy_simnet_stat_addr_9_w$[0:4]), .stat_table_id( _zy_simnet_dio_10), 
	.capability_lst( _zy_simnet_capability_lst_11_w$[0:15]), 
	.capability_type( _zy_simnet_capability_type_12_w$[0:3]), .enable( 
	_zy_simnet_dio_13), .addr_limit( _zy_simnet_addr_limit_14_w$[0:4]), 
	.wr_dat( _zy_simnet_cio_15[0:63]), .rd_dat( 
	_zy_simnet_rd_dat_16_w$[0:63]), .sw_cs( _zy_simnet_sw_cs_17_w$), 
	.sw_ce( _zy_simnet_dio_18), .sw_we( _zy_simnet_sw_we_19_w$), 
	.sw_add( _zy_simnet_sw_add_20_w$[0:4]), .sw_wdat( 
	_zy_simnet_sw_wdat_21_w$[0:63]), .sw_rdat( 
	_zy_simnet_sw_rdat_22_w$[0:63]), .sw_match( _zy_simnet_cio_23), 
	.sw_aindex( _zy_simnet_cio_24[0:3]), .grant( _zy_simnet_cio_25), 
	.yield( _zy_simnet_dio_26), .reset( _zy_simnet_reset_27_w$));
ixc_context_read_2048 _zzixc_ctxrd_0 ( { \_zyixc_ctx_rdata_29[0][63] , 
	\_zyixc_ctx_rdata_29[0][62] , \_zyixc_ctx_rdata_29[0][61] , 
	\_zyixc_ctx_rdata_29[0][60] , \_zyixc_ctx_rdata_29[0][59] , 
	\_zyixc_ctx_rdata_29[0][58] , \_zyixc_ctx_rdata_29[0][57] , 
	\_zyixc_ctx_rdata_29[0][56] , \_zyixc_ctx_rdata_29[0][55] , 
	\_zyixc_ctx_rdata_29[0][54] , \_zyixc_ctx_rdata_29[0][53] , 
	\_zyixc_ctx_rdata_29[0][52] , \_zyixc_ctx_rdata_29[0][51] , 
	\_zyixc_ctx_rdata_29[0][50] , \_zyixc_ctx_rdata_29[0][49] , 
	\_zyixc_ctx_rdata_29[0][48] , \_zyixc_ctx_rdata_29[0][47] , 
	\_zyixc_ctx_rdata_29[0][46] , \_zyixc_ctx_rdata_29[0][45] , 
	\_zyixc_ctx_rdata_29[0][44] , \_zyixc_ctx_rdata_29[0][43] , 
	\_zyixc_ctx_rdata_29[0][42] , \_zyixc_ctx_rdata_29[0][41] , 
	\_zyixc_ctx_rdata_29[0][40] , \_zyixc_ctx_rdata_29[0][39] , 
	\_zyixc_ctx_rdata_29[0][38] , \_zyixc_ctx_rdata_29[0][37] , 
	\_zyixc_ctx_rdata_29[0][36] , \_zyixc_ctx_rdata_29[0][35] , 
	\_zyixc_ctx_rdata_29[0][34] , \_zyixc_ctx_rdata_29[0][33] , 
	\_zyixc_ctx_rdata_29[0][32] , \_zyixc_ctx_rdata_29[0][31] , 
	\_zyixc_ctx_rdata_29[0][30] , \_zyixc_ctx_rdata_29[0][29] , 
	\_zyixc_ctx_rdata_29[0][28] , \_zyixc_ctx_rdata_29[0][27] , 
	\_zyixc_ctx_rdata_29[0][26] , \_zyixc_ctx_rdata_29[0][25] , 
	\_zyixc_ctx_rdata_29[0][24] , \_zyixc_ctx_rdata_29[0][23] , 
	\_zyixc_ctx_rdata_29[0][22] , \_zyixc_ctx_rdata_29[0][21] , 
	\_zyixc_ctx_rdata_29[0][20] , \_zyixc_ctx_rdata_29[0][19] , 
	\_zyixc_ctx_rdata_29[0][18] , \_zyixc_ctx_rdata_29[0][17] , 
	\_zyixc_ctx_rdata_29[0][16] , \_zyixc_ctx_rdata_29[0][15] , 
	\_zyixc_ctx_rdata_29[0][14] , \_zyixc_ctx_rdata_29[0][13] , 
	\_zyixc_ctx_rdata_29[0][12] , \_zyixc_ctx_rdata_29[0][11] , 
	\_zyixc_ctx_rdata_29[0][10] , \_zyixc_ctx_rdata_29[0][9] , 
	\_zyixc_ctx_rdata_29[0][8] , \_zyixc_ctx_rdata_29[0][7] , 
	\_zyixc_ctx_rdata_29[0][6] , \_zyixc_ctx_rdata_29[0][5] , 
	\_zyixc_ctx_rdata_29[0][4] , \_zyixc_ctx_rdata_29[0][3] , 
	\_zyixc_ctx_rdata_29[0][2] , \_zyixc_ctx_rdata_29[0][1] , 
	\_zyixc_ctx_rdata_29[0][0] , \_zyixc_ctx_rdata_29[1][63] , 
	\_zyixc_ctx_rdata_29[1][62] , \_zyixc_ctx_rdata_29[1][61] , 
	\_zyixc_ctx_rdata_29[1][60] , \_zyixc_ctx_rdata_29[1][59] , 
	\_zyixc_ctx_rdata_29[1][58] , \_zyixc_ctx_rdata_29[1][57] , 
	\_zyixc_ctx_rdata_29[1][56] , \_zyixc_ctx_rdata_29[1][55] , 
	\_zyixc_ctx_rdata_29[1][54] , \_zyixc_ctx_rdata_29[1][53] , 
	\_zyixc_ctx_rdata_29[1][52] , \_zyixc_ctx_rdata_29[1][51] , 
	\_zyixc_ctx_rdata_29[1][50] , \_zyixc_ctx_rdata_29[1][49] , 
	\_zyixc_ctx_rdata_29[1][48] , \_zyixc_ctx_rdata_29[1][47] , 
	\_zyixc_ctx_rdata_29[1][46] , \_zyixc_ctx_rdata_29[1][45] , 
	\_zyixc_ctx_rdata_29[1][44] , \_zyixc_ctx_rdata_29[1][43] , 
	\_zyixc_ctx_rdata_29[1][42] , \_zyixc_ctx_rdata_29[1][41] , 
	\_zyixc_ctx_rdata_29[1][40] , \_zyixc_ctx_rdata_29[1][39] , 
	\_zyixc_ctx_rdata_29[1][38] , \_zyixc_ctx_rdata_29[1][37] , 
	\_zyixc_ctx_rdata_29[1][36] , \_zyixc_ctx_rdata_29[1][35] , 
	\_zyixc_ctx_rdata_29[1][34] , \_zyixc_ctx_rdata_29[1][33] , 
	\_zyixc_ctx_rdata_29[1][32] , \_zyixc_ctx_rdata_29[1][31] , 
	\_zyixc_ctx_rdata_29[1][30] , \_zyixc_ctx_rdata_29[1][29] , 
	\_zyixc_ctx_rdata_29[1][28] , \_zyixc_ctx_rdata_29[1][27] , 
	\_zyixc_ctx_rdata_29[1][26] , \_zyixc_ctx_rdata_29[1][25] , 
	\_zyixc_ctx_rdata_29[1][24] , \_zyixc_ctx_rdata_29[1][23] , 
	\_zyixc_ctx_rdata_29[1][22] , \_zyixc_ctx_rdata_29[1][21] , 
	\_zyixc_ctx_rdata_29[1][20] , \_zyixc_ctx_rdata_29[1][19] , 
	\_zyixc_ctx_rdata_29[1][18] , \_zyixc_ctx_rdata_29[1][17] , 
	\_zyixc_ctx_rdata_29[1][16] , \_zyixc_ctx_rdata_29[1][15] , 
	\_zyixc_ctx_rdata_29[1][14] , \_zyixc_ctx_rdata_29[1][13] , 
	\_zyixc_ctx_rdata_29[1][12] , \_zyixc_ctx_rdata_29[1][11] , 
	\_zyixc_ctx_rdata_29[1][10] , \_zyixc_ctx_rdata_29[1][9] , 
	\_zyixc_ctx_rdata_29[1][8] , \_zyixc_ctx_rdata_29[1][7] , 
	\_zyixc_ctx_rdata_29[1][6] , \_zyixc_ctx_rdata_29[1][5] , 
	\_zyixc_ctx_rdata_29[1][4] , \_zyixc_ctx_rdata_29[1][3] , 
	\_zyixc_ctx_rdata_29[1][2] , \_zyixc_ctx_rdata_29[1][1] , 
	\_zyixc_ctx_rdata_29[1][0] , \_zyixc_ctx_rdata_29[2][63] , 
	\_zyixc_ctx_rdata_29[2][62] , \_zyixc_ctx_rdata_29[2][61] , 
	\_zyixc_ctx_rdata_29[2][60] , \_zyixc_ctx_rdata_29[2][59] , 
	\_zyixc_ctx_rdata_29[2][58] , \_zyixc_ctx_rdata_29[2][57] , 
	\_zyixc_ctx_rdata_29[2][56] , \_zyixc_ctx_rdata_29[2][55] , 
	\_zyixc_ctx_rdata_29[2][54] , \_zyixc_ctx_rdata_29[2][53] , 
	\_zyixc_ctx_rdata_29[2][52] , \_zyixc_ctx_rdata_29[2][51] , 
	\_zyixc_ctx_rdata_29[2][50] , \_zyixc_ctx_rdata_29[2][49] , 
	\_zyixc_ctx_rdata_29[2][48] , \_zyixc_ctx_rdata_29[2][47] , 
	\_zyixc_ctx_rdata_29[2][46] , \_zyixc_ctx_rdata_29[2][45] , 
	\_zyixc_ctx_rdata_29[2][44] , \_zyixc_ctx_rdata_29[2][43] , 
	\_zyixc_ctx_rdata_29[2][42] , \_zyixc_ctx_rdata_29[2][41] , 
	\_zyixc_ctx_rdata_29[2][40] , \_zyixc_ctx_rdata_29[2][39] , 
	\_zyixc_ctx_rdata_29[2][38] , \_zyixc_ctx_rdata_29[2][37] , 
	\_zyixc_ctx_rdata_29[2][36] , \_zyixc_ctx_rdata_29[2][35] , 
	\_zyixc_ctx_rdata_29[2][34] , \_zyixc_ctx_rdata_29[2][33] , 
	\_zyixc_ctx_rdata_29[2][32] , \_zyixc_ctx_rdata_29[2][31] , 
	\_zyixc_ctx_rdata_29[2][30] , \_zyixc_ctx_rdata_29[2][29] , 
	\_zyixc_ctx_rdata_29[2][28] , \_zyixc_ctx_rdata_29[2][27] , 
	\_zyixc_ctx_rdata_29[2][26] , \_zyixc_ctx_rdata_29[2][25] , 
	\_zyixc_ctx_rdata_29[2][24] , \_zyixc_ctx_rdata_29[2][23] , 
	\_zyixc_ctx_rdata_29[2][22] , \_zyixc_ctx_rdata_29[2][21] , 
	\_zyixc_ctx_rdata_29[2][20] , \_zyixc_ctx_rdata_29[2][19] , 
	\_zyixc_ctx_rdata_29[2][18] , \_zyixc_ctx_rdata_29[2][17] , 
	\_zyixc_ctx_rdata_29[2][16] , \_zyixc_ctx_rdata_29[2][15] , 
	\_zyixc_ctx_rdata_29[2][14] , \_zyixc_ctx_rdata_29[2][13] , 
	\_zyixc_ctx_rdata_29[2][12] , \_zyixc_ctx_rdata_29[2][11] , 
	\_zyixc_ctx_rdata_29[2][10] , \_zyixc_ctx_rdata_29[2][9] , 
	\_zyixc_ctx_rdata_29[2][8] , \_zyixc_ctx_rdata_29[2][7] , 
	\_zyixc_ctx_rdata_29[2][6] , \_zyixc_ctx_rdata_29[2][5] , 
	\_zyixc_ctx_rdata_29[2][4] , \_zyixc_ctx_rdata_29[2][3] , 
	\_zyixc_ctx_rdata_29[2][2] , \_zyixc_ctx_rdata_29[2][1] , 
	\_zyixc_ctx_rdata_29[2][0] , \_zyixc_ctx_rdata_29[3][63] , 
	\_zyixc_ctx_rdata_29[3][62] , \_zyixc_ctx_rdata_29[3][61] , 
	\_zyixc_ctx_rdata_29[3][60] , \_zyixc_ctx_rdata_29[3][59] , 
	\_zyixc_ctx_rdata_29[3][58] , \_zyixc_ctx_rdata_29[3][57] , 
	\_zyixc_ctx_rdata_29[3][56] , \_zyixc_ctx_rdata_29[3][55] , 
	\_zyixc_ctx_rdata_29[3][54] , \_zyixc_ctx_rdata_29[3][53] , 
	\_zyixc_ctx_rdata_29[3][52] , \_zyixc_ctx_rdata_29[3][51] , 
	\_zyixc_ctx_rdata_29[3][50] , \_zyixc_ctx_rdata_29[3][49] , 
	\_zyixc_ctx_rdata_29[3][48] , \_zyixc_ctx_rdata_29[3][47] , 
	\_zyixc_ctx_rdata_29[3][46] , \_zyixc_ctx_rdata_29[3][45] , 
	\_zyixc_ctx_rdata_29[3][44] , \_zyixc_ctx_rdata_29[3][43] , 
	\_zyixc_ctx_rdata_29[3][42] , \_zyixc_ctx_rdata_29[3][41] , 
	\_zyixc_ctx_rdata_29[3][40] , \_zyixc_ctx_rdata_29[3][39] , 
	\_zyixc_ctx_rdata_29[3][38] , \_zyixc_ctx_rdata_29[3][37] , 
	\_zyixc_ctx_rdata_29[3][36] , \_zyixc_ctx_rdata_29[3][35] , 
	\_zyixc_ctx_rdata_29[3][34] , \_zyixc_ctx_rdata_29[3][33] , 
	\_zyixc_ctx_rdata_29[3][32] , \_zyixc_ctx_rdata_29[3][31] , 
	\_zyixc_ctx_rdata_29[3][30] , \_zyixc_ctx_rdata_29[3][29] , 
	\_zyixc_ctx_rdata_29[3][28] , \_zyixc_ctx_rdata_29[3][27] , 
	\_zyixc_ctx_rdata_29[3][26] , \_zyixc_ctx_rdata_29[3][25] , 
	\_zyixc_ctx_rdata_29[3][24] , \_zyixc_ctx_rdata_29[3][23] , 
	\_zyixc_ctx_rdata_29[3][22] , \_zyixc_ctx_rdata_29[3][21] , 
	\_zyixc_ctx_rdata_29[3][20] , \_zyixc_ctx_rdata_29[3][19] , 
	\_zyixc_ctx_rdata_29[3][18] , \_zyixc_ctx_rdata_29[3][17] , 
	\_zyixc_ctx_rdata_29[3][16] , \_zyixc_ctx_rdata_29[3][15] , 
	\_zyixc_ctx_rdata_29[3][14] , \_zyixc_ctx_rdata_29[3][13] , 
	\_zyixc_ctx_rdata_29[3][12] , \_zyixc_ctx_rdata_29[3][11] , 
	\_zyixc_ctx_rdata_29[3][10] , \_zyixc_ctx_rdata_29[3][9] , 
	\_zyixc_ctx_rdata_29[3][8] , \_zyixc_ctx_rdata_29[3][7] , 
	\_zyixc_ctx_rdata_29[3][6] , \_zyixc_ctx_rdata_29[3][5] , 
	\_zyixc_ctx_rdata_29[3][4] , \_zyixc_ctx_rdata_29[3][3] , 
	\_zyixc_ctx_rdata_29[3][2] , \_zyixc_ctx_rdata_29[3][1] , 
	\_zyixc_ctx_rdata_29[3][0] , \_zyixc_ctx_rdata_29[4][63] , 
	\_zyixc_ctx_rdata_29[4][62] , \_zyixc_ctx_rdata_29[4][61] , 
	\_zyixc_ctx_rdata_29[4][60] , \_zyixc_ctx_rdata_29[4][59] , 
	\_zyixc_ctx_rdata_29[4][58] , \_zyixc_ctx_rdata_29[4][57] , 
	\_zyixc_ctx_rdata_29[4][56] , \_zyixc_ctx_rdata_29[4][55] , 
	\_zyixc_ctx_rdata_29[4][54] , \_zyixc_ctx_rdata_29[4][53] , 
	\_zyixc_ctx_rdata_29[4][52] , \_zyixc_ctx_rdata_29[4][51] , 
	\_zyixc_ctx_rdata_29[4][50] , \_zyixc_ctx_rdata_29[4][49] , 
	\_zyixc_ctx_rdata_29[4][48] , \_zyixc_ctx_rdata_29[4][47] , 
	\_zyixc_ctx_rdata_29[4][46] , \_zyixc_ctx_rdata_29[4][45] , 
	\_zyixc_ctx_rdata_29[4][44] , \_zyixc_ctx_rdata_29[4][43] , 
	\_zyixc_ctx_rdata_29[4][42] , \_zyixc_ctx_rdata_29[4][41] , 
	\_zyixc_ctx_rdata_29[4][40] , \_zyixc_ctx_rdata_29[4][39] , 
	\_zyixc_ctx_rdata_29[4][38] , \_zyixc_ctx_rdata_29[4][37] , 
	\_zyixc_ctx_rdata_29[4][36] , \_zyixc_ctx_rdata_29[4][35] , 
	\_zyixc_ctx_rdata_29[4][34] , \_zyixc_ctx_rdata_29[4][33] , 
	\_zyixc_ctx_rdata_29[4][32] , \_zyixc_ctx_rdata_29[4][31] , 
	\_zyixc_ctx_rdata_29[4][30] , \_zyixc_ctx_rdata_29[4][29] , 
	\_zyixc_ctx_rdata_29[4][28] , \_zyixc_ctx_rdata_29[4][27] , 
	\_zyixc_ctx_rdata_29[4][26] , \_zyixc_ctx_rdata_29[4][25] , 
	\_zyixc_ctx_rdata_29[4][24] , \_zyixc_ctx_rdata_29[4][23] , 
	\_zyixc_ctx_rdata_29[4][22] , \_zyixc_ctx_rdata_29[4][21] , 
	\_zyixc_ctx_rdata_29[4][20] , \_zyixc_ctx_rdata_29[4][19] , 
	\_zyixc_ctx_rdata_29[4][18] , \_zyixc_ctx_rdata_29[4][17] , 
	\_zyixc_ctx_rdata_29[4][16] , \_zyixc_ctx_rdata_29[4][15] , 
	\_zyixc_ctx_rdata_29[4][14] , \_zyixc_ctx_rdata_29[4][13] , 
	\_zyixc_ctx_rdata_29[4][12] , \_zyixc_ctx_rdata_29[4][11] , 
	\_zyixc_ctx_rdata_29[4][10] , \_zyixc_ctx_rdata_29[4][9] , 
	\_zyixc_ctx_rdata_29[4][8] , \_zyixc_ctx_rdata_29[4][7] , 
	\_zyixc_ctx_rdata_29[4][6] , \_zyixc_ctx_rdata_29[4][5] , 
	\_zyixc_ctx_rdata_29[4][4] , \_zyixc_ctx_rdata_29[4][3] , 
	\_zyixc_ctx_rdata_29[4][2] , \_zyixc_ctx_rdata_29[4][1] , 
	\_zyixc_ctx_rdata_29[4][0] , \_zyixc_ctx_rdata_29[5][63] , 
	\_zyixc_ctx_rdata_29[5][62] , \_zyixc_ctx_rdata_29[5][61] , 
	\_zyixc_ctx_rdata_29[5][60] , \_zyixc_ctx_rdata_29[5][59] , 
	\_zyixc_ctx_rdata_29[5][58] , \_zyixc_ctx_rdata_29[5][57] , 
	\_zyixc_ctx_rdata_29[5][56] , \_zyixc_ctx_rdata_29[5][55] , 
	\_zyixc_ctx_rdata_29[5][54] , \_zyixc_ctx_rdata_29[5][53] , 
	\_zyixc_ctx_rdata_29[5][52] , \_zyixc_ctx_rdata_29[5][51] , 
	\_zyixc_ctx_rdata_29[5][50] , \_zyixc_ctx_rdata_29[5][49] , 
	\_zyixc_ctx_rdata_29[5][48] , \_zyixc_ctx_rdata_29[5][47] , 
	\_zyixc_ctx_rdata_29[5][46] , \_zyixc_ctx_rdata_29[5][45] , 
	\_zyixc_ctx_rdata_29[5][44] , \_zyixc_ctx_rdata_29[5][43] , 
	\_zyixc_ctx_rdata_29[5][42] , \_zyixc_ctx_rdata_29[5][41] , 
	\_zyixc_ctx_rdata_29[5][40] , \_zyixc_ctx_rdata_29[5][39] , 
	\_zyixc_ctx_rdata_29[5][38] , \_zyixc_ctx_rdata_29[5][37] , 
	\_zyixc_ctx_rdata_29[5][36] , \_zyixc_ctx_rdata_29[5][35] , 
	\_zyixc_ctx_rdata_29[5][34] , \_zyixc_ctx_rdata_29[5][33] , 
	\_zyixc_ctx_rdata_29[5][32] , \_zyixc_ctx_rdata_29[5][31] , 
	\_zyixc_ctx_rdata_29[5][30] , \_zyixc_ctx_rdata_29[5][29] , 
	\_zyixc_ctx_rdata_29[5][28] , \_zyixc_ctx_rdata_29[5][27] , 
	\_zyixc_ctx_rdata_29[5][26] , \_zyixc_ctx_rdata_29[5][25] , 
	\_zyixc_ctx_rdata_29[5][24] , \_zyixc_ctx_rdata_29[5][23] , 
	\_zyixc_ctx_rdata_29[5][22] , \_zyixc_ctx_rdata_29[5][21] , 
	\_zyixc_ctx_rdata_29[5][20] , \_zyixc_ctx_rdata_29[5][19] , 
	\_zyixc_ctx_rdata_29[5][18] , \_zyixc_ctx_rdata_29[5][17] , 
	\_zyixc_ctx_rdata_29[5][16] , \_zyixc_ctx_rdata_29[5][15] , 
	\_zyixc_ctx_rdata_29[5][14] , \_zyixc_ctx_rdata_29[5][13] , 
	\_zyixc_ctx_rdata_29[5][12] , \_zyixc_ctx_rdata_29[5][11] , 
	\_zyixc_ctx_rdata_29[5][10] , \_zyixc_ctx_rdata_29[5][9] , 
	\_zyixc_ctx_rdata_29[5][8] , \_zyixc_ctx_rdata_29[5][7] , 
	\_zyixc_ctx_rdata_29[5][6] , \_zyixc_ctx_rdata_29[5][5] , 
	\_zyixc_ctx_rdata_29[5][4] , \_zyixc_ctx_rdata_29[5][3] , 
	\_zyixc_ctx_rdata_29[5][2] , \_zyixc_ctx_rdata_29[5][1] , 
	\_zyixc_ctx_rdata_29[5][0] , \_zyixc_ctx_rdata_29[6][63] , 
	\_zyixc_ctx_rdata_29[6][62] , \_zyixc_ctx_rdata_29[6][61] , 
	\_zyixc_ctx_rdata_29[6][60] , \_zyixc_ctx_rdata_29[6][59] , 
	\_zyixc_ctx_rdata_29[6][58] , \_zyixc_ctx_rdata_29[6][57] , 
	\_zyixc_ctx_rdata_29[6][56] , \_zyixc_ctx_rdata_29[6][55] , 
	\_zyixc_ctx_rdata_29[6][54] , \_zyixc_ctx_rdata_29[6][53] , 
	\_zyixc_ctx_rdata_29[6][52] , \_zyixc_ctx_rdata_29[6][51] , 
	\_zyixc_ctx_rdata_29[6][50] , \_zyixc_ctx_rdata_29[6][49] , 
	\_zyixc_ctx_rdata_29[6][48] , \_zyixc_ctx_rdata_29[6][47] , 
	\_zyixc_ctx_rdata_29[6][46] , \_zyixc_ctx_rdata_29[6][45] , 
	\_zyixc_ctx_rdata_29[6][44] , \_zyixc_ctx_rdata_29[6][43] , 
	\_zyixc_ctx_rdata_29[6][42] , \_zyixc_ctx_rdata_29[6][41] , 
	\_zyixc_ctx_rdata_29[6][40] , \_zyixc_ctx_rdata_29[6][39] , 
	\_zyixc_ctx_rdata_29[6][38] , \_zyixc_ctx_rdata_29[6][37] , 
	\_zyixc_ctx_rdata_29[6][36] , \_zyixc_ctx_rdata_29[6][35] , 
	\_zyixc_ctx_rdata_29[6][34] , \_zyixc_ctx_rdata_29[6][33] , 
	\_zyixc_ctx_rdata_29[6][32] , \_zyixc_ctx_rdata_29[6][31] , 
	\_zyixc_ctx_rdata_29[6][30] , \_zyixc_ctx_rdata_29[6][29] , 
	\_zyixc_ctx_rdata_29[6][28] , \_zyixc_ctx_rdata_29[6][27] , 
	\_zyixc_ctx_rdata_29[6][26] , \_zyixc_ctx_rdata_29[6][25] , 
	\_zyixc_ctx_rdata_29[6][24] , \_zyixc_ctx_rdata_29[6][23] , 
	\_zyixc_ctx_rdata_29[6][22] , \_zyixc_ctx_rdata_29[6][21] , 
	\_zyixc_ctx_rdata_29[6][20] , \_zyixc_ctx_rdata_29[6][19] , 
	\_zyixc_ctx_rdata_29[6][18] , \_zyixc_ctx_rdata_29[6][17] , 
	\_zyixc_ctx_rdata_29[6][16] , \_zyixc_ctx_rdata_29[6][15] , 
	\_zyixc_ctx_rdata_29[6][14] , \_zyixc_ctx_rdata_29[6][13] , 
	\_zyixc_ctx_rdata_29[6][12] , \_zyixc_ctx_rdata_29[6][11] , 
	\_zyixc_ctx_rdata_29[6][10] , \_zyixc_ctx_rdata_29[6][9] , 
	\_zyixc_ctx_rdata_29[6][8] , \_zyixc_ctx_rdata_29[6][7] , 
	\_zyixc_ctx_rdata_29[6][6] , \_zyixc_ctx_rdata_29[6][5] , 
	\_zyixc_ctx_rdata_29[6][4] , \_zyixc_ctx_rdata_29[6][3] , 
	\_zyixc_ctx_rdata_29[6][2] , \_zyixc_ctx_rdata_29[6][1] , 
	\_zyixc_ctx_rdata_29[6][0] , \_zyixc_ctx_rdata_29[7][63] , 
	\_zyixc_ctx_rdata_29[7][62] , \_zyixc_ctx_rdata_29[7][61] , 
	\_zyixc_ctx_rdata_29[7][60] , \_zyixc_ctx_rdata_29[7][59] , 
	\_zyixc_ctx_rdata_29[7][58] , \_zyixc_ctx_rdata_29[7][57] , 
	\_zyixc_ctx_rdata_29[7][56] , \_zyixc_ctx_rdata_29[7][55] , 
	\_zyixc_ctx_rdata_29[7][54] , \_zyixc_ctx_rdata_29[7][53] , 
	\_zyixc_ctx_rdata_29[7][52] , \_zyixc_ctx_rdata_29[7][51] , 
	\_zyixc_ctx_rdata_29[7][50] , \_zyixc_ctx_rdata_29[7][49] , 
	\_zyixc_ctx_rdata_29[7][48] , \_zyixc_ctx_rdata_29[7][47] , 
	\_zyixc_ctx_rdata_29[7][46] , \_zyixc_ctx_rdata_29[7][45] , 
	\_zyixc_ctx_rdata_29[7][44] , \_zyixc_ctx_rdata_29[7][43] , 
	\_zyixc_ctx_rdata_29[7][42] , \_zyixc_ctx_rdata_29[7][41] , 
	\_zyixc_ctx_rdata_29[7][40] , \_zyixc_ctx_rdata_29[7][39] , 
	\_zyixc_ctx_rdata_29[7][38] , \_zyixc_ctx_rdata_29[7][37] , 
	\_zyixc_ctx_rdata_29[7][36] , \_zyixc_ctx_rdata_29[7][35] , 
	\_zyixc_ctx_rdata_29[7][34] , \_zyixc_ctx_rdata_29[7][33] , 
	\_zyixc_ctx_rdata_29[7][32] , \_zyixc_ctx_rdata_29[7][31] , 
	\_zyixc_ctx_rdata_29[7][30] , \_zyixc_ctx_rdata_29[7][29] , 
	\_zyixc_ctx_rdata_29[7][28] , \_zyixc_ctx_rdata_29[7][27] , 
	\_zyixc_ctx_rdata_29[7][26] , \_zyixc_ctx_rdata_29[7][25] , 
	\_zyixc_ctx_rdata_29[7][24] , \_zyixc_ctx_rdata_29[7][23] , 
	\_zyixc_ctx_rdata_29[7][22] , \_zyixc_ctx_rdata_29[7][21] , 
	\_zyixc_ctx_rdata_29[7][20] , \_zyixc_ctx_rdata_29[7][19] , 
	\_zyixc_ctx_rdata_29[7][18] , \_zyixc_ctx_rdata_29[7][17] , 
	\_zyixc_ctx_rdata_29[7][16] , \_zyixc_ctx_rdata_29[7][15] , 
	\_zyixc_ctx_rdata_29[7][14] , \_zyixc_ctx_rdata_29[7][13] , 
	\_zyixc_ctx_rdata_29[7][12] , \_zyixc_ctx_rdata_29[7][11] , 
	\_zyixc_ctx_rdata_29[7][10] , \_zyixc_ctx_rdata_29[7][9] , 
	\_zyixc_ctx_rdata_29[7][8] , \_zyixc_ctx_rdata_29[7][7] , 
	\_zyixc_ctx_rdata_29[7][6] , \_zyixc_ctx_rdata_29[7][5] , 
	\_zyixc_ctx_rdata_29[7][4] , \_zyixc_ctx_rdata_29[7][3] , 
	\_zyixc_ctx_rdata_29[7][2] , \_zyixc_ctx_rdata_29[7][1] , 
	\_zyixc_ctx_rdata_29[7][0] , \_zyixc_ctx_rdata_29[8][63] , 
	\_zyixc_ctx_rdata_29[8][62] , \_zyixc_ctx_rdata_29[8][61] , 
	\_zyixc_ctx_rdata_29[8][60] , \_zyixc_ctx_rdata_29[8][59] , 
	\_zyixc_ctx_rdata_29[8][58] , \_zyixc_ctx_rdata_29[8][57] , 
	\_zyixc_ctx_rdata_29[8][56] , \_zyixc_ctx_rdata_29[8][55] , 
	\_zyixc_ctx_rdata_29[8][54] , \_zyixc_ctx_rdata_29[8][53] , 
	\_zyixc_ctx_rdata_29[8][52] , \_zyixc_ctx_rdata_29[8][51] , 
	\_zyixc_ctx_rdata_29[8][50] , \_zyixc_ctx_rdata_29[8][49] , 
	\_zyixc_ctx_rdata_29[8][48] , \_zyixc_ctx_rdata_29[8][47] , 
	\_zyixc_ctx_rdata_29[8][46] , \_zyixc_ctx_rdata_29[8][45] , 
	\_zyixc_ctx_rdata_29[8][44] , \_zyixc_ctx_rdata_29[8][43] , 
	\_zyixc_ctx_rdata_29[8][42] , \_zyixc_ctx_rdata_29[8][41] , 
	\_zyixc_ctx_rdata_29[8][40] , \_zyixc_ctx_rdata_29[8][39] , 
	\_zyixc_ctx_rdata_29[8][38] , \_zyixc_ctx_rdata_29[8][37] , 
	\_zyixc_ctx_rdata_29[8][36] , \_zyixc_ctx_rdata_29[8][35] , 
	\_zyixc_ctx_rdata_29[8][34] , \_zyixc_ctx_rdata_29[8][33] , 
	\_zyixc_ctx_rdata_29[8][32] , \_zyixc_ctx_rdata_29[8][31] , 
	\_zyixc_ctx_rdata_29[8][30] , \_zyixc_ctx_rdata_29[8][29] , 
	\_zyixc_ctx_rdata_29[8][28] , \_zyixc_ctx_rdata_29[8][27] , 
	\_zyixc_ctx_rdata_29[8][26] , \_zyixc_ctx_rdata_29[8][25] , 
	\_zyixc_ctx_rdata_29[8][24] , \_zyixc_ctx_rdata_29[8][23] , 
	\_zyixc_ctx_rdata_29[8][22] , \_zyixc_ctx_rdata_29[8][21] , 
	\_zyixc_ctx_rdata_29[8][20] , \_zyixc_ctx_rdata_29[8][19] , 
	\_zyixc_ctx_rdata_29[8][18] , \_zyixc_ctx_rdata_29[8][17] , 
	\_zyixc_ctx_rdata_29[8][16] , \_zyixc_ctx_rdata_29[8][15] , 
	\_zyixc_ctx_rdata_29[8][14] , \_zyixc_ctx_rdata_29[8][13] , 
	\_zyixc_ctx_rdata_29[8][12] , \_zyixc_ctx_rdata_29[8][11] , 
	\_zyixc_ctx_rdata_29[8][10] , \_zyixc_ctx_rdata_29[8][9] , 
	\_zyixc_ctx_rdata_29[8][8] , \_zyixc_ctx_rdata_29[8][7] , 
	\_zyixc_ctx_rdata_29[8][6] , \_zyixc_ctx_rdata_29[8][5] , 
	\_zyixc_ctx_rdata_29[8][4] , \_zyixc_ctx_rdata_29[8][3] , 
	\_zyixc_ctx_rdata_29[8][2] , \_zyixc_ctx_rdata_29[8][1] , 
	\_zyixc_ctx_rdata_29[8][0] , \_zyixc_ctx_rdata_29[9][63] , 
	\_zyixc_ctx_rdata_29[9][62] , \_zyixc_ctx_rdata_29[9][61] , 
	\_zyixc_ctx_rdata_29[9][60] , \_zyixc_ctx_rdata_29[9][59] , 
	\_zyixc_ctx_rdata_29[9][58] , \_zyixc_ctx_rdata_29[9][57] , 
	\_zyixc_ctx_rdata_29[9][56] , \_zyixc_ctx_rdata_29[9][55] , 
	\_zyixc_ctx_rdata_29[9][54] , \_zyixc_ctx_rdata_29[9][53] , 
	\_zyixc_ctx_rdata_29[9][52] , \_zyixc_ctx_rdata_29[9][51] , 
	\_zyixc_ctx_rdata_29[9][50] , \_zyixc_ctx_rdata_29[9][49] , 
	\_zyixc_ctx_rdata_29[9][48] , \_zyixc_ctx_rdata_29[9][47] , 
	\_zyixc_ctx_rdata_29[9][46] , \_zyixc_ctx_rdata_29[9][45] , 
	\_zyixc_ctx_rdata_29[9][44] , \_zyixc_ctx_rdata_29[9][43] , 
	\_zyixc_ctx_rdata_29[9][42] , \_zyixc_ctx_rdata_29[9][41] , 
	\_zyixc_ctx_rdata_29[9][40] , \_zyixc_ctx_rdata_29[9][39] , 
	\_zyixc_ctx_rdata_29[9][38] , \_zyixc_ctx_rdata_29[9][37] , 
	\_zyixc_ctx_rdata_29[9][36] , \_zyixc_ctx_rdata_29[9][35] , 
	\_zyixc_ctx_rdata_29[9][34] , \_zyixc_ctx_rdata_29[9][33] , 
	\_zyixc_ctx_rdata_29[9][32] , \_zyixc_ctx_rdata_29[9][31] , 
	\_zyixc_ctx_rdata_29[9][30] , \_zyixc_ctx_rdata_29[9][29] , 
	\_zyixc_ctx_rdata_29[9][28] , \_zyixc_ctx_rdata_29[9][27] , 
	\_zyixc_ctx_rdata_29[9][26] , \_zyixc_ctx_rdata_29[9][25] , 
	\_zyixc_ctx_rdata_29[9][24] , \_zyixc_ctx_rdata_29[9][23] , 
	\_zyixc_ctx_rdata_29[9][22] , \_zyixc_ctx_rdata_29[9][21] , 
	\_zyixc_ctx_rdata_29[9][20] , \_zyixc_ctx_rdata_29[9][19] , 
	\_zyixc_ctx_rdata_29[9][18] , \_zyixc_ctx_rdata_29[9][17] , 
	\_zyixc_ctx_rdata_29[9][16] , \_zyixc_ctx_rdata_29[9][15] , 
	\_zyixc_ctx_rdata_29[9][14] , \_zyixc_ctx_rdata_29[9][13] , 
	\_zyixc_ctx_rdata_29[9][12] , \_zyixc_ctx_rdata_29[9][11] , 
	\_zyixc_ctx_rdata_29[9][10] , \_zyixc_ctx_rdata_29[9][9] , 
	\_zyixc_ctx_rdata_29[9][8] , \_zyixc_ctx_rdata_29[9][7] , 
	\_zyixc_ctx_rdata_29[9][6] , \_zyixc_ctx_rdata_29[9][5] , 
	\_zyixc_ctx_rdata_29[9][4] , \_zyixc_ctx_rdata_29[9][3] , 
	\_zyixc_ctx_rdata_29[9][2] , \_zyixc_ctx_rdata_29[9][1] , 
	\_zyixc_ctx_rdata_29[9][0] , \_zyixc_ctx_rdata_29[10][63] , 
	\_zyixc_ctx_rdata_29[10][62] , \_zyixc_ctx_rdata_29[10][61] , 
	\_zyixc_ctx_rdata_29[10][60] , \_zyixc_ctx_rdata_29[10][59] , 
	\_zyixc_ctx_rdata_29[10][58] , \_zyixc_ctx_rdata_29[10][57] , 
	\_zyixc_ctx_rdata_29[10][56] , \_zyixc_ctx_rdata_29[10][55] , 
	\_zyixc_ctx_rdata_29[10][54] , \_zyixc_ctx_rdata_29[10][53] , 
	\_zyixc_ctx_rdata_29[10][52] , \_zyixc_ctx_rdata_29[10][51] , 
	\_zyixc_ctx_rdata_29[10][50] , \_zyixc_ctx_rdata_29[10][49] , 
	\_zyixc_ctx_rdata_29[10][48] , \_zyixc_ctx_rdata_29[10][47] , 
	\_zyixc_ctx_rdata_29[10][46] , \_zyixc_ctx_rdata_29[10][45] , 
	\_zyixc_ctx_rdata_29[10][44] , \_zyixc_ctx_rdata_29[10][43] , 
	\_zyixc_ctx_rdata_29[10][42] , \_zyixc_ctx_rdata_29[10][41] , 
	\_zyixc_ctx_rdata_29[10][40] , \_zyixc_ctx_rdata_29[10][39] , 
	\_zyixc_ctx_rdata_29[10][38] , \_zyixc_ctx_rdata_29[10][37] , 
	\_zyixc_ctx_rdata_29[10][36] , \_zyixc_ctx_rdata_29[10][35] , 
	\_zyixc_ctx_rdata_29[10][34] , \_zyixc_ctx_rdata_29[10][33] , 
	\_zyixc_ctx_rdata_29[10][32] , \_zyixc_ctx_rdata_29[10][31] , 
	\_zyixc_ctx_rdata_29[10][30] , \_zyixc_ctx_rdata_29[10][29] , 
	\_zyixc_ctx_rdata_29[10][28] , \_zyixc_ctx_rdata_29[10][27] , 
	\_zyixc_ctx_rdata_29[10][26] , \_zyixc_ctx_rdata_29[10][25] , 
	\_zyixc_ctx_rdata_29[10][24] , \_zyixc_ctx_rdata_29[10][23] , 
	\_zyixc_ctx_rdata_29[10][22] , \_zyixc_ctx_rdata_29[10][21] , 
	\_zyixc_ctx_rdata_29[10][20] , \_zyixc_ctx_rdata_29[10][19] , 
	\_zyixc_ctx_rdata_29[10][18] , \_zyixc_ctx_rdata_29[10][17] , 
	\_zyixc_ctx_rdata_29[10][16] , \_zyixc_ctx_rdata_29[10][15] , 
	\_zyixc_ctx_rdata_29[10][14] , \_zyixc_ctx_rdata_29[10][13] , 
	\_zyixc_ctx_rdata_29[10][12] , \_zyixc_ctx_rdata_29[10][11] , 
	\_zyixc_ctx_rdata_29[10][10] , \_zyixc_ctx_rdata_29[10][9] , 
	\_zyixc_ctx_rdata_29[10][8] , \_zyixc_ctx_rdata_29[10][7] , 
	\_zyixc_ctx_rdata_29[10][6] , \_zyixc_ctx_rdata_29[10][5] , 
	\_zyixc_ctx_rdata_29[10][4] , \_zyixc_ctx_rdata_29[10][3] , 
	\_zyixc_ctx_rdata_29[10][2] , \_zyixc_ctx_rdata_29[10][1] , 
	\_zyixc_ctx_rdata_29[10][0] , \_zyixc_ctx_rdata_29[11][63] , 
	\_zyixc_ctx_rdata_29[11][62] , \_zyixc_ctx_rdata_29[11][61] , 
	\_zyixc_ctx_rdata_29[11][60] , \_zyixc_ctx_rdata_29[11][59] , 
	\_zyixc_ctx_rdata_29[11][58] , \_zyixc_ctx_rdata_29[11][57] , 
	\_zyixc_ctx_rdata_29[11][56] , \_zyixc_ctx_rdata_29[11][55] , 
	\_zyixc_ctx_rdata_29[11][54] , \_zyixc_ctx_rdata_29[11][53] , 
	\_zyixc_ctx_rdata_29[11][52] , \_zyixc_ctx_rdata_29[11][51] , 
	\_zyixc_ctx_rdata_29[11][50] , \_zyixc_ctx_rdata_29[11][49] , 
	\_zyixc_ctx_rdata_29[11][48] , \_zyixc_ctx_rdata_29[11][47] , 
	\_zyixc_ctx_rdata_29[11][46] , \_zyixc_ctx_rdata_29[11][45] , 
	\_zyixc_ctx_rdata_29[11][44] , \_zyixc_ctx_rdata_29[11][43] , 
	\_zyixc_ctx_rdata_29[11][42] , \_zyixc_ctx_rdata_29[11][41] , 
	\_zyixc_ctx_rdata_29[11][40] , \_zyixc_ctx_rdata_29[11][39] , 
	\_zyixc_ctx_rdata_29[11][38] , \_zyixc_ctx_rdata_29[11][37] , 
	\_zyixc_ctx_rdata_29[11][36] , \_zyixc_ctx_rdata_29[11][35] , 
	\_zyixc_ctx_rdata_29[11][34] , \_zyixc_ctx_rdata_29[11][33] , 
	\_zyixc_ctx_rdata_29[11][32] , \_zyixc_ctx_rdata_29[11][31] , 
	\_zyixc_ctx_rdata_29[11][30] , \_zyixc_ctx_rdata_29[11][29] , 
	\_zyixc_ctx_rdata_29[11][28] , \_zyixc_ctx_rdata_29[11][27] , 
	\_zyixc_ctx_rdata_29[11][26] , \_zyixc_ctx_rdata_29[11][25] , 
	\_zyixc_ctx_rdata_29[11][24] , \_zyixc_ctx_rdata_29[11][23] , 
	\_zyixc_ctx_rdata_29[11][22] , \_zyixc_ctx_rdata_29[11][21] , 
	\_zyixc_ctx_rdata_29[11][20] , \_zyixc_ctx_rdata_29[11][19] , 
	\_zyixc_ctx_rdata_29[11][18] , \_zyixc_ctx_rdata_29[11][17] , 
	\_zyixc_ctx_rdata_29[11][16] , \_zyixc_ctx_rdata_29[11][15] , 
	\_zyixc_ctx_rdata_29[11][14] , \_zyixc_ctx_rdata_29[11][13] , 
	\_zyixc_ctx_rdata_29[11][12] , \_zyixc_ctx_rdata_29[11][11] , 
	\_zyixc_ctx_rdata_29[11][10] , \_zyixc_ctx_rdata_29[11][9] , 
	\_zyixc_ctx_rdata_29[11][8] , \_zyixc_ctx_rdata_29[11][7] , 
	\_zyixc_ctx_rdata_29[11][6] , \_zyixc_ctx_rdata_29[11][5] , 
	\_zyixc_ctx_rdata_29[11][4] , \_zyixc_ctx_rdata_29[11][3] , 
	\_zyixc_ctx_rdata_29[11][2] , \_zyixc_ctx_rdata_29[11][1] , 
	\_zyixc_ctx_rdata_29[11][0] , \_zyixc_ctx_rdata_29[12][63] , 
	\_zyixc_ctx_rdata_29[12][62] , \_zyixc_ctx_rdata_29[12][61] , 
	\_zyixc_ctx_rdata_29[12][60] , \_zyixc_ctx_rdata_29[12][59] , 
	\_zyixc_ctx_rdata_29[12][58] , \_zyixc_ctx_rdata_29[12][57] , 
	\_zyixc_ctx_rdata_29[12][56] , \_zyixc_ctx_rdata_29[12][55] , 
	\_zyixc_ctx_rdata_29[12][54] , \_zyixc_ctx_rdata_29[12][53] , 
	\_zyixc_ctx_rdata_29[12][52] , \_zyixc_ctx_rdata_29[12][51] , 
	\_zyixc_ctx_rdata_29[12][50] , \_zyixc_ctx_rdata_29[12][49] , 
	\_zyixc_ctx_rdata_29[12][48] , \_zyixc_ctx_rdata_29[12][47] , 
	\_zyixc_ctx_rdata_29[12][46] , \_zyixc_ctx_rdata_29[12][45] , 
	\_zyixc_ctx_rdata_29[12][44] , \_zyixc_ctx_rdata_29[12][43] , 
	\_zyixc_ctx_rdata_29[12][42] , \_zyixc_ctx_rdata_29[12][41] , 
	\_zyixc_ctx_rdata_29[12][40] , \_zyixc_ctx_rdata_29[12][39] , 
	\_zyixc_ctx_rdata_29[12][38] , \_zyixc_ctx_rdata_29[12][37] , 
	\_zyixc_ctx_rdata_29[12][36] , \_zyixc_ctx_rdata_29[12][35] , 
	\_zyixc_ctx_rdata_29[12][34] , \_zyixc_ctx_rdata_29[12][33] , 
	\_zyixc_ctx_rdata_29[12][32] , \_zyixc_ctx_rdata_29[12][31] , 
	\_zyixc_ctx_rdata_29[12][30] , \_zyixc_ctx_rdata_29[12][29] , 
	\_zyixc_ctx_rdata_29[12][28] , \_zyixc_ctx_rdata_29[12][27] , 
	\_zyixc_ctx_rdata_29[12][26] , \_zyixc_ctx_rdata_29[12][25] , 
	\_zyixc_ctx_rdata_29[12][24] , \_zyixc_ctx_rdata_29[12][23] , 
	\_zyixc_ctx_rdata_29[12][22] , \_zyixc_ctx_rdata_29[12][21] , 
	\_zyixc_ctx_rdata_29[12][20] , \_zyixc_ctx_rdata_29[12][19] , 
	\_zyixc_ctx_rdata_29[12][18] , \_zyixc_ctx_rdata_29[12][17] , 
	\_zyixc_ctx_rdata_29[12][16] , \_zyixc_ctx_rdata_29[12][15] , 
	\_zyixc_ctx_rdata_29[12][14] , \_zyixc_ctx_rdata_29[12][13] , 
	\_zyixc_ctx_rdata_29[12][12] , \_zyixc_ctx_rdata_29[12][11] , 
	\_zyixc_ctx_rdata_29[12][10] , \_zyixc_ctx_rdata_29[12][9] , 
	\_zyixc_ctx_rdata_29[12][8] , \_zyixc_ctx_rdata_29[12][7] , 
	\_zyixc_ctx_rdata_29[12][6] , \_zyixc_ctx_rdata_29[12][5] , 
	\_zyixc_ctx_rdata_29[12][4] , \_zyixc_ctx_rdata_29[12][3] , 
	\_zyixc_ctx_rdata_29[12][2] , \_zyixc_ctx_rdata_29[12][1] , 
	\_zyixc_ctx_rdata_29[12][0] , \_zyixc_ctx_rdata_29[13][63] , 
	\_zyixc_ctx_rdata_29[13][62] , \_zyixc_ctx_rdata_29[13][61] , 
	\_zyixc_ctx_rdata_29[13][60] , \_zyixc_ctx_rdata_29[13][59] , 
	\_zyixc_ctx_rdata_29[13][58] , \_zyixc_ctx_rdata_29[13][57] , 
	\_zyixc_ctx_rdata_29[13][56] , \_zyixc_ctx_rdata_29[13][55] , 
	\_zyixc_ctx_rdata_29[13][54] , \_zyixc_ctx_rdata_29[13][53] , 
	\_zyixc_ctx_rdata_29[13][52] , \_zyixc_ctx_rdata_29[13][51] , 
	\_zyixc_ctx_rdata_29[13][50] , \_zyixc_ctx_rdata_29[13][49] , 
	\_zyixc_ctx_rdata_29[13][48] , \_zyixc_ctx_rdata_29[13][47] , 
	\_zyixc_ctx_rdata_29[13][46] , \_zyixc_ctx_rdata_29[13][45] , 
	\_zyixc_ctx_rdata_29[13][44] , \_zyixc_ctx_rdata_29[13][43] , 
	\_zyixc_ctx_rdata_29[13][42] , \_zyixc_ctx_rdata_29[13][41] , 
	\_zyixc_ctx_rdata_29[13][40] , \_zyixc_ctx_rdata_29[13][39] , 
	\_zyixc_ctx_rdata_29[13][38] , \_zyixc_ctx_rdata_29[13][37] , 
	\_zyixc_ctx_rdata_29[13][36] , \_zyixc_ctx_rdata_29[13][35] , 
	\_zyixc_ctx_rdata_29[13][34] , \_zyixc_ctx_rdata_29[13][33] , 
	\_zyixc_ctx_rdata_29[13][32] , \_zyixc_ctx_rdata_29[13][31] , 
	\_zyixc_ctx_rdata_29[13][30] , \_zyixc_ctx_rdata_29[13][29] , 
	\_zyixc_ctx_rdata_29[13][28] , \_zyixc_ctx_rdata_29[13][27] , 
	\_zyixc_ctx_rdata_29[13][26] , \_zyixc_ctx_rdata_29[13][25] , 
	\_zyixc_ctx_rdata_29[13][24] , \_zyixc_ctx_rdata_29[13][23] , 
	\_zyixc_ctx_rdata_29[13][22] , \_zyixc_ctx_rdata_29[13][21] , 
	\_zyixc_ctx_rdata_29[13][20] , \_zyixc_ctx_rdata_29[13][19] , 
	\_zyixc_ctx_rdata_29[13][18] , \_zyixc_ctx_rdata_29[13][17] , 
	\_zyixc_ctx_rdata_29[13][16] , \_zyixc_ctx_rdata_29[13][15] , 
	\_zyixc_ctx_rdata_29[13][14] , \_zyixc_ctx_rdata_29[13][13] , 
	\_zyixc_ctx_rdata_29[13][12] , \_zyixc_ctx_rdata_29[13][11] , 
	\_zyixc_ctx_rdata_29[13][10] , \_zyixc_ctx_rdata_29[13][9] , 
	\_zyixc_ctx_rdata_29[13][8] , \_zyixc_ctx_rdata_29[13][7] , 
	\_zyixc_ctx_rdata_29[13][6] , \_zyixc_ctx_rdata_29[13][5] , 
	\_zyixc_ctx_rdata_29[13][4] , \_zyixc_ctx_rdata_29[13][3] , 
	\_zyixc_ctx_rdata_29[13][2] , \_zyixc_ctx_rdata_29[13][1] , 
	\_zyixc_ctx_rdata_29[13][0] , \_zyixc_ctx_rdata_29[14][63] , 
	\_zyixc_ctx_rdata_29[14][62] , \_zyixc_ctx_rdata_29[14][61] , 
	\_zyixc_ctx_rdata_29[14][60] , \_zyixc_ctx_rdata_29[14][59] , 
	\_zyixc_ctx_rdata_29[14][58] , \_zyixc_ctx_rdata_29[14][57] , 
	\_zyixc_ctx_rdata_29[14][56] , \_zyixc_ctx_rdata_29[14][55] , 
	\_zyixc_ctx_rdata_29[14][54] , \_zyixc_ctx_rdata_29[14][53] , 
	\_zyixc_ctx_rdata_29[14][52] , \_zyixc_ctx_rdata_29[14][51] , 
	\_zyixc_ctx_rdata_29[14][50] , \_zyixc_ctx_rdata_29[14][49] , 
	\_zyixc_ctx_rdata_29[14][48] , \_zyixc_ctx_rdata_29[14][47] , 
	\_zyixc_ctx_rdata_29[14][46] , \_zyixc_ctx_rdata_29[14][45] , 
	\_zyixc_ctx_rdata_29[14][44] , \_zyixc_ctx_rdata_29[14][43] , 
	\_zyixc_ctx_rdata_29[14][42] , \_zyixc_ctx_rdata_29[14][41] , 
	\_zyixc_ctx_rdata_29[14][40] , \_zyixc_ctx_rdata_29[14][39] , 
	\_zyixc_ctx_rdata_29[14][38] , \_zyixc_ctx_rdata_29[14][37] , 
	\_zyixc_ctx_rdata_29[14][36] , \_zyixc_ctx_rdata_29[14][35] , 
	\_zyixc_ctx_rdata_29[14][34] , \_zyixc_ctx_rdata_29[14][33] , 
	\_zyixc_ctx_rdata_29[14][32] , \_zyixc_ctx_rdata_29[14][31] , 
	\_zyixc_ctx_rdata_29[14][30] , \_zyixc_ctx_rdata_29[14][29] , 
	\_zyixc_ctx_rdata_29[14][28] , \_zyixc_ctx_rdata_29[14][27] , 
	\_zyixc_ctx_rdata_29[14][26] , \_zyixc_ctx_rdata_29[14][25] , 
	\_zyixc_ctx_rdata_29[14][24] , \_zyixc_ctx_rdata_29[14][23] , 
	\_zyixc_ctx_rdata_29[14][22] , \_zyixc_ctx_rdata_29[14][21] , 
	\_zyixc_ctx_rdata_29[14][20] , \_zyixc_ctx_rdata_29[14][19] , 
	\_zyixc_ctx_rdata_29[14][18] , \_zyixc_ctx_rdata_29[14][17] , 
	\_zyixc_ctx_rdata_29[14][16] , \_zyixc_ctx_rdata_29[14][15] , 
	\_zyixc_ctx_rdata_29[14][14] , \_zyixc_ctx_rdata_29[14][13] , 
	\_zyixc_ctx_rdata_29[14][12] , \_zyixc_ctx_rdata_29[14][11] , 
	\_zyixc_ctx_rdata_29[14][10] , \_zyixc_ctx_rdata_29[14][9] , 
	\_zyixc_ctx_rdata_29[14][8] , \_zyixc_ctx_rdata_29[14][7] , 
	\_zyixc_ctx_rdata_29[14][6] , \_zyixc_ctx_rdata_29[14][5] , 
	\_zyixc_ctx_rdata_29[14][4] , \_zyixc_ctx_rdata_29[14][3] , 
	\_zyixc_ctx_rdata_29[14][2] , \_zyixc_ctx_rdata_29[14][1] , 
	\_zyixc_ctx_rdata_29[14][0] , \_zyixc_ctx_rdata_29[15][63] , 
	\_zyixc_ctx_rdata_29[15][62] , \_zyixc_ctx_rdata_29[15][61] , 
	\_zyixc_ctx_rdata_29[15][60] , \_zyixc_ctx_rdata_29[15][59] , 
	\_zyixc_ctx_rdata_29[15][58] , \_zyixc_ctx_rdata_29[15][57] , 
	\_zyixc_ctx_rdata_29[15][56] , \_zyixc_ctx_rdata_29[15][55] , 
	\_zyixc_ctx_rdata_29[15][54] , \_zyixc_ctx_rdata_29[15][53] , 
	\_zyixc_ctx_rdata_29[15][52] , \_zyixc_ctx_rdata_29[15][51] , 
	\_zyixc_ctx_rdata_29[15][50] , \_zyixc_ctx_rdata_29[15][49] , 
	\_zyixc_ctx_rdata_29[15][48] , \_zyixc_ctx_rdata_29[15][47] , 
	\_zyixc_ctx_rdata_29[15][46] , \_zyixc_ctx_rdata_29[15][45] , 
	\_zyixc_ctx_rdata_29[15][44] , \_zyixc_ctx_rdata_29[15][43] , 
	\_zyixc_ctx_rdata_29[15][42] , \_zyixc_ctx_rdata_29[15][41] , 
	\_zyixc_ctx_rdata_29[15][40] , \_zyixc_ctx_rdata_29[15][39] , 
	\_zyixc_ctx_rdata_29[15][38] , \_zyixc_ctx_rdata_29[15][37] , 
	\_zyixc_ctx_rdata_29[15][36] , \_zyixc_ctx_rdata_29[15][35] , 
	\_zyixc_ctx_rdata_29[15][34] , \_zyixc_ctx_rdata_29[15][33] , 
	\_zyixc_ctx_rdata_29[15][32] , \_zyixc_ctx_rdata_29[15][31] , 
	\_zyixc_ctx_rdata_29[15][30] , \_zyixc_ctx_rdata_29[15][29] , 
	\_zyixc_ctx_rdata_29[15][28] , \_zyixc_ctx_rdata_29[15][27] , 
	\_zyixc_ctx_rdata_29[15][26] , \_zyixc_ctx_rdata_29[15][25] , 
	\_zyixc_ctx_rdata_29[15][24] , \_zyixc_ctx_rdata_29[15][23] , 
	\_zyixc_ctx_rdata_29[15][22] , \_zyixc_ctx_rdata_29[15][21] , 
	\_zyixc_ctx_rdata_29[15][20] , \_zyixc_ctx_rdata_29[15][19] , 
	\_zyixc_ctx_rdata_29[15][18] , \_zyixc_ctx_rdata_29[15][17] , 
	\_zyixc_ctx_rdata_29[15][16] , \_zyixc_ctx_rdata_29[15][15] , 
	\_zyixc_ctx_rdata_29[15][14] , \_zyixc_ctx_rdata_29[15][13] , 
	\_zyixc_ctx_rdata_29[15][12] , \_zyixc_ctx_rdata_29[15][11] , 
	\_zyixc_ctx_rdata_29[15][10] , \_zyixc_ctx_rdata_29[15][9] , 
	\_zyixc_ctx_rdata_29[15][8] , \_zyixc_ctx_rdata_29[15][7] , 
	\_zyixc_ctx_rdata_29[15][6] , \_zyixc_ctx_rdata_29[15][5] , 
	\_zyixc_ctx_rdata_29[15][4] , \_zyixc_ctx_rdata_29[15][3] , 
	\_zyixc_ctx_rdata_29[15][2] , \_zyixc_ctx_rdata_29[15][1] , 
	\_zyixc_ctx_rdata_29[15][0] , \_zyixc_ctx_rdata_29[16][63] , 
	\_zyixc_ctx_rdata_29[16][62] , \_zyixc_ctx_rdata_29[16][61] , 
	\_zyixc_ctx_rdata_29[16][60] , \_zyixc_ctx_rdata_29[16][59] , 
	\_zyixc_ctx_rdata_29[16][58] , \_zyixc_ctx_rdata_29[16][57] , 
	\_zyixc_ctx_rdata_29[16][56] , \_zyixc_ctx_rdata_29[16][55] , 
	\_zyixc_ctx_rdata_29[16][54] , \_zyixc_ctx_rdata_29[16][53] , 
	\_zyixc_ctx_rdata_29[16][52] , \_zyixc_ctx_rdata_29[16][51] , 
	\_zyixc_ctx_rdata_29[16][50] , \_zyixc_ctx_rdata_29[16][49] , 
	\_zyixc_ctx_rdata_29[16][48] , \_zyixc_ctx_rdata_29[16][47] , 
	\_zyixc_ctx_rdata_29[16][46] , \_zyixc_ctx_rdata_29[16][45] , 
	\_zyixc_ctx_rdata_29[16][44] , \_zyixc_ctx_rdata_29[16][43] , 
	\_zyixc_ctx_rdata_29[16][42] , \_zyixc_ctx_rdata_29[16][41] , 
	\_zyixc_ctx_rdata_29[16][40] , \_zyixc_ctx_rdata_29[16][39] , 
	\_zyixc_ctx_rdata_29[16][38] , \_zyixc_ctx_rdata_29[16][37] , 
	\_zyixc_ctx_rdata_29[16][36] , \_zyixc_ctx_rdata_29[16][35] , 
	\_zyixc_ctx_rdata_29[16][34] , \_zyixc_ctx_rdata_29[16][33] , 
	\_zyixc_ctx_rdata_29[16][32] , \_zyixc_ctx_rdata_29[16][31] , 
	\_zyixc_ctx_rdata_29[16][30] , \_zyixc_ctx_rdata_29[16][29] , 
	\_zyixc_ctx_rdata_29[16][28] , \_zyixc_ctx_rdata_29[16][27] , 
	\_zyixc_ctx_rdata_29[16][26] , \_zyixc_ctx_rdata_29[16][25] , 
	\_zyixc_ctx_rdata_29[16][24] , \_zyixc_ctx_rdata_29[16][23] , 
	\_zyixc_ctx_rdata_29[16][22] , \_zyixc_ctx_rdata_29[16][21] , 
	\_zyixc_ctx_rdata_29[16][20] , \_zyixc_ctx_rdata_29[16][19] , 
	\_zyixc_ctx_rdata_29[16][18] , \_zyixc_ctx_rdata_29[16][17] , 
	\_zyixc_ctx_rdata_29[16][16] , \_zyixc_ctx_rdata_29[16][15] , 
	\_zyixc_ctx_rdata_29[16][14] , \_zyixc_ctx_rdata_29[16][13] , 
	\_zyixc_ctx_rdata_29[16][12] , \_zyixc_ctx_rdata_29[16][11] , 
	\_zyixc_ctx_rdata_29[16][10] , \_zyixc_ctx_rdata_29[16][9] , 
	\_zyixc_ctx_rdata_29[16][8] , \_zyixc_ctx_rdata_29[16][7] , 
	\_zyixc_ctx_rdata_29[16][6] , \_zyixc_ctx_rdata_29[16][5] , 
	\_zyixc_ctx_rdata_29[16][4] , \_zyixc_ctx_rdata_29[16][3] , 
	\_zyixc_ctx_rdata_29[16][2] , \_zyixc_ctx_rdata_29[16][1] , 
	\_zyixc_ctx_rdata_29[16][0] , \_zyixc_ctx_rdata_29[17][63] , 
	\_zyixc_ctx_rdata_29[17][62] , \_zyixc_ctx_rdata_29[17][61] , 
	\_zyixc_ctx_rdata_29[17][60] , \_zyixc_ctx_rdata_29[17][59] , 
	\_zyixc_ctx_rdata_29[17][58] , \_zyixc_ctx_rdata_29[17][57] , 
	\_zyixc_ctx_rdata_29[17][56] , \_zyixc_ctx_rdata_29[17][55] , 
	\_zyixc_ctx_rdata_29[17][54] , \_zyixc_ctx_rdata_29[17][53] , 
	\_zyixc_ctx_rdata_29[17][52] , \_zyixc_ctx_rdata_29[17][51] , 
	\_zyixc_ctx_rdata_29[17][50] , \_zyixc_ctx_rdata_29[17][49] , 
	\_zyixc_ctx_rdata_29[17][48] , \_zyixc_ctx_rdata_29[17][47] , 
	\_zyixc_ctx_rdata_29[17][46] , \_zyixc_ctx_rdata_29[17][45] , 
	\_zyixc_ctx_rdata_29[17][44] , \_zyixc_ctx_rdata_29[17][43] , 
	\_zyixc_ctx_rdata_29[17][42] , \_zyixc_ctx_rdata_29[17][41] , 
	\_zyixc_ctx_rdata_29[17][40] , \_zyixc_ctx_rdata_29[17][39] , 
	\_zyixc_ctx_rdata_29[17][38] , \_zyixc_ctx_rdata_29[17][37] , 
	\_zyixc_ctx_rdata_29[17][36] , \_zyixc_ctx_rdata_29[17][35] , 
	\_zyixc_ctx_rdata_29[17][34] , \_zyixc_ctx_rdata_29[17][33] , 
	\_zyixc_ctx_rdata_29[17][32] , \_zyixc_ctx_rdata_29[17][31] , 
	\_zyixc_ctx_rdata_29[17][30] , \_zyixc_ctx_rdata_29[17][29] , 
	\_zyixc_ctx_rdata_29[17][28] , \_zyixc_ctx_rdata_29[17][27] , 
	\_zyixc_ctx_rdata_29[17][26] , \_zyixc_ctx_rdata_29[17][25] , 
	\_zyixc_ctx_rdata_29[17][24] , \_zyixc_ctx_rdata_29[17][23] , 
	\_zyixc_ctx_rdata_29[17][22] , \_zyixc_ctx_rdata_29[17][21] , 
	\_zyixc_ctx_rdata_29[17][20] , \_zyixc_ctx_rdata_29[17][19] , 
	\_zyixc_ctx_rdata_29[17][18] , \_zyixc_ctx_rdata_29[17][17] , 
	\_zyixc_ctx_rdata_29[17][16] , \_zyixc_ctx_rdata_29[17][15] , 
	\_zyixc_ctx_rdata_29[17][14] , \_zyixc_ctx_rdata_29[17][13] , 
	\_zyixc_ctx_rdata_29[17][12] , \_zyixc_ctx_rdata_29[17][11] , 
	\_zyixc_ctx_rdata_29[17][10] , \_zyixc_ctx_rdata_29[17][9] , 
	\_zyixc_ctx_rdata_29[17][8] , \_zyixc_ctx_rdata_29[17][7] , 
	\_zyixc_ctx_rdata_29[17][6] , \_zyixc_ctx_rdata_29[17][5] , 
	\_zyixc_ctx_rdata_29[17][4] , \_zyixc_ctx_rdata_29[17][3] , 
	\_zyixc_ctx_rdata_29[17][2] , \_zyixc_ctx_rdata_29[17][1] , 
	\_zyixc_ctx_rdata_29[17][0] , \_zyixc_ctx_rdata_29[18][63] , 
	\_zyixc_ctx_rdata_29[18][62] , \_zyixc_ctx_rdata_29[18][61] , 
	\_zyixc_ctx_rdata_29[18][60] , \_zyixc_ctx_rdata_29[18][59] , 
	\_zyixc_ctx_rdata_29[18][58] , \_zyixc_ctx_rdata_29[18][57] , 
	\_zyixc_ctx_rdata_29[18][56] , \_zyixc_ctx_rdata_29[18][55] , 
	\_zyixc_ctx_rdata_29[18][54] , \_zyixc_ctx_rdata_29[18][53] , 
	\_zyixc_ctx_rdata_29[18][52] , \_zyixc_ctx_rdata_29[18][51] , 
	\_zyixc_ctx_rdata_29[18][50] , \_zyixc_ctx_rdata_29[18][49] , 
	\_zyixc_ctx_rdata_29[18][48] , \_zyixc_ctx_rdata_29[18][47] , 
	\_zyixc_ctx_rdata_29[18][46] , \_zyixc_ctx_rdata_29[18][45] , 
	\_zyixc_ctx_rdata_29[18][44] , \_zyixc_ctx_rdata_29[18][43] , 
	\_zyixc_ctx_rdata_29[18][42] , \_zyixc_ctx_rdata_29[18][41] , 
	\_zyixc_ctx_rdata_29[18][40] , \_zyixc_ctx_rdata_29[18][39] , 
	\_zyixc_ctx_rdata_29[18][38] , \_zyixc_ctx_rdata_29[18][37] , 
	\_zyixc_ctx_rdata_29[18][36] , \_zyixc_ctx_rdata_29[18][35] , 
	\_zyixc_ctx_rdata_29[18][34] , \_zyixc_ctx_rdata_29[18][33] , 
	\_zyixc_ctx_rdata_29[18][32] , \_zyixc_ctx_rdata_29[18][31] , 
	\_zyixc_ctx_rdata_29[18][30] , \_zyixc_ctx_rdata_29[18][29] , 
	\_zyixc_ctx_rdata_29[18][28] , \_zyixc_ctx_rdata_29[18][27] , 
	\_zyixc_ctx_rdata_29[18][26] , \_zyixc_ctx_rdata_29[18][25] , 
	\_zyixc_ctx_rdata_29[18][24] , \_zyixc_ctx_rdata_29[18][23] , 
	\_zyixc_ctx_rdata_29[18][22] , \_zyixc_ctx_rdata_29[18][21] , 
	\_zyixc_ctx_rdata_29[18][20] , \_zyixc_ctx_rdata_29[18][19] , 
	\_zyixc_ctx_rdata_29[18][18] , \_zyixc_ctx_rdata_29[18][17] , 
	\_zyixc_ctx_rdata_29[18][16] , \_zyixc_ctx_rdata_29[18][15] , 
	\_zyixc_ctx_rdata_29[18][14] , \_zyixc_ctx_rdata_29[18][13] , 
	\_zyixc_ctx_rdata_29[18][12] , \_zyixc_ctx_rdata_29[18][11] , 
	\_zyixc_ctx_rdata_29[18][10] , \_zyixc_ctx_rdata_29[18][9] , 
	\_zyixc_ctx_rdata_29[18][8] , \_zyixc_ctx_rdata_29[18][7] , 
	\_zyixc_ctx_rdata_29[18][6] , \_zyixc_ctx_rdata_29[18][5] , 
	\_zyixc_ctx_rdata_29[18][4] , \_zyixc_ctx_rdata_29[18][3] , 
	\_zyixc_ctx_rdata_29[18][2] , \_zyixc_ctx_rdata_29[18][1] , 
	\_zyixc_ctx_rdata_29[18][0] , \_zyixc_ctx_rdata_29[19][63] , 
	\_zyixc_ctx_rdata_29[19][62] , \_zyixc_ctx_rdata_29[19][61] , 
	\_zyixc_ctx_rdata_29[19][60] , \_zyixc_ctx_rdata_29[19][59] , 
	\_zyixc_ctx_rdata_29[19][58] , \_zyixc_ctx_rdata_29[19][57] , 
	\_zyixc_ctx_rdata_29[19][56] , \_zyixc_ctx_rdata_29[19][55] , 
	\_zyixc_ctx_rdata_29[19][54] , \_zyixc_ctx_rdata_29[19][53] , 
	\_zyixc_ctx_rdata_29[19][52] , \_zyixc_ctx_rdata_29[19][51] , 
	\_zyixc_ctx_rdata_29[19][50] , \_zyixc_ctx_rdata_29[19][49] , 
	\_zyixc_ctx_rdata_29[19][48] , \_zyixc_ctx_rdata_29[19][47] , 
	\_zyixc_ctx_rdata_29[19][46] , \_zyixc_ctx_rdata_29[19][45] , 
	\_zyixc_ctx_rdata_29[19][44] , \_zyixc_ctx_rdata_29[19][43] , 
	\_zyixc_ctx_rdata_29[19][42] , \_zyixc_ctx_rdata_29[19][41] , 
	\_zyixc_ctx_rdata_29[19][40] , \_zyixc_ctx_rdata_29[19][39] , 
	\_zyixc_ctx_rdata_29[19][38] , \_zyixc_ctx_rdata_29[19][37] , 
	\_zyixc_ctx_rdata_29[19][36] , \_zyixc_ctx_rdata_29[19][35] , 
	\_zyixc_ctx_rdata_29[19][34] , \_zyixc_ctx_rdata_29[19][33] , 
	\_zyixc_ctx_rdata_29[19][32] , \_zyixc_ctx_rdata_29[19][31] , 
	\_zyixc_ctx_rdata_29[19][30] , \_zyixc_ctx_rdata_29[19][29] , 
	\_zyixc_ctx_rdata_29[19][28] , \_zyixc_ctx_rdata_29[19][27] , 
	\_zyixc_ctx_rdata_29[19][26] , \_zyixc_ctx_rdata_29[19][25] , 
	\_zyixc_ctx_rdata_29[19][24] , \_zyixc_ctx_rdata_29[19][23] , 
	\_zyixc_ctx_rdata_29[19][22] , \_zyixc_ctx_rdata_29[19][21] , 
	\_zyixc_ctx_rdata_29[19][20] , \_zyixc_ctx_rdata_29[19][19] , 
	\_zyixc_ctx_rdata_29[19][18] , \_zyixc_ctx_rdata_29[19][17] , 
	\_zyixc_ctx_rdata_29[19][16] , \_zyixc_ctx_rdata_29[19][15] , 
	\_zyixc_ctx_rdata_29[19][14] , \_zyixc_ctx_rdata_29[19][13] , 
	\_zyixc_ctx_rdata_29[19][12] , \_zyixc_ctx_rdata_29[19][11] , 
	\_zyixc_ctx_rdata_29[19][10] , \_zyixc_ctx_rdata_29[19][9] , 
	\_zyixc_ctx_rdata_29[19][8] , \_zyixc_ctx_rdata_29[19][7] , 
	\_zyixc_ctx_rdata_29[19][6] , \_zyixc_ctx_rdata_29[19][5] , 
	\_zyixc_ctx_rdata_29[19][4] , \_zyixc_ctx_rdata_29[19][3] , 
	\_zyixc_ctx_rdata_29[19][2] , \_zyixc_ctx_rdata_29[19][1] , 
	\_zyixc_ctx_rdata_29[19][0] , \_zyixc_ctx_rdata_29[20][63] , 
	\_zyixc_ctx_rdata_29[20][62] , \_zyixc_ctx_rdata_29[20][61] , 
	\_zyixc_ctx_rdata_29[20][60] , \_zyixc_ctx_rdata_29[20][59] , 
	\_zyixc_ctx_rdata_29[20][58] , \_zyixc_ctx_rdata_29[20][57] , 
	\_zyixc_ctx_rdata_29[20][56] , \_zyixc_ctx_rdata_29[20][55] , 
	\_zyixc_ctx_rdata_29[20][54] , \_zyixc_ctx_rdata_29[20][53] , 
	\_zyixc_ctx_rdata_29[20][52] , \_zyixc_ctx_rdata_29[20][51] , 
	\_zyixc_ctx_rdata_29[20][50] , \_zyixc_ctx_rdata_29[20][49] , 
	\_zyixc_ctx_rdata_29[20][48] , \_zyixc_ctx_rdata_29[20][47] , 
	\_zyixc_ctx_rdata_29[20][46] , \_zyixc_ctx_rdata_29[20][45] , 
	\_zyixc_ctx_rdata_29[20][44] , \_zyixc_ctx_rdata_29[20][43] , 
	\_zyixc_ctx_rdata_29[20][42] , \_zyixc_ctx_rdata_29[20][41] , 
	\_zyixc_ctx_rdata_29[20][40] , \_zyixc_ctx_rdata_29[20][39] , 
	\_zyixc_ctx_rdata_29[20][38] , \_zyixc_ctx_rdata_29[20][37] , 
	\_zyixc_ctx_rdata_29[20][36] , \_zyixc_ctx_rdata_29[20][35] , 
	\_zyixc_ctx_rdata_29[20][34] , \_zyixc_ctx_rdata_29[20][33] , 
	\_zyixc_ctx_rdata_29[20][32] , \_zyixc_ctx_rdata_29[20][31] , 
	\_zyixc_ctx_rdata_29[20][30] , \_zyixc_ctx_rdata_29[20][29] , 
	\_zyixc_ctx_rdata_29[20][28] , \_zyixc_ctx_rdata_29[20][27] , 
	\_zyixc_ctx_rdata_29[20][26] , \_zyixc_ctx_rdata_29[20][25] , 
	\_zyixc_ctx_rdata_29[20][24] , \_zyixc_ctx_rdata_29[20][23] , 
	\_zyixc_ctx_rdata_29[20][22] , \_zyixc_ctx_rdata_29[20][21] , 
	\_zyixc_ctx_rdata_29[20][20] , \_zyixc_ctx_rdata_29[20][19] , 
	\_zyixc_ctx_rdata_29[20][18] , \_zyixc_ctx_rdata_29[20][17] , 
	\_zyixc_ctx_rdata_29[20][16] , \_zyixc_ctx_rdata_29[20][15] , 
	\_zyixc_ctx_rdata_29[20][14] , \_zyixc_ctx_rdata_29[20][13] , 
	\_zyixc_ctx_rdata_29[20][12] , \_zyixc_ctx_rdata_29[20][11] , 
	\_zyixc_ctx_rdata_29[20][10] , \_zyixc_ctx_rdata_29[20][9] , 
	\_zyixc_ctx_rdata_29[20][8] , \_zyixc_ctx_rdata_29[20][7] , 
	\_zyixc_ctx_rdata_29[20][6] , \_zyixc_ctx_rdata_29[20][5] , 
	\_zyixc_ctx_rdata_29[20][4] , \_zyixc_ctx_rdata_29[20][3] , 
	\_zyixc_ctx_rdata_29[20][2] , \_zyixc_ctx_rdata_29[20][1] , 
	\_zyixc_ctx_rdata_29[20][0] , \_zyixc_ctx_rdata_29[21][63] , 
	\_zyixc_ctx_rdata_29[21][62] , \_zyixc_ctx_rdata_29[21][61] , 
	\_zyixc_ctx_rdata_29[21][60] , \_zyixc_ctx_rdata_29[21][59] , 
	\_zyixc_ctx_rdata_29[21][58] , \_zyixc_ctx_rdata_29[21][57] , 
	\_zyixc_ctx_rdata_29[21][56] , \_zyixc_ctx_rdata_29[21][55] , 
	\_zyixc_ctx_rdata_29[21][54] , \_zyixc_ctx_rdata_29[21][53] , 
	\_zyixc_ctx_rdata_29[21][52] , \_zyixc_ctx_rdata_29[21][51] , 
	\_zyixc_ctx_rdata_29[21][50] , \_zyixc_ctx_rdata_29[21][49] , 
	\_zyixc_ctx_rdata_29[21][48] , \_zyixc_ctx_rdata_29[21][47] , 
	\_zyixc_ctx_rdata_29[21][46] , \_zyixc_ctx_rdata_29[21][45] , 
	\_zyixc_ctx_rdata_29[21][44] , \_zyixc_ctx_rdata_29[21][43] , 
	\_zyixc_ctx_rdata_29[21][42] , \_zyixc_ctx_rdata_29[21][41] , 
	\_zyixc_ctx_rdata_29[21][40] , \_zyixc_ctx_rdata_29[21][39] , 
	\_zyixc_ctx_rdata_29[21][38] , \_zyixc_ctx_rdata_29[21][37] , 
	\_zyixc_ctx_rdata_29[21][36] , \_zyixc_ctx_rdata_29[21][35] , 
	\_zyixc_ctx_rdata_29[21][34] , \_zyixc_ctx_rdata_29[21][33] , 
	\_zyixc_ctx_rdata_29[21][32] , \_zyixc_ctx_rdata_29[21][31] , 
	\_zyixc_ctx_rdata_29[21][30] , \_zyixc_ctx_rdata_29[21][29] , 
	\_zyixc_ctx_rdata_29[21][28] , \_zyixc_ctx_rdata_29[21][27] , 
	\_zyixc_ctx_rdata_29[21][26] , \_zyixc_ctx_rdata_29[21][25] , 
	\_zyixc_ctx_rdata_29[21][24] , \_zyixc_ctx_rdata_29[21][23] , 
	\_zyixc_ctx_rdata_29[21][22] , \_zyixc_ctx_rdata_29[21][21] , 
	\_zyixc_ctx_rdata_29[21][20] , \_zyixc_ctx_rdata_29[21][19] , 
	\_zyixc_ctx_rdata_29[21][18] , \_zyixc_ctx_rdata_29[21][17] , 
	\_zyixc_ctx_rdata_29[21][16] , \_zyixc_ctx_rdata_29[21][15] , 
	\_zyixc_ctx_rdata_29[21][14] , \_zyixc_ctx_rdata_29[21][13] , 
	\_zyixc_ctx_rdata_29[21][12] , \_zyixc_ctx_rdata_29[21][11] , 
	\_zyixc_ctx_rdata_29[21][10] , \_zyixc_ctx_rdata_29[21][9] , 
	\_zyixc_ctx_rdata_29[21][8] , \_zyixc_ctx_rdata_29[21][7] , 
	\_zyixc_ctx_rdata_29[21][6] , \_zyixc_ctx_rdata_29[21][5] , 
	\_zyixc_ctx_rdata_29[21][4] , \_zyixc_ctx_rdata_29[21][3] , 
	\_zyixc_ctx_rdata_29[21][2] , \_zyixc_ctx_rdata_29[21][1] , 
	\_zyixc_ctx_rdata_29[21][0] , \_zyixc_ctx_rdata_29[22][63] , 
	\_zyixc_ctx_rdata_29[22][62] , \_zyixc_ctx_rdata_29[22][61] , 
	\_zyixc_ctx_rdata_29[22][60] , \_zyixc_ctx_rdata_29[22][59] , 
	\_zyixc_ctx_rdata_29[22][58] , \_zyixc_ctx_rdata_29[22][57] , 
	\_zyixc_ctx_rdata_29[22][56] , \_zyixc_ctx_rdata_29[22][55] , 
	\_zyixc_ctx_rdata_29[22][54] , \_zyixc_ctx_rdata_29[22][53] , 
	\_zyixc_ctx_rdata_29[22][52] , \_zyixc_ctx_rdata_29[22][51] , 
	\_zyixc_ctx_rdata_29[22][50] , \_zyixc_ctx_rdata_29[22][49] , 
	\_zyixc_ctx_rdata_29[22][48] , \_zyixc_ctx_rdata_29[22][47] , 
	\_zyixc_ctx_rdata_29[22][46] , \_zyixc_ctx_rdata_29[22][45] , 
	\_zyixc_ctx_rdata_29[22][44] , \_zyixc_ctx_rdata_29[22][43] , 
	\_zyixc_ctx_rdata_29[22][42] , \_zyixc_ctx_rdata_29[22][41] , 
	\_zyixc_ctx_rdata_29[22][40] , \_zyixc_ctx_rdata_29[22][39] , 
	\_zyixc_ctx_rdata_29[22][38] , \_zyixc_ctx_rdata_29[22][37] , 
	\_zyixc_ctx_rdata_29[22][36] , \_zyixc_ctx_rdata_29[22][35] , 
	\_zyixc_ctx_rdata_29[22][34] , \_zyixc_ctx_rdata_29[22][33] , 
	\_zyixc_ctx_rdata_29[22][32] , \_zyixc_ctx_rdata_29[22][31] , 
	\_zyixc_ctx_rdata_29[22][30] , \_zyixc_ctx_rdata_29[22][29] , 
	\_zyixc_ctx_rdata_29[22][28] , \_zyixc_ctx_rdata_29[22][27] , 
	\_zyixc_ctx_rdata_29[22][26] , \_zyixc_ctx_rdata_29[22][25] , 
	\_zyixc_ctx_rdata_29[22][24] , \_zyixc_ctx_rdata_29[22][23] , 
	\_zyixc_ctx_rdata_29[22][22] , \_zyixc_ctx_rdata_29[22][21] , 
	\_zyixc_ctx_rdata_29[22][20] , \_zyixc_ctx_rdata_29[22][19] , 
	\_zyixc_ctx_rdata_29[22][18] , \_zyixc_ctx_rdata_29[22][17] , 
	\_zyixc_ctx_rdata_29[22][16] , \_zyixc_ctx_rdata_29[22][15] , 
	\_zyixc_ctx_rdata_29[22][14] , \_zyixc_ctx_rdata_29[22][13] , 
	\_zyixc_ctx_rdata_29[22][12] , \_zyixc_ctx_rdata_29[22][11] , 
	\_zyixc_ctx_rdata_29[22][10] , \_zyixc_ctx_rdata_29[22][9] , 
	\_zyixc_ctx_rdata_29[22][8] , \_zyixc_ctx_rdata_29[22][7] , 
	\_zyixc_ctx_rdata_29[22][6] , \_zyixc_ctx_rdata_29[22][5] , 
	\_zyixc_ctx_rdata_29[22][4] , \_zyixc_ctx_rdata_29[22][3] , 
	\_zyixc_ctx_rdata_29[22][2] , \_zyixc_ctx_rdata_29[22][1] , 
	\_zyixc_ctx_rdata_29[22][0] , \_zyixc_ctx_rdata_29[23][63] , 
	\_zyixc_ctx_rdata_29[23][62] , \_zyixc_ctx_rdata_29[23][61] , 
	\_zyixc_ctx_rdata_29[23][60] , \_zyixc_ctx_rdata_29[23][59] , 
	\_zyixc_ctx_rdata_29[23][58] , \_zyixc_ctx_rdata_29[23][57] , 
	\_zyixc_ctx_rdata_29[23][56] , \_zyixc_ctx_rdata_29[23][55] , 
	\_zyixc_ctx_rdata_29[23][54] , \_zyixc_ctx_rdata_29[23][53] , 
	\_zyixc_ctx_rdata_29[23][52] , \_zyixc_ctx_rdata_29[23][51] , 
	\_zyixc_ctx_rdata_29[23][50] , \_zyixc_ctx_rdata_29[23][49] , 
	\_zyixc_ctx_rdata_29[23][48] , \_zyixc_ctx_rdata_29[23][47] , 
	\_zyixc_ctx_rdata_29[23][46] , \_zyixc_ctx_rdata_29[23][45] , 
	\_zyixc_ctx_rdata_29[23][44] , \_zyixc_ctx_rdata_29[23][43] , 
	\_zyixc_ctx_rdata_29[23][42] , \_zyixc_ctx_rdata_29[23][41] , 
	\_zyixc_ctx_rdata_29[23][40] , \_zyixc_ctx_rdata_29[23][39] , 
	\_zyixc_ctx_rdata_29[23][38] , \_zyixc_ctx_rdata_29[23][37] , 
	\_zyixc_ctx_rdata_29[23][36] , \_zyixc_ctx_rdata_29[23][35] , 
	\_zyixc_ctx_rdata_29[23][34] , \_zyixc_ctx_rdata_29[23][33] , 
	\_zyixc_ctx_rdata_29[23][32] , \_zyixc_ctx_rdata_29[23][31] , 
	\_zyixc_ctx_rdata_29[23][30] , \_zyixc_ctx_rdata_29[23][29] , 
	\_zyixc_ctx_rdata_29[23][28] , \_zyixc_ctx_rdata_29[23][27] , 
	\_zyixc_ctx_rdata_29[23][26] , \_zyixc_ctx_rdata_29[23][25] , 
	\_zyixc_ctx_rdata_29[23][24] , \_zyixc_ctx_rdata_29[23][23] , 
	\_zyixc_ctx_rdata_29[23][22] , \_zyixc_ctx_rdata_29[23][21] , 
	\_zyixc_ctx_rdata_29[23][20] , \_zyixc_ctx_rdata_29[23][19] , 
	\_zyixc_ctx_rdata_29[23][18] , \_zyixc_ctx_rdata_29[23][17] , 
	\_zyixc_ctx_rdata_29[23][16] , \_zyixc_ctx_rdata_29[23][15] , 
	\_zyixc_ctx_rdata_29[23][14] , \_zyixc_ctx_rdata_29[23][13] , 
	\_zyixc_ctx_rdata_29[23][12] , \_zyixc_ctx_rdata_29[23][11] , 
	\_zyixc_ctx_rdata_29[23][10] , \_zyixc_ctx_rdata_29[23][9] , 
	\_zyixc_ctx_rdata_29[23][8] , \_zyixc_ctx_rdata_29[23][7] , 
	\_zyixc_ctx_rdata_29[23][6] , \_zyixc_ctx_rdata_29[23][5] , 
	\_zyixc_ctx_rdata_29[23][4] , \_zyixc_ctx_rdata_29[23][3] , 
	\_zyixc_ctx_rdata_29[23][2] , \_zyixc_ctx_rdata_29[23][1] , 
	\_zyixc_ctx_rdata_29[23][0] , \_zyixc_ctx_rdata_29[24][63] , 
	\_zyixc_ctx_rdata_29[24][62] , \_zyixc_ctx_rdata_29[24][61] , 
	\_zyixc_ctx_rdata_29[24][60] , \_zyixc_ctx_rdata_29[24][59] , 
	\_zyixc_ctx_rdata_29[24][58] , \_zyixc_ctx_rdata_29[24][57] , 
	\_zyixc_ctx_rdata_29[24][56] , \_zyixc_ctx_rdata_29[24][55] , 
	\_zyixc_ctx_rdata_29[24][54] , \_zyixc_ctx_rdata_29[24][53] , 
	\_zyixc_ctx_rdata_29[24][52] , \_zyixc_ctx_rdata_29[24][51] , 
	\_zyixc_ctx_rdata_29[24][50] , \_zyixc_ctx_rdata_29[24][49] , 
	\_zyixc_ctx_rdata_29[24][48] , \_zyixc_ctx_rdata_29[24][47] , 
	\_zyixc_ctx_rdata_29[24][46] , \_zyixc_ctx_rdata_29[24][45] , 
	\_zyixc_ctx_rdata_29[24][44] , \_zyixc_ctx_rdata_29[24][43] , 
	\_zyixc_ctx_rdata_29[24][42] , \_zyixc_ctx_rdata_29[24][41] , 
	\_zyixc_ctx_rdata_29[24][40] , \_zyixc_ctx_rdata_29[24][39] , 
	\_zyixc_ctx_rdata_29[24][38] , \_zyixc_ctx_rdata_29[24][37] , 
	\_zyixc_ctx_rdata_29[24][36] , \_zyixc_ctx_rdata_29[24][35] , 
	\_zyixc_ctx_rdata_29[24][34] , \_zyixc_ctx_rdata_29[24][33] , 
	\_zyixc_ctx_rdata_29[24][32] , \_zyixc_ctx_rdata_29[24][31] , 
	\_zyixc_ctx_rdata_29[24][30] , \_zyixc_ctx_rdata_29[24][29] , 
	\_zyixc_ctx_rdata_29[24][28] , \_zyixc_ctx_rdata_29[24][27] , 
	\_zyixc_ctx_rdata_29[24][26] , \_zyixc_ctx_rdata_29[24][25] , 
	\_zyixc_ctx_rdata_29[24][24] , \_zyixc_ctx_rdata_29[24][23] , 
	\_zyixc_ctx_rdata_29[24][22] , \_zyixc_ctx_rdata_29[24][21] , 
	\_zyixc_ctx_rdata_29[24][20] , \_zyixc_ctx_rdata_29[24][19] , 
	\_zyixc_ctx_rdata_29[24][18] , \_zyixc_ctx_rdata_29[24][17] , 
	\_zyixc_ctx_rdata_29[24][16] , \_zyixc_ctx_rdata_29[24][15] , 
	\_zyixc_ctx_rdata_29[24][14] , \_zyixc_ctx_rdata_29[24][13] , 
	\_zyixc_ctx_rdata_29[24][12] , \_zyixc_ctx_rdata_29[24][11] , 
	\_zyixc_ctx_rdata_29[24][10] , \_zyixc_ctx_rdata_29[24][9] , 
	\_zyixc_ctx_rdata_29[24][8] , \_zyixc_ctx_rdata_29[24][7] , 
	\_zyixc_ctx_rdata_29[24][6] , \_zyixc_ctx_rdata_29[24][5] , 
	\_zyixc_ctx_rdata_29[24][4] , \_zyixc_ctx_rdata_29[24][3] , 
	\_zyixc_ctx_rdata_29[24][2] , \_zyixc_ctx_rdata_29[24][1] , 
	\_zyixc_ctx_rdata_29[24][0] , \_zyixc_ctx_rdata_29[25][63] , 
	\_zyixc_ctx_rdata_29[25][62] , \_zyixc_ctx_rdata_29[25][61] , 
	\_zyixc_ctx_rdata_29[25][60] , \_zyixc_ctx_rdata_29[25][59] , 
	\_zyixc_ctx_rdata_29[25][58] , \_zyixc_ctx_rdata_29[25][57] , 
	\_zyixc_ctx_rdata_29[25][56] , \_zyixc_ctx_rdata_29[25][55] , 
	\_zyixc_ctx_rdata_29[25][54] , \_zyixc_ctx_rdata_29[25][53] , 
	\_zyixc_ctx_rdata_29[25][52] , \_zyixc_ctx_rdata_29[25][51] , 
	\_zyixc_ctx_rdata_29[25][50] , \_zyixc_ctx_rdata_29[25][49] , 
	\_zyixc_ctx_rdata_29[25][48] , \_zyixc_ctx_rdata_29[25][47] , 
	\_zyixc_ctx_rdata_29[25][46] , \_zyixc_ctx_rdata_29[25][45] , 
	\_zyixc_ctx_rdata_29[25][44] , \_zyixc_ctx_rdata_29[25][43] , 
	\_zyixc_ctx_rdata_29[25][42] , \_zyixc_ctx_rdata_29[25][41] , 
	\_zyixc_ctx_rdata_29[25][40] , \_zyixc_ctx_rdata_29[25][39] , 
	\_zyixc_ctx_rdata_29[25][38] , \_zyixc_ctx_rdata_29[25][37] , 
	\_zyixc_ctx_rdata_29[25][36] , \_zyixc_ctx_rdata_29[25][35] , 
	\_zyixc_ctx_rdata_29[25][34] , \_zyixc_ctx_rdata_29[25][33] , 
	\_zyixc_ctx_rdata_29[25][32] , \_zyixc_ctx_rdata_29[25][31] , 
	\_zyixc_ctx_rdata_29[25][30] , \_zyixc_ctx_rdata_29[25][29] , 
	\_zyixc_ctx_rdata_29[25][28] , \_zyixc_ctx_rdata_29[25][27] , 
	\_zyixc_ctx_rdata_29[25][26] , \_zyixc_ctx_rdata_29[25][25] , 
	\_zyixc_ctx_rdata_29[25][24] , \_zyixc_ctx_rdata_29[25][23] , 
	\_zyixc_ctx_rdata_29[25][22] , \_zyixc_ctx_rdata_29[25][21] , 
	\_zyixc_ctx_rdata_29[25][20] , \_zyixc_ctx_rdata_29[25][19] , 
	\_zyixc_ctx_rdata_29[25][18] , \_zyixc_ctx_rdata_29[25][17] , 
	\_zyixc_ctx_rdata_29[25][16] , \_zyixc_ctx_rdata_29[25][15] , 
	\_zyixc_ctx_rdata_29[25][14] , \_zyixc_ctx_rdata_29[25][13] , 
	\_zyixc_ctx_rdata_29[25][12] , \_zyixc_ctx_rdata_29[25][11] , 
	\_zyixc_ctx_rdata_29[25][10] , \_zyixc_ctx_rdata_29[25][9] , 
	\_zyixc_ctx_rdata_29[25][8] , \_zyixc_ctx_rdata_29[25][7] , 
	\_zyixc_ctx_rdata_29[25][6] , \_zyixc_ctx_rdata_29[25][5] , 
	\_zyixc_ctx_rdata_29[25][4] , \_zyixc_ctx_rdata_29[25][3] , 
	\_zyixc_ctx_rdata_29[25][2] , \_zyixc_ctx_rdata_29[25][1] , 
	\_zyixc_ctx_rdata_29[25][0] , \_zyixc_ctx_rdata_29[26][63] , 
	\_zyixc_ctx_rdata_29[26][62] , \_zyixc_ctx_rdata_29[26][61] , 
	\_zyixc_ctx_rdata_29[26][60] , \_zyixc_ctx_rdata_29[26][59] , 
	\_zyixc_ctx_rdata_29[26][58] , \_zyixc_ctx_rdata_29[26][57] , 
	\_zyixc_ctx_rdata_29[26][56] , \_zyixc_ctx_rdata_29[26][55] , 
	\_zyixc_ctx_rdata_29[26][54] , \_zyixc_ctx_rdata_29[26][53] , 
	\_zyixc_ctx_rdata_29[26][52] , \_zyixc_ctx_rdata_29[26][51] , 
	\_zyixc_ctx_rdata_29[26][50] , \_zyixc_ctx_rdata_29[26][49] , 
	\_zyixc_ctx_rdata_29[26][48] , \_zyixc_ctx_rdata_29[26][47] , 
	\_zyixc_ctx_rdata_29[26][46] , \_zyixc_ctx_rdata_29[26][45] , 
	\_zyixc_ctx_rdata_29[26][44] , \_zyixc_ctx_rdata_29[26][43] , 
	\_zyixc_ctx_rdata_29[26][42] , \_zyixc_ctx_rdata_29[26][41] , 
	\_zyixc_ctx_rdata_29[26][40] , \_zyixc_ctx_rdata_29[26][39] , 
	\_zyixc_ctx_rdata_29[26][38] , \_zyixc_ctx_rdata_29[26][37] , 
	\_zyixc_ctx_rdata_29[26][36] , \_zyixc_ctx_rdata_29[26][35] , 
	\_zyixc_ctx_rdata_29[26][34] , \_zyixc_ctx_rdata_29[26][33] , 
	\_zyixc_ctx_rdata_29[26][32] , \_zyixc_ctx_rdata_29[26][31] , 
	\_zyixc_ctx_rdata_29[26][30] , \_zyixc_ctx_rdata_29[26][29] , 
	\_zyixc_ctx_rdata_29[26][28] , \_zyixc_ctx_rdata_29[26][27] , 
	\_zyixc_ctx_rdata_29[26][26] , \_zyixc_ctx_rdata_29[26][25] , 
	\_zyixc_ctx_rdata_29[26][24] , \_zyixc_ctx_rdata_29[26][23] , 
	\_zyixc_ctx_rdata_29[26][22] , \_zyixc_ctx_rdata_29[26][21] , 
	\_zyixc_ctx_rdata_29[26][20] , \_zyixc_ctx_rdata_29[26][19] , 
	\_zyixc_ctx_rdata_29[26][18] , \_zyixc_ctx_rdata_29[26][17] , 
	\_zyixc_ctx_rdata_29[26][16] , \_zyixc_ctx_rdata_29[26][15] , 
	\_zyixc_ctx_rdata_29[26][14] , \_zyixc_ctx_rdata_29[26][13] , 
	\_zyixc_ctx_rdata_29[26][12] , \_zyixc_ctx_rdata_29[26][11] , 
	\_zyixc_ctx_rdata_29[26][10] , \_zyixc_ctx_rdata_29[26][9] , 
	\_zyixc_ctx_rdata_29[26][8] , \_zyixc_ctx_rdata_29[26][7] , 
	\_zyixc_ctx_rdata_29[26][6] , \_zyixc_ctx_rdata_29[26][5] , 
	\_zyixc_ctx_rdata_29[26][4] , \_zyixc_ctx_rdata_29[26][3] , 
	\_zyixc_ctx_rdata_29[26][2] , \_zyixc_ctx_rdata_29[26][1] , 
	\_zyixc_ctx_rdata_29[26][0] , \_zyixc_ctx_rdata_29[27][63] , 
	\_zyixc_ctx_rdata_29[27][62] , \_zyixc_ctx_rdata_29[27][61] , 
	\_zyixc_ctx_rdata_29[27][60] , \_zyixc_ctx_rdata_29[27][59] , 
	\_zyixc_ctx_rdata_29[27][58] , \_zyixc_ctx_rdata_29[27][57] , 
	\_zyixc_ctx_rdata_29[27][56] , \_zyixc_ctx_rdata_29[27][55] , 
	\_zyixc_ctx_rdata_29[27][54] , \_zyixc_ctx_rdata_29[27][53] , 
	\_zyixc_ctx_rdata_29[27][52] , \_zyixc_ctx_rdata_29[27][51] , 
	\_zyixc_ctx_rdata_29[27][50] , \_zyixc_ctx_rdata_29[27][49] , 
	\_zyixc_ctx_rdata_29[27][48] , \_zyixc_ctx_rdata_29[27][47] , 
	\_zyixc_ctx_rdata_29[27][46] , \_zyixc_ctx_rdata_29[27][45] , 
	\_zyixc_ctx_rdata_29[27][44] , \_zyixc_ctx_rdata_29[27][43] , 
	\_zyixc_ctx_rdata_29[27][42] , \_zyixc_ctx_rdata_29[27][41] , 
	\_zyixc_ctx_rdata_29[27][40] , \_zyixc_ctx_rdata_29[27][39] , 
	\_zyixc_ctx_rdata_29[27][38] , \_zyixc_ctx_rdata_29[27][37] , 
	\_zyixc_ctx_rdata_29[27][36] , \_zyixc_ctx_rdata_29[27][35] , 
	\_zyixc_ctx_rdata_29[27][34] , \_zyixc_ctx_rdata_29[27][33] , 
	\_zyixc_ctx_rdata_29[27][32] , \_zyixc_ctx_rdata_29[27][31] , 
	\_zyixc_ctx_rdata_29[27][30] , \_zyixc_ctx_rdata_29[27][29] , 
	\_zyixc_ctx_rdata_29[27][28] , \_zyixc_ctx_rdata_29[27][27] , 
	\_zyixc_ctx_rdata_29[27][26] , \_zyixc_ctx_rdata_29[27][25] , 
	\_zyixc_ctx_rdata_29[27][24] , \_zyixc_ctx_rdata_29[27][23] , 
	\_zyixc_ctx_rdata_29[27][22] , \_zyixc_ctx_rdata_29[27][21] , 
	\_zyixc_ctx_rdata_29[27][20] , \_zyixc_ctx_rdata_29[27][19] , 
	\_zyixc_ctx_rdata_29[27][18] , \_zyixc_ctx_rdata_29[27][17] , 
	\_zyixc_ctx_rdata_29[27][16] , \_zyixc_ctx_rdata_29[27][15] , 
	\_zyixc_ctx_rdata_29[27][14] , \_zyixc_ctx_rdata_29[27][13] , 
	\_zyixc_ctx_rdata_29[27][12] , \_zyixc_ctx_rdata_29[27][11] , 
	\_zyixc_ctx_rdata_29[27][10] , \_zyixc_ctx_rdata_29[27][9] , 
	\_zyixc_ctx_rdata_29[27][8] , \_zyixc_ctx_rdata_29[27][7] , 
	\_zyixc_ctx_rdata_29[27][6] , \_zyixc_ctx_rdata_29[27][5] , 
	\_zyixc_ctx_rdata_29[27][4] , \_zyixc_ctx_rdata_29[27][3] , 
	\_zyixc_ctx_rdata_29[27][2] , \_zyixc_ctx_rdata_29[27][1] , 
	\_zyixc_ctx_rdata_29[27][0] , \_zyixc_ctx_rdata_29[28][63] , 
	\_zyixc_ctx_rdata_29[28][62] , \_zyixc_ctx_rdata_29[28][61] , 
	\_zyixc_ctx_rdata_29[28][60] , \_zyixc_ctx_rdata_29[28][59] , 
	\_zyixc_ctx_rdata_29[28][58] , \_zyixc_ctx_rdata_29[28][57] , 
	\_zyixc_ctx_rdata_29[28][56] , \_zyixc_ctx_rdata_29[28][55] , 
	\_zyixc_ctx_rdata_29[28][54] , \_zyixc_ctx_rdata_29[28][53] , 
	\_zyixc_ctx_rdata_29[28][52] , \_zyixc_ctx_rdata_29[28][51] , 
	\_zyixc_ctx_rdata_29[28][50] , \_zyixc_ctx_rdata_29[28][49] , 
	\_zyixc_ctx_rdata_29[28][48] , \_zyixc_ctx_rdata_29[28][47] , 
	\_zyixc_ctx_rdata_29[28][46] , \_zyixc_ctx_rdata_29[28][45] , 
	\_zyixc_ctx_rdata_29[28][44] , \_zyixc_ctx_rdata_29[28][43] , 
	\_zyixc_ctx_rdata_29[28][42] , \_zyixc_ctx_rdata_29[28][41] , 
	\_zyixc_ctx_rdata_29[28][40] , \_zyixc_ctx_rdata_29[28][39] , 
	\_zyixc_ctx_rdata_29[28][38] , \_zyixc_ctx_rdata_29[28][37] , 
	\_zyixc_ctx_rdata_29[28][36] , \_zyixc_ctx_rdata_29[28][35] , 
	\_zyixc_ctx_rdata_29[28][34] , \_zyixc_ctx_rdata_29[28][33] , 
	\_zyixc_ctx_rdata_29[28][32] , \_zyixc_ctx_rdata_29[28][31] , 
	\_zyixc_ctx_rdata_29[28][30] , \_zyixc_ctx_rdata_29[28][29] , 
	\_zyixc_ctx_rdata_29[28][28] , \_zyixc_ctx_rdata_29[28][27] , 
	\_zyixc_ctx_rdata_29[28][26] , \_zyixc_ctx_rdata_29[28][25] , 
	\_zyixc_ctx_rdata_29[28][24] , \_zyixc_ctx_rdata_29[28][23] , 
	\_zyixc_ctx_rdata_29[28][22] , \_zyixc_ctx_rdata_29[28][21] , 
	\_zyixc_ctx_rdata_29[28][20] , \_zyixc_ctx_rdata_29[28][19] , 
	\_zyixc_ctx_rdata_29[28][18] , \_zyixc_ctx_rdata_29[28][17] , 
	\_zyixc_ctx_rdata_29[28][16] , \_zyixc_ctx_rdata_29[28][15] , 
	\_zyixc_ctx_rdata_29[28][14] , \_zyixc_ctx_rdata_29[28][13] , 
	\_zyixc_ctx_rdata_29[28][12] , \_zyixc_ctx_rdata_29[28][11] , 
	\_zyixc_ctx_rdata_29[28][10] , \_zyixc_ctx_rdata_29[28][9] , 
	\_zyixc_ctx_rdata_29[28][8] , \_zyixc_ctx_rdata_29[28][7] , 
	\_zyixc_ctx_rdata_29[28][6] , \_zyixc_ctx_rdata_29[28][5] , 
	\_zyixc_ctx_rdata_29[28][4] , \_zyixc_ctx_rdata_29[28][3] , 
	\_zyixc_ctx_rdata_29[28][2] , \_zyixc_ctx_rdata_29[28][1] , 
	\_zyixc_ctx_rdata_29[28][0] , \_zyixc_ctx_rdata_29[29][63] , 
	\_zyixc_ctx_rdata_29[29][62] , \_zyixc_ctx_rdata_29[29][61] , 
	\_zyixc_ctx_rdata_29[29][60] , \_zyixc_ctx_rdata_29[29][59] , 
	\_zyixc_ctx_rdata_29[29][58] , \_zyixc_ctx_rdata_29[29][57] , 
	\_zyixc_ctx_rdata_29[29][56] , \_zyixc_ctx_rdata_29[29][55] , 
	\_zyixc_ctx_rdata_29[29][54] , \_zyixc_ctx_rdata_29[29][53] , 
	\_zyixc_ctx_rdata_29[29][52] , \_zyixc_ctx_rdata_29[29][51] , 
	\_zyixc_ctx_rdata_29[29][50] , \_zyixc_ctx_rdata_29[29][49] , 
	\_zyixc_ctx_rdata_29[29][48] , \_zyixc_ctx_rdata_29[29][47] , 
	\_zyixc_ctx_rdata_29[29][46] , \_zyixc_ctx_rdata_29[29][45] , 
	\_zyixc_ctx_rdata_29[29][44] , \_zyixc_ctx_rdata_29[29][43] , 
	\_zyixc_ctx_rdata_29[29][42] , \_zyixc_ctx_rdata_29[29][41] , 
	\_zyixc_ctx_rdata_29[29][40] , \_zyixc_ctx_rdata_29[29][39] , 
	\_zyixc_ctx_rdata_29[29][38] , \_zyixc_ctx_rdata_29[29][37] , 
	\_zyixc_ctx_rdata_29[29][36] , \_zyixc_ctx_rdata_29[29][35] , 
	\_zyixc_ctx_rdata_29[29][34] , \_zyixc_ctx_rdata_29[29][33] , 
	\_zyixc_ctx_rdata_29[29][32] , \_zyixc_ctx_rdata_29[29][31] , 
	\_zyixc_ctx_rdata_29[29][30] , \_zyixc_ctx_rdata_29[29][29] , 
	\_zyixc_ctx_rdata_29[29][28] , \_zyixc_ctx_rdata_29[29][27] , 
	\_zyixc_ctx_rdata_29[29][26] , \_zyixc_ctx_rdata_29[29][25] , 
	\_zyixc_ctx_rdata_29[29][24] , \_zyixc_ctx_rdata_29[29][23] , 
	\_zyixc_ctx_rdata_29[29][22] , \_zyixc_ctx_rdata_29[29][21] , 
	\_zyixc_ctx_rdata_29[29][20] , \_zyixc_ctx_rdata_29[29][19] , 
	\_zyixc_ctx_rdata_29[29][18] , \_zyixc_ctx_rdata_29[29][17] , 
	\_zyixc_ctx_rdata_29[29][16] , \_zyixc_ctx_rdata_29[29][15] , 
	\_zyixc_ctx_rdata_29[29][14] , \_zyixc_ctx_rdata_29[29][13] , 
	\_zyixc_ctx_rdata_29[29][12] , \_zyixc_ctx_rdata_29[29][11] , 
	\_zyixc_ctx_rdata_29[29][10] , \_zyixc_ctx_rdata_29[29][9] , 
	\_zyixc_ctx_rdata_29[29][8] , \_zyixc_ctx_rdata_29[29][7] , 
	\_zyixc_ctx_rdata_29[29][6] , \_zyixc_ctx_rdata_29[29][5] , 
	\_zyixc_ctx_rdata_29[29][4] , \_zyixc_ctx_rdata_29[29][3] , 
	\_zyixc_ctx_rdata_29[29][2] , \_zyixc_ctx_rdata_29[29][1] , 
	\_zyixc_ctx_rdata_29[29][0] , \_zyixc_ctx_rdata_29[30][63] , 
	\_zyixc_ctx_rdata_29[30][62] , \_zyixc_ctx_rdata_29[30][61] , 
	\_zyixc_ctx_rdata_29[30][60] , \_zyixc_ctx_rdata_29[30][59] , 
	\_zyixc_ctx_rdata_29[30][58] , \_zyixc_ctx_rdata_29[30][57] , 
	\_zyixc_ctx_rdata_29[30][56] , \_zyixc_ctx_rdata_29[30][55] , 
	\_zyixc_ctx_rdata_29[30][54] , \_zyixc_ctx_rdata_29[30][53] , 
	\_zyixc_ctx_rdata_29[30][52] , \_zyixc_ctx_rdata_29[30][51] , 
	\_zyixc_ctx_rdata_29[30][50] , \_zyixc_ctx_rdata_29[30][49] , 
	\_zyixc_ctx_rdata_29[30][48] , \_zyixc_ctx_rdata_29[30][47] , 
	\_zyixc_ctx_rdata_29[30][46] , \_zyixc_ctx_rdata_29[30][45] , 
	\_zyixc_ctx_rdata_29[30][44] , \_zyixc_ctx_rdata_29[30][43] , 
	\_zyixc_ctx_rdata_29[30][42] , \_zyixc_ctx_rdata_29[30][41] , 
	\_zyixc_ctx_rdata_29[30][40] , \_zyixc_ctx_rdata_29[30][39] , 
	\_zyixc_ctx_rdata_29[30][38] , \_zyixc_ctx_rdata_29[30][37] , 
	\_zyixc_ctx_rdata_29[30][36] , \_zyixc_ctx_rdata_29[30][35] , 
	\_zyixc_ctx_rdata_29[30][34] , \_zyixc_ctx_rdata_29[30][33] , 
	\_zyixc_ctx_rdata_29[30][32] , \_zyixc_ctx_rdata_29[30][31] , 
	\_zyixc_ctx_rdata_29[30][30] , \_zyixc_ctx_rdata_29[30][29] , 
	\_zyixc_ctx_rdata_29[30][28] , \_zyixc_ctx_rdata_29[30][27] , 
	\_zyixc_ctx_rdata_29[30][26] , \_zyixc_ctx_rdata_29[30][25] , 
	\_zyixc_ctx_rdata_29[30][24] , \_zyixc_ctx_rdata_29[30][23] , 
	\_zyixc_ctx_rdata_29[30][22] , \_zyixc_ctx_rdata_29[30][21] , 
	\_zyixc_ctx_rdata_29[30][20] , \_zyixc_ctx_rdata_29[30][19] , 
	\_zyixc_ctx_rdata_29[30][18] , \_zyixc_ctx_rdata_29[30][17] , 
	\_zyixc_ctx_rdata_29[30][16] , \_zyixc_ctx_rdata_29[30][15] , 
	\_zyixc_ctx_rdata_29[30][14] , \_zyixc_ctx_rdata_29[30][13] , 
	\_zyixc_ctx_rdata_29[30][12] , \_zyixc_ctx_rdata_29[30][11] , 
	\_zyixc_ctx_rdata_29[30][10] , \_zyixc_ctx_rdata_29[30][9] , 
	\_zyixc_ctx_rdata_29[30][8] , \_zyixc_ctx_rdata_29[30][7] , 
	\_zyixc_ctx_rdata_29[30][6] , \_zyixc_ctx_rdata_29[30][5] , 
	\_zyixc_ctx_rdata_29[30][4] , \_zyixc_ctx_rdata_29[30][3] , 
	\_zyixc_ctx_rdata_29[30][2] , \_zyixc_ctx_rdata_29[30][1] , 
	\_zyixc_ctx_rdata_29[30][0] , \_zyixc_ctx_rdata_29[31][63] , 
	\_zyixc_ctx_rdata_29[31][62] , \_zyixc_ctx_rdata_29[31][61] , 
	\_zyixc_ctx_rdata_29[31][60] , \_zyixc_ctx_rdata_29[31][59] , 
	\_zyixc_ctx_rdata_29[31][58] , \_zyixc_ctx_rdata_29[31][57] , 
	\_zyixc_ctx_rdata_29[31][56] , \_zyixc_ctx_rdata_29[31][55] , 
	\_zyixc_ctx_rdata_29[31][54] , \_zyixc_ctx_rdata_29[31][53] , 
	\_zyixc_ctx_rdata_29[31][52] , \_zyixc_ctx_rdata_29[31][51] , 
	\_zyixc_ctx_rdata_29[31][50] , \_zyixc_ctx_rdata_29[31][49] , 
	\_zyixc_ctx_rdata_29[31][48] , \_zyixc_ctx_rdata_29[31][47] , 
	\_zyixc_ctx_rdata_29[31][46] , \_zyixc_ctx_rdata_29[31][45] , 
	\_zyixc_ctx_rdata_29[31][44] , \_zyixc_ctx_rdata_29[31][43] , 
	\_zyixc_ctx_rdata_29[31][42] , \_zyixc_ctx_rdata_29[31][41] , 
	\_zyixc_ctx_rdata_29[31][40] , \_zyixc_ctx_rdata_29[31][39] , 
	\_zyixc_ctx_rdata_29[31][38] , \_zyixc_ctx_rdata_29[31][37] , 
	\_zyixc_ctx_rdata_29[31][36] , \_zyixc_ctx_rdata_29[31][35] , 
	\_zyixc_ctx_rdata_29[31][34] , \_zyixc_ctx_rdata_29[31][33] , 
	\_zyixc_ctx_rdata_29[31][32] , \_zyixc_ctx_rdata_29[31][31] , 
	\_zyixc_ctx_rdata_29[31][30] , \_zyixc_ctx_rdata_29[31][29] , 
	\_zyixc_ctx_rdata_29[31][28] , \_zyixc_ctx_rdata_29[31][27] , 
	\_zyixc_ctx_rdata_29[31][26] , \_zyixc_ctx_rdata_29[31][25] , 
	\_zyixc_ctx_rdata_29[31][24] , \_zyixc_ctx_rdata_29[31][23] , 
	\_zyixc_ctx_rdata_29[31][22] , \_zyixc_ctx_rdata_29[31][21] , 
	\_zyixc_ctx_rdata_29[31][20] , \_zyixc_ctx_rdata_29[31][19] , 
	\_zyixc_ctx_rdata_29[31][18] , \_zyixc_ctx_rdata_29[31][17] , 
	\_zyixc_ctx_rdata_29[31][16] , \_zyixc_ctx_rdata_29[31][15] , 
	\_zyixc_ctx_rdata_29[31][14] , \_zyixc_ctx_rdata_29[31][13] , 
	\_zyixc_ctx_rdata_29[31][12] , \_zyixc_ctx_rdata_29[31][11] , 
	\_zyixc_ctx_rdata_29[31][10] , \_zyixc_ctx_rdata_29[31][9] , 
	\_zyixc_ctx_rdata_29[31][8] , \_zyixc_ctx_rdata_29[31][7] , 
	\_zyixc_ctx_rdata_29[31][6] , \_zyixc_ctx_rdata_29[31][5] , 
	\_zyixc_ctx_rdata_29[31][4] , \_zyixc_ctx_rdata_29[31][3] , 
	\_zyixc_ctx_rdata_29[31][2] , \_zyixc_ctx_rdata_29[31][1] , 
	\_zyixc_ctx_rdata_29[31][0] });
ixc_assign _zz_strnp_20 ( reset, _zy_simnet_reset_27_w$);
ixc_assign_64 _zz_strnp_19 ( _zy_simnet_sw_rdat_22_w$[0:63], sw_rdat[63:0]);
ixc_assign_64 _zz_strnp_18 ( sw_wdat[63:0], _zy_simnet_sw_wdat_21_w$[0:63]);
ixc_assign_5 _zz_strnp_17 ( sw_add[4:0], _zy_simnet_sw_add_20_w$[0:4]);
ixc_assign _zz_strnp_16 ( sw_we, _zy_simnet_sw_we_19_w$);
ixc_assign _zz_strnp_15 ( sw_cs, _zy_simnet_sw_cs_17_w$);
ixc_assign_64 _zz_strnp_14 ( rd_dat[63:0], _zy_simnet_rd_dat_16_w$[0:63]);
ixc_assign_5 _zz_strnp_13 ( _zy_simnet_addr_limit_14_w$[0:4], addr_limit[4:0]);
ixc_assign_4 _zz_strnp_12 ( capability_type[3:0], 
	_zy_simnet_capability_type_12_w$[0:3]);
ixc_assign_16 _zz_strnp_11 ( capability_lst[15:0], 
	_zy_simnet_capability_lst_11_w$[0:15]);
ixc_assign_5 _zz_strnp_10 ( stat_addr[4:0], _zy_simnet_stat_addr_9_w$[0:4]);
ixc_assign_5 _zz_strnp_9 ( stat_datawords[4:0], 
	_zy_simnet_stat_datawords_8_w$[0:4]);
ixc_assign_3 _zz_strnp_8 ( stat_code[2:0], _zy_simnet_stat_code_7_w$[0:2]);
ixc_assign_64 _zz_strnp_7 ( _zy_simnet_rd_dat_5_w$[0:63], rd_dat[63:0]);
ixc_assign_4 _zz_strnp_6 ( _zy_simnet_capability_type_4_w$[0:3], 
	capability_type[3:0]);
ixc_assign_16 _zz_strnp_5 ( _zy_simnet_capability_lst_3_w$[0:15], 
	capability_lst[15:0]);
ixc_assign_5 _zz_strnp_4 ( _zy_simnet_stat_addr_2_w$[0:4], stat_addr[4:0]);
ixc_assign_5 _zz_strnp_3 ( _zy_simnet_stat_datawords_1_w$[0:4], 
	stat_datawords[4:0]);
ixc_assign_3 _zz_strnp_2 ( _zy_simnet_stat_code_0_w$[0:2], stat_code[2:0]);
Q_MX08 U97 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][0] ), .A1(\mem_a[25][0] ), .A2(\mem_a[26][0] ), .A3(\mem_a[27][0] ), .A4(\mem_a[28][0] ), .A5(\mem_a[29][0] ), .A6(\mem_a[30][0] ), .A7(\mem_a[31][0] ), .Z(n3));
Q_MX08 U98 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][0] ), .A1(\mem_a[17][0] ), .A2(\mem_a[18][0] ), .A3(\mem_a[19][0] ), .A4(\mem_a[20][0] ), .A5(\mem_a[21][0] ), .A6(\mem_a[22][0] ), .A7(\mem_a[23][0] ), .Z(n4));
Q_MX08 U99 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][0] ), .A1(\mem_a[9][0] ), .A2(\mem_a[10][0] ), .A3(\mem_a[11][0] ), .A4(\mem_a[12][0] ), .A5(\mem_a[13][0] ), .A6(\mem_a[14][0] ), .A7(\mem_a[15][0] ), .Z(n5));
Q_MX08 U100 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][0] ), .A1(\mem_a[1][0] ), .A2(\mem_a[2][0] ), .A3(\mem_a[3][0] ), .A4(\mem_a[4][0] ), .A5(\mem_a[5][0] ), .A6(\mem_a[6][0] ), .A7(\mem_a[7][0] ), .Z(n6));
Q_MX04 U101 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n6), .A1(n5), .A2(n4), .A3(n3), .Z(n7));
Q_MX08 U102 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][1] ), .A1(\mem_a[25][1] ), .A2(\mem_a[26][1] ), .A3(\mem_a[27][1] ), .A4(\mem_a[28][1] ), .A5(\mem_a[29][1] ), .A6(\mem_a[30][1] ), .A7(\mem_a[31][1] ), .Z(n8));
Q_MX08 U103 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][1] ), .A1(\mem_a[17][1] ), .A2(\mem_a[18][1] ), .A3(\mem_a[19][1] ), .A4(\mem_a[20][1] ), .A5(\mem_a[21][1] ), .A6(\mem_a[22][1] ), .A7(\mem_a[23][1] ), .Z(n9));
Q_MX08 U104 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][1] ), .A1(\mem_a[9][1] ), .A2(\mem_a[10][1] ), .A3(\mem_a[11][1] ), .A4(\mem_a[12][1] ), .A5(\mem_a[13][1] ), .A6(\mem_a[14][1] ), .A7(\mem_a[15][1] ), .Z(n10));
Q_MX08 U105 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][1] ), .A1(\mem_a[1][1] ), .A2(\mem_a[2][1] ), .A3(\mem_a[3][1] ), .A4(\mem_a[4][1] ), .A5(\mem_a[5][1] ), .A6(\mem_a[6][1] ), .A7(\mem_a[7][1] ), .Z(n11));
Q_MX04 U106 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n11), .A1(n10), .A2(n9), .A3(n8), .Z(n12));
Q_MX08 U107 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][2] ), .A1(\mem_a[25][2] ), .A2(\mem_a[26][2] ), .A3(\mem_a[27][2] ), .A4(\mem_a[28][2] ), .A5(\mem_a[29][2] ), .A6(\mem_a[30][2] ), .A7(\mem_a[31][2] ), .Z(n13));
Q_MX08 U108 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][2] ), .A1(\mem_a[17][2] ), .A2(\mem_a[18][2] ), .A3(\mem_a[19][2] ), .A4(\mem_a[20][2] ), .A5(\mem_a[21][2] ), .A6(\mem_a[22][2] ), .A7(\mem_a[23][2] ), .Z(n14));
Q_MX08 U109 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][2] ), .A1(\mem_a[9][2] ), .A2(\mem_a[10][2] ), .A3(\mem_a[11][2] ), .A4(\mem_a[12][2] ), .A5(\mem_a[13][2] ), .A6(\mem_a[14][2] ), .A7(\mem_a[15][2] ), .Z(n15));
Q_MX08 U110 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][2] ), .A1(\mem_a[1][2] ), .A2(\mem_a[2][2] ), .A3(\mem_a[3][2] ), .A4(\mem_a[4][2] ), .A5(\mem_a[5][2] ), .A6(\mem_a[6][2] ), .A7(\mem_a[7][2] ), .Z(n16));
Q_MX04 U111 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n16), .A1(n15), .A2(n14), .A3(n13), .Z(n17));
Q_MX08 U112 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][3] ), .A1(\mem_a[25][3] ), .A2(\mem_a[26][3] ), .A3(\mem_a[27][3] ), .A4(\mem_a[28][3] ), .A5(\mem_a[29][3] ), .A6(\mem_a[30][3] ), .A7(\mem_a[31][3] ), .Z(n18));
Q_MX08 U113 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][3] ), .A1(\mem_a[17][3] ), .A2(\mem_a[18][3] ), .A3(\mem_a[19][3] ), .A4(\mem_a[20][3] ), .A5(\mem_a[21][3] ), .A6(\mem_a[22][3] ), .A7(\mem_a[23][3] ), .Z(n19));
Q_MX08 U114 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][3] ), .A1(\mem_a[9][3] ), .A2(\mem_a[10][3] ), .A3(\mem_a[11][3] ), .A4(\mem_a[12][3] ), .A5(\mem_a[13][3] ), .A6(\mem_a[14][3] ), .A7(\mem_a[15][3] ), .Z(n20));
Q_MX08 U115 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][3] ), .A1(\mem_a[1][3] ), .A2(\mem_a[2][3] ), .A3(\mem_a[3][3] ), .A4(\mem_a[4][3] ), .A5(\mem_a[5][3] ), .A6(\mem_a[6][3] ), .A7(\mem_a[7][3] ), .Z(n21));
Q_MX04 U116 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n21), .A1(n20), .A2(n19), .A3(n18), .Z(n22));
Q_MX08 U117 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][4] ), .A1(\mem_a[25][4] ), .A2(\mem_a[26][4] ), .A3(\mem_a[27][4] ), .A4(\mem_a[28][4] ), .A5(\mem_a[29][4] ), .A6(\mem_a[30][4] ), .A7(\mem_a[31][4] ), .Z(n23));
Q_MX08 U118 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][4] ), .A1(\mem_a[17][4] ), .A2(\mem_a[18][4] ), .A3(\mem_a[19][4] ), .A4(\mem_a[20][4] ), .A5(\mem_a[21][4] ), .A6(\mem_a[22][4] ), .A7(\mem_a[23][4] ), .Z(n24));
Q_MX08 U119 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][4] ), .A1(\mem_a[9][4] ), .A2(\mem_a[10][4] ), .A3(\mem_a[11][4] ), .A4(\mem_a[12][4] ), .A5(\mem_a[13][4] ), .A6(\mem_a[14][4] ), .A7(\mem_a[15][4] ), .Z(n25));
Q_MX08 U120 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][4] ), .A1(\mem_a[1][4] ), .A2(\mem_a[2][4] ), .A3(\mem_a[3][4] ), .A4(\mem_a[4][4] ), .A5(\mem_a[5][4] ), .A6(\mem_a[6][4] ), .A7(\mem_a[7][4] ), .Z(n26));
Q_MX04 U121 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n26), .A1(n25), .A2(n24), .A3(n23), .Z(n27));
Q_MX08 U122 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][5] ), .A1(\mem_a[25][5] ), .A2(\mem_a[26][5] ), .A3(\mem_a[27][5] ), .A4(\mem_a[28][5] ), .A5(\mem_a[29][5] ), .A6(\mem_a[30][5] ), .A7(\mem_a[31][5] ), .Z(n28));
Q_MX08 U123 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][5] ), .A1(\mem_a[17][5] ), .A2(\mem_a[18][5] ), .A3(\mem_a[19][5] ), .A4(\mem_a[20][5] ), .A5(\mem_a[21][5] ), .A6(\mem_a[22][5] ), .A7(\mem_a[23][5] ), .Z(n29));
Q_MX08 U124 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][5] ), .A1(\mem_a[9][5] ), .A2(\mem_a[10][5] ), .A3(\mem_a[11][5] ), .A4(\mem_a[12][5] ), .A5(\mem_a[13][5] ), .A6(\mem_a[14][5] ), .A7(\mem_a[15][5] ), .Z(n30));
Q_MX08 U125 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][5] ), .A1(\mem_a[1][5] ), .A2(\mem_a[2][5] ), .A3(\mem_a[3][5] ), .A4(\mem_a[4][5] ), .A5(\mem_a[5][5] ), .A6(\mem_a[6][5] ), .A7(\mem_a[7][5] ), .Z(n31));
Q_MX04 U126 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n31), .A1(n30), .A2(n29), .A3(n28), .Z(n32));
Q_MX08 U127 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][6] ), .A1(\mem_a[25][6] ), .A2(\mem_a[26][6] ), .A3(\mem_a[27][6] ), .A4(\mem_a[28][6] ), .A5(\mem_a[29][6] ), .A6(\mem_a[30][6] ), .A7(\mem_a[31][6] ), .Z(n33));
Q_MX08 U128 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][6] ), .A1(\mem_a[17][6] ), .A2(\mem_a[18][6] ), .A3(\mem_a[19][6] ), .A4(\mem_a[20][6] ), .A5(\mem_a[21][6] ), .A6(\mem_a[22][6] ), .A7(\mem_a[23][6] ), .Z(n34));
Q_MX08 U129 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][6] ), .A1(\mem_a[9][6] ), .A2(\mem_a[10][6] ), .A3(\mem_a[11][6] ), .A4(\mem_a[12][6] ), .A5(\mem_a[13][6] ), .A6(\mem_a[14][6] ), .A7(\mem_a[15][6] ), .Z(n35));
Q_MX08 U130 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][6] ), .A1(\mem_a[1][6] ), .A2(\mem_a[2][6] ), .A3(\mem_a[3][6] ), .A4(\mem_a[4][6] ), .A5(\mem_a[5][6] ), .A6(\mem_a[6][6] ), .A7(\mem_a[7][6] ), .Z(n36));
Q_MX04 U131 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n36), .A1(n35), .A2(n34), .A3(n33), .Z(n37));
Q_MX08 U132 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][7] ), .A1(\mem_a[25][7] ), .A2(\mem_a[26][7] ), .A3(\mem_a[27][7] ), .A4(\mem_a[28][7] ), .A5(\mem_a[29][7] ), .A6(\mem_a[30][7] ), .A7(\mem_a[31][7] ), .Z(n38));
Q_MX08 U133 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][7] ), .A1(\mem_a[17][7] ), .A2(\mem_a[18][7] ), .A3(\mem_a[19][7] ), .A4(\mem_a[20][7] ), .A5(\mem_a[21][7] ), .A6(\mem_a[22][7] ), .A7(\mem_a[23][7] ), .Z(n39));
Q_MX08 U134 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][7] ), .A1(\mem_a[9][7] ), .A2(\mem_a[10][7] ), .A3(\mem_a[11][7] ), .A4(\mem_a[12][7] ), .A5(\mem_a[13][7] ), .A6(\mem_a[14][7] ), .A7(\mem_a[15][7] ), .Z(n40));
Q_MX08 U135 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][7] ), .A1(\mem_a[1][7] ), .A2(\mem_a[2][7] ), .A3(\mem_a[3][7] ), .A4(\mem_a[4][7] ), .A5(\mem_a[5][7] ), .A6(\mem_a[6][7] ), .A7(\mem_a[7][7] ), .Z(n41));
Q_MX04 U136 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n41), .A1(n40), .A2(n39), .A3(n38), .Z(n42));
Q_MX08 U137 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][8] ), .A1(\mem_a[25][8] ), .A2(\mem_a[26][8] ), .A3(\mem_a[27][8] ), .A4(\mem_a[28][8] ), .A5(\mem_a[29][8] ), .A6(\mem_a[30][8] ), .A7(\mem_a[31][8] ), .Z(n43));
Q_MX08 U138 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][8] ), .A1(\mem_a[17][8] ), .A2(\mem_a[18][8] ), .A3(\mem_a[19][8] ), .A4(\mem_a[20][8] ), .A5(\mem_a[21][8] ), .A6(\mem_a[22][8] ), .A7(\mem_a[23][8] ), .Z(n44));
Q_MX08 U139 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][8] ), .A1(\mem_a[9][8] ), .A2(\mem_a[10][8] ), .A3(\mem_a[11][8] ), .A4(\mem_a[12][8] ), .A5(\mem_a[13][8] ), .A6(\mem_a[14][8] ), .A7(\mem_a[15][8] ), .Z(n45));
Q_MX08 U140 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][8] ), .A1(\mem_a[1][8] ), .A2(\mem_a[2][8] ), .A3(\mem_a[3][8] ), .A4(\mem_a[4][8] ), .A5(\mem_a[5][8] ), .A6(\mem_a[6][8] ), .A7(\mem_a[7][8] ), .Z(n46));
Q_MX04 U141 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n46), .A1(n45), .A2(n44), .A3(n43), .Z(n47));
Q_MX08 U142 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][9] ), .A1(\mem_a[25][9] ), .A2(\mem_a[26][9] ), .A3(\mem_a[27][9] ), .A4(\mem_a[28][9] ), .A5(\mem_a[29][9] ), .A6(\mem_a[30][9] ), .A7(\mem_a[31][9] ), .Z(n48));
Q_MX08 U143 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][9] ), .A1(\mem_a[17][9] ), .A2(\mem_a[18][9] ), .A3(\mem_a[19][9] ), .A4(\mem_a[20][9] ), .A5(\mem_a[21][9] ), .A6(\mem_a[22][9] ), .A7(\mem_a[23][9] ), .Z(n49));
Q_MX08 U144 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][9] ), .A1(\mem_a[9][9] ), .A2(\mem_a[10][9] ), .A3(\mem_a[11][9] ), .A4(\mem_a[12][9] ), .A5(\mem_a[13][9] ), .A6(\mem_a[14][9] ), .A7(\mem_a[15][9] ), .Z(n50));
Q_MX08 U145 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][9] ), .A1(\mem_a[1][9] ), .A2(\mem_a[2][9] ), .A3(\mem_a[3][9] ), .A4(\mem_a[4][9] ), .A5(\mem_a[5][9] ), .A6(\mem_a[6][9] ), .A7(\mem_a[7][9] ), .Z(n51));
Q_MX04 U146 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n51), .A1(n50), .A2(n49), .A3(n48), .Z(n52));
Q_MX08 U147 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][10] ), .A1(\mem_a[25][10] ), .A2(\mem_a[26][10] ), .A3(\mem_a[27][10] ), .A4(\mem_a[28][10] ), .A5(\mem_a[29][10] ), .A6(\mem_a[30][10] ), .A7(\mem_a[31][10] ), .Z(n53));
Q_MX08 U148 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][10] ), .A1(\mem_a[17][10] ), .A2(\mem_a[18][10] ), .A3(\mem_a[19][10] ), .A4(\mem_a[20][10] ), .A5(\mem_a[21][10] ), .A6(\mem_a[22][10] ), .A7(\mem_a[23][10] ), .Z(n54));
Q_MX08 U149 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][10] ), .A1(\mem_a[9][10] ), .A2(\mem_a[10][10] ), .A3(\mem_a[11][10] ), .A4(\mem_a[12][10] ), .A5(\mem_a[13][10] ), .A6(\mem_a[14][10] ), .A7(\mem_a[15][10] ), .Z(n55));
Q_MX08 U150 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][10] ), .A1(\mem_a[1][10] ), .A2(\mem_a[2][10] ), .A3(\mem_a[3][10] ), .A4(\mem_a[4][10] ), .A5(\mem_a[5][10] ), .A6(\mem_a[6][10] ), .A7(\mem_a[7][10] ), .Z(n56));
Q_MX04 U151 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n56), .A1(n55), .A2(n54), .A3(n53), .Z(n57));
Q_MX08 U152 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][11] ), .A1(\mem_a[25][11] ), .A2(\mem_a[26][11] ), .A3(\mem_a[27][11] ), .A4(\mem_a[28][11] ), .A5(\mem_a[29][11] ), .A6(\mem_a[30][11] ), .A7(\mem_a[31][11] ), .Z(n58));
Q_MX08 U153 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][11] ), .A1(\mem_a[17][11] ), .A2(\mem_a[18][11] ), .A3(\mem_a[19][11] ), .A4(\mem_a[20][11] ), .A5(\mem_a[21][11] ), .A6(\mem_a[22][11] ), .A7(\mem_a[23][11] ), .Z(n59));
Q_MX08 U154 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][11] ), .A1(\mem_a[9][11] ), .A2(\mem_a[10][11] ), .A3(\mem_a[11][11] ), .A4(\mem_a[12][11] ), .A5(\mem_a[13][11] ), .A6(\mem_a[14][11] ), .A7(\mem_a[15][11] ), .Z(n60));
Q_MX08 U155 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][11] ), .A1(\mem_a[1][11] ), .A2(\mem_a[2][11] ), .A3(\mem_a[3][11] ), .A4(\mem_a[4][11] ), .A5(\mem_a[5][11] ), .A6(\mem_a[6][11] ), .A7(\mem_a[7][11] ), .Z(n61));
Q_MX04 U156 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n61), .A1(n60), .A2(n59), .A3(n58), .Z(n62));
Q_MX08 U157 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][12] ), .A1(\mem_a[25][12] ), .A2(\mem_a[26][12] ), .A3(\mem_a[27][12] ), .A4(\mem_a[28][12] ), .A5(\mem_a[29][12] ), .A6(\mem_a[30][12] ), .A7(\mem_a[31][12] ), .Z(n63));
Q_MX08 U158 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][12] ), .A1(\mem_a[17][12] ), .A2(\mem_a[18][12] ), .A3(\mem_a[19][12] ), .A4(\mem_a[20][12] ), .A5(\mem_a[21][12] ), .A6(\mem_a[22][12] ), .A7(\mem_a[23][12] ), .Z(n64));
Q_MX08 U159 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][12] ), .A1(\mem_a[9][12] ), .A2(\mem_a[10][12] ), .A3(\mem_a[11][12] ), .A4(\mem_a[12][12] ), .A5(\mem_a[13][12] ), .A6(\mem_a[14][12] ), .A7(\mem_a[15][12] ), .Z(n65));
Q_MX08 U160 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][12] ), .A1(\mem_a[1][12] ), .A2(\mem_a[2][12] ), .A3(\mem_a[3][12] ), .A4(\mem_a[4][12] ), .A5(\mem_a[5][12] ), .A6(\mem_a[6][12] ), .A7(\mem_a[7][12] ), .Z(n66));
Q_MX04 U161 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n66), .A1(n65), .A2(n64), .A3(n63), .Z(n67));
Q_MX08 U162 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][13] ), .A1(\mem_a[25][13] ), .A2(\mem_a[26][13] ), .A3(\mem_a[27][13] ), .A4(\mem_a[28][13] ), .A5(\mem_a[29][13] ), .A6(\mem_a[30][13] ), .A7(\mem_a[31][13] ), .Z(n68));
Q_MX08 U163 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][13] ), .A1(\mem_a[17][13] ), .A2(\mem_a[18][13] ), .A3(\mem_a[19][13] ), .A4(\mem_a[20][13] ), .A5(\mem_a[21][13] ), .A6(\mem_a[22][13] ), .A7(\mem_a[23][13] ), .Z(n69));
Q_MX08 U164 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][13] ), .A1(\mem_a[9][13] ), .A2(\mem_a[10][13] ), .A3(\mem_a[11][13] ), .A4(\mem_a[12][13] ), .A5(\mem_a[13][13] ), .A6(\mem_a[14][13] ), .A7(\mem_a[15][13] ), .Z(n70));
Q_MX08 U165 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][13] ), .A1(\mem_a[1][13] ), .A2(\mem_a[2][13] ), .A3(\mem_a[3][13] ), .A4(\mem_a[4][13] ), .A5(\mem_a[5][13] ), .A6(\mem_a[6][13] ), .A7(\mem_a[7][13] ), .Z(n71));
Q_MX04 U166 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n71), .A1(n70), .A2(n69), .A3(n68), .Z(n72));
Q_MX08 U167 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][14] ), .A1(\mem_a[25][14] ), .A2(\mem_a[26][14] ), .A3(\mem_a[27][14] ), .A4(\mem_a[28][14] ), .A5(\mem_a[29][14] ), .A6(\mem_a[30][14] ), .A7(\mem_a[31][14] ), .Z(n73));
Q_MX08 U168 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][14] ), .A1(\mem_a[17][14] ), .A2(\mem_a[18][14] ), .A3(\mem_a[19][14] ), .A4(\mem_a[20][14] ), .A5(\mem_a[21][14] ), .A6(\mem_a[22][14] ), .A7(\mem_a[23][14] ), .Z(n74));
Q_MX08 U169 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][14] ), .A1(\mem_a[9][14] ), .A2(\mem_a[10][14] ), .A3(\mem_a[11][14] ), .A4(\mem_a[12][14] ), .A5(\mem_a[13][14] ), .A6(\mem_a[14][14] ), .A7(\mem_a[15][14] ), .Z(n75));
Q_MX08 U170 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][14] ), .A1(\mem_a[1][14] ), .A2(\mem_a[2][14] ), .A3(\mem_a[3][14] ), .A4(\mem_a[4][14] ), .A5(\mem_a[5][14] ), .A6(\mem_a[6][14] ), .A7(\mem_a[7][14] ), .Z(n76));
Q_MX04 U171 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n76), .A1(n75), .A2(n74), .A3(n73), .Z(n77));
Q_MX08 U172 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][15] ), .A1(\mem_a[25][15] ), .A2(\mem_a[26][15] ), .A3(\mem_a[27][15] ), .A4(\mem_a[28][15] ), .A5(\mem_a[29][15] ), .A6(\mem_a[30][15] ), .A7(\mem_a[31][15] ), .Z(n78));
Q_MX08 U173 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][15] ), .A1(\mem_a[17][15] ), .A2(\mem_a[18][15] ), .A3(\mem_a[19][15] ), .A4(\mem_a[20][15] ), .A5(\mem_a[21][15] ), .A6(\mem_a[22][15] ), .A7(\mem_a[23][15] ), .Z(n79));
Q_MX08 U174 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][15] ), .A1(\mem_a[9][15] ), .A2(\mem_a[10][15] ), .A3(\mem_a[11][15] ), .A4(\mem_a[12][15] ), .A5(\mem_a[13][15] ), .A6(\mem_a[14][15] ), .A7(\mem_a[15][15] ), .Z(n80));
Q_MX08 U175 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][15] ), .A1(\mem_a[1][15] ), .A2(\mem_a[2][15] ), .A3(\mem_a[3][15] ), .A4(\mem_a[4][15] ), .A5(\mem_a[5][15] ), .A6(\mem_a[6][15] ), .A7(\mem_a[7][15] ), .Z(n81));
Q_MX04 U176 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n81), .A1(n80), .A2(n79), .A3(n78), .Z(n82));
Q_MX08 U177 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][16] ), .A1(\mem_a[25][16] ), .A2(\mem_a[26][16] ), .A3(\mem_a[27][16] ), .A4(\mem_a[28][16] ), .A5(\mem_a[29][16] ), .A6(\mem_a[30][16] ), .A7(\mem_a[31][16] ), .Z(n83));
Q_MX08 U178 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][16] ), .A1(\mem_a[17][16] ), .A2(\mem_a[18][16] ), .A3(\mem_a[19][16] ), .A4(\mem_a[20][16] ), .A5(\mem_a[21][16] ), .A6(\mem_a[22][16] ), .A7(\mem_a[23][16] ), .Z(n84));
Q_MX08 U179 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][16] ), .A1(\mem_a[9][16] ), .A2(\mem_a[10][16] ), .A3(\mem_a[11][16] ), .A4(\mem_a[12][16] ), .A5(\mem_a[13][16] ), .A6(\mem_a[14][16] ), .A7(\mem_a[15][16] ), .Z(n85));
Q_MX08 U180 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][16] ), .A1(\mem_a[1][16] ), .A2(\mem_a[2][16] ), .A3(\mem_a[3][16] ), .A4(\mem_a[4][16] ), .A5(\mem_a[5][16] ), .A6(\mem_a[6][16] ), .A7(\mem_a[7][16] ), .Z(n86));
Q_MX04 U181 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n86), .A1(n85), .A2(n84), .A3(n83), .Z(n87));
Q_MX08 U182 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][17] ), .A1(\mem_a[25][17] ), .A2(\mem_a[26][17] ), .A3(\mem_a[27][17] ), .A4(\mem_a[28][17] ), .A5(\mem_a[29][17] ), .A6(\mem_a[30][17] ), .A7(\mem_a[31][17] ), .Z(n88));
Q_MX08 U183 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][17] ), .A1(\mem_a[17][17] ), .A2(\mem_a[18][17] ), .A3(\mem_a[19][17] ), .A4(\mem_a[20][17] ), .A5(\mem_a[21][17] ), .A6(\mem_a[22][17] ), .A7(\mem_a[23][17] ), .Z(n89));
Q_MX08 U184 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][17] ), .A1(\mem_a[9][17] ), .A2(\mem_a[10][17] ), .A3(\mem_a[11][17] ), .A4(\mem_a[12][17] ), .A5(\mem_a[13][17] ), .A6(\mem_a[14][17] ), .A7(\mem_a[15][17] ), .Z(n90));
Q_MX08 U185 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][17] ), .A1(\mem_a[1][17] ), .A2(\mem_a[2][17] ), .A3(\mem_a[3][17] ), .A4(\mem_a[4][17] ), .A5(\mem_a[5][17] ), .A6(\mem_a[6][17] ), .A7(\mem_a[7][17] ), .Z(n91));
Q_MX04 U186 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n91), .A1(n90), .A2(n89), .A3(n88), .Z(n92));
Q_MX08 U187 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][18] ), .A1(\mem_a[25][18] ), .A2(\mem_a[26][18] ), .A3(\mem_a[27][18] ), .A4(\mem_a[28][18] ), .A5(\mem_a[29][18] ), .A6(\mem_a[30][18] ), .A7(\mem_a[31][18] ), .Z(n93));
Q_MX08 U188 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][18] ), .A1(\mem_a[17][18] ), .A2(\mem_a[18][18] ), .A3(\mem_a[19][18] ), .A4(\mem_a[20][18] ), .A5(\mem_a[21][18] ), .A6(\mem_a[22][18] ), .A7(\mem_a[23][18] ), .Z(n94));
Q_MX08 U189 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][18] ), .A1(\mem_a[9][18] ), .A2(\mem_a[10][18] ), .A3(\mem_a[11][18] ), .A4(\mem_a[12][18] ), .A5(\mem_a[13][18] ), .A6(\mem_a[14][18] ), .A7(\mem_a[15][18] ), .Z(n95));
Q_MX08 U190 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][18] ), .A1(\mem_a[1][18] ), .A2(\mem_a[2][18] ), .A3(\mem_a[3][18] ), .A4(\mem_a[4][18] ), .A5(\mem_a[5][18] ), .A6(\mem_a[6][18] ), .A7(\mem_a[7][18] ), .Z(n96));
Q_MX04 U191 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n96), .A1(n95), .A2(n94), .A3(n93), .Z(n97));
Q_MX08 U192 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][19] ), .A1(\mem_a[25][19] ), .A2(\mem_a[26][19] ), .A3(\mem_a[27][19] ), .A4(\mem_a[28][19] ), .A5(\mem_a[29][19] ), .A6(\mem_a[30][19] ), .A7(\mem_a[31][19] ), .Z(n98));
Q_MX08 U193 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][19] ), .A1(\mem_a[17][19] ), .A2(\mem_a[18][19] ), .A3(\mem_a[19][19] ), .A4(\mem_a[20][19] ), .A5(\mem_a[21][19] ), .A6(\mem_a[22][19] ), .A7(\mem_a[23][19] ), .Z(n99));
Q_MX08 U194 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][19] ), .A1(\mem_a[9][19] ), .A2(\mem_a[10][19] ), .A3(\mem_a[11][19] ), .A4(\mem_a[12][19] ), .A5(\mem_a[13][19] ), .A6(\mem_a[14][19] ), .A7(\mem_a[15][19] ), .Z(n100));
Q_MX08 U195 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][19] ), .A1(\mem_a[1][19] ), .A2(\mem_a[2][19] ), .A3(\mem_a[3][19] ), .A4(\mem_a[4][19] ), .A5(\mem_a[5][19] ), .A6(\mem_a[6][19] ), .A7(\mem_a[7][19] ), .Z(n101));
Q_MX04 U196 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n101), .A1(n100), .A2(n99), .A3(n98), .Z(n102));
Q_MX08 U197 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][20] ), .A1(\mem_a[25][20] ), .A2(\mem_a[26][20] ), .A3(\mem_a[27][20] ), .A4(\mem_a[28][20] ), .A5(\mem_a[29][20] ), .A6(\mem_a[30][20] ), .A7(\mem_a[31][20] ), .Z(n103));
Q_MX08 U198 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][20] ), .A1(\mem_a[17][20] ), .A2(\mem_a[18][20] ), .A3(\mem_a[19][20] ), .A4(\mem_a[20][20] ), .A5(\mem_a[21][20] ), .A6(\mem_a[22][20] ), .A7(\mem_a[23][20] ), .Z(n104));
Q_MX08 U199 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][20] ), .A1(\mem_a[9][20] ), .A2(\mem_a[10][20] ), .A3(\mem_a[11][20] ), .A4(\mem_a[12][20] ), .A5(\mem_a[13][20] ), .A6(\mem_a[14][20] ), .A7(\mem_a[15][20] ), .Z(n105));
Q_MX08 U200 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][20] ), .A1(\mem_a[1][20] ), .A2(\mem_a[2][20] ), .A3(\mem_a[3][20] ), .A4(\mem_a[4][20] ), .A5(\mem_a[5][20] ), .A6(\mem_a[6][20] ), .A7(\mem_a[7][20] ), .Z(n106));
Q_MX04 U201 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n106), .A1(n105), .A2(n104), .A3(n103), .Z(n107));
Q_MX08 U202 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][21] ), .A1(\mem_a[25][21] ), .A2(\mem_a[26][21] ), .A3(\mem_a[27][21] ), .A4(\mem_a[28][21] ), .A5(\mem_a[29][21] ), .A6(\mem_a[30][21] ), .A7(\mem_a[31][21] ), .Z(n108));
Q_MX08 U203 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][21] ), .A1(\mem_a[17][21] ), .A2(\mem_a[18][21] ), .A3(\mem_a[19][21] ), .A4(\mem_a[20][21] ), .A5(\mem_a[21][21] ), .A6(\mem_a[22][21] ), .A7(\mem_a[23][21] ), .Z(n109));
Q_MX08 U204 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][21] ), .A1(\mem_a[9][21] ), .A2(\mem_a[10][21] ), .A3(\mem_a[11][21] ), .A4(\mem_a[12][21] ), .A5(\mem_a[13][21] ), .A6(\mem_a[14][21] ), .A7(\mem_a[15][21] ), .Z(n110));
Q_MX08 U205 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][21] ), .A1(\mem_a[1][21] ), .A2(\mem_a[2][21] ), .A3(\mem_a[3][21] ), .A4(\mem_a[4][21] ), .A5(\mem_a[5][21] ), .A6(\mem_a[6][21] ), .A7(\mem_a[7][21] ), .Z(n111));
Q_MX04 U206 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n111), .A1(n110), .A2(n109), .A3(n108), .Z(n112));
Q_MX08 U207 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][22] ), .A1(\mem_a[25][22] ), .A2(\mem_a[26][22] ), .A3(\mem_a[27][22] ), .A4(\mem_a[28][22] ), .A5(\mem_a[29][22] ), .A6(\mem_a[30][22] ), .A7(\mem_a[31][22] ), .Z(n113));
Q_MX08 U208 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][22] ), .A1(\mem_a[17][22] ), .A2(\mem_a[18][22] ), .A3(\mem_a[19][22] ), .A4(\mem_a[20][22] ), .A5(\mem_a[21][22] ), .A6(\mem_a[22][22] ), .A7(\mem_a[23][22] ), .Z(n114));
Q_MX08 U209 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][22] ), .A1(\mem_a[9][22] ), .A2(\mem_a[10][22] ), .A3(\mem_a[11][22] ), .A4(\mem_a[12][22] ), .A5(\mem_a[13][22] ), .A6(\mem_a[14][22] ), .A7(\mem_a[15][22] ), .Z(n115));
Q_MX08 U210 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][22] ), .A1(\mem_a[1][22] ), .A2(\mem_a[2][22] ), .A3(\mem_a[3][22] ), .A4(\mem_a[4][22] ), .A5(\mem_a[5][22] ), .A6(\mem_a[6][22] ), .A7(\mem_a[7][22] ), .Z(n116));
Q_MX04 U211 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n116), .A1(n115), .A2(n114), .A3(n113), .Z(n117));
Q_MX08 U212 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][23] ), .A1(\mem_a[25][23] ), .A2(\mem_a[26][23] ), .A3(\mem_a[27][23] ), .A4(\mem_a[28][23] ), .A5(\mem_a[29][23] ), .A6(\mem_a[30][23] ), .A7(\mem_a[31][23] ), .Z(n118));
Q_MX08 U213 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][23] ), .A1(\mem_a[17][23] ), .A2(\mem_a[18][23] ), .A3(\mem_a[19][23] ), .A4(\mem_a[20][23] ), .A5(\mem_a[21][23] ), .A6(\mem_a[22][23] ), .A7(\mem_a[23][23] ), .Z(n119));
Q_MX08 U214 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][23] ), .A1(\mem_a[9][23] ), .A2(\mem_a[10][23] ), .A3(\mem_a[11][23] ), .A4(\mem_a[12][23] ), .A5(\mem_a[13][23] ), .A6(\mem_a[14][23] ), .A7(\mem_a[15][23] ), .Z(n120));
Q_MX08 U215 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][23] ), .A1(\mem_a[1][23] ), .A2(\mem_a[2][23] ), .A3(\mem_a[3][23] ), .A4(\mem_a[4][23] ), .A5(\mem_a[5][23] ), .A6(\mem_a[6][23] ), .A7(\mem_a[7][23] ), .Z(n121));
Q_MX04 U216 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n121), .A1(n120), .A2(n119), .A3(n118), .Z(n122));
Q_MX08 U217 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][24] ), .A1(\mem_a[25][24] ), .A2(\mem_a[26][24] ), .A3(\mem_a[27][24] ), .A4(\mem_a[28][24] ), .A5(\mem_a[29][24] ), .A6(\mem_a[30][24] ), .A7(\mem_a[31][24] ), .Z(n123));
Q_MX08 U218 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][24] ), .A1(\mem_a[17][24] ), .A2(\mem_a[18][24] ), .A3(\mem_a[19][24] ), .A4(\mem_a[20][24] ), .A5(\mem_a[21][24] ), .A6(\mem_a[22][24] ), .A7(\mem_a[23][24] ), .Z(n124));
Q_MX08 U219 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][24] ), .A1(\mem_a[9][24] ), .A2(\mem_a[10][24] ), .A3(\mem_a[11][24] ), .A4(\mem_a[12][24] ), .A5(\mem_a[13][24] ), .A6(\mem_a[14][24] ), .A7(\mem_a[15][24] ), .Z(n125));
Q_MX08 U220 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][24] ), .A1(\mem_a[1][24] ), .A2(\mem_a[2][24] ), .A3(\mem_a[3][24] ), .A4(\mem_a[4][24] ), .A5(\mem_a[5][24] ), .A6(\mem_a[6][24] ), .A7(\mem_a[7][24] ), .Z(n126));
Q_MX04 U221 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n126), .A1(n125), .A2(n124), .A3(n123), .Z(n127));
Q_MX08 U222 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][25] ), .A1(\mem_a[25][25] ), .A2(\mem_a[26][25] ), .A3(\mem_a[27][25] ), .A4(\mem_a[28][25] ), .A5(\mem_a[29][25] ), .A6(\mem_a[30][25] ), .A7(\mem_a[31][25] ), .Z(n128));
Q_MX08 U223 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][25] ), .A1(\mem_a[17][25] ), .A2(\mem_a[18][25] ), .A3(\mem_a[19][25] ), .A4(\mem_a[20][25] ), .A5(\mem_a[21][25] ), .A6(\mem_a[22][25] ), .A7(\mem_a[23][25] ), .Z(n129));
Q_MX08 U224 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][25] ), .A1(\mem_a[9][25] ), .A2(\mem_a[10][25] ), .A3(\mem_a[11][25] ), .A4(\mem_a[12][25] ), .A5(\mem_a[13][25] ), .A6(\mem_a[14][25] ), .A7(\mem_a[15][25] ), .Z(n130));
Q_MX08 U225 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][25] ), .A1(\mem_a[1][25] ), .A2(\mem_a[2][25] ), .A3(\mem_a[3][25] ), .A4(\mem_a[4][25] ), .A5(\mem_a[5][25] ), .A6(\mem_a[6][25] ), .A7(\mem_a[7][25] ), .Z(n131));
Q_MX04 U226 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n131), .A1(n130), .A2(n129), .A3(n128), .Z(n132));
Q_MX08 U227 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][26] ), .A1(\mem_a[25][26] ), .A2(\mem_a[26][26] ), .A3(\mem_a[27][26] ), .A4(\mem_a[28][26] ), .A5(\mem_a[29][26] ), .A6(\mem_a[30][26] ), .A7(\mem_a[31][26] ), .Z(n133));
Q_MX08 U228 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][26] ), .A1(\mem_a[17][26] ), .A2(\mem_a[18][26] ), .A3(\mem_a[19][26] ), .A4(\mem_a[20][26] ), .A5(\mem_a[21][26] ), .A6(\mem_a[22][26] ), .A7(\mem_a[23][26] ), .Z(n134));
Q_MX08 U229 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][26] ), .A1(\mem_a[9][26] ), .A2(\mem_a[10][26] ), .A3(\mem_a[11][26] ), .A4(\mem_a[12][26] ), .A5(\mem_a[13][26] ), .A6(\mem_a[14][26] ), .A7(\mem_a[15][26] ), .Z(n135));
Q_MX08 U230 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][26] ), .A1(\mem_a[1][26] ), .A2(\mem_a[2][26] ), .A3(\mem_a[3][26] ), .A4(\mem_a[4][26] ), .A5(\mem_a[5][26] ), .A6(\mem_a[6][26] ), .A7(\mem_a[7][26] ), .Z(n136));
Q_MX04 U231 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n136), .A1(n135), .A2(n134), .A3(n133), .Z(n137));
Q_MX08 U232 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][27] ), .A1(\mem_a[25][27] ), .A2(\mem_a[26][27] ), .A3(\mem_a[27][27] ), .A4(\mem_a[28][27] ), .A5(\mem_a[29][27] ), .A6(\mem_a[30][27] ), .A7(\mem_a[31][27] ), .Z(n138));
Q_MX08 U233 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][27] ), .A1(\mem_a[17][27] ), .A2(\mem_a[18][27] ), .A3(\mem_a[19][27] ), .A4(\mem_a[20][27] ), .A5(\mem_a[21][27] ), .A6(\mem_a[22][27] ), .A7(\mem_a[23][27] ), .Z(n139));
Q_MX08 U234 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][27] ), .A1(\mem_a[9][27] ), .A2(\mem_a[10][27] ), .A3(\mem_a[11][27] ), .A4(\mem_a[12][27] ), .A5(\mem_a[13][27] ), .A6(\mem_a[14][27] ), .A7(\mem_a[15][27] ), .Z(n140));
Q_MX08 U235 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][27] ), .A1(\mem_a[1][27] ), .A2(\mem_a[2][27] ), .A3(\mem_a[3][27] ), .A4(\mem_a[4][27] ), .A5(\mem_a[5][27] ), .A6(\mem_a[6][27] ), .A7(\mem_a[7][27] ), .Z(n141));
Q_MX04 U236 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n141), .A1(n140), .A2(n139), .A3(n138), .Z(n142));
Q_MX08 U237 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][28] ), .A1(\mem_a[25][28] ), .A2(\mem_a[26][28] ), .A3(\mem_a[27][28] ), .A4(\mem_a[28][28] ), .A5(\mem_a[29][28] ), .A6(\mem_a[30][28] ), .A7(\mem_a[31][28] ), .Z(n143));
Q_MX08 U238 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][28] ), .A1(\mem_a[17][28] ), .A2(\mem_a[18][28] ), .A3(\mem_a[19][28] ), .A4(\mem_a[20][28] ), .A5(\mem_a[21][28] ), .A6(\mem_a[22][28] ), .A7(\mem_a[23][28] ), .Z(n144));
Q_MX08 U239 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][28] ), .A1(\mem_a[9][28] ), .A2(\mem_a[10][28] ), .A3(\mem_a[11][28] ), .A4(\mem_a[12][28] ), .A5(\mem_a[13][28] ), .A6(\mem_a[14][28] ), .A7(\mem_a[15][28] ), .Z(n145));
Q_MX08 U240 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][28] ), .A1(\mem_a[1][28] ), .A2(\mem_a[2][28] ), .A3(\mem_a[3][28] ), .A4(\mem_a[4][28] ), .A5(\mem_a[5][28] ), .A6(\mem_a[6][28] ), .A7(\mem_a[7][28] ), .Z(n146));
Q_MX04 U241 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n146), .A1(n145), .A2(n144), .A3(n143), .Z(n147));
Q_MX08 U242 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][29] ), .A1(\mem_a[25][29] ), .A2(\mem_a[26][29] ), .A3(\mem_a[27][29] ), .A4(\mem_a[28][29] ), .A5(\mem_a[29][29] ), .A6(\mem_a[30][29] ), .A7(\mem_a[31][29] ), .Z(n148));
Q_MX08 U243 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][29] ), .A1(\mem_a[17][29] ), .A2(\mem_a[18][29] ), .A3(\mem_a[19][29] ), .A4(\mem_a[20][29] ), .A5(\mem_a[21][29] ), .A6(\mem_a[22][29] ), .A7(\mem_a[23][29] ), .Z(n149));
Q_MX08 U244 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][29] ), .A1(\mem_a[9][29] ), .A2(\mem_a[10][29] ), .A3(\mem_a[11][29] ), .A4(\mem_a[12][29] ), .A5(\mem_a[13][29] ), .A6(\mem_a[14][29] ), .A7(\mem_a[15][29] ), .Z(n150));
Q_MX08 U245 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][29] ), .A1(\mem_a[1][29] ), .A2(\mem_a[2][29] ), .A3(\mem_a[3][29] ), .A4(\mem_a[4][29] ), .A5(\mem_a[5][29] ), .A6(\mem_a[6][29] ), .A7(\mem_a[7][29] ), .Z(n151));
Q_MX04 U246 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n151), .A1(n150), .A2(n149), .A3(n148), .Z(n152));
Q_MX08 U247 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][30] ), .A1(\mem_a[25][30] ), .A2(\mem_a[26][30] ), .A3(\mem_a[27][30] ), .A4(\mem_a[28][30] ), .A5(\mem_a[29][30] ), .A6(\mem_a[30][30] ), .A7(\mem_a[31][30] ), .Z(n153));
Q_MX08 U248 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][30] ), .A1(\mem_a[17][30] ), .A2(\mem_a[18][30] ), .A3(\mem_a[19][30] ), .A4(\mem_a[20][30] ), .A5(\mem_a[21][30] ), .A6(\mem_a[22][30] ), .A7(\mem_a[23][30] ), .Z(n154));
Q_MX08 U249 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][30] ), .A1(\mem_a[9][30] ), .A2(\mem_a[10][30] ), .A3(\mem_a[11][30] ), .A4(\mem_a[12][30] ), .A5(\mem_a[13][30] ), .A6(\mem_a[14][30] ), .A7(\mem_a[15][30] ), .Z(n155));
Q_MX08 U250 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][30] ), .A1(\mem_a[1][30] ), .A2(\mem_a[2][30] ), .A3(\mem_a[3][30] ), .A4(\mem_a[4][30] ), .A5(\mem_a[5][30] ), .A6(\mem_a[6][30] ), .A7(\mem_a[7][30] ), .Z(n156));
Q_MX04 U251 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n156), .A1(n155), .A2(n154), .A3(n153), .Z(n157));
Q_MX08 U252 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][31] ), .A1(\mem_a[25][31] ), .A2(\mem_a[26][31] ), .A3(\mem_a[27][31] ), .A4(\mem_a[28][31] ), .A5(\mem_a[29][31] ), .A6(\mem_a[30][31] ), .A7(\mem_a[31][31] ), .Z(n158));
Q_MX08 U253 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][31] ), .A1(\mem_a[17][31] ), .A2(\mem_a[18][31] ), .A3(\mem_a[19][31] ), .A4(\mem_a[20][31] ), .A5(\mem_a[21][31] ), .A6(\mem_a[22][31] ), .A7(\mem_a[23][31] ), .Z(n159));
Q_MX08 U254 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][31] ), .A1(\mem_a[9][31] ), .A2(\mem_a[10][31] ), .A3(\mem_a[11][31] ), .A4(\mem_a[12][31] ), .A5(\mem_a[13][31] ), .A6(\mem_a[14][31] ), .A7(\mem_a[15][31] ), .Z(n160));
Q_MX08 U255 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][31] ), .A1(\mem_a[1][31] ), .A2(\mem_a[2][31] ), .A3(\mem_a[3][31] ), .A4(\mem_a[4][31] ), .A5(\mem_a[5][31] ), .A6(\mem_a[6][31] ), .A7(\mem_a[7][31] ), .Z(n161));
Q_MX04 U256 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n161), .A1(n160), .A2(n159), .A3(n158), .Z(n162));
Q_MX08 U257 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][32] ), .A1(\mem_a[25][32] ), .A2(\mem_a[26][32] ), .A3(\mem_a[27][32] ), .A4(\mem_a[28][32] ), .A5(\mem_a[29][32] ), .A6(\mem_a[30][32] ), .A7(\mem_a[31][32] ), .Z(n163));
Q_MX08 U258 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][32] ), .A1(\mem_a[17][32] ), .A2(\mem_a[18][32] ), .A3(\mem_a[19][32] ), .A4(\mem_a[20][32] ), .A5(\mem_a[21][32] ), .A6(\mem_a[22][32] ), .A7(\mem_a[23][32] ), .Z(n164));
Q_MX08 U259 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][32] ), .A1(\mem_a[9][32] ), .A2(\mem_a[10][32] ), .A3(\mem_a[11][32] ), .A4(\mem_a[12][32] ), .A5(\mem_a[13][32] ), .A6(\mem_a[14][32] ), .A7(\mem_a[15][32] ), .Z(n165));
Q_MX08 U260 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][32] ), .A1(\mem_a[1][32] ), .A2(\mem_a[2][32] ), .A3(\mem_a[3][32] ), .A4(\mem_a[4][32] ), .A5(\mem_a[5][32] ), .A6(\mem_a[6][32] ), .A7(\mem_a[7][32] ), .Z(n166));
Q_MX04 U261 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n166), .A1(n165), .A2(n164), .A3(n163), .Z(n167));
Q_MX08 U262 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][33] ), .A1(\mem_a[25][33] ), .A2(\mem_a[26][33] ), .A3(\mem_a[27][33] ), .A4(\mem_a[28][33] ), .A5(\mem_a[29][33] ), .A6(\mem_a[30][33] ), .A7(\mem_a[31][33] ), .Z(n168));
Q_MX08 U263 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][33] ), .A1(\mem_a[17][33] ), .A2(\mem_a[18][33] ), .A3(\mem_a[19][33] ), .A4(\mem_a[20][33] ), .A5(\mem_a[21][33] ), .A6(\mem_a[22][33] ), .A7(\mem_a[23][33] ), .Z(n169));
Q_MX08 U264 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][33] ), .A1(\mem_a[9][33] ), .A2(\mem_a[10][33] ), .A3(\mem_a[11][33] ), .A4(\mem_a[12][33] ), .A5(\mem_a[13][33] ), .A6(\mem_a[14][33] ), .A7(\mem_a[15][33] ), .Z(n170));
Q_MX08 U265 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][33] ), .A1(\mem_a[1][33] ), .A2(\mem_a[2][33] ), .A3(\mem_a[3][33] ), .A4(\mem_a[4][33] ), .A5(\mem_a[5][33] ), .A6(\mem_a[6][33] ), .A7(\mem_a[7][33] ), .Z(n171));
Q_MX04 U266 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n171), .A1(n170), .A2(n169), .A3(n168), .Z(n172));
Q_MX08 U267 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][34] ), .A1(\mem_a[25][34] ), .A2(\mem_a[26][34] ), .A3(\mem_a[27][34] ), .A4(\mem_a[28][34] ), .A5(\mem_a[29][34] ), .A6(\mem_a[30][34] ), .A7(\mem_a[31][34] ), .Z(n173));
Q_MX08 U268 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][34] ), .A1(\mem_a[17][34] ), .A2(\mem_a[18][34] ), .A3(\mem_a[19][34] ), .A4(\mem_a[20][34] ), .A5(\mem_a[21][34] ), .A6(\mem_a[22][34] ), .A7(\mem_a[23][34] ), .Z(n174));
Q_MX08 U269 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][34] ), .A1(\mem_a[9][34] ), .A2(\mem_a[10][34] ), .A3(\mem_a[11][34] ), .A4(\mem_a[12][34] ), .A5(\mem_a[13][34] ), .A6(\mem_a[14][34] ), .A7(\mem_a[15][34] ), .Z(n175));
Q_MX08 U270 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][34] ), .A1(\mem_a[1][34] ), .A2(\mem_a[2][34] ), .A3(\mem_a[3][34] ), .A4(\mem_a[4][34] ), .A5(\mem_a[5][34] ), .A6(\mem_a[6][34] ), .A7(\mem_a[7][34] ), .Z(n176));
Q_MX04 U271 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n176), .A1(n175), .A2(n174), .A3(n173), .Z(n177));
Q_MX08 U272 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][35] ), .A1(\mem_a[25][35] ), .A2(\mem_a[26][35] ), .A3(\mem_a[27][35] ), .A4(\mem_a[28][35] ), .A5(\mem_a[29][35] ), .A6(\mem_a[30][35] ), .A7(\mem_a[31][35] ), .Z(n178));
Q_MX08 U273 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][35] ), .A1(\mem_a[17][35] ), .A2(\mem_a[18][35] ), .A3(\mem_a[19][35] ), .A4(\mem_a[20][35] ), .A5(\mem_a[21][35] ), .A6(\mem_a[22][35] ), .A7(\mem_a[23][35] ), .Z(n179));
Q_MX08 U274 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][35] ), .A1(\mem_a[9][35] ), .A2(\mem_a[10][35] ), .A3(\mem_a[11][35] ), .A4(\mem_a[12][35] ), .A5(\mem_a[13][35] ), .A6(\mem_a[14][35] ), .A7(\mem_a[15][35] ), .Z(n180));
Q_MX08 U275 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][35] ), .A1(\mem_a[1][35] ), .A2(\mem_a[2][35] ), .A3(\mem_a[3][35] ), .A4(\mem_a[4][35] ), .A5(\mem_a[5][35] ), .A6(\mem_a[6][35] ), .A7(\mem_a[7][35] ), .Z(n181));
Q_MX04 U276 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n181), .A1(n180), .A2(n179), .A3(n178), .Z(n182));
Q_MX08 U277 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][36] ), .A1(\mem_a[25][36] ), .A2(\mem_a[26][36] ), .A3(\mem_a[27][36] ), .A4(\mem_a[28][36] ), .A5(\mem_a[29][36] ), .A6(\mem_a[30][36] ), .A7(\mem_a[31][36] ), .Z(n183));
Q_MX08 U278 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][36] ), .A1(\mem_a[17][36] ), .A2(\mem_a[18][36] ), .A3(\mem_a[19][36] ), .A4(\mem_a[20][36] ), .A5(\mem_a[21][36] ), .A6(\mem_a[22][36] ), .A7(\mem_a[23][36] ), .Z(n184));
Q_MX08 U279 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][36] ), .A1(\mem_a[9][36] ), .A2(\mem_a[10][36] ), .A3(\mem_a[11][36] ), .A4(\mem_a[12][36] ), .A5(\mem_a[13][36] ), .A6(\mem_a[14][36] ), .A7(\mem_a[15][36] ), .Z(n185));
Q_MX08 U280 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][36] ), .A1(\mem_a[1][36] ), .A2(\mem_a[2][36] ), .A3(\mem_a[3][36] ), .A4(\mem_a[4][36] ), .A5(\mem_a[5][36] ), .A6(\mem_a[6][36] ), .A7(\mem_a[7][36] ), .Z(n186));
Q_MX04 U281 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n186), .A1(n185), .A2(n184), .A3(n183), .Z(n187));
Q_MX08 U282 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][37] ), .A1(\mem_a[25][37] ), .A2(\mem_a[26][37] ), .A3(\mem_a[27][37] ), .A4(\mem_a[28][37] ), .A5(\mem_a[29][37] ), .A6(\mem_a[30][37] ), .A7(\mem_a[31][37] ), .Z(n188));
Q_MX08 U283 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][37] ), .A1(\mem_a[17][37] ), .A2(\mem_a[18][37] ), .A3(\mem_a[19][37] ), .A4(\mem_a[20][37] ), .A5(\mem_a[21][37] ), .A6(\mem_a[22][37] ), .A7(\mem_a[23][37] ), .Z(n189));
Q_MX08 U284 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][37] ), .A1(\mem_a[9][37] ), .A2(\mem_a[10][37] ), .A3(\mem_a[11][37] ), .A4(\mem_a[12][37] ), .A5(\mem_a[13][37] ), .A6(\mem_a[14][37] ), .A7(\mem_a[15][37] ), .Z(n190));
Q_MX08 U285 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][37] ), .A1(\mem_a[1][37] ), .A2(\mem_a[2][37] ), .A3(\mem_a[3][37] ), .A4(\mem_a[4][37] ), .A5(\mem_a[5][37] ), .A6(\mem_a[6][37] ), .A7(\mem_a[7][37] ), .Z(n191));
Q_MX04 U286 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n191), .A1(n190), .A2(n189), .A3(n188), .Z(n192));
Q_MX08 U287 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][38] ), .A1(\mem_a[25][38] ), .A2(\mem_a[26][38] ), .A3(\mem_a[27][38] ), .A4(\mem_a[28][38] ), .A5(\mem_a[29][38] ), .A6(\mem_a[30][38] ), .A7(\mem_a[31][38] ), .Z(n193));
Q_MX08 U288 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][38] ), .A1(\mem_a[17][38] ), .A2(\mem_a[18][38] ), .A3(\mem_a[19][38] ), .A4(\mem_a[20][38] ), .A5(\mem_a[21][38] ), .A6(\mem_a[22][38] ), .A7(\mem_a[23][38] ), .Z(n194));
Q_MX08 U289 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][38] ), .A1(\mem_a[9][38] ), .A2(\mem_a[10][38] ), .A3(\mem_a[11][38] ), .A4(\mem_a[12][38] ), .A5(\mem_a[13][38] ), .A6(\mem_a[14][38] ), .A7(\mem_a[15][38] ), .Z(n195));
Q_MX08 U290 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][38] ), .A1(\mem_a[1][38] ), .A2(\mem_a[2][38] ), .A3(\mem_a[3][38] ), .A4(\mem_a[4][38] ), .A5(\mem_a[5][38] ), .A6(\mem_a[6][38] ), .A7(\mem_a[7][38] ), .Z(n196));
Q_MX04 U291 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n196), .A1(n195), .A2(n194), .A3(n193), .Z(n197));
Q_MX08 U292 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][39] ), .A1(\mem_a[25][39] ), .A2(\mem_a[26][39] ), .A3(\mem_a[27][39] ), .A4(\mem_a[28][39] ), .A5(\mem_a[29][39] ), .A6(\mem_a[30][39] ), .A7(\mem_a[31][39] ), .Z(n198));
Q_MX08 U293 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][39] ), .A1(\mem_a[17][39] ), .A2(\mem_a[18][39] ), .A3(\mem_a[19][39] ), .A4(\mem_a[20][39] ), .A5(\mem_a[21][39] ), .A6(\mem_a[22][39] ), .A7(\mem_a[23][39] ), .Z(n199));
Q_MX08 U294 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][39] ), .A1(\mem_a[9][39] ), .A2(\mem_a[10][39] ), .A3(\mem_a[11][39] ), .A4(\mem_a[12][39] ), .A5(\mem_a[13][39] ), .A6(\mem_a[14][39] ), .A7(\mem_a[15][39] ), .Z(n200));
Q_MX08 U295 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][39] ), .A1(\mem_a[1][39] ), .A2(\mem_a[2][39] ), .A3(\mem_a[3][39] ), .A4(\mem_a[4][39] ), .A5(\mem_a[5][39] ), .A6(\mem_a[6][39] ), .A7(\mem_a[7][39] ), .Z(n201));
Q_MX04 U296 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n201), .A1(n200), .A2(n199), .A3(n198), .Z(n202));
Q_MX08 U297 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][40] ), .A1(\mem_a[25][40] ), .A2(\mem_a[26][40] ), .A3(\mem_a[27][40] ), .A4(\mem_a[28][40] ), .A5(\mem_a[29][40] ), .A6(\mem_a[30][40] ), .A7(\mem_a[31][40] ), .Z(n203));
Q_MX08 U298 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][40] ), .A1(\mem_a[17][40] ), .A2(\mem_a[18][40] ), .A3(\mem_a[19][40] ), .A4(\mem_a[20][40] ), .A5(\mem_a[21][40] ), .A6(\mem_a[22][40] ), .A7(\mem_a[23][40] ), .Z(n204));
Q_MX08 U299 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][40] ), .A1(\mem_a[9][40] ), .A2(\mem_a[10][40] ), .A3(\mem_a[11][40] ), .A4(\mem_a[12][40] ), .A5(\mem_a[13][40] ), .A6(\mem_a[14][40] ), .A7(\mem_a[15][40] ), .Z(n205));
Q_MX08 U300 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][40] ), .A1(\mem_a[1][40] ), .A2(\mem_a[2][40] ), .A3(\mem_a[3][40] ), .A4(\mem_a[4][40] ), .A5(\mem_a[5][40] ), .A6(\mem_a[6][40] ), .A7(\mem_a[7][40] ), .Z(n206));
Q_MX04 U301 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n206), .A1(n205), .A2(n204), .A3(n203), .Z(n207));
Q_MX08 U302 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][41] ), .A1(\mem_a[25][41] ), .A2(\mem_a[26][41] ), .A3(\mem_a[27][41] ), .A4(\mem_a[28][41] ), .A5(\mem_a[29][41] ), .A6(\mem_a[30][41] ), .A7(\mem_a[31][41] ), .Z(n208));
Q_MX08 U303 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][41] ), .A1(\mem_a[17][41] ), .A2(\mem_a[18][41] ), .A3(\mem_a[19][41] ), .A4(\mem_a[20][41] ), .A5(\mem_a[21][41] ), .A6(\mem_a[22][41] ), .A7(\mem_a[23][41] ), .Z(n209));
Q_MX08 U304 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][41] ), .A1(\mem_a[9][41] ), .A2(\mem_a[10][41] ), .A3(\mem_a[11][41] ), .A4(\mem_a[12][41] ), .A5(\mem_a[13][41] ), .A6(\mem_a[14][41] ), .A7(\mem_a[15][41] ), .Z(n210));
Q_MX08 U305 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][41] ), .A1(\mem_a[1][41] ), .A2(\mem_a[2][41] ), .A3(\mem_a[3][41] ), .A4(\mem_a[4][41] ), .A5(\mem_a[5][41] ), .A6(\mem_a[6][41] ), .A7(\mem_a[7][41] ), .Z(n211));
Q_MX04 U306 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n211), .A1(n210), .A2(n209), .A3(n208), .Z(n212));
Q_MX08 U307 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][42] ), .A1(\mem_a[25][42] ), .A2(\mem_a[26][42] ), .A3(\mem_a[27][42] ), .A4(\mem_a[28][42] ), .A5(\mem_a[29][42] ), .A6(\mem_a[30][42] ), .A7(\mem_a[31][42] ), .Z(n213));
Q_MX08 U308 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][42] ), .A1(\mem_a[17][42] ), .A2(\mem_a[18][42] ), .A3(\mem_a[19][42] ), .A4(\mem_a[20][42] ), .A5(\mem_a[21][42] ), .A6(\mem_a[22][42] ), .A7(\mem_a[23][42] ), .Z(n214));
Q_MX08 U309 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][42] ), .A1(\mem_a[9][42] ), .A2(\mem_a[10][42] ), .A3(\mem_a[11][42] ), .A4(\mem_a[12][42] ), .A5(\mem_a[13][42] ), .A6(\mem_a[14][42] ), .A7(\mem_a[15][42] ), .Z(n215));
Q_MX08 U310 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][42] ), .A1(\mem_a[1][42] ), .A2(\mem_a[2][42] ), .A3(\mem_a[3][42] ), .A4(\mem_a[4][42] ), .A5(\mem_a[5][42] ), .A6(\mem_a[6][42] ), .A7(\mem_a[7][42] ), .Z(n216));
Q_MX04 U311 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n216), .A1(n215), .A2(n214), .A3(n213), .Z(n217));
Q_MX08 U312 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][43] ), .A1(\mem_a[25][43] ), .A2(\mem_a[26][43] ), .A3(\mem_a[27][43] ), .A4(\mem_a[28][43] ), .A5(\mem_a[29][43] ), .A6(\mem_a[30][43] ), .A7(\mem_a[31][43] ), .Z(n218));
Q_MX08 U313 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][43] ), .A1(\mem_a[17][43] ), .A2(\mem_a[18][43] ), .A3(\mem_a[19][43] ), .A4(\mem_a[20][43] ), .A5(\mem_a[21][43] ), .A6(\mem_a[22][43] ), .A7(\mem_a[23][43] ), .Z(n219));
Q_MX08 U314 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][43] ), .A1(\mem_a[9][43] ), .A2(\mem_a[10][43] ), .A3(\mem_a[11][43] ), .A4(\mem_a[12][43] ), .A5(\mem_a[13][43] ), .A6(\mem_a[14][43] ), .A7(\mem_a[15][43] ), .Z(n220));
Q_MX08 U315 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][43] ), .A1(\mem_a[1][43] ), .A2(\mem_a[2][43] ), .A3(\mem_a[3][43] ), .A4(\mem_a[4][43] ), .A5(\mem_a[5][43] ), .A6(\mem_a[6][43] ), .A7(\mem_a[7][43] ), .Z(n221));
Q_MX04 U316 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n221), .A1(n220), .A2(n219), .A3(n218), .Z(n222));
Q_MX08 U317 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][44] ), .A1(\mem_a[25][44] ), .A2(\mem_a[26][44] ), .A3(\mem_a[27][44] ), .A4(\mem_a[28][44] ), .A5(\mem_a[29][44] ), .A6(\mem_a[30][44] ), .A7(\mem_a[31][44] ), .Z(n223));
Q_MX08 U318 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][44] ), .A1(\mem_a[17][44] ), .A2(\mem_a[18][44] ), .A3(\mem_a[19][44] ), .A4(\mem_a[20][44] ), .A5(\mem_a[21][44] ), .A6(\mem_a[22][44] ), .A7(\mem_a[23][44] ), .Z(n224));
Q_MX08 U319 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][44] ), .A1(\mem_a[9][44] ), .A2(\mem_a[10][44] ), .A3(\mem_a[11][44] ), .A4(\mem_a[12][44] ), .A5(\mem_a[13][44] ), .A6(\mem_a[14][44] ), .A7(\mem_a[15][44] ), .Z(n225));
Q_MX08 U320 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][44] ), .A1(\mem_a[1][44] ), .A2(\mem_a[2][44] ), .A3(\mem_a[3][44] ), .A4(\mem_a[4][44] ), .A5(\mem_a[5][44] ), .A6(\mem_a[6][44] ), .A7(\mem_a[7][44] ), .Z(n226));
Q_MX04 U321 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n226), .A1(n225), .A2(n224), .A3(n223), .Z(n227));
Q_MX08 U322 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][45] ), .A1(\mem_a[25][45] ), .A2(\mem_a[26][45] ), .A3(\mem_a[27][45] ), .A4(\mem_a[28][45] ), .A5(\mem_a[29][45] ), .A6(\mem_a[30][45] ), .A7(\mem_a[31][45] ), .Z(n228));
Q_MX08 U323 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][45] ), .A1(\mem_a[17][45] ), .A2(\mem_a[18][45] ), .A3(\mem_a[19][45] ), .A4(\mem_a[20][45] ), .A5(\mem_a[21][45] ), .A6(\mem_a[22][45] ), .A7(\mem_a[23][45] ), .Z(n229));
Q_MX08 U324 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][45] ), .A1(\mem_a[9][45] ), .A2(\mem_a[10][45] ), .A3(\mem_a[11][45] ), .A4(\mem_a[12][45] ), .A5(\mem_a[13][45] ), .A6(\mem_a[14][45] ), .A7(\mem_a[15][45] ), .Z(n230));
Q_MX08 U325 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][45] ), .A1(\mem_a[1][45] ), .A2(\mem_a[2][45] ), .A3(\mem_a[3][45] ), .A4(\mem_a[4][45] ), .A5(\mem_a[5][45] ), .A6(\mem_a[6][45] ), .A7(\mem_a[7][45] ), .Z(n231));
Q_MX04 U326 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n231), .A1(n230), .A2(n229), .A3(n228), .Z(n232));
Q_MX08 U327 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][46] ), .A1(\mem_a[25][46] ), .A2(\mem_a[26][46] ), .A3(\mem_a[27][46] ), .A4(\mem_a[28][46] ), .A5(\mem_a[29][46] ), .A6(\mem_a[30][46] ), .A7(\mem_a[31][46] ), .Z(n233));
Q_MX08 U328 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][46] ), .A1(\mem_a[17][46] ), .A2(\mem_a[18][46] ), .A3(\mem_a[19][46] ), .A4(\mem_a[20][46] ), .A5(\mem_a[21][46] ), .A6(\mem_a[22][46] ), .A7(\mem_a[23][46] ), .Z(n234));
Q_MX08 U329 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][46] ), .A1(\mem_a[9][46] ), .A2(\mem_a[10][46] ), .A3(\mem_a[11][46] ), .A4(\mem_a[12][46] ), .A5(\mem_a[13][46] ), .A6(\mem_a[14][46] ), .A7(\mem_a[15][46] ), .Z(n235));
Q_MX08 U330 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][46] ), .A1(\mem_a[1][46] ), .A2(\mem_a[2][46] ), .A3(\mem_a[3][46] ), .A4(\mem_a[4][46] ), .A5(\mem_a[5][46] ), .A6(\mem_a[6][46] ), .A7(\mem_a[7][46] ), .Z(n236));
Q_MX04 U331 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n236), .A1(n235), .A2(n234), .A3(n233), .Z(n237));
Q_MX08 U332 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][47] ), .A1(\mem_a[25][47] ), .A2(\mem_a[26][47] ), .A3(\mem_a[27][47] ), .A4(\mem_a[28][47] ), .A5(\mem_a[29][47] ), .A6(\mem_a[30][47] ), .A7(\mem_a[31][47] ), .Z(n238));
Q_MX08 U333 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][47] ), .A1(\mem_a[17][47] ), .A2(\mem_a[18][47] ), .A3(\mem_a[19][47] ), .A4(\mem_a[20][47] ), .A5(\mem_a[21][47] ), .A6(\mem_a[22][47] ), .A7(\mem_a[23][47] ), .Z(n239));
Q_MX08 U334 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][47] ), .A1(\mem_a[9][47] ), .A2(\mem_a[10][47] ), .A3(\mem_a[11][47] ), .A4(\mem_a[12][47] ), .A5(\mem_a[13][47] ), .A6(\mem_a[14][47] ), .A7(\mem_a[15][47] ), .Z(n240));
Q_MX08 U335 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][47] ), .A1(\mem_a[1][47] ), .A2(\mem_a[2][47] ), .A3(\mem_a[3][47] ), .A4(\mem_a[4][47] ), .A5(\mem_a[5][47] ), .A6(\mem_a[6][47] ), .A7(\mem_a[7][47] ), .Z(n241));
Q_MX04 U336 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n241), .A1(n240), .A2(n239), .A3(n238), .Z(n242));
Q_MX08 U337 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][48] ), .A1(\mem_a[25][48] ), .A2(\mem_a[26][48] ), .A3(\mem_a[27][48] ), .A4(\mem_a[28][48] ), .A5(\mem_a[29][48] ), .A6(\mem_a[30][48] ), .A7(\mem_a[31][48] ), .Z(n243));
Q_MX08 U338 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][48] ), .A1(\mem_a[17][48] ), .A2(\mem_a[18][48] ), .A3(\mem_a[19][48] ), .A4(\mem_a[20][48] ), .A5(\mem_a[21][48] ), .A6(\mem_a[22][48] ), .A7(\mem_a[23][48] ), .Z(n244));
Q_MX08 U339 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][48] ), .A1(\mem_a[9][48] ), .A2(\mem_a[10][48] ), .A3(\mem_a[11][48] ), .A4(\mem_a[12][48] ), .A5(\mem_a[13][48] ), .A6(\mem_a[14][48] ), .A7(\mem_a[15][48] ), .Z(n245));
Q_MX08 U340 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][48] ), .A1(\mem_a[1][48] ), .A2(\mem_a[2][48] ), .A3(\mem_a[3][48] ), .A4(\mem_a[4][48] ), .A5(\mem_a[5][48] ), .A6(\mem_a[6][48] ), .A7(\mem_a[7][48] ), .Z(n246));
Q_MX04 U341 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n246), .A1(n245), .A2(n244), .A3(n243), .Z(n247));
Q_MX08 U342 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][49] ), .A1(\mem_a[25][49] ), .A2(\mem_a[26][49] ), .A3(\mem_a[27][49] ), .A4(\mem_a[28][49] ), .A5(\mem_a[29][49] ), .A6(\mem_a[30][49] ), .A7(\mem_a[31][49] ), .Z(n248));
Q_MX08 U343 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][49] ), .A1(\mem_a[17][49] ), .A2(\mem_a[18][49] ), .A3(\mem_a[19][49] ), .A4(\mem_a[20][49] ), .A5(\mem_a[21][49] ), .A6(\mem_a[22][49] ), .A7(\mem_a[23][49] ), .Z(n249));
Q_MX08 U344 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][49] ), .A1(\mem_a[9][49] ), .A2(\mem_a[10][49] ), .A3(\mem_a[11][49] ), .A4(\mem_a[12][49] ), .A5(\mem_a[13][49] ), .A6(\mem_a[14][49] ), .A7(\mem_a[15][49] ), .Z(n250));
Q_MX08 U345 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][49] ), .A1(\mem_a[1][49] ), .A2(\mem_a[2][49] ), .A3(\mem_a[3][49] ), .A4(\mem_a[4][49] ), .A5(\mem_a[5][49] ), .A6(\mem_a[6][49] ), .A7(\mem_a[7][49] ), .Z(n251));
Q_MX04 U346 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n251), .A1(n250), .A2(n249), .A3(n248), .Z(n252));
Q_MX08 U347 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][50] ), .A1(\mem_a[25][50] ), .A2(\mem_a[26][50] ), .A3(\mem_a[27][50] ), .A4(\mem_a[28][50] ), .A5(\mem_a[29][50] ), .A6(\mem_a[30][50] ), .A7(\mem_a[31][50] ), .Z(n253));
Q_MX08 U348 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][50] ), .A1(\mem_a[17][50] ), .A2(\mem_a[18][50] ), .A3(\mem_a[19][50] ), .A4(\mem_a[20][50] ), .A5(\mem_a[21][50] ), .A6(\mem_a[22][50] ), .A7(\mem_a[23][50] ), .Z(n254));
Q_MX08 U349 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][50] ), .A1(\mem_a[9][50] ), .A2(\mem_a[10][50] ), .A3(\mem_a[11][50] ), .A4(\mem_a[12][50] ), .A5(\mem_a[13][50] ), .A6(\mem_a[14][50] ), .A7(\mem_a[15][50] ), .Z(n255));
Q_MX08 U350 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][50] ), .A1(\mem_a[1][50] ), .A2(\mem_a[2][50] ), .A3(\mem_a[3][50] ), .A4(\mem_a[4][50] ), .A5(\mem_a[5][50] ), .A6(\mem_a[6][50] ), .A7(\mem_a[7][50] ), .Z(n256));
Q_MX04 U351 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n256), .A1(n255), .A2(n254), .A3(n253), .Z(n257));
Q_MX08 U352 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][51] ), .A1(\mem_a[25][51] ), .A2(\mem_a[26][51] ), .A3(\mem_a[27][51] ), .A4(\mem_a[28][51] ), .A5(\mem_a[29][51] ), .A6(\mem_a[30][51] ), .A7(\mem_a[31][51] ), .Z(n258));
Q_MX08 U353 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][51] ), .A1(\mem_a[17][51] ), .A2(\mem_a[18][51] ), .A3(\mem_a[19][51] ), .A4(\mem_a[20][51] ), .A5(\mem_a[21][51] ), .A6(\mem_a[22][51] ), .A7(\mem_a[23][51] ), .Z(n259));
Q_MX08 U354 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][51] ), .A1(\mem_a[9][51] ), .A2(\mem_a[10][51] ), .A3(\mem_a[11][51] ), .A4(\mem_a[12][51] ), .A5(\mem_a[13][51] ), .A6(\mem_a[14][51] ), .A7(\mem_a[15][51] ), .Z(n260));
Q_MX08 U355 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][51] ), .A1(\mem_a[1][51] ), .A2(\mem_a[2][51] ), .A3(\mem_a[3][51] ), .A4(\mem_a[4][51] ), .A5(\mem_a[5][51] ), .A6(\mem_a[6][51] ), .A7(\mem_a[7][51] ), .Z(n261));
Q_MX04 U356 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n261), .A1(n260), .A2(n259), .A3(n258), .Z(n262));
Q_MX08 U357 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][52] ), .A1(\mem_a[25][52] ), .A2(\mem_a[26][52] ), .A3(\mem_a[27][52] ), .A4(\mem_a[28][52] ), .A5(\mem_a[29][52] ), .A6(\mem_a[30][52] ), .A7(\mem_a[31][52] ), .Z(n263));
Q_MX08 U358 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][52] ), .A1(\mem_a[17][52] ), .A2(\mem_a[18][52] ), .A3(\mem_a[19][52] ), .A4(\mem_a[20][52] ), .A5(\mem_a[21][52] ), .A6(\mem_a[22][52] ), .A7(\mem_a[23][52] ), .Z(n264));
Q_MX08 U359 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][52] ), .A1(\mem_a[9][52] ), .A2(\mem_a[10][52] ), .A3(\mem_a[11][52] ), .A4(\mem_a[12][52] ), .A5(\mem_a[13][52] ), .A6(\mem_a[14][52] ), .A7(\mem_a[15][52] ), .Z(n265));
Q_MX08 U360 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][52] ), .A1(\mem_a[1][52] ), .A2(\mem_a[2][52] ), .A3(\mem_a[3][52] ), .A4(\mem_a[4][52] ), .A5(\mem_a[5][52] ), .A6(\mem_a[6][52] ), .A7(\mem_a[7][52] ), .Z(n266));
Q_MX04 U361 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n266), .A1(n265), .A2(n264), .A3(n263), .Z(n267));
Q_MX08 U362 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][53] ), .A1(\mem_a[25][53] ), .A2(\mem_a[26][53] ), .A3(\mem_a[27][53] ), .A4(\mem_a[28][53] ), .A5(\mem_a[29][53] ), .A6(\mem_a[30][53] ), .A7(\mem_a[31][53] ), .Z(n268));
Q_MX08 U363 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][53] ), .A1(\mem_a[17][53] ), .A2(\mem_a[18][53] ), .A3(\mem_a[19][53] ), .A4(\mem_a[20][53] ), .A5(\mem_a[21][53] ), .A6(\mem_a[22][53] ), .A7(\mem_a[23][53] ), .Z(n269));
Q_MX08 U364 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][53] ), .A1(\mem_a[9][53] ), .A2(\mem_a[10][53] ), .A3(\mem_a[11][53] ), .A4(\mem_a[12][53] ), .A5(\mem_a[13][53] ), .A6(\mem_a[14][53] ), .A7(\mem_a[15][53] ), .Z(n270));
Q_MX08 U365 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][53] ), .A1(\mem_a[1][53] ), .A2(\mem_a[2][53] ), .A3(\mem_a[3][53] ), .A4(\mem_a[4][53] ), .A5(\mem_a[5][53] ), .A6(\mem_a[6][53] ), .A7(\mem_a[7][53] ), .Z(n271));
Q_MX04 U366 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n271), .A1(n270), .A2(n269), .A3(n268), .Z(n272));
Q_MX08 U367 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][54] ), .A1(\mem_a[25][54] ), .A2(\mem_a[26][54] ), .A3(\mem_a[27][54] ), .A4(\mem_a[28][54] ), .A5(\mem_a[29][54] ), .A6(\mem_a[30][54] ), .A7(\mem_a[31][54] ), .Z(n273));
Q_MX08 U368 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][54] ), .A1(\mem_a[17][54] ), .A2(\mem_a[18][54] ), .A3(\mem_a[19][54] ), .A4(\mem_a[20][54] ), .A5(\mem_a[21][54] ), .A6(\mem_a[22][54] ), .A7(\mem_a[23][54] ), .Z(n274));
Q_MX08 U369 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][54] ), .A1(\mem_a[9][54] ), .A2(\mem_a[10][54] ), .A3(\mem_a[11][54] ), .A4(\mem_a[12][54] ), .A5(\mem_a[13][54] ), .A6(\mem_a[14][54] ), .A7(\mem_a[15][54] ), .Z(n275));
Q_MX08 U370 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][54] ), .A1(\mem_a[1][54] ), .A2(\mem_a[2][54] ), .A3(\mem_a[3][54] ), .A4(\mem_a[4][54] ), .A5(\mem_a[5][54] ), .A6(\mem_a[6][54] ), .A7(\mem_a[7][54] ), .Z(n276));
Q_MX04 U371 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n276), .A1(n275), .A2(n274), .A3(n273), .Z(n277));
Q_MX08 U372 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][55] ), .A1(\mem_a[25][55] ), .A2(\mem_a[26][55] ), .A3(\mem_a[27][55] ), .A4(\mem_a[28][55] ), .A5(\mem_a[29][55] ), .A6(\mem_a[30][55] ), .A7(\mem_a[31][55] ), .Z(n278));
Q_MX08 U373 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][55] ), .A1(\mem_a[17][55] ), .A2(\mem_a[18][55] ), .A3(\mem_a[19][55] ), .A4(\mem_a[20][55] ), .A5(\mem_a[21][55] ), .A6(\mem_a[22][55] ), .A7(\mem_a[23][55] ), .Z(n279));
Q_MX08 U374 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][55] ), .A1(\mem_a[9][55] ), .A2(\mem_a[10][55] ), .A3(\mem_a[11][55] ), .A4(\mem_a[12][55] ), .A5(\mem_a[13][55] ), .A6(\mem_a[14][55] ), .A7(\mem_a[15][55] ), .Z(n280));
Q_MX08 U375 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][55] ), .A1(\mem_a[1][55] ), .A2(\mem_a[2][55] ), .A3(\mem_a[3][55] ), .A4(\mem_a[4][55] ), .A5(\mem_a[5][55] ), .A6(\mem_a[6][55] ), .A7(\mem_a[7][55] ), .Z(n281));
Q_MX04 U376 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n281), .A1(n280), .A2(n279), .A3(n278), .Z(n282));
Q_MX08 U377 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][56] ), .A1(\mem_a[25][56] ), .A2(\mem_a[26][56] ), .A3(\mem_a[27][56] ), .A4(\mem_a[28][56] ), .A5(\mem_a[29][56] ), .A6(\mem_a[30][56] ), .A7(\mem_a[31][56] ), .Z(n283));
Q_MX08 U378 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][56] ), .A1(\mem_a[17][56] ), .A2(\mem_a[18][56] ), .A3(\mem_a[19][56] ), .A4(\mem_a[20][56] ), .A5(\mem_a[21][56] ), .A6(\mem_a[22][56] ), .A7(\mem_a[23][56] ), .Z(n284));
Q_MX08 U379 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][56] ), .A1(\mem_a[9][56] ), .A2(\mem_a[10][56] ), .A3(\mem_a[11][56] ), .A4(\mem_a[12][56] ), .A5(\mem_a[13][56] ), .A6(\mem_a[14][56] ), .A7(\mem_a[15][56] ), .Z(n285));
Q_MX08 U380 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][56] ), .A1(\mem_a[1][56] ), .A2(\mem_a[2][56] ), .A3(\mem_a[3][56] ), .A4(\mem_a[4][56] ), .A5(\mem_a[5][56] ), .A6(\mem_a[6][56] ), .A7(\mem_a[7][56] ), .Z(n286));
Q_MX04 U381 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n286), .A1(n285), .A2(n284), .A3(n283), .Z(n287));
Q_MX08 U382 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][57] ), .A1(\mem_a[25][57] ), .A2(\mem_a[26][57] ), .A3(\mem_a[27][57] ), .A4(\mem_a[28][57] ), .A5(\mem_a[29][57] ), .A6(\mem_a[30][57] ), .A7(\mem_a[31][57] ), .Z(n288));
Q_MX08 U383 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][57] ), .A1(\mem_a[17][57] ), .A2(\mem_a[18][57] ), .A3(\mem_a[19][57] ), .A4(\mem_a[20][57] ), .A5(\mem_a[21][57] ), .A6(\mem_a[22][57] ), .A7(\mem_a[23][57] ), .Z(n289));
Q_MX08 U384 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][57] ), .A1(\mem_a[9][57] ), .A2(\mem_a[10][57] ), .A3(\mem_a[11][57] ), .A4(\mem_a[12][57] ), .A5(\mem_a[13][57] ), .A6(\mem_a[14][57] ), .A7(\mem_a[15][57] ), .Z(n290));
Q_MX08 U385 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][57] ), .A1(\mem_a[1][57] ), .A2(\mem_a[2][57] ), .A3(\mem_a[3][57] ), .A4(\mem_a[4][57] ), .A5(\mem_a[5][57] ), .A6(\mem_a[6][57] ), .A7(\mem_a[7][57] ), .Z(n291));
Q_MX04 U386 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n291), .A1(n290), .A2(n289), .A3(n288), .Z(n292));
Q_MX08 U387 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][58] ), .A1(\mem_a[25][58] ), .A2(\mem_a[26][58] ), .A3(\mem_a[27][58] ), .A4(\mem_a[28][58] ), .A5(\mem_a[29][58] ), .A6(\mem_a[30][58] ), .A7(\mem_a[31][58] ), .Z(n293));
Q_MX08 U388 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][58] ), .A1(\mem_a[17][58] ), .A2(\mem_a[18][58] ), .A3(\mem_a[19][58] ), .A4(\mem_a[20][58] ), .A5(\mem_a[21][58] ), .A6(\mem_a[22][58] ), .A7(\mem_a[23][58] ), .Z(n294));
Q_MX08 U389 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][58] ), .A1(\mem_a[9][58] ), .A2(\mem_a[10][58] ), .A3(\mem_a[11][58] ), .A4(\mem_a[12][58] ), .A5(\mem_a[13][58] ), .A6(\mem_a[14][58] ), .A7(\mem_a[15][58] ), .Z(n295));
Q_MX08 U390 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][58] ), .A1(\mem_a[1][58] ), .A2(\mem_a[2][58] ), .A3(\mem_a[3][58] ), .A4(\mem_a[4][58] ), .A5(\mem_a[5][58] ), .A6(\mem_a[6][58] ), .A7(\mem_a[7][58] ), .Z(n296));
Q_MX04 U391 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n296), .A1(n295), .A2(n294), .A3(n293), .Z(n297));
Q_MX08 U392 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][59] ), .A1(\mem_a[25][59] ), .A2(\mem_a[26][59] ), .A3(\mem_a[27][59] ), .A4(\mem_a[28][59] ), .A5(\mem_a[29][59] ), .A6(\mem_a[30][59] ), .A7(\mem_a[31][59] ), .Z(n298));
Q_MX08 U393 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][59] ), .A1(\mem_a[17][59] ), .A2(\mem_a[18][59] ), .A3(\mem_a[19][59] ), .A4(\mem_a[20][59] ), .A5(\mem_a[21][59] ), .A6(\mem_a[22][59] ), .A7(\mem_a[23][59] ), .Z(n299));
Q_MX08 U394 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][59] ), .A1(\mem_a[9][59] ), .A2(\mem_a[10][59] ), .A3(\mem_a[11][59] ), .A4(\mem_a[12][59] ), .A5(\mem_a[13][59] ), .A6(\mem_a[14][59] ), .A7(\mem_a[15][59] ), .Z(n300));
Q_MX08 U395 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][59] ), .A1(\mem_a[1][59] ), .A2(\mem_a[2][59] ), .A3(\mem_a[3][59] ), .A4(\mem_a[4][59] ), .A5(\mem_a[5][59] ), .A6(\mem_a[6][59] ), .A7(\mem_a[7][59] ), .Z(n301));
Q_MX04 U396 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n301), .A1(n300), .A2(n299), .A3(n298), .Z(n302));
Q_MX08 U397 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][60] ), .A1(\mem_a[25][60] ), .A2(\mem_a[26][60] ), .A3(\mem_a[27][60] ), .A4(\mem_a[28][60] ), .A5(\mem_a[29][60] ), .A6(\mem_a[30][60] ), .A7(\mem_a[31][60] ), .Z(n303));
Q_MX08 U398 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][60] ), .A1(\mem_a[17][60] ), .A2(\mem_a[18][60] ), .A3(\mem_a[19][60] ), .A4(\mem_a[20][60] ), .A5(\mem_a[21][60] ), .A6(\mem_a[22][60] ), .A7(\mem_a[23][60] ), .Z(n304));
Q_MX08 U399 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][60] ), .A1(\mem_a[9][60] ), .A2(\mem_a[10][60] ), .A3(\mem_a[11][60] ), .A4(\mem_a[12][60] ), .A5(\mem_a[13][60] ), .A6(\mem_a[14][60] ), .A7(\mem_a[15][60] ), .Z(n305));
Q_MX08 U400 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][60] ), .A1(\mem_a[1][60] ), .A2(\mem_a[2][60] ), .A3(\mem_a[3][60] ), .A4(\mem_a[4][60] ), .A5(\mem_a[5][60] ), .A6(\mem_a[6][60] ), .A7(\mem_a[7][60] ), .Z(n306));
Q_MX04 U401 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n306), .A1(n305), .A2(n304), .A3(n303), .Z(n307));
Q_MX08 U402 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][61] ), .A1(\mem_a[25][61] ), .A2(\mem_a[26][61] ), .A3(\mem_a[27][61] ), .A4(\mem_a[28][61] ), .A5(\mem_a[29][61] ), .A6(\mem_a[30][61] ), .A7(\mem_a[31][61] ), .Z(n308));
Q_MX08 U403 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][61] ), .A1(\mem_a[17][61] ), .A2(\mem_a[18][61] ), .A3(\mem_a[19][61] ), .A4(\mem_a[20][61] ), .A5(\mem_a[21][61] ), .A6(\mem_a[22][61] ), .A7(\mem_a[23][61] ), .Z(n309));
Q_MX08 U404 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][61] ), .A1(\mem_a[9][61] ), .A2(\mem_a[10][61] ), .A3(\mem_a[11][61] ), .A4(\mem_a[12][61] ), .A5(\mem_a[13][61] ), .A6(\mem_a[14][61] ), .A7(\mem_a[15][61] ), .Z(n310));
Q_MX08 U405 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][61] ), .A1(\mem_a[1][61] ), .A2(\mem_a[2][61] ), .A3(\mem_a[3][61] ), .A4(\mem_a[4][61] ), .A5(\mem_a[5][61] ), .A6(\mem_a[6][61] ), .A7(\mem_a[7][61] ), .Z(n311));
Q_MX04 U406 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n311), .A1(n310), .A2(n309), .A3(n308), .Z(n312));
Q_MX08 U407 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][62] ), .A1(\mem_a[25][62] ), .A2(\mem_a[26][62] ), .A3(\mem_a[27][62] ), .A4(\mem_a[28][62] ), .A5(\mem_a[29][62] ), .A6(\mem_a[30][62] ), .A7(\mem_a[31][62] ), .Z(n313));
Q_MX08 U408 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][62] ), .A1(\mem_a[17][62] ), .A2(\mem_a[18][62] ), .A3(\mem_a[19][62] ), .A4(\mem_a[20][62] ), .A5(\mem_a[21][62] ), .A6(\mem_a[22][62] ), .A7(\mem_a[23][62] ), .Z(n314));
Q_MX08 U409 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][62] ), .A1(\mem_a[9][62] ), .A2(\mem_a[10][62] ), .A3(\mem_a[11][62] ), .A4(\mem_a[12][62] ), .A5(\mem_a[13][62] ), .A6(\mem_a[14][62] ), .A7(\mem_a[15][62] ), .Z(n315));
Q_MX08 U410 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][62] ), .A1(\mem_a[1][62] ), .A2(\mem_a[2][62] ), .A3(\mem_a[3][62] ), .A4(\mem_a[4][62] ), .A5(\mem_a[5][62] ), .A6(\mem_a[6][62] ), .A7(\mem_a[7][62] ), .Z(n316));
Q_MX04 U411 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n316), .A1(n315), .A2(n314), .A3(n313), .Z(n317));
Q_MX08 U412 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[24][63] ), .A1(\mem_a[25][63] ), .A2(\mem_a[26][63] ), .A3(\mem_a[27][63] ), .A4(\mem_a[28][63] ), .A5(\mem_a[29][63] ), .A6(\mem_a[30][63] ), .A7(\mem_a[31][63] ), .Z(n318));
Q_MX08 U413 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[16][63] ), .A1(\mem_a[17][63] ), .A2(\mem_a[18][63] ), .A3(\mem_a[19][63] ), .A4(\mem_a[20][63] ), .A5(\mem_a[21][63] ), .A6(\mem_a[22][63] ), .A7(\mem_a[23][63] ), .Z(n319));
Q_MX08 U414 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[8][63] ), .A1(\mem_a[9][63] ), .A2(\mem_a[10][63] ), .A3(\mem_a[11][63] ), .A4(\mem_a[12][63] ), .A5(\mem_a[13][63] ), .A6(\mem_a[14][63] ), .A7(\mem_a[15][63] ), .Z(n320));
Q_MX08 U415 ( .S0(sw_add[0]), .S1(sw_add[1]), .S2(sw_add[2]), .A0(\mem_a[0][63] ), .A1(\mem_a[1][63] ), .A2(\mem_a[2][63] ), .A3(\mem_a[3][63] ), .A4(\mem_a[4][63] ), .A5(\mem_a[5][63] ), .A6(\mem_a[6][63] ), .A7(\mem_a[7][63] ), .Z(n321));
Q_MX04 U416 ( .S0(sw_add[3]), .S1(sw_add[4]), .A0(n321), .A1(n320), .A2(n319), .A3(n318), .Z(n322));
Q_ASSIGN U417 ( .B(\mem_a[0][0] ), .A(\_zyixc_ctx_rdata_29[0][0] ));
Q_ASSIGN U418 ( .B(\mem_a[0][1] ), .A(\_zyixc_ctx_rdata_29[0][1] ));
Q_ASSIGN U419 ( .B(\mem_a[0][2] ), .A(\_zyixc_ctx_rdata_29[0][2] ));
Q_ASSIGN U420 ( .B(\mem_a[0][3] ), .A(\_zyixc_ctx_rdata_29[0][3] ));
Q_ASSIGN U421 ( .B(\mem_a[0][4] ), .A(\_zyixc_ctx_rdata_29[0][4] ));
Q_ASSIGN U422 ( .B(\mem_a[0][5] ), .A(\_zyixc_ctx_rdata_29[0][5] ));
Q_ASSIGN U423 ( .B(\mem_a[0][6] ), .A(\_zyixc_ctx_rdata_29[0][6] ));
Q_ASSIGN U424 ( .B(\mem_a[0][7] ), .A(\_zyixc_ctx_rdata_29[0][7] ));
Q_ASSIGN U425 ( .B(\mem_a[0][8] ), .A(\_zyixc_ctx_rdata_29[0][8] ));
Q_ASSIGN U426 ( .B(\mem_a[0][9] ), .A(\_zyixc_ctx_rdata_29[0][9] ));
Q_ASSIGN U427 ( .B(\mem_a[0][10] ), .A(\_zyixc_ctx_rdata_29[0][10] ));
Q_ASSIGN U428 ( .B(\mem_a[0][11] ), .A(\_zyixc_ctx_rdata_29[0][11] ));
Q_ASSIGN U429 ( .B(\mem_a[0][12] ), .A(\_zyixc_ctx_rdata_29[0][12] ));
Q_ASSIGN U430 ( .B(\mem_a[0][13] ), .A(\_zyixc_ctx_rdata_29[0][13] ));
Q_ASSIGN U431 ( .B(\mem_a[0][14] ), .A(\_zyixc_ctx_rdata_29[0][14] ));
Q_ASSIGN U432 ( .B(\mem_a[0][15] ), .A(\_zyixc_ctx_rdata_29[0][15] ));
Q_ASSIGN U433 ( .B(\mem_a[0][16] ), .A(\_zyixc_ctx_rdata_29[0][16] ));
Q_ASSIGN U434 ( .B(\mem_a[0][17] ), .A(\_zyixc_ctx_rdata_29[0][17] ));
Q_ASSIGN U435 ( .B(\mem_a[0][18] ), .A(\_zyixc_ctx_rdata_29[0][18] ));
Q_ASSIGN U436 ( .B(\mem_a[0][19] ), .A(\_zyixc_ctx_rdata_29[0][19] ));
Q_ASSIGN U437 ( .B(\mem_a[0][20] ), .A(\_zyixc_ctx_rdata_29[0][20] ));
Q_ASSIGN U438 ( .B(\mem_a[0][21] ), .A(\_zyixc_ctx_rdata_29[0][21] ));
Q_ASSIGN U439 ( .B(\mem_a[0][22] ), .A(\_zyixc_ctx_rdata_29[0][22] ));
Q_ASSIGN U440 ( .B(\mem_a[0][23] ), .A(\_zyixc_ctx_rdata_29[0][23] ));
Q_ASSIGN U441 ( .B(\mem_a[0][24] ), .A(\_zyixc_ctx_rdata_29[0][24] ));
Q_ASSIGN U442 ( .B(\mem_a[0][25] ), .A(\_zyixc_ctx_rdata_29[0][25] ));
Q_ASSIGN U443 ( .B(\mem_a[0][26] ), .A(\_zyixc_ctx_rdata_29[0][26] ));
Q_ASSIGN U444 ( .B(\mem_a[0][27] ), .A(\_zyixc_ctx_rdata_29[0][27] ));
Q_ASSIGN U445 ( .B(\mem_a[0][28] ), .A(\_zyixc_ctx_rdata_29[0][28] ));
Q_ASSIGN U446 ( .B(\mem_a[0][29] ), .A(\_zyixc_ctx_rdata_29[0][29] ));
Q_ASSIGN U447 ( .B(\mem_a[0][30] ), .A(\_zyixc_ctx_rdata_29[0][30] ));
Q_ASSIGN U448 ( .B(\mem_a[0][31] ), .A(\_zyixc_ctx_rdata_29[0][31] ));
Q_ASSIGN U449 ( .B(\mem_a[0][32] ), .A(\_zyixc_ctx_rdata_29[0][32] ));
Q_ASSIGN U450 ( .B(\mem_a[0][33] ), .A(\_zyixc_ctx_rdata_29[0][33] ));
Q_ASSIGN U451 ( .B(\mem_a[0][34] ), .A(\_zyixc_ctx_rdata_29[0][34] ));
Q_ASSIGN U452 ( .B(\mem_a[0][35] ), .A(\_zyixc_ctx_rdata_29[0][35] ));
Q_ASSIGN U453 ( .B(\mem_a[0][36] ), .A(\_zyixc_ctx_rdata_29[0][36] ));
Q_ASSIGN U454 ( .B(\mem_a[0][37] ), .A(\_zyixc_ctx_rdata_29[0][37] ));
Q_ASSIGN U455 ( .B(\mem_a[0][38] ), .A(\_zyixc_ctx_rdata_29[0][38] ));
Q_ASSIGN U456 ( .B(\mem_a[0][39] ), .A(\_zyixc_ctx_rdata_29[0][39] ));
Q_ASSIGN U457 ( .B(\mem_a[0][40] ), .A(\_zyixc_ctx_rdata_29[0][40] ));
Q_ASSIGN U458 ( .B(\mem_a[0][41] ), .A(\_zyixc_ctx_rdata_29[0][41] ));
Q_ASSIGN U459 ( .B(\mem_a[0][42] ), .A(\_zyixc_ctx_rdata_29[0][42] ));
Q_ASSIGN U460 ( .B(\mem_a[0][43] ), .A(\_zyixc_ctx_rdata_29[0][43] ));
Q_ASSIGN U461 ( .B(\mem_a[0][44] ), .A(\_zyixc_ctx_rdata_29[0][44] ));
Q_ASSIGN U462 ( .B(\mem_a[0][45] ), .A(\_zyixc_ctx_rdata_29[0][45] ));
Q_ASSIGN U463 ( .B(\mem_a[0][46] ), .A(\_zyixc_ctx_rdata_29[0][46] ));
Q_ASSIGN U464 ( .B(\mem_a[0][47] ), .A(\_zyixc_ctx_rdata_29[0][47] ));
Q_ASSIGN U465 ( .B(\mem_a[0][48] ), .A(\_zyixc_ctx_rdata_29[0][48] ));
Q_ASSIGN U466 ( .B(\mem_a[0][49] ), .A(\_zyixc_ctx_rdata_29[0][49] ));
Q_ASSIGN U467 ( .B(\mem_a[0][50] ), .A(\_zyixc_ctx_rdata_29[0][50] ));
Q_ASSIGN U468 ( .B(\mem_a[0][51] ), .A(\_zyixc_ctx_rdata_29[0][51] ));
Q_ASSIGN U469 ( .B(\mem_a[0][52] ), .A(\_zyixc_ctx_rdata_29[0][52] ));
Q_ASSIGN U470 ( .B(\mem_a[0][53] ), .A(\_zyixc_ctx_rdata_29[0][53] ));
Q_ASSIGN U471 ( .B(\mem_a[0][54] ), .A(\_zyixc_ctx_rdata_29[0][54] ));
Q_ASSIGN U472 ( .B(\mem_a[0][55] ), .A(\_zyixc_ctx_rdata_29[0][55] ));
Q_ASSIGN U473 ( .B(\mem_a[0][56] ), .A(\_zyixc_ctx_rdata_29[0][56] ));
Q_ASSIGN U474 ( .B(\mem_a[0][57] ), .A(\_zyixc_ctx_rdata_29[0][57] ));
Q_ASSIGN U475 ( .B(\mem_a[0][58] ), .A(\_zyixc_ctx_rdata_29[0][58] ));
Q_ASSIGN U476 ( .B(\mem_a[0][59] ), .A(\_zyixc_ctx_rdata_29[0][59] ));
Q_ASSIGN U477 ( .B(\mem_a[0][60] ), .A(\_zyixc_ctx_rdata_29[0][60] ));
Q_ASSIGN U478 ( .B(\mem_a[0][61] ), .A(\_zyixc_ctx_rdata_29[0][61] ));
Q_ASSIGN U479 ( .B(\mem_a[0][62] ), .A(\_zyixc_ctx_rdata_29[0][62] ));
Q_ASSIGN U480 ( .B(\mem_a[0][63] ), .A(\_zyixc_ctx_rdata_29[0][63] ));
Q_ASSIGN U481 ( .B(\mem_a[1][0] ), .A(\_zyixc_ctx_rdata_29[1][0] ));
Q_ASSIGN U482 ( .B(\mem_a[1][1] ), .A(\_zyixc_ctx_rdata_29[1][1] ));
Q_ASSIGN U483 ( .B(\mem_a[1][2] ), .A(\_zyixc_ctx_rdata_29[1][2] ));
Q_ASSIGN U484 ( .B(\mem_a[1][3] ), .A(\_zyixc_ctx_rdata_29[1][3] ));
Q_ASSIGN U485 ( .B(\mem_a[1][4] ), .A(\_zyixc_ctx_rdata_29[1][4] ));
Q_ASSIGN U486 ( .B(\mem_a[1][5] ), .A(\_zyixc_ctx_rdata_29[1][5] ));
Q_ASSIGN U487 ( .B(\mem_a[1][6] ), .A(\_zyixc_ctx_rdata_29[1][6] ));
Q_ASSIGN U488 ( .B(\mem_a[1][7] ), .A(\_zyixc_ctx_rdata_29[1][7] ));
Q_ASSIGN U489 ( .B(\mem_a[1][8] ), .A(\_zyixc_ctx_rdata_29[1][8] ));
Q_ASSIGN U490 ( .B(\mem_a[1][9] ), .A(\_zyixc_ctx_rdata_29[1][9] ));
Q_ASSIGN U491 ( .B(\mem_a[1][10] ), .A(\_zyixc_ctx_rdata_29[1][10] ));
Q_ASSIGN U492 ( .B(\mem_a[1][11] ), .A(\_zyixc_ctx_rdata_29[1][11] ));
Q_ASSIGN U493 ( .B(\mem_a[1][12] ), .A(\_zyixc_ctx_rdata_29[1][12] ));
Q_ASSIGN U494 ( .B(\mem_a[1][13] ), .A(\_zyixc_ctx_rdata_29[1][13] ));
Q_ASSIGN U495 ( .B(\mem_a[1][14] ), .A(\_zyixc_ctx_rdata_29[1][14] ));
Q_ASSIGN U496 ( .B(\mem_a[1][15] ), .A(\_zyixc_ctx_rdata_29[1][15] ));
Q_ASSIGN U497 ( .B(\mem_a[1][16] ), .A(\_zyixc_ctx_rdata_29[1][16] ));
Q_ASSIGN U498 ( .B(\mem_a[1][17] ), .A(\_zyixc_ctx_rdata_29[1][17] ));
Q_ASSIGN U499 ( .B(\mem_a[1][18] ), .A(\_zyixc_ctx_rdata_29[1][18] ));
Q_ASSIGN U500 ( .B(\mem_a[1][19] ), .A(\_zyixc_ctx_rdata_29[1][19] ));
Q_ASSIGN U501 ( .B(\mem_a[1][20] ), .A(\_zyixc_ctx_rdata_29[1][20] ));
Q_ASSIGN U502 ( .B(\mem_a[1][21] ), .A(\_zyixc_ctx_rdata_29[1][21] ));
Q_ASSIGN U503 ( .B(\mem_a[1][22] ), .A(\_zyixc_ctx_rdata_29[1][22] ));
Q_ASSIGN U504 ( .B(\mem_a[1][23] ), .A(\_zyixc_ctx_rdata_29[1][23] ));
Q_ASSIGN U505 ( .B(\mem_a[1][24] ), .A(\_zyixc_ctx_rdata_29[1][24] ));
Q_ASSIGN U506 ( .B(\mem_a[1][25] ), .A(\_zyixc_ctx_rdata_29[1][25] ));
Q_ASSIGN U507 ( .B(\mem_a[1][26] ), .A(\_zyixc_ctx_rdata_29[1][26] ));
Q_ASSIGN U508 ( .B(\mem_a[1][27] ), .A(\_zyixc_ctx_rdata_29[1][27] ));
Q_ASSIGN U509 ( .B(\mem_a[1][28] ), .A(\_zyixc_ctx_rdata_29[1][28] ));
Q_ASSIGN U510 ( .B(\mem_a[1][29] ), .A(\_zyixc_ctx_rdata_29[1][29] ));
Q_ASSIGN U511 ( .B(\mem_a[1][30] ), .A(\_zyixc_ctx_rdata_29[1][30] ));
Q_ASSIGN U512 ( .B(\mem_a[1][31] ), .A(\_zyixc_ctx_rdata_29[1][31] ));
Q_ASSIGN U513 ( .B(\mem_a[1][32] ), .A(\_zyixc_ctx_rdata_29[1][32] ));
Q_ASSIGN U514 ( .B(\mem_a[1][33] ), .A(\_zyixc_ctx_rdata_29[1][33] ));
Q_ASSIGN U515 ( .B(\mem_a[1][34] ), .A(\_zyixc_ctx_rdata_29[1][34] ));
Q_ASSIGN U516 ( .B(\mem_a[1][35] ), .A(\_zyixc_ctx_rdata_29[1][35] ));
Q_ASSIGN U517 ( .B(\mem_a[1][36] ), .A(\_zyixc_ctx_rdata_29[1][36] ));
Q_ASSIGN U518 ( .B(\mem_a[1][37] ), .A(\_zyixc_ctx_rdata_29[1][37] ));
Q_ASSIGN U519 ( .B(\mem_a[1][38] ), .A(\_zyixc_ctx_rdata_29[1][38] ));
Q_ASSIGN U520 ( .B(\mem_a[1][39] ), .A(\_zyixc_ctx_rdata_29[1][39] ));
Q_ASSIGN U521 ( .B(\mem_a[1][40] ), .A(\_zyixc_ctx_rdata_29[1][40] ));
Q_ASSIGN U522 ( .B(\mem_a[1][41] ), .A(\_zyixc_ctx_rdata_29[1][41] ));
Q_ASSIGN U523 ( .B(\mem_a[1][42] ), .A(\_zyixc_ctx_rdata_29[1][42] ));
Q_ASSIGN U524 ( .B(\mem_a[1][43] ), .A(\_zyixc_ctx_rdata_29[1][43] ));
Q_ASSIGN U525 ( .B(\mem_a[1][44] ), .A(\_zyixc_ctx_rdata_29[1][44] ));
Q_ASSIGN U526 ( .B(\mem_a[1][45] ), .A(\_zyixc_ctx_rdata_29[1][45] ));
Q_ASSIGN U527 ( .B(\mem_a[1][46] ), .A(\_zyixc_ctx_rdata_29[1][46] ));
Q_ASSIGN U528 ( .B(\mem_a[1][47] ), .A(\_zyixc_ctx_rdata_29[1][47] ));
Q_ASSIGN U529 ( .B(\mem_a[1][48] ), .A(\_zyixc_ctx_rdata_29[1][48] ));
Q_ASSIGN U530 ( .B(\mem_a[1][49] ), .A(\_zyixc_ctx_rdata_29[1][49] ));
Q_ASSIGN U531 ( .B(\mem_a[1][50] ), .A(\_zyixc_ctx_rdata_29[1][50] ));
Q_ASSIGN U532 ( .B(\mem_a[1][51] ), .A(\_zyixc_ctx_rdata_29[1][51] ));
Q_ASSIGN U533 ( .B(\mem_a[1][52] ), .A(\_zyixc_ctx_rdata_29[1][52] ));
Q_ASSIGN U534 ( .B(\mem_a[1][53] ), .A(\_zyixc_ctx_rdata_29[1][53] ));
Q_ASSIGN U535 ( .B(\mem_a[1][54] ), .A(\_zyixc_ctx_rdata_29[1][54] ));
Q_ASSIGN U536 ( .B(\mem_a[1][55] ), .A(\_zyixc_ctx_rdata_29[1][55] ));
Q_ASSIGN U537 ( .B(\mem_a[1][56] ), .A(\_zyixc_ctx_rdata_29[1][56] ));
Q_ASSIGN U538 ( .B(\mem_a[1][57] ), .A(\_zyixc_ctx_rdata_29[1][57] ));
Q_ASSIGN U539 ( .B(\mem_a[1][58] ), .A(\_zyixc_ctx_rdata_29[1][58] ));
Q_ASSIGN U540 ( .B(\mem_a[1][59] ), .A(\_zyixc_ctx_rdata_29[1][59] ));
Q_ASSIGN U541 ( .B(\mem_a[1][60] ), .A(\_zyixc_ctx_rdata_29[1][60] ));
Q_ASSIGN U542 ( .B(\mem_a[1][61] ), .A(\_zyixc_ctx_rdata_29[1][61] ));
Q_ASSIGN U543 ( .B(\mem_a[1][62] ), .A(\_zyixc_ctx_rdata_29[1][62] ));
Q_ASSIGN U544 ( .B(\mem_a[1][63] ), .A(\_zyixc_ctx_rdata_29[1][63] ));
Q_ASSIGN U545 ( .B(\mem_a[2][0] ), .A(\_zyixc_ctx_rdata_29[2][0] ));
Q_ASSIGN U546 ( .B(\mem_a[2][1] ), .A(\_zyixc_ctx_rdata_29[2][1] ));
Q_ASSIGN U547 ( .B(\mem_a[2][2] ), .A(\_zyixc_ctx_rdata_29[2][2] ));
Q_ASSIGN U548 ( .B(\mem_a[2][3] ), .A(\_zyixc_ctx_rdata_29[2][3] ));
Q_ASSIGN U549 ( .B(\mem_a[2][4] ), .A(\_zyixc_ctx_rdata_29[2][4] ));
Q_ASSIGN U550 ( .B(\mem_a[2][5] ), .A(\_zyixc_ctx_rdata_29[2][5] ));
Q_ASSIGN U551 ( .B(\mem_a[2][6] ), .A(\_zyixc_ctx_rdata_29[2][6] ));
Q_ASSIGN U552 ( .B(\mem_a[2][7] ), .A(\_zyixc_ctx_rdata_29[2][7] ));
Q_ASSIGN U553 ( .B(\mem_a[2][8] ), .A(\_zyixc_ctx_rdata_29[2][8] ));
Q_ASSIGN U554 ( .B(\mem_a[2][9] ), .A(\_zyixc_ctx_rdata_29[2][9] ));
Q_ASSIGN U555 ( .B(\mem_a[2][10] ), .A(\_zyixc_ctx_rdata_29[2][10] ));
Q_ASSIGN U556 ( .B(\mem_a[2][11] ), .A(\_zyixc_ctx_rdata_29[2][11] ));
Q_ASSIGN U557 ( .B(\mem_a[2][12] ), .A(\_zyixc_ctx_rdata_29[2][12] ));
Q_ASSIGN U558 ( .B(\mem_a[2][13] ), .A(\_zyixc_ctx_rdata_29[2][13] ));
Q_ASSIGN U559 ( .B(\mem_a[2][14] ), .A(\_zyixc_ctx_rdata_29[2][14] ));
Q_ASSIGN U560 ( .B(\mem_a[2][15] ), .A(\_zyixc_ctx_rdata_29[2][15] ));
Q_ASSIGN U561 ( .B(\mem_a[2][16] ), .A(\_zyixc_ctx_rdata_29[2][16] ));
Q_ASSIGN U562 ( .B(\mem_a[2][17] ), .A(\_zyixc_ctx_rdata_29[2][17] ));
Q_ASSIGN U563 ( .B(\mem_a[2][18] ), .A(\_zyixc_ctx_rdata_29[2][18] ));
Q_ASSIGN U564 ( .B(\mem_a[2][19] ), .A(\_zyixc_ctx_rdata_29[2][19] ));
Q_ASSIGN U565 ( .B(\mem_a[2][20] ), .A(\_zyixc_ctx_rdata_29[2][20] ));
Q_ASSIGN U566 ( .B(\mem_a[2][21] ), .A(\_zyixc_ctx_rdata_29[2][21] ));
Q_ASSIGN U567 ( .B(\mem_a[2][22] ), .A(\_zyixc_ctx_rdata_29[2][22] ));
Q_ASSIGN U568 ( .B(\mem_a[2][23] ), .A(\_zyixc_ctx_rdata_29[2][23] ));
Q_ASSIGN U569 ( .B(\mem_a[2][24] ), .A(\_zyixc_ctx_rdata_29[2][24] ));
Q_ASSIGN U570 ( .B(\mem_a[2][25] ), .A(\_zyixc_ctx_rdata_29[2][25] ));
Q_ASSIGN U571 ( .B(\mem_a[2][26] ), .A(\_zyixc_ctx_rdata_29[2][26] ));
Q_ASSIGN U572 ( .B(\mem_a[2][27] ), .A(\_zyixc_ctx_rdata_29[2][27] ));
Q_ASSIGN U573 ( .B(\mem_a[2][28] ), .A(\_zyixc_ctx_rdata_29[2][28] ));
Q_ASSIGN U574 ( .B(\mem_a[2][29] ), .A(\_zyixc_ctx_rdata_29[2][29] ));
Q_ASSIGN U575 ( .B(\mem_a[2][30] ), .A(\_zyixc_ctx_rdata_29[2][30] ));
Q_ASSIGN U576 ( .B(\mem_a[2][31] ), .A(\_zyixc_ctx_rdata_29[2][31] ));
Q_ASSIGN U577 ( .B(\mem_a[2][32] ), .A(\_zyixc_ctx_rdata_29[2][32] ));
Q_ASSIGN U578 ( .B(\mem_a[2][33] ), .A(\_zyixc_ctx_rdata_29[2][33] ));
Q_ASSIGN U579 ( .B(\mem_a[2][34] ), .A(\_zyixc_ctx_rdata_29[2][34] ));
Q_ASSIGN U580 ( .B(\mem_a[2][35] ), .A(\_zyixc_ctx_rdata_29[2][35] ));
Q_ASSIGN U581 ( .B(\mem_a[2][36] ), .A(\_zyixc_ctx_rdata_29[2][36] ));
Q_ASSIGN U582 ( .B(\mem_a[2][37] ), .A(\_zyixc_ctx_rdata_29[2][37] ));
Q_ASSIGN U583 ( .B(\mem_a[2][38] ), .A(\_zyixc_ctx_rdata_29[2][38] ));
Q_ASSIGN U584 ( .B(\mem_a[2][39] ), .A(\_zyixc_ctx_rdata_29[2][39] ));
Q_ASSIGN U585 ( .B(\mem_a[2][40] ), .A(\_zyixc_ctx_rdata_29[2][40] ));
Q_ASSIGN U586 ( .B(\mem_a[2][41] ), .A(\_zyixc_ctx_rdata_29[2][41] ));
Q_ASSIGN U587 ( .B(\mem_a[2][42] ), .A(\_zyixc_ctx_rdata_29[2][42] ));
Q_ASSIGN U588 ( .B(\mem_a[2][43] ), .A(\_zyixc_ctx_rdata_29[2][43] ));
Q_ASSIGN U589 ( .B(\mem_a[2][44] ), .A(\_zyixc_ctx_rdata_29[2][44] ));
Q_ASSIGN U590 ( .B(\mem_a[2][45] ), .A(\_zyixc_ctx_rdata_29[2][45] ));
Q_ASSIGN U591 ( .B(\mem_a[2][46] ), .A(\_zyixc_ctx_rdata_29[2][46] ));
Q_ASSIGN U592 ( .B(\mem_a[2][47] ), .A(\_zyixc_ctx_rdata_29[2][47] ));
Q_ASSIGN U593 ( .B(\mem_a[2][48] ), .A(\_zyixc_ctx_rdata_29[2][48] ));
Q_ASSIGN U594 ( .B(\mem_a[2][49] ), .A(\_zyixc_ctx_rdata_29[2][49] ));
Q_ASSIGN U595 ( .B(\mem_a[2][50] ), .A(\_zyixc_ctx_rdata_29[2][50] ));
Q_ASSIGN U596 ( .B(\mem_a[2][51] ), .A(\_zyixc_ctx_rdata_29[2][51] ));
Q_ASSIGN U597 ( .B(\mem_a[2][52] ), .A(\_zyixc_ctx_rdata_29[2][52] ));
Q_ASSIGN U598 ( .B(\mem_a[2][53] ), .A(\_zyixc_ctx_rdata_29[2][53] ));
Q_ASSIGN U599 ( .B(\mem_a[2][54] ), .A(\_zyixc_ctx_rdata_29[2][54] ));
Q_ASSIGN U600 ( .B(\mem_a[2][55] ), .A(\_zyixc_ctx_rdata_29[2][55] ));
Q_ASSIGN U601 ( .B(\mem_a[2][56] ), .A(\_zyixc_ctx_rdata_29[2][56] ));
Q_ASSIGN U602 ( .B(\mem_a[2][57] ), .A(\_zyixc_ctx_rdata_29[2][57] ));
Q_ASSIGN U603 ( .B(\mem_a[2][58] ), .A(\_zyixc_ctx_rdata_29[2][58] ));
Q_ASSIGN U604 ( .B(\mem_a[2][59] ), .A(\_zyixc_ctx_rdata_29[2][59] ));
Q_ASSIGN U605 ( .B(\mem_a[2][60] ), .A(\_zyixc_ctx_rdata_29[2][60] ));
Q_ASSIGN U606 ( .B(\mem_a[2][61] ), .A(\_zyixc_ctx_rdata_29[2][61] ));
Q_ASSIGN U607 ( .B(\mem_a[2][62] ), .A(\_zyixc_ctx_rdata_29[2][62] ));
Q_ASSIGN U608 ( .B(\mem_a[2][63] ), .A(\_zyixc_ctx_rdata_29[2][63] ));
Q_ASSIGN U609 ( .B(\mem_a[3][0] ), .A(\_zyixc_ctx_rdata_29[3][0] ));
Q_ASSIGN U610 ( .B(\mem_a[3][1] ), .A(\_zyixc_ctx_rdata_29[3][1] ));
Q_ASSIGN U611 ( .B(\mem_a[3][2] ), .A(\_zyixc_ctx_rdata_29[3][2] ));
Q_ASSIGN U612 ( .B(\mem_a[3][3] ), .A(\_zyixc_ctx_rdata_29[3][3] ));
Q_ASSIGN U613 ( .B(\mem_a[3][4] ), .A(\_zyixc_ctx_rdata_29[3][4] ));
Q_ASSIGN U614 ( .B(\mem_a[3][5] ), .A(\_zyixc_ctx_rdata_29[3][5] ));
Q_ASSIGN U615 ( .B(\mem_a[3][6] ), .A(\_zyixc_ctx_rdata_29[3][6] ));
Q_ASSIGN U616 ( .B(\mem_a[3][7] ), .A(\_zyixc_ctx_rdata_29[3][7] ));
Q_ASSIGN U617 ( .B(\mem_a[3][8] ), .A(\_zyixc_ctx_rdata_29[3][8] ));
Q_ASSIGN U618 ( .B(\mem_a[3][9] ), .A(\_zyixc_ctx_rdata_29[3][9] ));
Q_ASSIGN U619 ( .B(\mem_a[3][10] ), .A(\_zyixc_ctx_rdata_29[3][10] ));
Q_ASSIGN U620 ( .B(\mem_a[3][11] ), .A(\_zyixc_ctx_rdata_29[3][11] ));
Q_ASSIGN U621 ( .B(\mem_a[3][12] ), .A(\_zyixc_ctx_rdata_29[3][12] ));
Q_ASSIGN U622 ( .B(\mem_a[3][13] ), .A(\_zyixc_ctx_rdata_29[3][13] ));
Q_ASSIGN U623 ( .B(\mem_a[3][14] ), .A(\_zyixc_ctx_rdata_29[3][14] ));
Q_ASSIGN U624 ( .B(\mem_a[3][15] ), .A(\_zyixc_ctx_rdata_29[3][15] ));
Q_ASSIGN U625 ( .B(\mem_a[3][16] ), .A(\_zyixc_ctx_rdata_29[3][16] ));
Q_ASSIGN U626 ( .B(\mem_a[3][17] ), .A(\_zyixc_ctx_rdata_29[3][17] ));
Q_ASSIGN U627 ( .B(\mem_a[3][18] ), .A(\_zyixc_ctx_rdata_29[3][18] ));
Q_ASSIGN U628 ( .B(\mem_a[3][19] ), .A(\_zyixc_ctx_rdata_29[3][19] ));
Q_ASSIGN U629 ( .B(\mem_a[3][20] ), .A(\_zyixc_ctx_rdata_29[3][20] ));
Q_ASSIGN U630 ( .B(\mem_a[3][21] ), .A(\_zyixc_ctx_rdata_29[3][21] ));
Q_ASSIGN U631 ( .B(\mem_a[3][22] ), .A(\_zyixc_ctx_rdata_29[3][22] ));
Q_ASSIGN U632 ( .B(\mem_a[3][23] ), .A(\_zyixc_ctx_rdata_29[3][23] ));
Q_ASSIGN U633 ( .B(\mem_a[3][24] ), .A(\_zyixc_ctx_rdata_29[3][24] ));
Q_ASSIGN U634 ( .B(\mem_a[3][25] ), .A(\_zyixc_ctx_rdata_29[3][25] ));
Q_ASSIGN U635 ( .B(\mem_a[3][26] ), .A(\_zyixc_ctx_rdata_29[3][26] ));
Q_ASSIGN U636 ( .B(\mem_a[3][27] ), .A(\_zyixc_ctx_rdata_29[3][27] ));
Q_ASSIGN U637 ( .B(\mem_a[3][28] ), .A(\_zyixc_ctx_rdata_29[3][28] ));
Q_ASSIGN U638 ( .B(\mem_a[3][29] ), .A(\_zyixc_ctx_rdata_29[3][29] ));
Q_ASSIGN U639 ( .B(\mem_a[3][30] ), .A(\_zyixc_ctx_rdata_29[3][30] ));
Q_ASSIGN U640 ( .B(\mem_a[3][31] ), .A(\_zyixc_ctx_rdata_29[3][31] ));
Q_ASSIGN U641 ( .B(\mem_a[3][32] ), .A(\_zyixc_ctx_rdata_29[3][32] ));
Q_ASSIGN U642 ( .B(\mem_a[3][33] ), .A(\_zyixc_ctx_rdata_29[3][33] ));
Q_ASSIGN U643 ( .B(\mem_a[3][34] ), .A(\_zyixc_ctx_rdata_29[3][34] ));
Q_ASSIGN U644 ( .B(\mem_a[3][35] ), .A(\_zyixc_ctx_rdata_29[3][35] ));
Q_ASSIGN U645 ( .B(\mem_a[3][36] ), .A(\_zyixc_ctx_rdata_29[3][36] ));
Q_ASSIGN U646 ( .B(\mem_a[3][37] ), .A(\_zyixc_ctx_rdata_29[3][37] ));
Q_ASSIGN U647 ( .B(\mem_a[3][38] ), .A(\_zyixc_ctx_rdata_29[3][38] ));
Q_ASSIGN U648 ( .B(\mem_a[3][39] ), .A(\_zyixc_ctx_rdata_29[3][39] ));
Q_ASSIGN U649 ( .B(\mem_a[3][40] ), .A(\_zyixc_ctx_rdata_29[3][40] ));
Q_ASSIGN U650 ( .B(\mem_a[3][41] ), .A(\_zyixc_ctx_rdata_29[3][41] ));
Q_ASSIGN U651 ( .B(\mem_a[3][42] ), .A(\_zyixc_ctx_rdata_29[3][42] ));
Q_ASSIGN U652 ( .B(\mem_a[3][43] ), .A(\_zyixc_ctx_rdata_29[3][43] ));
Q_ASSIGN U653 ( .B(\mem_a[3][44] ), .A(\_zyixc_ctx_rdata_29[3][44] ));
Q_ASSIGN U654 ( .B(\mem_a[3][45] ), .A(\_zyixc_ctx_rdata_29[3][45] ));
Q_ASSIGN U655 ( .B(\mem_a[3][46] ), .A(\_zyixc_ctx_rdata_29[3][46] ));
Q_ASSIGN U656 ( .B(\mem_a[3][47] ), .A(\_zyixc_ctx_rdata_29[3][47] ));
Q_ASSIGN U657 ( .B(\mem_a[3][48] ), .A(\_zyixc_ctx_rdata_29[3][48] ));
Q_ASSIGN U658 ( .B(\mem_a[3][49] ), .A(\_zyixc_ctx_rdata_29[3][49] ));
Q_ASSIGN U659 ( .B(\mem_a[3][50] ), .A(\_zyixc_ctx_rdata_29[3][50] ));
Q_ASSIGN U660 ( .B(\mem_a[3][51] ), .A(\_zyixc_ctx_rdata_29[3][51] ));
Q_ASSIGN U661 ( .B(\mem_a[3][52] ), .A(\_zyixc_ctx_rdata_29[3][52] ));
Q_ASSIGN U662 ( .B(\mem_a[3][53] ), .A(\_zyixc_ctx_rdata_29[3][53] ));
Q_ASSIGN U663 ( .B(\mem_a[3][54] ), .A(\_zyixc_ctx_rdata_29[3][54] ));
Q_ASSIGN U664 ( .B(\mem_a[3][55] ), .A(\_zyixc_ctx_rdata_29[3][55] ));
Q_ASSIGN U665 ( .B(\mem_a[3][56] ), .A(\_zyixc_ctx_rdata_29[3][56] ));
Q_ASSIGN U666 ( .B(\mem_a[3][57] ), .A(\_zyixc_ctx_rdata_29[3][57] ));
Q_ASSIGN U667 ( .B(\mem_a[3][58] ), .A(\_zyixc_ctx_rdata_29[3][58] ));
Q_ASSIGN U668 ( .B(\mem_a[3][59] ), .A(\_zyixc_ctx_rdata_29[3][59] ));
Q_ASSIGN U669 ( .B(\mem_a[3][60] ), .A(\_zyixc_ctx_rdata_29[3][60] ));
Q_ASSIGN U670 ( .B(\mem_a[3][61] ), .A(\_zyixc_ctx_rdata_29[3][61] ));
Q_ASSIGN U671 ( .B(\mem_a[3][62] ), .A(\_zyixc_ctx_rdata_29[3][62] ));
Q_ASSIGN U672 ( .B(\mem_a[3][63] ), .A(\_zyixc_ctx_rdata_29[3][63] ));
Q_ASSIGN U673 ( .B(\mem_a[4][0] ), .A(\_zyixc_ctx_rdata_29[4][0] ));
Q_ASSIGN U674 ( .B(\mem_a[4][1] ), .A(\_zyixc_ctx_rdata_29[4][1] ));
Q_ASSIGN U675 ( .B(\mem_a[4][2] ), .A(\_zyixc_ctx_rdata_29[4][2] ));
Q_ASSIGN U676 ( .B(\mem_a[4][3] ), .A(\_zyixc_ctx_rdata_29[4][3] ));
Q_ASSIGN U677 ( .B(\mem_a[4][4] ), .A(\_zyixc_ctx_rdata_29[4][4] ));
Q_ASSIGN U678 ( .B(\mem_a[4][5] ), .A(\_zyixc_ctx_rdata_29[4][5] ));
Q_ASSIGN U679 ( .B(\mem_a[4][6] ), .A(\_zyixc_ctx_rdata_29[4][6] ));
Q_ASSIGN U680 ( .B(\mem_a[4][7] ), .A(\_zyixc_ctx_rdata_29[4][7] ));
Q_ASSIGN U681 ( .B(\mem_a[4][8] ), .A(\_zyixc_ctx_rdata_29[4][8] ));
Q_ASSIGN U682 ( .B(\mem_a[4][9] ), .A(\_zyixc_ctx_rdata_29[4][9] ));
Q_ASSIGN U683 ( .B(\mem_a[4][10] ), .A(\_zyixc_ctx_rdata_29[4][10] ));
Q_ASSIGN U684 ( .B(\mem_a[4][11] ), .A(\_zyixc_ctx_rdata_29[4][11] ));
Q_ASSIGN U685 ( .B(\mem_a[4][12] ), .A(\_zyixc_ctx_rdata_29[4][12] ));
Q_ASSIGN U686 ( .B(\mem_a[4][13] ), .A(\_zyixc_ctx_rdata_29[4][13] ));
Q_ASSIGN U687 ( .B(\mem_a[4][14] ), .A(\_zyixc_ctx_rdata_29[4][14] ));
Q_ASSIGN U688 ( .B(\mem_a[4][15] ), .A(\_zyixc_ctx_rdata_29[4][15] ));
Q_ASSIGN U689 ( .B(\mem_a[4][16] ), .A(\_zyixc_ctx_rdata_29[4][16] ));
Q_ASSIGN U690 ( .B(\mem_a[4][17] ), .A(\_zyixc_ctx_rdata_29[4][17] ));
Q_ASSIGN U691 ( .B(\mem_a[4][18] ), .A(\_zyixc_ctx_rdata_29[4][18] ));
Q_ASSIGN U692 ( .B(\mem_a[4][19] ), .A(\_zyixc_ctx_rdata_29[4][19] ));
Q_ASSIGN U693 ( .B(\mem_a[4][20] ), .A(\_zyixc_ctx_rdata_29[4][20] ));
Q_ASSIGN U694 ( .B(\mem_a[4][21] ), .A(\_zyixc_ctx_rdata_29[4][21] ));
Q_ASSIGN U695 ( .B(\mem_a[4][22] ), .A(\_zyixc_ctx_rdata_29[4][22] ));
Q_ASSIGN U696 ( .B(\mem_a[4][23] ), .A(\_zyixc_ctx_rdata_29[4][23] ));
Q_ASSIGN U697 ( .B(\mem_a[4][24] ), .A(\_zyixc_ctx_rdata_29[4][24] ));
Q_ASSIGN U698 ( .B(\mem_a[4][25] ), .A(\_zyixc_ctx_rdata_29[4][25] ));
Q_ASSIGN U699 ( .B(\mem_a[4][26] ), .A(\_zyixc_ctx_rdata_29[4][26] ));
Q_ASSIGN U700 ( .B(\mem_a[4][27] ), .A(\_zyixc_ctx_rdata_29[4][27] ));
Q_ASSIGN U701 ( .B(\mem_a[4][28] ), .A(\_zyixc_ctx_rdata_29[4][28] ));
Q_ASSIGN U702 ( .B(\mem_a[4][29] ), .A(\_zyixc_ctx_rdata_29[4][29] ));
Q_ASSIGN U703 ( .B(\mem_a[4][30] ), .A(\_zyixc_ctx_rdata_29[4][30] ));
Q_ASSIGN U704 ( .B(\mem_a[4][31] ), .A(\_zyixc_ctx_rdata_29[4][31] ));
Q_ASSIGN U705 ( .B(\mem_a[4][32] ), .A(\_zyixc_ctx_rdata_29[4][32] ));
Q_ASSIGN U706 ( .B(\mem_a[4][33] ), .A(\_zyixc_ctx_rdata_29[4][33] ));
Q_ASSIGN U707 ( .B(\mem_a[4][34] ), .A(\_zyixc_ctx_rdata_29[4][34] ));
Q_ASSIGN U708 ( .B(\mem_a[4][35] ), .A(\_zyixc_ctx_rdata_29[4][35] ));
Q_ASSIGN U709 ( .B(\mem_a[4][36] ), .A(\_zyixc_ctx_rdata_29[4][36] ));
Q_ASSIGN U710 ( .B(\mem_a[4][37] ), .A(\_zyixc_ctx_rdata_29[4][37] ));
Q_ASSIGN U711 ( .B(\mem_a[4][38] ), .A(\_zyixc_ctx_rdata_29[4][38] ));
Q_ASSIGN U712 ( .B(\mem_a[4][39] ), .A(\_zyixc_ctx_rdata_29[4][39] ));
Q_ASSIGN U713 ( .B(\mem_a[4][40] ), .A(\_zyixc_ctx_rdata_29[4][40] ));
Q_ASSIGN U714 ( .B(\mem_a[4][41] ), .A(\_zyixc_ctx_rdata_29[4][41] ));
Q_ASSIGN U715 ( .B(\mem_a[4][42] ), .A(\_zyixc_ctx_rdata_29[4][42] ));
Q_ASSIGN U716 ( .B(\mem_a[4][43] ), .A(\_zyixc_ctx_rdata_29[4][43] ));
Q_ASSIGN U717 ( .B(\mem_a[4][44] ), .A(\_zyixc_ctx_rdata_29[4][44] ));
Q_ASSIGN U718 ( .B(\mem_a[4][45] ), .A(\_zyixc_ctx_rdata_29[4][45] ));
Q_ASSIGN U719 ( .B(\mem_a[4][46] ), .A(\_zyixc_ctx_rdata_29[4][46] ));
Q_ASSIGN U720 ( .B(\mem_a[4][47] ), .A(\_zyixc_ctx_rdata_29[4][47] ));
Q_ASSIGN U721 ( .B(\mem_a[4][48] ), .A(\_zyixc_ctx_rdata_29[4][48] ));
Q_ASSIGN U722 ( .B(\mem_a[4][49] ), .A(\_zyixc_ctx_rdata_29[4][49] ));
Q_ASSIGN U723 ( .B(\mem_a[4][50] ), .A(\_zyixc_ctx_rdata_29[4][50] ));
Q_ASSIGN U724 ( .B(\mem_a[4][51] ), .A(\_zyixc_ctx_rdata_29[4][51] ));
Q_ASSIGN U725 ( .B(\mem_a[4][52] ), .A(\_zyixc_ctx_rdata_29[4][52] ));
Q_ASSIGN U726 ( .B(\mem_a[4][53] ), .A(\_zyixc_ctx_rdata_29[4][53] ));
Q_ASSIGN U727 ( .B(\mem_a[4][54] ), .A(\_zyixc_ctx_rdata_29[4][54] ));
Q_ASSIGN U728 ( .B(\mem_a[4][55] ), .A(\_zyixc_ctx_rdata_29[4][55] ));
Q_ASSIGN U729 ( .B(\mem_a[4][56] ), .A(\_zyixc_ctx_rdata_29[4][56] ));
Q_ASSIGN U730 ( .B(\mem_a[4][57] ), .A(\_zyixc_ctx_rdata_29[4][57] ));
Q_ASSIGN U731 ( .B(\mem_a[4][58] ), .A(\_zyixc_ctx_rdata_29[4][58] ));
Q_ASSIGN U732 ( .B(\mem_a[4][59] ), .A(\_zyixc_ctx_rdata_29[4][59] ));
Q_ASSIGN U733 ( .B(\mem_a[4][60] ), .A(\_zyixc_ctx_rdata_29[4][60] ));
Q_ASSIGN U734 ( .B(\mem_a[4][61] ), .A(\_zyixc_ctx_rdata_29[4][61] ));
Q_ASSIGN U735 ( .B(\mem_a[4][62] ), .A(\_zyixc_ctx_rdata_29[4][62] ));
Q_ASSIGN U736 ( .B(\mem_a[4][63] ), .A(\_zyixc_ctx_rdata_29[4][63] ));
Q_ASSIGN U737 ( .B(\mem_a[5][0] ), .A(\_zyixc_ctx_rdata_29[5][0] ));
Q_ASSIGN U738 ( .B(\mem_a[5][1] ), .A(\_zyixc_ctx_rdata_29[5][1] ));
Q_ASSIGN U739 ( .B(\mem_a[5][2] ), .A(\_zyixc_ctx_rdata_29[5][2] ));
Q_ASSIGN U740 ( .B(\mem_a[5][3] ), .A(\_zyixc_ctx_rdata_29[5][3] ));
Q_ASSIGN U741 ( .B(\mem_a[5][4] ), .A(\_zyixc_ctx_rdata_29[5][4] ));
Q_ASSIGN U742 ( .B(\mem_a[5][5] ), .A(\_zyixc_ctx_rdata_29[5][5] ));
Q_ASSIGN U743 ( .B(\mem_a[5][6] ), .A(\_zyixc_ctx_rdata_29[5][6] ));
Q_ASSIGN U744 ( .B(\mem_a[5][7] ), .A(\_zyixc_ctx_rdata_29[5][7] ));
Q_ASSIGN U745 ( .B(\mem_a[5][8] ), .A(\_zyixc_ctx_rdata_29[5][8] ));
Q_ASSIGN U746 ( .B(\mem_a[5][9] ), .A(\_zyixc_ctx_rdata_29[5][9] ));
Q_ASSIGN U747 ( .B(\mem_a[5][10] ), .A(\_zyixc_ctx_rdata_29[5][10] ));
Q_ASSIGN U748 ( .B(\mem_a[5][11] ), .A(\_zyixc_ctx_rdata_29[5][11] ));
Q_ASSIGN U749 ( .B(\mem_a[5][12] ), .A(\_zyixc_ctx_rdata_29[5][12] ));
Q_ASSIGN U750 ( .B(\mem_a[5][13] ), .A(\_zyixc_ctx_rdata_29[5][13] ));
Q_ASSIGN U751 ( .B(\mem_a[5][14] ), .A(\_zyixc_ctx_rdata_29[5][14] ));
Q_ASSIGN U752 ( .B(\mem_a[5][15] ), .A(\_zyixc_ctx_rdata_29[5][15] ));
Q_ASSIGN U753 ( .B(\mem_a[5][16] ), .A(\_zyixc_ctx_rdata_29[5][16] ));
Q_ASSIGN U754 ( .B(\mem_a[5][17] ), .A(\_zyixc_ctx_rdata_29[5][17] ));
Q_ASSIGN U755 ( .B(\mem_a[5][18] ), .A(\_zyixc_ctx_rdata_29[5][18] ));
Q_ASSIGN U756 ( .B(\mem_a[5][19] ), .A(\_zyixc_ctx_rdata_29[5][19] ));
Q_ASSIGN U757 ( .B(\mem_a[5][20] ), .A(\_zyixc_ctx_rdata_29[5][20] ));
Q_ASSIGN U758 ( .B(\mem_a[5][21] ), .A(\_zyixc_ctx_rdata_29[5][21] ));
Q_ASSIGN U759 ( .B(\mem_a[5][22] ), .A(\_zyixc_ctx_rdata_29[5][22] ));
Q_ASSIGN U760 ( .B(\mem_a[5][23] ), .A(\_zyixc_ctx_rdata_29[5][23] ));
Q_ASSIGN U761 ( .B(\mem_a[5][24] ), .A(\_zyixc_ctx_rdata_29[5][24] ));
Q_ASSIGN U762 ( .B(\mem_a[5][25] ), .A(\_zyixc_ctx_rdata_29[5][25] ));
Q_ASSIGN U763 ( .B(\mem_a[5][26] ), .A(\_zyixc_ctx_rdata_29[5][26] ));
Q_ASSIGN U764 ( .B(\mem_a[5][27] ), .A(\_zyixc_ctx_rdata_29[5][27] ));
Q_ASSIGN U765 ( .B(\mem_a[5][28] ), .A(\_zyixc_ctx_rdata_29[5][28] ));
Q_ASSIGN U766 ( .B(\mem_a[5][29] ), .A(\_zyixc_ctx_rdata_29[5][29] ));
Q_ASSIGN U767 ( .B(\mem_a[5][30] ), .A(\_zyixc_ctx_rdata_29[5][30] ));
Q_ASSIGN U768 ( .B(\mem_a[5][31] ), .A(\_zyixc_ctx_rdata_29[5][31] ));
Q_ASSIGN U769 ( .B(\mem_a[5][32] ), .A(\_zyixc_ctx_rdata_29[5][32] ));
Q_ASSIGN U770 ( .B(\mem_a[5][33] ), .A(\_zyixc_ctx_rdata_29[5][33] ));
Q_ASSIGN U771 ( .B(\mem_a[5][34] ), .A(\_zyixc_ctx_rdata_29[5][34] ));
Q_ASSIGN U772 ( .B(\mem_a[5][35] ), .A(\_zyixc_ctx_rdata_29[5][35] ));
Q_ASSIGN U773 ( .B(\mem_a[5][36] ), .A(\_zyixc_ctx_rdata_29[5][36] ));
Q_ASSIGN U774 ( .B(\mem_a[5][37] ), .A(\_zyixc_ctx_rdata_29[5][37] ));
Q_ASSIGN U775 ( .B(\mem_a[5][38] ), .A(\_zyixc_ctx_rdata_29[5][38] ));
Q_ASSIGN U776 ( .B(\mem_a[5][39] ), .A(\_zyixc_ctx_rdata_29[5][39] ));
Q_ASSIGN U777 ( .B(\mem_a[5][40] ), .A(\_zyixc_ctx_rdata_29[5][40] ));
Q_ASSIGN U778 ( .B(\mem_a[5][41] ), .A(\_zyixc_ctx_rdata_29[5][41] ));
Q_ASSIGN U779 ( .B(\mem_a[5][42] ), .A(\_zyixc_ctx_rdata_29[5][42] ));
Q_ASSIGN U780 ( .B(\mem_a[5][43] ), .A(\_zyixc_ctx_rdata_29[5][43] ));
Q_ASSIGN U781 ( .B(\mem_a[5][44] ), .A(\_zyixc_ctx_rdata_29[5][44] ));
Q_ASSIGN U782 ( .B(\mem_a[5][45] ), .A(\_zyixc_ctx_rdata_29[5][45] ));
Q_ASSIGN U783 ( .B(\mem_a[5][46] ), .A(\_zyixc_ctx_rdata_29[5][46] ));
Q_ASSIGN U784 ( .B(\mem_a[5][47] ), .A(\_zyixc_ctx_rdata_29[5][47] ));
Q_ASSIGN U785 ( .B(\mem_a[5][48] ), .A(\_zyixc_ctx_rdata_29[5][48] ));
Q_ASSIGN U786 ( .B(\mem_a[5][49] ), .A(\_zyixc_ctx_rdata_29[5][49] ));
Q_ASSIGN U787 ( .B(\mem_a[5][50] ), .A(\_zyixc_ctx_rdata_29[5][50] ));
Q_ASSIGN U788 ( .B(\mem_a[5][51] ), .A(\_zyixc_ctx_rdata_29[5][51] ));
Q_ASSIGN U789 ( .B(\mem_a[5][52] ), .A(\_zyixc_ctx_rdata_29[5][52] ));
Q_ASSIGN U790 ( .B(\mem_a[5][53] ), .A(\_zyixc_ctx_rdata_29[5][53] ));
Q_ASSIGN U791 ( .B(\mem_a[5][54] ), .A(\_zyixc_ctx_rdata_29[5][54] ));
Q_ASSIGN U792 ( .B(\mem_a[5][55] ), .A(\_zyixc_ctx_rdata_29[5][55] ));
Q_ASSIGN U793 ( .B(\mem_a[5][56] ), .A(\_zyixc_ctx_rdata_29[5][56] ));
Q_ASSIGN U794 ( .B(\mem_a[5][57] ), .A(\_zyixc_ctx_rdata_29[5][57] ));
Q_ASSIGN U795 ( .B(\mem_a[5][58] ), .A(\_zyixc_ctx_rdata_29[5][58] ));
Q_ASSIGN U796 ( .B(\mem_a[5][59] ), .A(\_zyixc_ctx_rdata_29[5][59] ));
Q_ASSIGN U797 ( .B(\mem_a[5][60] ), .A(\_zyixc_ctx_rdata_29[5][60] ));
Q_ASSIGN U798 ( .B(\mem_a[5][61] ), .A(\_zyixc_ctx_rdata_29[5][61] ));
Q_ASSIGN U799 ( .B(\mem_a[5][62] ), .A(\_zyixc_ctx_rdata_29[5][62] ));
Q_ASSIGN U800 ( .B(\mem_a[5][63] ), .A(\_zyixc_ctx_rdata_29[5][63] ));
Q_ASSIGN U801 ( .B(\mem_a[6][0] ), .A(\_zyixc_ctx_rdata_29[6][0] ));
Q_ASSIGN U802 ( .B(\mem_a[6][1] ), .A(\_zyixc_ctx_rdata_29[6][1] ));
Q_ASSIGN U803 ( .B(\mem_a[6][2] ), .A(\_zyixc_ctx_rdata_29[6][2] ));
Q_ASSIGN U804 ( .B(\mem_a[6][3] ), .A(\_zyixc_ctx_rdata_29[6][3] ));
Q_ASSIGN U805 ( .B(\mem_a[6][4] ), .A(\_zyixc_ctx_rdata_29[6][4] ));
Q_ASSIGN U806 ( .B(\mem_a[6][5] ), .A(\_zyixc_ctx_rdata_29[6][5] ));
Q_ASSIGN U807 ( .B(\mem_a[6][6] ), .A(\_zyixc_ctx_rdata_29[6][6] ));
Q_ASSIGN U808 ( .B(\mem_a[6][7] ), .A(\_zyixc_ctx_rdata_29[6][7] ));
Q_ASSIGN U809 ( .B(\mem_a[6][8] ), .A(\_zyixc_ctx_rdata_29[6][8] ));
Q_ASSIGN U810 ( .B(\mem_a[6][9] ), .A(\_zyixc_ctx_rdata_29[6][9] ));
Q_ASSIGN U811 ( .B(\mem_a[6][10] ), .A(\_zyixc_ctx_rdata_29[6][10] ));
Q_ASSIGN U812 ( .B(\mem_a[6][11] ), .A(\_zyixc_ctx_rdata_29[6][11] ));
Q_ASSIGN U813 ( .B(\mem_a[6][12] ), .A(\_zyixc_ctx_rdata_29[6][12] ));
Q_ASSIGN U814 ( .B(\mem_a[6][13] ), .A(\_zyixc_ctx_rdata_29[6][13] ));
Q_ASSIGN U815 ( .B(\mem_a[6][14] ), .A(\_zyixc_ctx_rdata_29[6][14] ));
Q_ASSIGN U816 ( .B(\mem_a[6][15] ), .A(\_zyixc_ctx_rdata_29[6][15] ));
Q_ASSIGN U817 ( .B(\mem_a[6][16] ), .A(\_zyixc_ctx_rdata_29[6][16] ));
Q_ASSIGN U818 ( .B(\mem_a[6][17] ), .A(\_zyixc_ctx_rdata_29[6][17] ));
Q_ASSIGN U819 ( .B(\mem_a[6][18] ), .A(\_zyixc_ctx_rdata_29[6][18] ));
Q_ASSIGN U820 ( .B(\mem_a[6][19] ), .A(\_zyixc_ctx_rdata_29[6][19] ));
Q_ASSIGN U821 ( .B(\mem_a[6][20] ), .A(\_zyixc_ctx_rdata_29[6][20] ));
Q_ASSIGN U822 ( .B(\mem_a[6][21] ), .A(\_zyixc_ctx_rdata_29[6][21] ));
Q_ASSIGN U823 ( .B(\mem_a[6][22] ), .A(\_zyixc_ctx_rdata_29[6][22] ));
Q_ASSIGN U824 ( .B(\mem_a[6][23] ), .A(\_zyixc_ctx_rdata_29[6][23] ));
Q_ASSIGN U825 ( .B(\mem_a[6][24] ), .A(\_zyixc_ctx_rdata_29[6][24] ));
Q_ASSIGN U826 ( .B(\mem_a[6][25] ), .A(\_zyixc_ctx_rdata_29[6][25] ));
Q_ASSIGN U827 ( .B(\mem_a[6][26] ), .A(\_zyixc_ctx_rdata_29[6][26] ));
Q_ASSIGN U828 ( .B(\mem_a[6][27] ), .A(\_zyixc_ctx_rdata_29[6][27] ));
Q_ASSIGN U829 ( .B(\mem_a[6][28] ), .A(\_zyixc_ctx_rdata_29[6][28] ));
Q_ASSIGN U830 ( .B(\mem_a[6][29] ), .A(\_zyixc_ctx_rdata_29[6][29] ));
Q_ASSIGN U831 ( .B(\mem_a[6][30] ), .A(\_zyixc_ctx_rdata_29[6][30] ));
Q_ASSIGN U832 ( .B(\mem_a[6][31] ), .A(\_zyixc_ctx_rdata_29[6][31] ));
Q_ASSIGN U833 ( .B(\mem_a[6][32] ), .A(\_zyixc_ctx_rdata_29[6][32] ));
Q_ASSIGN U834 ( .B(\mem_a[6][33] ), .A(\_zyixc_ctx_rdata_29[6][33] ));
Q_ASSIGN U835 ( .B(\mem_a[6][34] ), .A(\_zyixc_ctx_rdata_29[6][34] ));
Q_ASSIGN U836 ( .B(\mem_a[6][35] ), .A(\_zyixc_ctx_rdata_29[6][35] ));
Q_ASSIGN U837 ( .B(\mem_a[6][36] ), .A(\_zyixc_ctx_rdata_29[6][36] ));
Q_ASSIGN U838 ( .B(\mem_a[6][37] ), .A(\_zyixc_ctx_rdata_29[6][37] ));
Q_ASSIGN U839 ( .B(\mem_a[6][38] ), .A(\_zyixc_ctx_rdata_29[6][38] ));
Q_ASSIGN U840 ( .B(\mem_a[6][39] ), .A(\_zyixc_ctx_rdata_29[6][39] ));
Q_ASSIGN U841 ( .B(\mem_a[6][40] ), .A(\_zyixc_ctx_rdata_29[6][40] ));
Q_ASSIGN U842 ( .B(\mem_a[6][41] ), .A(\_zyixc_ctx_rdata_29[6][41] ));
Q_ASSIGN U843 ( .B(\mem_a[6][42] ), .A(\_zyixc_ctx_rdata_29[6][42] ));
Q_ASSIGN U844 ( .B(\mem_a[6][43] ), .A(\_zyixc_ctx_rdata_29[6][43] ));
Q_ASSIGN U845 ( .B(\mem_a[6][44] ), .A(\_zyixc_ctx_rdata_29[6][44] ));
Q_ASSIGN U846 ( .B(\mem_a[6][45] ), .A(\_zyixc_ctx_rdata_29[6][45] ));
Q_ASSIGN U847 ( .B(\mem_a[6][46] ), .A(\_zyixc_ctx_rdata_29[6][46] ));
Q_ASSIGN U848 ( .B(\mem_a[6][47] ), .A(\_zyixc_ctx_rdata_29[6][47] ));
Q_ASSIGN U849 ( .B(\mem_a[6][48] ), .A(\_zyixc_ctx_rdata_29[6][48] ));
Q_ASSIGN U850 ( .B(\mem_a[6][49] ), .A(\_zyixc_ctx_rdata_29[6][49] ));
Q_ASSIGN U851 ( .B(\mem_a[6][50] ), .A(\_zyixc_ctx_rdata_29[6][50] ));
Q_ASSIGN U852 ( .B(\mem_a[6][51] ), .A(\_zyixc_ctx_rdata_29[6][51] ));
Q_ASSIGN U853 ( .B(\mem_a[6][52] ), .A(\_zyixc_ctx_rdata_29[6][52] ));
Q_ASSIGN U854 ( .B(\mem_a[6][53] ), .A(\_zyixc_ctx_rdata_29[6][53] ));
Q_ASSIGN U855 ( .B(\mem_a[6][54] ), .A(\_zyixc_ctx_rdata_29[6][54] ));
Q_ASSIGN U856 ( .B(\mem_a[6][55] ), .A(\_zyixc_ctx_rdata_29[6][55] ));
Q_ASSIGN U857 ( .B(\mem_a[6][56] ), .A(\_zyixc_ctx_rdata_29[6][56] ));
Q_ASSIGN U858 ( .B(\mem_a[6][57] ), .A(\_zyixc_ctx_rdata_29[6][57] ));
Q_ASSIGN U859 ( .B(\mem_a[6][58] ), .A(\_zyixc_ctx_rdata_29[6][58] ));
Q_ASSIGN U860 ( .B(\mem_a[6][59] ), .A(\_zyixc_ctx_rdata_29[6][59] ));
Q_ASSIGN U861 ( .B(\mem_a[6][60] ), .A(\_zyixc_ctx_rdata_29[6][60] ));
Q_ASSIGN U862 ( .B(\mem_a[6][61] ), .A(\_zyixc_ctx_rdata_29[6][61] ));
Q_ASSIGN U863 ( .B(\mem_a[6][62] ), .A(\_zyixc_ctx_rdata_29[6][62] ));
Q_ASSIGN U864 ( .B(\mem_a[6][63] ), .A(\_zyixc_ctx_rdata_29[6][63] ));
Q_ASSIGN U865 ( .B(\mem_a[7][0] ), .A(\_zyixc_ctx_rdata_29[7][0] ));
Q_ASSIGN U866 ( .B(\mem_a[7][1] ), .A(\_zyixc_ctx_rdata_29[7][1] ));
Q_ASSIGN U867 ( .B(\mem_a[7][2] ), .A(\_zyixc_ctx_rdata_29[7][2] ));
Q_ASSIGN U868 ( .B(\mem_a[7][3] ), .A(\_zyixc_ctx_rdata_29[7][3] ));
Q_ASSIGN U869 ( .B(\mem_a[7][4] ), .A(\_zyixc_ctx_rdata_29[7][4] ));
Q_ASSIGN U870 ( .B(\mem_a[7][5] ), .A(\_zyixc_ctx_rdata_29[7][5] ));
Q_ASSIGN U871 ( .B(\mem_a[7][6] ), .A(\_zyixc_ctx_rdata_29[7][6] ));
Q_ASSIGN U872 ( .B(\mem_a[7][7] ), .A(\_zyixc_ctx_rdata_29[7][7] ));
Q_ASSIGN U873 ( .B(\mem_a[7][8] ), .A(\_zyixc_ctx_rdata_29[7][8] ));
Q_ASSIGN U874 ( .B(\mem_a[7][9] ), .A(\_zyixc_ctx_rdata_29[7][9] ));
Q_ASSIGN U875 ( .B(\mem_a[7][10] ), .A(\_zyixc_ctx_rdata_29[7][10] ));
Q_ASSIGN U876 ( .B(\mem_a[7][11] ), .A(\_zyixc_ctx_rdata_29[7][11] ));
Q_ASSIGN U877 ( .B(\mem_a[7][12] ), .A(\_zyixc_ctx_rdata_29[7][12] ));
Q_ASSIGN U878 ( .B(\mem_a[7][13] ), .A(\_zyixc_ctx_rdata_29[7][13] ));
Q_ASSIGN U879 ( .B(\mem_a[7][14] ), .A(\_zyixc_ctx_rdata_29[7][14] ));
Q_ASSIGN U880 ( .B(\mem_a[7][15] ), .A(\_zyixc_ctx_rdata_29[7][15] ));
Q_ASSIGN U881 ( .B(\mem_a[7][16] ), .A(\_zyixc_ctx_rdata_29[7][16] ));
Q_ASSIGN U882 ( .B(\mem_a[7][17] ), .A(\_zyixc_ctx_rdata_29[7][17] ));
Q_ASSIGN U883 ( .B(\mem_a[7][18] ), .A(\_zyixc_ctx_rdata_29[7][18] ));
Q_ASSIGN U884 ( .B(\mem_a[7][19] ), .A(\_zyixc_ctx_rdata_29[7][19] ));
Q_ASSIGN U885 ( .B(\mem_a[7][20] ), .A(\_zyixc_ctx_rdata_29[7][20] ));
Q_ASSIGN U886 ( .B(\mem_a[7][21] ), .A(\_zyixc_ctx_rdata_29[7][21] ));
Q_ASSIGN U887 ( .B(\mem_a[7][22] ), .A(\_zyixc_ctx_rdata_29[7][22] ));
Q_ASSIGN U888 ( .B(\mem_a[7][23] ), .A(\_zyixc_ctx_rdata_29[7][23] ));
Q_ASSIGN U889 ( .B(\mem_a[7][24] ), .A(\_zyixc_ctx_rdata_29[7][24] ));
Q_ASSIGN U890 ( .B(\mem_a[7][25] ), .A(\_zyixc_ctx_rdata_29[7][25] ));
Q_ASSIGN U891 ( .B(\mem_a[7][26] ), .A(\_zyixc_ctx_rdata_29[7][26] ));
Q_ASSIGN U892 ( .B(\mem_a[7][27] ), .A(\_zyixc_ctx_rdata_29[7][27] ));
Q_ASSIGN U893 ( .B(\mem_a[7][28] ), .A(\_zyixc_ctx_rdata_29[7][28] ));
Q_ASSIGN U894 ( .B(\mem_a[7][29] ), .A(\_zyixc_ctx_rdata_29[7][29] ));
Q_ASSIGN U895 ( .B(\mem_a[7][30] ), .A(\_zyixc_ctx_rdata_29[7][30] ));
Q_ASSIGN U896 ( .B(\mem_a[7][31] ), .A(\_zyixc_ctx_rdata_29[7][31] ));
Q_ASSIGN U897 ( .B(\mem_a[7][32] ), .A(\_zyixc_ctx_rdata_29[7][32] ));
Q_ASSIGN U898 ( .B(\mem_a[7][33] ), .A(\_zyixc_ctx_rdata_29[7][33] ));
Q_ASSIGN U899 ( .B(\mem_a[7][34] ), .A(\_zyixc_ctx_rdata_29[7][34] ));
Q_ASSIGN U900 ( .B(\mem_a[7][35] ), .A(\_zyixc_ctx_rdata_29[7][35] ));
Q_ASSIGN U901 ( .B(\mem_a[7][36] ), .A(\_zyixc_ctx_rdata_29[7][36] ));
Q_ASSIGN U902 ( .B(\mem_a[7][37] ), .A(\_zyixc_ctx_rdata_29[7][37] ));
Q_ASSIGN U903 ( .B(\mem_a[7][38] ), .A(\_zyixc_ctx_rdata_29[7][38] ));
Q_ASSIGN U904 ( .B(\mem_a[7][39] ), .A(\_zyixc_ctx_rdata_29[7][39] ));
Q_ASSIGN U905 ( .B(\mem_a[7][40] ), .A(\_zyixc_ctx_rdata_29[7][40] ));
Q_ASSIGN U906 ( .B(\mem_a[7][41] ), .A(\_zyixc_ctx_rdata_29[7][41] ));
Q_ASSIGN U907 ( .B(\mem_a[7][42] ), .A(\_zyixc_ctx_rdata_29[7][42] ));
Q_ASSIGN U908 ( .B(\mem_a[7][43] ), .A(\_zyixc_ctx_rdata_29[7][43] ));
Q_ASSIGN U909 ( .B(\mem_a[7][44] ), .A(\_zyixc_ctx_rdata_29[7][44] ));
Q_ASSIGN U910 ( .B(\mem_a[7][45] ), .A(\_zyixc_ctx_rdata_29[7][45] ));
Q_ASSIGN U911 ( .B(\mem_a[7][46] ), .A(\_zyixc_ctx_rdata_29[7][46] ));
Q_ASSIGN U912 ( .B(\mem_a[7][47] ), .A(\_zyixc_ctx_rdata_29[7][47] ));
Q_ASSIGN U913 ( .B(\mem_a[7][48] ), .A(\_zyixc_ctx_rdata_29[7][48] ));
Q_ASSIGN U914 ( .B(\mem_a[7][49] ), .A(\_zyixc_ctx_rdata_29[7][49] ));
Q_ASSIGN U915 ( .B(\mem_a[7][50] ), .A(\_zyixc_ctx_rdata_29[7][50] ));
Q_ASSIGN U916 ( .B(\mem_a[7][51] ), .A(\_zyixc_ctx_rdata_29[7][51] ));
Q_ASSIGN U917 ( .B(\mem_a[7][52] ), .A(\_zyixc_ctx_rdata_29[7][52] ));
Q_ASSIGN U918 ( .B(\mem_a[7][53] ), .A(\_zyixc_ctx_rdata_29[7][53] ));
Q_ASSIGN U919 ( .B(\mem_a[7][54] ), .A(\_zyixc_ctx_rdata_29[7][54] ));
Q_ASSIGN U920 ( .B(\mem_a[7][55] ), .A(\_zyixc_ctx_rdata_29[7][55] ));
Q_ASSIGN U921 ( .B(\mem_a[7][56] ), .A(\_zyixc_ctx_rdata_29[7][56] ));
Q_ASSIGN U922 ( .B(\mem_a[7][57] ), .A(\_zyixc_ctx_rdata_29[7][57] ));
Q_ASSIGN U923 ( .B(\mem_a[7][58] ), .A(\_zyixc_ctx_rdata_29[7][58] ));
Q_ASSIGN U924 ( .B(\mem_a[7][59] ), .A(\_zyixc_ctx_rdata_29[7][59] ));
Q_ASSIGN U925 ( .B(\mem_a[7][60] ), .A(\_zyixc_ctx_rdata_29[7][60] ));
Q_ASSIGN U926 ( .B(\mem_a[7][61] ), .A(\_zyixc_ctx_rdata_29[7][61] ));
Q_ASSIGN U927 ( .B(\mem_a[7][62] ), .A(\_zyixc_ctx_rdata_29[7][62] ));
Q_ASSIGN U928 ( .B(\mem_a[7][63] ), .A(\_zyixc_ctx_rdata_29[7][63] ));
Q_ASSIGN U929 ( .B(\mem_a[8][0] ), .A(\_zyixc_ctx_rdata_29[8][0] ));
Q_ASSIGN U930 ( .B(\mem_a[8][1] ), .A(\_zyixc_ctx_rdata_29[8][1] ));
Q_ASSIGN U931 ( .B(\mem_a[8][2] ), .A(\_zyixc_ctx_rdata_29[8][2] ));
Q_ASSIGN U932 ( .B(\mem_a[8][3] ), .A(\_zyixc_ctx_rdata_29[8][3] ));
Q_ASSIGN U933 ( .B(\mem_a[8][4] ), .A(\_zyixc_ctx_rdata_29[8][4] ));
Q_ASSIGN U934 ( .B(\mem_a[8][5] ), .A(\_zyixc_ctx_rdata_29[8][5] ));
Q_ASSIGN U935 ( .B(\mem_a[8][6] ), .A(\_zyixc_ctx_rdata_29[8][6] ));
Q_ASSIGN U936 ( .B(\mem_a[8][7] ), .A(\_zyixc_ctx_rdata_29[8][7] ));
Q_ASSIGN U937 ( .B(\mem_a[8][8] ), .A(\_zyixc_ctx_rdata_29[8][8] ));
Q_ASSIGN U938 ( .B(\mem_a[8][9] ), .A(\_zyixc_ctx_rdata_29[8][9] ));
Q_ASSIGN U939 ( .B(\mem_a[8][10] ), .A(\_zyixc_ctx_rdata_29[8][10] ));
Q_ASSIGN U940 ( .B(\mem_a[8][11] ), .A(\_zyixc_ctx_rdata_29[8][11] ));
Q_ASSIGN U941 ( .B(\mem_a[8][12] ), .A(\_zyixc_ctx_rdata_29[8][12] ));
Q_ASSIGN U942 ( .B(\mem_a[8][13] ), .A(\_zyixc_ctx_rdata_29[8][13] ));
Q_ASSIGN U943 ( .B(\mem_a[8][14] ), .A(\_zyixc_ctx_rdata_29[8][14] ));
Q_ASSIGN U944 ( .B(\mem_a[8][15] ), .A(\_zyixc_ctx_rdata_29[8][15] ));
Q_ASSIGN U945 ( .B(\mem_a[8][16] ), .A(\_zyixc_ctx_rdata_29[8][16] ));
Q_ASSIGN U946 ( .B(\mem_a[8][17] ), .A(\_zyixc_ctx_rdata_29[8][17] ));
Q_ASSIGN U947 ( .B(\mem_a[8][18] ), .A(\_zyixc_ctx_rdata_29[8][18] ));
Q_ASSIGN U948 ( .B(\mem_a[8][19] ), .A(\_zyixc_ctx_rdata_29[8][19] ));
Q_ASSIGN U949 ( .B(\mem_a[8][20] ), .A(\_zyixc_ctx_rdata_29[8][20] ));
Q_ASSIGN U950 ( .B(\mem_a[8][21] ), .A(\_zyixc_ctx_rdata_29[8][21] ));
Q_ASSIGN U951 ( .B(\mem_a[8][22] ), .A(\_zyixc_ctx_rdata_29[8][22] ));
Q_ASSIGN U952 ( .B(\mem_a[8][23] ), .A(\_zyixc_ctx_rdata_29[8][23] ));
Q_ASSIGN U953 ( .B(\mem_a[8][24] ), .A(\_zyixc_ctx_rdata_29[8][24] ));
Q_ASSIGN U954 ( .B(\mem_a[8][25] ), .A(\_zyixc_ctx_rdata_29[8][25] ));
Q_ASSIGN U955 ( .B(\mem_a[8][26] ), .A(\_zyixc_ctx_rdata_29[8][26] ));
Q_ASSIGN U956 ( .B(\mem_a[8][27] ), .A(\_zyixc_ctx_rdata_29[8][27] ));
Q_ASSIGN U957 ( .B(\mem_a[8][28] ), .A(\_zyixc_ctx_rdata_29[8][28] ));
Q_ASSIGN U958 ( .B(\mem_a[8][29] ), .A(\_zyixc_ctx_rdata_29[8][29] ));
Q_ASSIGN U959 ( .B(\mem_a[8][30] ), .A(\_zyixc_ctx_rdata_29[8][30] ));
Q_ASSIGN U960 ( .B(\mem_a[8][31] ), .A(\_zyixc_ctx_rdata_29[8][31] ));
Q_ASSIGN U961 ( .B(\mem_a[8][32] ), .A(\_zyixc_ctx_rdata_29[8][32] ));
Q_ASSIGN U962 ( .B(\mem_a[8][33] ), .A(\_zyixc_ctx_rdata_29[8][33] ));
Q_ASSIGN U963 ( .B(\mem_a[8][34] ), .A(\_zyixc_ctx_rdata_29[8][34] ));
Q_ASSIGN U964 ( .B(\mem_a[8][35] ), .A(\_zyixc_ctx_rdata_29[8][35] ));
Q_ASSIGN U965 ( .B(\mem_a[8][36] ), .A(\_zyixc_ctx_rdata_29[8][36] ));
Q_ASSIGN U966 ( .B(\mem_a[8][37] ), .A(\_zyixc_ctx_rdata_29[8][37] ));
Q_ASSIGN U967 ( .B(\mem_a[8][38] ), .A(\_zyixc_ctx_rdata_29[8][38] ));
Q_ASSIGN U968 ( .B(\mem_a[8][39] ), .A(\_zyixc_ctx_rdata_29[8][39] ));
Q_ASSIGN U969 ( .B(\mem_a[8][40] ), .A(\_zyixc_ctx_rdata_29[8][40] ));
Q_ASSIGN U970 ( .B(\mem_a[8][41] ), .A(\_zyixc_ctx_rdata_29[8][41] ));
Q_ASSIGN U971 ( .B(\mem_a[8][42] ), .A(\_zyixc_ctx_rdata_29[8][42] ));
Q_ASSIGN U972 ( .B(\mem_a[8][43] ), .A(\_zyixc_ctx_rdata_29[8][43] ));
Q_ASSIGN U973 ( .B(\mem_a[8][44] ), .A(\_zyixc_ctx_rdata_29[8][44] ));
Q_ASSIGN U974 ( .B(\mem_a[8][45] ), .A(\_zyixc_ctx_rdata_29[8][45] ));
Q_ASSIGN U975 ( .B(\mem_a[8][46] ), .A(\_zyixc_ctx_rdata_29[8][46] ));
Q_ASSIGN U976 ( .B(\mem_a[8][47] ), .A(\_zyixc_ctx_rdata_29[8][47] ));
Q_ASSIGN U977 ( .B(\mem_a[8][48] ), .A(\_zyixc_ctx_rdata_29[8][48] ));
Q_ASSIGN U978 ( .B(\mem_a[8][49] ), .A(\_zyixc_ctx_rdata_29[8][49] ));
Q_ASSIGN U979 ( .B(\mem_a[8][50] ), .A(\_zyixc_ctx_rdata_29[8][50] ));
Q_ASSIGN U980 ( .B(\mem_a[8][51] ), .A(\_zyixc_ctx_rdata_29[8][51] ));
Q_ASSIGN U981 ( .B(\mem_a[8][52] ), .A(\_zyixc_ctx_rdata_29[8][52] ));
Q_ASSIGN U982 ( .B(\mem_a[8][53] ), .A(\_zyixc_ctx_rdata_29[8][53] ));
Q_ASSIGN U983 ( .B(\mem_a[8][54] ), .A(\_zyixc_ctx_rdata_29[8][54] ));
Q_ASSIGN U984 ( .B(\mem_a[8][55] ), .A(\_zyixc_ctx_rdata_29[8][55] ));
Q_ASSIGN U985 ( .B(\mem_a[8][56] ), .A(\_zyixc_ctx_rdata_29[8][56] ));
Q_ASSIGN U986 ( .B(\mem_a[8][57] ), .A(\_zyixc_ctx_rdata_29[8][57] ));
Q_ASSIGN U987 ( .B(\mem_a[8][58] ), .A(\_zyixc_ctx_rdata_29[8][58] ));
Q_ASSIGN U988 ( .B(\mem_a[8][59] ), .A(\_zyixc_ctx_rdata_29[8][59] ));
Q_ASSIGN U989 ( .B(\mem_a[8][60] ), .A(\_zyixc_ctx_rdata_29[8][60] ));
Q_ASSIGN U990 ( .B(\mem_a[8][61] ), .A(\_zyixc_ctx_rdata_29[8][61] ));
Q_ASSIGN U991 ( .B(\mem_a[8][62] ), .A(\_zyixc_ctx_rdata_29[8][62] ));
Q_ASSIGN U992 ( .B(\mem_a[8][63] ), .A(\_zyixc_ctx_rdata_29[8][63] ));
Q_ASSIGN U993 ( .B(\mem_a[9][0] ), .A(\_zyixc_ctx_rdata_29[9][0] ));
Q_ASSIGN U994 ( .B(\mem_a[9][1] ), .A(\_zyixc_ctx_rdata_29[9][1] ));
Q_ASSIGN U995 ( .B(\mem_a[9][2] ), .A(\_zyixc_ctx_rdata_29[9][2] ));
Q_ASSIGN U996 ( .B(\mem_a[9][3] ), .A(\_zyixc_ctx_rdata_29[9][3] ));
Q_ASSIGN U997 ( .B(\mem_a[9][4] ), .A(\_zyixc_ctx_rdata_29[9][4] ));
Q_ASSIGN U998 ( .B(\mem_a[9][5] ), .A(\_zyixc_ctx_rdata_29[9][5] ));
Q_ASSIGN U999 ( .B(\mem_a[9][6] ), .A(\_zyixc_ctx_rdata_29[9][6] ));
Q_ASSIGN U1000 ( .B(\mem_a[9][7] ), .A(\_zyixc_ctx_rdata_29[9][7] ));
Q_ASSIGN U1001 ( .B(\mem_a[9][8] ), .A(\_zyixc_ctx_rdata_29[9][8] ));
Q_ASSIGN U1002 ( .B(\mem_a[9][9] ), .A(\_zyixc_ctx_rdata_29[9][9] ));
Q_ASSIGN U1003 ( .B(\mem_a[9][10] ), .A(\_zyixc_ctx_rdata_29[9][10] ));
Q_ASSIGN U1004 ( .B(\mem_a[9][11] ), .A(\_zyixc_ctx_rdata_29[9][11] ));
Q_ASSIGN U1005 ( .B(\mem_a[9][12] ), .A(\_zyixc_ctx_rdata_29[9][12] ));
Q_ASSIGN U1006 ( .B(\mem_a[9][13] ), .A(\_zyixc_ctx_rdata_29[9][13] ));
Q_ASSIGN U1007 ( .B(\mem_a[9][14] ), .A(\_zyixc_ctx_rdata_29[9][14] ));
Q_ASSIGN U1008 ( .B(\mem_a[9][15] ), .A(\_zyixc_ctx_rdata_29[9][15] ));
Q_ASSIGN U1009 ( .B(\mem_a[9][16] ), .A(\_zyixc_ctx_rdata_29[9][16] ));
Q_ASSIGN U1010 ( .B(\mem_a[9][17] ), .A(\_zyixc_ctx_rdata_29[9][17] ));
Q_ASSIGN U1011 ( .B(\mem_a[9][18] ), .A(\_zyixc_ctx_rdata_29[9][18] ));
Q_ASSIGN U1012 ( .B(\mem_a[9][19] ), .A(\_zyixc_ctx_rdata_29[9][19] ));
Q_ASSIGN U1013 ( .B(\mem_a[9][20] ), .A(\_zyixc_ctx_rdata_29[9][20] ));
Q_ASSIGN U1014 ( .B(\mem_a[9][21] ), .A(\_zyixc_ctx_rdata_29[9][21] ));
Q_ASSIGN U1015 ( .B(\mem_a[9][22] ), .A(\_zyixc_ctx_rdata_29[9][22] ));
Q_ASSIGN U1016 ( .B(\mem_a[9][23] ), .A(\_zyixc_ctx_rdata_29[9][23] ));
Q_ASSIGN U1017 ( .B(\mem_a[9][24] ), .A(\_zyixc_ctx_rdata_29[9][24] ));
Q_ASSIGN U1018 ( .B(\mem_a[9][25] ), .A(\_zyixc_ctx_rdata_29[9][25] ));
Q_ASSIGN U1019 ( .B(\mem_a[9][26] ), .A(\_zyixc_ctx_rdata_29[9][26] ));
Q_ASSIGN U1020 ( .B(\mem_a[9][27] ), .A(\_zyixc_ctx_rdata_29[9][27] ));
Q_ASSIGN U1021 ( .B(\mem_a[9][28] ), .A(\_zyixc_ctx_rdata_29[9][28] ));
Q_ASSIGN U1022 ( .B(\mem_a[9][29] ), .A(\_zyixc_ctx_rdata_29[9][29] ));
Q_ASSIGN U1023 ( .B(\mem_a[9][30] ), .A(\_zyixc_ctx_rdata_29[9][30] ));
Q_ASSIGN U1024 ( .B(\mem_a[9][31] ), .A(\_zyixc_ctx_rdata_29[9][31] ));
Q_ASSIGN U1025 ( .B(\mem_a[9][32] ), .A(\_zyixc_ctx_rdata_29[9][32] ));
Q_ASSIGN U1026 ( .B(\mem_a[9][33] ), .A(\_zyixc_ctx_rdata_29[9][33] ));
Q_ASSIGN U1027 ( .B(\mem_a[9][34] ), .A(\_zyixc_ctx_rdata_29[9][34] ));
Q_ASSIGN U1028 ( .B(\mem_a[9][35] ), .A(\_zyixc_ctx_rdata_29[9][35] ));
Q_ASSIGN U1029 ( .B(\mem_a[9][36] ), .A(\_zyixc_ctx_rdata_29[9][36] ));
Q_ASSIGN U1030 ( .B(\mem_a[9][37] ), .A(\_zyixc_ctx_rdata_29[9][37] ));
Q_ASSIGN U1031 ( .B(\mem_a[9][38] ), .A(\_zyixc_ctx_rdata_29[9][38] ));
Q_ASSIGN U1032 ( .B(\mem_a[9][39] ), .A(\_zyixc_ctx_rdata_29[9][39] ));
Q_ASSIGN U1033 ( .B(\mem_a[9][40] ), .A(\_zyixc_ctx_rdata_29[9][40] ));
Q_ASSIGN U1034 ( .B(\mem_a[9][41] ), .A(\_zyixc_ctx_rdata_29[9][41] ));
Q_ASSIGN U1035 ( .B(\mem_a[9][42] ), .A(\_zyixc_ctx_rdata_29[9][42] ));
Q_ASSIGN U1036 ( .B(\mem_a[9][43] ), .A(\_zyixc_ctx_rdata_29[9][43] ));
Q_ASSIGN U1037 ( .B(\mem_a[9][44] ), .A(\_zyixc_ctx_rdata_29[9][44] ));
Q_ASSIGN U1038 ( .B(\mem_a[9][45] ), .A(\_zyixc_ctx_rdata_29[9][45] ));
Q_ASSIGN U1039 ( .B(\mem_a[9][46] ), .A(\_zyixc_ctx_rdata_29[9][46] ));
Q_ASSIGN U1040 ( .B(\mem_a[9][47] ), .A(\_zyixc_ctx_rdata_29[9][47] ));
Q_ASSIGN U1041 ( .B(\mem_a[9][48] ), .A(\_zyixc_ctx_rdata_29[9][48] ));
Q_ASSIGN U1042 ( .B(\mem_a[9][49] ), .A(\_zyixc_ctx_rdata_29[9][49] ));
Q_ASSIGN U1043 ( .B(\mem_a[9][50] ), .A(\_zyixc_ctx_rdata_29[9][50] ));
Q_ASSIGN U1044 ( .B(\mem_a[9][51] ), .A(\_zyixc_ctx_rdata_29[9][51] ));
Q_ASSIGN U1045 ( .B(\mem_a[9][52] ), .A(\_zyixc_ctx_rdata_29[9][52] ));
Q_ASSIGN U1046 ( .B(\mem_a[9][53] ), .A(\_zyixc_ctx_rdata_29[9][53] ));
Q_ASSIGN U1047 ( .B(\mem_a[9][54] ), .A(\_zyixc_ctx_rdata_29[9][54] ));
Q_ASSIGN U1048 ( .B(\mem_a[9][55] ), .A(\_zyixc_ctx_rdata_29[9][55] ));
Q_ASSIGN U1049 ( .B(\mem_a[9][56] ), .A(\_zyixc_ctx_rdata_29[9][56] ));
Q_ASSIGN U1050 ( .B(\mem_a[9][57] ), .A(\_zyixc_ctx_rdata_29[9][57] ));
Q_ASSIGN U1051 ( .B(\mem_a[9][58] ), .A(\_zyixc_ctx_rdata_29[9][58] ));
Q_ASSIGN U1052 ( .B(\mem_a[9][59] ), .A(\_zyixc_ctx_rdata_29[9][59] ));
Q_ASSIGN U1053 ( .B(\mem_a[9][60] ), .A(\_zyixc_ctx_rdata_29[9][60] ));
Q_ASSIGN U1054 ( .B(\mem_a[9][61] ), .A(\_zyixc_ctx_rdata_29[9][61] ));
Q_ASSIGN U1055 ( .B(\mem_a[9][62] ), .A(\_zyixc_ctx_rdata_29[9][62] ));
Q_ASSIGN U1056 ( .B(\mem_a[9][63] ), .A(\_zyixc_ctx_rdata_29[9][63] ));
Q_ASSIGN U1057 ( .B(\mem_a[10][0] ), .A(\_zyixc_ctx_rdata_29[10][0] ));
Q_ASSIGN U1058 ( .B(\mem_a[10][1] ), .A(\_zyixc_ctx_rdata_29[10][1] ));
Q_ASSIGN U1059 ( .B(\mem_a[10][2] ), .A(\_zyixc_ctx_rdata_29[10][2] ));
Q_ASSIGN U1060 ( .B(\mem_a[10][3] ), .A(\_zyixc_ctx_rdata_29[10][3] ));
Q_ASSIGN U1061 ( .B(\mem_a[10][4] ), .A(\_zyixc_ctx_rdata_29[10][4] ));
Q_ASSIGN U1062 ( .B(\mem_a[10][5] ), .A(\_zyixc_ctx_rdata_29[10][5] ));
Q_ASSIGN U1063 ( .B(\mem_a[10][6] ), .A(\_zyixc_ctx_rdata_29[10][6] ));
Q_ASSIGN U1064 ( .B(\mem_a[10][7] ), .A(\_zyixc_ctx_rdata_29[10][7] ));
Q_ASSIGN U1065 ( .B(\mem_a[10][8] ), .A(\_zyixc_ctx_rdata_29[10][8] ));
Q_ASSIGN U1066 ( .B(\mem_a[10][9] ), .A(\_zyixc_ctx_rdata_29[10][9] ));
Q_ASSIGN U1067 ( .B(\mem_a[10][10] ), .A(\_zyixc_ctx_rdata_29[10][10] ));
Q_ASSIGN U1068 ( .B(\mem_a[10][11] ), .A(\_zyixc_ctx_rdata_29[10][11] ));
Q_ASSIGN U1069 ( .B(\mem_a[10][12] ), .A(\_zyixc_ctx_rdata_29[10][12] ));
Q_ASSIGN U1070 ( .B(\mem_a[10][13] ), .A(\_zyixc_ctx_rdata_29[10][13] ));
Q_ASSIGN U1071 ( .B(\mem_a[10][14] ), .A(\_zyixc_ctx_rdata_29[10][14] ));
Q_ASSIGN U1072 ( .B(\mem_a[10][15] ), .A(\_zyixc_ctx_rdata_29[10][15] ));
Q_ASSIGN U1073 ( .B(\mem_a[10][16] ), .A(\_zyixc_ctx_rdata_29[10][16] ));
Q_ASSIGN U1074 ( .B(\mem_a[10][17] ), .A(\_zyixc_ctx_rdata_29[10][17] ));
Q_ASSIGN U1075 ( .B(\mem_a[10][18] ), .A(\_zyixc_ctx_rdata_29[10][18] ));
Q_ASSIGN U1076 ( .B(\mem_a[10][19] ), .A(\_zyixc_ctx_rdata_29[10][19] ));
Q_ASSIGN U1077 ( .B(\mem_a[10][20] ), .A(\_zyixc_ctx_rdata_29[10][20] ));
Q_ASSIGN U1078 ( .B(\mem_a[10][21] ), .A(\_zyixc_ctx_rdata_29[10][21] ));
Q_ASSIGN U1079 ( .B(\mem_a[10][22] ), .A(\_zyixc_ctx_rdata_29[10][22] ));
Q_ASSIGN U1080 ( .B(\mem_a[10][23] ), .A(\_zyixc_ctx_rdata_29[10][23] ));
Q_ASSIGN U1081 ( .B(\mem_a[10][24] ), .A(\_zyixc_ctx_rdata_29[10][24] ));
Q_ASSIGN U1082 ( .B(\mem_a[10][25] ), .A(\_zyixc_ctx_rdata_29[10][25] ));
Q_ASSIGN U1083 ( .B(\mem_a[10][26] ), .A(\_zyixc_ctx_rdata_29[10][26] ));
Q_ASSIGN U1084 ( .B(\mem_a[10][27] ), .A(\_zyixc_ctx_rdata_29[10][27] ));
Q_ASSIGN U1085 ( .B(\mem_a[10][28] ), .A(\_zyixc_ctx_rdata_29[10][28] ));
Q_ASSIGN U1086 ( .B(\mem_a[10][29] ), .A(\_zyixc_ctx_rdata_29[10][29] ));
Q_ASSIGN U1087 ( .B(\mem_a[10][30] ), .A(\_zyixc_ctx_rdata_29[10][30] ));
Q_ASSIGN U1088 ( .B(\mem_a[10][31] ), .A(\_zyixc_ctx_rdata_29[10][31] ));
Q_ASSIGN U1089 ( .B(\mem_a[10][32] ), .A(\_zyixc_ctx_rdata_29[10][32] ));
Q_ASSIGN U1090 ( .B(\mem_a[10][33] ), .A(\_zyixc_ctx_rdata_29[10][33] ));
Q_ASSIGN U1091 ( .B(\mem_a[10][34] ), .A(\_zyixc_ctx_rdata_29[10][34] ));
Q_ASSIGN U1092 ( .B(\mem_a[10][35] ), .A(\_zyixc_ctx_rdata_29[10][35] ));
Q_ASSIGN U1093 ( .B(\mem_a[10][36] ), .A(\_zyixc_ctx_rdata_29[10][36] ));
Q_ASSIGN U1094 ( .B(\mem_a[10][37] ), .A(\_zyixc_ctx_rdata_29[10][37] ));
Q_ASSIGN U1095 ( .B(\mem_a[10][38] ), .A(\_zyixc_ctx_rdata_29[10][38] ));
Q_ASSIGN U1096 ( .B(\mem_a[10][39] ), .A(\_zyixc_ctx_rdata_29[10][39] ));
Q_ASSIGN U1097 ( .B(\mem_a[10][40] ), .A(\_zyixc_ctx_rdata_29[10][40] ));
Q_ASSIGN U1098 ( .B(\mem_a[10][41] ), .A(\_zyixc_ctx_rdata_29[10][41] ));
Q_ASSIGN U1099 ( .B(\mem_a[10][42] ), .A(\_zyixc_ctx_rdata_29[10][42] ));
Q_ASSIGN U1100 ( .B(\mem_a[10][43] ), .A(\_zyixc_ctx_rdata_29[10][43] ));
Q_ASSIGN U1101 ( .B(\mem_a[10][44] ), .A(\_zyixc_ctx_rdata_29[10][44] ));
Q_ASSIGN U1102 ( .B(\mem_a[10][45] ), .A(\_zyixc_ctx_rdata_29[10][45] ));
Q_ASSIGN U1103 ( .B(\mem_a[10][46] ), .A(\_zyixc_ctx_rdata_29[10][46] ));
Q_ASSIGN U1104 ( .B(\mem_a[10][47] ), .A(\_zyixc_ctx_rdata_29[10][47] ));
Q_ASSIGN U1105 ( .B(\mem_a[10][48] ), .A(\_zyixc_ctx_rdata_29[10][48] ));
Q_ASSIGN U1106 ( .B(\mem_a[10][49] ), .A(\_zyixc_ctx_rdata_29[10][49] ));
Q_ASSIGN U1107 ( .B(\mem_a[10][50] ), .A(\_zyixc_ctx_rdata_29[10][50] ));
Q_ASSIGN U1108 ( .B(\mem_a[10][51] ), .A(\_zyixc_ctx_rdata_29[10][51] ));
Q_ASSIGN U1109 ( .B(\mem_a[10][52] ), .A(\_zyixc_ctx_rdata_29[10][52] ));
Q_ASSIGN U1110 ( .B(\mem_a[10][53] ), .A(\_zyixc_ctx_rdata_29[10][53] ));
Q_ASSIGN U1111 ( .B(\mem_a[10][54] ), .A(\_zyixc_ctx_rdata_29[10][54] ));
Q_ASSIGN U1112 ( .B(\mem_a[10][55] ), .A(\_zyixc_ctx_rdata_29[10][55] ));
Q_ASSIGN U1113 ( .B(\mem_a[10][56] ), .A(\_zyixc_ctx_rdata_29[10][56] ));
Q_ASSIGN U1114 ( .B(\mem_a[10][57] ), .A(\_zyixc_ctx_rdata_29[10][57] ));
Q_ASSIGN U1115 ( .B(\mem_a[10][58] ), .A(\_zyixc_ctx_rdata_29[10][58] ));
Q_ASSIGN U1116 ( .B(\mem_a[10][59] ), .A(\_zyixc_ctx_rdata_29[10][59] ));
Q_ASSIGN U1117 ( .B(\mem_a[10][60] ), .A(\_zyixc_ctx_rdata_29[10][60] ));
Q_ASSIGN U1118 ( .B(\mem_a[10][61] ), .A(\_zyixc_ctx_rdata_29[10][61] ));
Q_ASSIGN U1119 ( .B(\mem_a[10][62] ), .A(\_zyixc_ctx_rdata_29[10][62] ));
Q_ASSIGN U1120 ( .B(\mem_a[10][63] ), .A(\_zyixc_ctx_rdata_29[10][63] ));
Q_ASSIGN U1121 ( .B(\mem_a[11][0] ), .A(\_zyixc_ctx_rdata_29[11][0] ));
Q_ASSIGN U1122 ( .B(\mem_a[11][1] ), .A(\_zyixc_ctx_rdata_29[11][1] ));
Q_ASSIGN U1123 ( .B(\mem_a[11][2] ), .A(\_zyixc_ctx_rdata_29[11][2] ));
Q_ASSIGN U1124 ( .B(\mem_a[11][3] ), .A(\_zyixc_ctx_rdata_29[11][3] ));
Q_ASSIGN U1125 ( .B(\mem_a[11][4] ), .A(\_zyixc_ctx_rdata_29[11][4] ));
Q_ASSIGN U1126 ( .B(\mem_a[11][5] ), .A(\_zyixc_ctx_rdata_29[11][5] ));
Q_ASSIGN U1127 ( .B(\mem_a[11][6] ), .A(\_zyixc_ctx_rdata_29[11][6] ));
Q_ASSIGN U1128 ( .B(\mem_a[11][7] ), .A(\_zyixc_ctx_rdata_29[11][7] ));
Q_ASSIGN U1129 ( .B(\mem_a[11][8] ), .A(\_zyixc_ctx_rdata_29[11][8] ));
Q_ASSIGN U1130 ( .B(\mem_a[11][9] ), .A(\_zyixc_ctx_rdata_29[11][9] ));
Q_ASSIGN U1131 ( .B(\mem_a[11][10] ), .A(\_zyixc_ctx_rdata_29[11][10] ));
Q_ASSIGN U1132 ( .B(\mem_a[11][11] ), .A(\_zyixc_ctx_rdata_29[11][11] ));
Q_ASSIGN U1133 ( .B(\mem_a[11][12] ), .A(\_zyixc_ctx_rdata_29[11][12] ));
Q_ASSIGN U1134 ( .B(\mem_a[11][13] ), .A(\_zyixc_ctx_rdata_29[11][13] ));
Q_ASSIGN U1135 ( .B(\mem_a[11][14] ), .A(\_zyixc_ctx_rdata_29[11][14] ));
Q_ASSIGN U1136 ( .B(\mem_a[11][15] ), .A(\_zyixc_ctx_rdata_29[11][15] ));
Q_ASSIGN U1137 ( .B(\mem_a[11][16] ), .A(\_zyixc_ctx_rdata_29[11][16] ));
Q_ASSIGN U1138 ( .B(\mem_a[11][17] ), .A(\_zyixc_ctx_rdata_29[11][17] ));
Q_ASSIGN U1139 ( .B(\mem_a[11][18] ), .A(\_zyixc_ctx_rdata_29[11][18] ));
Q_ASSIGN U1140 ( .B(\mem_a[11][19] ), .A(\_zyixc_ctx_rdata_29[11][19] ));
Q_ASSIGN U1141 ( .B(\mem_a[11][20] ), .A(\_zyixc_ctx_rdata_29[11][20] ));
Q_ASSIGN U1142 ( .B(\mem_a[11][21] ), .A(\_zyixc_ctx_rdata_29[11][21] ));
Q_ASSIGN U1143 ( .B(\mem_a[11][22] ), .A(\_zyixc_ctx_rdata_29[11][22] ));
Q_ASSIGN U1144 ( .B(\mem_a[11][23] ), .A(\_zyixc_ctx_rdata_29[11][23] ));
Q_ASSIGN U1145 ( .B(\mem_a[11][24] ), .A(\_zyixc_ctx_rdata_29[11][24] ));
Q_ASSIGN U1146 ( .B(\mem_a[11][25] ), .A(\_zyixc_ctx_rdata_29[11][25] ));
Q_ASSIGN U1147 ( .B(\mem_a[11][26] ), .A(\_zyixc_ctx_rdata_29[11][26] ));
Q_ASSIGN U1148 ( .B(\mem_a[11][27] ), .A(\_zyixc_ctx_rdata_29[11][27] ));
Q_ASSIGN U1149 ( .B(\mem_a[11][28] ), .A(\_zyixc_ctx_rdata_29[11][28] ));
Q_ASSIGN U1150 ( .B(\mem_a[11][29] ), .A(\_zyixc_ctx_rdata_29[11][29] ));
Q_ASSIGN U1151 ( .B(\mem_a[11][30] ), .A(\_zyixc_ctx_rdata_29[11][30] ));
Q_ASSIGN U1152 ( .B(\mem_a[11][31] ), .A(\_zyixc_ctx_rdata_29[11][31] ));
Q_ASSIGN U1153 ( .B(\mem_a[11][32] ), .A(\_zyixc_ctx_rdata_29[11][32] ));
Q_ASSIGN U1154 ( .B(\mem_a[11][33] ), .A(\_zyixc_ctx_rdata_29[11][33] ));
Q_ASSIGN U1155 ( .B(\mem_a[11][34] ), .A(\_zyixc_ctx_rdata_29[11][34] ));
Q_ASSIGN U1156 ( .B(\mem_a[11][35] ), .A(\_zyixc_ctx_rdata_29[11][35] ));
Q_ASSIGN U1157 ( .B(\mem_a[11][36] ), .A(\_zyixc_ctx_rdata_29[11][36] ));
Q_ASSIGN U1158 ( .B(\mem_a[11][37] ), .A(\_zyixc_ctx_rdata_29[11][37] ));
Q_ASSIGN U1159 ( .B(\mem_a[11][38] ), .A(\_zyixc_ctx_rdata_29[11][38] ));
Q_ASSIGN U1160 ( .B(\mem_a[11][39] ), .A(\_zyixc_ctx_rdata_29[11][39] ));
Q_ASSIGN U1161 ( .B(\mem_a[11][40] ), .A(\_zyixc_ctx_rdata_29[11][40] ));
Q_ASSIGN U1162 ( .B(\mem_a[11][41] ), .A(\_zyixc_ctx_rdata_29[11][41] ));
Q_ASSIGN U1163 ( .B(\mem_a[11][42] ), .A(\_zyixc_ctx_rdata_29[11][42] ));
Q_ASSIGN U1164 ( .B(\mem_a[11][43] ), .A(\_zyixc_ctx_rdata_29[11][43] ));
Q_ASSIGN U1165 ( .B(\mem_a[11][44] ), .A(\_zyixc_ctx_rdata_29[11][44] ));
Q_ASSIGN U1166 ( .B(\mem_a[11][45] ), .A(\_zyixc_ctx_rdata_29[11][45] ));
Q_ASSIGN U1167 ( .B(\mem_a[11][46] ), .A(\_zyixc_ctx_rdata_29[11][46] ));
Q_ASSIGN U1168 ( .B(\mem_a[11][47] ), .A(\_zyixc_ctx_rdata_29[11][47] ));
Q_ASSIGN U1169 ( .B(\mem_a[11][48] ), .A(\_zyixc_ctx_rdata_29[11][48] ));
Q_ASSIGN U1170 ( .B(\mem_a[11][49] ), .A(\_zyixc_ctx_rdata_29[11][49] ));
Q_ASSIGN U1171 ( .B(\mem_a[11][50] ), .A(\_zyixc_ctx_rdata_29[11][50] ));
Q_ASSIGN U1172 ( .B(\mem_a[11][51] ), .A(\_zyixc_ctx_rdata_29[11][51] ));
Q_ASSIGN U1173 ( .B(\mem_a[11][52] ), .A(\_zyixc_ctx_rdata_29[11][52] ));
Q_ASSIGN U1174 ( .B(\mem_a[11][53] ), .A(\_zyixc_ctx_rdata_29[11][53] ));
Q_ASSIGN U1175 ( .B(\mem_a[11][54] ), .A(\_zyixc_ctx_rdata_29[11][54] ));
Q_ASSIGN U1176 ( .B(\mem_a[11][55] ), .A(\_zyixc_ctx_rdata_29[11][55] ));
Q_ASSIGN U1177 ( .B(\mem_a[11][56] ), .A(\_zyixc_ctx_rdata_29[11][56] ));
Q_ASSIGN U1178 ( .B(\mem_a[11][57] ), .A(\_zyixc_ctx_rdata_29[11][57] ));
Q_ASSIGN U1179 ( .B(\mem_a[11][58] ), .A(\_zyixc_ctx_rdata_29[11][58] ));
Q_ASSIGN U1180 ( .B(\mem_a[11][59] ), .A(\_zyixc_ctx_rdata_29[11][59] ));
Q_ASSIGN U1181 ( .B(\mem_a[11][60] ), .A(\_zyixc_ctx_rdata_29[11][60] ));
Q_ASSIGN U1182 ( .B(\mem_a[11][61] ), .A(\_zyixc_ctx_rdata_29[11][61] ));
Q_ASSIGN U1183 ( .B(\mem_a[11][62] ), .A(\_zyixc_ctx_rdata_29[11][62] ));
Q_ASSIGN U1184 ( .B(\mem_a[11][63] ), .A(\_zyixc_ctx_rdata_29[11][63] ));
Q_ASSIGN U1185 ( .B(\mem_a[12][0] ), .A(\_zyixc_ctx_rdata_29[12][0] ));
Q_ASSIGN U1186 ( .B(\mem_a[12][1] ), .A(\_zyixc_ctx_rdata_29[12][1] ));
Q_ASSIGN U1187 ( .B(\mem_a[12][2] ), .A(\_zyixc_ctx_rdata_29[12][2] ));
Q_ASSIGN U1188 ( .B(\mem_a[12][3] ), .A(\_zyixc_ctx_rdata_29[12][3] ));
Q_ASSIGN U1189 ( .B(\mem_a[12][4] ), .A(\_zyixc_ctx_rdata_29[12][4] ));
Q_ASSIGN U1190 ( .B(\mem_a[12][5] ), .A(\_zyixc_ctx_rdata_29[12][5] ));
Q_ASSIGN U1191 ( .B(\mem_a[12][6] ), .A(\_zyixc_ctx_rdata_29[12][6] ));
Q_ASSIGN U1192 ( .B(\mem_a[12][7] ), .A(\_zyixc_ctx_rdata_29[12][7] ));
Q_ASSIGN U1193 ( .B(\mem_a[12][8] ), .A(\_zyixc_ctx_rdata_29[12][8] ));
Q_ASSIGN U1194 ( .B(\mem_a[12][9] ), .A(\_zyixc_ctx_rdata_29[12][9] ));
Q_ASSIGN U1195 ( .B(\mem_a[12][10] ), .A(\_zyixc_ctx_rdata_29[12][10] ));
Q_ASSIGN U1196 ( .B(\mem_a[12][11] ), .A(\_zyixc_ctx_rdata_29[12][11] ));
Q_ASSIGN U1197 ( .B(\mem_a[12][12] ), .A(\_zyixc_ctx_rdata_29[12][12] ));
Q_ASSIGN U1198 ( .B(\mem_a[12][13] ), .A(\_zyixc_ctx_rdata_29[12][13] ));
Q_ASSIGN U1199 ( .B(\mem_a[12][14] ), .A(\_zyixc_ctx_rdata_29[12][14] ));
Q_ASSIGN U1200 ( .B(\mem_a[12][15] ), .A(\_zyixc_ctx_rdata_29[12][15] ));
Q_ASSIGN U1201 ( .B(\mem_a[12][16] ), .A(\_zyixc_ctx_rdata_29[12][16] ));
Q_ASSIGN U1202 ( .B(\mem_a[12][17] ), .A(\_zyixc_ctx_rdata_29[12][17] ));
Q_ASSIGN U1203 ( .B(\mem_a[12][18] ), .A(\_zyixc_ctx_rdata_29[12][18] ));
Q_ASSIGN U1204 ( .B(\mem_a[12][19] ), .A(\_zyixc_ctx_rdata_29[12][19] ));
Q_ASSIGN U1205 ( .B(\mem_a[12][20] ), .A(\_zyixc_ctx_rdata_29[12][20] ));
Q_ASSIGN U1206 ( .B(\mem_a[12][21] ), .A(\_zyixc_ctx_rdata_29[12][21] ));
Q_ASSIGN U1207 ( .B(\mem_a[12][22] ), .A(\_zyixc_ctx_rdata_29[12][22] ));
Q_ASSIGN U1208 ( .B(\mem_a[12][23] ), .A(\_zyixc_ctx_rdata_29[12][23] ));
Q_ASSIGN U1209 ( .B(\mem_a[12][24] ), .A(\_zyixc_ctx_rdata_29[12][24] ));
Q_ASSIGN U1210 ( .B(\mem_a[12][25] ), .A(\_zyixc_ctx_rdata_29[12][25] ));
Q_ASSIGN U1211 ( .B(\mem_a[12][26] ), .A(\_zyixc_ctx_rdata_29[12][26] ));
Q_ASSIGN U1212 ( .B(\mem_a[12][27] ), .A(\_zyixc_ctx_rdata_29[12][27] ));
Q_ASSIGN U1213 ( .B(\mem_a[12][28] ), .A(\_zyixc_ctx_rdata_29[12][28] ));
Q_ASSIGN U1214 ( .B(\mem_a[12][29] ), .A(\_zyixc_ctx_rdata_29[12][29] ));
Q_ASSIGN U1215 ( .B(\mem_a[12][30] ), .A(\_zyixc_ctx_rdata_29[12][30] ));
Q_ASSIGN U1216 ( .B(\mem_a[12][31] ), .A(\_zyixc_ctx_rdata_29[12][31] ));
Q_ASSIGN U1217 ( .B(\mem_a[12][32] ), .A(\_zyixc_ctx_rdata_29[12][32] ));
Q_ASSIGN U1218 ( .B(\mem_a[12][33] ), .A(\_zyixc_ctx_rdata_29[12][33] ));
Q_ASSIGN U1219 ( .B(\mem_a[12][34] ), .A(\_zyixc_ctx_rdata_29[12][34] ));
Q_ASSIGN U1220 ( .B(\mem_a[12][35] ), .A(\_zyixc_ctx_rdata_29[12][35] ));
Q_ASSIGN U1221 ( .B(\mem_a[12][36] ), .A(\_zyixc_ctx_rdata_29[12][36] ));
Q_ASSIGN U1222 ( .B(\mem_a[12][37] ), .A(\_zyixc_ctx_rdata_29[12][37] ));
Q_ASSIGN U1223 ( .B(\mem_a[12][38] ), .A(\_zyixc_ctx_rdata_29[12][38] ));
Q_ASSIGN U1224 ( .B(\mem_a[12][39] ), .A(\_zyixc_ctx_rdata_29[12][39] ));
Q_ASSIGN U1225 ( .B(\mem_a[12][40] ), .A(\_zyixc_ctx_rdata_29[12][40] ));
Q_ASSIGN U1226 ( .B(\mem_a[12][41] ), .A(\_zyixc_ctx_rdata_29[12][41] ));
Q_ASSIGN U1227 ( .B(\mem_a[12][42] ), .A(\_zyixc_ctx_rdata_29[12][42] ));
Q_ASSIGN U1228 ( .B(\mem_a[12][43] ), .A(\_zyixc_ctx_rdata_29[12][43] ));
Q_ASSIGN U1229 ( .B(\mem_a[12][44] ), .A(\_zyixc_ctx_rdata_29[12][44] ));
Q_ASSIGN U1230 ( .B(\mem_a[12][45] ), .A(\_zyixc_ctx_rdata_29[12][45] ));
Q_ASSIGN U1231 ( .B(\mem_a[12][46] ), .A(\_zyixc_ctx_rdata_29[12][46] ));
Q_ASSIGN U1232 ( .B(\mem_a[12][47] ), .A(\_zyixc_ctx_rdata_29[12][47] ));
Q_ASSIGN U1233 ( .B(\mem_a[12][48] ), .A(\_zyixc_ctx_rdata_29[12][48] ));
Q_ASSIGN U1234 ( .B(\mem_a[12][49] ), .A(\_zyixc_ctx_rdata_29[12][49] ));
Q_ASSIGN U1235 ( .B(\mem_a[12][50] ), .A(\_zyixc_ctx_rdata_29[12][50] ));
Q_ASSIGN U1236 ( .B(\mem_a[12][51] ), .A(\_zyixc_ctx_rdata_29[12][51] ));
Q_ASSIGN U1237 ( .B(\mem_a[12][52] ), .A(\_zyixc_ctx_rdata_29[12][52] ));
Q_ASSIGN U1238 ( .B(\mem_a[12][53] ), .A(\_zyixc_ctx_rdata_29[12][53] ));
Q_ASSIGN U1239 ( .B(\mem_a[12][54] ), .A(\_zyixc_ctx_rdata_29[12][54] ));
Q_ASSIGN U1240 ( .B(\mem_a[12][55] ), .A(\_zyixc_ctx_rdata_29[12][55] ));
Q_ASSIGN U1241 ( .B(\mem_a[12][56] ), .A(\_zyixc_ctx_rdata_29[12][56] ));
Q_ASSIGN U1242 ( .B(\mem_a[12][57] ), .A(\_zyixc_ctx_rdata_29[12][57] ));
Q_ASSIGN U1243 ( .B(\mem_a[12][58] ), .A(\_zyixc_ctx_rdata_29[12][58] ));
Q_ASSIGN U1244 ( .B(\mem_a[12][59] ), .A(\_zyixc_ctx_rdata_29[12][59] ));
Q_ASSIGN U1245 ( .B(\mem_a[12][60] ), .A(\_zyixc_ctx_rdata_29[12][60] ));
Q_ASSIGN U1246 ( .B(\mem_a[12][61] ), .A(\_zyixc_ctx_rdata_29[12][61] ));
Q_ASSIGN U1247 ( .B(\mem_a[12][62] ), .A(\_zyixc_ctx_rdata_29[12][62] ));
Q_ASSIGN U1248 ( .B(\mem_a[12][63] ), .A(\_zyixc_ctx_rdata_29[12][63] ));
Q_ASSIGN U1249 ( .B(\mem_a[13][0] ), .A(\_zyixc_ctx_rdata_29[13][0] ));
Q_ASSIGN U1250 ( .B(\mem_a[13][1] ), .A(\_zyixc_ctx_rdata_29[13][1] ));
Q_ASSIGN U1251 ( .B(\mem_a[13][2] ), .A(\_zyixc_ctx_rdata_29[13][2] ));
Q_ASSIGN U1252 ( .B(\mem_a[13][3] ), .A(\_zyixc_ctx_rdata_29[13][3] ));
Q_ASSIGN U1253 ( .B(\mem_a[13][4] ), .A(\_zyixc_ctx_rdata_29[13][4] ));
Q_ASSIGN U1254 ( .B(\mem_a[13][5] ), .A(\_zyixc_ctx_rdata_29[13][5] ));
Q_ASSIGN U1255 ( .B(\mem_a[13][6] ), .A(\_zyixc_ctx_rdata_29[13][6] ));
Q_ASSIGN U1256 ( .B(\mem_a[13][7] ), .A(\_zyixc_ctx_rdata_29[13][7] ));
Q_ASSIGN U1257 ( .B(\mem_a[13][8] ), .A(\_zyixc_ctx_rdata_29[13][8] ));
Q_ASSIGN U1258 ( .B(\mem_a[13][9] ), .A(\_zyixc_ctx_rdata_29[13][9] ));
Q_ASSIGN U1259 ( .B(\mem_a[13][10] ), .A(\_zyixc_ctx_rdata_29[13][10] ));
Q_ASSIGN U1260 ( .B(\mem_a[13][11] ), .A(\_zyixc_ctx_rdata_29[13][11] ));
Q_ASSIGN U1261 ( .B(\mem_a[13][12] ), .A(\_zyixc_ctx_rdata_29[13][12] ));
Q_ASSIGN U1262 ( .B(\mem_a[13][13] ), .A(\_zyixc_ctx_rdata_29[13][13] ));
Q_ASSIGN U1263 ( .B(\mem_a[13][14] ), .A(\_zyixc_ctx_rdata_29[13][14] ));
Q_ASSIGN U1264 ( .B(\mem_a[13][15] ), .A(\_zyixc_ctx_rdata_29[13][15] ));
Q_ASSIGN U1265 ( .B(\mem_a[13][16] ), .A(\_zyixc_ctx_rdata_29[13][16] ));
Q_ASSIGN U1266 ( .B(\mem_a[13][17] ), .A(\_zyixc_ctx_rdata_29[13][17] ));
Q_ASSIGN U1267 ( .B(\mem_a[13][18] ), .A(\_zyixc_ctx_rdata_29[13][18] ));
Q_ASSIGN U1268 ( .B(\mem_a[13][19] ), .A(\_zyixc_ctx_rdata_29[13][19] ));
Q_ASSIGN U1269 ( .B(\mem_a[13][20] ), .A(\_zyixc_ctx_rdata_29[13][20] ));
Q_ASSIGN U1270 ( .B(\mem_a[13][21] ), .A(\_zyixc_ctx_rdata_29[13][21] ));
Q_ASSIGN U1271 ( .B(\mem_a[13][22] ), .A(\_zyixc_ctx_rdata_29[13][22] ));
Q_ASSIGN U1272 ( .B(\mem_a[13][23] ), .A(\_zyixc_ctx_rdata_29[13][23] ));
Q_ASSIGN U1273 ( .B(\mem_a[13][24] ), .A(\_zyixc_ctx_rdata_29[13][24] ));
Q_ASSIGN U1274 ( .B(\mem_a[13][25] ), .A(\_zyixc_ctx_rdata_29[13][25] ));
Q_ASSIGN U1275 ( .B(\mem_a[13][26] ), .A(\_zyixc_ctx_rdata_29[13][26] ));
Q_ASSIGN U1276 ( .B(\mem_a[13][27] ), .A(\_zyixc_ctx_rdata_29[13][27] ));
Q_ASSIGN U1277 ( .B(\mem_a[13][28] ), .A(\_zyixc_ctx_rdata_29[13][28] ));
Q_ASSIGN U1278 ( .B(\mem_a[13][29] ), .A(\_zyixc_ctx_rdata_29[13][29] ));
Q_ASSIGN U1279 ( .B(\mem_a[13][30] ), .A(\_zyixc_ctx_rdata_29[13][30] ));
Q_ASSIGN U1280 ( .B(\mem_a[13][31] ), .A(\_zyixc_ctx_rdata_29[13][31] ));
Q_ASSIGN U1281 ( .B(\mem_a[13][32] ), .A(\_zyixc_ctx_rdata_29[13][32] ));
Q_ASSIGN U1282 ( .B(\mem_a[13][33] ), .A(\_zyixc_ctx_rdata_29[13][33] ));
Q_ASSIGN U1283 ( .B(\mem_a[13][34] ), .A(\_zyixc_ctx_rdata_29[13][34] ));
Q_ASSIGN U1284 ( .B(\mem_a[13][35] ), .A(\_zyixc_ctx_rdata_29[13][35] ));
Q_ASSIGN U1285 ( .B(\mem_a[13][36] ), .A(\_zyixc_ctx_rdata_29[13][36] ));
Q_ASSIGN U1286 ( .B(\mem_a[13][37] ), .A(\_zyixc_ctx_rdata_29[13][37] ));
Q_ASSIGN U1287 ( .B(\mem_a[13][38] ), .A(\_zyixc_ctx_rdata_29[13][38] ));
Q_ASSIGN U1288 ( .B(\mem_a[13][39] ), .A(\_zyixc_ctx_rdata_29[13][39] ));
Q_ASSIGN U1289 ( .B(\mem_a[13][40] ), .A(\_zyixc_ctx_rdata_29[13][40] ));
Q_ASSIGN U1290 ( .B(\mem_a[13][41] ), .A(\_zyixc_ctx_rdata_29[13][41] ));
Q_ASSIGN U1291 ( .B(\mem_a[13][42] ), .A(\_zyixc_ctx_rdata_29[13][42] ));
Q_ASSIGN U1292 ( .B(\mem_a[13][43] ), .A(\_zyixc_ctx_rdata_29[13][43] ));
Q_ASSIGN U1293 ( .B(\mem_a[13][44] ), .A(\_zyixc_ctx_rdata_29[13][44] ));
Q_ASSIGN U1294 ( .B(\mem_a[13][45] ), .A(\_zyixc_ctx_rdata_29[13][45] ));
Q_ASSIGN U1295 ( .B(\mem_a[13][46] ), .A(\_zyixc_ctx_rdata_29[13][46] ));
Q_ASSIGN U1296 ( .B(\mem_a[13][47] ), .A(\_zyixc_ctx_rdata_29[13][47] ));
Q_ASSIGN U1297 ( .B(\mem_a[13][48] ), .A(\_zyixc_ctx_rdata_29[13][48] ));
Q_ASSIGN U1298 ( .B(\mem_a[13][49] ), .A(\_zyixc_ctx_rdata_29[13][49] ));
Q_ASSIGN U1299 ( .B(\mem_a[13][50] ), .A(\_zyixc_ctx_rdata_29[13][50] ));
Q_ASSIGN U1300 ( .B(\mem_a[13][51] ), .A(\_zyixc_ctx_rdata_29[13][51] ));
Q_ASSIGN U1301 ( .B(\mem_a[13][52] ), .A(\_zyixc_ctx_rdata_29[13][52] ));
Q_ASSIGN U1302 ( .B(\mem_a[13][53] ), .A(\_zyixc_ctx_rdata_29[13][53] ));
Q_ASSIGN U1303 ( .B(\mem_a[13][54] ), .A(\_zyixc_ctx_rdata_29[13][54] ));
Q_ASSIGN U1304 ( .B(\mem_a[13][55] ), .A(\_zyixc_ctx_rdata_29[13][55] ));
Q_ASSIGN U1305 ( .B(\mem_a[13][56] ), .A(\_zyixc_ctx_rdata_29[13][56] ));
Q_ASSIGN U1306 ( .B(\mem_a[13][57] ), .A(\_zyixc_ctx_rdata_29[13][57] ));
Q_ASSIGN U1307 ( .B(\mem_a[13][58] ), .A(\_zyixc_ctx_rdata_29[13][58] ));
Q_ASSIGN U1308 ( .B(\mem_a[13][59] ), .A(\_zyixc_ctx_rdata_29[13][59] ));
Q_ASSIGN U1309 ( .B(\mem_a[13][60] ), .A(\_zyixc_ctx_rdata_29[13][60] ));
Q_ASSIGN U1310 ( .B(\mem_a[13][61] ), .A(\_zyixc_ctx_rdata_29[13][61] ));
Q_ASSIGN U1311 ( .B(\mem_a[13][62] ), .A(\_zyixc_ctx_rdata_29[13][62] ));
Q_ASSIGN U1312 ( .B(\mem_a[13][63] ), .A(\_zyixc_ctx_rdata_29[13][63] ));
Q_ASSIGN U1313 ( .B(\mem_a[14][0] ), .A(\_zyixc_ctx_rdata_29[14][0] ));
Q_ASSIGN U1314 ( .B(\mem_a[14][1] ), .A(\_zyixc_ctx_rdata_29[14][1] ));
Q_ASSIGN U1315 ( .B(\mem_a[14][2] ), .A(\_zyixc_ctx_rdata_29[14][2] ));
Q_ASSIGN U1316 ( .B(\mem_a[14][3] ), .A(\_zyixc_ctx_rdata_29[14][3] ));
Q_ASSIGN U1317 ( .B(\mem_a[14][4] ), .A(\_zyixc_ctx_rdata_29[14][4] ));
Q_ASSIGN U1318 ( .B(\mem_a[14][5] ), .A(\_zyixc_ctx_rdata_29[14][5] ));
Q_ASSIGN U1319 ( .B(\mem_a[14][6] ), .A(\_zyixc_ctx_rdata_29[14][6] ));
Q_ASSIGN U1320 ( .B(\mem_a[14][7] ), .A(\_zyixc_ctx_rdata_29[14][7] ));
Q_ASSIGN U1321 ( .B(\mem_a[14][8] ), .A(\_zyixc_ctx_rdata_29[14][8] ));
Q_ASSIGN U1322 ( .B(\mem_a[14][9] ), .A(\_zyixc_ctx_rdata_29[14][9] ));
Q_ASSIGN U1323 ( .B(\mem_a[14][10] ), .A(\_zyixc_ctx_rdata_29[14][10] ));
Q_ASSIGN U1324 ( .B(\mem_a[14][11] ), .A(\_zyixc_ctx_rdata_29[14][11] ));
Q_ASSIGN U1325 ( .B(\mem_a[14][12] ), .A(\_zyixc_ctx_rdata_29[14][12] ));
Q_ASSIGN U1326 ( .B(\mem_a[14][13] ), .A(\_zyixc_ctx_rdata_29[14][13] ));
Q_ASSIGN U1327 ( .B(\mem_a[14][14] ), .A(\_zyixc_ctx_rdata_29[14][14] ));
Q_ASSIGN U1328 ( .B(\mem_a[14][15] ), .A(\_zyixc_ctx_rdata_29[14][15] ));
Q_ASSIGN U1329 ( .B(\mem_a[14][16] ), .A(\_zyixc_ctx_rdata_29[14][16] ));
Q_ASSIGN U1330 ( .B(\mem_a[14][17] ), .A(\_zyixc_ctx_rdata_29[14][17] ));
Q_ASSIGN U1331 ( .B(\mem_a[14][18] ), .A(\_zyixc_ctx_rdata_29[14][18] ));
Q_ASSIGN U1332 ( .B(\mem_a[14][19] ), .A(\_zyixc_ctx_rdata_29[14][19] ));
Q_ASSIGN U1333 ( .B(\mem_a[14][20] ), .A(\_zyixc_ctx_rdata_29[14][20] ));
Q_ASSIGN U1334 ( .B(\mem_a[14][21] ), .A(\_zyixc_ctx_rdata_29[14][21] ));
Q_ASSIGN U1335 ( .B(\mem_a[14][22] ), .A(\_zyixc_ctx_rdata_29[14][22] ));
Q_ASSIGN U1336 ( .B(\mem_a[14][23] ), .A(\_zyixc_ctx_rdata_29[14][23] ));
Q_ASSIGN U1337 ( .B(\mem_a[14][24] ), .A(\_zyixc_ctx_rdata_29[14][24] ));
Q_ASSIGN U1338 ( .B(\mem_a[14][25] ), .A(\_zyixc_ctx_rdata_29[14][25] ));
Q_ASSIGN U1339 ( .B(\mem_a[14][26] ), .A(\_zyixc_ctx_rdata_29[14][26] ));
Q_ASSIGN U1340 ( .B(\mem_a[14][27] ), .A(\_zyixc_ctx_rdata_29[14][27] ));
Q_ASSIGN U1341 ( .B(\mem_a[14][28] ), .A(\_zyixc_ctx_rdata_29[14][28] ));
Q_ASSIGN U1342 ( .B(\mem_a[14][29] ), .A(\_zyixc_ctx_rdata_29[14][29] ));
Q_ASSIGN U1343 ( .B(\mem_a[14][30] ), .A(\_zyixc_ctx_rdata_29[14][30] ));
Q_ASSIGN U1344 ( .B(\mem_a[14][31] ), .A(\_zyixc_ctx_rdata_29[14][31] ));
Q_ASSIGN U1345 ( .B(\mem_a[14][32] ), .A(\_zyixc_ctx_rdata_29[14][32] ));
Q_ASSIGN U1346 ( .B(\mem_a[14][33] ), .A(\_zyixc_ctx_rdata_29[14][33] ));
Q_ASSIGN U1347 ( .B(\mem_a[14][34] ), .A(\_zyixc_ctx_rdata_29[14][34] ));
Q_ASSIGN U1348 ( .B(\mem_a[14][35] ), .A(\_zyixc_ctx_rdata_29[14][35] ));
Q_ASSIGN U1349 ( .B(\mem_a[14][36] ), .A(\_zyixc_ctx_rdata_29[14][36] ));
Q_ASSIGN U1350 ( .B(\mem_a[14][37] ), .A(\_zyixc_ctx_rdata_29[14][37] ));
Q_ASSIGN U1351 ( .B(\mem_a[14][38] ), .A(\_zyixc_ctx_rdata_29[14][38] ));
Q_ASSIGN U1352 ( .B(\mem_a[14][39] ), .A(\_zyixc_ctx_rdata_29[14][39] ));
Q_ASSIGN U1353 ( .B(\mem_a[14][40] ), .A(\_zyixc_ctx_rdata_29[14][40] ));
Q_ASSIGN U1354 ( .B(\mem_a[14][41] ), .A(\_zyixc_ctx_rdata_29[14][41] ));
Q_ASSIGN U1355 ( .B(\mem_a[14][42] ), .A(\_zyixc_ctx_rdata_29[14][42] ));
Q_ASSIGN U1356 ( .B(\mem_a[14][43] ), .A(\_zyixc_ctx_rdata_29[14][43] ));
Q_ASSIGN U1357 ( .B(\mem_a[14][44] ), .A(\_zyixc_ctx_rdata_29[14][44] ));
Q_ASSIGN U1358 ( .B(\mem_a[14][45] ), .A(\_zyixc_ctx_rdata_29[14][45] ));
Q_ASSIGN U1359 ( .B(\mem_a[14][46] ), .A(\_zyixc_ctx_rdata_29[14][46] ));
Q_ASSIGN U1360 ( .B(\mem_a[14][47] ), .A(\_zyixc_ctx_rdata_29[14][47] ));
Q_ASSIGN U1361 ( .B(\mem_a[14][48] ), .A(\_zyixc_ctx_rdata_29[14][48] ));
Q_ASSIGN U1362 ( .B(\mem_a[14][49] ), .A(\_zyixc_ctx_rdata_29[14][49] ));
Q_ASSIGN U1363 ( .B(\mem_a[14][50] ), .A(\_zyixc_ctx_rdata_29[14][50] ));
Q_ASSIGN U1364 ( .B(\mem_a[14][51] ), .A(\_zyixc_ctx_rdata_29[14][51] ));
Q_ASSIGN U1365 ( .B(\mem_a[14][52] ), .A(\_zyixc_ctx_rdata_29[14][52] ));
Q_ASSIGN U1366 ( .B(\mem_a[14][53] ), .A(\_zyixc_ctx_rdata_29[14][53] ));
Q_ASSIGN U1367 ( .B(\mem_a[14][54] ), .A(\_zyixc_ctx_rdata_29[14][54] ));
Q_ASSIGN U1368 ( .B(\mem_a[14][55] ), .A(\_zyixc_ctx_rdata_29[14][55] ));
Q_ASSIGN U1369 ( .B(\mem_a[14][56] ), .A(\_zyixc_ctx_rdata_29[14][56] ));
Q_ASSIGN U1370 ( .B(\mem_a[14][57] ), .A(\_zyixc_ctx_rdata_29[14][57] ));
Q_ASSIGN U1371 ( .B(\mem_a[14][58] ), .A(\_zyixc_ctx_rdata_29[14][58] ));
Q_ASSIGN U1372 ( .B(\mem_a[14][59] ), .A(\_zyixc_ctx_rdata_29[14][59] ));
Q_ASSIGN U1373 ( .B(\mem_a[14][60] ), .A(\_zyixc_ctx_rdata_29[14][60] ));
Q_ASSIGN U1374 ( .B(\mem_a[14][61] ), .A(\_zyixc_ctx_rdata_29[14][61] ));
Q_ASSIGN U1375 ( .B(\mem_a[14][62] ), .A(\_zyixc_ctx_rdata_29[14][62] ));
Q_ASSIGN U1376 ( .B(\mem_a[14][63] ), .A(\_zyixc_ctx_rdata_29[14][63] ));
Q_ASSIGN U1377 ( .B(\mem_a[15][0] ), .A(\_zyixc_ctx_rdata_29[15][0] ));
Q_ASSIGN U1378 ( .B(\mem_a[15][1] ), .A(\_zyixc_ctx_rdata_29[15][1] ));
Q_ASSIGN U1379 ( .B(\mem_a[15][2] ), .A(\_zyixc_ctx_rdata_29[15][2] ));
Q_ASSIGN U1380 ( .B(\mem_a[15][3] ), .A(\_zyixc_ctx_rdata_29[15][3] ));
Q_ASSIGN U1381 ( .B(\mem_a[15][4] ), .A(\_zyixc_ctx_rdata_29[15][4] ));
Q_ASSIGN U1382 ( .B(\mem_a[15][5] ), .A(\_zyixc_ctx_rdata_29[15][5] ));
Q_ASSIGN U1383 ( .B(\mem_a[15][6] ), .A(\_zyixc_ctx_rdata_29[15][6] ));
Q_ASSIGN U1384 ( .B(\mem_a[15][7] ), .A(\_zyixc_ctx_rdata_29[15][7] ));
Q_ASSIGN U1385 ( .B(\mem_a[15][8] ), .A(\_zyixc_ctx_rdata_29[15][8] ));
Q_ASSIGN U1386 ( .B(\mem_a[15][9] ), .A(\_zyixc_ctx_rdata_29[15][9] ));
Q_ASSIGN U1387 ( .B(\mem_a[15][10] ), .A(\_zyixc_ctx_rdata_29[15][10] ));
Q_ASSIGN U1388 ( .B(\mem_a[15][11] ), .A(\_zyixc_ctx_rdata_29[15][11] ));
Q_ASSIGN U1389 ( .B(\mem_a[15][12] ), .A(\_zyixc_ctx_rdata_29[15][12] ));
Q_ASSIGN U1390 ( .B(\mem_a[15][13] ), .A(\_zyixc_ctx_rdata_29[15][13] ));
Q_ASSIGN U1391 ( .B(\mem_a[15][14] ), .A(\_zyixc_ctx_rdata_29[15][14] ));
Q_ASSIGN U1392 ( .B(\mem_a[15][15] ), .A(\_zyixc_ctx_rdata_29[15][15] ));
Q_ASSIGN U1393 ( .B(\mem_a[15][16] ), .A(\_zyixc_ctx_rdata_29[15][16] ));
Q_ASSIGN U1394 ( .B(\mem_a[15][17] ), .A(\_zyixc_ctx_rdata_29[15][17] ));
Q_ASSIGN U1395 ( .B(\mem_a[15][18] ), .A(\_zyixc_ctx_rdata_29[15][18] ));
Q_ASSIGN U1396 ( .B(\mem_a[15][19] ), .A(\_zyixc_ctx_rdata_29[15][19] ));
Q_ASSIGN U1397 ( .B(\mem_a[15][20] ), .A(\_zyixc_ctx_rdata_29[15][20] ));
Q_ASSIGN U1398 ( .B(\mem_a[15][21] ), .A(\_zyixc_ctx_rdata_29[15][21] ));
Q_ASSIGN U1399 ( .B(\mem_a[15][22] ), .A(\_zyixc_ctx_rdata_29[15][22] ));
Q_ASSIGN U1400 ( .B(\mem_a[15][23] ), .A(\_zyixc_ctx_rdata_29[15][23] ));
Q_ASSIGN U1401 ( .B(\mem_a[15][24] ), .A(\_zyixc_ctx_rdata_29[15][24] ));
Q_ASSIGN U1402 ( .B(\mem_a[15][25] ), .A(\_zyixc_ctx_rdata_29[15][25] ));
Q_ASSIGN U1403 ( .B(\mem_a[15][26] ), .A(\_zyixc_ctx_rdata_29[15][26] ));
Q_ASSIGN U1404 ( .B(\mem_a[15][27] ), .A(\_zyixc_ctx_rdata_29[15][27] ));
Q_ASSIGN U1405 ( .B(\mem_a[15][28] ), .A(\_zyixc_ctx_rdata_29[15][28] ));
Q_ASSIGN U1406 ( .B(\mem_a[15][29] ), .A(\_zyixc_ctx_rdata_29[15][29] ));
Q_ASSIGN U1407 ( .B(\mem_a[15][30] ), .A(\_zyixc_ctx_rdata_29[15][30] ));
Q_ASSIGN U1408 ( .B(\mem_a[15][31] ), .A(\_zyixc_ctx_rdata_29[15][31] ));
Q_ASSIGN U1409 ( .B(\mem_a[15][32] ), .A(\_zyixc_ctx_rdata_29[15][32] ));
Q_ASSIGN U1410 ( .B(\mem_a[15][33] ), .A(\_zyixc_ctx_rdata_29[15][33] ));
Q_ASSIGN U1411 ( .B(\mem_a[15][34] ), .A(\_zyixc_ctx_rdata_29[15][34] ));
Q_ASSIGN U1412 ( .B(\mem_a[15][35] ), .A(\_zyixc_ctx_rdata_29[15][35] ));
Q_ASSIGN U1413 ( .B(\mem_a[15][36] ), .A(\_zyixc_ctx_rdata_29[15][36] ));
Q_ASSIGN U1414 ( .B(\mem_a[15][37] ), .A(\_zyixc_ctx_rdata_29[15][37] ));
Q_ASSIGN U1415 ( .B(\mem_a[15][38] ), .A(\_zyixc_ctx_rdata_29[15][38] ));
Q_ASSIGN U1416 ( .B(\mem_a[15][39] ), .A(\_zyixc_ctx_rdata_29[15][39] ));
Q_ASSIGN U1417 ( .B(\mem_a[15][40] ), .A(\_zyixc_ctx_rdata_29[15][40] ));
Q_ASSIGN U1418 ( .B(\mem_a[15][41] ), .A(\_zyixc_ctx_rdata_29[15][41] ));
Q_ASSIGN U1419 ( .B(\mem_a[15][42] ), .A(\_zyixc_ctx_rdata_29[15][42] ));
Q_ASSIGN U1420 ( .B(\mem_a[15][43] ), .A(\_zyixc_ctx_rdata_29[15][43] ));
Q_ASSIGN U1421 ( .B(\mem_a[15][44] ), .A(\_zyixc_ctx_rdata_29[15][44] ));
Q_ASSIGN U1422 ( .B(\mem_a[15][45] ), .A(\_zyixc_ctx_rdata_29[15][45] ));
Q_ASSIGN U1423 ( .B(\mem_a[15][46] ), .A(\_zyixc_ctx_rdata_29[15][46] ));
Q_ASSIGN U1424 ( .B(\mem_a[15][47] ), .A(\_zyixc_ctx_rdata_29[15][47] ));
Q_ASSIGN U1425 ( .B(\mem_a[15][48] ), .A(\_zyixc_ctx_rdata_29[15][48] ));
Q_ASSIGN U1426 ( .B(\mem_a[15][49] ), .A(\_zyixc_ctx_rdata_29[15][49] ));
Q_ASSIGN U1427 ( .B(\mem_a[15][50] ), .A(\_zyixc_ctx_rdata_29[15][50] ));
Q_ASSIGN U1428 ( .B(\mem_a[15][51] ), .A(\_zyixc_ctx_rdata_29[15][51] ));
Q_ASSIGN U1429 ( .B(\mem_a[15][52] ), .A(\_zyixc_ctx_rdata_29[15][52] ));
Q_ASSIGN U1430 ( .B(\mem_a[15][53] ), .A(\_zyixc_ctx_rdata_29[15][53] ));
Q_ASSIGN U1431 ( .B(\mem_a[15][54] ), .A(\_zyixc_ctx_rdata_29[15][54] ));
Q_ASSIGN U1432 ( .B(\mem_a[15][55] ), .A(\_zyixc_ctx_rdata_29[15][55] ));
Q_ASSIGN U1433 ( .B(\mem_a[15][56] ), .A(\_zyixc_ctx_rdata_29[15][56] ));
Q_ASSIGN U1434 ( .B(\mem_a[15][57] ), .A(\_zyixc_ctx_rdata_29[15][57] ));
Q_ASSIGN U1435 ( .B(\mem_a[15][58] ), .A(\_zyixc_ctx_rdata_29[15][58] ));
Q_ASSIGN U1436 ( .B(\mem_a[15][59] ), .A(\_zyixc_ctx_rdata_29[15][59] ));
Q_ASSIGN U1437 ( .B(\mem_a[15][60] ), .A(\_zyixc_ctx_rdata_29[15][60] ));
Q_ASSIGN U1438 ( .B(\mem_a[15][61] ), .A(\_zyixc_ctx_rdata_29[15][61] ));
Q_ASSIGN U1439 ( .B(\mem_a[15][62] ), .A(\_zyixc_ctx_rdata_29[15][62] ));
Q_ASSIGN U1440 ( .B(\mem_a[15][63] ), .A(\_zyixc_ctx_rdata_29[15][63] ));
Q_ASSIGN U1441 ( .B(\mem_a[16][0] ), .A(\_zyixc_ctx_rdata_29[16][0] ));
Q_ASSIGN U1442 ( .B(\mem_a[16][1] ), .A(\_zyixc_ctx_rdata_29[16][1] ));
Q_ASSIGN U1443 ( .B(\mem_a[16][2] ), .A(\_zyixc_ctx_rdata_29[16][2] ));
Q_ASSIGN U1444 ( .B(\mem_a[16][3] ), .A(\_zyixc_ctx_rdata_29[16][3] ));
Q_ASSIGN U1445 ( .B(\mem_a[16][4] ), .A(\_zyixc_ctx_rdata_29[16][4] ));
Q_ASSIGN U1446 ( .B(\mem_a[16][5] ), .A(\_zyixc_ctx_rdata_29[16][5] ));
Q_ASSIGN U1447 ( .B(\mem_a[16][6] ), .A(\_zyixc_ctx_rdata_29[16][6] ));
Q_ASSIGN U1448 ( .B(\mem_a[16][7] ), .A(\_zyixc_ctx_rdata_29[16][7] ));
Q_ASSIGN U1449 ( .B(\mem_a[16][8] ), .A(\_zyixc_ctx_rdata_29[16][8] ));
Q_ASSIGN U1450 ( .B(\mem_a[16][9] ), .A(\_zyixc_ctx_rdata_29[16][9] ));
Q_ASSIGN U1451 ( .B(\mem_a[16][10] ), .A(\_zyixc_ctx_rdata_29[16][10] ));
Q_ASSIGN U1452 ( .B(\mem_a[16][11] ), .A(\_zyixc_ctx_rdata_29[16][11] ));
Q_ASSIGN U1453 ( .B(\mem_a[16][12] ), .A(\_zyixc_ctx_rdata_29[16][12] ));
Q_ASSIGN U1454 ( .B(\mem_a[16][13] ), .A(\_zyixc_ctx_rdata_29[16][13] ));
Q_ASSIGN U1455 ( .B(\mem_a[16][14] ), .A(\_zyixc_ctx_rdata_29[16][14] ));
Q_ASSIGN U1456 ( .B(\mem_a[16][15] ), .A(\_zyixc_ctx_rdata_29[16][15] ));
Q_ASSIGN U1457 ( .B(\mem_a[16][16] ), .A(\_zyixc_ctx_rdata_29[16][16] ));
Q_ASSIGN U1458 ( .B(\mem_a[16][17] ), .A(\_zyixc_ctx_rdata_29[16][17] ));
Q_ASSIGN U1459 ( .B(\mem_a[16][18] ), .A(\_zyixc_ctx_rdata_29[16][18] ));
Q_ASSIGN U1460 ( .B(\mem_a[16][19] ), .A(\_zyixc_ctx_rdata_29[16][19] ));
Q_ASSIGN U1461 ( .B(\mem_a[16][20] ), .A(\_zyixc_ctx_rdata_29[16][20] ));
Q_ASSIGN U1462 ( .B(\mem_a[16][21] ), .A(\_zyixc_ctx_rdata_29[16][21] ));
Q_ASSIGN U1463 ( .B(\mem_a[16][22] ), .A(\_zyixc_ctx_rdata_29[16][22] ));
Q_ASSIGN U1464 ( .B(\mem_a[16][23] ), .A(\_zyixc_ctx_rdata_29[16][23] ));
Q_ASSIGN U1465 ( .B(\mem_a[16][24] ), .A(\_zyixc_ctx_rdata_29[16][24] ));
Q_ASSIGN U1466 ( .B(\mem_a[16][25] ), .A(\_zyixc_ctx_rdata_29[16][25] ));
Q_ASSIGN U1467 ( .B(\mem_a[16][26] ), .A(\_zyixc_ctx_rdata_29[16][26] ));
Q_ASSIGN U1468 ( .B(\mem_a[16][27] ), .A(\_zyixc_ctx_rdata_29[16][27] ));
Q_ASSIGN U1469 ( .B(\mem_a[16][28] ), .A(\_zyixc_ctx_rdata_29[16][28] ));
Q_ASSIGN U1470 ( .B(\mem_a[16][29] ), .A(\_zyixc_ctx_rdata_29[16][29] ));
Q_ASSIGN U1471 ( .B(\mem_a[16][30] ), .A(\_zyixc_ctx_rdata_29[16][30] ));
Q_ASSIGN U1472 ( .B(\mem_a[16][31] ), .A(\_zyixc_ctx_rdata_29[16][31] ));
Q_ASSIGN U1473 ( .B(\mem_a[16][32] ), .A(\_zyixc_ctx_rdata_29[16][32] ));
Q_ASSIGN U1474 ( .B(\mem_a[16][33] ), .A(\_zyixc_ctx_rdata_29[16][33] ));
Q_ASSIGN U1475 ( .B(\mem_a[16][34] ), .A(\_zyixc_ctx_rdata_29[16][34] ));
Q_ASSIGN U1476 ( .B(\mem_a[16][35] ), .A(\_zyixc_ctx_rdata_29[16][35] ));
Q_ASSIGN U1477 ( .B(\mem_a[16][36] ), .A(\_zyixc_ctx_rdata_29[16][36] ));
Q_ASSIGN U1478 ( .B(\mem_a[16][37] ), .A(\_zyixc_ctx_rdata_29[16][37] ));
Q_ASSIGN U1479 ( .B(\mem_a[16][38] ), .A(\_zyixc_ctx_rdata_29[16][38] ));
Q_ASSIGN U1480 ( .B(\mem_a[16][39] ), .A(\_zyixc_ctx_rdata_29[16][39] ));
Q_ASSIGN U1481 ( .B(\mem_a[16][40] ), .A(\_zyixc_ctx_rdata_29[16][40] ));
Q_ASSIGN U1482 ( .B(\mem_a[16][41] ), .A(\_zyixc_ctx_rdata_29[16][41] ));
Q_ASSIGN U1483 ( .B(\mem_a[16][42] ), .A(\_zyixc_ctx_rdata_29[16][42] ));
Q_ASSIGN U1484 ( .B(\mem_a[16][43] ), .A(\_zyixc_ctx_rdata_29[16][43] ));
Q_ASSIGN U1485 ( .B(\mem_a[16][44] ), .A(\_zyixc_ctx_rdata_29[16][44] ));
Q_ASSIGN U1486 ( .B(\mem_a[16][45] ), .A(\_zyixc_ctx_rdata_29[16][45] ));
Q_ASSIGN U1487 ( .B(\mem_a[16][46] ), .A(\_zyixc_ctx_rdata_29[16][46] ));
Q_ASSIGN U1488 ( .B(\mem_a[16][47] ), .A(\_zyixc_ctx_rdata_29[16][47] ));
Q_ASSIGN U1489 ( .B(\mem_a[16][48] ), .A(\_zyixc_ctx_rdata_29[16][48] ));
Q_ASSIGN U1490 ( .B(\mem_a[16][49] ), .A(\_zyixc_ctx_rdata_29[16][49] ));
Q_ASSIGN U1491 ( .B(\mem_a[16][50] ), .A(\_zyixc_ctx_rdata_29[16][50] ));
Q_ASSIGN U1492 ( .B(\mem_a[16][51] ), .A(\_zyixc_ctx_rdata_29[16][51] ));
Q_ASSIGN U1493 ( .B(\mem_a[16][52] ), .A(\_zyixc_ctx_rdata_29[16][52] ));
Q_ASSIGN U1494 ( .B(\mem_a[16][53] ), .A(\_zyixc_ctx_rdata_29[16][53] ));
Q_ASSIGN U1495 ( .B(\mem_a[16][54] ), .A(\_zyixc_ctx_rdata_29[16][54] ));
Q_ASSIGN U1496 ( .B(\mem_a[16][55] ), .A(\_zyixc_ctx_rdata_29[16][55] ));
Q_ASSIGN U1497 ( .B(\mem_a[16][56] ), .A(\_zyixc_ctx_rdata_29[16][56] ));
Q_ASSIGN U1498 ( .B(\mem_a[16][57] ), .A(\_zyixc_ctx_rdata_29[16][57] ));
Q_ASSIGN U1499 ( .B(\mem_a[16][58] ), .A(\_zyixc_ctx_rdata_29[16][58] ));
Q_ASSIGN U1500 ( .B(\mem_a[16][59] ), .A(\_zyixc_ctx_rdata_29[16][59] ));
Q_ASSIGN U1501 ( .B(\mem_a[16][60] ), .A(\_zyixc_ctx_rdata_29[16][60] ));
Q_ASSIGN U1502 ( .B(\mem_a[16][61] ), .A(\_zyixc_ctx_rdata_29[16][61] ));
Q_ASSIGN U1503 ( .B(\mem_a[16][62] ), .A(\_zyixc_ctx_rdata_29[16][62] ));
Q_ASSIGN U1504 ( .B(\mem_a[16][63] ), .A(\_zyixc_ctx_rdata_29[16][63] ));
Q_ASSIGN U1505 ( .B(\mem_a[17][0] ), .A(\_zyixc_ctx_rdata_29[17][0] ));
Q_ASSIGN U1506 ( .B(\mem_a[17][1] ), .A(\_zyixc_ctx_rdata_29[17][1] ));
Q_ASSIGN U1507 ( .B(\mem_a[17][2] ), .A(\_zyixc_ctx_rdata_29[17][2] ));
Q_ASSIGN U1508 ( .B(\mem_a[17][3] ), .A(\_zyixc_ctx_rdata_29[17][3] ));
Q_ASSIGN U1509 ( .B(\mem_a[17][4] ), .A(\_zyixc_ctx_rdata_29[17][4] ));
Q_ASSIGN U1510 ( .B(\mem_a[17][5] ), .A(\_zyixc_ctx_rdata_29[17][5] ));
Q_ASSIGN U1511 ( .B(\mem_a[17][6] ), .A(\_zyixc_ctx_rdata_29[17][6] ));
Q_ASSIGN U1512 ( .B(\mem_a[17][7] ), .A(\_zyixc_ctx_rdata_29[17][7] ));
Q_ASSIGN U1513 ( .B(\mem_a[17][8] ), .A(\_zyixc_ctx_rdata_29[17][8] ));
Q_ASSIGN U1514 ( .B(\mem_a[17][9] ), .A(\_zyixc_ctx_rdata_29[17][9] ));
Q_ASSIGN U1515 ( .B(\mem_a[17][10] ), .A(\_zyixc_ctx_rdata_29[17][10] ));
Q_ASSIGN U1516 ( .B(\mem_a[17][11] ), .A(\_zyixc_ctx_rdata_29[17][11] ));
Q_ASSIGN U1517 ( .B(\mem_a[17][12] ), .A(\_zyixc_ctx_rdata_29[17][12] ));
Q_ASSIGN U1518 ( .B(\mem_a[17][13] ), .A(\_zyixc_ctx_rdata_29[17][13] ));
Q_ASSIGN U1519 ( .B(\mem_a[17][14] ), .A(\_zyixc_ctx_rdata_29[17][14] ));
Q_ASSIGN U1520 ( .B(\mem_a[17][15] ), .A(\_zyixc_ctx_rdata_29[17][15] ));
Q_ASSIGN U1521 ( .B(\mem_a[17][16] ), .A(\_zyixc_ctx_rdata_29[17][16] ));
Q_ASSIGN U1522 ( .B(\mem_a[17][17] ), .A(\_zyixc_ctx_rdata_29[17][17] ));
Q_ASSIGN U1523 ( .B(\mem_a[17][18] ), .A(\_zyixc_ctx_rdata_29[17][18] ));
Q_ASSIGN U1524 ( .B(\mem_a[17][19] ), .A(\_zyixc_ctx_rdata_29[17][19] ));
Q_ASSIGN U1525 ( .B(\mem_a[17][20] ), .A(\_zyixc_ctx_rdata_29[17][20] ));
Q_ASSIGN U1526 ( .B(\mem_a[17][21] ), .A(\_zyixc_ctx_rdata_29[17][21] ));
Q_ASSIGN U1527 ( .B(\mem_a[17][22] ), .A(\_zyixc_ctx_rdata_29[17][22] ));
Q_ASSIGN U1528 ( .B(\mem_a[17][23] ), .A(\_zyixc_ctx_rdata_29[17][23] ));
Q_ASSIGN U1529 ( .B(\mem_a[17][24] ), .A(\_zyixc_ctx_rdata_29[17][24] ));
Q_ASSIGN U1530 ( .B(\mem_a[17][25] ), .A(\_zyixc_ctx_rdata_29[17][25] ));
Q_ASSIGN U1531 ( .B(\mem_a[17][26] ), .A(\_zyixc_ctx_rdata_29[17][26] ));
Q_ASSIGN U1532 ( .B(\mem_a[17][27] ), .A(\_zyixc_ctx_rdata_29[17][27] ));
Q_ASSIGN U1533 ( .B(\mem_a[17][28] ), .A(\_zyixc_ctx_rdata_29[17][28] ));
Q_ASSIGN U1534 ( .B(\mem_a[17][29] ), .A(\_zyixc_ctx_rdata_29[17][29] ));
Q_ASSIGN U1535 ( .B(\mem_a[17][30] ), .A(\_zyixc_ctx_rdata_29[17][30] ));
Q_ASSIGN U1536 ( .B(\mem_a[17][31] ), .A(\_zyixc_ctx_rdata_29[17][31] ));
Q_ASSIGN U1537 ( .B(\mem_a[17][32] ), .A(\_zyixc_ctx_rdata_29[17][32] ));
Q_ASSIGN U1538 ( .B(\mem_a[17][33] ), .A(\_zyixc_ctx_rdata_29[17][33] ));
Q_ASSIGN U1539 ( .B(\mem_a[17][34] ), .A(\_zyixc_ctx_rdata_29[17][34] ));
Q_ASSIGN U1540 ( .B(\mem_a[17][35] ), .A(\_zyixc_ctx_rdata_29[17][35] ));
Q_ASSIGN U1541 ( .B(\mem_a[17][36] ), .A(\_zyixc_ctx_rdata_29[17][36] ));
Q_ASSIGN U1542 ( .B(\mem_a[17][37] ), .A(\_zyixc_ctx_rdata_29[17][37] ));
Q_ASSIGN U1543 ( .B(\mem_a[17][38] ), .A(\_zyixc_ctx_rdata_29[17][38] ));
Q_ASSIGN U1544 ( .B(\mem_a[17][39] ), .A(\_zyixc_ctx_rdata_29[17][39] ));
Q_ASSIGN U1545 ( .B(\mem_a[17][40] ), .A(\_zyixc_ctx_rdata_29[17][40] ));
Q_ASSIGN U1546 ( .B(\mem_a[17][41] ), .A(\_zyixc_ctx_rdata_29[17][41] ));
Q_ASSIGN U1547 ( .B(\mem_a[17][42] ), .A(\_zyixc_ctx_rdata_29[17][42] ));
Q_ASSIGN U1548 ( .B(\mem_a[17][43] ), .A(\_zyixc_ctx_rdata_29[17][43] ));
Q_ASSIGN U1549 ( .B(\mem_a[17][44] ), .A(\_zyixc_ctx_rdata_29[17][44] ));
Q_ASSIGN U1550 ( .B(\mem_a[17][45] ), .A(\_zyixc_ctx_rdata_29[17][45] ));
Q_ASSIGN U1551 ( .B(\mem_a[17][46] ), .A(\_zyixc_ctx_rdata_29[17][46] ));
Q_ASSIGN U1552 ( .B(\mem_a[17][47] ), .A(\_zyixc_ctx_rdata_29[17][47] ));
Q_ASSIGN U1553 ( .B(\mem_a[17][48] ), .A(\_zyixc_ctx_rdata_29[17][48] ));
Q_ASSIGN U1554 ( .B(\mem_a[17][49] ), .A(\_zyixc_ctx_rdata_29[17][49] ));
Q_ASSIGN U1555 ( .B(\mem_a[17][50] ), .A(\_zyixc_ctx_rdata_29[17][50] ));
Q_ASSIGN U1556 ( .B(\mem_a[17][51] ), .A(\_zyixc_ctx_rdata_29[17][51] ));
Q_ASSIGN U1557 ( .B(\mem_a[17][52] ), .A(\_zyixc_ctx_rdata_29[17][52] ));
Q_ASSIGN U1558 ( .B(\mem_a[17][53] ), .A(\_zyixc_ctx_rdata_29[17][53] ));
Q_ASSIGN U1559 ( .B(\mem_a[17][54] ), .A(\_zyixc_ctx_rdata_29[17][54] ));
Q_ASSIGN U1560 ( .B(\mem_a[17][55] ), .A(\_zyixc_ctx_rdata_29[17][55] ));
Q_ASSIGN U1561 ( .B(\mem_a[17][56] ), .A(\_zyixc_ctx_rdata_29[17][56] ));
Q_ASSIGN U1562 ( .B(\mem_a[17][57] ), .A(\_zyixc_ctx_rdata_29[17][57] ));
Q_ASSIGN U1563 ( .B(\mem_a[17][58] ), .A(\_zyixc_ctx_rdata_29[17][58] ));
Q_ASSIGN U1564 ( .B(\mem_a[17][59] ), .A(\_zyixc_ctx_rdata_29[17][59] ));
Q_ASSIGN U1565 ( .B(\mem_a[17][60] ), .A(\_zyixc_ctx_rdata_29[17][60] ));
Q_ASSIGN U1566 ( .B(\mem_a[17][61] ), .A(\_zyixc_ctx_rdata_29[17][61] ));
Q_ASSIGN U1567 ( .B(\mem_a[17][62] ), .A(\_zyixc_ctx_rdata_29[17][62] ));
Q_ASSIGN U1568 ( .B(\mem_a[17][63] ), .A(\_zyixc_ctx_rdata_29[17][63] ));
Q_ASSIGN U1569 ( .B(\mem_a[18][0] ), .A(\_zyixc_ctx_rdata_29[18][0] ));
Q_ASSIGN U1570 ( .B(\mem_a[18][1] ), .A(\_zyixc_ctx_rdata_29[18][1] ));
Q_ASSIGN U1571 ( .B(\mem_a[18][2] ), .A(\_zyixc_ctx_rdata_29[18][2] ));
Q_ASSIGN U1572 ( .B(\mem_a[18][3] ), .A(\_zyixc_ctx_rdata_29[18][3] ));
Q_ASSIGN U1573 ( .B(\mem_a[18][4] ), .A(\_zyixc_ctx_rdata_29[18][4] ));
Q_ASSIGN U1574 ( .B(\mem_a[18][5] ), .A(\_zyixc_ctx_rdata_29[18][5] ));
Q_ASSIGN U1575 ( .B(\mem_a[18][6] ), .A(\_zyixc_ctx_rdata_29[18][6] ));
Q_ASSIGN U1576 ( .B(\mem_a[18][7] ), .A(\_zyixc_ctx_rdata_29[18][7] ));
Q_ASSIGN U1577 ( .B(\mem_a[18][8] ), .A(\_zyixc_ctx_rdata_29[18][8] ));
Q_ASSIGN U1578 ( .B(\mem_a[18][9] ), .A(\_zyixc_ctx_rdata_29[18][9] ));
Q_ASSIGN U1579 ( .B(\mem_a[18][10] ), .A(\_zyixc_ctx_rdata_29[18][10] ));
Q_ASSIGN U1580 ( .B(\mem_a[18][11] ), .A(\_zyixc_ctx_rdata_29[18][11] ));
Q_ASSIGN U1581 ( .B(\mem_a[18][12] ), .A(\_zyixc_ctx_rdata_29[18][12] ));
Q_ASSIGN U1582 ( .B(\mem_a[18][13] ), .A(\_zyixc_ctx_rdata_29[18][13] ));
Q_ASSIGN U1583 ( .B(\mem_a[18][14] ), .A(\_zyixc_ctx_rdata_29[18][14] ));
Q_ASSIGN U1584 ( .B(\mem_a[18][15] ), .A(\_zyixc_ctx_rdata_29[18][15] ));
Q_ASSIGN U1585 ( .B(\mem_a[18][16] ), .A(\_zyixc_ctx_rdata_29[18][16] ));
Q_ASSIGN U1586 ( .B(\mem_a[18][17] ), .A(\_zyixc_ctx_rdata_29[18][17] ));
Q_ASSIGN U1587 ( .B(\mem_a[18][18] ), .A(\_zyixc_ctx_rdata_29[18][18] ));
Q_ASSIGN U1588 ( .B(\mem_a[18][19] ), .A(\_zyixc_ctx_rdata_29[18][19] ));
Q_ASSIGN U1589 ( .B(\mem_a[18][20] ), .A(\_zyixc_ctx_rdata_29[18][20] ));
Q_ASSIGN U1590 ( .B(\mem_a[18][21] ), .A(\_zyixc_ctx_rdata_29[18][21] ));
Q_ASSIGN U1591 ( .B(\mem_a[18][22] ), .A(\_zyixc_ctx_rdata_29[18][22] ));
Q_ASSIGN U1592 ( .B(\mem_a[18][23] ), .A(\_zyixc_ctx_rdata_29[18][23] ));
Q_ASSIGN U1593 ( .B(\mem_a[18][24] ), .A(\_zyixc_ctx_rdata_29[18][24] ));
Q_ASSIGN U1594 ( .B(\mem_a[18][25] ), .A(\_zyixc_ctx_rdata_29[18][25] ));
Q_ASSIGN U1595 ( .B(\mem_a[18][26] ), .A(\_zyixc_ctx_rdata_29[18][26] ));
Q_ASSIGN U1596 ( .B(\mem_a[18][27] ), .A(\_zyixc_ctx_rdata_29[18][27] ));
Q_ASSIGN U1597 ( .B(\mem_a[18][28] ), .A(\_zyixc_ctx_rdata_29[18][28] ));
Q_ASSIGN U1598 ( .B(\mem_a[18][29] ), .A(\_zyixc_ctx_rdata_29[18][29] ));
Q_ASSIGN U1599 ( .B(\mem_a[18][30] ), .A(\_zyixc_ctx_rdata_29[18][30] ));
Q_ASSIGN U1600 ( .B(\mem_a[18][31] ), .A(\_zyixc_ctx_rdata_29[18][31] ));
Q_ASSIGN U1601 ( .B(\mem_a[18][32] ), .A(\_zyixc_ctx_rdata_29[18][32] ));
Q_ASSIGN U1602 ( .B(\mem_a[18][33] ), .A(\_zyixc_ctx_rdata_29[18][33] ));
Q_ASSIGN U1603 ( .B(\mem_a[18][34] ), .A(\_zyixc_ctx_rdata_29[18][34] ));
Q_ASSIGN U1604 ( .B(\mem_a[18][35] ), .A(\_zyixc_ctx_rdata_29[18][35] ));
Q_ASSIGN U1605 ( .B(\mem_a[18][36] ), .A(\_zyixc_ctx_rdata_29[18][36] ));
Q_ASSIGN U1606 ( .B(\mem_a[18][37] ), .A(\_zyixc_ctx_rdata_29[18][37] ));
Q_ASSIGN U1607 ( .B(\mem_a[18][38] ), .A(\_zyixc_ctx_rdata_29[18][38] ));
Q_ASSIGN U1608 ( .B(\mem_a[18][39] ), .A(\_zyixc_ctx_rdata_29[18][39] ));
Q_ASSIGN U1609 ( .B(\mem_a[18][40] ), .A(\_zyixc_ctx_rdata_29[18][40] ));
Q_ASSIGN U1610 ( .B(\mem_a[18][41] ), .A(\_zyixc_ctx_rdata_29[18][41] ));
Q_ASSIGN U1611 ( .B(\mem_a[18][42] ), .A(\_zyixc_ctx_rdata_29[18][42] ));
Q_ASSIGN U1612 ( .B(\mem_a[18][43] ), .A(\_zyixc_ctx_rdata_29[18][43] ));
Q_ASSIGN U1613 ( .B(\mem_a[18][44] ), .A(\_zyixc_ctx_rdata_29[18][44] ));
Q_ASSIGN U1614 ( .B(\mem_a[18][45] ), .A(\_zyixc_ctx_rdata_29[18][45] ));
Q_ASSIGN U1615 ( .B(\mem_a[18][46] ), .A(\_zyixc_ctx_rdata_29[18][46] ));
Q_ASSIGN U1616 ( .B(\mem_a[18][47] ), .A(\_zyixc_ctx_rdata_29[18][47] ));
Q_ASSIGN U1617 ( .B(\mem_a[18][48] ), .A(\_zyixc_ctx_rdata_29[18][48] ));
Q_ASSIGN U1618 ( .B(\mem_a[18][49] ), .A(\_zyixc_ctx_rdata_29[18][49] ));
Q_ASSIGN U1619 ( .B(\mem_a[18][50] ), .A(\_zyixc_ctx_rdata_29[18][50] ));
Q_ASSIGN U1620 ( .B(\mem_a[18][51] ), .A(\_zyixc_ctx_rdata_29[18][51] ));
Q_ASSIGN U1621 ( .B(\mem_a[18][52] ), .A(\_zyixc_ctx_rdata_29[18][52] ));
Q_ASSIGN U1622 ( .B(\mem_a[18][53] ), .A(\_zyixc_ctx_rdata_29[18][53] ));
Q_ASSIGN U1623 ( .B(\mem_a[18][54] ), .A(\_zyixc_ctx_rdata_29[18][54] ));
Q_ASSIGN U1624 ( .B(\mem_a[18][55] ), .A(\_zyixc_ctx_rdata_29[18][55] ));
Q_ASSIGN U1625 ( .B(\mem_a[18][56] ), .A(\_zyixc_ctx_rdata_29[18][56] ));
Q_ASSIGN U1626 ( .B(\mem_a[18][57] ), .A(\_zyixc_ctx_rdata_29[18][57] ));
Q_ASSIGN U1627 ( .B(\mem_a[18][58] ), .A(\_zyixc_ctx_rdata_29[18][58] ));
Q_ASSIGN U1628 ( .B(\mem_a[18][59] ), .A(\_zyixc_ctx_rdata_29[18][59] ));
Q_ASSIGN U1629 ( .B(\mem_a[18][60] ), .A(\_zyixc_ctx_rdata_29[18][60] ));
Q_ASSIGN U1630 ( .B(\mem_a[18][61] ), .A(\_zyixc_ctx_rdata_29[18][61] ));
Q_ASSIGN U1631 ( .B(\mem_a[18][62] ), .A(\_zyixc_ctx_rdata_29[18][62] ));
Q_ASSIGN U1632 ( .B(\mem_a[18][63] ), .A(\_zyixc_ctx_rdata_29[18][63] ));
Q_ASSIGN U1633 ( .B(\mem_a[19][0] ), .A(\_zyixc_ctx_rdata_29[19][0] ));
Q_ASSIGN U1634 ( .B(\mem_a[19][1] ), .A(\_zyixc_ctx_rdata_29[19][1] ));
Q_ASSIGN U1635 ( .B(\mem_a[19][2] ), .A(\_zyixc_ctx_rdata_29[19][2] ));
Q_ASSIGN U1636 ( .B(\mem_a[19][3] ), .A(\_zyixc_ctx_rdata_29[19][3] ));
Q_ASSIGN U1637 ( .B(\mem_a[19][4] ), .A(\_zyixc_ctx_rdata_29[19][4] ));
Q_ASSIGN U1638 ( .B(\mem_a[19][5] ), .A(\_zyixc_ctx_rdata_29[19][5] ));
Q_ASSIGN U1639 ( .B(\mem_a[19][6] ), .A(\_zyixc_ctx_rdata_29[19][6] ));
Q_ASSIGN U1640 ( .B(\mem_a[19][7] ), .A(\_zyixc_ctx_rdata_29[19][7] ));
Q_ASSIGN U1641 ( .B(\mem_a[19][8] ), .A(\_zyixc_ctx_rdata_29[19][8] ));
Q_ASSIGN U1642 ( .B(\mem_a[19][9] ), .A(\_zyixc_ctx_rdata_29[19][9] ));
Q_ASSIGN U1643 ( .B(\mem_a[19][10] ), .A(\_zyixc_ctx_rdata_29[19][10] ));
Q_ASSIGN U1644 ( .B(\mem_a[19][11] ), .A(\_zyixc_ctx_rdata_29[19][11] ));
Q_ASSIGN U1645 ( .B(\mem_a[19][12] ), .A(\_zyixc_ctx_rdata_29[19][12] ));
Q_ASSIGN U1646 ( .B(\mem_a[19][13] ), .A(\_zyixc_ctx_rdata_29[19][13] ));
Q_ASSIGN U1647 ( .B(\mem_a[19][14] ), .A(\_zyixc_ctx_rdata_29[19][14] ));
Q_ASSIGN U1648 ( .B(\mem_a[19][15] ), .A(\_zyixc_ctx_rdata_29[19][15] ));
Q_ASSIGN U1649 ( .B(\mem_a[19][16] ), .A(\_zyixc_ctx_rdata_29[19][16] ));
Q_ASSIGN U1650 ( .B(\mem_a[19][17] ), .A(\_zyixc_ctx_rdata_29[19][17] ));
Q_ASSIGN U1651 ( .B(\mem_a[19][18] ), .A(\_zyixc_ctx_rdata_29[19][18] ));
Q_ASSIGN U1652 ( .B(\mem_a[19][19] ), .A(\_zyixc_ctx_rdata_29[19][19] ));
Q_ASSIGN U1653 ( .B(\mem_a[19][20] ), .A(\_zyixc_ctx_rdata_29[19][20] ));
Q_ASSIGN U1654 ( .B(\mem_a[19][21] ), .A(\_zyixc_ctx_rdata_29[19][21] ));
Q_ASSIGN U1655 ( .B(\mem_a[19][22] ), .A(\_zyixc_ctx_rdata_29[19][22] ));
Q_ASSIGN U1656 ( .B(\mem_a[19][23] ), .A(\_zyixc_ctx_rdata_29[19][23] ));
Q_ASSIGN U1657 ( .B(\mem_a[19][24] ), .A(\_zyixc_ctx_rdata_29[19][24] ));
Q_ASSIGN U1658 ( .B(\mem_a[19][25] ), .A(\_zyixc_ctx_rdata_29[19][25] ));
Q_ASSIGN U1659 ( .B(\mem_a[19][26] ), .A(\_zyixc_ctx_rdata_29[19][26] ));
Q_ASSIGN U1660 ( .B(\mem_a[19][27] ), .A(\_zyixc_ctx_rdata_29[19][27] ));
Q_ASSIGN U1661 ( .B(\mem_a[19][28] ), .A(\_zyixc_ctx_rdata_29[19][28] ));
Q_ASSIGN U1662 ( .B(\mem_a[19][29] ), .A(\_zyixc_ctx_rdata_29[19][29] ));
Q_ASSIGN U1663 ( .B(\mem_a[19][30] ), .A(\_zyixc_ctx_rdata_29[19][30] ));
Q_ASSIGN U1664 ( .B(\mem_a[19][31] ), .A(\_zyixc_ctx_rdata_29[19][31] ));
Q_ASSIGN U1665 ( .B(\mem_a[19][32] ), .A(\_zyixc_ctx_rdata_29[19][32] ));
Q_ASSIGN U1666 ( .B(\mem_a[19][33] ), .A(\_zyixc_ctx_rdata_29[19][33] ));
Q_ASSIGN U1667 ( .B(\mem_a[19][34] ), .A(\_zyixc_ctx_rdata_29[19][34] ));
Q_ASSIGN U1668 ( .B(\mem_a[19][35] ), .A(\_zyixc_ctx_rdata_29[19][35] ));
Q_ASSIGN U1669 ( .B(\mem_a[19][36] ), .A(\_zyixc_ctx_rdata_29[19][36] ));
Q_ASSIGN U1670 ( .B(\mem_a[19][37] ), .A(\_zyixc_ctx_rdata_29[19][37] ));
Q_ASSIGN U1671 ( .B(\mem_a[19][38] ), .A(\_zyixc_ctx_rdata_29[19][38] ));
Q_ASSIGN U1672 ( .B(\mem_a[19][39] ), .A(\_zyixc_ctx_rdata_29[19][39] ));
Q_ASSIGN U1673 ( .B(\mem_a[19][40] ), .A(\_zyixc_ctx_rdata_29[19][40] ));
Q_ASSIGN U1674 ( .B(\mem_a[19][41] ), .A(\_zyixc_ctx_rdata_29[19][41] ));
Q_ASSIGN U1675 ( .B(\mem_a[19][42] ), .A(\_zyixc_ctx_rdata_29[19][42] ));
Q_ASSIGN U1676 ( .B(\mem_a[19][43] ), .A(\_zyixc_ctx_rdata_29[19][43] ));
Q_ASSIGN U1677 ( .B(\mem_a[19][44] ), .A(\_zyixc_ctx_rdata_29[19][44] ));
Q_ASSIGN U1678 ( .B(\mem_a[19][45] ), .A(\_zyixc_ctx_rdata_29[19][45] ));
Q_ASSIGN U1679 ( .B(\mem_a[19][46] ), .A(\_zyixc_ctx_rdata_29[19][46] ));
Q_ASSIGN U1680 ( .B(\mem_a[19][47] ), .A(\_zyixc_ctx_rdata_29[19][47] ));
Q_ASSIGN U1681 ( .B(\mem_a[19][48] ), .A(\_zyixc_ctx_rdata_29[19][48] ));
Q_ASSIGN U1682 ( .B(\mem_a[19][49] ), .A(\_zyixc_ctx_rdata_29[19][49] ));
Q_ASSIGN U1683 ( .B(\mem_a[19][50] ), .A(\_zyixc_ctx_rdata_29[19][50] ));
Q_ASSIGN U1684 ( .B(\mem_a[19][51] ), .A(\_zyixc_ctx_rdata_29[19][51] ));
Q_ASSIGN U1685 ( .B(\mem_a[19][52] ), .A(\_zyixc_ctx_rdata_29[19][52] ));
Q_ASSIGN U1686 ( .B(\mem_a[19][53] ), .A(\_zyixc_ctx_rdata_29[19][53] ));
Q_ASSIGN U1687 ( .B(\mem_a[19][54] ), .A(\_zyixc_ctx_rdata_29[19][54] ));
Q_ASSIGN U1688 ( .B(\mem_a[19][55] ), .A(\_zyixc_ctx_rdata_29[19][55] ));
Q_ASSIGN U1689 ( .B(\mem_a[19][56] ), .A(\_zyixc_ctx_rdata_29[19][56] ));
Q_ASSIGN U1690 ( .B(\mem_a[19][57] ), .A(\_zyixc_ctx_rdata_29[19][57] ));
Q_ASSIGN U1691 ( .B(\mem_a[19][58] ), .A(\_zyixc_ctx_rdata_29[19][58] ));
Q_ASSIGN U1692 ( .B(\mem_a[19][59] ), .A(\_zyixc_ctx_rdata_29[19][59] ));
Q_ASSIGN U1693 ( .B(\mem_a[19][60] ), .A(\_zyixc_ctx_rdata_29[19][60] ));
Q_ASSIGN U1694 ( .B(\mem_a[19][61] ), .A(\_zyixc_ctx_rdata_29[19][61] ));
Q_ASSIGN U1695 ( .B(\mem_a[19][62] ), .A(\_zyixc_ctx_rdata_29[19][62] ));
Q_ASSIGN U1696 ( .B(\mem_a[19][63] ), .A(\_zyixc_ctx_rdata_29[19][63] ));
Q_ASSIGN U1697 ( .B(\mem_a[20][0] ), .A(\_zyixc_ctx_rdata_29[20][0] ));
Q_ASSIGN U1698 ( .B(\mem_a[20][1] ), .A(\_zyixc_ctx_rdata_29[20][1] ));
Q_ASSIGN U1699 ( .B(\mem_a[20][2] ), .A(\_zyixc_ctx_rdata_29[20][2] ));
Q_ASSIGN U1700 ( .B(\mem_a[20][3] ), .A(\_zyixc_ctx_rdata_29[20][3] ));
Q_ASSIGN U1701 ( .B(\mem_a[20][4] ), .A(\_zyixc_ctx_rdata_29[20][4] ));
Q_ASSIGN U1702 ( .B(\mem_a[20][5] ), .A(\_zyixc_ctx_rdata_29[20][5] ));
Q_ASSIGN U1703 ( .B(\mem_a[20][6] ), .A(\_zyixc_ctx_rdata_29[20][6] ));
Q_ASSIGN U1704 ( .B(\mem_a[20][7] ), .A(\_zyixc_ctx_rdata_29[20][7] ));
Q_ASSIGN U1705 ( .B(\mem_a[20][8] ), .A(\_zyixc_ctx_rdata_29[20][8] ));
Q_ASSIGN U1706 ( .B(\mem_a[20][9] ), .A(\_zyixc_ctx_rdata_29[20][9] ));
Q_ASSIGN U1707 ( .B(\mem_a[20][10] ), .A(\_zyixc_ctx_rdata_29[20][10] ));
Q_ASSIGN U1708 ( .B(\mem_a[20][11] ), .A(\_zyixc_ctx_rdata_29[20][11] ));
Q_ASSIGN U1709 ( .B(\mem_a[20][12] ), .A(\_zyixc_ctx_rdata_29[20][12] ));
Q_ASSIGN U1710 ( .B(\mem_a[20][13] ), .A(\_zyixc_ctx_rdata_29[20][13] ));
Q_ASSIGN U1711 ( .B(\mem_a[20][14] ), .A(\_zyixc_ctx_rdata_29[20][14] ));
Q_ASSIGN U1712 ( .B(\mem_a[20][15] ), .A(\_zyixc_ctx_rdata_29[20][15] ));
Q_ASSIGN U1713 ( .B(\mem_a[20][16] ), .A(\_zyixc_ctx_rdata_29[20][16] ));
Q_ASSIGN U1714 ( .B(\mem_a[20][17] ), .A(\_zyixc_ctx_rdata_29[20][17] ));
Q_ASSIGN U1715 ( .B(\mem_a[20][18] ), .A(\_zyixc_ctx_rdata_29[20][18] ));
Q_ASSIGN U1716 ( .B(\mem_a[20][19] ), .A(\_zyixc_ctx_rdata_29[20][19] ));
Q_ASSIGN U1717 ( .B(\mem_a[20][20] ), .A(\_zyixc_ctx_rdata_29[20][20] ));
Q_ASSIGN U1718 ( .B(\mem_a[20][21] ), .A(\_zyixc_ctx_rdata_29[20][21] ));
Q_ASSIGN U1719 ( .B(\mem_a[20][22] ), .A(\_zyixc_ctx_rdata_29[20][22] ));
Q_ASSIGN U1720 ( .B(\mem_a[20][23] ), .A(\_zyixc_ctx_rdata_29[20][23] ));
Q_ASSIGN U1721 ( .B(\mem_a[20][24] ), .A(\_zyixc_ctx_rdata_29[20][24] ));
Q_ASSIGN U1722 ( .B(\mem_a[20][25] ), .A(\_zyixc_ctx_rdata_29[20][25] ));
Q_ASSIGN U1723 ( .B(\mem_a[20][26] ), .A(\_zyixc_ctx_rdata_29[20][26] ));
Q_ASSIGN U1724 ( .B(\mem_a[20][27] ), .A(\_zyixc_ctx_rdata_29[20][27] ));
Q_ASSIGN U1725 ( .B(\mem_a[20][28] ), .A(\_zyixc_ctx_rdata_29[20][28] ));
Q_ASSIGN U1726 ( .B(\mem_a[20][29] ), .A(\_zyixc_ctx_rdata_29[20][29] ));
Q_ASSIGN U1727 ( .B(\mem_a[20][30] ), .A(\_zyixc_ctx_rdata_29[20][30] ));
Q_ASSIGN U1728 ( .B(\mem_a[20][31] ), .A(\_zyixc_ctx_rdata_29[20][31] ));
Q_ASSIGN U1729 ( .B(\mem_a[20][32] ), .A(\_zyixc_ctx_rdata_29[20][32] ));
Q_ASSIGN U1730 ( .B(\mem_a[20][33] ), .A(\_zyixc_ctx_rdata_29[20][33] ));
Q_ASSIGN U1731 ( .B(\mem_a[20][34] ), .A(\_zyixc_ctx_rdata_29[20][34] ));
Q_ASSIGN U1732 ( .B(\mem_a[20][35] ), .A(\_zyixc_ctx_rdata_29[20][35] ));
Q_ASSIGN U1733 ( .B(\mem_a[20][36] ), .A(\_zyixc_ctx_rdata_29[20][36] ));
Q_ASSIGN U1734 ( .B(\mem_a[20][37] ), .A(\_zyixc_ctx_rdata_29[20][37] ));
Q_ASSIGN U1735 ( .B(\mem_a[20][38] ), .A(\_zyixc_ctx_rdata_29[20][38] ));
Q_ASSIGN U1736 ( .B(\mem_a[20][39] ), .A(\_zyixc_ctx_rdata_29[20][39] ));
Q_ASSIGN U1737 ( .B(\mem_a[20][40] ), .A(\_zyixc_ctx_rdata_29[20][40] ));
Q_ASSIGN U1738 ( .B(\mem_a[20][41] ), .A(\_zyixc_ctx_rdata_29[20][41] ));
Q_ASSIGN U1739 ( .B(\mem_a[20][42] ), .A(\_zyixc_ctx_rdata_29[20][42] ));
Q_ASSIGN U1740 ( .B(\mem_a[20][43] ), .A(\_zyixc_ctx_rdata_29[20][43] ));
Q_ASSIGN U1741 ( .B(\mem_a[20][44] ), .A(\_zyixc_ctx_rdata_29[20][44] ));
Q_ASSIGN U1742 ( .B(\mem_a[20][45] ), .A(\_zyixc_ctx_rdata_29[20][45] ));
Q_ASSIGN U1743 ( .B(\mem_a[20][46] ), .A(\_zyixc_ctx_rdata_29[20][46] ));
Q_ASSIGN U1744 ( .B(\mem_a[20][47] ), .A(\_zyixc_ctx_rdata_29[20][47] ));
Q_ASSIGN U1745 ( .B(\mem_a[20][48] ), .A(\_zyixc_ctx_rdata_29[20][48] ));
Q_ASSIGN U1746 ( .B(\mem_a[20][49] ), .A(\_zyixc_ctx_rdata_29[20][49] ));
Q_ASSIGN U1747 ( .B(\mem_a[20][50] ), .A(\_zyixc_ctx_rdata_29[20][50] ));
Q_ASSIGN U1748 ( .B(\mem_a[20][51] ), .A(\_zyixc_ctx_rdata_29[20][51] ));
Q_ASSIGN U1749 ( .B(\mem_a[20][52] ), .A(\_zyixc_ctx_rdata_29[20][52] ));
Q_ASSIGN U1750 ( .B(\mem_a[20][53] ), .A(\_zyixc_ctx_rdata_29[20][53] ));
Q_ASSIGN U1751 ( .B(\mem_a[20][54] ), .A(\_zyixc_ctx_rdata_29[20][54] ));
Q_ASSIGN U1752 ( .B(\mem_a[20][55] ), .A(\_zyixc_ctx_rdata_29[20][55] ));
Q_ASSIGN U1753 ( .B(\mem_a[20][56] ), .A(\_zyixc_ctx_rdata_29[20][56] ));
Q_ASSIGN U1754 ( .B(\mem_a[20][57] ), .A(\_zyixc_ctx_rdata_29[20][57] ));
Q_ASSIGN U1755 ( .B(\mem_a[20][58] ), .A(\_zyixc_ctx_rdata_29[20][58] ));
Q_ASSIGN U1756 ( .B(\mem_a[20][59] ), .A(\_zyixc_ctx_rdata_29[20][59] ));
Q_ASSIGN U1757 ( .B(\mem_a[20][60] ), .A(\_zyixc_ctx_rdata_29[20][60] ));
Q_ASSIGN U1758 ( .B(\mem_a[20][61] ), .A(\_zyixc_ctx_rdata_29[20][61] ));
Q_ASSIGN U1759 ( .B(\mem_a[20][62] ), .A(\_zyixc_ctx_rdata_29[20][62] ));
Q_ASSIGN U1760 ( .B(\mem_a[20][63] ), .A(\_zyixc_ctx_rdata_29[20][63] ));
Q_ASSIGN U1761 ( .B(\mem_a[21][0] ), .A(\_zyixc_ctx_rdata_29[21][0] ));
Q_ASSIGN U1762 ( .B(\mem_a[21][1] ), .A(\_zyixc_ctx_rdata_29[21][1] ));
Q_ASSIGN U1763 ( .B(\mem_a[21][2] ), .A(\_zyixc_ctx_rdata_29[21][2] ));
Q_ASSIGN U1764 ( .B(\mem_a[21][3] ), .A(\_zyixc_ctx_rdata_29[21][3] ));
Q_ASSIGN U1765 ( .B(\mem_a[21][4] ), .A(\_zyixc_ctx_rdata_29[21][4] ));
Q_ASSIGN U1766 ( .B(\mem_a[21][5] ), .A(\_zyixc_ctx_rdata_29[21][5] ));
Q_ASSIGN U1767 ( .B(\mem_a[21][6] ), .A(\_zyixc_ctx_rdata_29[21][6] ));
Q_ASSIGN U1768 ( .B(\mem_a[21][7] ), .A(\_zyixc_ctx_rdata_29[21][7] ));
Q_ASSIGN U1769 ( .B(\mem_a[21][8] ), .A(\_zyixc_ctx_rdata_29[21][8] ));
Q_ASSIGN U1770 ( .B(\mem_a[21][9] ), .A(\_zyixc_ctx_rdata_29[21][9] ));
Q_ASSIGN U1771 ( .B(\mem_a[21][10] ), .A(\_zyixc_ctx_rdata_29[21][10] ));
Q_ASSIGN U1772 ( .B(\mem_a[21][11] ), .A(\_zyixc_ctx_rdata_29[21][11] ));
Q_ASSIGN U1773 ( .B(\mem_a[21][12] ), .A(\_zyixc_ctx_rdata_29[21][12] ));
Q_ASSIGN U1774 ( .B(\mem_a[21][13] ), .A(\_zyixc_ctx_rdata_29[21][13] ));
Q_ASSIGN U1775 ( .B(\mem_a[21][14] ), .A(\_zyixc_ctx_rdata_29[21][14] ));
Q_ASSIGN U1776 ( .B(\mem_a[21][15] ), .A(\_zyixc_ctx_rdata_29[21][15] ));
Q_ASSIGN U1777 ( .B(\mem_a[21][16] ), .A(\_zyixc_ctx_rdata_29[21][16] ));
Q_ASSIGN U1778 ( .B(\mem_a[21][17] ), .A(\_zyixc_ctx_rdata_29[21][17] ));
Q_ASSIGN U1779 ( .B(\mem_a[21][18] ), .A(\_zyixc_ctx_rdata_29[21][18] ));
Q_ASSIGN U1780 ( .B(\mem_a[21][19] ), .A(\_zyixc_ctx_rdata_29[21][19] ));
Q_ASSIGN U1781 ( .B(\mem_a[21][20] ), .A(\_zyixc_ctx_rdata_29[21][20] ));
Q_ASSIGN U1782 ( .B(\mem_a[21][21] ), .A(\_zyixc_ctx_rdata_29[21][21] ));
Q_ASSIGN U1783 ( .B(\mem_a[21][22] ), .A(\_zyixc_ctx_rdata_29[21][22] ));
Q_ASSIGN U1784 ( .B(\mem_a[21][23] ), .A(\_zyixc_ctx_rdata_29[21][23] ));
Q_ASSIGN U1785 ( .B(\mem_a[21][24] ), .A(\_zyixc_ctx_rdata_29[21][24] ));
Q_ASSIGN U1786 ( .B(\mem_a[21][25] ), .A(\_zyixc_ctx_rdata_29[21][25] ));
Q_ASSIGN U1787 ( .B(\mem_a[21][26] ), .A(\_zyixc_ctx_rdata_29[21][26] ));
Q_ASSIGN U1788 ( .B(\mem_a[21][27] ), .A(\_zyixc_ctx_rdata_29[21][27] ));
Q_ASSIGN U1789 ( .B(\mem_a[21][28] ), .A(\_zyixc_ctx_rdata_29[21][28] ));
Q_ASSIGN U1790 ( .B(\mem_a[21][29] ), .A(\_zyixc_ctx_rdata_29[21][29] ));
Q_ASSIGN U1791 ( .B(\mem_a[21][30] ), .A(\_zyixc_ctx_rdata_29[21][30] ));
Q_ASSIGN U1792 ( .B(\mem_a[21][31] ), .A(\_zyixc_ctx_rdata_29[21][31] ));
Q_ASSIGN U1793 ( .B(\mem_a[21][32] ), .A(\_zyixc_ctx_rdata_29[21][32] ));
Q_ASSIGN U1794 ( .B(\mem_a[21][33] ), .A(\_zyixc_ctx_rdata_29[21][33] ));
Q_ASSIGN U1795 ( .B(\mem_a[21][34] ), .A(\_zyixc_ctx_rdata_29[21][34] ));
Q_ASSIGN U1796 ( .B(\mem_a[21][35] ), .A(\_zyixc_ctx_rdata_29[21][35] ));
Q_ASSIGN U1797 ( .B(\mem_a[21][36] ), .A(\_zyixc_ctx_rdata_29[21][36] ));
Q_ASSIGN U1798 ( .B(\mem_a[21][37] ), .A(\_zyixc_ctx_rdata_29[21][37] ));
Q_ASSIGN U1799 ( .B(\mem_a[21][38] ), .A(\_zyixc_ctx_rdata_29[21][38] ));
Q_ASSIGN U1800 ( .B(\mem_a[21][39] ), .A(\_zyixc_ctx_rdata_29[21][39] ));
Q_ASSIGN U1801 ( .B(\mem_a[21][40] ), .A(\_zyixc_ctx_rdata_29[21][40] ));
Q_ASSIGN U1802 ( .B(\mem_a[21][41] ), .A(\_zyixc_ctx_rdata_29[21][41] ));
Q_ASSIGN U1803 ( .B(\mem_a[21][42] ), .A(\_zyixc_ctx_rdata_29[21][42] ));
Q_ASSIGN U1804 ( .B(\mem_a[21][43] ), .A(\_zyixc_ctx_rdata_29[21][43] ));
Q_ASSIGN U1805 ( .B(\mem_a[21][44] ), .A(\_zyixc_ctx_rdata_29[21][44] ));
Q_ASSIGN U1806 ( .B(\mem_a[21][45] ), .A(\_zyixc_ctx_rdata_29[21][45] ));
Q_ASSIGN U1807 ( .B(\mem_a[21][46] ), .A(\_zyixc_ctx_rdata_29[21][46] ));
Q_ASSIGN U1808 ( .B(\mem_a[21][47] ), .A(\_zyixc_ctx_rdata_29[21][47] ));
Q_ASSIGN U1809 ( .B(\mem_a[21][48] ), .A(\_zyixc_ctx_rdata_29[21][48] ));
Q_ASSIGN U1810 ( .B(\mem_a[21][49] ), .A(\_zyixc_ctx_rdata_29[21][49] ));
Q_ASSIGN U1811 ( .B(\mem_a[21][50] ), .A(\_zyixc_ctx_rdata_29[21][50] ));
Q_ASSIGN U1812 ( .B(\mem_a[21][51] ), .A(\_zyixc_ctx_rdata_29[21][51] ));
Q_ASSIGN U1813 ( .B(\mem_a[21][52] ), .A(\_zyixc_ctx_rdata_29[21][52] ));
Q_ASSIGN U1814 ( .B(\mem_a[21][53] ), .A(\_zyixc_ctx_rdata_29[21][53] ));
Q_ASSIGN U1815 ( .B(\mem_a[21][54] ), .A(\_zyixc_ctx_rdata_29[21][54] ));
Q_ASSIGN U1816 ( .B(\mem_a[21][55] ), .A(\_zyixc_ctx_rdata_29[21][55] ));
Q_ASSIGN U1817 ( .B(\mem_a[21][56] ), .A(\_zyixc_ctx_rdata_29[21][56] ));
Q_ASSIGN U1818 ( .B(\mem_a[21][57] ), .A(\_zyixc_ctx_rdata_29[21][57] ));
Q_ASSIGN U1819 ( .B(\mem_a[21][58] ), .A(\_zyixc_ctx_rdata_29[21][58] ));
Q_ASSIGN U1820 ( .B(\mem_a[21][59] ), .A(\_zyixc_ctx_rdata_29[21][59] ));
Q_ASSIGN U1821 ( .B(\mem_a[21][60] ), .A(\_zyixc_ctx_rdata_29[21][60] ));
Q_ASSIGN U1822 ( .B(\mem_a[21][61] ), .A(\_zyixc_ctx_rdata_29[21][61] ));
Q_ASSIGN U1823 ( .B(\mem_a[21][62] ), .A(\_zyixc_ctx_rdata_29[21][62] ));
Q_ASSIGN U1824 ( .B(\mem_a[21][63] ), .A(\_zyixc_ctx_rdata_29[21][63] ));
Q_ASSIGN U1825 ( .B(\mem_a[22][0] ), .A(\_zyixc_ctx_rdata_29[22][0] ));
Q_ASSIGN U1826 ( .B(\mem_a[22][1] ), .A(\_zyixc_ctx_rdata_29[22][1] ));
Q_ASSIGN U1827 ( .B(\mem_a[22][2] ), .A(\_zyixc_ctx_rdata_29[22][2] ));
Q_ASSIGN U1828 ( .B(\mem_a[22][3] ), .A(\_zyixc_ctx_rdata_29[22][3] ));
Q_ASSIGN U1829 ( .B(\mem_a[22][4] ), .A(\_zyixc_ctx_rdata_29[22][4] ));
Q_ASSIGN U1830 ( .B(\mem_a[22][5] ), .A(\_zyixc_ctx_rdata_29[22][5] ));
Q_ASSIGN U1831 ( .B(\mem_a[22][6] ), .A(\_zyixc_ctx_rdata_29[22][6] ));
Q_ASSIGN U1832 ( .B(\mem_a[22][7] ), .A(\_zyixc_ctx_rdata_29[22][7] ));
Q_ASSIGN U1833 ( .B(\mem_a[22][8] ), .A(\_zyixc_ctx_rdata_29[22][8] ));
Q_ASSIGN U1834 ( .B(\mem_a[22][9] ), .A(\_zyixc_ctx_rdata_29[22][9] ));
Q_ASSIGN U1835 ( .B(\mem_a[22][10] ), .A(\_zyixc_ctx_rdata_29[22][10] ));
Q_ASSIGN U1836 ( .B(\mem_a[22][11] ), .A(\_zyixc_ctx_rdata_29[22][11] ));
Q_ASSIGN U1837 ( .B(\mem_a[22][12] ), .A(\_zyixc_ctx_rdata_29[22][12] ));
Q_ASSIGN U1838 ( .B(\mem_a[22][13] ), .A(\_zyixc_ctx_rdata_29[22][13] ));
Q_ASSIGN U1839 ( .B(\mem_a[22][14] ), .A(\_zyixc_ctx_rdata_29[22][14] ));
Q_ASSIGN U1840 ( .B(\mem_a[22][15] ), .A(\_zyixc_ctx_rdata_29[22][15] ));
Q_ASSIGN U1841 ( .B(\mem_a[22][16] ), .A(\_zyixc_ctx_rdata_29[22][16] ));
Q_ASSIGN U1842 ( .B(\mem_a[22][17] ), .A(\_zyixc_ctx_rdata_29[22][17] ));
Q_ASSIGN U1843 ( .B(\mem_a[22][18] ), .A(\_zyixc_ctx_rdata_29[22][18] ));
Q_ASSIGN U1844 ( .B(\mem_a[22][19] ), .A(\_zyixc_ctx_rdata_29[22][19] ));
Q_ASSIGN U1845 ( .B(\mem_a[22][20] ), .A(\_zyixc_ctx_rdata_29[22][20] ));
Q_ASSIGN U1846 ( .B(\mem_a[22][21] ), .A(\_zyixc_ctx_rdata_29[22][21] ));
Q_ASSIGN U1847 ( .B(\mem_a[22][22] ), .A(\_zyixc_ctx_rdata_29[22][22] ));
Q_ASSIGN U1848 ( .B(\mem_a[22][23] ), .A(\_zyixc_ctx_rdata_29[22][23] ));
Q_ASSIGN U1849 ( .B(\mem_a[22][24] ), .A(\_zyixc_ctx_rdata_29[22][24] ));
Q_ASSIGN U1850 ( .B(\mem_a[22][25] ), .A(\_zyixc_ctx_rdata_29[22][25] ));
Q_ASSIGN U1851 ( .B(\mem_a[22][26] ), .A(\_zyixc_ctx_rdata_29[22][26] ));
Q_ASSIGN U1852 ( .B(\mem_a[22][27] ), .A(\_zyixc_ctx_rdata_29[22][27] ));
Q_ASSIGN U1853 ( .B(\mem_a[22][28] ), .A(\_zyixc_ctx_rdata_29[22][28] ));
Q_ASSIGN U1854 ( .B(\mem_a[22][29] ), .A(\_zyixc_ctx_rdata_29[22][29] ));
Q_ASSIGN U1855 ( .B(\mem_a[22][30] ), .A(\_zyixc_ctx_rdata_29[22][30] ));
Q_ASSIGN U1856 ( .B(\mem_a[22][31] ), .A(\_zyixc_ctx_rdata_29[22][31] ));
Q_ASSIGN U1857 ( .B(\mem_a[22][32] ), .A(\_zyixc_ctx_rdata_29[22][32] ));
Q_ASSIGN U1858 ( .B(\mem_a[22][33] ), .A(\_zyixc_ctx_rdata_29[22][33] ));
Q_ASSIGN U1859 ( .B(\mem_a[22][34] ), .A(\_zyixc_ctx_rdata_29[22][34] ));
Q_ASSIGN U1860 ( .B(\mem_a[22][35] ), .A(\_zyixc_ctx_rdata_29[22][35] ));
Q_ASSIGN U1861 ( .B(\mem_a[22][36] ), .A(\_zyixc_ctx_rdata_29[22][36] ));
Q_ASSIGN U1862 ( .B(\mem_a[22][37] ), .A(\_zyixc_ctx_rdata_29[22][37] ));
Q_ASSIGN U1863 ( .B(\mem_a[22][38] ), .A(\_zyixc_ctx_rdata_29[22][38] ));
Q_ASSIGN U1864 ( .B(\mem_a[22][39] ), .A(\_zyixc_ctx_rdata_29[22][39] ));
Q_ASSIGN U1865 ( .B(\mem_a[22][40] ), .A(\_zyixc_ctx_rdata_29[22][40] ));
Q_ASSIGN U1866 ( .B(\mem_a[22][41] ), .A(\_zyixc_ctx_rdata_29[22][41] ));
Q_ASSIGN U1867 ( .B(\mem_a[22][42] ), .A(\_zyixc_ctx_rdata_29[22][42] ));
Q_ASSIGN U1868 ( .B(\mem_a[22][43] ), .A(\_zyixc_ctx_rdata_29[22][43] ));
Q_ASSIGN U1869 ( .B(\mem_a[22][44] ), .A(\_zyixc_ctx_rdata_29[22][44] ));
Q_ASSIGN U1870 ( .B(\mem_a[22][45] ), .A(\_zyixc_ctx_rdata_29[22][45] ));
Q_ASSIGN U1871 ( .B(\mem_a[22][46] ), .A(\_zyixc_ctx_rdata_29[22][46] ));
Q_ASSIGN U1872 ( .B(\mem_a[22][47] ), .A(\_zyixc_ctx_rdata_29[22][47] ));
Q_ASSIGN U1873 ( .B(\mem_a[22][48] ), .A(\_zyixc_ctx_rdata_29[22][48] ));
Q_ASSIGN U1874 ( .B(\mem_a[22][49] ), .A(\_zyixc_ctx_rdata_29[22][49] ));
Q_ASSIGN U1875 ( .B(\mem_a[22][50] ), .A(\_zyixc_ctx_rdata_29[22][50] ));
Q_ASSIGN U1876 ( .B(\mem_a[22][51] ), .A(\_zyixc_ctx_rdata_29[22][51] ));
Q_ASSIGN U1877 ( .B(\mem_a[22][52] ), .A(\_zyixc_ctx_rdata_29[22][52] ));
Q_ASSIGN U1878 ( .B(\mem_a[22][53] ), .A(\_zyixc_ctx_rdata_29[22][53] ));
Q_ASSIGN U1879 ( .B(\mem_a[22][54] ), .A(\_zyixc_ctx_rdata_29[22][54] ));
Q_ASSIGN U1880 ( .B(\mem_a[22][55] ), .A(\_zyixc_ctx_rdata_29[22][55] ));
Q_ASSIGN U1881 ( .B(\mem_a[22][56] ), .A(\_zyixc_ctx_rdata_29[22][56] ));
Q_ASSIGN U1882 ( .B(\mem_a[22][57] ), .A(\_zyixc_ctx_rdata_29[22][57] ));
Q_ASSIGN U1883 ( .B(\mem_a[22][58] ), .A(\_zyixc_ctx_rdata_29[22][58] ));
Q_ASSIGN U1884 ( .B(\mem_a[22][59] ), .A(\_zyixc_ctx_rdata_29[22][59] ));
Q_ASSIGN U1885 ( .B(\mem_a[22][60] ), .A(\_zyixc_ctx_rdata_29[22][60] ));
Q_ASSIGN U1886 ( .B(\mem_a[22][61] ), .A(\_zyixc_ctx_rdata_29[22][61] ));
Q_ASSIGN U1887 ( .B(\mem_a[22][62] ), .A(\_zyixc_ctx_rdata_29[22][62] ));
Q_ASSIGN U1888 ( .B(\mem_a[22][63] ), .A(\_zyixc_ctx_rdata_29[22][63] ));
Q_ASSIGN U1889 ( .B(\mem_a[23][0] ), .A(\_zyixc_ctx_rdata_29[23][0] ));
Q_ASSIGN U1890 ( .B(\mem_a[23][1] ), .A(\_zyixc_ctx_rdata_29[23][1] ));
Q_ASSIGN U1891 ( .B(\mem_a[23][2] ), .A(\_zyixc_ctx_rdata_29[23][2] ));
Q_ASSIGN U1892 ( .B(\mem_a[23][3] ), .A(\_zyixc_ctx_rdata_29[23][3] ));
Q_ASSIGN U1893 ( .B(\mem_a[23][4] ), .A(\_zyixc_ctx_rdata_29[23][4] ));
Q_ASSIGN U1894 ( .B(\mem_a[23][5] ), .A(\_zyixc_ctx_rdata_29[23][5] ));
Q_ASSIGN U1895 ( .B(\mem_a[23][6] ), .A(\_zyixc_ctx_rdata_29[23][6] ));
Q_ASSIGN U1896 ( .B(\mem_a[23][7] ), .A(\_zyixc_ctx_rdata_29[23][7] ));
Q_ASSIGN U1897 ( .B(\mem_a[23][8] ), .A(\_zyixc_ctx_rdata_29[23][8] ));
Q_ASSIGN U1898 ( .B(\mem_a[23][9] ), .A(\_zyixc_ctx_rdata_29[23][9] ));
Q_ASSIGN U1899 ( .B(\mem_a[23][10] ), .A(\_zyixc_ctx_rdata_29[23][10] ));
Q_ASSIGN U1900 ( .B(\mem_a[23][11] ), .A(\_zyixc_ctx_rdata_29[23][11] ));
Q_ASSIGN U1901 ( .B(\mem_a[23][12] ), .A(\_zyixc_ctx_rdata_29[23][12] ));
Q_ASSIGN U1902 ( .B(\mem_a[23][13] ), .A(\_zyixc_ctx_rdata_29[23][13] ));
Q_ASSIGN U1903 ( .B(\mem_a[23][14] ), .A(\_zyixc_ctx_rdata_29[23][14] ));
Q_ASSIGN U1904 ( .B(\mem_a[23][15] ), .A(\_zyixc_ctx_rdata_29[23][15] ));
Q_ASSIGN U1905 ( .B(\mem_a[23][16] ), .A(\_zyixc_ctx_rdata_29[23][16] ));
Q_ASSIGN U1906 ( .B(\mem_a[23][17] ), .A(\_zyixc_ctx_rdata_29[23][17] ));
Q_ASSIGN U1907 ( .B(\mem_a[23][18] ), .A(\_zyixc_ctx_rdata_29[23][18] ));
Q_ASSIGN U1908 ( .B(\mem_a[23][19] ), .A(\_zyixc_ctx_rdata_29[23][19] ));
Q_ASSIGN U1909 ( .B(\mem_a[23][20] ), .A(\_zyixc_ctx_rdata_29[23][20] ));
Q_ASSIGN U1910 ( .B(\mem_a[23][21] ), .A(\_zyixc_ctx_rdata_29[23][21] ));
Q_ASSIGN U1911 ( .B(\mem_a[23][22] ), .A(\_zyixc_ctx_rdata_29[23][22] ));
Q_ASSIGN U1912 ( .B(\mem_a[23][23] ), .A(\_zyixc_ctx_rdata_29[23][23] ));
Q_ASSIGN U1913 ( .B(\mem_a[23][24] ), .A(\_zyixc_ctx_rdata_29[23][24] ));
Q_ASSIGN U1914 ( .B(\mem_a[23][25] ), .A(\_zyixc_ctx_rdata_29[23][25] ));
Q_ASSIGN U1915 ( .B(\mem_a[23][26] ), .A(\_zyixc_ctx_rdata_29[23][26] ));
Q_ASSIGN U1916 ( .B(\mem_a[23][27] ), .A(\_zyixc_ctx_rdata_29[23][27] ));
Q_ASSIGN U1917 ( .B(\mem_a[23][28] ), .A(\_zyixc_ctx_rdata_29[23][28] ));
Q_ASSIGN U1918 ( .B(\mem_a[23][29] ), .A(\_zyixc_ctx_rdata_29[23][29] ));
Q_ASSIGN U1919 ( .B(\mem_a[23][30] ), .A(\_zyixc_ctx_rdata_29[23][30] ));
Q_ASSIGN U1920 ( .B(\mem_a[23][31] ), .A(\_zyixc_ctx_rdata_29[23][31] ));
Q_ASSIGN U1921 ( .B(\mem_a[23][32] ), .A(\_zyixc_ctx_rdata_29[23][32] ));
Q_ASSIGN U1922 ( .B(\mem_a[23][33] ), .A(\_zyixc_ctx_rdata_29[23][33] ));
Q_ASSIGN U1923 ( .B(\mem_a[23][34] ), .A(\_zyixc_ctx_rdata_29[23][34] ));
Q_ASSIGN U1924 ( .B(\mem_a[23][35] ), .A(\_zyixc_ctx_rdata_29[23][35] ));
Q_ASSIGN U1925 ( .B(\mem_a[23][36] ), .A(\_zyixc_ctx_rdata_29[23][36] ));
Q_ASSIGN U1926 ( .B(\mem_a[23][37] ), .A(\_zyixc_ctx_rdata_29[23][37] ));
Q_ASSIGN U1927 ( .B(\mem_a[23][38] ), .A(\_zyixc_ctx_rdata_29[23][38] ));
Q_ASSIGN U1928 ( .B(\mem_a[23][39] ), .A(\_zyixc_ctx_rdata_29[23][39] ));
Q_ASSIGN U1929 ( .B(\mem_a[23][40] ), .A(\_zyixc_ctx_rdata_29[23][40] ));
Q_ASSIGN U1930 ( .B(\mem_a[23][41] ), .A(\_zyixc_ctx_rdata_29[23][41] ));
Q_ASSIGN U1931 ( .B(\mem_a[23][42] ), .A(\_zyixc_ctx_rdata_29[23][42] ));
Q_ASSIGN U1932 ( .B(\mem_a[23][43] ), .A(\_zyixc_ctx_rdata_29[23][43] ));
Q_ASSIGN U1933 ( .B(\mem_a[23][44] ), .A(\_zyixc_ctx_rdata_29[23][44] ));
Q_ASSIGN U1934 ( .B(\mem_a[23][45] ), .A(\_zyixc_ctx_rdata_29[23][45] ));
Q_ASSIGN U1935 ( .B(\mem_a[23][46] ), .A(\_zyixc_ctx_rdata_29[23][46] ));
Q_ASSIGN U1936 ( .B(\mem_a[23][47] ), .A(\_zyixc_ctx_rdata_29[23][47] ));
Q_ASSIGN U1937 ( .B(\mem_a[23][48] ), .A(\_zyixc_ctx_rdata_29[23][48] ));
Q_ASSIGN U1938 ( .B(\mem_a[23][49] ), .A(\_zyixc_ctx_rdata_29[23][49] ));
Q_ASSIGN U1939 ( .B(\mem_a[23][50] ), .A(\_zyixc_ctx_rdata_29[23][50] ));
Q_ASSIGN U1940 ( .B(\mem_a[23][51] ), .A(\_zyixc_ctx_rdata_29[23][51] ));
Q_ASSIGN U1941 ( .B(\mem_a[23][52] ), .A(\_zyixc_ctx_rdata_29[23][52] ));
Q_ASSIGN U1942 ( .B(\mem_a[23][53] ), .A(\_zyixc_ctx_rdata_29[23][53] ));
Q_ASSIGN U1943 ( .B(\mem_a[23][54] ), .A(\_zyixc_ctx_rdata_29[23][54] ));
Q_ASSIGN U1944 ( .B(\mem_a[23][55] ), .A(\_zyixc_ctx_rdata_29[23][55] ));
Q_ASSIGN U1945 ( .B(\mem_a[23][56] ), .A(\_zyixc_ctx_rdata_29[23][56] ));
Q_ASSIGN U1946 ( .B(\mem_a[23][57] ), .A(\_zyixc_ctx_rdata_29[23][57] ));
Q_ASSIGN U1947 ( .B(\mem_a[23][58] ), .A(\_zyixc_ctx_rdata_29[23][58] ));
Q_ASSIGN U1948 ( .B(\mem_a[23][59] ), .A(\_zyixc_ctx_rdata_29[23][59] ));
Q_ASSIGN U1949 ( .B(\mem_a[23][60] ), .A(\_zyixc_ctx_rdata_29[23][60] ));
Q_ASSIGN U1950 ( .B(\mem_a[23][61] ), .A(\_zyixc_ctx_rdata_29[23][61] ));
Q_ASSIGN U1951 ( .B(\mem_a[23][62] ), .A(\_zyixc_ctx_rdata_29[23][62] ));
Q_ASSIGN U1952 ( .B(\mem_a[23][63] ), .A(\_zyixc_ctx_rdata_29[23][63] ));
Q_ASSIGN U1953 ( .B(\mem_a[24][0] ), .A(\_zyixc_ctx_rdata_29[24][0] ));
Q_ASSIGN U1954 ( .B(\mem_a[24][1] ), .A(\_zyixc_ctx_rdata_29[24][1] ));
Q_ASSIGN U1955 ( .B(\mem_a[24][2] ), .A(\_zyixc_ctx_rdata_29[24][2] ));
Q_ASSIGN U1956 ( .B(\mem_a[24][3] ), .A(\_zyixc_ctx_rdata_29[24][3] ));
Q_ASSIGN U1957 ( .B(\mem_a[24][4] ), .A(\_zyixc_ctx_rdata_29[24][4] ));
Q_ASSIGN U1958 ( .B(\mem_a[24][5] ), .A(\_zyixc_ctx_rdata_29[24][5] ));
Q_ASSIGN U1959 ( .B(\mem_a[24][6] ), .A(\_zyixc_ctx_rdata_29[24][6] ));
Q_ASSIGN U1960 ( .B(\mem_a[24][7] ), .A(\_zyixc_ctx_rdata_29[24][7] ));
Q_ASSIGN U1961 ( .B(\mem_a[24][8] ), .A(\_zyixc_ctx_rdata_29[24][8] ));
Q_ASSIGN U1962 ( .B(\mem_a[24][9] ), .A(\_zyixc_ctx_rdata_29[24][9] ));
Q_ASSIGN U1963 ( .B(\mem_a[24][10] ), .A(\_zyixc_ctx_rdata_29[24][10] ));
Q_ASSIGN U1964 ( .B(\mem_a[24][11] ), .A(\_zyixc_ctx_rdata_29[24][11] ));
Q_ASSIGN U1965 ( .B(\mem_a[24][12] ), .A(\_zyixc_ctx_rdata_29[24][12] ));
Q_ASSIGN U1966 ( .B(\mem_a[24][13] ), .A(\_zyixc_ctx_rdata_29[24][13] ));
Q_ASSIGN U1967 ( .B(\mem_a[24][14] ), .A(\_zyixc_ctx_rdata_29[24][14] ));
Q_ASSIGN U1968 ( .B(\mem_a[24][15] ), .A(\_zyixc_ctx_rdata_29[24][15] ));
Q_ASSIGN U1969 ( .B(\mem_a[24][16] ), .A(\_zyixc_ctx_rdata_29[24][16] ));
Q_ASSIGN U1970 ( .B(\mem_a[24][17] ), .A(\_zyixc_ctx_rdata_29[24][17] ));
Q_ASSIGN U1971 ( .B(\mem_a[24][18] ), .A(\_zyixc_ctx_rdata_29[24][18] ));
Q_ASSIGN U1972 ( .B(\mem_a[24][19] ), .A(\_zyixc_ctx_rdata_29[24][19] ));
Q_ASSIGN U1973 ( .B(\mem_a[24][20] ), .A(\_zyixc_ctx_rdata_29[24][20] ));
Q_ASSIGN U1974 ( .B(\mem_a[24][21] ), .A(\_zyixc_ctx_rdata_29[24][21] ));
Q_ASSIGN U1975 ( .B(\mem_a[24][22] ), .A(\_zyixc_ctx_rdata_29[24][22] ));
Q_ASSIGN U1976 ( .B(\mem_a[24][23] ), .A(\_zyixc_ctx_rdata_29[24][23] ));
Q_ASSIGN U1977 ( .B(\mem_a[24][24] ), .A(\_zyixc_ctx_rdata_29[24][24] ));
Q_ASSIGN U1978 ( .B(\mem_a[24][25] ), .A(\_zyixc_ctx_rdata_29[24][25] ));
Q_ASSIGN U1979 ( .B(\mem_a[24][26] ), .A(\_zyixc_ctx_rdata_29[24][26] ));
Q_ASSIGN U1980 ( .B(\mem_a[24][27] ), .A(\_zyixc_ctx_rdata_29[24][27] ));
Q_ASSIGN U1981 ( .B(\mem_a[24][28] ), .A(\_zyixc_ctx_rdata_29[24][28] ));
Q_ASSIGN U1982 ( .B(\mem_a[24][29] ), .A(\_zyixc_ctx_rdata_29[24][29] ));
Q_ASSIGN U1983 ( .B(\mem_a[24][30] ), .A(\_zyixc_ctx_rdata_29[24][30] ));
Q_ASSIGN U1984 ( .B(\mem_a[24][31] ), .A(\_zyixc_ctx_rdata_29[24][31] ));
Q_ASSIGN U1985 ( .B(\mem_a[24][32] ), .A(\_zyixc_ctx_rdata_29[24][32] ));
Q_ASSIGN U1986 ( .B(\mem_a[24][33] ), .A(\_zyixc_ctx_rdata_29[24][33] ));
Q_ASSIGN U1987 ( .B(\mem_a[24][34] ), .A(\_zyixc_ctx_rdata_29[24][34] ));
Q_ASSIGN U1988 ( .B(\mem_a[24][35] ), .A(\_zyixc_ctx_rdata_29[24][35] ));
Q_ASSIGN U1989 ( .B(\mem_a[24][36] ), .A(\_zyixc_ctx_rdata_29[24][36] ));
Q_ASSIGN U1990 ( .B(\mem_a[24][37] ), .A(\_zyixc_ctx_rdata_29[24][37] ));
Q_ASSIGN U1991 ( .B(\mem_a[24][38] ), .A(\_zyixc_ctx_rdata_29[24][38] ));
Q_ASSIGN U1992 ( .B(\mem_a[24][39] ), .A(\_zyixc_ctx_rdata_29[24][39] ));
Q_ASSIGN U1993 ( .B(\mem_a[24][40] ), .A(\_zyixc_ctx_rdata_29[24][40] ));
Q_ASSIGN U1994 ( .B(\mem_a[24][41] ), .A(\_zyixc_ctx_rdata_29[24][41] ));
Q_ASSIGN U1995 ( .B(\mem_a[24][42] ), .A(\_zyixc_ctx_rdata_29[24][42] ));
Q_ASSIGN U1996 ( .B(\mem_a[24][43] ), .A(\_zyixc_ctx_rdata_29[24][43] ));
Q_ASSIGN U1997 ( .B(\mem_a[24][44] ), .A(\_zyixc_ctx_rdata_29[24][44] ));
Q_ASSIGN U1998 ( .B(\mem_a[24][45] ), .A(\_zyixc_ctx_rdata_29[24][45] ));
Q_ASSIGN U1999 ( .B(\mem_a[24][46] ), .A(\_zyixc_ctx_rdata_29[24][46] ));
Q_ASSIGN U2000 ( .B(\mem_a[24][47] ), .A(\_zyixc_ctx_rdata_29[24][47] ));
Q_ASSIGN U2001 ( .B(\mem_a[24][48] ), .A(\_zyixc_ctx_rdata_29[24][48] ));
Q_ASSIGN U2002 ( .B(\mem_a[24][49] ), .A(\_zyixc_ctx_rdata_29[24][49] ));
Q_ASSIGN U2003 ( .B(\mem_a[24][50] ), .A(\_zyixc_ctx_rdata_29[24][50] ));
Q_ASSIGN U2004 ( .B(\mem_a[24][51] ), .A(\_zyixc_ctx_rdata_29[24][51] ));
Q_ASSIGN U2005 ( .B(\mem_a[24][52] ), .A(\_zyixc_ctx_rdata_29[24][52] ));
Q_ASSIGN U2006 ( .B(\mem_a[24][53] ), .A(\_zyixc_ctx_rdata_29[24][53] ));
Q_ASSIGN U2007 ( .B(\mem_a[24][54] ), .A(\_zyixc_ctx_rdata_29[24][54] ));
Q_ASSIGN U2008 ( .B(\mem_a[24][55] ), .A(\_zyixc_ctx_rdata_29[24][55] ));
Q_ASSIGN U2009 ( .B(\mem_a[24][56] ), .A(\_zyixc_ctx_rdata_29[24][56] ));
Q_ASSIGN U2010 ( .B(\mem_a[24][57] ), .A(\_zyixc_ctx_rdata_29[24][57] ));
Q_ASSIGN U2011 ( .B(\mem_a[24][58] ), .A(\_zyixc_ctx_rdata_29[24][58] ));
Q_ASSIGN U2012 ( .B(\mem_a[24][59] ), .A(\_zyixc_ctx_rdata_29[24][59] ));
Q_ASSIGN U2013 ( .B(\mem_a[24][60] ), .A(\_zyixc_ctx_rdata_29[24][60] ));
Q_ASSIGN U2014 ( .B(\mem_a[24][61] ), .A(\_zyixc_ctx_rdata_29[24][61] ));
Q_ASSIGN U2015 ( .B(\mem_a[24][62] ), .A(\_zyixc_ctx_rdata_29[24][62] ));
Q_ASSIGN U2016 ( .B(\mem_a[24][63] ), .A(\_zyixc_ctx_rdata_29[24][63] ));
Q_ASSIGN U2017 ( .B(\mem_a[25][0] ), .A(\_zyixc_ctx_rdata_29[25][0] ));
Q_ASSIGN U2018 ( .B(\mem_a[25][1] ), .A(\_zyixc_ctx_rdata_29[25][1] ));
Q_ASSIGN U2019 ( .B(\mem_a[25][2] ), .A(\_zyixc_ctx_rdata_29[25][2] ));
Q_ASSIGN U2020 ( .B(\mem_a[25][3] ), .A(\_zyixc_ctx_rdata_29[25][3] ));
Q_ASSIGN U2021 ( .B(\mem_a[25][4] ), .A(\_zyixc_ctx_rdata_29[25][4] ));
Q_ASSIGN U2022 ( .B(\mem_a[25][5] ), .A(\_zyixc_ctx_rdata_29[25][5] ));
Q_ASSIGN U2023 ( .B(\mem_a[25][6] ), .A(\_zyixc_ctx_rdata_29[25][6] ));
Q_ASSIGN U2024 ( .B(\mem_a[25][7] ), .A(\_zyixc_ctx_rdata_29[25][7] ));
Q_ASSIGN U2025 ( .B(\mem_a[25][8] ), .A(\_zyixc_ctx_rdata_29[25][8] ));
Q_ASSIGN U2026 ( .B(\mem_a[25][9] ), .A(\_zyixc_ctx_rdata_29[25][9] ));
Q_ASSIGN U2027 ( .B(\mem_a[25][10] ), .A(\_zyixc_ctx_rdata_29[25][10] ));
Q_ASSIGN U2028 ( .B(\mem_a[25][11] ), .A(\_zyixc_ctx_rdata_29[25][11] ));
Q_ASSIGN U2029 ( .B(\mem_a[25][12] ), .A(\_zyixc_ctx_rdata_29[25][12] ));
Q_ASSIGN U2030 ( .B(\mem_a[25][13] ), .A(\_zyixc_ctx_rdata_29[25][13] ));
Q_ASSIGN U2031 ( .B(\mem_a[25][14] ), .A(\_zyixc_ctx_rdata_29[25][14] ));
Q_ASSIGN U2032 ( .B(\mem_a[25][15] ), .A(\_zyixc_ctx_rdata_29[25][15] ));
Q_ASSIGN U2033 ( .B(\mem_a[25][16] ), .A(\_zyixc_ctx_rdata_29[25][16] ));
Q_ASSIGN U2034 ( .B(\mem_a[25][17] ), .A(\_zyixc_ctx_rdata_29[25][17] ));
Q_ASSIGN U2035 ( .B(\mem_a[25][18] ), .A(\_zyixc_ctx_rdata_29[25][18] ));
Q_ASSIGN U2036 ( .B(\mem_a[25][19] ), .A(\_zyixc_ctx_rdata_29[25][19] ));
Q_ASSIGN U2037 ( .B(\mem_a[25][20] ), .A(\_zyixc_ctx_rdata_29[25][20] ));
Q_ASSIGN U2038 ( .B(\mem_a[25][21] ), .A(\_zyixc_ctx_rdata_29[25][21] ));
Q_ASSIGN U2039 ( .B(\mem_a[25][22] ), .A(\_zyixc_ctx_rdata_29[25][22] ));
Q_ASSIGN U2040 ( .B(\mem_a[25][23] ), .A(\_zyixc_ctx_rdata_29[25][23] ));
Q_ASSIGN U2041 ( .B(\mem_a[25][24] ), .A(\_zyixc_ctx_rdata_29[25][24] ));
Q_ASSIGN U2042 ( .B(\mem_a[25][25] ), .A(\_zyixc_ctx_rdata_29[25][25] ));
Q_ASSIGN U2043 ( .B(\mem_a[25][26] ), .A(\_zyixc_ctx_rdata_29[25][26] ));
Q_ASSIGN U2044 ( .B(\mem_a[25][27] ), .A(\_zyixc_ctx_rdata_29[25][27] ));
Q_ASSIGN U2045 ( .B(\mem_a[25][28] ), .A(\_zyixc_ctx_rdata_29[25][28] ));
Q_ASSIGN U2046 ( .B(\mem_a[25][29] ), .A(\_zyixc_ctx_rdata_29[25][29] ));
Q_ASSIGN U2047 ( .B(\mem_a[25][30] ), .A(\_zyixc_ctx_rdata_29[25][30] ));
Q_ASSIGN U2048 ( .B(\mem_a[25][31] ), .A(\_zyixc_ctx_rdata_29[25][31] ));
Q_ASSIGN U2049 ( .B(\mem_a[25][32] ), .A(\_zyixc_ctx_rdata_29[25][32] ));
Q_ASSIGN U2050 ( .B(\mem_a[25][33] ), .A(\_zyixc_ctx_rdata_29[25][33] ));
Q_ASSIGN U2051 ( .B(\mem_a[25][34] ), .A(\_zyixc_ctx_rdata_29[25][34] ));
Q_ASSIGN U2052 ( .B(\mem_a[25][35] ), .A(\_zyixc_ctx_rdata_29[25][35] ));
Q_ASSIGN U2053 ( .B(\mem_a[25][36] ), .A(\_zyixc_ctx_rdata_29[25][36] ));
Q_ASSIGN U2054 ( .B(\mem_a[25][37] ), .A(\_zyixc_ctx_rdata_29[25][37] ));
Q_ASSIGN U2055 ( .B(\mem_a[25][38] ), .A(\_zyixc_ctx_rdata_29[25][38] ));
Q_ASSIGN U2056 ( .B(\mem_a[25][39] ), .A(\_zyixc_ctx_rdata_29[25][39] ));
Q_ASSIGN U2057 ( .B(\mem_a[25][40] ), .A(\_zyixc_ctx_rdata_29[25][40] ));
Q_ASSIGN U2058 ( .B(\mem_a[25][41] ), .A(\_zyixc_ctx_rdata_29[25][41] ));
Q_ASSIGN U2059 ( .B(\mem_a[25][42] ), .A(\_zyixc_ctx_rdata_29[25][42] ));
Q_ASSIGN U2060 ( .B(\mem_a[25][43] ), .A(\_zyixc_ctx_rdata_29[25][43] ));
Q_ASSIGN U2061 ( .B(\mem_a[25][44] ), .A(\_zyixc_ctx_rdata_29[25][44] ));
Q_ASSIGN U2062 ( .B(\mem_a[25][45] ), .A(\_zyixc_ctx_rdata_29[25][45] ));
Q_ASSIGN U2063 ( .B(\mem_a[25][46] ), .A(\_zyixc_ctx_rdata_29[25][46] ));
Q_ASSIGN U2064 ( .B(\mem_a[25][47] ), .A(\_zyixc_ctx_rdata_29[25][47] ));
Q_ASSIGN U2065 ( .B(\mem_a[25][48] ), .A(\_zyixc_ctx_rdata_29[25][48] ));
Q_ASSIGN U2066 ( .B(\mem_a[25][49] ), .A(\_zyixc_ctx_rdata_29[25][49] ));
Q_ASSIGN U2067 ( .B(\mem_a[25][50] ), .A(\_zyixc_ctx_rdata_29[25][50] ));
Q_ASSIGN U2068 ( .B(\mem_a[25][51] ), .A(\_zyixc_ctx_rdata_29[25][51] ));
Q_ASSIGN U2069 ( .B(\mem_a[25][52] ), .A(\_zyixc_ctx_rdata_29[25][52] ));
Q_ASSIGN U2070 ( .B(\mem_a[25][53] ), .A(\_zyixc_ctx_rdata_29[25][53] ));
Q_ASSIGN U2071 ( .B(\mem_a[25][54] ), .A(\_zyixc_ctx_rdata_29[25][54] ));
Q_ASSIGN U2072 ( .B(\mem_a[25][55] ), .A(\_zyixc_ctx_rdata_29[25][55] ));
Q_ASSIGN U2073 ( .B(\mem_a[25][56] ), .A(\_zyixc_ctx_rdata_29[25][56] ));
Q_ASSIGN U2074 ( .B(\mem_a[25][57] ), .A(\_zyixc_ctx_rdata_29[25][57] ));
Q_ASSIGN U2075 ( .B(\mem_a[25][58] ), .A(\_zyixc_ctx_rdata_29[25][58] ));
Q_ASSIGN U2076 ( .B(\mem_a[25][59] ), .A(\_zyixc_ctx_rdata_29[25][59] ));
Q_ASSIGN U2077 ( .B(\mem_a[25][60] ), .A(\_zyixc_ctx_rdata_29[25][60] ));
Q_ASSIGN U2078 ( .B(\mem_a[25][61] ), .A(\_zyixc_ctx_rdata_29[25][61] ));
Q_ASSIGN U2079 ( .B(\mem_a[25][62] ), .A(\_zyixc_ctx_rdata_29[25][62] ));
Q_ASSIGN U2080 ( .B(\mem_a[25][63] ), .A(\_zyixc_ctx_rdata_29[25][63] ));
Q_ASSIGN U2081 ( .B(\mem_a[26][0] ), .A(\_zyixc_ctx_rdata_29[26][0] ));
Q_ASSIGN U2082 ( .B(\mem_a[26][1] ), .A(\_zyixc_ctx_rdata_29[26][1] ));
Q_ASSIGN U2083 ( .B(\mem_a[26][2] ), .A(\_zyixc_ctx_rdata_29[26][2] ));
Q_ASSIGN U2084 ( .B(\mem_a[26][3] ), .A(\_zyixc_ctx_rdata_29[26][3] ));
Q_ASSIGN U2085 ( .B(\mem_a[26][4] ), .A(\_zyixc_ctx_rdata_29[26][4] ));
Q_ASSIGN U2086 ( .B(\mem_a[26][5] ), .A(\_zyixc_ctx_rdata_29[26][5] ));
Q_ASSIGN U2087 ( .B(\mem_a[26][6] ), .A(\_zyixc_ctx_rdata_29[26][6] ));
Q_ASSIGN U2088 ( .B(\mem_a[26][7] ), .A(\_zyixc_ctx_rdata_29[26][7] ));
Q_ASSIGN U2089 ( .B(\mem_a[26][8] ), .A(\_zyixc_ctx_rdata_29[26][8] ));
Q_ASSIGN U2090 ( .B(\mem_a[26][9] ), .A(\_zyixc_ctx_rdata_29[26][9] ));
Q_ASSIGN U2091 ( .B(\mem_a[26][10] ), .A(\_zyixc_ctx_rdata_29[26][10] ));
Q_ASSIGN U2092 ( .B(\mem_a[26][11] ), .A(\_zyixc_ctx_rdata_29[26][11] ));
Q_ASSIGN U2093 ( .B(\mem_a[26][12] ), .A(\_zyixc_ctx_rdata_29[26][12] ));
Q_ASSIGN U2094 ( .B(\mem_a[26][13] ), .A(\_zyixc_ctx_rdata_29[26][13] ));
Q_ASSIGN U2095 ( .B(\mem_a[26][14] ), .A(\_zyixc_ctx_rdata_29[26][14] ));
Q_ASSIGN U2096 ( .B(\mem_a[26][15] ), .A(\_zyixc_ctx_rdata_29[26][15] ));
Q_ASSIGN U2097 ( .B(\mem_a[26][16] ), .A(\_zyixc_ctx_rdata_29[26][16] ));
Q_ASSIGN U2098 ( .B(\mem_a[26][17] ), .A(\_zyixc_ctx_rdata_29[26][17] ));
Q_ASSIGN U2099 ( .B(\mem_a[26][18] ), .A(\_zyixc_ctx_rdata_29[26][18] ));
Q_ASSIGN U2100 ( .B(\mem_a[26][19] ), .A(\_zyixc_ctx_rdata_29[26][19] ));
Q_ASSIGN U2101 ( .B(\mem_a[26][20] ), .A(\_zyixc_ctx_rdata_29[26][20] ));
Q_ASSIGN U2102 ( .B(\mem_a[26][21] ), .A(\_zyixc_ctx_rdata_29[26][21] ));
Q_ASSIGN U2103 ( .B(\mem_a[26][22] ), .A(\_zyixc_ctx_rdata_29[26][22] ));
Q_ASSIGN U2104 ( .B(\mem_a[26][23] ), .A(\_zyixc_ctx_rdata_29[26][23] ));
Q_ASSIGN U2105 ( .B(\mem_a[26][24] ), .A(\_zyixc_ctx_rdata_29[26][24] ));
Q_ASSIGN U2106 ( .B(\mem_a[26][25] ), .A(\_zyixc_ctx_rdata_29[26][25] ));
Q_ASSIGN U2107 ( .B(\mem_a[26][26] ), .A(\_zyixc_ctx_rdata_29[26][26] ));
Q_ASSIGN U2108 ( .B(\mem_a[26][27] ), .A(\_zyixc_ctx_rdata_29[26][27] ));
Q_ASSIGN U2109 ( .B(\mem_a[26][28] ), .A(\_zyixc_ctx_rdata_29[26][28] ));
Q_ASSIGN U2110 ( .B(\mem_a[26][29] ), .A(\_zyixc_ctx_rdata_29[26][29] ));
Q_ASSIGN U2111 ( .B(\mem_a[26][30] ), .A(\_zyixc_ctx_rdata_29[26][30] ));
Q_ASSIGN U2112 ( .B(\mem_a[26][31] ), .A(\_zyixc_ctx_rdata_29[26][31] ));
Q_ASSIGN U2113 ( .B(\mem_a[26][32] ), .A(\_zyixc_ctx_rdata_29[26][32] ));
Q_ASSIGN U2114 ( .B(\mem_a[26][33] ), .A(\_zyixc_ctx_rdata_29[26][33] ));
Q_ASSIGN U2115 ( .B(\mem_a[26][34] ), .A(\_zyixc_ctx_rdata_29[26][34] ));
Q_ASSIGN U2116 ( .B(\mem_a[26][35] ), .A(\_zyixc_ctx_rdata_29[26][35] ));
Q_ASSIGN U2117 ( .B(\mem_a[26][36] ), .A(\_zyixc_ctx_rdata_29[26][36] ));
Q_ASSIGN U2118 ( .B(\mem_a[26][37] ), .A(\_zyixc_ctx_rdata_29[26][37] ));
Q_ASSIGN U2119 ( .B(\mem_a[26][38] ), .A(\_zyixc_ctx_rdata_29[26][38] ));
Q_ASSIGN U2120 ( .B(\mem_a[26][39] ), .A(\_zyixc_ctx_rdata_29[26][39] ));
Q_ASSIGN U2121 ( .B(\mem_a[26][40] ), .A(\_zyixc_ctx_rdata_29[26][40] ));
Q_ASSIGN U2122 ( .B(\mem_a[26][41] ), .A(\_zyixc_ctx_rdata_29[26][41] ));
Q_ASSIGN U2123 ( .B(\mem_a[26][42] ), .A(\_zyixc_ctx_rdata_29[26][42] ));
Q_ASSIGN U2124 ( .B(\mem_a[26][43] ), .A(\_zyixc_ctx_rdata_29[26][43] ));
Q_ASSIGN U2125 ( .B(\mem_a[26][44] ), .A(\_zyixc_ctx_rdata_29[26][44] ));
Q_ASSIGN U2126 ( .B(\mem_a[26][45] ), .A(\_zyixc_ctx_rdata_29[26][45] ));
Q_ASSIGN U2127 ( .B(\mem_a[26][46] ), .A(\_zyixc_ctx_rdata_29[26][46] ));
Q_ASSIGN U2128 ( .B(\mem_a[26][47] ), .A(\_zyixc_ctx_rdata_29[26][47] ));
Q_ASSIGN U2129 ( .B(\mem_a[26][48] ), .A(\_zyixc_ctx_rdata_29[26][48] ));
Q_ASSIGN U2130 ( .B(\mem_a[26][49] ), .A(\_zyixc_ctx_rdata_29[26][49] ));
Q_ASSIGN U2131 ( .B(\mem_a[26][50] ), .A(\_zyixc_ctx_rdata_29[26][50] ));
Q_ASSIGN U2132 ( .B(\mem_a[26][51] ), .A(\_zyixc_ctx_rdata_29[26][51] ));
Q_ASSIGN U2133 ( .B(\mem_a[26][52] ), .A(\_zyixc_ctx_rdata_29[26][52] ));
Q_ASSIGN U2134 ( .B(\mem_a[26][53] ), .A(\_zyixc_ctx_rdata_29[26][53] ));
Q_ASSIGN U2135 ( .B(\mem_a[26][54] ), .A(\_zyixc_ctx_rdata_29[26][54] ));
Q_ASSIGN U2136 ( .B(\mem_a[26][55] ), .A(\_zyixc_ctx_rdata_29[26][55] ));
Q_ASSIGN U2137 ( .B(\mem_a[26][56] ), .A(\_zyixc_ctx_rdata_29[26][56] ));
Q_ASSIGN U2138 ( .B(\mem_a[26][57] ), .A(\_zyixc_ctx_rdata_29[26][57] ));
Q_ASSIGN U2139 ( .B(\mem_a[26][58] ), .A(\_zyixc_ctx_rdata_29[26][58] ));
Q_ASSIGN U2140 ( .B(\mem_a[26][59] ), .A(\_zyixc_ctx_rdata_29[26][59] ));
Q_ASSIGN U2141 ( .B(\mem_a[26][60] ), .A(\_zyixc_ctx_rdata_29[26][60] ));
Q_ASSIGN U2142 ( .B(\mem_a[26][61] ), .A(\_zyixc_ctx_rdata_29[26][61] ));
Q_ASSIGN U2143 ( .B(\mem_a[26][62] ), .A(\_zyixc_ctx_rdata_29[26][62] ));
Q_ASSIGN U2144 ( .B(\mem_a[26][63] ), .A(\_zyixc_ctx_rdata_29[26][63] ));
Q_ASSIGN U2145 ( .B(\mem_a[27][0] ), .A(\_zyixc_ctx_rdata_29[27][0] ));
Q_ASSIGN U2146 ( .B(\mem_a[27][1] ), .A(\_zyixc_ctx_rdata_29[27][1] ));
Q_ASSIGN U2147 ( .B(\mem_a[27][2] ), .A(\_zyixc_ctx_rdata_29[27][2] ));
Q_ASSIGN U2148 ( .B(\mem_a[27][3] ), .A(\_zyixc_ctx_rdata_29[27][3] ));
Q_ASSIGN U2149 ( .B(\mem_a[27][4] ), .A(\_zyixc_ctx_rdata_29[27][4] ));
Q_ASSIGN U2150 ( .B(\mem_a[27][5] ), .A(\_zyixc_ctx_rdata_29[27][5] ));
Q_ASSIGN U2151 ( .B(\mem_a[27][6] ), .A(\_zyixc_ctx_rdata_29[27][6] ));
Q_ASSIGN U2152 ( .B(\mem_a[27][7] ), .A(\_zyixc_ctx_rdata_29[27][7] ));
Q_ASSIGN U2153 ( .B(\mem_a[27][8] ), .A(\_zyixc_ctx_rdata_29[27][8] ));
Q_ASSIGN U2154 ( .B(\mem_a[27][9] ), .A(\_zyixc_ctx_rdata_29[27][9] ));
Q_ASSIGN U2155 ( .B(\mem_a[27][10] ), .A(\_zyixc_ctx_rdata_29[27][10] ));
Q_ASSIGN U2156 ( .B(\mem_a[27][11] ), .A(\_zyixc_ctx_rdata_29[27][11] ));
Q_ASSIGN U2157 ( .B(\mem_a[27][12] ), .A(\_zyixc_ctx_rdata_29[27][12] ));
Q_ASSIGN U2158 ( .B(\mem_a[27][13] ), .A(\_zyixc_ctx_rdata_29[27][13] ));
Q_ASSIGN U2159 ( .B(\mem_a[27][14] ), .A(\_zyixc_ctx_rdata_29[27][14] ));
Q_ASSIGN U2160 ( .B(\mem_a[27][15] ), .A(\_zyixc_ctx_rdata_29[27][15] ));
Q_ASSIGN U2161 ( .B(\mem_a[27][16] ), .A(\_zyixc_ctx_rdata_29[27][16] ));
Q_ASSIGN U2162 ( .B(\mem_a[27][17] ), .A(\_zyixc_ctx_rdata_29[27][17] ));
Q_ASSIGN U2163 ( .B(\mem_a[27][18] ), .A(\_zyixc_ctx_rdata_29[27][18] ));
Q_ASSIGN U2164 ( .B(\mem_a[27][19] ), .A(\_zyixc_ctx_rdata_29[27][19] ));
Q_ASSIGN U2165 ( .B(\mem_a[27][20] ), .A(\_zyixc_ctx_rdata_29[27][20] ));
Q_ASSIGN U2166 ( .B(\mem_a[27][21] ), .A(\_zyixc_ctx_rdata_29[27][21] ));
Q_ASSIGN U2167 ( .B(\mem_a[27][22] ), .A(\_zyixc_ctx_rdata_29[27][22] ));
Q_ASSIGN U2168 ( .B(\mem_a[27][23] ), .A(\_zyixc_ctx_rdata_29[27][23] ));
Q_ASSIGN U2169 ( .B(\mem_a[27][24] ), .A(\_zyixc_ctx_rdata_29[27][24] ));
Q_ASSIGN U2170 ( .B(\mem_a[27][25] ), .A(\_zyixc_ctx_rdata_29[27][25] ));
Q_ASSIGN U2171 ( .B(\mem_a[27][26] ), .A(\_zyixc_ctx_rdata_29[27][26] ));
Q_ASSIGN U2172 ( .B(\mem_a[27][27] ), .A(\_zyixc_ctx_rdata_29[27][27] ));
Q_ASSIGN U2173 ( .B(\mem_a[27][28] ), .A(\_zyixc_ctx_rdata_29[27][28] ));
Q_ASSIGN U2174 ( .B(\mem_a[27][29] ), .A(\_zyixc_ctx_rdata_29[27][29] ));
Q_ASSIGN U2175 ( .B(\mem_a[27][30] ), .A(\_zyixc_ctx_rdata_29[27][30] ));
Q_ASSIGN U2176 ( .B(\mem_a[27][31] ), .A(\_zyixc_ctx_rdata_29[27][31] ));
Q_ASSIGN U2177 ( .B(\mem_a[27][32] ), .A(\_zyixc_ctx_rdata_29[27][32] ));
Q_ASSIGN U2178 ( .B(\mem_a[27][33] ), .A(\_zyixc_ctx_rdata_29[27][33] ));
Q_ASSIGN U2179 ( .B(\mem_a[27][34] ), .A(\_zyixc_ctx_rdata_29[27][34] ));
Q_ASSIGN U2180 ( .B(\mem_a[27][35] ), .A(\_zyixc_ctx_rdata_29[27][35] ));
Q_ASSIGN U2181 ( .B(\mem_a[27][36] ), .A(\_zyixc_ctx_rdata_29[27][36] ));
Q_ASSIGN U2182 ( .B(\mem_a[27][37] ), .A(\_zyixc_ctx_rdata_29[27][37] ));
Q_ASSIGN U2183 ( .B(\mem_a[27][38] ), .A(\_zyixc_ctx_rdata_29[27][38] ));
Q_ASSIGN U2184 ( .B(\mem_a[27][39] ), .A(\_zyixc_ctx_rdata_29[27][39] ));
Q_ASSIGN U2185 ( .B(\mem_a[27][40] ), .A(\_zyixc_ctx_rdata_29[27][40] ));
Q_ASSIGN U2186 ( .B(\mem_a[27][41] ), .A(\_zyixc_ctx_rdata_29[27][41] ));
Q_ASSIGN U2187 ( .B(\mem_a[27][42] ), .A(\_zyixc_ctx_rdata_29[27][42] ));
Q_ASSIGN U2188 ( .B(\mem_a[27][43] ), .A(\_zyixc_ctx_rdata_29[27][43] ));
Q_ASSIGN U2189 ( .B(\mem_a[27][44] ), .A(\_zyixc_ctx_rdata_29[27][44] ));
Q_ASSIGN U2190 ( .B(\mem_a[27][45] ), .A(\_zyixc_ctx_rdata_29[27][45] ));
Q_ASSIGN U2191 ( .B(\mem_a[27][46] ), .A(\_zyixc_ctx_rdata_29[27][46] ));
Q_ASSIGN U2192 ( .B(\mem_a[27][47] ), .A(\_zyixc_ctx_rdata_29[27][47] ));
Q_ASSIGN U2193 ( .B(\mem_a[27][48] ), .A(\_zyixc_ctx_rdata_29[27][48] ));
Q_ASSIGN U2194 ( .B(\mem_a[27][49] ), .A(\_zyixc_ctx_rdata_29[27][49] ));
Q_ASSIGN U2195 ( .B(\mem_a[27][50] ), .A(\_zyixc_ctx_rdata_29[27][50] ));
Q_ASSIGN U2196 ( .B(\mem_a[27][51] ), .A(\_zyixc_ctx_rdata_29[27][51] ));
Q_ASSIGN U2197 ( .B(\mem_a[27][52] ), .A(\_zyixc_ctx_rdata_29[27][52] ));
Q_ASSIGN U2198 ( .B(\mem_a[27][53] ), .A(\_zyixc_ctx_rdata_29[27][53] ));
Q_ASSIGN U2199 ( .B(\mem_a[27][54] ), .A(\_zyixc_ctx_rdata_29[27][54] ));
Q_ASSIGN U2200 ( .B(\mem_a[27][55] ), .A(\_zyixc_ctx_rdata_29[27][55] ));
Q_ASSIGN U2201 ( .B(\mem_a[27][56] ), .A(\_zyixc_ctx_rdata_29[27][56] ));
Q_ASSIGN U2202 ( .B(\mem_a[27][57] ), .A(\_zyixc_ctx_rdata_29[27][57] ));
Q_ASSIGN U2203 ( .B(\mem_a[27][58] ), .A(\_zyixc_ctx_rdata_29[27][58] ));
Q_ASSIGN U2204 ( .B(\mem_a[27][59] ), .A(\_zyixc_ctx_rdata_29[27][59] ));
Q_ASSIGN U2205 ( .B(\mem_a[27][60] ), .A(\_zyixc_ctx_rdata_29[27][60] ));
Q_ASSIGN U2206 ( .B(\mem_a[27][61] ), .A(\_zyixc_ctx_rdata_29[27][61] ));
Q_ASSIGN U2207 ( .B(\mem_a[27][62] ), .A(\_zyixc_ctx_rdata_29[27][62] ));
Q_ASSIGN U2208 ( .B(\mem_a[27][63] ), .A(\_zyixc_ctx_rdata_29[27][63] ));
Q_ASSIGN U2209 ( .B(\mem_a[28][0] ), .A(\_zyixc_ctx_rdata_29[28][0] ));
Q_ASSIGN U2210 ( .B(\mem_a[28][1] ), .A(\_zyixc_ctx_rdata_29[28][1] ));
Q_ASSIGN U2211 ( .B(\mem_a[28][2] ), .A(\_zyixc_ctx_rdata_29[28][2] ));
Q_ASSIGN U2212 ( .B(\mem_a[28][3] ), .A(\_zyixc_ctx_rdata_29[28][3] ));
Q_ASSIGN U2213 ( .B(\mem_a[28][4] ), .A(\_zyixc_ctx_rdata_29[28][4] ));
Q_ASSIGN U2214 ( .B(\mem_a[28][5] ), .A(\_zyixc_ctx_rdata_29[28][5] ));
Q_ASSIGN U2215 ( .B(\mem_a[28][6] ), .A(\_zyixc_ctx_rdata_29[28][6] ));
Q_ASSIGN U2216 ( .B(\mem_a[28][7] ), .A(\_zyixc_ctx_rdata_29[28][7] ));
Q_ASSIGN U2217 ( .B(\mem_a[28][8] ), .A(\_zyixc_ctx_rdata_29[28][8] ));
Q_ASSIGN U2218 ( .B(\mem_a[28][9] ), .A(\_zyixc_ctx_rdata_29[28][9] ));
Q_ASSIGN U2219 ( .B(\mem_a[28][10] ), .A(\_zyixc_ctx_rdata_29[28][10] ));
Q_ASSIGN U2220 ( .B(\mem_a[28][11] ), .A(\_zyixc_ctx_rdata_29[28][11] ));
Q_ASSIGN U2221 ( .B(\mem_a[28][12] ), .A(\_zyixc_ctx_rdata_29[28][12] ));
Q_ASSIGN U2222 ( .B(\mem_a[28][13] ), .A(\_zyixc_ctx_rdata_29[28][13] ));
Q_ASSIGN U2223 ( .B(\mem_a[28][14] ), .A(\_zyixc_ctx_rdata_29[28][14] ));
Q_ASSIGN U2224 ( .B(\mem_a[28][15] ), .A(\_zyixc_ctx_rdata_29[28][15] ));
Q_ASSIGN U2225 ( .B(\mem_a[28][16] ), .A(\_zyixc_ctx_rdata_29[28][16] ));
Q_ASSIGN U2226 ( .B(\mem_a[28][17] ), .A(\_zyixc_ctx_rdata_29[28][17] ));
Q_ASSIGN U2227 ( .B(\mem_a[28][18] ), .A(\_zyixc_ctx_rdata_29[28][18] ));
Q_ASSIGN U2228 ( .B(\mem_a[28][19] ), .A(\_zyixc_ctx_rdata_29[28][19] ));
Q_ASSIGN U2229 ( .B(\mem_a[28][20] ), .A(\_zyixc_ctx_rdata_29[28][20] ));
Q_ASSIGN U2230 ( .B(\mem_a[28][21] ), .A(\_zyixc_ctx_rdata_29[28][21] ));
Q_ASSIGN U2231 ( .B(\mem_a[28][22] ), .A(\_zyixc_ctx_rdata_29[28][22] ));
Q_ASSIGN U2232 ( .B(\mem_a[28][23] ), .A(\_zyixc_ctx_rdata_29[28][23] ));
Q_ASSIGN U2233 ( .B(\mem_a[28][24] ), .A(\_zyixc_ctx_rdata_29[28][24] ));
Q_ASSIGN U2234 ( .B(\mem_a[28][25] ), .A(\_zyixc_ctx_rdata_29[28][25] ));
Q_ASSIGN U2235 ( .B(\mem_a[28][26] ), .A(\_zyixc_ctx_rdata_29[28][26] ));
Q_ASSIGN U2236 ( .B(\mem_a[28][27] ), .A(\_zyixc_ctx_rdata_29[28][27] ));
Q_ASSIGN U2237 ( .B(\mem_a[28][28] ), .A(\_zyixc_ctx_rdata_29[28][28] ));
Q_ASSIGN U2238 ( .B(\mem_a[28][29] ), .A(\_zyixc_ctx_rdata_29[28][29] ));
Q_ASSIGN U2239 ( .B(\mem_a[28][30] ), .A(\_zyixc_ctx_rdata_29[28][30] ));
Q_ASSIGN U2240 ( .B(\mem_a[28][31] ), .A(\_zyixc_ctx_rdata_29[28][31] ));
Q_ASSIGN U2241 ( .B(\mem_a[28][32] ), .A(\_zyixc_ctx_rdata_29[28][32] ));
Q_ASSIGN U2242 ( .B(\mem_a[28][33] ), .A(\_zyixc_ctx_rdata_29[28][33] ));
Q_ASSIGN U2243 ( .B(\mem_a[28][34] ), .A(\_zyixc_ctx_rdata_29[28][34] ));
Q_ASSIGN U2244 ( .B(\mem_a[28][35] ), .A(\_zyixc_ctx_rdata_29[28][35] ));
Q_ASSIGN U2245 ( .B(\mem_a[28][36] ), .A(\_zyixc_ctx_rdata_29[28][36] ));
Q_ASSIGN U2246 ( .B(\mem_a[28][37] ), .A(\_zyixc_ctx_rdata_29[28][37] ));
Q_ASSIGN U2247 ( .B(\mem_a[28][38] ), .A(\_zyixc_ctx_rdata_29[28][38] ));
Q_ASSIGN U2248 ( .B(\mem_a[28][39] ), .A(\_zyixc_ctx_rdata_29[28][39] ));
Q_ASSIGN U2249 ( .B(\mem_a[28][40] ), .A(\_zyixc_ctx_rdata_29[28][40] ));
Q_ASSIGN U2250 ( .B(\mem_a[28][41] ), .A(\_zyixc_ctx_rdata_29[28][41] ));
Q_ASSIGN U2251 ( .B(\mem_a[28][42] ), .A(\_zyixc_ctx_rdata_29[28][42] ));
Q_ASSIGN U2252 ( .B(\mem_a[28][43] ), .A(\_zyixc_ctx_rdata_29[28][43] ));
Q_ASSIGN U2253 ( .B(\mem_a[28][44] ), .A(\_zyixc_ctx_rdata_29[28][44] ));
Q_ASSIGN U2254 ( .B(\mem_a[28][45] ), .A(\_zyixc_ctx_rdata_29[28][45] ));
Q_ASSIGN U2255 ( .B(\mem_a[28][46] ), .A(\_zyixc_ctx_rdata_29[28][46] ));
Q_ASSIGN U2256 ( .B(\mem_a[28][47] ), .A(\_zyixc_ctx_rdata_29[28][47] ));
Q_ASSIGN U2257 ( .B(\mem_a[28][48] ), .A(\_zyixc_ctx_rdata_29[28][48] ));
Q_ASSIGN U2258 ( .B(\mem_a[28][49] ), .A(\_zyixc_ctx_rdata_29[28][49] ));
Q_ASSIGN U2259 ( .B(\mem_a[28][50] ), .A(\_zyixc_ctx_rdata_29[28][50] ));
Q_ASSIGN U2260 ( .B(\mem_a[28][51] ), .A(\_zyixc_ctx_rdata_29[28][51] ));
Q_ASSIGN U2261 ( .B(\mem_a[28][52] ), .A(\_zyixc_ctx_rdata_29[28][52] ));
Q_ASSIGN U2262 ( .B(\mem_a[28][53] ), .A(\_zyixc_ctx_rdata_29[28][53] ));
Q_ASSIGN U2263 ( .B(\mem_a[28][54] ), .A(\_zyixc_ctx_rdata_29[28][54] ));
Q_ASSIGN U2264 ( .B(\mem_a[28][55] ), .A(\_zyixc_ctx_rdata_29[28][55] ));
Q_ASSIGN U2265 ( .B(\mem_a[28][56] ), .A(\_zyixc_ctx_rdata_29[28][56] ));
Q_ASSIGN U2266 ( .B(\mem_a[28][57] ), .A(\_zyixc_ctx_rdata_29[28][57] ));
Q_ASSIGN U2267 ( .B(\mem_a[28][58] ), .A(\_zyixc_ctx_rdata_29[28][58] ));
Q_ASSIGN U2268 ( .B(\mem_a[28][59] ), .A(\_zyixc_ctx_rdata_29[28][59] ));
Q_ASSIGN U2269 ( .B(\mem_a[28][60] ), .A(\_zyixc_ctx_rdata_29[28][60] ));
Q_ASSIGN U2270 ( .B(\mem_a[28][61] ), .A(\_zyixc_ctx_rdata_29[28][61] ));
Q_ASSIGN U2271 ( .B(\mem_a[28][62] ), .A(\_zyixc_ctx_rdata_29[28][62] ));
Q_ASSIGN U2272 ( .B(\mem_a[28][63] ), .A(\_zyixc_ctx_rdata_29[28][63] ));
Q_ASSIGN U2273 ( .B(\mem_a[29][0] ), .A(\_zyixc_ctx_rdata_29[29][0] ));
Q_ASSIGN U2274 ( .B(\mem_a[29][1] ), .A(\_zyixc_ctx_rdata_29[29][1] ));
Q_ASSIGN U2275 ( .B(\mem_a[29][2] ), .A(\_zyixc_ctx_rdata_29[29][2] ));
Q_ASSIGN U2276 ( .B(\mem_a[29][3] ), .A(\_zyixc_ctx_rdata_29[29][3] ));
Q_ASSIGN U2277 ( .B(\mem_a[29][4] ), .A(\_zyixc_ctx_rdata_29[29][4] ));
Q_ASSIGN U2278 ( .B(\mem_a[29][5] ), .A(\_zyixc_ctx_rdata_29[29][5] ));
Q_ASSIGN U2279 ( .B(\mem_a[29][6] ), .A(\_zyixc_ctx_rdata_29[29][6] ));
Q_ASSIGN U2280 ( .B(\mem_a[29][7] ), .A(\_zyixc_ctx_rdata_29[29][7] ));
Q_ASSIGN U2281 ( .B(\mem_a[29][8] ), .A(\_zyixc_ctx_rdata_29[29][8] ));
Q_ASSIGN U2282 ( .B(\mem_a[29][9] ), .A(\_zyixc_ctx_rdata_29[29][9] ));
Q_ASSIGN U2283 ( .B(\mem_a[29][10] ), .A(\_zyixc_ctx_rdata_29[29][10] ));
Q_ASSIGN U2284 ( .B(\mem_a[29][11] ), .A(\_zyixc_ctx_rdata_29[29][11] ));
Q_ASSIGN U2285 ( .B(\mem_a[29][12] ), .A(\_zyixc_ctx_rdata_29[29][12] ));
Q_ASSIGN U2286 ( .B(\mem_a[29][13] ), .A(\_zyixc_ctx_rdata_29[29][13] ));
Q_ASSIGN U2287 ( .B(\mem_a[29][14] ), .A(\_zyixc_ctx_rdata_29[29][14] ));
Q_ASSIGN U2288 ( .B(\mem_a[29][15] ), .A(\_zyixc_ctx_rdata_29[29][15] ));
Q_ASSIGN U2289 ( .B(\mem_a[29][16] ), .A(\_zyixc_ctx_rdata_29[29][16] ));
Q_ASSIGN U2290 ( .B(\mem_a[29][17] ), .A(\_zyixc_ctx_rdata_29[29][17] ));
Q_ASSIGN U2291 ( .B(\mem_a[29][18] ), .A(\_zyixc_ctx_rdata_29[29][18] ));
Q_ASSIGN U2292 ( .B(\mem_a[29][19] ), .A(\_zyixc_ctx_rdata_29[29][19] ));
Q_ASSIGN U2293 ( .B(\mem_a[29][20] ), .A(\_zyixc_ctx_rdata_29[29][20] ));
Q_ASSIGN U2294 ( .B(\mem_a[29][21] ), .A(\_zyixc_ctx_rdata_29[29][21] ));
Q_ASSIGN U2295 ( .B(\mem_a[29][22] ), .A(\_zyixc_ctx_rdata_29[29][22] ));
Q_ASSIGN U2296 ( .B(\mem_a[29][23] ), .A(\_zyixc_ctx_rdata_29[29][23] ));
Q_ASSIGN U2297 ( .B(\mem_a[29][24] ), .A(\_zyixc_ctx_rdata_29[29][24] ));
Q_ASSIGN U2298 ( .B(\mem_a[29][25] ), .A(\_zyixc_ctx_rdata_29[29][25] ));
Q_ASSIGN U2299 ( .B(\mem_a[29][26] ), .A(\_zyixc_ctx_rdata_29[29][26] ));
Q_ASSIGN U2300 ( .B(\mem_a[29][27] ), .A(\_zyixc_ctx_rdata_29[29][27] ));
Q_ASSIGN U2301 ( .B(\mem_a[29][28] ), .A(\_zyixc_ctx_rdata_29[29][28] ));
Q_ASSIGN U2302 ( .B(\mem_a[29][29] ), .A(\_zyixc_ctx_rdata_29[29][29] ));
Q_ASSIGN U2303 ( .B(\mem_a[29][30] ), .A(\_zyixc_ctx_rdata_29[29][30] ));
Q_ASSIGN U2304 ( .B(\mem_a[29][31] ), .A(\_zyixc_ctx_rdata_29[29][31] ));
Q_ASSIGN U2305 ( .B(\mem_a[29][32] ), .A(\_zyixc_ctx_rdata_29[29][32] ));
Q_ASSIGN U2306 ( .B(\mem_a[29][33] ), .A(\_zyixc_ctx_rdata_29[29][33] ));
Q_ASSIGN U2307 ( .B(\mem_a[29][34] ), .A(\_zyixc_ctx_rdata_29[29][34] ));
Q_ASSIGN U2308 ( .B(\mem_a[29][35] ), .A(\_zyixc_ctx_rdata_29[29][35] ));
Q_ASSIGN U2309 ( .B(\mem_a[29][36] ), .A(\_zyixc_ctx_rdata_29[29][36] ));
Q_ASSIGN U2310 ( .B(\mem_a[29][37] ), .A(\_zyixc_ctx_rdata_29[29][37] ));
Q_ASSIGN U2311 ( .B(\mem_a[29][38] ), .A(\_zyixc_ctx_rdata_29[29][38] ));
Q_ASSIGN U2312 ( .B(\mem_a[29][39] ), .A(\_zyixc_ctx_rdata_29[29][39] ));
Q_ASSIGN U2313 ( .B(\mem_a[29][40] ), .A(\_zyixc_ctx_rdata_29[29][40] ));
Q_ASSIGN U2314 ( .B(\mem_a[29][41] ), .A(\_zyixc_ctx_rdata_29[29][41] ));
Q_ASSIGN U2315 ( .B(\mem_a[29][42] ), .A(\_zyixc_ctx_rdata_29[29][42] ));
Q_ASSIGN U2316 ( .B(\mem_a[29][43] ), .A(\_zyixc_ctx_rdata_29[29][43] ));
Q_ASSIGN U2317 ( .B(\mem_a[29][44] ), .A(\_zyixc_ctx_rdata_29[29][44] ));
Q_ASSIGN U2318 ( .B(\mem_a[29][45] ), .A(\_zyixc_ctx_rdata_29[29][45] ));
Q_ASSIGN U2319 ( .B(\mem_a[29][46] ), .A(\_zyixc_ctx_rdata_29[29][46] ));
Q_ASSIGN U2320 ( .B(\mem_a[29][47] ), .A(\_zyixc_ctx_rdata_29[29][47] ));
Q_ASSIGN U2321 ( .B(\mem_a[29][48] ), .A(\_zyixc_ctx_rdata_29[29][48] ));
Q_ASSIGN U2322 ( .B(\mem_a[29][49] ), .A(\_zyixc_ctx_rdata_29[29][49] ));
Q_ASSIGN U2323 ( .B(\mem_a[29][50] ), .A(\_zyixc_ctx_rdata_29[29][50] ));
Q_ASSIGN U2324 ( .B(\mem_a[29][51] ), .A(\_zyixc_ctx_rdata_29[29][51] ));
Q_ASSIGN U2325 ( .B(\mem_a[29][52] ), .A(\_zyixc_ctx_rdata_29[29][52] ));
Q_ASSIGN U2326 ( .B(\mem_a[29][53] ), .A(\_zyixc_ctx_rdata_29[29][53] ));
Q_ASSIGN U2327 ( .B(\mem_a[29][54] ), .A(\_zyixc_ctx_rdata_29[29][54] ));
Q_ASSIGN U2328 ( .B(\mem_a[29][55] ), .A(\_zyixc_ctx_rdata_29[29][55] ));
Q_ASSIGN U2329 ( .B(\mem_a[29][56] ), .A(\_zyixc_ctx_rdata_29[29][56] ));
Q_ASSIGN U2330 ( .B(\mem_a[29][57] ), .A(\_zyixc_ctx_rdata_29[29][57] ));
Q_ASSIGN U2331 ( .B(\mem_a[29][58] ), .A(\_zyixc_ctx_rdata_29[29][58] ));
Q_ASSIGN U2332 ( .B(\mem_a[29][59] ), .A(\_zyixc_ctx_rdata_29[29][59] ));
Q_ASSIGN U2333 ( .B(\mem_a[29][60] ), .A(\_zyixc_ctx_rdata_29[29][60] ));
Q_ASSIGN U2334 ( .B(\mem_a[29][61] ), .A(\_zyixc_ctx_rdata_29[29][61] ));
Q_ASSIGN U2335 ( .B(\mem_a[29][62] ), .A(\_zyixc_ctx_rdata_29[29][62] ));
Q_ASSIGN U2336 ( .B(\mem_a[29][63] ), .A(\_zyixc_ctx_rdata_29[29][63] ));
Q_ASSIGN U2337 ( .B(\mem_a[30][0] ), .A(\_zyixc_ctx_rdata_29[30][0] ));
Q_ASSIGN U2338 ( .B(\mem_a[30][1] ), .A(\_zyixc_ctx_rdata_29[30][1] ));
Q_ASSIGN U2339 ( .B(\mem_a[30][2] ), .A(\_zyixc_ctx_rdata_29[30][2] ));
Q_ASSIGN U2340 ( .B(\mem_a[30][3] ), .A(\_zyixc_ctx_rdata_29[30][3] ));
Q_ASSIGN U2341 ( .B(\mem_a[30][4] ), .A(\_zyixc_ctx_rdata_29[30][4] ));
Q_ASSIGN U2342 ( .B(\mem_a[30][5] ), .A(\_zyixc_ctx_rdata_29[30][5] ));
Q_ASSIGN U2343 ( .B(\mem_a[30][6] ), .A(\_zyixc_ctx_rdata_29[30][6] ));
Q_ASSIGN U2344 ( .B(\mem_a[30][7] ), .A(\_zyixc_ctx_rdata_29[30][7] ));
Q_ASSIGN U2345 ( .B(\mem_a[30][8] ), .A(\_zyixc_ctx_rdata_29[30][8] ));
Q_ASSIGN U2346 ( .B(\mem_a[30][9] ), .A(\_zyixc_ctx_rdata_29[30][9] ));
Q_ASSIGN U2347 ( .B(\mem_a[30][10] ), .A(\_zyixc_ctx_rdata_29[30][10] ));
Q_ASSIGN U2348 ( .B(\mem_a[30][11] ), .A(\_zyixc_ctx_rdata_29[30][11] ));
Q_ASSIGN U2349 ( .B(\mem_a[30][12] ), .A(\_zyixc_ctx_rdata_29[30][12] ));
Q_ASSIGN U2350 ( .B(\mem_a[30][13] ), .A(\_zyixc_ctx_rdata_29[30][13] ));
Q_ASSIGN U2351 ( .B(\mem_a[30][14] ), .A(\_zyixc_ctx_rdata_29[30][14] ));
Q_ASSIGN U2352 ( .B(\mem_a[30][15] ), .A(\_zyixc_ctx_rdata_29[30][15] ));
Q_ASSIGN U2353 ( .B(\mem_a[30][16] ), .A(\_zyixc_ctx_rdata_29[30][16] ));
Q_ASSIGN U2354 ( .B(\mem_a[30][17] ), .A(\_zyixc_ctx_rdata_29[30][17] ));
Q_ASSIGN U2355 ( .B(\mem_a[30][18] ), .A(\_zyixc_ctx_rdata_29[30][18] ));
Q_ASSIGN U2356 ( .B(\mem_a[30][19] ), .A(\_zyixc_ctx_rdata_29[30][19] ));
Q_ASSIGN U2357 ( .B(\mem_a[30][20] ), .A(\_zyixc_ctx_rdata_29[30][20] ));
Q_ASSIGN U2358 ( .B(\mem_a[30][21] ), .A(\_zyixc_ctx_rdata_29[30][21] ));
Q_ASSIGN U2359 ( .B(\mem_a[30][22] ), .A(\_zyixc_ctx_rdata_29[30][22] ));
Q_ASSIGN U2360 ( .B(\mem_a[30][23] ), .A(\_zyixc_ctx_rdata_29[30][23] ));
Q_ASSIGN U2361 ( .B(\mem_a[30][24] ), .A(\_zyixc_ctx_rdata_29[30][24] ));
Q_ASSIGN U2362 ( .B(\mem_a[30][25] ), .A(\_zyixc_ctx_rdata_29[30][25] ));
Q_ASSIGN U2363 ( .B(\mem_a[30][26] ), .A(\_zyixc_ctx_rdata_29[30][26] ));
Q_ASSIGN U2364 ( .B(\mem_a[30][27] ), .A(\_zyixc_ctx_rdata_29[30][27] ));
Q_ASSIGN U2365 ( .B(\mem_a[30][28] ), .A(\_zyixc_ctx_rdata_29[30][28] ));
Q_ASSIGN U2366 ( .B(\mem_a[30][29] ), .A(\_zyixc_ctx_rdata_29[30][29] ));
Q_ASSIGN U2367 ( .B(\mem_a[30][30] ), .A(\_zyixc_ctx_rdata_29[30][30] ));
Q_ASSIGN U2368 ( .B(\mem_a[30][31] ), .A(\_zyixc_ctx_rdata_29[30][31] ));
Q_ASSIGN U2369 ( .B(\mem_a[30][32] ), .A(\_zyixc_ctx_rdata_29[30][32] ));
Q_ASSIGN U2370 ( .B(\mem_a[30][33] ), .A(\_zyixc_ctx_rdata_29[30][33] ));
Q_ASSIGN U2371 ( .B(\mem_a[30][34] ), .A(\_zyixc_ctx_rdata_29[30][34] ));
Q_ASSIGN U2372 ( .B(\mem_a[30][35] ), .A(\_zyixc_ctx_rdata_29[30][35] ));
Q_ASSIGN U2373 ( .B(\mem_a[30][36] ), .A(\_zyixc_ctx_rdata_29[30][36] ));
Q_ASSIGN U2374 ( .B(\mem_a[30][37] ), .A(\_zyixc_ctx_rdata_29[30][37] ));
Q_ASSIGN U2375 ( .B(\mem_a[30][38] ), .A(\_zyixc_ctx_rdata_29[30][38] ));
Q_ASSIGN U2376 ( .B(\mem_a[30][39] ), .A(\_zyixc_ctx_rdata_29[30][39] ));
Q_ASSIGN U2377 ( .B(\mem_a[30][40] ), .A(\_zyixc_ctx_rdata_29[30][40] ));
Q_ASSIGN U2378 ( .B(\mem_a[30][41] ), .A(\_zyixc_ctx_rdata_29[30][41] ));
Q_ASSIGN U2379 ( .B(\mem_a[30][42] ), .A(\_zyixc_ctx_rdata_29[30][42] ));
Q_ASSIGN U2380 ( .B(\mem_a[30][43] ), .A(\_zyixc_ctx_rdata_29[30][43] ));
Q_ASSIGN U2381 ( .B(\mem_a[30][44] ), .A(\_zyixc_ctx_rdata_29[30][44] ));
Q_ASSIGN U2382 ( .B(\mem_a[30][45] ), .A(\_zyixc_ctx_rdata_29[30][45] ));
Q_ASSIGN U2383 ( .B(\mem_a[30][46] ), .A(\_zyixc_ctx_rdata_29[30][46] ));
Q_ASSIGN U2384 ( .B(\mem_a[30][47] ), .A(\_zyixc_ctx_rdata_29[30][47] ));
Q_ASSIGN U2385 ( .B(\mem_a[30][48] ), .A(\_zyixc_ctx_rdata_29[30][48] ));
Q_ASSIGN U2386 ( .B(\mem_a[30][49] ), .A(\_zyixc_ctx_rdata_29[30][49] ));
Q_ASSIGN U2387 ( .B(\mem_a[30][50] ), .A(\_zyixc_ctx_rdata_29[30][50] ));
Q_ASSIGN U2388 ( .B(\mem_a[30][51] ), .A(\_zyixc_ctx_rdata_29[30][51] ));
Q_ASSIGN U2389 ( .B(\mem_a[30][52] ), .A(\_zyixc_ctx_rdata_29[30][52] ));
Q_ASSIGN U2390 ( .B(\mem_a[30][53] ), .A(\_zyixc_ctx_rdata_29[30][53] ));
Q_ASSIGN U2391 ( .B(\mem_a[30][54] ), .A(\_zyixc_ctx_rdata_29[30][54] ));
Q_ASSIGN U2392 ( .B(\mem_a[30][55] ), .A(\_zyixc_ctx_rdata_29[30][55] ));
Q_ASSIGN U2393 ( .B(\mem_a[30][56] ), .A(\_zyixc_ctx_rdata_29[30][56] ));
Q_ASSIGN U2394 ( .B(\mem_a[30][57] ), .A(\_zyixc_ctx_rdata_29[30][57] ));
Q_ASSIGN U2395 ( .B(\mem_a[30][58] ), .A(\_zyixc_ctx_rdata_29[30][58] ));
Q_ASSIGN U2396 ( .B(\mem_a[30][59] ), .A(\_zyixc_ctx_rdata_29[30][59] ));
Q_ASSIGN U2397 ( .B(\mem_a[30][60] ), .A(\_zyixc_ctx_rdata_29[30][60] ));
Q_ASSIGN U2398 ( .B(\mem_a[30][61] ), .A(\_zyixc_ctx_rdata_29[30][61] ));
Q_ASSIGN U2399 ( .B(\mem_a[30][62] ), .A(\_zyixc_ctx_rdata_29[30][62] ));
Q_ASSIGN U2400 ( .B(\mem_a[30][63] ), .A(\_zyixc_ctx_rdata_29[30][63] ));
Q_ASSIGN U2401 ( .B(\mem_a[31][0] ), .A(\_zyixc_ctx_rdata_29[31][0] ));
Q_ASSIGN U2402 ( .B(\mem_a[31][1] ), .A(\_zyixc_ctx_rdata_29[31][1] ));
Q_ASSIGN U2403 ( .B(\mem_a[31][2] ), .A(\_zyixc_ctx_rdata_29[31][2] ));
Q_ASSIGN U2404 ( .B(\mem_a[31][3] ), .A(\_zyixc_ctx_rdata_29[31][3] ));
Q_ASSIGN U2405 ( .B(\mem_a[31][4] ), .A(\_zyixc_ctx_rdata_29[31][4] ));
Q_ASSIGN U2406 ( .B(\mem_a[31][5] ), .A(\_zyixc_ctx_rdata_29[31][5] ));
Q_ASSIGN U2407 ( .B(\mem_a[31][6] ), .A(\_zyixc_ctx_rdata_29[31][6] ));
Q_ASSIGN U2408 ( .B(\mem_a[31][7] ), .A(\_zyixc_ctx_rdata_29[31][7] ));
Q_ASSIGN U2409 ( .B(\mem_a[31][8] ), .A(\_zyixc_ctx_rdata_29[31][8] ));
Q_ASSIGN U2410 ( .B(\mem_a[31][9] ), .A(\_zyixc_ctx_rdata_29[31][9] ));
Q_ASSIGN U2411 ( .B(\mem_a[31][10] ), .A(\_zyixc_ctx_rdata_29[31][10] ));
Q_ASSIGN U2412 ( .B(\mem_a[31][11] ), .A(\_zyixc_ctx_rdata_29[31][11] ));
Q_ASSIGN U2413 ( .B(\mem_a[31][12] ), .A(\_zyixc_ctx_rdata_29[31][12] ));
Q_ASSIGN U2414 ( .B(\mem_a[31][13] ), .A(\_zyixc_ctx_rdata_29[31][13] ));
Q_ASSIGN U2415 ( .B(\mem_a[31][14] ), .A(\_zyixc_ctx_rdata_29[31][14] ));
Q_ASSIGN U2416 ( .B(\mem_a[31][15] ), .A(\_zyixc_ctx_rdata_29[31][15] ));
Q_ASSIGN U2417 ( .B(\mem_a[31][16] ), .A(\_zyixc_ctx_rdata_29[31][16] ));
Q_ASSIGN U2418 ( .B(\mem_a[31][17] ), .A(\_zyixc_ctx_rdata_29[31][17] ));
Q_ASSIGN U2419 ( .B(\mem_a[31][18] ), .A(\_zyixc_ctx_rdata_29[31][18] ));
Q_ASSIGN U2420 ( .B(\mem_a[31][19] ), .A(\_zyixc_ctx_rdata_29[31][19] ));
Q_ASSIGN U2421 ( .B(\mem_a[31][20] ), .A(\_zyixc_ctx_rdata_29[31][20] ));
Q_ASSIGN U2422 ( .B(\mem_a[31][21] ), .A(\_zyixc_ctx_rdata_29[31][21] ));
Q_ASSIGN U2423 ( .B(\mem_a[31][22] ), .A(\_zyixc_ctx_rdata_29[31][22] ));
Q_ASSIGN U2424 ( .B(\mem_a[31][23] ), .A(\_zyixc_ctx_rdata_29[31][23] ));
Q_ASSIGN U2425 ( .B(\mem_a[31][24] ), .A(\_zyixc_ctx_rdata_29[31][24] ));
Q_ASSIGN U2426 ( .B(\mem_a[31][25] ), .A(\_zyixc_ctx_rdata_29[31][25] ));
Q_ASSIGN U2427 ( .B(\mem_a[31][26] ), .A(\_zyixc_ctx_rdata_29[31][26] ));
Q_ASSIGN U2428 ( .B(\mem_a[31][27] ), .A(\_zyixc_ctx_rdata_29[31][27] ));
Q_ASSIGN U2429 ( .B(\mem_a[31][28] ), .A(\_zyixc_ctx_rdata_29[31][28] ));
Q_ASSIGN U2430 ( .B(\mem_a[31][29] ), .A(\_zyixc_ctx_rdata_29[31][29] ));
Q_ASSIGN U2431 ( .B(\mem_a[31][30] ), .A(\_zyixc_ctx_rdata_29[31][30] ));
Q_ASSIGN U2432 ( .B(\mem_a[31][31] ), .A(\_zyixc_ctx_rdata_29[31][31] ));
Q_ASSIGN U2433 ( .B(\mem_a[31][32] ), .A(\_zyixc_ctx_rdata_29[31][32] ));
Q_ASSIGN U2434 ( .B(\mem_a[31][33] ), .A(\_zyixc_ctx_rdata_29[31][33] ));
Q_ASSIGN U2435 ( .B(\mem_a[31][34] ), .A(\_zyixc_ctx_rdata_29[31][34] ));
Q_ASSIGN U2436 ( .B(\mem_a[31][35] ), .A(\_zyixc_ctx_rdata_29[31][35] ));
Q_ASSIGN U2437 ( .B(\mem_a[31][36] ), .A(\_zyixc_ctx_rdata_29[31][36] ));
Q_ASSIGN U2438 ( .B(\mem_a[31][37] ), .A(\_zyixc_ctx_rdata_29[31][37] ));
Q_ASSIGN U2439 ( .B(\mem_a[31][38] ), .A(\_zyixc_ctx_rdata_29[31][38] ));
Q_ASSIGN U2440 ( .B(\mem_a[31][39] ), .A(\_zyixc_ctx_rdata_29[31][39] ));
Q_ASSIGN U2441 ( .B(\mem_a[31][40] ), .A(\_zyixc_ctx_rdata_29[31][40] ));
Q_ASSIGN U2442 ( .B(\mem_a[31][41] ), .A(\_zyixc_ctx_rdata_29[31][41] ));
Q_ASSIGN U2443 ( .B(\mem_a[31][42] ), .A(\_zyixc_ctx_rdata_29[31][42] ));
Q_ASSIGN U2444 ( .B(\mem_a[31][43] ), .A(\_zyixc_ctx_rdata_29[31][43] ));
Q_ASSIGN U2445 ( .B(\mem_a[31][44] ), .A(\_zyixc_ctx_rdata_29[31][44] ));
Q_ASSIGN U2446 ( .B(\mem_a[31][45] ), .A(\_zyixc_ctx_rdata_29[31][45] ));
Q_ASSIGN U2447 ( .B(\mem_a[31][46] ), .A(\_zyixc_ctx_rdata_29[31][46] ));
Q_ASSIGN U2448 ( .B(\mem_a[31][47] ), .A(\_zyixc_ctx_rdata_29[31][47] ));
Q_ASSIGN U2449 ( .B(\mem_a[31][48] ), .A(\_zyixc_ctx_rdata_29[31][48] ));
Q_ASSIGN U2450 ( .B(\mem_a[31][49] ), .A(\_zyixc_ctx_rdata_29[31][49] ));
Q_ASSIGN U2451 ( .B(\mem_a[31][50] ), .A(\_zyixc_ctx_rdata_29[31][50] ));
Q_ASSIGN U2452 ( .B(\mem_a[31][51] ), .A(\_zyixc_ctx_rdata_29[31][51] ));
Q_ASSIGN U2453 ( .B(\mem_a[31][52] ), .A(\_zyixc_ctx_rdata_29[31][52] ));
Q_ASSIGN U2454 ( .B(\mem_a[31][53] ), .A(\_zyixc_ctx_rdata_29[31][53] ));
Q_ASSIGN U2455 ( .B(\mem_a[31][54] ), .A(\_zyixc_ctx_rdata_29[31][54] ));
Q_ASSIGN U2456 ( .B(\mem_a[31][55] ), .A(\_zyixc_ctx_rdata_29[31][55] ));
Q_ASSIGN U2457 ( .B(\mem_a[31][56] ), .A(\_zyixc_ctx_rdata_29[31][56] ));
Q_ASSIGN U2458 ( .B(\mem_a[31][57] ), .A(\_zyixc_ctx_rdata_29[31][57] ));
Q_ASSIGN U2459 ( .B(\mem_a[31][58] ), .A(\_zyixc_ctx_rdata_29[31][58] ));
Q_ASSIGN U2460 ( .B(\mem_a[31][59] ), .A(\_zyixc_ctx_rdata_29[31][59] ));
Q_ASSIGN U2461 ( .B(\mem_a[31][60] ), .A(\_zyixc_ctx_rdata_29[31][60] ));
Q_ASSIGN U2462 ( .B(\mem_a[31][61] ), .A(\_zyixc_ctx_rdata_29[31][61] ));
Q_ASSIGN U2463 ( .B(\mem_a[31][62] ), .A(\_zyixc_ctx_rdata_29[31][62] ));
Q_ASSIGN U2464 ( .B(\mem_a[31][63] ), .A(\_zyixc_ctx_rdata_29[31][63] ));
Q_FDP4EP \sw_rdat_REG[0] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n7), .Q(sw_rdat[0]));
Q_INV U2466 ( .A(rst_n), .Z(n323));
Q_FDP4EP \sw_rdat_REG[1] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n12), .Q(sw_rdat[1]));
Q_FDP4EP \sw_rdat_REG[2] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n17), .Q(sw_rdat[2]));
Q_FDP4EP \sw_rdat_REG[3] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n22), .Q(sw_rdat[3]));
Q_FDP4EP \sw_rdat_REG[4] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n27), .Q(sw_rdat[4]));
Q_FDP4EP \sw_rdat_REG[5] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n32), .Q(sw_rdat[5]));
Q_FDP4EP \sw_rdat_REG[6] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n37), .Q(sw_rdat[6]));
Q_FDP4EP \sw_rdat_REG[7] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n42), .Q(sw_rdat[7]));
Q_FDP4EP \sw_rdat_REG[8] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n47), .Q(sw_rdat[8]));
Q_FDP4EP \sw_rdat_REG[9] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n52), .Q(sw_rdat[9]));
Q_FDP4EP \sw_rdat_REG[10] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n57), .Q(sw_rdat[10]));
Q_FDP4EP \sw_rdat_REG[11] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n62), .Q(sw_rdat[11]));
Q_FDP4EP \sw_rdat_REG[12] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n67), .Q(sw_rdat[12]));
Q_FDP4EP \sw_rdat_REG[13] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n72), .Q(sw_rdat[13]));
Q_FDP4EP \sw_rdat_REG[14] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n77), .Q(sw_rdat[14]));
Q_FDP4EP \sw_rdat_REG[15] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n82), .Q(sw_rdat[15]));
Q_FDP4EP \sw_rdat_REG[16] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n87), .Q(sw_rdat[16]));
Q_FDP4EP \sw_rdat_REG[17] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n92), .Q(sw_rdat[17]));
Q_FDP4EP \sw_rdat_REG[18] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n97), .Q(sw_rdat[18]));
Q_FDP4EP \sw_rdat_REG[19] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n102), .Q(sw_rdat[19]));
Q_FDP4EP \sw_rdat_REG[20] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n107), .Q(sw_rdat[20]));
Q_FDP4EP \sw_rdat_REG[21] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n112), .Q(sw_rdat[21]));
Q_FDP4EP \sw_rdat_REG[22] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n117), .Q(sw_rdat[22]));
Q_FDP4EP \sw_rdat_REG[23] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n122), .Q(sw_rdat[23]));
Q_FDP4EP \sw_rdat_REG[24] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n127), .Q(sw_rdat[24]));
Q_FDP4EP \sw_rdat_REG[25] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n132), .Q(sw_rdat[25]));
Q_FDP4EP \sw_rdat_REG[26] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n137), .Q(sw_rdat[26]));
Q_FDP4EP \sw_rdat_REG[27] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n142), .Q(sw_rdat[27]));
Q_FDP4EP \sw_rdat_REG[28] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n147), .Q(sw_rdat[28]));
Q_FDP4EP \sw_rdat_REG[29] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n152), .Q(sw_rdat[29]));
Q_FDP4EP \sw_rdat_REG[30] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n157), .Q(sw_rdat[30]));
Q_FDP4EP \sw_rdat_REG[31] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n162), .Q(sw_rdat[31]));
Q_FDP4EP \sw_rdat_REG[32] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n167), .Q(sw_rdat[32]));
Q_FDP4EP \sw_rdat_REG[33] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n172), .Q(sw_rdat[33]));
Q_FDP4EP \sw_rdat_REG[34] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n177), .Q(sw_rdat[34]));
Q_FDP4EP \sw_rdat_REG[35] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n182), .Q(sw_rdat[35]));
Q_FDP4EP \sw_rdat_REG[36] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n187), .Q(sw_rdat[36]));
Q_FDP4EP \sw_rdat_REG[37] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n192), .Q(sw_rdat[37]));
Q_FDP4EP \sw_rdat_REG[38] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n197), .Q(sw_rdat[38]));
Q_FDP4EP \sw_rdat_REG[39] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n202), .Q(sw_rdat[39]));
Q_FDP4EP \sw_rdat_REG[40] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n207), .Q(sw_rdat[40]));
Q_FDP4EP \sw_rdat_REG[41] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n212), .Q(sw_rdat[41]));
Q_FDP4EP \sw_rdat_REG[42] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n217), .Q(sw_rdat[42]));
Q_FDP4EP \sw_rdat_REG[43] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n222), .Q(sw_rdat[43]));
Q_FDP4EP \sw_rdat_REG[44] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n227), .Q(sw_rdat[44]));
Q_FDP4EP \sw_rdat_REG[45] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n232), .Q(sw_rdat[45]));
Q_FDP4EP \sw_rdat_REG[46] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n237), .Q(sw_rdat[46]));
Q_FDP4EP \sw_rdat_REG[47] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n242), .Q(sw_rdat[47]));
Q_FDP4EP \sw_rdat_REG[48] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n247), .Q(sw_rdat[48]));
Q_FDP4EP \sw_rdat_REG[49] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n252), .Q(sw_rdat[49]));
Q_FDP4EP \sw_rdat_REG[50] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n257), .Q(sw_rdat[50]));
Q_FDP4EP \sw_rdat_REG[51] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n262), .Q(sw_rdat[51]));
Q_FDP4EP \sw_rdat_REG[52] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n267), .Q(sw_rdat[52]));
Q_FDP4EP \sw_rdat_REG[53] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n272), .Q(sw_rdat[53]));
Q_FDP4EP \sw_rdat_REG[54] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n277), .Q(sw_rdat[54]));
Q_FDP4EP \sw_rdat_REG[55] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n282), .Q(sw_rdat[55]));
Q_FDP4EP \sw_rdat_REG[56] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n287), .Q(sw_rdat[56]));
Q_FDP4EP \sw_rdat_REG[57] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n292), .Q(sw_rdat[57]));
Q_FDP4EP \sw_rdat_REG[58] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n297), .Q(sw_rdat[58]));
Q_FDP4EP \sw_rdat_REG[59] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n302), .Q(sw_rdat[59]));
Q_FDP4EP \sw_rdat_REG[60] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n307), .Q(sw_rdat[60]));
Q_FDP4EP \sw_rdat_REG[61] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n312), .Q(sw_rdat[61]));
Q_FDP4EP \sw_rdat_REG[62] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n317), .Q(sw_rdat[62]));
Q_FDP4EP \sw_rdat_REG[63] ( .CK(clk), .CE(sw_cs), .R(n323), .D(n322), .Q(sw_rdat[63]));
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m1 "_zyixc_ctx_rdata_29 1 63 0 0 31"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_NON_CMM "1"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "mem_a 1 63 0 0 31"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "1"
// pragma CVASTRPROP MODULE HDLICE PROP_RANOFF TRUE
endmodule
