
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module apb_xactor ( psel, penable, paddr, pwdata, pwrite, clk, reset_n, prdata, 
	pready, pslverr);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output psel;
output penable;
output [19:0] paddr;
output [31:0] pwdata;
output pwrite;
input clk;
input reset_n;
input [31:0] prdata;
input pready;
input pslverr;
wire _zy_simnet_psel_0_w$;
wire _zy_simnet_penable_1_w$;
wire [0:19] _zy_simnet_paddr_2_w$;
wire [0:31] _zy_simnet_pwdata_3_w$;
wire _zy_simnet_pwrite_4_w$;
wire [95:0] _zyixc_port_0_0_s2hW;
wire [63:0] _zyixc_port_0_1_s2hW;
wire _zyM2L61_pbcMevClk4;
wire _zyM2L61_pbcReq4;
wire _zyM2L61_pbcBusy4;
wire _zyM2L61_pbcWait4;
wire _zyM2L94_pbcMevClk9;
wire _zyM2L94_pbcReq9;
wire _zyM2L94_pbcBusy9;
wire _zyM2L94_pbcWait9;
wire _zzM2_bcBehEvalClk;
wire _zzM2_bcBehHalt;
wire _zzmdxOne;
wire _zzM2L46_mdxP0_EnNxt;
wire _zzM2L46_mdxP0_On;
wire _zzM2L61_mdxP1_EnNxt;
wire _zzM2L61_mdxP1_On;
wire _zzM2L94_mdxP2_EnNxt;
wire _zzM2L94_mdxP2_On;
wire [7:0] bus_timer;
`_2_ wire [7:0] _zyixc_port_0_0_h2s;
`_2_ wire [95:0] _zyixc_port_0_0_s2h;
`_2_ wire _zyixc_port_0_0_req;
`_2_ wire _zyixc_port_0_0_ack;
`_2_ wire _zyixc_port_0_0_isf;
`_2_ wire _zyixc_port_0_0_osf;
`_2_ wire [39:0] _zyixc_port_0_1_h2s;
`_2_ wire [63:0] _zyixc_port_0_1_s2h;
`_2_ wire _zyixc_port_0_1_req;
`_2_ wire _zyixc_port_0_1_ack;
`_2_ wire _zyixc_port_0_1_isf;
`_2_ wire _zyixc_port_0_1_osf;
wire [63:0] _zyaddr_L62_tfiV0_M2_pbcG0;
wire [31:0] _zydata_L63_tfiV1_M2_pbcG1;
wire _zyresponse_L64_tfiV2_M2_pbcG2;
wire [63:0] _zyaddr_L95_tfiV3_M2_pbcG3;
wire [31:0] _zydata_L96_tfiV4_M2_pbcG4;
wire _zyresponse_L97_tfiV5_M2_pbcG5;
wire _zyM2L61_pbcCapEn0;
wire _zyM2L73_pbcCapEn1;
wire _zyM2L79_pbcCapEn2;
wire _zyM2L90_pbcCapEn3;
wire _zyM2L94_pbcCapEn5;
wire _zyM2L104_pbcCapEn6;
wire _zyM2L110_pbcCapEn7;
wire _zyM2L121_pbcCapEn8;
wire [2:0] _zyM2L61_pbcFsm0_s;
wire _zyM2L61_pbcEn10;
wire [2:0] _zyM2L94_pbcFsm3_s;
wire _zyM2L94_pbcEn11;
wire [31:0] _zzM2_bcBehEval;
wire _zzM2L19_psel_mdxTmp0;
wire _zzM2L20_penable_mdxTmp1;
wire _zzM2L23_pwrite_mdxTmp2;
wire [19:0] _zzM2L21_paddr_mdxTmp3;
wire [31:0] _zzM2L22_pwdata_mdxTmp4;
wire [7:0] _zzM2L29_bus_timer_mdxTmp5;
wire _zzM2L46_mdxP0_En;
wire _zzM2L46_mdxP0_psel_wr0;
wire _zzM2L46_mdxP0_psel_Dwen0;
wire _zzM2L46_mdxP0_psel_DwenOn0;
wire _zzM2L46_mdxP0_penable_wr1;
wire _zzM2L46_mdxP0_penable_Dwen1;
wire _zzM2L46_mdxP0_penable_DwenOn1;
wire _zzM2L46_mdxP0_pwrite_wr2;
wire _zzM2L46_mdxP0_pwrite_Dwen2;
wire _zzM2L46_mdxP0_pwrite_DwenOn2;
wire [19:0] _zzM2L46_mdxP0_paddr_wr3;
wire _zzM2L46_mdxP0_paddr_Dwen3;
wire _zzM2L46_mdxP0_paddr_DwenOn3;
wire [31:0] _zzM2L46_mdxP0_pwdata_wr4;
wire _zzM2L46_mdxP0_pwdata_Dwen4;
wire _zzM2L46_mdxP0_pwdata_DwenOn4;
wire [7:0] _zzM2L46_mdxP0_bus_timer_wr5;
wire _zzM2L46_mdxP0_bus_timer_Dwen5;
wire _zzM2L46_mdxP0_bus_timer_DwenOn5;
wire _zzM2L61_mdxP1_En;
wire _zzM2L61_mdxP1_psel_wr0;
wire _zzM2L61_mdxP1_psel_Dwen0;
wire _zzM2L61_mdxP1_psel_DwenOn0;
wire _zzM2L61_mdxP1_penable_wr1;
wire _zzM2L61_mdxP1_penable_Dwen1;
wire _zzM2L61_mdxP1_penable_DwenOn1;
wire _zzM2L61_mdxP1_pwrite_wr2;
wire _zzM2L61_mdxP1_pwrite_Dwen2;
wire _zzM2L61_mdxP1_pwrite_DwenOn2;
wire [19:0] _zzM2L61_mdxP1_paddr_wr3;
wire _zzM2L61_mdxP1_paddr_Dwen3;
wire _zzM2L61_mdxP1_paddr_DwenOn3;
wire [31:0] _zzM2L61_mdxP1_pwdata_wr4;
wire _zzM2L61_mdxP1_pwdata_Dwen4;
wire _zzM2L61_mdxP1_pwdata_DwenOn4;
wire [7:0] _zzM2L61_mdxP1_bus_timer_wr5;
wire _zzM2L61_mdxP1_bus_timer_Dwen5;
wire _zzM2L61_mdxP1_bus_timer_DwenOn5;
wire _zzM2L94_mdxP2_En;
wire _zzM2L94_mdxP2_psel_wr0;
wire _zzM2L94_mdxP2_psel_Dwen0;
wire _zzM2L94_mdxP2_psel_DwenOn0;
wire _zzM2L94_mdxP2_penable_wr1;
wire _zzM2L94_mdxP2_penable_Dwen1;
wire _zzM2L94_mdxP2_penable_DwenOn1;
wire _zzM2L94_mdxP2_pwrite_wr2;
wire _zzM2L94_mdxP2_pwrite_Dwen2;
wire _zzM2L94_mdxP2_pwrite_DwenOn2;
wire [19:0] _zzM2L94_mdxP2_paddr_wr3;
wire _zzM2L94_mdxP2_paddr_Dwen3;
wire _zzM2L94_mdxP2_paddr_DwenOn3;
wire [7:0] _zzM2L94_mdxP2_bus_timer_wr4;
wire _zzM2L94_mdxP2_bus_timer_Dwen4;
wire _zzM2L94_mdxP2_bus_timer_DwenOn4;
wire _zzpsel_M2L19_mdxSvLt6;
wire _zzpenable_M2L20_mdxSvLt7;
wire _zzpwrite_M2L23_mdxSvLt8;
wire [19:0] _zzpaddr_M2L21_mdxSvLt9;
wire [31:0] _zzpwdata_M2L22_mdxSvLt10;
wire [7:0] _zzbus_timer_M2L29_mdxSvLt11;
supply1 n303;
supply0 n304;
supply0 n305;
supply0 n306;
supply0 n308;
supply0 n309;
supply0 n311;
supply0 n312;
supply0 n313;
supply0 n314;
Q_BUF U0 ( .A(n304), .Z(n1));
Q_AN02 U1 ( .A0(n27), .A1(n25), .Z(n2));
Q_OR02 U2 ( .A0(_zzM2L94_mdxP2_bus_timer_DwenOn4), .A1(_zzM2L61_mdxP1_bus_timer_DwenOn5), .Z(n3));
Q_INV U3 ( .A(_zzM2L46_mdxP0_bus_timer_DwenOn5), .Z(n5));
Q_NR02 U4 ( .A0(_zzM2L61_mdxP1_bus_timer_DwenOn5), .A1(n5), .Z(n6));
Q_OR02 U5 ( .A0(_zzM2L94_mdxP2_bus_timer_DwenOn4), .A1(n6), .Z(n4));
Q_LDP0 \bus_timer_REG[0] ( .G(_zzmdxOne), .D(_zzM2L29_bus_timer_mdxTmp5[0]), .Q(bus_timer[0]), .QN(n286));
Q_LDP0 \bus_timer_REG[1] ( .G(_zzmdxOne), .D(_zzM2L29_bus_timer_mdxTmp5[1]), .Q(bus_timer[1]), .QN( ));
Q_LDP0 \bus_timer_REG[2] ( .G(_zzmdxOne), .D(_zzM2L29_bus_timer_mdxTmp5[2]), .Q(bus_timer[2]), .QN(n294));
Q_LDP0 \bus_timer_REG[3] ( .G(_zzmdxOne), .D(_zzM2L29_bus_timer_mdxTmp5[3]), .Q(bus_timer[3]), .QN( ));
Q_LDP0 \bus_timer_REG[4] ( .G(_zzmdxOne), .D(_zzM2L29_bus_timer_mdxTmp5[4]), .Q(bus_timer[4]), .QN(n298));
Q_LDP0 \bus_timer_REG[5] ( .G(_zzmdxOne), .D(_zzM2L29_bus_timer_mdxTmp5[5]), .Q(bus_timer[5]), .QN(n299));
Q_LDP0 \bus_timer_REG[6] ( .G(_zzmdxOne), .D(_zzM2L29_bus_timer_mdxTmp5[6]), .Q(bus_timer[6]), .QN(n300));
Q_LDP0 \bus_timer_REG[7] ( .G(_zzmdxOne), .D(_zzM2L29_bus_timer_mdxTmp5[7]), .Q(bus_timer[7]), .QN(n301));
Q_MX04 U14 ( .S0(n4), .S1(n3), .A0(_zzbus_timer_M2L29_mdxSvLt11[7]), .A1(_zzM2L46_mdxP0_bus_timer_wr5[7]), .A2(_zzM2L61_mdxP1_bus_timer_wr5[7]), .A3(_zzM2L94_mdxP2_bus_timer_wr4[7]), .Z(_zzM2L29_bus_timer_mdxTmp5[7]));
Q_MX04 U15 ( .S0(n4), .S1(n3), .A0(_zzbus_timer_M2L29_mdxSvLt11[6]), .A1(_zzM2L46_mdxP0_bus_timer_wr5[6]), .A2(_zzM2L61_mdxP1_bus_timer_wr5[6]), .A3(_zzM2L94_mdxP2_bus_timer_wr4[6]), .Z(_zzM2L29_bus_timer_mdxTmp5[6]));
Q_MX04 U16 ( .S0(n4), .S1(n3), .A0(_zzbus_timer_M2L29_mdxSvLt11[5]), .A1(_zzM2L46_mdxP0_bus_timer_wr5[5]), .A2(_zzM2L61_mdxP1_bus_timer_wr5[5]), .A3(_zzM2L94_mdxP2_bus_timer_wr4[5]), .Z(_zzM2L29_bus_timer_mdxTmp5[5]));
Q_MX04 U17 ( .S0(n4), .S1(n3), .A0(_zzbus_timer_M2L29_mdxSvLt11[4]), .A1(_zzM2L46_mdxP0_bus_timer_wr5[4]), .A2(_zzM2L61_mdxP1_bus_timer_wr5[4]), .A3(_zzM2L94_mdxP2_bus_timer_wr4[4]), .Z(_zzM2L29_bus_timer_mdxTmp5[4]));
Q_MX04 U18 ( .S0(n4), .S1(n3), .A0(_zzbus_timer_M2L29_mdxSvLt11[3]), .A1(_zzM2L46_mdxP0_bus_timer_wr5[3]), .A2(_zzM2L61_mdxP1_bus_timer_wr5[3]), .A3(_zzM2L94_mdxP2_bus_timer_wr4[3]), .Z(_zzM2L29_bus_timer_mdxTmp5[3]));
Q_MX04 U19 ( .S0(n4), .S1(n3), .A0(_zzbus_timer_M2L29_mdxSvLt11[2]), .A1(_zzM2L46_mdxP0_bus_timer_wr5[2]), .A2(_zzM2L61_mdxP1_bus_timer_wr5[2]), .A3(_zzM2L94_mdxP2_bus_timer_wr4[2]), .Z(_zzM2L29_bus_timer_mdxTmp5[2]));
Q_MX04 U20 ( .S0(n4), .S1(n3), .A0(_zzbus_timer_M2L29_mdxSvLt11[1]), .A1(_zzM2L46_mdxP0_bus_timer_wr5[1]), .A2(_zzM2L61_mdxP1_bus_timer_wr5[1]), .A3(_zzM2L94_mdxP2_bus_timer_wr4[1]), .Z(_zzM2L29_bus_timer_mdxTmp5[1]));
Q_MX04 U21 ( .S0(n4), .S1(n3), .A0(_zzbus_timer_M2L29_mdxSvLt11[0]), .A1(_zzM2L46_mdxP0_bus_timer_wr5[0]), .A2(_zzM2L61_mdxP1_bus_timer_wr5[0]), .A3(_zzM2L94_mdxP2_bus_timer_wr4[0]), .Z(_zzM2L29_bus_timer_mdxTmp5[0]));
Q_AN02 U22 ( .A0(_zzM2L94_mdxP2_On), .A1(_zzM2L94_mdxP2_bus_timer_Dwen4), .Z(_zzM2L94_mdxP2_bus_timer_DwenOn4));
Q_AN02 U23 ( .A0(_zzM2L61_mdxP1_On), .A1(_zzM2L61_mdxP1_bus_timer_Dwen5), .Z(_zzM2L61_mdxP1_bus_timer_DwenOn5));
Q_AN02 U24 ( .A0(_zzM2L46_mdxP0_On), .A1(_zzM2L46_mdxP0_bus_timer_Dwen5), .Z(_zzM2L46_mdxP0_bus_timer_DwenOn5));
Q_INV U25 ( .A(_zzM2L61_mdxP1_pwdata_DwenOn4), .Z(n8));
Q_AN02 U26 ( .A0(_zzM2L46_mdxP0_pwdata_DwenOn4), .A1(n8), .Z(n7));
Q_LDP0 \pwdata_REG[0] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[0]), .Q(pwdata[0]), .QN( ));
Q_LDP0 \pwdata_REG[1] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[1]), .Q(pwdata[1]), .QN( ));
Q_LDP0 \pwdata_REG[2] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[2]), .Q(pwdata[2]), .QN( ));
Q_LDP0 \pwdata_REG[3] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[3]), .Q(pwdata[3]), .QN( ));
Q_LDP0 \pwdata_REG[4] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[4]), .Q(pwdata[4]), .QN( ));
Q_LDP0 \pwdata_REG[5] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[5]), .Q(pwdata[5]), .QN( ));
Q_LDP0 \pwdata_REG[6] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[6]), .Q(pwdata[6]), .QN( ));
Q_LDP0 \pwdata_REG[7] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[7]), .Q(pwdata[7]), .QN( ));
Q_LDP0 \pwdata_REG[8] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[8]), .Q(pwdata[8]), .QN( ));
Q_LDP0 \pwdata_REG[9] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[9]), .Q(pwdata[9]), .QN( ));
Q_LDP0 \pwdata_REG[10] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[10]), .Q(pwdata[10]), .QN( ));
Q_LDP0 \pwdata_REG[11] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[11]), .Q(pwdata[11]), .QN( ));
Q_LDP0 \pwdata_REG[12] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[12]), .Q(pwdata[12]), .QN( ));
Q_LDP0 \pwdata_REG[13] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[13]), .Q(pwdata[13]), .QN( ));
Q_LDP0 \pwdata_REG[14] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[14]), .Q(pwdata[14]), .QN( ));
Q_LDP0 \pwdata_REG[15] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[15]), .Q(pwdata[15]), .QN( ));
Q_LDP0 \pwdata_REG[16] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[16]), .Q(pwdata[16]), .QN( ));
Q_LDP0 \pwdata_REG[17] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[17]), .Q(pwdata[17]), .QN( ));
Q_LDP0 \pwdata_REG[18] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[18]), .Q(pwdata[18]), .QN( ));
Q_LDP0 \pwdata_REG[19] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[19]), .Q(pwdata[19]), .QN( ));
Q_LDP0 \pwdata_REG[20] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[20]), .Q(pwdata[20]), .QN( ));
Q_LDP0 \pwdata_REG[21] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[21]), .Q(pwdata[21]), .QN( ));
Q_LDP0 \pwdata_REG[22] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[22]), .Q(pwdata[22]), .QN( ));
Q_LDP0 \pwdata_REG[23] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[23]), .Q(pwdata[23]), .QN( ));
Q_LDP0 \pwdata_REG[24] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[24]), .Q(pwdata[24]), .QN( ));
Q_LDP0 \pwdata_REG[25] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[25]), .Q(pwdata[25]), .QN( ));
Q_LDP0 \pwdata_REG[26] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[26]), .Q(pwdata[26]), .QN( ));
Q_LDP0 \pwdata_REG[27] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[27]), .Q(pwdata[27]), .QN( ));
Q_LDP0 \pwdata_REG[28] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[28]), .Q(pwdata[28]), .QN( ));
Q_LDP0 \pwdata_REG[29] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[29]), .Q(pwdata[29]), .QN( ));
Q_LDP0 \pwdata_REG[30] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[30]), .Q(pwdata[30]), .QN( ));
Q_LDP0 \pwdata_REG[31] ( .G(_zzmdxOne), .D(_zzM2L22_pwdata_mdxTmp4[31]), .Q(pwdata[31]), .QN( ));
Q_MX03 U59 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[31]), .A1(_zzM2L46_mdxP0_pwdata_wr4[31]), .A2(_zzM2L61_mdxP1_pwdata_wr4[31]), .Z(_zzM2L22_pwdata_mdxTmp4[31]));
Q_MX03 U60 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[30]), .A1(_zzM2L46_mdxP0_pwdata_wr4[30]), .A2(_zzM2L61_mdxP1_pwdata_wr4[30]), .Z(_zzM2L22_pwdata_mdxTmp4[30]));
Q_MX03 U61 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[29]), .A1(_zzM2L46_mdxP0_pwdata_wr4[29]), .A2(_zzM2L61_mdxP1_pwdata_wr4[29]), .Z(_zzM2L22_pwdata_mdxTmp4[29]));
Q_MX03 U62 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[28]), .A1(_zzM2L46_mdxP0_pwdata_wr4[28]), .A2(_zzM2L61_mdxP1_pwdata_wr4[28]), .Z(_zzM2L22_pwdata_mdxTmp4[28]));
Q_MX03 U63 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[27]), .A1(_zzM2L46_mdxP0_pwdata_wr4[27]), .A2(_zzM2L61_mdxP1_pwdata_wr4[27]), .Z(_zzM2L22_pwdata_mdxTmp4[27]));
Q_MX03 U64 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[26]), .A1(_zzM2L46_mdxP0_pwdata_wr4[26]), .A2(_zzM2L61_mdxP1_pwdata_wr4[26]), .Z(_zzM2L22_pwdata_mdxTmp4[26]));
Q_MX03 U65 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[25]), .A1(_zzM2L46_mdxP0_pwdata_wr4[25]), .A2(_zzM2L61_mdxP1_pwdata_wr4[25]), .Z(_zzM2L22_pwdata_mdxTmp4[25]));
Q_MX03 U66 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[24]), .A1(_zzM2L46_mdxP0_pwdata_wr4[24]), .A2(_zzM2L61_mdxP1_pwdata_wr4[24]), .Z(_zzM2L22_pwdata_mdxTmp4[24]));
Q_MX03 U67 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[23]), .A1(_zzM2L46_mdxP0_pwdata_wr4[23]), .A2(_zzM2L61_mdxP1_pwdata_wr4[23]), .Z(_zzM2L22_pwdata_mdxTmp4[23]));
Q_MX03 U68 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[22]), .A1(_zzM2L46_mdxP0_pwdata_wr4[22]), .A2(_zzM2L61_mdxP1_pwdata_wr4[22]), .Z(_zzM2L22_pwdata_mdxTmp4[22]));
Q_MX03 U69 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[21]), .A1(_zzM2L46_mdxP0_pwdata_wr4[21]), .A2(_zzM2L61_mdxP1_pwdata_wr4[21]), .Z(_zzM2L22_pwdata_mdxTmp4[21]));
Q_MX03 U70 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[20]), .A1(_zzM2L46_mdxP0_pwdata_wr4[20]), .A2(_zzM2L61_mdxP1_pwdata_wr4[20]), .Z(_zzM2L22_pwdata_mdxTmp4[20]));
Q_MX03 U71 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[19]), .A1(_zzM2L46_mdxP0_pwdata_wr4[19]), .A2(_zzM2L61_mdxP1_pwdata_wr4[19]), .Z(_zzM2L22_pwdata_mdxTmp4[19]));
Q_MX03 U72 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[18]), .A1(_zzM2L46_mdxP0_pwdata_wr4[18]), .A2(_zzM2L61_mdxP1_pwdata_wr4[18]), .Z(_zzM2L22_pwdata_mdxTmp4[18]));
Q_MX03 U73 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[17]), .A1(_zzM2L46_mdxP0_pwdata_wr4[17]), .A2(_zzM2L61_mdxP1_pwdata_wr4[17]), .Z(_zzM2L22_pwdata_mdxTmp4[17]));
Q_MX03 U74 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[16]), .A1(_zzM2L46_mdxP0_pwdata_wr4[16]), .A2(_zzM2L61_mdxP1_pwdata_wr4[16]), .Z(_zzM2L22_pwdata_mdxTmp4[16]));
Q_MX03 U75 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[15]), .A1(_zzM2L46_mdxP0_pwdata_wr4[15]), .A2(_zzM2L61_mdxP1_pwdata_wr4[15]), .Z(_zzM2L22_pwdata_mdxTmp4[15]));
Q_MX03 U76 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[14]), .A1(_zzM2L46_mdxP0_pwdata_wr4[14]), .A2(_zzM2L61_mdxP1_pwdata_wr4[14]), .Z(_zzM2L22_pwdata_mdxTmp4[14]));
Q_MX03 U77 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[13]), .A1(_zzM2L46_mdxP0_pwdata_wr4[13]), .A2(_zzM2L61_mdxP1_pwdata_wr4[13]), .Z(_zzM2L22_pwdata_mdxTmp4[13]));
Q_MX03 U78 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[12]), .A1(_zzM2L46_mdxP0_pwdata_wr4[12]), .A2(_zzM2L61_mdxP1_pwdata_wr4[12]), .Z(_zzM2L22_pwdata_mdxTmp4[12]));
Q_MX03 U79 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[11]), .A1(_zzM2L46_mdxP0_pwdata_wr4[11]), .A2(_zzM2L61_mdxP1_pwdata_wr4[11]), .Z(_zzM2L22_pwdata_mdxTmp4[11]));
Q_MX03 U80 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[10]), .A1(_zzM2L46_mdxP0_pwdata_wr4[10]), .A2(_zzM2L61_mdxP1_pwdata_wr4[10]), .Z(_zzM2L22_pwdata_mdxTmp4[10]));
Q_MX03 U81 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[9]), .A1(_zzM2L46_mdxP0_pwdata_wr4[9]), .A2(_zzM2L61_mdxP1_pwdata_wr4[9]), .Z(_zzM2L22_pwdata_mdxTmp4[9]));
Q_MX03 U82 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[8]), .A1(_zzM2L46_mdxP0_pwdata_wr4[8]), .A2(_zzM2L61_mdxP1_pwdata_wr4[8]), .Z(_zzM2L22_pwdata_mdxTmp4[8]));
Q_MX03 U83 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[7]), .A1(_zzM2L46_mdxP0_pwdata_wr4[7]), .A2(_zzM2L61_mdxP1_pwdata_wr4[7]), .Z(_zzM2L22_pwdata_mdxTmp4[7]));
Q_MX03 U84 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[6]), .A1(_zzM2L46_mdxP0_pwdata_wr4[6]), .A2(_zzM2L61_mdxP1_pwdata_wr4[6]), .Z(_zzM2L22_pwdata_mdxTmp4[6]));
Q_MX03 U85 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[5]), .A1(_zzM2L46_mdxP0_pwdata_wr4[5]), .A2(_zzM2L61_mdxP1_pwdata_wr4[5]), .Z(_zzM2L22_pwdata_mdxTmp4[5]));
Q_MX03 U86 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[4]), .A1(_zzM2L46_mdxP0_pwdata_wr4[4]), .A2(_zzM2L61_mdxP1_pwdata_wr4[4]), .Z(_zzM2L22_pwdata_mdxTmp4[4]));
Q_MX03 U87 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[3]), .A1(_zzM2L46_mdxP0_pwdata_wr4[3]), .A2(_zzM2L61_mdxP1_pwdata_wr4[3]), .Z(_zzM2L22_pwdata_mdxTmp4[3]));
Q_MX03 U88 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[2]), .A1(_zzM2L46_mdxP0_pwdata_wr4[2]), .A2(_zzM2L61_mdxP1_pwdata_wr4[2]), .Z(_zzM2L22_pwdata_mdxTmp4[2]));
Q_MX03 U89 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[1]), .A1(_zzM2L46_mdxP0_pwdata_wr4[1]), .A2(_zzM2L61_mdxP1_pwdata_wr4[1]), .Z(_zzM2L22_pwdata_mdxTmp4[1]));
Q_MX03 U90 ( .S0(n7), .S1(_zzM2L61_mdxP1_pwdata_DwenOn4), .A0(_zzpwdata_M2L22_mdxSvLt10[0]), .A1(_zzM2L46_mdxP0_pwdata_wr4[0]), .A2(_zzM2L61_mdxP1_pwdata_wr4[0]), .Z(_zzM2L22_pwdata_mdxTmp4[0]));
Q_AN02 U91 ( .A0(_zzM2L61_mdxP1_On), .A1(_zzM2L61_mdxP1_pwdata_Dwen4), .Z(_zzM2L61_mdxP1_pwdata_DwenOn4));
Q_AN02 U92 ( .A0(_zzM2L46_mdxP0_On), .A1(_zzM2L46_mdxP0_pwdata_Dwen4), .Z(_zzM2L46_mdxP0_pwdata_DwenOn4));
Q_OR02 U93 ( .A0(_zzM2L94_mdxP2_paddr_DwenOn3), .A1(_zzM2L61_mdxP1_paddr_DwenOn3), .Z(n9));
Q_INV U94 ( .A(_zzM2L46_mdxP0_paddr_DwenOn3), .Z(n11));
Q_NR02 U95 ( .A0(_zzM2L61_mdxP1_paddr_DwenOn3), .A1(n11), .Z(n12));
Q_OR02 U96 ( .A0(_zzM2L94_mdxP2_paddr_DwenOn3), .A1(n12), .Z(n10));
Q_LDP0 \paddr_REG[0] ( .G(_zzmdxOne), .D(_zzM2L21_paddr_mdxTmp3[0]), .Q(paddr[0]), .QN( ));
Q_LDP0 \paddr_REG[1] ( .G(_zzmdxOne), .D(_zzM2L21_paddr_mdxTmp3[1]), .Q(paddr[1]), .QN( ));
Q_LDP0 \paddr_REG[2] ( .G(_zzmdxOne), .D(_zzM2L21_paddr_mdxTmp3[2]), .Q(paddr[2]), .QN( ));
Q_LDP0 \paddr_REG[3] ( .G(_zzmdxOne), .D(_zzM2L21_paddr_mdxTmp3[3]), .Q(paddr[3]), .QN( ));
Q_LDP0 \paddr_REG[4] ( .G(_zzmdxOne), .D(_zzM2L21_paddr_mdxTmp3[4]), .Q(paddr[4]), .QN( ));
Q_LDP0 \paddr_REG[5] ( .G(_zzmdxOne), .D(_zzM2L21_paddr_mdxTmp3[5]), .Q(paddr[5]), .QN( ));
Q_LDP0 \paddr_REG[6] ( .G(_zzmdxOne), .D(_zzM2L21_paddr_mdxTmp3[6]), .Q(paddr[6]), .QN( ));
Q_LDP0 \paddr_REG[7] ( .G(_zzmdxOne), .D(_zzM2L21_paddr_mdxTmp3[7]), .Q(paddr[7]), .QN( ));
Q_LDP0 \paddr_REG[8] ( .G(_zzmdxOne), .D(_zzM2L21_paddr_mdxTmp3[8]), .Q(paddr[8]), .QN( ));
Q_LDP0 \paddr_REG[9] ( .G(_zzmdxOne), .D(_zzM2L21_paddr_mdxTmp3[9]), .Q(paddr[9]), .QN( ));
Q_LDP0 \paddr_REG[10] ( .G(_zzmdxOne), .D(_zzM2L21_paddr_mdxTmp3[10]), .Q(paddr[10]), .QN( ));
Q_LDP0 \paddr_REG[11] ( .G(_zzmdxOne), .D(_zzM2L21_paddr_mdxTmp3[11]), .Q(paddr[11]), .QN( ));
Q_LDP0 \paddr_REG[12] ( .G(_zzmdxOne), .D(_zzM2L21_paddr_mdxTmp3[12]), .Q(paddr[12]), .QN( ));
Q_LDP0 \paddr_REG[13] ( .G(_zzmdxOne), .D(_zzM2L21_paddr_mdxTmp3[13]), .Q(paddr[13]), .QN( ));
Q_LDP0 \paddr_REG[14] ( .G(_zzmdxOne), .D(_zzM2L21_paddr_mdxTmp3[14]), .Q(paddr[14]), .QN( ));
Q_LDP0 \paddr_REG[15] ( .G(_zzmdxOne), .D(_zzM2L21_paddr_mdxTmp3[15]), .Q(paddr[15]), .QN( ));
Q_LDP0 \paddr_REG[16] ( .G(_zzmdxOne), .D(_zzM2L21_paddr_mdxTmp3[16]), .Q(paddr[16]), .QN( ));
Q_LDP0 \paddr_REG[17] ( .G(_zzmdxOne), .D(_zzM2L21_paddr_mdxTmp3[17]), .Q(paddr[17]), .QN( ));
Q_LDP0 \paddr_REG[18] ( .G(_zzmdxOne), .D(_zzM2L21_paddr_mdxTmp3[18]), .Q(paddr[18]), .QN( ));
Q_LDP0 \paddr_REG[19] ( .G(_zzmdxOne), .D(_zzM2L21_paddr_mdxTmp3[19]), .Q(paddr[19]), .QN( ));
Q_MX04 U117 ( .S0(n10), .S1(n9), .A0(_zzpaddr_M2L21_mdxSvLt9[19]), .A1(_zzM2L46_mdxP0_paddr_wr3[19]), .A2(_zzM2L61_mdxP1_paddr_wr3[19]), .A3(_zzM2L94_mdxP2_paddr_wr3[19]), .Z(_zzM2L21_paddr_mdxTmp3[19]));
Q_MX04 U118 ( .S0(n10), .S1(n9), .A0(_zzpaddr_M2L21_mdxSvLt9[18]), .A1(_zzM2L46_mdxP0_paddr_wr3[18]), .A2(_zzM2L61_mdxP1_paddr_wr3[18]), .A3(_zzM2L94_mdxP2_paddr_wr3[18]), .Z(_zzM2L21_paddr_mdxTmp3[18]));
Q_MX04 U119 ( .S0(n10), .S1(n9), .A0(_zzpaddr_M2L21_mdxSvLt9[17]), .A1(_zzM2L46_mdxP0_paddr_wr3[17]), .A2(_zzM2L61_mdxP1_paddr_wr3[17]), .A3(_zzM2L94_mdxP2_paddr_wr3[17]), .Z(_zzM2L21_paddr_mdxTmp3[17]));
Q_MX04 U120 ( .S0(n10), .S1(n9), .A0(_zzpaddr_M2L21_mdxSvLt9[16]), .A1(_zzM2L46_mdxP0_paddr_wr3[16]), .A2(_zzM2L61_mdxP1_paddr_wr3[16]), .A3(_zzM2L94_mdxP2_paddr_wr3[16]), .Z(_zzM2L21_paddr_mdxTmp3[16]));
Q_MX04 U121 ( .S0(n10), .S1(n9), .A0(_zzpaddr_M2L21_mdxSvLt9[15]), .A1(_zzM2L46_mdxP0_paddr_wr3[15]), .A2(_zzM2L61_mdxP1_paddr_wr3[15]), .A3(_zzM2L94_mdxP2_paddr_wr3[15]), .Z(_zzM2L21_paddr_mdxTmp3[15]));
Q_MX04 U122 ( .S0(n10), .S1(n9), .A0(_zzpaddr_M2L21_mdxSvLt9[14]), .A1(_zzM2L46_mdxP0_paddr_wr3[14]), .A2(_zzM2L61_mdxP1_paddr_wr3[14]), .A3(_zzM2L94_mdxP2_paddr_wr3[14]), .Z(_zzM2L21_paddr_mdxTmp3[14]));
Q_MX04 U123 ( .S0(n10), .S1(n9), .A0(_zzpaddr_M2L21_mdxSvLt9[13]), .A1(_zzM2L46_mdxP0_paddr_wr3[13]), .A2(_zzM2L61_mdxP1_paddr_wr3[13]), .A3(_zzM2L94_mdxP2_paddr_wr3[13]), .Z(_zzM2L21_paddr_mdxTmp3[13]));
Q_MX04 U124 ( .S0(n10), .S1(n9), .A0(_zzpaddr_M2L21_mdxSvLt9[12]), .A1(_zzM2L46_mdxP0_paddr_wr3[12]), .A2(_zzM2L61_mdxP1_paddr_wr3[12]), .A3(_zzM2L94_mdxP2_paddr_wr3[12]), .Z(_zzM2L21_paddr_mdxTmp3[12]));
Q_MX04 U125 ( .S0(n10), .S1(n9), .A0(_zzpaddr_M2L21_mdxSvLt9[11]), .A1(_zzM2L46_mdxP0_paddr_wr3[11]), .A2(_zzM2L61_mdxP1_paddr_wr3[11]), .A3(_zzM2L94_mdxP2_paddr_wr3[11]), .Z(_zzM2L21_paddr_mdxTmp3[11]));
Q_MX04 U126 ( .S0(n10), .S1(n9), .A0(_zzpaddr_M2L21_mdxSvLt9[10]), .A1(_zzM2L46_mdxP0_paddr_wr3[10]), .A2(_zzM2L61_mdxP1_paddr_wr3[10]), .A3(_zzM2L94_mdxP2_paddr_wr3[10]), .Z(_zzM2L21_paddr_mdxTmp3[10]));
Q_MX04 U127 ( .S0(n10), .S1(n9), .A0(_zzpaddr_M2L21_mdxSvLt9[9]), .A1(_zzM2L46_mdxP0_paddr_wr3[9]), .A2(_zzM2L61_mdxP1_paddr_wr3[9]), .A3(_zzM2L94_mdxP2_paddr_wr3[9]), .Z(_zzM2L21_paddr_mdxTmp3[9]));
Q_MX04 U128 ( .S0(n10), .S1(n9), .A0(_zzpaddr_M2L21_mdxSvLt9[8]), .A1(_zzM2L46_mdxP0_paddr_wr3[8]), .A2(_zzM2L61_mdxP1_paddr_wr3[8]), .A3(_zzM2L94_mdxP2_paddr_wr3[8]), .Z(_zzM2L21_paddr_mdxTmp3[8]));
Q_MX04 U129 ( .S0(n10), .S1(n9), .A0(_zzpaddr_M2L21_mdxSvLt9[7]), .A1(_zzM2L46_mdxP0_paddr_wr3[7]), .A2(_zzM2L61_mdxP1_paddr_wr3[7]), .A3(_zzM2L94_mdxP2_paddr_wr3[7]), .Z(_zzM2L21_paddr_mdxTmp3[7]));
Q_MX04 U130 ( .S0(n10), .S1(n9), .A0(_zzpaddr_M2L21_mdxSvLt9[6]), .A1(_zzM2L46_mdxP0_paddr_wr3[6]), .A2(_zzM2L61_mdxP1_paddr_wr3[6]), .A3(_zzM2L94_mdxP2_paddr_wr3[6]), .Z(_zzM2L21_paddr_mdxTmp3[6]));
Q_MX04 U131 ( .S0(n10), .S1(n9), .A0(_zzpaddr_M2L21_mdxSvLt9[5]), .A1(_zzM2L46_mdxP0_paddr_wr3[5]), .A2(_zzM2L61_mdxP1_paddr_wr3[5]), .A3(_zzM2L94_mdxP2_paddr_wr3[5]), .Z(_zzM2L21_paddr_mdxTmp3[5]));
Q_MX04 U132 ( .S0(n10), .S1(n9), .A0(_zzpaddr_M2L21_mdxSvLt9[4]), .A1(_zzM2L46_mdxP0_paddr_wr3[4]), .A2(_zzM2L61_mdxP1_paddr_wr3[4]), .A3(_zzM2L94_mdxP2_paddr_wr3[4]), .Z(_zzM2L21_paddr_mdxTmp3[4]));
Q_MX04 U133 ( .S0(n10), .S1(n9), .A0(_zzpaddr_M2L21_mdxSvLt9[3]), .A1(_zzM2L46_mdxP0_paddr_wr3[3]), .A2(_zzM2L61_mdxP1_paddr_wr3[3]), .A3(_zzM2L94_mdxP2_paddr_wr3[3]), .Z(_zzM2L21_paddr_mdxTmp3[3]));
Q_MX04 U134 ( .S0(n10), .S1(n9), .A0(_zzpaddr_M2L21_mdxSvLt9[2]), .A1(_zzM2L46_mdxP0_paddr_wr3[2]), .A2(_zzM2L61_mdxP1_paddr_wr3[2]), .A3(_zzM2L94_mdxP2_paddr_wr3[2]), .Z(_zzM2L21_paddr_mdxTmp3[2]));
Q_MX04 U135 ( .S0(n10), .S1(n9), .A0(_zzpaddr_M2L21_mdxSvLt9[1]), .A1(_zzM2L46_mdxP0_paddr_wr3[1]), .A2(_zzM2L61_mdxP1_paddr_wr3[1]), .A3(_zzM2L94_mdxP2_paddr_wr3[1]), .Z(_zzM2L21_paddr_mdxTmp3[1]));
Q_MX04 U136 ( .S0(n10), .S1(n9), .A0(_zzpaddr_M2L21_mdxSvLt9[0]), .A1(_zzM2L46_mdxP0_paddr_wr3[0]), .A2(_zzM2L61_mdxP1_paddr_wr3[0]), .A3(_zzM2L94_mdxP2_paddr_wr3[0]), .Z(_zzM2L21_paddr_mdxTmp3[0]));
Q_AN02 U137 ( .A0(_zzM2L94_mdxP2_On), .A1(_zzM2L94_mdxP2_paddr_Dwen3), .Z(_zzM2L94_mdxP2_paddr_DwenOn3));
Q_AN02 U138 ( .A0(_zzM2L61_mdxP1_On), .A1(_zzM2L61_mdxP1_paddr_Dwen3), .Z(_zzM2L61_mdxP1_paddr_DwenOn3));
Q_AN02 U139 ( .A0(_zzM2L46_mdxP0_On), .A1(_zzM2L46_mdxP0_paddr_Dwen3), .Z(_zzM2L46_mdxP0_paddr_DwenOn3));
Q_OR02 U140 ( .A0(_zzM2L94_mdxP2_pwrite_DwenOn2), .A1(_zzM2L61_mdxP1_pwrite_DwenOn2), .Z(n13));
Q_INV U141 ( .A(_zzM2L46_mdxP0_pwrite_DwenOn2), .Z(n15));
Q_NR02 U142 ( .A0(_zzM2L61_mdxP1_pwrite_DwenOn2), .A1(n15), .Z(n16));
Q_OR02 U143 ( .A0(_zzM2L94_mdxP2_pwrite_DwenOn2), .A1(n16), .Z(n14));
Q_LDP0 pwrite_REG  ( .G(_zzmdxOne), .D(_zzM2L23_pwrite_mdxTmp2), .Q(pwrite), .QN( ));
Q_MX04 U145 ( .S0(n14), .S1(n13), .A0(_zzpwrite_M2L23_mdxSvLt8), .A1(_zzM2L46_mdxP0_pwrite_wr2), .A2(_zzM2L61_mdxP1_pwrite_wr2), .A3(_zzM2L94_mdxP2_pwrite_wr2), .Z(_zzM2L23_pwrite_mdxTmp2));
Q_AN02 U146 ( .A0(_zzM2L94_mdxP2_On), .A1(_zzM2L94_mdxP2_pwrite_Dwen2), .Z(_zzM2L94_mdxP2_pwrite_DwenOn2));
Q_AN02 U147 ( .A0(_zzM2L61_mdxP1_On), .A1(_zzM2L61_mdxP1_pwrite_Dwen2), .Z(_zzM2L61_mdxP1_pwrite_DwenOn2));
Q_AN02 U148 ( .A0(_zzM2L46_mdxP0_On), .A1(_zzM2L46_mdxP0_pwrite_Dwen2), .Z(_zzM2L46_mdxP0_pwrite_DwenOn2));
Q_OR02 U149 ( .A0(_zzM2L94_mdxP2_penable_DwenOn1), .A1(_zzM2L61_mdxP1_penable_DwenOn1), .Z(n17));
Q_INV U150 ( .A(_zzM2L46_mdxP0_penable_DwenOn1), .Z(n19));
Q_NR02 U151 ( .A0(_zzM2L61_mdxP1_penable_DwenOn1), .A1(n19), .Z(n20));
Q_OR02 U152 ( .A0(_zzM2L94_mdxP2_penable_DwenOn1), .A1(n20), .Z(n18));
Q_LDP0 penable_REG  ( .G(_zzmdxOne), .D(_zzM2L20_penable_mdxTmp1), .Q(penable), .QN( ));
Q_MX04 U154 ( .S0(n18), .S1(n17), .A0(_zzpenable_M2L20_mdxSvLt7), .A1(_zzM2L46_mdxP0_penable_wr1), .A2(_zzM2L61_mdxP1_penable_wr1), .A3(_zzM2L94_mdxP2_penable_wr1), .Z(_zzM2L20_penable_mdxTmp1));
Q_AN02 U155 ( .A0(_zzM2L94_mdxP2_On), .A1(_zzM2L94_mdxP2_penable_Dwen1), .Z(_zzM2L94_mdxP2_penable_DwenOn1));
Q_AN02 U156 ( .A0(_zzM2L61_mdxP1_On), .A1(_zzM2L61_mdxP1_penable_Dwen1), .Z(_zzM2L61_mdxP1_penable_DwenOn1));
Q_AN02 U157 ( .A0(_zzM2L46_mdxP0_On), .A1(_zzM2L46_mdxP0_penable_Dwen1), .Z(_zzM2L46_mdxP0_penable_DwenOn1));
Q_OR02 U158 ( .A0(_zzM2L94_mdxP2_psel_DwenOn0), .A1(_zzM2L61_mdxP1_psel_DwenOn0), .Z(n21));
Q_INV U159 ( .A(_zzM2L46_mdxP0_psel_DwenOn0), .Z(n23));
Q_NR02 U160 ( .A0(_zzM2L61_mdxP1_psel_DwenOn0), .A1(n23), .Z(n24));
Q_OR02 U161 ( .A0(_zzM2L94_mdxP2_psel_DwenOn0), .A1(n24), .Z(n22));
Q_LDP0 psel_REG  ( .G(_zzmdxOne), .D(_zzM2L19_psel_mdxTmp0), .Q(psel), .QN( ));
Q_MX04 U163 ( .S0(n22), .S1(n21), .A0(_zzpsel_M2L19_mdxSvLt6), .A1(_zzM2L46_mdxP0_psel_wr0), .A2(_zzM2L61_mdxP1_psel_wr0), .A3(_zzM2L94_mdxP2_psel_wr0), .Z(_zzM2L19_psel_mdxTmp0));
Q_AN02 U164 ( .A0(_zzM2L94_mdxP2_On), .A1(_zzM2L94_mdxP2_psel_Dwen0), .Z(_zzM2L94_mdxP2_psel_DwenOn0));
Q_AN02 U165 ( .A0(_zzM2L61_mdxP1_On), .A1(_zzM2L61_mdxP1_psel_Dwen0), .Z(_zzM2L61_mdxP1_psel_DwenOn0));
Q_AN02 U166 ( .A0(_zzM2L46_mdxP0_On), .A1(_zzM2L46_mdxP0_psel_Dwen0), .Z(_zzM2L46_mdxP0_psel_DwenOn0));
Q_AN02 U167 ( .A0(n26), .A1(n85), .Z(n25));
Q_AD01HF U168 ( .A0(_zzM2_bcBehEval[29]), .B0(n29), .S(n28), .CO(n27));
Q_AD01HF U169 ( .A0(_zzM2_bcBehEval[28]), .B0(n31), .S(n30), .CO(n29));
Q_AD01HF U170 ( .A0(_zzM2_bcBehEval[27]), .B0(n33), .S(n32), .CO(n31));
Q_AD01HF U171 ( .A0(_zzM2_bcBehEval[26]), .B0(n35), .S(n34), .CO(n33));
Q_AD01HF U172 ( .A0(_zzM2_bcBehEval[25]), .B0(n37), .S(n36), .CO(n35));
Q_AD01HF U173 ( .A0(_zzM2_bcBehEval[24]), .B0(n39), .S(n38), .CO(n37));
Q_AD01HF U174 ( .A0(_zzM2_bcBehEval[23]), .B0(n41), .S(n40), .CO(n39));
Q_AD01HF U175 ( .A0(_zzM2_bcBehEval[22]), .B0(n43), .S(n42), .CO(n41));
Q_AD01HF U176 ( .A0(_zzM2_bcBehEval[21]), .B0(n45), .S(n44), .CO(n43));
Q_AD01HF U177 ( .A0(_zzM2_bcBehEval[20]), .B0(n47), .S(n46), .CO(n45));
Q_AD01HF U178 ( .A0(_zzM2_bcBehEval[19]), .B0(n49), .S(n48), .CO(n47));
Q_AD01HF U179 ( .A0(_zzM2_bcBehEval[18]), .B0(n51), .S(n50), .CO(n49));
Q_AD01HF U180 ( .A0(_zzM2_bcBehEval[17]), .B0(n53), .S(n52), .CO(n51));
Q_AD01HF U181 ( .A0(_zzM2_bcBehEval[16]), .B0(n55), .S(n54), .CO(n53));
Q_AD01HF U182 ( .A0(_zzM2_bcBehEval[15]), .B0(n57), .S(n56), .CO(n55));
Q_AD01HF U183 ( .A0(_zzM2_bcBehEval[14]), .B0(n59), .S(n58), .CO(n57));
Q_AD01HF U184 ( .A0(_zzM2_bcBehEval[13]), .B0(n61), .S(n60), .CO(n59));
Q_AD01HF U185 ( .A0(_zzM2_bcBehEval[12]), .B0(n63), .S(n62), .CO(n61));
Q_AD01HF U186 ( .A0(_zzM2_bcBehEval[11]), .B0(n65), .S(n64), .CO(n63));
Q_AD01HF U187 ( .A0(_zzM2_bcBehEval[10]), .B0(n67), .S(n66), .CO(n65));
Q_AD01HF U188 ( .A0(_zzM2_bcBehEval[9]), .B0(n69), .S(n68), .CO(n67));
Q_AD01HF U189 ( .A0(_zzM2_bcBehEval[8]), .B0(n71), .S(n70), .CO(n69));
Q_AD01HF U190 ( .A0(_zzM2_bcBehEval[7]), .B0(n73), .S(n72), .CO(n71));
Q_AD01HF U191 ( .A0(_zzM2_bcBehEval[6]), .B0(n75), .S(n74), .CO(n73));
Q_AD01HF U192 ( .A0(_zzM2_bcBehEval[5]), .B0(n77), .S(n76), .CO(n75));
Q_AD01HF U193 ( .A0(_zzM2_bcBehEval[4]), .B0(n79), .S(n78), .CO(n77));
Q_AD01HF U194 ( .A0(_zzM2_bcBehEval[3]), .B0(n81), .S(n80), .CO(n79));
Q_AD01HF U195 ( .A0(_zzM2_bcBehEval[2]), .B0(n83), .S(n82), .CO(n81));
Q_AD01HF U196 ( .A0(_zzM2_bcBehEval[1]), .B0(_zzM2_bcBehEval[0]), .S(n84), .CO(n83));
Q_OR02 U197 ( .A0(_zyM2L61_pbcWait4), .A1(_zyM2L94_pbcWait9), .Z(n26));
Q_ND03 U198 ( .A0(n88), .A1(n87), .A2(n86), .Z(n85));
Q_AN03 U199 ( .A0(n91), .A1(n90), .A2(n89), .Z(n86));
Q_AN03 U200 ( .A0(n94), .A1(n93), .A2(n92), .Z(n87));
Q_AN03 U201 ( .A0(n97), .A1(n96), .A2(n95), .Z(n88));
Q_AN03 U202 ( .A0(_zzM2_bcBehEval[0]), .A1(n99), .A2(n98), .Z(n89));
Q_AN03 U203 ( .A0(_zzM2_bcBehEval[3]), .A1(_zzM2_bcBehEval[2]), .A2(_zzM2_bcBehEval[1]), .Z(n90));
Q_AN03 U204 ( .A0(_zzM2_bcBehEval[6]), .A1(_zzM2_bcBehEval[5]), .A2(_zzM2_bcBehEval[4]), .Z(n91));
Q_AN03 U205 ( .A0(_zzM2_bcBehEval[9]), .A1(_zzM2_bcBehEval[8]), .A2(_zzM2_bcBehEval[7]), .Z(n92));
Q_AN03 U206 ( .A0(_zzM2_bcBehEval[12]), .A1(_zzM2_bcBehEval[11]), .A2(_zzM2_bcBehEval[10]), .Z(n93));
Q_AN03 U207 ( .A0(_zzM2_bcBehEval[15]), .A1(_zzM2_bcBehEval[14]), .A2(_zzM2_bcBehEval[13]), .Z(n94));
Q_AN03 U208 ( .A0(_zzM2_bcBehEval[18]), .A1(_zzM2_bcBehEval[17]), .A2(_zzM2_bcBehEval[16]), .Z(n95));
Q_AN03 U209 ( .A0(_zzM2_bcBehEval[21]), .A1(_zzM2_bcBehEval[20]), .A2(_zzM2_bcBehEval[19]), .Z(n96));
Q_AN03 U210 ( .A0(_zzM2_bcBehEval[24]), .A1(_zzM2_bcBehEval[23]), .A2(_zzM2_bcBehEval[22]), .Z(n97));
Q_AN03 U211 ( .A0(_zzM2_bcBehEval[27]), .A1(_zzM2_bcBehEval[26]), .A2(_zzM2_bcBehEval[25]), .Z(n98));
Q_AN03 U212 ( .A0(_zzM2_bcBehEval[30]), .A1(_zzM2_bcBehEval[29]), .A2(_zzM2_bcBehEval[28]), .Z(n99));
Q_AO21 U213 ( .A0(n127), .A1(_zyM2L94_pbcFsm3_s[0]), .B0(n125), .Z(n131));
Q_AN02 U214 ( .A0(_zyM2L94_pbcFsm3_s[1]), .A1(n108), .Z(n125));
Q_AN02 U215 ( .A0(n101), .A1(n131), .Z(n117));
Q_OR02 U216 ( .A0(_zyM2L94_pbcFsm3_s[1]), .A1(_zyM2L94_pbcFsm3_s[0]), .Z(n107));
Q_INV U217 ( .A(pready), .Z(n124));
Q_AN02 U218 ( .A0(n124), .A1(n100), .Z(n132));
Q_AO21 U219 ( .A0(n107), .A1(n132), .B0(n122), .Z(n133));
Q_AN02 U220 ( .A0(_zyM2L94_pbcFsm3_s[1]), .A1(_zyM2L94_pbcFsm3_s[0]), .Z(n122));
Q_OR02 U221 ( .A0(n133), .A1(_zyM2L94_pbcFsm3_s[2]), .Z(n119));
Q_INV U222 ( .A(n119), .Z(n115));
Q_OA21 U223 ( .A0(n132), .A1(_zyM2L94_pbcFsm3_s[0]), .B0(_zyM2L94_pbcFsm3_s[1]), .Z(n120));
Q_OR02 U224 ( .A0(n120), .A1(_zyM2L94_pbcFsm3_s[2]), .Z(n121));
Q_INV U225 ( .A(n121), .Z(n113));
Q_OR02 U226 ( .A0(n122), .A1(_zyM2L94_pbcFsm3_s[2]), .Z(n129));
Q_INV U227 ( .A(n122), .Z(n109));
Q_INV U228 ( .A(n107), .Z(n114));
Q_AO21 U229 ( .A0(n109), .A1(n132), .B0(n114), .Z(n111));
Q_OR02 U230 ( .A0(n111), .A1(_zyM2L94_pbcFsm3_s[2]), .Z(n123));
Q_AN03 U231 ( .A0(_zyM2L94_pbcFsm3_s[0]), .A1(n124), .A2(n100), .Z(n112));
Q_AO21 U232 ( .A0(n127), .A1(n112), .B0(n125), .Z(n126));
Q_AN02 U233 ( .A0(n101), .A1(n126), .Z(n102));
Q_AN02 U234 ( .A0(n101), .A1(n127), .Z(n103));
Q_INV U235 ( .A(n131), .Z(n128));
Q_AN02 U236 ( .A0(n101), .A1(n128), .Z(n104));
Q_OR03 U237 ( .A0(n114), .A1(n132), .A2(n129), .Z(n130));
Q_AN03 U238 ( .A0(n101), .A1(_zyM2L94_pbcFsm3_s[1]), .A2(_zyM2L94_pbcFsm3_s[0]), .Z(n105));
Q_AN02 U239 ( .A0(n103), .A1(n108), .Z(n106));
Q_AN02 U240 ( .A0(n132), .A1(n131), .Z(n116));
Q_INV U241 ( .A(n133), .Z(n110));
Q_INV U242 ( .A(n116), .Z(n118));
Q_FDP0 _zzM2L94_mdxP2_bus_timer_Dwen4_REG  ( .CK(_zyM2L94_pbcMevClk9), .D(n117), .Q(_zzM2L94_mdxP2_bus_timer_Dwen4), .QN( ));
Q_FDP0 _zzM2L94_mdxP2_paddr_Dwen3_REG  ( .CK(_zyM2L94_pbcMevClk9), .D(n115), .Q(_zzM2L94_mdxP2_paddr_Dwen3), .QN( ));
Q_FDP0 _zzM2L94_mdxP2_pwrite_Dwen2_REG  ( .CK(_zyM2L94_pbcMevClk9), .D(n115), .Q(_zzM2L94_mdxP2_pwrite_Dwen2), .QN( ));
Q_FDP0 _zzM2L94_mdxP2_penable_Dwen1_REG  ( .CK(_zyM2L94_pbcMevClk9), .D(n113), .Q(_zzM2L94_mdxP2_penable_Dwen1), .QN( ));
Q_FDP0 _zzM2L94_mdxP2_psel_Dwen0_REG  ( .CK(_zyM2L94_pbcMevClk9), .D(n115), .Q(_zzM2L94_mdxP2_psel_Dwen0), .QN( ));
Q_FDP0 \_zyM2L94_pbcFsm3_s_REG[2] ( .CK(_zyM2L94_pbcMevClk9), .D(_zyM2L94_pbcFsm3_s[2]), .Q(_zyM2L94_pbcFsm3_s[2]), .QN(n101));
Q_XNR2 U249 ( .A0(n111), .A1(n133), .Z(n134));
Q_AN02 U250 ( .A0(n114), .A1(_zyixc_port_0_1_s2h[19]), .Z(n135));
Q_AN02 U251 ( .A0(n114), .A1(_zyixc_port_0_1_s2h[18]), .Z(n136));
Q_AN02 U252 ( .A0(n114), .A1(_zyixc_port_0_1_s2h[17]), .Z(n137));
Q_AN02 U253 ( .A0(n114), .A1(_zyixc_port_0_1_s2h[16]), .Z(n138));
Q_AN02 U254 ( .A0(n114), .A1(_zyixc_port_0_1_s2h[15]), .Z(n139));
Q_AN02 U255 ( .A0(n114), .A1(_zyixc_port_0_1_s2h[14]), .Z(n140));
Q_AN02 U256 ( .A0(n114), .A1(_zyixc_port_0_1_s2h[13]), .Z(n141));
Q_AN02 U257 ( .A0(n114), .A1(_zyixc_port_0_1_s2h[12]), .Z(n142));
Q_AN02 U258 ( .A0(n114), .A1(_zyixc_port_0_1_s2h[11]), .Z(n143));
Q_AN02 U259 ( .A0(n114), .A1(_zyixc_port_0_1_s2h[10]), .Z(n144));
Q_AN02 U260 ( .A0(n114), .A1(_zyixc_port_0_1_s2h[9]), .Z(n145));
Q_AN02 U261 ( .A0(n114), .A1(_zyixc_port_0_1_s2h[8]), .Z(n146));
Q_AN02 U262 ( .A0(n114), .A1(_zyixc_port_0_1_s2h[7]), .Z(n147));
Q_AN02 U263 ( .A0(n114), .A1(_zyixc_port_0_1_s2h[6]), .Z(n148));
Q_AN02 U264 ( .A0(n114), .A1(_zyixc_port_0_1_s2h[5]), .Z(n149));
Q_AN02 U265 ( .A0(n114), .A1(_zyixc_port_0_1_s2h[4]), .Z(n150));
Q_AN02 U266 ( .A0(n114), .A1(_zyixc_port_0_1_s2h[3]), .Z(n151));
Q_AN02 U267 ( .A0(n114), .A1(_zyixc_port_0_1_s2h[2]), .Z(n152));
Q_AN02 U268 ( .A0(n114), .A1(_zyixc_port_0_1_s2h[1]), .Z(n153));
Q_AN02 U269 ( .A0(n114), .A1(_zyixc_port_0_1_s2h[0]), .Z(n154));
Q_AN02 U270 ( .A0(n116), .A1(n163), .Z(n155));
Q_AN02 U271 ( .A0(n116), .A1(n165), .Z(n156));
Q_AN02 U272 ( .A0(n116), .A1(n167), .Z(n157));
Q_AN02 U273 ( .A0(n116), .A1(n169), .Z(n158));
Q_AN02 U274 ( .A0(n116), .A1(n171), .Z(n159));
Q_AN02 U275 ( .A0(n116), .A1(n173), .Z(n160));
Q_AN02 U276 ( .A0(n116), .A1(n175), .Z(n161));
Q_AN02 U277 ( .A0(n116), .A1(n176), .Z(n162));
Q_XOR2 U278 ( .A0(bus_timer[7]), .A1(n164), .Z(n163));
Q_AD01HF U279 ( .A0(bus_timer[6]), .B0(n166), .S(n165), .CO(n164));
Q_AD01HF U280 ( .A0(bus_timer[5]), .B0(n168), .S(n167), .CO(n166));
Q_AD01HF U281 ( .A0(bus_timer[4]), .B0(n170), .S(n169), .CO(n168));
Q_AD01HF U282 ( .A0(bus_timer[3]), .B0(n172), .S(n171), .CO(n170));
Q_AD01HF U283 ( .A0(bus_timer[2]), .B0(n174), .S(n173), .CO(n172));
Q_AD01HF U284 ( .A0(bus_timer[1]), .B0(bus_timer[0]), .S(n175), .CO(n174));
Q_INV U285 ( .A(bus_timer[0]), .Z(n176));
Q_OR02 U286 ( .A0(pslverr), .A1(n178), .Z(n177));
Q_NR02 U287 ( .A0(n180), .A1(n179), .Z(n178));
Q_OR03 U288 ( .A0(bus_timer[1]), .A1(bus_timer[0]), .A2(n181), .Z(n179));
Q_OR03 U289 ( .A0(bus_timer[4]), .A1(bus_timer[3]), .A2(n184), .Z(n180));
Q_OR03 U290 ( .A0(bus_timer[7]), .A1(n182), .A2(n183), .Z(n181));
Q_INV U291 ( .A(bus_timer[6]), .Z(n182));
Q_INV U292 ( .A(bus_timer[5]), .Z(n183));
Q_INV U293 ( .A(bus_timer[2]), .Z(n184));
Q_AO21 U294 ( .A0(n186), .A1(n185), .B0(n187), .Z(n100));
Q_NR02 U295 ( .A0(bus_timer[3]), .A1(bus_timer[2]), .Z(n185));
Q_AN02 U296 ( .A0(n191), .A1(n188), .Z(n186));
Q_OA21 U297 ( .A0(n190), .A1(n189), .B0(n191), .Z(n187));
Q_INV U298 ( .A(bus_timer[4]), .Z(n188));
Q_INV U299 ( .A(bus_timer[5]), .Z(n189));
Q_INV U300 ( .A(bus_timer[6]), .Z(n190));
Q_INV U301 ( .A(bus_timer[7]), .Z(n191));
Q_AO21 U302 ( .A0(n218), .A1(_zyM2L61_pbcFsm0_s[0]), .B0(n216), .Z(n222));
Q_AN02 U303 ( .A0(_zyM2L61_pbcFsm0_s[1]), .A1(n200), .Z(n216));
Q_AN02 U304 ( .A0(n193), .A1(n222), .Z(n209));
Q_OR02 U305 ( .A0(_zyM2L61_pbcFsm0_s[1]), .A1(_zyM2L61_pbcFsm0_s[0]), .Z(n199));
Q_AN02 U306 ( .A0(n124), .A1(n192), .Z(n223));
Q_AO21 U307 ( .A0(n199), .A1(n223), .B0(n214), .Z(n224));
Q_AN02 U308 ( .A0(_zyM2L61_pbcFsm0_s[1]), .A1(_zyM2L61_pbcFsm0_s[0]), .Z(n214));
Q_OR02 U309 ( .A0(n224), .A1(_zyM2L61_pbcFsm0_s[2]), .Z(n211));
Q_INV U310 ( .A(n211), .Z(n207));
Q_OA21 U311 ( .A0(n223), .A1(_zyM2L61_pbcFsm0_s[0]), .B0(_zyM2L61_pbcFsm0_s[1]), .Z(n212));
Q_OR02 U312 ( .A0(n212), .A1(_zyM2L61_pbcFsm0_s[2]), .Z(n213));
Q_INV U313 ( .A(n213), .Z(n205));
Q_OR02 U314 ( .A0(n214), .A1(_zyM2L61_pbcFsm0_s[2]), .Z(n220));
Q_INV U315 ( .A(n214), .Z(n201));
Q_INV U316 ( .A(n199), .Z(n206));
Q_AO21 U317 ( .A0(n201), .A1(n223), .B0(n206), .Z(n203));
Q_OR02 U318 ( .A0(n203), .A1(_zyM2L61_pbcFsm0_s[2]), .Z(n215));
Q_AN03 U319 ( .A0(_zyM2L61_pbcFsm0_s[0]), .A1(n124), .A2(n192), .Z(n204));
Q_AO21 U320 ( .A0(n218), .A1(n204), .B0(n216), .Z(n217));
Q_AN02 U321 ( .A0(n193), .A1(n217), .Z(n194));
Q_AN02 U322 ( .A0(n193), .A1(n218), .Z(n195));
Q_INV U323 ( .A(n222), .Z(n219));
Q_AN02 U324 ( .A0(n193), .A1(n219), .Z(n196));
Q_OR03 U325 ( .A0(n206), .A1(n223), .A2(n220), .Z(n221));
Q_AN03 U326 ( .A0(n193), .A1(_zyM2L61_pbcFsm0_s[1]), .A2(_zyM2L61_pbcFsm0_s[0]), .Z(n197));
Q_AN02 U327 ( .A0(n195), .A1(n200), .Z(n198));
Q_AN02 U328 ( .A0(n223), .A1(n222), .Z(n208));
Q_INV U329 ( .A(n224), .Z(n202));
Q_INV U330 ( .A(n208), .Z(n210));
Q_FDP0 _zzM2L61_mdxP1_bus_timer_Dwen5_REG  ( .CK(_zyM2L61_pbcMevClk4), .D(n209), .Q(_zzM2L61_mdxP1_bus_timer_Dwen5), .QN( ));
Q_FDP0 _zzM2L61_mdxP1_pwdata_Dwen4_REG  ( .CK(_zyM2L61_pbcMevClk4), .D(n207), .Q(_zzM2L61_mdxP1_pwdata_Dwen4), .QN( ));
Q_FDP0 _zzM2L61_mdxP1_paddr_Dwen3_REG  ( .CK(_zyM2L61_pbcMevClk4), .D(n207), .Q(_zzM2L61_mdxP1_paddr_Dwen3), .QN( ));
Q_FDP0 _zzM2L61_mdxP1_pwrite_Dwen2_REG  ( .CK(_zyM2L61_pbcMevClk4), .D(n207), .Q(_zzM2L61_mdxP1_pwrite_Dwen2), .QN( ));
Q_FDP0 _zzM2L61_mdxP1_penable_Dwen1_REG  ( .CK(_zyM2L61_pbcMevClk4), .D(n205), .Q(_zzM2L61_mdxP1_penable_Dwen1), .QN( ));
Q_FDP0 _zzM2L61_mdxP1_psel_Dwen0_REG  ( .CK(_zyM2L61_pbcMevClk4), .D(n207), .Q(_zzM2L61_mdxP1_psel_Dwen0), .QN( ));
Q_FDP0 \_zyM2L61_pbcFsm0_s_REG[2] ( .CK(_zyM2L61_pbcMevClk4), .D(_zyM2L61_pbcFsm0_s[2]), .Q(_zyM2L61_pbcFsm0_s[2]), .QN(n193));
Q_XNR2 U338 ( .A0(n203), .A1(n224), .Z(n225));
Q_AN02 U339 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[19]), .Z(n226));
Q_AN02 U340 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[18]), .Z(n227));
Q_AN02 U341 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[17]), .Z(n228));
Q_AN02 U342 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[16]), .Z(n229));
Q_AN02 U343 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[15]), .Z(n230));
Q_AN02 U344 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[14]), .Z(n231));
Q_AN02 U345 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[13]), .Z(n232));
Q_AN02 U346 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[12]), .Z(n233));
Q_AN02 U347 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[11]), .Z(n234));
Q_AN02 U348 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[10]), .Z(n235));
Q_AN02 U349 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[9]), .Z(n236));
Q_AN02 U350 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[8]), .Z(n237));
Q_AN02 U351 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[7]), .Z(n238));
Q_AN02 U352 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[6]), .Z(n239));
Q_AN02 U353 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[5]), .Z(n240));
Q_AN02 U354 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[4]), .Z(n241));
Q_AN02 U355 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[3]), .Z(n242));
Q_AN02 U356 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[2]), .Z(n243));
Q_AN02 U357 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[1]), .Z(n244));
Q_AN02 U358 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[0]), .Z(n245));
Q_AN02 U359 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[95]), .Z(n246));
Q_AN02 U360 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[94]), .Z(n247));
Q_AN02 U361 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[93]), .Z(n248));
Q_AN02 U362 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[92]), .Z(n249));
Q_AN02 U363 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[91]), .Z(n250));
Q_AN02 U364 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[90]), .Z(n251));
Q_AN02 U365 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[89]), .Z(n252));
Q_AN02 U366 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[88]), .Z(n253));
Q_AN02 U367 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[87]), .Z(n254));
Q_AN02 U368 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[86]), .Z(n255));
Q_AN02 U369 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[85]), .Z(n256));
Q_AN02 U370 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[84]), .Z(n257));
Q_AN02 U371 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[83]), .Z(n258));
Q_AN02 U372 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[82]), .Z(n259));
Q_AN02 U373 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[81]), .Z(n260));
Q_AN02 U374 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[80]), .Z(n261));
Q_AN02 U375 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[79]), .Z(n262));
Q_AN02 U376 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[78]), .Z(n263));
Q_AN02 U377 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[77]), .Z(n264));
Q_AN02 U378 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[76]), .Z(n265));
Q_AN02 U379 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[75]), .Z(n266));
Q_AN02 U380 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[74]), .Z(n267));
Q_AN02 U381 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[73]), .Z(n268));
Q_AN02 U382 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[72]), .Z(n269));
Q_AN02 U383 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[71]), .Z(n270));
Q_AN02 U384 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[70]), .Z(n271));
Q_AN02 U385 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[69]), .Z(n272));
Q_AN02 U386 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[68]), .Z(n273));
Q_AN02 U387 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[67]), .Z(n274));
Q_AN02 U388 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[66]), .Z(n275));
Q_AN02 U389 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[65]), .Z(n276));
Q_AN02 U390 ( .A0(n206), .A1(_zyixc_port_0_0_s2h[64]), .Z(n277));
Q_AN02 U391 ( .A0(n208), .A1(n163), .Z(n278));
Q_AN02 U392 ( .A0(n208), .A1(n165), .Z(n279));
Q_AN02 U393 ( .A0(n208), .A1(n167), .Z(n280));
Q_AN02 U394 ( .A0(n208), .A1(n169), .Z(n281));
Q_AN02 U395 ( .A0(n208), .A1(n171), .Z(n282));
Q_AN02 U396 ( .A0(n208), .A1(n173), .Z(n283));
Q_AN02 U397 ( .A0(n208), .A1(n175), .Z(n284));
Q_AN02 U398 ( .A0(n208), .A1(n286), .Z(n285));
Q_OR02 U399 ( .A0(pslverr), .A1(n288), .Z(n287));
Q_NR02 U400 ( .A0(n290), .A1(n289), .Z(n288));
Q_OR03 U401 ( .A0(bus_timer[1]), .A1(bus_timer[0]), .A2(n291), .Z(n289));
Q_OR03 U402 ( .A0(bus_timer[4]), .A1(bus_timer[3]), .A2(n294), .Z(n290));
Q_OR03 U403 ( .A0(bus_timer[7]), .A1(n292), .A2(n293), .Z(n291));
Q_INV U404 ( .A(bus_timer[6]), .Z(n292));
Q_INV U405 ( .A(bus_timer[5]), .Z(n293));
Q_AO21 U406 ( .A0(n296), .A1(n295), .B0(n297), .Z(n192));
Q_NR02 U407 ( .A0(bus_timer[3]), .A1(bus_timer[2]), .Z(n295));
Q_AN02 U408 ( .A0(n301), .A1(n298), .Z(n296));
Q_OA21 U409 ( .A0(n300), .A1(n299), .B0(n301), .Z(n297));
Q_INV U410 ( .A(reset_n), .Z(n302));
Q_FDP0 _zzM2L46_mdxP0_bus_timer_Dwen5_REG  ( .CK(clk), .D(n302), .Q(_zzM2L46_mdxP0_bus_timer_Dwen5), .QN( ));
Q_FDP0 _zzM2L46_mdxP0_pwdata_Dwen4_REG  ( .CK(clk), .D(n302), .Q(_zzM2L46_mdxP0_pwdata_Dwen4), .QN( ));
Q_FDP0 _zzM2L46_mdxP0_paddr_Dwen3_REG  ( .CK(clk), .D(n302), .Q(_zzM2L46_mdxP0_paddr_Dwen3), .QN( ));
Q_FDP0 _zzM2L46_mdxP0_pwrite_Dwen2_REG  ( .CK(clk), .D(n302), .Q(_zzM2L46_mdxP0_pwrite_Dwen2), .QN( ));
Q_FDP0 _zzM2L46_mdxP0_penable_Dwen1_REG  ( .CK(clk), .D(n302), .Q(_zzM2L46_mdxP0_penable_Dwen1), .QN( ));
Q_FDP0 _zzM2L46_mdxP0_psel_Dwen0_REG  ( .CK(clk), .D(n302), .Q(_zzM2L46_mdxP0_psel_Dwen0), .QN( ));
Q_NOT_TOUCH _zzqnt ( .sig());
ixc_assign _zz_strnp_0 ( _zy_simnet_psel_0_w$, psel);
ixc_assign _zz_strnp_1 ( _zy_simnet_penable_1_w$, penable);
ixc_assign_20 _zz_strnp_2 ( _zy_simnet_paddr_2_w$[0:19], paddr[19:0]);
ixc_assign_32 _zz_strnp_3 ( _zy_simnet_pwdata_3_w$[0:31], pwdata[31:0]);
ixc_assign _zz_strnp_4 ( _zy_simnet_pwrite_4_w$, pwrite);
ixc_mem_call_96_8 _zzixc_tfport_0_0 ( _zyixc_port_0_0_req, 
	_zyixc_port_0_0_s2h[95:0], _zyixc_port_0_0_isf, _zyixc_port_0_0_ack, 
	_zyixc_port_0_0_h2s[7:0], _zyixc_port_0_0_osf, n314, n313);
ixc_mem_call_64_40 _zzixc_tfport_0_1 ( _zyixc_port_0_1_req, 
	_zyixc_port_0_1_s2h[63:0], _zyixc_port_0_1_isf, _zyixc_port_0_1_ack, 
	_zyixc_port_0_1_h2s[39:0], _zyixc_port_0_1_osf, n312, n311);
Q_OR03 U425 ( .A0(_zyM2L73_pbcCapEn1), .A1(_zyM2L79_pbcCapEn2), .A2(_zyM2L90_pbcCapEn3), .Z(n310));
ixc_mevClk_2_0_0_1 _zzM2L61_pbcMevClk4 ( _zyM2L61_pbcMevClk4, { 
	_zyixc_port_0_0_req, clk}, { _zyM2L61_pbcCapEn0, n310}, n309, n308, 
	_zyM2L61_pbcReq4, _zyM2L61_pbcBusy4, _zyM2L61_pbcWait4);
Q_OR03 U427 ( .A0(_zyM2L104_pbcCapEn6), .A1(_zyM2L110_pbcCapEn7), .A2(_zyM2L121_pbcCapEn8), .Z(n307));
ixc_mevClk_2_0_0_1 _zzM2L94_pbcMevClk9 ( _zyM2L94_pbcMevClk9, { 
	_zyixc_port_0_1_req, clk}, { _zyM2L94_pbcCapEn5, n307}, n306, n305, 
	_zyM2L94_pbcReq9, _zyM2L94_pbcBusy9, _zyM2L94_pbcWait9);
ixc_capLoopXp _zzM2L10_bcBehEvalP0 ( _zzM2_bcBehEvalClk, n1,, _zzM2_bcBehHalt);
ixc_mdrOn _zzM2L46_mdxP0_OnP ( _zzM2L46_mdxP0_On, _zzM2L46_mdxP0_EnNxt, 
	_zzM2L46_mdxP0_En);
ixc_mdrOn _zzM2L61_mdxP1_OnP ( _zzM2L61_mdxP1_On, _zzM2L61_mdxP1_EnNxt, 
	_zzM2L61_mdxP1_En);
ixc_mdrOn _zzM2L94_mdxP2_OnP ( _zzM2L94_mdxP2_On, _zzM2L94_mdxP2_EnNxt, 
	_zzM2L94_mdxP2_En);
ixc_sampleLT _zzpsel_M2L19_mdxSpLt6 ( _zzpsel_M2L19_mdxSvLt6, psel);
ixc_sampleLT _zzpenable_M2L20_mdxSpLt7 ( _zzpenable_M2L20_mdxSvLt7, penable);
ixc_sampleLT _zzpwrite_M2L23_mdxSpLt8 ( _zzpwrite_M2L23_mdxSvLt8, pwrite);
ixc_sampleLT_20 _zzpaddr_M2L21_mdxSpLt9 ( _zzpaddr_M2L21_mdxSvLt9[19:0], 
	paddr[19:0]);
ixc_sampleLT_32 _zzpwdata_M2L22_mdxSpLt10 ( _zzpwdata_M2L22_mdxSvLt10[31:0], 
	pwdata[31:0]);
ixc_sampleLT_8 _zzbus_timer_M2L29_mdxSpLt11 ( 
	_zzbus_timer_M2L29_mdxSvLt11[7:0], bus_timer[7:0]);
ixc_assign _zzmdx1 ( _zzmdxOne, n303);
Q_FDP4EP _zzM2L46_mdxP0_En_REG  ( .CK(clk), .CE(n302), .R(n304), .D(_zzM2L46_mdxP0_EnNxt), .Q(_zzM2L46_mdxP0_En));
Q_FDP4EP _zzM2L46_mdxP0_psel_wr0_REG  ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_psel_wr0));
Q_FDP4EP _zzM2L46_mdxP0_penable_wr1_REG  ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_penable_wr1));
Q_FDP4EP _zzM2L46_mdxP0_pwrite_wr2_REG  ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwrite_wr2));
Q_FDP4EP \_zzM2L46_mdxP0_paddr_wr3_REG[19] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_paddr_wr3[19]));
Q_FDP4EP \_zzM2L46_mdxP0_paddr_wr3_REG[18] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_paddr_wr3[18]));
Q_FDP4EP \_zzM2L46_mdxP0_paddr_wr3_REG[17] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_paddr_wr3[17]));
Q_FDP4EP \_zzM2L46_mdxP0_paddr_wr3_REG[16] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_paddr_wr3[16]));
Q_FDP4EP \_zzM2L46_mdxP0_paddr_wr3_REG[15] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_paddr_wr3[15]));
Q_FDP4EP \_zzM2L46_mdxP0_paddr_wr3_REG[14] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_paddr_wr3[14]));
Q_FDP4EP \_zzM2L46_mdxP0_paddr_wr3_REG[13] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_paddr_wr3[13]));
Q_FDP4EP \_zzM2L46_mdxP0_paddr_wr3_REG[12] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_paddr_wr3[12]));
Q_FDP4EP \_zzM2L46_mdxP0_paddr_wr3_REG[11] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_paddr_wr3[11]));
Q_FDP4EP \_zzM2L46_mdxP0_paddr_wr3_REG[10] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_paddr_wr3[10]));
Q_FDP4EP \_zzM2L46_mdxP0_paddr_wr3_REG[9] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_paddr_wr3[9]));
Q_FDP4EP \_zzM2L46_mdxP0_paddr_wr3_REG[8] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_paddr_wr3[8]));
Q_FDP4EP \_zzM2L46_mdxP0_paddr_wr3_REG[7] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_paddr_wr3[7]));
Q_FDP4EP \_zzM2L46_mdxP0_paddr_wr3_REG[6] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_paddr_wr3[6]));
Q_FDP4EP \_zzM2L46_mdxP0_paddr_wr3_REG[5] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_paddr_wr3[5]));
Q_FDP4EP \_zzM2L46_mdxP0_paddr_wr3_REG[4] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_paddr_wr3[4]));
Q_FDP4EP \_zzM2L46_mdxP0_paddr_wr3_REG[3] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_paddr_wr3[3]));
Q_FDP4EP \_zzM2L46_mdxP0_paddr_wr3_REG[2] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_paddr_wr3[2]));
Q_FDP4EP \_zzM2L46_mdxP0_paddr_wr3_REG[1] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_paddr_wr3[1]));
Q_FDP4EP \_zzM2L46_mdxP0_paddr_wr3_REG[0] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_paddr_wr3[0]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[31] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[31]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[30] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[30]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[29] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[29]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[28] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[28]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[27] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[27]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[26] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[26]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[25] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[25]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[24] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[24]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[23] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[23]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[22] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[22]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[21] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[21]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[20] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[20]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[19] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[19]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[18] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[18]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[17] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[17]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[16] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[16]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[15] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[15]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[14] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[14]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[13] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[13]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[12] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[12]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[11] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[11]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[10] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[10]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[9] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[9]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[8] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[8]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[7] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[7]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[6] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[6]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[5] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[5]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[4] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[4]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[3] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[3]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[2] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[2]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[1] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[1]));
Q_FDP4EP \_zzM2L46_mdxP0_pwdata_wr4_REG[0] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_pwdata_wr4[0]));
Q_FDP4EP \_zzM2L46_mdxP0_bus_timer_wr5_REG[7] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_bus_timer_wr5[7]));
Q_FDP4EP \_zzM2L46_mdxP0_bus_timer_wr5_REG[6] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_bus_timer_wr5[6]));
Q_FDP4EP \_zzM2L46_mdxP0_bus_timer_wr5_REG[5] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_bus_timer_wr5[5]));
Q_FDP4EP \_zzM2L46_mdxP0_bus_timer_wr5_REG[4] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_bus_timer_wr5[4]));
Q_FDP4EP \_zzM2L46_mdxP0_bus_timer_wr5_REG[3] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_bus_timer_wr5[3]));
Q_FDP4EP \_zzM2L46_mdxP0_bus_timer_wr5_REG[2] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_bus_timer_wr5[2]));
Q_FDP4EP \_zzM2L46_mdxP0_bus_timer_wr5_REG[1] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_bus_timer_wr5[1]));
Q_FDP4EP \_zzM2L46_mdxP0_bus_timer_wr5_REG[0] ( .CK(clk), .CE(n302), .R(n304), .D(n304), .Q(_zzM2L46_mdxP0_bus_timer_wr5[0]));
Q_INV U504 ( .A(n220), .Z(n316));
Q_FDP4EP _zzM2L61_mdxP1_En_REG  ( .CK(_zyM2L61_pbcMevClk4), .CE(n316), .R(n304), .D(_zzM2L61_mdxP1_EnNxt), .Q(_zzM2L61_mdxP1_En));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[63] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[63]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[63]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[62] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[62]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[62]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[61] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[61]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[61]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[60] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[60]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[60]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[59] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[59]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[59]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[58] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[58]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[58]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[57] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[57]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[57]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[56] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[56]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[56]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[55] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[55]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[55]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[54] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[54]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[54]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[53] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[53]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[53]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[52] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[52]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[52]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[51] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[51]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[51]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[50] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[50]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[50]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[49] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[49]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[49]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[48] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[48]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[48]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[47] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[47]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[47]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[46] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[46]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[46]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[45] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[45]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[45]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[44] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[44]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[44]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[43] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[43]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[43]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[42] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[42]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[42]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[41] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[41]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[41]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[40] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[40]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[40]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[39] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[39]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[39]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[38] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[38]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[38]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[37] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[37]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[37]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[36] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[36]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[36]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[35] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[35]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[35]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[34] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[34]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[34]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[33] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[33]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[33]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[32] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[32]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[32]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[31] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[31]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[31]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[30] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[30]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[30]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[29] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[29]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[29]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[28] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[28]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[28]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[27] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[27]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[27]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[26] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[26]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[26]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[25] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[25]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[25]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[24] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[24]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[24]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[23] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[23]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[23]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[22] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[22]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[22]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[21] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[21]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[21]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[20] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[20]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[20]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[19] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[19]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[19]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[18] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[18]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[18]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[17] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[17]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[17]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[16] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[16]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[16]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[15] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[15]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[15]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[14] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[14]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[14]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[13] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[13]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[13]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[12] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[12]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[12]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[11] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[11]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[11]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[10] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[10]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[10]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[9] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[9]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[9]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[8] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[8]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[8]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[7] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[7]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[7]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[6] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[6]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[6]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[5] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[5]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[5]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[4] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[4]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[4]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[3] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[3]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[3]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[2] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[2]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[2]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[1] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[1]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[1]));
Q_FDP4EP \_zyaddr_L62_tfiV0_M2_pbcG0_REG[0] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[0]), .Q(_zyaddr_L62_tfiV0_M2_pbcG0[0]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[31] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[95]), .Q(_zydata_L63_tfiV1_M2_pbcG1[31]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[30] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[94]), .Q(_zydata_L63_tfiV1_M2_pbcG1[30]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[29] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[93]), .Q(_zydata_L63_tfiV1_M2_pbcG1[29]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[28] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[92]), .Q(_zydata_L63_tfiV1_M2_pbcG1[28]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[27] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[91]), .Q(_zydata_L63_tfiV1_M2_pbcG1[27]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[26] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[90]), .Q(_zydata_L63_tfiV1_M2_pbcG1[26]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[25] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[89]), .Q(_zydata_L63_tfiV1_M2_pbcG1[25]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[24] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[88]), .Q(_zydata_L63_tfiV1_M2_pbcG1[24]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[23] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[87]), .Q(_zydata_L63_tfiV1_M2_pbcG1[23]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[22] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[86]), .Q(_zydata_L63_tfiV1_M2_pbcG1[22]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[21] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[85]), .Q(_zydata_L63_tfiV1_M2_pbcG1[21]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[20] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[84]), .Q(_zydata_L63_tfiV1_M2_pbcG1[20]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[19] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[83]), .Q(_zydata_L63_tfiV1_M2_pbcG1[19]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[18] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[82]), .Q(_zydata_L63_tfiV1_M2_pbcG1[18]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[17] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[81]), .Q(_zydata_L63_tfiV1_M2_pbcG1[17]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[16] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[80]), .Q(_zydata_L63_tfiV1_M2_pbcG1[16]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[15] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[79]), .Q(_zydata_L63_tfiV1_M2_pbcG1[15]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[14] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[78]), .Q(_zydata_L63_tfiV1_M2_pbcG1[14]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[13] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[77]), .Q(_zydata_L63_tfiV1_M2_pbcG1[13]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[12] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[76]), .Q(_zydata_L63_tfiV1_M2_pbcG1[12]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[11] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[75]), .Q(_zydata_L63_tfiV1_M2_pbcG1[11]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[10] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[74]), .Q(_zydata_L63_tfiV1_M2_pbcG1[10]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[9] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[73]), .Q(_zydata_L63_tfiV1_M2_pbcG1[9]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[8] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[72]), .Q(_zydata_L63_tfiV1_M2_pbcG1[8]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[7] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[71]), .Q(_zydata_L63_tfiV1_M2_pbcG1[7]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[6] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[70]), .Q(_zydata_L63_tfiV1_M2_pbcG1[6]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[5] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[69]), .Q(_zydata_L63_tfiV1_M2_pbcG1[5]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[4] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[68]), .Q(_zydata_L63_tfiV1_M2_pbcG1[4]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[3] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[67]), .Q(_zydata_L63_tfiV1_M2_pbcG1[3]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[2] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[66]), .Q(_zydata_L63_tfiV1_M2_pbcG1[2]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[1] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[65]), .Q(_zydata_L63_tfiV1_M2_pbcG1[1]));
Q_FDP4EP \_zydata_L63_tfiV1_M2_pbcG1_REG[0] ( .CK(_zyM2L61_pbcMevClk4), .CE(n198), .R(n304), .D(_zyixc_port_0_0_s2h[64]), .Q(_zydata_L63_tfiV1_M2_pbcG1[0]));
Q_FDP4EP \_zyixc_port_0_0_h2s_REG[7] ( .CK(_zyM2L61_pbcMevClk4), .CE(n197), .R(n304), .D(n304), .Q(_zyixc_port_0_0_h2s[7]));
Q_FDP4EP \_zyixc_port_0_0_h2s_REG[6] ( .CK(_zyM2L61_pbcMevClk4), .CE(n197), .R(n304), .D(n304), .Q(_zyixc_port_0_0_h2s[6]));
Q_FDP4EP \_zyixc_port_0_0_h2s_REG[5] ( .CK(_zyM2L61_pbcMevClk4), .CE(n197), .R(n304), .D(n304), .Q(_zyixc_port_0_0_h2s[5]));
Q_FDP4EP \_zyixc_port_0_0_h2s_REG[4] ( .CK(_zyM2L61_pbcMevClk4), .CE(n197), .R(n304), .D(n304), .Q(_zyixc_port_0_0_h2s[4]));
Q_FDP4EP \_zyixc_port_0_0_h2s_REG[3] ( .CK(_zyM2L61_pbcMevClk4), .CE(n197), .R(n304), .D(n304), .Q(_zyixc_port_0_0_h2s[3]));
Q_FDP4EP \_zyixc_port_0_0_h2s_REG[2] ( .CK(_zyM2L61_pbcMevClk4), .CE(n197), .R(n304), .D(n304), .Q(_zyixc_port_0_0_h2s[2]));
Q_FDP4EP \_zyixc_port_0_0_h2s_REG[1] ( .CK(_zyM2L61_pbcMevClk4), .CE(n197), .R(n304), .D(n304), .Q(_zyixc_port_0_0_h2s[1]));
Q_FDP4EP \_zyixc_port_0_0_h2s_REG[0] ( .CK(_zyM2L61_pbcMevClk4), .CE(n197), .R(n304), .D(_zyresponse_L64_tfiV2_M2_pbcG2), .Q(_zyixc_port_0_0_h2s[0]));
Q_INV U610 ( .A(_zyixc_port_0_0_ack), .Z(n317));
Q_FDP4EP _zyixc_port_0_0_ack_REG  ( .CK(_zyM2L61_pbcMevClk4), .CE(n197), .R(n304), .D(n317), .Q(_zyixc_port_0_0_ack));
Q_INV U612 ( .A(n221), .Z(n318));
Q_FDP4EP _zyresponse_L64_tfiV2_M2_pbcG2_REG  ( .CK(_zyM2L61_pbcMevClk4), .CE(n318), .R(n304), .D(n287), .Q(_zyresponse_L64_tfiV2_M2_pbcG2));
Q_FDP4EP \_zzM2L61_mdxP1_paddr_wr3_REG[19] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n226), .Q(_zzM2L61_mdxP1_paddr_wr3[19]));
Q_FDP4EP \_zzM2L61_mdxP1_paddr_wr3_REG[18] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n227), .Q(_zzM2L61_mdxP1_paddr_wr3[18]));
Q_FDP4EP \_zzM2L61_mdxP1_paddr_wr3_REG[17] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n228), .Q(_zzM2L61_mdxP1_paddr_wr3[17]));
Q_FDP4EP \_zzM2L61_mdxP1_paddr_wr3_REG[16] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n229), .Q(_zzM2L61_mdxP1_paddr_wr3[16]));
Q_FDP4EP \_zzM2L61_mdxP1_paddr_wr3_REG[15] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n230), .Q(_zzM2L61_mdxP1_paddr_wr3[15]));
Q_FDP4EP \_zzM2L61_mdxP1_paddr_wr3_REG[14] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n231), .Q(_zzM2L61_mdxP1_paddr_wr3[14]));
Q_FDP4EP \_zzM2L61_mdxP1_paddr_wr3_REG[13] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n232), .Q(_zzM2L61_mdxP1_paddr_wr3[13]));
Q_FDP4EP \_zzM2L61_mdxP1_paddr_wr3_REG[12] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n233), .Q(_zzM2L61_mdxP1_paddr_wr3[12]));
Q_FDP4EP \_zzM2L61_mdxP1_paddr_wr3_REG[11] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n234), .Q(_zzM2L61_mdxP1_paddr_wr3[11]));
Q_FDP4EP \_zzM2L61_mdxP1_paddr_wr3_REG[10] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n235), .Q(_zzM2L61_mdxP1_paddr_wr3[10]));
Q_FDP4EP \_zzM2L61_mdxP1_paddr_wr3_REG[9] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n236), .Q(_zzM2L61_mdxP1_paddr_wr3[9]));
Q_FDP4EP \_zzM2L61_mdxP1_paddr_wr3_REG[8] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n237), .Q(_zzM2L61_mdxP1_paddr_wr3[8]));
Q_FDP4EP \_zzM2L61_mdxP1_paddr_wr3_REG[7] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n238), .Q(_zzM2L61_mdxP1_paddr_wr3[7]));
Q_FDP4EP \_zzM2L61_mdxP1_paddr_wr3_REG[6] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n239), .Q(_zzM2L61_mdxP1_paddr_wr3[6]));
Q_FDP4EP \_zzM2L61_mdxP1_paddr_wr3_REG[5] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n240), .Q(_zzM2L61_mdxP1_paddr_wr3[5]));
Q_FDP4EP \_zzM2L61_mdxP1_paddr_wr3_REG[4] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n241), .Q(_zzM2L61_mdxP1_paddr_wr3[4]));
Q_FDP4EP \_zzM2L61_mdxP1_paddr_wr3_REG[3] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n242), .Q(_zzM2L61_mdxP1_paddr_wr3[3]));
Q_FDP4EP \_zzM2L61_mdxP1_paddr_wr3_REG[2] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n243), .Q(_zzM2L61_mdxP1_paddr_wr3[2]));
Q_FDP4EP \_zzM2L61_mdxP1_paddr_wr3_REG[1] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n244), .Q(_zzM2L61_mdxP1_paddr_wr3[1]));
Q_FDP4EP \_zzM2L61_mdxP1_paddr_wr3_REG[0] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n245), .Q(_zzM2L61_mdxP1_paddr_wr3[0]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[31] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n246), .Q(_zzM2L61_mdxP1_pwdata_wr4[31]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[30] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n247), .Q(_zzM2L61_mdxP1_pwdata_wr4[30]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[29] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n248), .Q(_zzM2L61_mdxP1_pwdata_wr4[29]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[28] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n249), .Q(_zzM2L61_mdxP1_pwdata_wr4[28]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[27] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n250), .Q(_zzM2L61_mdxP1_pwdata_wr4[27]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[26] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n251), .Q(_zzM2L61_mdxP1_pwdata_wr4[26]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[25] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n252), .Q(_zzM2L61_mdxP1_pwdata_wr4[25]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[24] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n253), .Q(_zzM2L61_mdxP1_pwdata_wr4[24]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[23] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n254), .Q(_zzM2L61_mdxP1_pwdata_wr4[23]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[22] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n255), .Q(_zzM2L61_mdxP1_pwdata_wr4[22]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[21] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n256), .Q(_zzM2L61_mdxP1_pwdata_wr4[21]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[20] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n257), .Q(_zzM2L61_mdxP1_pwdata_wr4[20]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[19] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n258), .Q(_zzM2L61_mdxP1_pwdata_wr4[19]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[18] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n259), .Q(_zzM2L61_mdxP1_pwdata_wr4[18]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[17] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n260), .Q(_zzM2L61_mdxP1_pwdata_wr4[17]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[16] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n261), .Q(_zzM2L61_mdxP1_pwdata_wr4[16]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[15] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n262), .Q(_zzM2L61_mdxP1_pwdata_wr4[15]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[14] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n263), .Q(_zzM2L61_mdxP1_pwdata_wr4[14]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[13] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n264), .Q(_zzM2L61_mdxP1_pwdata_wr4[13]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[12] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n265), .Q(_zzM2L61_mdxP1_pwdata_wr4[12]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[11] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n266), .Q(_zzM2L61_mdxP1_pwdata_wr4[11]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[10] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n267), .Q(_zzM2L61_mdxP1_pwdata_wr4[10]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[9] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n268), .Q(_zzM2L61_mdxP1_pwdata_wr4[9]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[8] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n269), .Q(_zzM2L61_mdxP1_pwdata_wr4[8]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[7] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n270), .Q(_zzM2L61_mdxP1_pwdata_wr4[7]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[6] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n271), .Q(_zzM2L61_mdxP1_pwdata_wr4[6]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[5] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n272), .Q(_zzM2L61_mdxP1_pwdata_wr4[5]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[4] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n273), .Q(_zzM2L61_mdxP1_pwdata_wr4[4]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[3] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n274), .Q(_zzM2L61_mdxP1_pwdata_wr4[3]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[2] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n275), .Q(_zzM2L61_mdxP1_pwdata_wr4[2]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[1] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n276), .Q(_zzM2L61_mdxP1_pwdata_wr4[1]));
Q_FDP4EP \_zzM2L61_mdxP1_pwdata_wr4_REG[0] ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n277), .Q(_zzM2L61_mdxP1_pwdata_wr4[0]));
Q_FDP4EP \_zzM2L61_mdxP1_bus_timer_wr5_REG[7] ( .CK(_zyM2L61_pbcMevClk4), .CE(n209), .R(n304), .D(n278), .Q(_zzM2L61_mdxP1_bus_timer_wr5[7]));
Q_FDP4EP \_zzM2L61_mdxP1_bus_timer_wr5_REG[6] ( .CK(_zyM2L61_pbcMevClk4), .CE(n209), .R(n304), .D(n279), .Q(_zzM2L61_mdxP1_bus_timer_wr5[6]));
Q_FDP4EP \_zzM2L61_mdxP1_bus_timer_wr5_REG[5] ( .CK(_zyM2L61_pbcMevClk4), .CE(n209), .R(n304), .D(n280), .Q(_zzM2L61_mdxP1_bus_timer_wr5[5]));
Q_FDP4EP \_zzM2L61_mdxP1_bus_timer_wr5_REG[4] ( .CK(_zyM2L61_pbcMevClk4), .CE(n209), .R(n304), .D(n281), .Q(_zzM2L61_mdxP1_bus_timer_wr5[4]));
Q_FDP4EP \_zzM2L61_mdxP1_bus_timer_wr5_REG[3] ( .CK(_zyM2L61_pbcMevClk4), .CE(n209), .R(n304), .D(n282), .Q(_zzM2L61_mdxP1_bus_timer_wr5[3]));
Q_FDP4EP \_zzM2L61_mdxP1_bus_timer_wr5_REG[2] ( .CK(_zyM2L61_pbcMevClk4), .CE(n209), .R(n304), .D(n283), .Q(_zzM2L61_mdxP1_bus_timer_wr5[2]));
Q_FDP4EP \_zzM2L61_mdxP1_bus_timer_wr5_REG[1] ( .CK(_zyM2L61_pbcMevClk4), .CE(n209), .R(n304), .D(n284), .Q(_zzM2L61_mdxP1_bus_timer_wr5[1]));
Q_FDP4EP \_zzM2L61_mdxP1_bus_timer_wr5_REG[0] ( .CK(_zyM2L61_pbcMevClk4), .CE(n209), .R(n304), .D(n285), .Q(_zzM2L61_mdxP1_bus_timer_wr5[0]));
Q_FDP4EP _zyM2L61_pbcCapEn0_REG  ( .CK(_zyM2L61_pbcMevClk4), .CE(n196), .R(n304), .D(n199), .Q(_zyM2L61_pbcCapEn0));
Q_FDP4EP _zyM2L73_pbcCapEn1_REG  ( .CK(_zyM2L61_pbcMevClk4), .CE(n195), .R(n304), .D(n200), .Q(_zyM2L73_pbcCapEn1));
Q_FDP4EP _zyM2L79_pbcCapEn2_REG  ( .CK(_zyM2L61_pbcMevClk4), .CE(n194), .R(n304), .D(n208), .Q(_zyM2L79_pbcCapEn2));
Q_INV U677 ( .A(n215), .Z(n319));
Q_FDP4EP _zyM2L90_pbcCapEn3_REG  ( .CK(_zyM2L61_pbcMevClk4), .CE(n319), .R(n304), .D(n201), .Q(_zyM2L90_pbcCapEn3));
Q_FDP4EP \_zyM2L61_pbcFsm0_s_REG[1] ( .CK(_zyM2L61_pbcMevClk4), .CE(n193), .R(n304), .D(n225), .Q(_zyM2L61_pbcFsm0_s[1]));
Q_INV U680 ( .A(_zyM2L61_pbcFsm0_s[1]), .Z(n218));
Q_FDP4EP \_zyM2L61_pbcFsm0_s_REG[0] ( .CK(_zyM2L61_pbcMevClk4), .CE(n193), .R(n304), .D(n202), .Q(_zyM2L61_pbcFsm0_s[0]));
Q_INV U682 ( .A(_zyM2L61_pbcFsm0_s[0]), .Z(n200));
Q_FDP4EP _zzM2L61_mdxP1_psel_wr0_REG  ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n206), .Q(_zzM2L61_mdxP1_psel_wr0));
Q_FDP4EP _zzM2L61_mdxP1_penable_wr1_REG  ( .CK(_zyM2L61_pbcMevClk4), .CE(n205), .R(n304), .D(n204), .Q(_zzM2L61_mdxP1_penable_wr1));
Q_FDP4EP _zzM2L61_mdxP1_pwrite_wr2_REG  ( .CK(_zyM2L61_pbcMevClk4), .CE(n207), .R(n304), .D(n206), .Q(_zzM2L61_mdxP1_pwrite_wr2));
Q_FDP4EP _zyM2L61_pbcEn10_REG  ( .CK(_zyM2L61_pbcMevClk4), .CE(n209), .R(n304), .D(n210), .Q(_zyM2L61_pbcEn10));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[31] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[31]), .Q(_zyixc_port_0_1_h2s[31]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[30] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[30]), .Q(_zyixc_port_0_1_h2s[30]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[29] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[29]), .Q(_zyixc_port_0_1_h2s[29]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[28] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[28]), .Q(_zyixc_port_0_1_h2s[28]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[27] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[27]), .Q(_zyixc_port_0_1_h2s[27]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[26] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[26]), .Q(_zyixc_port_0_1_h2s[26]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[25] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[25]), .Q(_zyixc_port_0_1_h2s[25]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[24] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[24]), .Q(_zyixc_port_0_1_h2s[24]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[23] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[23]), .Q(_zyixc_port_0_1_h2s[23]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[22] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[22]), .Q(_zyixc_port_0_1_h2s[22]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[21] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[21]), .Q(_zyixc_port_0_1_h2s[21]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[20] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[20]), .Q(_zyixc_port_0_1_h2s[20]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[19] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[19]), .Q(_zyixc_port_0_1_h2s[19]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[18] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[18]), .Q(_zyixc_port_0_1_h2s[18]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[17] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[17]), .Q(_zyixc_port_0_1_h2s[17]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[16] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[16]), .Q(_zyixc_port_0_1_h2s[16]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[15] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[15]), .Q(_zyixc_port_0_1_h2s[15]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[14] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[14]), .Q(_zyixc_port_0_1_h2s[14]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[13] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[13]), .Q(_zyixc_port_0_1_h2s[13]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[12] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[12]), .Q(_zyixc_port_0_1_h2s[12]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[11] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[11]), .Q(_zyixc_port_0_1_h2s[11]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[10] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[10]), .Q(_zyixc_port_0_1_h2s[10]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[9] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[9]), .Q(_zyixc_port_0_1_h2s[9]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[8] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[8]), .Q(_zyixc_port_0_1_h2s[8]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[7] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[7]), .Q(_zyixc_port_0_1_h2s[7]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[6] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[6]), .Q(_zyixc_port_0_1_h2s[6]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[5] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[5]), .Q(_zyixc_port_0_1_h2s[5]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[4] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[4]), .Q(_zyixc_port_0_1_h2s[4]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[3] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[3]), .Q(_zyixc_port_0_1_h2s[3]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[2] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[2]), .Q(_zyixc_port_0_1_h2s[2]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[1] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[1]), .Q(_zyixc_port_0_1_h2s[1]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[0] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zydata_L96_tfiV4_M2_pbcG4[0]), .Q(_zyixc_port_0_1_h2s[0]));
Q_INV U719 ( .A(n130), .Z(n320));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[31] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[31]), .Q(_zydata_L96_tfiV4_M2_pbcG4[31]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[30] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[30]), .Q(_zydata_L96_tfiV4_M2_pbcG4[30]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[29] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[29]), .Q(_zydata_L96_tfiV4_M2_pbcG4[29]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[28] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[28]), .Q(_zydata_L96_tfiV4_M2_pbcG4[28]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[27] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[27]), .Q(_zydata_L96_tfiV4_M2_pbcG4[27]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[26] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[26]), .Q(_zydata_L96_tfiV4_M2_pbcG4[26]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[25] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[25]), .Q(_zydata_L96_tfiV4_M2_pbcG4[25]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[24] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[24]), .Q(_zydata_L96_tfiV4_M2_pbcG4[24]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[23] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[23]), .Q(_zydata_L96_tfiV4_M2_pbcG4[23]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[22] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[22]), .Q(_zydata_L96_tfiV4_M2_pbcG4[22]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[21] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[21]), .Q(_zydata_L96_tfiV4_M2_pbcG4[21]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[20] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[20]), .Q(_zydata_L96_tfiV4_M2_pbcG4[20]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[19] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[19]), .Q(_zydata_L96_tfiV4_M2_pbcG4[19]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[18] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[18]), .Q(_zydata_L96_tfiV4_M2_pbcG4[18]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[17] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[17]), .Q(_zydata_L96_tfiV4_M2_pbcG4[17]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[16] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[16]), .Q(_zydata_L96_tfiV4_M2_pbcG4[16]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[15] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[15]), .Q(_zydata_L96_tfiV4_M2_pbcG4[15]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[14] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[14]), .Q(_zydata_L96_tfiV4_M2_pbcG4[14]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[13] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[13]), .Q(_zydata_L96_tfiV4_M2_pbcG4[13]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[12] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[12]), .Q(_zydata_L96_tfiV4_M2_pbcG4[12]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[11] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[11]), .Q(_zydata_L96_tfiV4_M2_pbcG4[11]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[10] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[10]), .Q(_zydata_L96_tfiV4_M2_pbcG4[10]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[9] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[9]), .Q(_zydata_L96_tfiV4_M2_pbcG4[9]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[8] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[8]), .Q(_zydata_L96_tfiV4_M2_pbcG4[8]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[7] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[7]), .Q(_zydata_L96_tfiV4_M2_pbcG4[7]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[6] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[6]), .Q(_zydata_L96_tfiV4_M2_pbcG4[6]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[5] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[5]), .Q(_zydata_L96_tfiV4_M2_pbcG4[5]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[4] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[4]), .Q(_zydata_L96_tfiV4_M2_pbcG4[4]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[3] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[3]), .Q(_zydata_L96_tfiV4_M2_pbcG4[3]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[2] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[2]), .Q(_zydata_L96_tfiV4_M2_pbcG4[2]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[1] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[1]), .Q(_zydata_L96_tfiV4_M2_pbcG4[1]));
Q_FDP4EP \_zydata_L96_tfiV4_M2_pbcG4_REG[0] ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(prdata[0]), .Q(_zydata_L96_tfiV4_M2_pbcG4[0]));
Q_INV U752 ( .A(n129), .Z(n321));
Q_FDP4EP _zzM2L94_mdxP2_En_REG  ( .CK(_zyM2L94_pbcMevClk9), .CE(n321), .R(n304), .D(_zzM2L94_mdxP2_EnNxt), .Q(_zzM2L94_mdxP2_En));
Q_FDP4EP _zzM2L94_mdxP2_pwrite_wr2_REG  ( .CK(_zyM2L94_pbcMevClk9), .CE(n115), .R(n304), .D(n304), .Q(_zzM2L94_mdxP2_pwrite_wr2));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[63] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[63]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[63]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[62] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[62]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[62]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[61] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[61]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[61]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[60] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[60]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[60]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[59] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[59]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[59]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[58] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[58]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[58]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[57] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[57]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[57]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[56] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[56]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[56]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[55] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[55]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[55]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[54] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[54]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[54]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[53] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[53]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[53]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[52] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[52]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[52]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[51] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[51]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[51]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[50] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[50]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[50]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[49] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[49]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[49]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[48] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[48]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[48]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[47] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[47]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[47]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[46] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[46]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[46]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[45] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[45]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[45]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[44] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[44]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[44]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[43] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[43]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[43]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[42] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[42]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[42]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[41] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[41]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[41]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[40] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[40]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[40]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[39] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[39]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[39]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[38] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[38]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[38]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[37] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[37]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[37]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[36] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[36]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[36]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[35] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[35]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[35]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[34] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[34]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[34]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[33] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[33]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[33]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[32] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[32]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[32]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[31] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[31]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[31]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[30] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[30]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[30]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[29] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[29]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[29]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[28] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[28]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[28]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[27] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[27]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[27]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[26] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[26]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[26]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[25] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[25]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[25]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[24] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[24]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[24]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[23] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[23]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[23]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[22] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[22]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[22]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[21] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[21]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[21]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[20] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[20]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[20]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[19] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[19]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[19]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[18] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[18]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[18]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[17] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[17]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[17]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[16] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[16]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[16]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[15] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[15]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[15]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[14] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[14]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[14]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[13] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[13]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[13]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[12] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[12]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[12]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[11] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[11]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[11]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[10] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[10]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[10]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[9] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[9]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[9]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[8] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[8]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[8]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[7] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[7]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[7]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[6] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[6]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[6]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[5] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[5]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[5]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[4] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[4]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[4]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[3] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[3]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[3]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[2] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[2]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[2]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[1] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[1]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[1]));
Q_FDP4EP \_zyaddr_L95_tfiV3_M2_pbcG3_REG[0] ( .CK(_zyM2L94_pbcMevClk9), .CE(n106), .R(n304), .D(_zyixc_port_0_1_s2h[0]), .Q(_zyaddr_L95_tfiV3_M2_pbcG3[0]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[39] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(n304), .Q(_zyixc_port_0_1_h2s[39]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[38] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(n304), .Q(_zyixc_port_0_1_h2s[38]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[37] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(n304), .Q(_zyixc_port_0_1_h2s[37]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[36] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(n304), .Q(_zyixc_port_0_1_h2s[36]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[35] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(n304), .Q(_zyixc_port_0_1_h2s[35]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[34] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(n304), .Q(_zyixc_port_0_1_h2s[34]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[33] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(n304), .Q(_zyixc_port_0_1_h2s[33]));
Q_FDP4EP \_zyixc_port_0_1_h2s_REG[32] ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(_zyresponse_L97_tfiV5_M2_pbcG5), .Q(_zyixc_port_0_1_h2s[32]));
Q_INV U827 ( .A(_zyixc_port_0_1_ack), .Z(n322));
Q_FDP4EP _zyixc_port_0_1_ack_REG  ( .CK(_zyM2L94_pbcMevClk9), .CE(n105), .R(n304), .D(n322), .Q(_zyixc_port_0_1_ack));
Q_FDP4EP _zyresponse_L97_tfiV5_M2_pbcG5_REG  ( .CK(_zyM2L94_pbcMevClk9), .CE(n320), .R(n304), .D(n177), .Q(_zyresponse_L97_tfiV5_M2_pbcG5));
Q_FDP4EP \_zzM2L94_mdxP2_paddr_wr3_REG[19] ( .CK(_zyM2L94_pbcMevClk9), .CE(n115), .R(n304), .D(n135), .Q(_zzM2L94_mdxP2_paddr_wr3[19]));
Q_FDP4EP \_zzM2L94_mdxP2_paddr_wr3_REG[18] ( .CK(_zyM2L94_pbcMevClk9), .CE(n115), .R(n304), .D(n136), .Q(_zzM2L94_mdxP2_paddr_wr3[18]));
Q_FDP4EP \_zzM2L94_mdxP2_paddr_wr3_REG[17] ( .CK(_zyM2L94_pbcMevClk9), .CE(n115), .R(n304), .D(n137), .Q(_zzM2L94_mdxP2_paddr_wr3[17]));
Q_FDP4EP \_zzM2L94_mdxP2_paddr_wr3_REG[16] ( .CK(_zyM2L94_pbcMevClk9), .CE(n115), .R(n304), .D(n138), .Q(_zzM2L94_mdxP2_paddr_wr3[16]));
Q_FDP4EP \_zzM2L94_mdxP2_paddr_wr3_REG[15] ( .CK(_zyM2L94_pbcMevClk9), .CE(n115), .R(n304), .D(n139), .Q(_zzM2L94_mdxP2_paddr_wr3[15]));
Q_FDP4EP \_zzM2L94_mdxP2_paddr_wr3_REG[14] ( .CK(_zyM2L94_pbcMevClk9), .CE(n115), .R(n304), .D(n140), .Q(_zzM2L94_mdxP2_paddr_wr3[14]));
Q_FDP4EP \_zzM2L94_mdxP2_paddr_wr3_REG[13] ( .CK(_zyM2L94_pbcMevClk9), .CE(n115), .R(n304), .D(n141), .Q(_zzM2L94_mdxP2_paddr_wr3[13]));
Q_FDP4EP \_zzM2L94_mdxP2_paddr_wr3_REG[12] ( .CK(_zyM2L94_pbcMevClk9), .CE(n115), .R(n304), .D(n142), .Q(_zzM2L94_mdxP2_paddr_wr3[12]));
Q_FDP4EP \_zzM2L94_mdxP2_paddr_wr3_REG[11] ( .CK(_zyM2L94_pbcMevClk9), .CE(n115), .R(n304), .D(n143), .Q(_zzM2L94_mdxP2_paddr_wr3[11]));
Q_FDP4EP \_zzM2L94_mdxP2_paddr_wr3_REG[10] ( .CK(_zyM2L94_pbcMevClk9), .CE(n115), .R(n304), .D(n144), .Q(_zzM2L94_mdxP2_paddr_wr3[10]));
Q_FDP4EP \_zzM2L94_mdxP2_paddr_wr3_REG[9] ( .CK(_zyM2L94_pbcMevClk9), .CE(n115), .R(n304), .D(n145), .Q(_zzM2L94_mdxP2_paddr_wr3[9]));
Q_FDP4EP \_zzM2L94_mdxP2_paddr_wr3_REG[8] ( .CK(_zyM2L94_pbcMevClk9), .CE(n115), .R(n304), .D(n146), .Q(_zzM2L94_mdxP2_paddr_wr3[8]));
Q_FDP4EP \_zzM2L94_mdxP2_paddr_wr3_REG[7] ( .CK(_zyM2L94_pbcMevClk9), .CE(n115), .R(n304), .D(n147), .Q(_zzM2L94_mdxP2_paddr_wr3[7]));
Q_FDP4EP \_zzM2L94_mdxP2_paddr_wr3_REG[6] ( .CK(_zyM2L94_pbcMevClk9), .CE(n115), .R(n304), .D(n148), .Q(_zzM2L94_mdxP2_paddr_wr3[6]));
Q_FDP4EP \_zzM2L94_mdxP2_paddr_wr3_REG[5] ( .CK(_zyM2L94_pbcMevClk9), .CE(n115), .R(n304), .D(n149), .Q(_zzM2L94_mdxP2_paddr_wr3[5]));
Q_FDP4EP \_zzM2L94_mdxP2_paddr_wr3_REG[4] ( .CK(_zyM2L94_pbcMevClk9), .CE(n115), .R(n304), .D(n150), .Q(_zzM2L94_mdxP2_paddr_wr3[4]));
Q_FDP4EP \_zzM2L94_mdxP2_paddr_wr3_REG[3] ( .CK(_zyM2L94_pbcMevClk9), .CE(n115), .R(n304), .D(n151), .Q(_zzM2L94_mdxP2_paddr_wr3[3]));
Q_FDP4EP \_zzM2L94_mdxP2_paddr_wr3_REG[2] ( .CK(_zyM2L94_pbcMevClk9), .CE(n115), .R(n304), .D(n152), .Q(_zzM2L94_mdxP2_paddr_wr3[2]));
Q_FDP4EP \_zzM2L94_mdxP2_paddr_wr3_REG[1] ( .CK(_zyM2L94_pbcMevClk9), .CE(n115), .R(n304), .D(n153), .Q(_zzM2L94_mdxP2_paddr_wr3[1]));
Q_FDP4EP \_zzM2L94_mdxP2_paddr_wr3_REG[0] ( .CK(_zyM2L94_pbcMevClk9), .CE(n115), .R(n304), .D(n154), .Q(_zzM2L94_mdxP2_paddr_wr3[0]));
Q_FDP4EP \_zzM2L94_mdxP2_bus_timer_wr4_REG[7] ( .CK(_zyM2L94_pbcMevClk9), .CE(n117), .R(n304), .D(n155), .Q(_zzM2L94_mdxP2_bus_timer_wr4[7]));
Q_FDP4EP \_zzM2L94_mdxP2_bus_timer_wr4_REG[6] ( .CK(_zyM2L94_pbcMevClk9), .CE(n117), .R(n304), .D(n156), .Q(_zzM2L94_mdxP2_bus_timer_wr4[6]));
Q_FDP4EP \_zzM2L94_mdxP2_bus_timer_wr4_REG[5] ( .CK(_zyM2L94_pbcMevClk9), .CE(n117), .R(n304), .D(n157), .Q(_zzM2L94_mdxP2_bus_timer_wr4[5]));
Q_FDP4EP \_zzM2L94_mdxP2_bus_timer_wr4_REG[4] ( .CK(_zyM2L94_pbcMevClk9), .CE(n117), .R(n304), .D(n158), .Q(_zzM2L94_mdxP2_bus_timer_wr4[4]));
Q_FDP4EP \_zzM2L94_mdxP2_bus_timer_wr4_REG[3] ( .CK(_zyM2L94_pbcMevClk9), .CE(n117), .R(n304), .D(n159), .Q(_zzM2L94_mdxP2_bus_timer_wr4[3]));
Q_FDP4EP \_zzM2L94_mdxP2_bus_timer_wr4_REG[2] ( .CK(_zyM2L94_pbcMevClk9), .CE(n117), .R(n304), .D(n160), .Q(_zzM2L94_mdxP2_bus_timer_wr4[2]));
Q_FDP4EP \_zzM2L94_mdxP2_bus_timer_wr4_REG[1] ( .CK(_zyM2L94_pbcMevClk9), .CE(n117), .R(n304), .D(n161), .Q(_zzM2L94_mdxP2_bus_timer_wr4[1]));
Q_FDP4EP \_zzM2L94_mdxP2_bus_timer_wr4_REG[0] ( .CK(_zyM2L94_pbcMevClk9), .CE(n117), .R(n304), .D(n162), .Q(_zzM2L94_mdxP2_bus_timer_wr4[0]));
Q_FDP4EP _zyM2L94_pbcCapEn5_REG  ( .CK(_zyM2L94_pbcMevClk9), .CE(n104), .R(n304), .D(n107), .Q(_zyM2L94_pbcCapEn5));
Q_FDP4EP _zyM2L104_pbcCapEn6_REG  ( .CK(_zyM2L94_pbcMevClk9), .CE(n103), .R(n304), .D(n108), .Q(_zyM2L104_pbcCapEn6));
Q_FDP4EP _zyM2L110_pbcCapEn7_REG  ( .CK(_zyM2L94_pbcMevClk9), .CE(n102), .R(n304), .D(n116), .Q(_zyM2L110_pbcCapEn7));
Q_INV U861 ( .A(n123), .Z(n323));
Q_FDP4EP _zyM2L121_pbcCapEn8_REG  ( .CK(_zyM2L94_pbcMevClk9), .CE(n323), .R(n304), .D(n109), .Q(_zyM2L121_pbcCapEn8));
Q_FDP4EP \_zyM2L94_pbcFsm3_s_REG[1] ( .CK(_zyM2L94_pbcMevClk9), .CE(n101), .R(n304), .D(n134), .Q(_zyM2L94_pbcFsm3_s[1]));
Q_INV U864 ( .A(_zyM2L94_pbcFsm3_s[1]), .Z(n127));
Q_FDP4EP \_zyM2L94_pbcFsm3_s_REG[0] ( .CK(_zyM2L94_pbcMevClk9), .CE(n101), .R(n304), .D(n110), .Q(_zyM2L94_pbcFsm3_s[0]));
Q_INV U866 ( .A(_zyM2L94_pbcFsm3_s[0]), .Z(n108));
Q_FDP4EP _zzM2L94_mdxP2_psel_wr0_REG  ( .CK(_zyM2L94_pbcMevClk9), .CE(n115), .R(n304), .D(n114), .Q(_zzM2L94_mdxP2_psel_wr0));
Q_FDP4EP _zzM2L94_mdxP2_penable_wr1_REG  ( .CK(_zyM2L94_pbcMevClk9), .CE(n113), .R(n304), .D(n112), .Q(_zzM2L94_mdxP2_penable_wr1));
Q_FDP4EP _zyM2L94_pbcEn11_REG  ( .CK(_zyM2L94_pbcMevClk9), .CE(n117), .R(n304), .D(n118), .Q(_zyM2L94_pbcEn11));
Q_FDP4EP \_zzM2_bcBehEval_REG[31] ( .CK(_zzM2_bcBehEvalClk), .CE(n26), .R(n304), .D(_zzM2_bcBehHalt), .Q(_zzM2_bcBehEval[31]));
Q_INV U871 ( .A(_zzM2_bcBehEval[30]), .Z(n324));
Q_FDP4EP \_zzM2_bcBehEval_REG[30] ( .CK(_zzM2_bcBehEvalClk), .CE(n2), .R(n304), .D(n324), .Q(_zzM2_bcBehEval[30]));
Q_FDP4EP \_zzM2_bcBehEval_REG[29] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n28), .Q(_zzM2_bcBehEval[29]));
Q_FDP4EP \_zzM2_bcBehEval_REG[28] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n30), .Q(_zzM2_bcBehEval[28]));
Q_FDP4EP \_zzM2_bcBehEval_REG[27] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n32), .Q(_zzM2_bcBehEval[27]));
Q_FDP4EP \_zzM2_bcBehEval_REG[26] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n34), .Q(_zzM2_bcBehEval[26]));
Q_FDP4EP \_zzM2_bcBehEval_REG[25] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n36), .Q(_zzM2_bcBehEval[25]));
Q_FDP4EP \_zzM2_bcBehEval_REG[24] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n38), .Q(_zzM2_bcBehEval[24]));
Q_FDP4EP \_zzM2_bcBehEval_REG[23] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n40), .Q(_zzM2_bcBehEval[23]));
Q_FDP4EP \_zzM2_bcBehEval_REG[22] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n42), .Q(_zzM2_bcBehEval[22]));
Q_FDP4EP \_zzM2_bcBehEval_REG[21] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n44), .Q(_zzM2_bcBehEval[21]));
Q_FDP4EP \_zzM2_bcBehEval_REG[20] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n46), .Q(_zzM2_bcBehEval[20]));
Q_FDP4EP \_zzM2_bcBehEval_REG[19] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n48), .Q(_zzM2_bcBehEval[19]));
Q_FDP4EP \_zzM2_bcBehEval_REG[18] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n50), .Q(_zzM2_bcBehEval[18]));
Q_FDP4EP \_zzM2_bcBehEval_REG[17] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n52), .Q(_zzM2_bcBehEval[17]));
Q_FDP4EP \_zzM2_bcBehEval_REG[16] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n54), .Q(_zzM2_bcBehEval[16]));
Q_FDP4EP \_zzM2_bcBehEval_REG[15] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n56), .Q(_zzM2_bcBehEval[15]));
Q_FDP4EP \_zzM2_bcBehEval_REG[14] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n58), .Q(_zzM2_bcBehEval[14]));
Q_FDP4EP \_zzM2_bcBehEval_REG[13] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n60), .Q(_zzM2_bcBehEval[13]));
Q_FDP4EP \_zzM2_bcBehEval_REG[12] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n62), .Q(_zzM2_bcBehEval[12]));
Q_FDP4EP \_zzM2_bcBehEval_REG[11] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n64), .Q(_zzM2_bcBehEval[11]));
Q_FDP4EP \_zzM2_bcBehEval_REG[10] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n66), .Q(_zzM2_bcBehEval[10]));
Q_FDP4EP \_zzM2_bcBehEval_REG[9] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n68), .Q(_zzM2_bcBehEval[9]));
Q_FDP4EP \_zzM2_bcBehEval_REG[8] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n70), .Q(_zzM2_bcBehEval[8]));
Q_FDP4EP \_zzM2_bcBehEval_REG[7] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n72), .Q(_zzM2_bcBehEval[7]));
Q_FDP4EP \_zzM2_bcBehEval_REG[6] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n74), .Q(_zzM2_bcBehEval[6]));
Q_FDP4EP \_zzM2_bcBehEval_REG[5] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n76), .Q(_zzM2_bcBehEval[5]));
Q_FDP4EP \_zzM2_bcBehEval_REG[4] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n78), .Q(_zzM2_bcBehEval[4]));
Q_FDP4EP \_zzM2_bcBehEval_REG[3] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n80), .Q(_zzM2_bcBehEval[3]));
Q_FDP4EP \_zzM2_bcBehEval_REG[2] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n82), .Q(_zzM2_bcBehEval[2]));
Q_FDP4EP \_zzM2_bcBehEval_REG[1] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n84), .Q(_zzM2_bcBehEval[1]));
Q_INV U902 ( .A(_zzM2_bcBehEval[0]), .Z(n325));
Q_FDP4EP \_zzM2_bcBehEval_REG[0] ( .CK(_zzM2_bcBehEvalClk), .CE(n25), .R(n304), .D(n325), .Q(_zzM2_bcBehEval[0]));
// pragma CVASTRPROP MODULE HDLICE PROP_RANOFF TRUE
endmodule
