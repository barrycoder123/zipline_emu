// xc_work/v/2n.sv
// /home/ibarry/Project-Zipline-master/dv/KME/run/kme_tb.sv:10
// NOTE: This file corresponds to a module in the Hardware/DUT partition.
`timescale 1ns/1ns
module kme_tb;
// external : apb_xactor.read (resolved )  (task)  
// external : apb_xactor.write (resolved )  (task)  
// external : apb_xactor._zyL94_iscX1c0_s (resolved )  (var)  
// external : apb_xactor._zyL94_iscX1c0_f (resolved )  (var)  
// external : apb_xactor._zyL94_iscX1c0_i0 (resolved )  (var)  
// external : apb_xactor._zyL94_iscX1c0_o1 (resolved )  (var)  
// external : apb_xactor._zyL94_iscX1c0_o2 (resolved )  (var)  
// external : apb_xactor._zyL61_iscX2c0_s (resolved )  (var)  
// external : apb_xactor._zyL61_iscX2c0_f (resolved )  (var)  
// external : apb_xactor._zyL61_iscX2c0_i0 (resolved )  (var)  
// external : apb_xactor._zyL61_iscX2c0_i1 (resolved )  (var)  
// external : apb_xactor._zyL61_iscX2c0_o2 (resolved )  (var)  
// exported object:  (scope) tb_task 
// exported object:  (var) my_clk (R)  
// exported object:  (var) _zyixc_port_0_0_isf (R)  
// exported object:  (var) _zyixc_port_0_0_osf (R)  
// exported object:  (var) _zyL94_iscX1c0_s (R)  
// exported object:  (var) _zyL94_iscX1c0_f (R)  
// exported object:  (var) _zyL94_iscX1c0_i0 (R)  
// exported object:  (var) _zyL94_iscX1c0_o1 (R)  
// exported object:  (var) _zyL94_iscX1c0_o2 (R)  
// exported object:  (var) _zyL61_iscX2c0_s (R)  
// exported object:  (var) _zyL61_iscX2c0_f (R)  
// exported object:  (var) _zyL61_iscX2c0_i0 (R)  
// exported object:  (var) _zyL61_iscX2c0_i1 (R)  
// exported object:  (var) _zyL61_iscX2c0_o2 (R)  
// exported object:  (var) _zyGfifo_mod2_dflt_ci (R)  
// exported object:  (var) _zyGfifo_mod2_dflt_co (R)  
reg [279:0] testname ;
reg [279:0] seed ;
reg [31:0] initial_seed ;
int error_cntr;
string fsdbFilename;
logic clk;
logic rst_n;
logic kme_ib_tready;
logic [0:0] kme_ib_tid ;
logic [63:0] kme_ib_tdata ;
logic [7:0] kme_ib_tstrb ;
logic [7:0] kme_ib_tuser ;
logic kme_ib_tvalid;
logic kme_ib_tlast;
logic kme_ob_tready;
logic [0:0] kme_ob_tid ;
logic [63:0] kme_ob_tdata ;
logic [7:0] kme_ob_tstrb ;
logic [7:0] kme_ob_tuser ;
logic kme_ob_tvalid;
logic kme_ob_tlast;
logic [19:0] kme_apb_paddr ;
logic kme_apb_psel;
logic kme_apb_penable;
logic kme_apb_pwrite;
logic [31:0] kme_apb_pwdata ;
logic [31:0] kme_apb_prdata ;
logic kme_apb_pready;
logic kme_apb_pslverr;
logic my_clk;
logic config_done = 0;
bit [7:0] tstrb_ib ;
bit [63:0] tdata_ib ;
bit [31:0] tuser_string_ib ;
bit [31:0] str_get_ib ;
reg [24:0] user_string_ib  = 25'b0;
int retval_ib;
logic ready_ib = 0;
logic saw_mega;
logic saw_guid_tlv;
logic have_guid_tlv;
int mega_tlv_word_count;
bit [7:0] tstrb_ob ;
bit [63:0] tdata_ob ;
bit [31:0] tuser_string_ob ;
reg [24:0] user_string_ob ;
bit [31:0] str_get_ob ;
int retval_ob;
logic ready_ob = 0;
reg [7:0] tuser ;
reg tlast;
logic saw_cqe;
logic saw_stats;
logic ignore_compare_result;
integer watchdog_timer;
reg [31:0] returned_data ;
reg response;
bit [7:0] operation ;
bit [31:0] address ;
bit [31:0] data ;
int retval;
logic config_ready = 0;
integer _zz_58_258_2;
integer _zz_58_264_3;
wire  _zy_simnet_kme_apb_psel_0_w$;
wire  _zy_simnet_kme_apb_penable_1_w$;
wire  [0:19] _zy_simnet_kme_apb_paddr_2_w$ ;
wire  [0:31] _zy_simnet_kme_apb_pwdata_3_w$ ;
wire  _zy_simnet_kme_apb_pwrite_4_w$;
wire  _zy_simnet_clk_5_w$;
wire  _zy_simnet_rst_n_6_w$;
wire  [0:31] _zy_simnet_kme_apb_prdata_7_w$ ;
wire  _zy_simnet_kme_apb_pready_8_w$;
wire  _zy_simnet_kme_apb_pslverr_9_w$;
wire  _zy_simnet_dio_10;
wire  _zy_simnet_kme_ib_tready_11_w$;
wire  _zy_simnet_kme_ob_tvalid_12_w$;
wire  _zy_simnet_kme_ob_tlast_13_w$;
wire  _zy_simnet_kme_ob_tid_14_w$;
wire  [0:7] _zy_simnet_kme_ob_tstrb_15_w$ ;
wire  [0:7] _zy_simnet_kme_ob_tuser_16_w$ ;
wire  [0:63] _zy_simnet_kme_ob_tdata_17_w$ ;
wire  [0:31] _zy_simnet_kme_apb_prdata_18_w$ ;
wire  _zy_simnet_kme_apb_pready_19_w$;
wire  _zy_simnet_kme_apb_pslverr_20_w$;
wire  _zy_simnet_dio_21;
wire  _zy_simnet_clk_22_w$;
wire  _zy_simnet_rst_n_23_w$;
wire  _zy_simnet_cio_24;
wire  _zy_simnet_cio_25;
wire  _zy_simnet_cio_26;
wire  _zy_simnet_cio_27;
wire  _zy_simnet_cio_28;
wire  _zy_simnet_cio_29;
wire  _zy_simnet_cio_30;
wire  _zy_simnet_cio_31;
wire  _zy_simnet_kme_ib_tvalid_32_w$;
wire  _zy_simnet_kme_ib_tlast_33_w$;
wire  _zy_simnet_kme_ib_tid_34_w$;
wire  [0:7] _zy_simnet_kme_ib_tstrb_35_w$ ;
wire  [0:7] _zy_simnet_kme_ib_tuser_36_w$ ;
wire  [0:63] _zy_simnet_kme_ib_tdata_37_w$ ;
wire  _zy_simnet_kme_ob_tready_38_w$;
wire  [0:15] _zy_simnet_kme_apb_paddr_39_w$ ;
wire  _zy_simnet_kme_apb_psel_40_w$;
wire  _zy_simnet_kme_apb_penable_41_w$;
wire  _zy_simnet_kme_apb_pwrite_42_w$;
wire  [0:31] _zy_simnet_kme_apb_pwdata_43_w$ ;
bit [71:0] _zygsfis_get_config_data_fifo [0:31];
bit [4:0] _zygsfis_get_config_data_wptr ;
bit [4:0] _zygsfis_get_config_data_rptr ;
bit [4:0] _zygsfis_get_config_data_req ;
bit [4:0] _zygsfis_get_config_data_ack ;
bit _zygsfis_get_config_data_eos;
bit [4:0] _zygsfis_get_config_data_space ;
bit [135:0] _zygsfis_ib_service_data_fifo [0:31];
bit [4:0] _zygsfis_ib_service_data_wptr ;
bit [4:0] _zygsfis_ib_service_data_rptr ;
bit [4:0] _zygsfis_ib_service_data_req ;
bit [4:0] _zygsfis_ib_service_data_ack ;
bit _zygsfis_ib_service_data_eos;
bit [4:0] _zygsfis_ib_service_data_space ;
bit [135:0] _zygsfis_ob_service_data_fifo [0:31];
bit [4:0] _zygsfis_ob_service_data_wptr ;
bit [4:0] _zygsfis_ob_service_data_rptr ;
bit [4:0] _zygsfis_ob_service_data_req ;
bit [4:0] _zygsfis_ob_service_data_ack ;
bit _zygsfis_ob_service_data_eos;
bit [4:0] _zygsfis_ob_service_data_space ;
wire  _zyixc_port_0_0_s2h;
wire  _zyixc_port_0_0_s2hW;
bit _zyixc_port_0_0_req;
bit _zyixc_port_0_0_ack;
bit _zyixc_port_0_0_isf;
bit _zyixc_port_0_0_osf;
bit [21:0] _zySfifoF0_get_config_data_zyackf_tid ;
wire  _zySfifoF0_call;
wire  _zySfifoF0_fen;
wire  [31:0] _zySfifoF0_iarg ;
wire  [511:0] _zyGfifo_SiData ;
wire  [21:0] _zyGfifo_StId ;
wire  [511:0] _zyGfifo_SoData ;
wire  _zyGfifo_SoDataEn;
wire  [3:0] _zyGfifo_SoDataLen ;
bit [21:0] _zySfifoF1_get_config_data_zyputf_tid ;
wire  _zySfifoF1_call;
wire  _zySfifoF1_fen;
wire  [71:0] _zySfifoF1_iarg ;
bit [21:0] _zySfifoF2_ib_service_data_zyackf_tid ;
wire  _zySfifoF2_call;
wire  _zySfifoF2_fen;
wire  [31:0] _zySfifoF2_iarg ;
bit [21:0] _zySfifoF3_ib_service_data_zyputf_tid ;
wire  _zySfifoF3_call;
wire  _zySfifoF3_fen;
wire  [135:0] _zySfifoF3_iarg ;
bit [21:0] _zySfifoF4_ob_service_data_zyackf_tid ;
wire  _zySfifoF4_call;
wire  _zySfifoF4_fen;
wire  [31:0] _zySfifoF4_iarg ;
bit [21:0] _zySfifoF5_ob_service_data_zyputf_tid ;
wire  _zySfifoF5_call;
wire  _zySfifoF5_fen;
wire  [135:0] _zySfifoF5_iarg ;
reg _zyL94_iscX1c0_s;
wire  _zyL94_iscX1c0_f;
reg _zyL94_iscX1c0_n;
reg [63:0]  _zyL94_iscX1c0_i0;
wire [31:0]  _zyL94_iscX1c0_o1;
wire  _zyL94_iscX1c0_o2;
reg _zyL61_iscX2c0_s;
wire  _zyL61_iscX2c0_f;
reg _zyL61_iscX2c0_n;
reg [63:0]  _zyL61_iscX2c0_i0;
reg [31:0]  _zyL61_iscX2c0_i1;
wire  _zyL61_iscX2c0_o2;
logic [24:0] _zyL372_tfiRv5 ;
logic [7:0] _zyL406_tfiRv6 ;
logic [24:0] _zyL443_tfiRv7 ;
logic [7:0] _zyL462_tfiRv8 ;
reg [279:0] _zyictd_sysfunc_36_L258_0 ;
const integer _zyictd_sysfunc_36_L258_1 = $value$plusargs("SEED=%d",_zyictd_sysfunc_36_L258_0);
const integer _zyictd_sysfunc_11_L257_2 = $test$plusargs("SEED");
reg [279:0] _zyictd_sysfunc_36_L264_3 ;
const integer _zyictd_sysfunc_36_L264_4 = $value$plusargs("TESTNAME=%s",_zyictd_sysfunc_36_L264_3);
const integer _zyictd_sysfunc_11_L263_5 = $test$plusargs("TESTNAME");
bit _zyictd_finish_L320_0;
bit _zyictd_finish_L338_1;
bit _zyictd_finish_L454_2;
wire  _zyictd_finish_mgr;
int _zyL326_tfiRv17;
int _zyL370_tfiRv18;
int _zyL441_tfiRv19;
wire  _zyGfifo_mod2_dflt_ci;
wire  _zyGfifo_mod2_dflt_co;
wire  [26:0] _zyGfifo_dflt_ci ;
wire  [26:0] _zyGfifo_dflt_co ;
bit [0:0] _zyGfifo_mod2_simData ;
bit _zyGfifo__gfdL435_34_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL435_34_P0_m2_cbid ;
bit _zyGfifo__gfdL513_33_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL513_33_P0_m2_cbid ;
bit _zyGfifo__gfdL316_32_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL316_32_P0_m2_cbid ;
bit _zyGfifo__gfdL318_31_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL318_31_P0_m2_cbid ;
bit _zyGfifo_get_config_data_2_zyprefetch_m2_gfOff;
bit [19:0] _zyGfifo_get_config_data_2_zyprefetch_m2_cbid ;
bit _zyGfifo__gfdL327_30_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL327_30_P0_m2_cbid ;
bit _zyGfifo__gfdL330_29_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL330_29_P0_m2_cbid ;
bit _zyGfifo__gfdL334_28_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL334_28_P0_m2_cbid ;
bit _zyGfifo__gfdL336_27_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL336_27_P0_m2_cbid ;
bit _zyGfifo__gfdL341_26_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL341_26_P0_m2_cbid ;
bit _zyGfifo__gfdL351_25_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL351_25_P0_m2_cbid ;
bit _zyGfifo_ib_service_data_2_zyprefetch_m2_gfOff;
bit [19:0] _zyGfifo_ib_service_data_2_zyprefetch_m2_cbid ;
bit _zyGfifo__gfdL519_24_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL519_24_P0_m2_cbid ;
bit _zyGfifo__gfdL522_23_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL522_23_P0_m2_cbid ;
bit _zyGfifo__gfdL373_22_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL373_22_P0_m2_cbid ;
bit _zyGfifo__gfdL375_21_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL375_21_P0_m2_cbid ;
bit _zyGfifo__gfdL381_20_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL381_20_P0_m2_cbid ;
bit _zyGfifo__gfdL390_19_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL390_19_P0_m2_cbid ;
bit _zyGfifo__gfdL530_18_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL530_18_P0_m2_cbid ;
bit _zyGfifo__gfdL412_17_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL412_17_P0_m2_cbid ;
bit _zyGfifo_ob_service_data_2_zyprefetch_m2_gfOff;
bit [19:0] _zyGfifo_ob_service_data_2_zyprefetch_m2_cbid ;
bit _zyGfifo__gfdL519_16_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL519_16_P0_m2_cbid ;
bit _zyGfifo__gfdL522_15_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL522_15_P0_m2_cbid ;
bit _zyGfifo__gfdL444_14_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL444_14_P0_m2_cbid ;
bit _zyGfifo__gfdL446_13_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL446_13_P0_m2_cbid ;
bit _zyGfifo__gfdL460_12_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL460_12_P0_m2_cbid ;
bit _zyGfifo__gfdL530_11_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL530_11_P0_m2_cbid ;
bit _zyGfifo__gfdL480_10_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL480_10_P0_m2_cbid ;
bit _zyGfifo__gfdL482_9_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL482_9_P0_m2_cbid ;
bit _zyGfifo__gfdL487_8_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL487_8_P0_m2_cbid ;
bit _zyGfifo__gfdL491_7_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL491_7_P0_m2_cbid ;
bit _zyGfifo__gfdL496_6_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL496_6_P0_m2_cbid ;
bit _zyGfifo__gfdL265_5_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL265_5_P0_m2_cbid ;
bit _zyGfifo__gfdL268_4_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL268_4_P0_m2_cbid ;
bit _zyGfifo__gfdL271_3_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL271_3_P0_m2_cbid ;
bit _zyGfifo__gfdL276_2_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL276_2_P0_m2_cbid ;
bit _zyGfifo__gfdL289_1_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL289_1_P0_m2_cbid ;
bit _zyGfifo__gfdL365_0_P0_m2_gfOff;
bit [19:0] _zyGfifo__gfdL365_0_P0_m2_cbid ;
bit _zyGfifoF0_L435_req_0;
wire  _zyGfifo_SGFtsReq;
wire  [19:0] _zyGfifo_SGFcbid ;
wire  [11:0] _zyGfifo_SGFlen ;
wire  [511:0] _zyGfifo_SGFidata ;
wire  _zyGfifo_SGFfull;
wire  _zyGfifo_SLBreq;
wire  [3:0] _zyGfifo_SLBrd ;
wire  [3:0] _zyGfifo_SLBwr ;
wire  _zyGfifo_SLBfull;
wire  _zyGfifo_SRtkin;
bit _zyGfifoF1_L513_req_0;
bit _zyGfifoF0_L312_s2_req_0;
bit [279:0] _zyGfifoF0_L312_s2_data_0 ;
bit [19:0] _zyGfifoF0_L312_s2_cbid_0 ;
bit _zyGfifoF0_L324_s3_req_1;
bit [95:0] _zyGfifoF0_L324_s3_data_1 ;
bit [19:0] _zyGfifoF0_L324_s3_cbid_1 ;
bit [11:0] _zyGfifoF0_L324_s3_len_1 ;
bit _zyGfifoF1_L324_s2_req_2;
bit [31:0] _zyGfifoF1_L324_s2_data_2 ;
bit [19:0] _zyGfifoF1_L324_s2_cbid_2 ;
bit _zyGfifoF2_L324_s2_req_3;
bit [71:0] _zyGfifoF2_L324_s2_data_3 ;
bit [19:0] _zyGfifoF2_L324_s2_cbid_3 ;
bit [11:0] _zyGfifoF2_L324_s2_len_3 ;
bit _zyGfifoF11_L207_req_0;
bit [31:0] _zyGfifoF11_L207_data_0 ;
bit _zyGfifoF0_L368_s2_req_4;
bit [19:0] _zyGfifoF0_L368_s2_cbid_4 ;
bit _zyGfifoF14_L373_req_0;
bit [31:0] _zyGfifoF14_L373_data_0 ;
bit _zyGfifoF15_L375_req_0;
bit [135:0] _zyGfifoF15_L375_data_0 ;
bit _zyGfifoF16_L381_req_0;
bit _zyGfifoF17_L390_req_0;
bit [63:0] _zyGfifoF17_L390_data_0 ;
bit _zyGfifoF18_L530_req_0;
bit [31:0] _zyGfifoF18_L530_data_0 ;
bit _zyGfifoF19_L412_req_0;
bit [7:0] _zyGfifoF19_L412_data_0 ;
bit _zyGfifoF20_L209_req_0;
bit [31:0] _zyGfifoF20_L209_data_0 ;
bit _zyGfifoF0_L439_s2_req_5;
bit [19:0] _zyGfifoF0_L439_s2_cbid_5 ;
bit _zyGfifoF23_L444_req_0;
bit [31:0] _zyGfifoF23_L444_data_0 ;
bit _zyGfifoF24_L446_req_0;
bit [135:0] _zyGfifoF24_L446_data_0 ;
bit _zyGfifoF25_L460_req_0;
bit [63:0] _zyGfifoF25_L460_data_0 ;
bit _zyGfifoF26_L530_req_0;
bit [31:0] _zyGfifoF26_L530_data_0 ;
bit _zyGfifoF27_L480_req_0;
bit [7:0] _zyGfifoF27_L480_data_0 ;
bit _zyGfifoF28_L482_req_0;
bit [127:0] _zyGfifoF28_L482_data_0 ;
bit _zyGfifoF29_L487_req_0;
bit [15:0] _zyGfifoF29_L487_data_0 ;
bit _zyGfifoF30_L491_req_0;
bit [15:0] _zyGfifoF30_L491_data_0 ;
bit _zyGfifoF31_L496_req_0;
bit [15:0] _zyGfifoF31_L496_data_0 ;
bit _zyGfifoF0_L253_s4_req_6;
bit [559:0] _zyGfifoF0_L253_s4_data_6 ;
bit [19:0] _zyGfifoF0_L253_s4_cbid_6 ;
bit [11:0] _zyGfifoF0_L253_s4_len_6 ;
bit _zyGfifoF1_L253_s2_req_7;
bit [19:0] _zyGfifoF1_L253_s2_cbid_7 ;
bit [7:0] _zyoperation_L206_tfiV0_M2_pbcG0 ;
bit [31:0] _zyaddress_L206_tfiV1_M2_pbcG1 ;
bit [31:0] _zydata_L206_tfiV2_M2_pbcG2 ;
int _zyxr_L206_tfiV3_M2_pbcG3;
reg signed [31:0]  _zyM2L273_pbcT0;
reg signed [31:0]  _zyM2L286_pbcT1;
reg signed [31:0]  _zyM2L292_pbcT2;
reg signed [31:0]  _zyM2L299_pbcT3;
reg _zyM2L324_pbcCapEn0;
reg _zyM2L333_pbcCapEn1;
reg _zyM2L349_pbcCapEn2;
reg _zyM2L355_pbcCapEn3;
wire  _zyM2L324_pbcMevClk4;
wire  _zyM2L324_pbcReq4;
wire  _zyM2L324_pbcBusy4;
wire  _zyM2L324_pbcWait4;
reg _zyM2L253_pbcCapEn5;
reg _zyM2L274_pbcCapEn6;
reg _zyM2L287_pbcCapEn7;
reg _zyM2L293_pbcCapEn8;
reg _zyM2L295_pbcCapEn9;
reg _zyM2L364_pbcCapEn10;
reg _zyM2L300_pbcCapEn11;
wire  _zyM2L253_pbcMevClk12;
wire  _zyM2L253_pbcReq12;
wire  _zyM2L253_pbcBusy12;
wire  _zyM2L253_pbcWait12;
reg [2:0]  _zyM2L324_pbcFsm0_s;
reg _zyM2L324_pbcEn13;
reg [2:0]  _zyM2L253_pbcFsm2_s;
reg _zyM2L253_pbcEn14;
reg [0:0]  _zyL306_meState0;
reg [0:0]  _zyL312_meState2;
reg [0:0]  _zyL368_meState4;
reg [1:0]  _zyL439_meState8;
wire  _zyictd_finish_mgr_x$tbc;
// F1, L91
assign  clk = my_clk;
// F1, L99
assign  kme_apb_psel = _zy_simnet_kme_apb_psel_0_w$;
// F1, L100
assign  kme_apb_penable = _zy_simnet_kme_apb_penable_1_w$;
// F1, L101
assign  kme_apb_paddr = _zy_simnet_kme_apb_paddr_2_w$;
// F1, L102
assign  kme_apb_pwdata = _zy_simnet_kme_apb_pwdata_3_w$;
// F1, L103
assign  kme_apb_pwrite = _zy_simnet_kme_apb_pwrite_4_w$;
// F1, L26
assign  _zy_simnet_clk_5_w$ = clk;
// F1, L27
assign  _zy_simnet_rst_n_6_w$ = rst_n;
// F1, L65
assign  _zy_simnet_kme_apb_prdata_7_w$ = kme_apb_prdata;
// F1, L66
assign  _zy_simnet_kme_apb_pready_8_w$ = kme_apb_pready;
// F1, L67
assign  _zy_simnet_kme_apb_pslverr_9_w$ = kme_apb_pslverr;
// F1, L107
assign  kme_ib_tready = _zy_simnet_kme_ib_tready_11_w$;
// F1, L116
assign  kme_ob_tvalid = _zy_simnet_kme_ob_tvalid_12_w$;
// F1, L117
assign  kme_ob_tlast = _zy_simnet_kme_ob_tlast_13_w$;
// F1, L118
assign  kme_ob_tid = _zy_simnet_kme_ob_tid_14_w$;
// F1, L119
assign  kme_ob_tstrb = _zy_simnet_kme_ob_tstrb_15_w$;
// F1, L120
assign  kme_ob_tuser = _zy_simnet_kme_ob_tuser_16_w$;
// F1, L121
assign  kme_ob_tdata = _zy_simnet_kme_ob_tdata_17_w$;
// F1, L186
assign  kme_apb_prdata = _zy_simnet_kme_apb_prdata_18_w$;
// F1, L187
assign  kme_apb_pready = _zy_simnet_kme_apb_pready_19_w$;
// F1, L188
assign  kme_apb_pslverr = _zy_simnet_kme_apb_pslverr_20_w$;
// F1, L26
assign  _zy_simnet_clk_22_w$ = clk;
// F1, L27
assign  _zy_simnet_rst_n_23_w$ = rst_n;
// F1, L192
assign  _zy_simnet_cio_24 = 1'b0;
// F1, L193
assign  _zy_simnet_cio_25 = 1'b0;
// F1, L194
assign  _zy_simnet_cio_26 = 1'b0;
// F1, L196
assign  _zy_simnet_cio_27 = 1'b1;
// F1, L197
assign  _zy_simnet_cio_28 = 1'b0;
// F1, L198
assign  _zy_simnet_cio_29 = 1'b0;
// F1, L201
assign  _zy_simnet_cio_30 = 1'b0;
// F1, L203
assign  _zy_simnet_cio_31 = 1'b0;
// F1, L36
assign  _zy_simnet_kme_ib_tvalid_32_w$ = kme_ib_tvalid;
// F1, L37
assign  _zy_simnet_kme_ib_tlast_33_w$ = kme_ib_tlast;
// F1, L32
assign  _zy_simnet_kme_ib_tid_34_w$ = kme_ib_tid;
// F1, L34
assign  _zy_simnet_kme_ib_tstrb_35_w$ = kme_ib_tstrb;
// F1, L35
assign  _zy_simnet_kme_ib_tuser_36_w$ = kme_ib_tuser;
// F1, L33
assign  _zy_simnet_kme_ib_tdata_37_w$ = kme_ib_tdata;
// F1, L45
assign  _zy_simnet_kme_ob_tready_38_w$ = kme_ob_tready;
// F1, L60
assign  _zy_simnet_kme_apb_paddr_39_w$ = kme_apb_paddr[15:0];
// F1, L61
assign  _zy_simnet_kme_apb_psel_40_w$ = kme_apb_psel;
// F1, L62
assign  _zy_simnet_kme_apb_penable_41_w$ = kme_apb_penable;
// F1, L63
assign  _zy_simnet_kme_apb_pwrite_42_w$ = kme_apb_pwrite;
// F1, L64
assign  _zy_simnet_kme_apb_pwdata_43_w$ = kme_apb_pwdata;
// F1, L10
ixc_mem_call #(0,0,0,0) _zzixc_tfport_0_0 (_zyixc_port_0_0_req,_zyixc_port_0_0_s2h,_zyixc_port_0_0_isf,_zyixc_port_0_0_ack,1'b0,_zyixc_port_0_0_osf,1'b0,1'b0);
// F1, L206
ixc_sfifo_port #(32,0) _zzSfifoF0_L206_p (_zySfifoF0_call,_zySfifoF0_iarg,1'b0,_zySfifoF0_get_config_data_zyackf_tid,_zySfifoF0_fen,_zyGfifo_SiData,_zyGfifo_StId,_zyGfifo_SoData,_zyGfifo_SoDataEn,_zyGfifo_SoDataLen);
// F1, L206
ixc_sfifo_port #(72,0) _zzSfifoF1_L206_p (_zySfifoF1_call,_zySfifoF1_iarg,1'b0,_zySfifoF1_get_config_data_zyputf_tid,_zySfifoF1_fen,_zyGfifo_SiData,_zyGfifo_StId,_zyGfifo_SoData,_zyGfifo_SoDataEn,_zyGfifo_SoDataLen);
// F1, L207
ixc_sfifo_port #(32,0) _zzSfifoF2_L207_p (_zySfifoF2_call,_zySfifoF2_iarg,1'b0,_zySfifoF2_ib_service_data_zyackf_tid,_zySfifoF2_fen,_zyGfifo_SiData,_zyGfifo_StId,_zyGfifo_SoData,_zyGfifo_SoDataEn,_zyGfifo_SoDataLen);
// F1, L207
ixc_sfifo_port #(136,0) _zzSfifoF3_L207_p (_zySfifoF3_call,_zySfifoF3_iarg,1'b0,_zySfifoF3_ib_service_data_zyputf_tid,_zySfifoF3_fen,_zyGfifo_SiData,_zyGfifo_StId,_zyGfifo_SoData,_zyGfifo_SoDataEn,_zyGfifo_SoDataLen);
// F1, L209
ixc_sfifo_port #(32,0) _zzSfifoF4_L209_p (_zySfifoF4_call,_zySfifoF4_iarg,1'b0,_zySfifoF4_ob_service_data_zyackf_tid,_zySfifoF4_fen,_zyGfifo_SiData,_zyGfifo_StId,_zyGfifo_SoData,_zyGfifo_SoDataEn,_zyGfifo_SoDataLen);
// F1, L209
ixc_sfifo_port #(136,0) _zzSfifoF5_L209_p (_zySfifoF5_call,_zySfifoF5_iarg,1'b0,_zySfifoF5_ob_service_data_zyputf_tid,_zySfifoF5_fen,_zyGfifo_SiData,_zyGfifo_StId,_zyGfifo_SoData,_zyGfifo_SoDataEn,_zyGfifo_SoDataLen);
// F1, L10
assign  apb_xactor._zyL94_iscX1c0_s = _zyL94_iscX1c0_s;
// F1, L10
assign  _zyL94_iscX1c0_f = apb_xactor._zyL94_iscX1c0_f;
// F1, L10
assign  apb_xactor._zyL94_iscX1c0_i0[63:0] = _zyL94_iscX1c0_i0;
// F1, L10
assign  _zyL94_iscX1c0_o1 = apb_xactor._zyL94_iscX1c0_o1[31:0];
// F1, L10
assign  _zyL94_iscX1c0_o2 = apb_xactor._zyL94_iscX1c0_o2;
// F1, L10
assign  apb_xactor._zyL61_iscX2c0_s = _zyL61_iscX2c0_s;
// F1, L10
assign  _zyL61_iscX2c0_f = apb_xactor._zyL61_iscX2c0_f;
// F1, L10
assign  apb_xactor._zyL61_iscX2c0_i0[63:0] = _zyL61_iscX2c0_i0;
// F1, L10
assign  apb_xactor._zyL61_iscX2c0_i1[31:0] = _zyL61_iscX2c0_i1;
// F1, L10
assign  _zyL61_iscX2c0_o2 = apb_xactor._zyL61_iscX2c0_o2;
// F1, L10
initial begin
 #(1'b0)
  forever
   @(posedge _zyictd_finish_mgr)
    if (!(xc_top.hwOutInit && 1'b1))
     begin
      xc_top.xcSchPulseQ;
      @(xc_top.pulseQEvent) ;
      _zzictd_finishT_L10_0;
     end
end

// F1, L10
assign  _zyictd_finish_mgr = ((_zyictd_finish_L454_2 | _zyictd_finish_L320_0) | _zyictd_finish_L338_1);
// F1, L435
ixc_gfifo_port #(1,0,1,4,1) _zzGfifoF0_L435_p_0 (_zyGfifo_dflt_co[0],_zyGfifo_dflt_ci[0],_zyGfifoF0_L435_req_0,_zyGfifo__gfdL435_34_P0_m2_cbid,12'b0,1'b0,_zyGfifo_SGFtsReq,_zyGfifo_SGFcbid,_zyGfifo_SGFlen,_zyGfifo_SGFidata,
_zyGfifo_SGFfull,_zyGfifo_SLBreq,_zyGfifo_SLBrd,_zyGfifo_SLBwr,_zyGfifo_SLBfull,_zyGfifo_SRtkin);
// F1, L513
ixc_gfifo_port #(1,0,1,4,1) _zzGfifoF1_L513_p_0 (_zyGfifo_dflt_co[1],_zyGfifo_dflt_ci[1],_zyGfifoF1_L513_req_0,_zyGfifo__gfdL513_33_P0_m2_cbid,12'b0,1'b0,_zyGfifo_SGFtsReq,_zyGfifo_SGFcbid,_zyGfifo_SGFlen,_zyGfifo_SGFidata,
_zyGfifo_SGFfull,_zyGfifo_SLBreq,_zyGfifo_SLBrd,_zyGfifo_SLBwr,_zyGfifo_SLBfull,_zyGfifo_SRtkin);
// F1, L312
ixc_gfifo_port #(280,2,0,4,1) _zzGfifoF0_L312_s2_p_0 (_zyGfifo_dflt_co[2],_zyGfifo_dflt_ci[2],_zyGfifoF0_L312_s2_req_0,_zyGfifoF0_L312_s2_cbid_0,12'b01001,_zyGfifoF0_L312_s2_data_0,_zyGfifo_SGFtsReq,_zyGfifo_SGFcbid,_zyGfifo_SGFlen,_zyGfifo_SGFidata,
_zyGfifo_SGFfull,_zyGfifo_SLBreq,_zyGfifo_SLBrd,_zyGfifo_SLBwr,_zyGfifo_SLBfull,_zyGfifo_SRtkin);
// F1, L324
ixc_gfifo_port #(96,3,1,4,1) _zzGfifoF0_L324_s3_p_1 (_zyGfifo_dflt_co[3],_zyGfifo_dflt_ci[3],_zyGfifoF0_L324_s3_req_1,_zyGfifoF0_L324_s3_cbid_1,_zyGfifoF0_L324_s3_len_1,_zyGfifoF0_L324_s3_data_1,_zyGfifo_SGFtsReq,_zyGfifo_SGFcbid,_zyGfifo_SGFlen,_zyGfifo_SGFidata,
_zyGfifo_SGFfull,_zyGfifo_SLBreq,_zyGfifo_SLBrd,_zyGfifo_SLBwr,_zyGfifo_SLBfull,_zyGfifo_SRtkin);
// F1, L324
ixc_gfifo_port #(32,2,1,4,1) _zzGfifoF1_L324_s2_p_2 (_zyGfifo_dflt_co[4],_zyGfifo_dflt_ci[4],_zyGfifoF1_L324_s2_req_2,_zyGfifoF1_L324_s2_cbid_2,12'b01,_zyGfifoF1_L324_s2_data_2,_zyGfifo_SGFtsReq,_zyGfifo_SGFcbid,_zyGfifo_SGFlen,_zyGfifo_SGFidata,
_zyGfifo_SGFfull,_zyGfifo_SLBreq,_zyGfifo_SLBrd,_zyGfifo_SLBwr,_zyGfifo_SLBfull,_zyGfifo_SRtkin);
// F1, L324
ixc_gfifo_port #(72,3,1,4,1) _zzGfifoF2_L324_s2_p_3 (_zyGfifo_dflt_co[5],_zyGfifo_dflt_ci[5],_zyGfifoF2_L324_s2_req_3,_zyGfifoF2_L324_s2_cbid_3,_zyGfifoF2_L324_s2_len_3,_zyGfifoF2_L324_s2_data_3,_zyGfifo_SGFtsReq,_zyGfifo_SGFcbid,_zyGfifo_SGFlen,_zyGfifo_SGFidata,
_zyGfifo_SGFfull,_zyGfifo_SLBreq,_zyGfifo_SLBrd,_zyGfifo_SLBwr,_zyGfifo_SLBfull,_zyGfifo_SRtkin);
// F1, L207
ixc_gfifo_port #(32,0,0,4,1) _zzGfifoF11_L207_p_0 (_zyGfifo_dflt_co[6],_zyGfifo_dflt_ci[6],_zyGfifoF11_L207_req_0,_zyGfifo_ib_service_data_2_zyprefetch_m2_cbid,12'b01,_zyGfifoF11_L207_data_0,_zyGfifo_SGFtsReq,_zyGfifo_SGFcbid,_zyGfifo_SGFlen,_zyGfifo_SGFidata,
_zyGfifo_SGFfull,_zyGfifo_SLBreq,_zyGfifo_SLBrd,_zyGfifo_SLBwr,_zyGfifo_SLBfull,_zyGfifo_SRtkin);
// F1, L368
ixc_gfifo_port #(1,2,0,4,1) _zzGfifoF0_L368_s2_p_4 (_zyGfifo_dflt_co[7],_zyGfifo_dflt_ci[7],_zyGfifoF0_L368_s2_req_4,_zyGfifoF0_L368_s2_cbid_4,12'b0,1'b0,_zyGfifo_SGFtsReq,_zyGfifo_SGFcbid,_zyGfifo_SGFlen,_zyGfifo_SGFidata,
_zyGfifo_SGFfull,_zyGfifo_SLBreq,_zyGfifo_SLBrd,_zyGfifo_SLBwr,_zyGfifo_SLBfull,_zyGfifo_SRtkin);
// F1, L373
ixc_gfifo_port #(32,0,0,4,1) _zzGfifoF14_L373_p_0 (_zyGfifo_dflt_co[8],_zyGfifo_dflt_ci[8],_zyGfifoF14_L373_req_0,_zyGfifo__gfdL373_22_P0_m2_cbid,12'b01,_zyGfifoF14_L373_data_0,_zyGfifo_SGFtsReq,_zyGfifo_SGFcbid,_zyGfifo_SGFlen,_zyGfifo_SGFidata,
_zyGfifo_SGFfull,_zyGfifo_SLBreq,_zyGfifo_SLBrd,_zyGfifo_SLBwr,_zyGfifo_SLBfull,_zyGfifo_SRtkin);
// F1, L375
ixc_gfifo_port #(136,0,0,4,1) _zzGfifoF15_L375_p_0 (_zyGfifo_dflt_co[9],_zyGfifo_dflt_ci[9],_zyGfifoF15_L375_req_0,_zyGfifo__gfdL375_21_P0_m2_cbid,12'b0101,_zyGfifoF15_L375_data_0,_zyGfifo_SGFtsReq,_zyGfifo_SGFcbid,_zyGfifo_SGFlen,_zyGfifo_SGFidata,
_zyGfifo_SGFfull,_zyGfifo_SLBreq,_zyGfifo_SLBrd,_zyGfifo_SLBwr,_zyGfifo_SLBfull,_zyGfifo_SRtkin);
// F1, L381
ixc_gfifo_port #(1,0,0,4,1) _zzGfifoF16_L381_p_0 (_zyGfifo_dflt_co[10],_zyGfifo_dflt_ci[10],_zyGfifoF16_L381_req_0,_zyGfifo__gfdL381_20_P0_m2_cbid,12'b0,1'b0,_zyGfifo_SGFtsReq,_zyGfifo_SGFcbid,_zyGfifo_SGFlen,_zyGfifo_SGFidata,
_zyGfifo_SGFfull,_zyGfifo_SLBreq,_zyGfifo_SLBrd,_zyGfifo_SLBwr,_zyGfifo_SLBfull,_zyGfifo_SRtkin);
// F1, L390
ixc_gfifo_port #(64,0,0,4,1) _zzGfifoF17_L390_p_0 (_zyGfifo_dflt_co[11],_zyGfifo_dflt_ci[11],_zyGfifoF17_L390_req_0,_zyGfifo__gfdL390_19_P0_m2_cbid,12'b010,_zyGfifoF17_L390_data_0,_zyGfifo_SGFtsReq,_zyGfifo_SGFcbid,_zyGfifo_SGFlen,_zyGfifo_SGFidata,
_zyGfifo_SGFfull,_zyGfifo_SLBreq,_zyGfifo_SLBrd,_zyGfifo_SLBwr,_zyGfifo_SLBfull,_zyGfifo_SRtkin);
// F1, L530
ixc_gfifo_port #(32,0,0,4,1) _zzGfifoF18_L530_p_0 (_zyGfifo_dflt_co[12],_zyGfifo_dflt_ci[12],_zyGfifoF18_L530_req_0,_zyGfifo__gfdL530_18_P0_m2_cbid,12'b01,_zyGfifoF18_L530_data_0,_zyGfifo_SGFtsReq,_zyGfifo_SGFcbid,_zyGfifo_SGFlen,_zyGfifo_SGFidata,
_zyGfifo_SGFfull,_zyGfifo_SLBreq,_zyGfifo_SLBrd,_zyGfifo_SLBwr,_zyGfifo_SLBfull,_zyGfifo_SRtkin);
// F1, L412
ixc_gfifo_port #(8,0,0,4,1) _zzGfifoF19_L412_p_0 (_zyGfifo_dflt_co[13],_zyGfifo_dflt_ci[13],_zyGfifoF19_L412_req_0,_zyGfifo__gfdL412_17_P0_m2_cbid,12'b01,_zyGfifoF19_L412_data_0,_zyGfifo_SGFtsReq,_zyGfifo_SGFcbid,_zyGfifo_SGFlen,_zyGfifo_SGFidata,
_zyGfifo_SGFfull,_zyGfifo_SLBreq,_zyGfifo_SLBrd,_zyGfifo_SLBwr,_zyGfifo_SLBfull,_zyGfifo_SRtkin);
// F1, L209
ixc_gfifo_port #(32,0,0,4,1) _zzGfifoF20_L209_p_0 (_zyGfifo_dflt_co[14],_zyGfifo_dflt_ci[14],_zyGfifoF20_L209_req_0,_zyGfifo_ob_service_data_2_zyprefetch_m2_cbid,12'b01,_zyGfifoF20_L209_data_0,_zyGfifo_SGFtsReq,_zyGfifo_SGFcbid,_zyGfifo_SGFlen,_zyGfifo_SGFidata,
_zyGfifo_SGFfull,_zyGfifo_SLBreq,_zyGfifo_SLBrd,_zyGfifo_SLBwr,_zyGfifo_SLBfull,_zyGfifo_SRtkin);
// F1, L439
ixc_gfifo_port #(1,2,0,4,1) _zzGfifoF0_L439_s2_p_5 (_zyGfifo_dflt_co[15],_zyGfifo_dflt_ci[15],_zyGfifoF0_L439_s2_req_5,_zyGfifoF0_L439_s2_cbid_5,12'b0,1'b0,_zyGfifo_SGFtsReq,_zyGfifo_SGFcbid,_zyGfifo_SGFlen,_zyGfifo_SGFidata,
_zyGfifo_SGFfull,_zyGfifo_SLBreq,_zyGfifo_SLBrd,_zyGfifo_SLBwr,_zyGfifo_SLBfull,_zyGfifo_SRtkin);
// F1, L444
ixc_gfifo_port #(32,0,0,4,1) _zzGfifoF23_L444_p_0 (_zyGfifo_dflt_co[16],_zyGfifo_dflt_ci[16],_zyGfifoF23_L444_req_0,_zyGfifo__gfdL444_14_P0_m2_cbid,12'b01,_zyGfifoF23_L444_data_0,_zyGfifo_SGFtsReq,_zyGfifo_SGFcbid,_zyGfifo_SGFlen,_zyGfifo_SGFidata,
_zyGfifo_SGFfull,_zyGfifo_SLBreq,_zyGfifo_SLBrd,_zyGfifo_SLBwr,_zyGfifo_SLBfull,_zyGfifo_SRtkin);
// F1, L446
ixc_gfifo_port #(136,0,0,4,1) _zzGfifoF24_L446_p_0 (_zyGfifo_dflt_co[17],_zyGfifo_dflt_ci[17],_zyGfifoF24_L446_req_0,_zyGfifo__gfdL446_13_P0_m2_cbid,12'b0101,_zyGfifoF24_L446_data_0,_zyGfifo_SGFtsReq,_zyGfifo_SGFcbid,_zyGfifo_SGFlen,_zyGfifo_SGFidata,
_zyGfifo_SGFfull,_zyGfifo_SLBreq,_zyGfifo_SLBrd,_zyGfifo_SLBwr,_zyGfifo_SLBfull,_zyGfifo_SRtkin);
// F1, L460
ixc_gfifo_port #(64,0,1,4,1) _zzGfifoF25_L460_p_0 (_zyGfifo_dflt_co[18],_zyGfifo_dflt_ci[18],_zyGfifoF25_L460_req_0,_zyGfifo__gfdL460_12_P0_m2_cbid,12'b010,_zyGfifoF25_L460_data_0,_zyGfifo_SGFtsReq,_zyGfifo_SGFcbid,_zyGfifo_SGFlen,_zyGfifo_SGFidata,
_zyGfifo_SGFfull,_zyGfifo_SLBreq,_zyGfifo_SLBrd,_zyGfifo_SLBwr,_zyGfifo_SLBfull,_zyGfifo_SRtkin);
// F1, L530
ixc_gfifo_port #(32,0,0,4,1) _zzGfifoF26_L530_p_0 (_zyGfifo_dflt_co[19],_zyGfifo_dflt_ci[19],_zyGfifoF26_L530_req_0,_zyGfifo__gfdL530_11_P0_m2_cbid,12'b01,_zyGfifoF26_L530_data_0,_zyGfifo_SGFtsReq,_zyGfifo_SGFcbid,_zyGfifo_SGFlen,_zyGfifo_SGFidata,
_zyGfifo_SGFfull,_zyGfifo_SLBreq,_zyGfifo_SLBrd,_zyGfifo_SLBwr,_zyGfifo_SLBfull,_zyGfifo_SRtkin);
// F1, L480
ixc_gfifo_port #(8,0,0,4,1) _zzGfifoF27_L480_p_0 (_zyGfifo_dflt_co[20],_zyGfifo_dflt_ci[20],_zyGfifoF27_L480_req_0,_zyGfifo__gfdL480_10_P0_m2_cbid,12'b01,_zyGfifoF27_L480_data_0,_zyGfifo_SGFtsReq,_zyGfifo_SGFcbid,_zyGfifo_SGFlen,_zyGfifo_SGFidata,
_zyGfifo_SGFfull,_zyGfifo_SLBreq,_zyGfifo_SLBrd,_zyGfifo_SLBwr,_zyGfifo_SLBfull,_zyGfifo_SRtkin);
// F1, L482
ixc_gfifo_port #(128,0,1,4,1) _zzGfifoF28_L482_p_0 (_zyGfifo_dflt_co[21],_zyGfifo_dflt_ci[21],_zyGfifoF28_L482_req_0,_zyGfifo__gfdL482_9_P0_m2_cbid,12'b0100,_zyGfifoF28_L482_data_0,_zyGfifo_SGFtsReq,_zyGfifo_SGFcbid,_zyGfifo_SGFlen,_zyGfifo_SGFidata,
_zyGfifo_SGFfull,_zyGfifo_SLBreq,_zyGfifo_SLBrd,_zyGfifo_SLBwr,_zyGfifo_SLBfull,_zyGfifo_SRtkin);
// F1, L487
ixc_gfifo_port #(16,0,1,4,1) _zzGfifoF29_L487_p_0 (_zyGfifo_dflt_co[22],_zyGfifo_dflt_ci[22],_zyGfifoF29_L487_req_0,_zyGfifo__gfdL487_8_P0_m2_cbid,12'b01,_zyGfifoF29_L487_data_0,_zyGfifo_SGFtsReq,_zyGfifo_SGFcbid,_zyGfifo_SGFlen,_zyGfifo_SGFidata,
_zyGfifo_SGFfull,_zyGfifo_SLBreq,_zyGfifo_SLBrd,_zyGfifo_SLBwr,_zyGfifo_SLBfull,_zyGfifo_SRtkin);
// F1, L491
ixc_gfifo_port #(16,0,1,4,1) _zzGfifoF30_L491_p_0 (_zyGfifo_dflt_co[23],_zyGfifo_dflt_ci[23],_zyGfifoF30_L491_req_0,_zyGfifo__gfdL491_7_P0_m2_cbid,12'b01,_zyGfifoF30_L491_data_0,_zyGfifo_SGFtsReq,_zyGfifo_SGFcbid,_zyGfifo_SGFlen,_zyGfifo_SGFidata,
_zyGfifo_SGFfull,_zyGfifo_SLBreq,_zyGfifo_SLBrd,_zyGfifo_SLBwr,_zyGfifo_SLBfull,_zyGfifo_SRtkin);
// F1, L496
ixc_gfifo_port #(16,0,1,4,1) _zzGfifoF31_L496_p_0 (_zyGfifo_dflt_co[24],_zyGfifo_dflt_ci[24],_zyGfifoF31_L496_req_0,_zyGfifo__gfdL496_6_P0_m2_cbid,12'b01,_zyGfifoF31_L496_data_0,_zyGfifo_SGFtsReq,_zyGfifo_SGFcbid,_zyGfifo_SGFlen,_zyGfifo_SGFidata,
_zyGfifo_SGFfull,_zyGfifo_SLBreq,_zyGfifo_SLBrd,_zyGfifo_SLBwr,_zyGfifo_SLBfull,_zyGfifo_SRtkin);
// F1, L253
ixc_gfifo_port #(560,3,1,4,1) _zzGfifoF0_L253_s4_p_6 (_zyGfifo_dflt_co[25],_zyGfifo_dflt_ci[25],_zyGfifoF0_L253_s4_req_6,_zyGfifoF0_L253_s4_cbid_6,_zyGfifoF0_L253_s4_len_6,_zyGfifoF0_L253_s4_data_6,_zyGfifo_SGFtsReq,_zyGfifo_SGFcbid,_zyGfifo_SGFlen,_zyGfifo_SGFidata,
_zyGfifo_SGFfull,_zyGfifo_SLBreq,_zyGfifo_SLBrd,_zyGfifo_SLBwr,_zyGfifo_SLBfull,_zyGfifo_SRtkin);
// F1, L253
ixc_gfifo_port #(1,2,0,4,1) _zzGfifoF1_L253_s2_p_7 (_zyGfifo_dflt_co[26],_zyGfifo_dflt_ci[26],_zyGfifoF1_L253_s2_req_7,_zyGfifoF1_L253_s2_cbid_7,12'b0,1'b0,_zyGfifo_SGFtsReq,_zyGfifo_SGFcbid,_zyGfifo_SGFlen,_zyGfifo_SGFidata,
_zyGfifo_SGFfull,_zyGfifo_SLBreq,_zyGfifo_SLBrd,_zyGfifo_SLBwr,_zyGfifo_SLBfull,_zyGfifo_SRtkin);
// F1, L10
assign  _zyGfifo_dflt_ci[0] = _zyGfifo_mod2_dflt_ci;
// F1, L10
assign  _zyGfifo_dflt_ci[1] = (_zyGfifo_dflt_co[0] | _zyGfifo_mod2_dflt_ci);
// F1, L10
assign  _zyGfifo_dflt_ci[2] = (( | _zyGfifo_dflt_co[1:0] ) | _zyGfifo_mod2_dflt_ci);
// F1, L10
assign  _zyGfifo_dflt_ci[3] = (( | _zyGfifo_dflt_co[2:0] ) | _zyGfifo_mod2_dflt_ci);
// F1, L10
assign  _zyGfifo_dflt_ci[4] = (( | _zyGfifo_dflt_co[3:0] ) | _zyGfifo_mod2_dflt_ci);
// F1, L10
assign  _zyGfifo_dflt_ci[5] = (( | _zyGfifo_dflt_co[4:0] ) | _zyGfifo_mod2_dflt_ci);
// F1, L10
assign  _zyGfifo_dflt_ci[6] = (( | _zyGfifo_dflt_co[5:0] ) | _zyGfifo_mod2_dflt_ci);
// F1, L10
assign  _zyGfifo_dflt_ci[7] = (( | _zyGfifo_dflt_co[6:0] ) | _zyGfifo_mod2_dflt_ci);
// F1, L10
assign  _zyGfifo_dflt_ci[8] = (( | _zyGfifo_dflt_co[7:0] ) | _zyGfifo_mod2_dflt_ci);
// F1, L10
assign  _zyGfifo_dflt_ci[9] = (( | _zyGfifo_dflt_co[8:0] ) | _zyGfifo_mod2_dflt_ci);
// F1, L10
assign  _zyGfifo_dflt_ci[10] = (( | _zyGfifo_dflt_co[9:0] ) | _zyGfifo_mod2_dflt_ci);
// F1, L10
assign  _zyGfifo_dflt_ci[11] = (( | _zyGfifo_dflt_co[10:0] ) | _zyGfifo_mod2_dflt_ci);
// F1, L10
assign  _zyGfifo_dflt_ci[12] = (( | _zyGfifo_dflt_co[11:0] ) | _zyGfifo_mod2_dflt_ci);
// F1, L10
assign  _zyGfifo_dflt_ci[13] = (( | _zyGfifo_dflt_co[12:0] ) | _zyGfifo_mod2_dflt_ci);
// F1, L10
assign  _zyGfifo_dflt_ci[14] = (( | _zyGfifo_dflt_co[13:0] ) | _zyGfifo_mod2_dflt_ci);
// F1, L10
assign  _zyGfifo_dflt_ci[15] = (( | _zyGfifo_dflt_co[14:0] ) | _zyGfifo_mod2_dflt_ci);
// F1, L10
assign  _zyGfifo_dflt_ci[16] = (( | _zyGfifo_dflt_co[15:0] ) | _zyGfifo_mod2_dflt_ci);
// F1, L10
assign  _zyGfifo_dflt_ci[17] = (( | _zyGfifo_dflt_co[16:0] ) | _zyGfifo_mod2_dflt_ci);
// F1, L10
assign  _zyGfifo_dflt_ci[18] = (( | _zyGfifo_dflt_co[17:0] ) | _zyGfifo_mod2_dflt_ci);
// F1, L10
assign  _zyGfifo_dflt_ci[19] = (( | _zyGfifo_dflt_co[18:0] ) | _zyGfifo_mod2_dflt_ci);
// F1, L10
assign  _zyGfifo_dflt_ci[20] = (( | _zyGfifo_dflt_co[19:0] ) | _zyGfifo_mod2_dflt_ci);
// F1, L10
assign  _zyGfifo_dflt_ci[21] = (( | _zyGfifo_dflt_co[20:0] ) | _zyGfifo_mod2_dflt_ci);
// F1, L10
assign  _zyGfifo_dflt_ci[22] = (( | _zyGfifo_dflt_co[21:0] ) | _zyGfifo_mod2_dflt_ci);
// F1, L10
assign  _zyGfifo_dflt_ci[23] = (( | _zyGfifo_dflt_co[22:0] ) | _zyGfifo_mod2_dflt_ci);
// F1, L10
assign  _zyGfifo_dflt_ci[24] = (( | _zyGfifo_dflt_co[23:0] ) | _zyGfifo_mod2_dflt_ci);
// F1, L10
assign  _zyGfifo_dflt_ci[25] = (( | _zyGfifo_dflt_co[24:0] ) | _zyGfifo_mod2_dflt_ci);
// F1, L10
assign  _zyGfifo_dflt_ci[26] = (( | _zyGfifo_dflt_co[25:0] ) | _zyGfifo_mod2_dflt_ci);
// F1, L10
assign  _zyGfifo_mod2_dflt_co = ( | _zyGfifo_dflt_co );
// F1, L324
ixc_mevClk #(3,0,0,3'b100,3'b0,3'b011,3'b0,3'b0,3'b0) _zzM2L324_pbcMevClk4 (_zyM2L324_pbcMevClk4,{clk,_zyL94_iscX1c0_f,_zyL61_iscX2c0_f},{(_zyM2L324_pbcCapEn0 | _zyM2L355_pbcCapEn3),_zyM2L333_pbcCapEn1,_zyM2L349_pbcCapEn2},1'b0,1'b0,_zyM2L324_pbcReq4,_zyM2L324_pbcBusy4,_zyM2L324_pbcWait4);
// F1, L253
ixc_mevClk #(2,0,0,2'b01,2'b0,2'b0,2'b0,2'b0,2'b0) _zzM2L253_pbcMevClk12 (_zyM2L253_pbcMevClk12,{_zyixc_port_0_0_req,clk},{_zyM2L253_pbcCapEn5,(((((_zyM2L274_pbcCapEn6 | _zyM2L287_pbcCapEn7) | _zyM2L293_pbcCapEn8) | _zyM2L295_pbcCapEn9) | _zyM2L364_pbcCapEn10) | _zyM2L300_pbcCapEn11)},1'b0,1'b0,_zyM2L253_pbcReq12,_zyM2L253_pbcBusy12,_zyM2L253_pbcWait12);
apb_xactor apb_xactor(
  .psel(_zy_simnet_kme_apb_psel_0_w$) ,
  .penable(_zy_simnet_kme_apb_penable_1_w$) ,
  .paddr(_zy_simnet_kme_apb_paddr_2_w$) ,
  .pwdata(_zy_simnet_kme_apb_pwdata_3_w$) ,
  .pwrite(_zy_simnet_kme_apb_pwrite_4_w$) ,
  .clk(_zy_simnet_clk_5_w$) ,
  .reset_n(_zy_simnet_rst_n_6_w$) ,
  .prdata(_zy_simnet_kme_apb_prdata_7_w$) ,
  .pready(_zy_simnet_kme_apb_pready_8_w$) ,
  .pslverr(_zy_simnet_kme_apb_pslverr_9_w$) ); 
cr_kme kme_dut(
  .kme_interrupt(_zy_simnet_dio_10) ,
  .kme_ib_tready(_zy_simnet_kme_ib_tready_11_w$) ,
  .kme_cceip0_ob_tvalid(_zy_simnet_kme_ob_tvalid_12_w$) ,
  .kme_cceip0_ob_tlast(_zy_simnet_kme_ob_tlast_13_w$) ,
  .kme_cceip0_ob_tid(_zy_simnet_kme_ob_tid_14_w$) ,
  .kme_cceip0_ob_tstrb(_zy_simnet_kme_ob_tstrb_15_w$) ,
  .kme_cceip0_ob_tuser(_zy_simnet_kme_ob_tuser_16_w$) ,
  .kme_cceip0_ob_tdata(_zy_simnet_kme_ob_tdata_17_w$) ,
  .apb_prdata(_zy_simnet_kme_apb_prdata_18_w$) ,
  .apb_pready(_zy_simnet_kme_apb_pready_19_w$) ,
  .apb_pslverr(_zy_simnet_kme_apb_pslverr_20_w$) ,
  .kme_idle(_zy_simnet_dio_21) ,
  .clk(_zy_simnet_clk_22_w$) ,
  .rst_n(_zy_simnet_rst_n_23_w$) ,
  .scan_en(_zy_simnet_cio_24) ,
  .scan_mode(_zy_simnet_cio_25) ,
  .scan_rst_n(_zy_simnet_cio_26) ,
  .ovstb(_zy_simnet_cio_27) ,
  .lvm(_zy_simnet_cio_28) ,
  .mlvm(_zy_simnet_cio_29) ,
  .disable_debug_cmd(_zy_simnet_cio_30) ,
  .disable_unencrypted_keys(_zy_simnet_cio_31) ,
  .kme_ib_tvalid(_zy_simnet_kme_ib_tvalid_32_w$) ,
  .kme_ib_tlast(_zy_simnet_kme_ib_tlast_33_w$) ,
  .kme_ib_tid(_zy_simnet_kme_ib_tid_34_w$) ,
  .kme_ib_tstrb(_zy_simnet_kme_ib_tstrb_35_w$) ,
  .kme_ib_tuser(_zy_simnet_kme_ib_tuser_36_w$) ,
  .kme_ib_tdata(_zy_simnet_kme_ib_tdata_37_w$) ,
  .kme_cceip0_ob_tready(_zy_simnet_kme_ob_tready_38_w$) ,
  .apb_paddr(_zy_simnet_kme_apb_paddr_39_w$) ,
  .apb_psel(_zy_simnet_kme_apb_psel_40_w$) ,
  .apb_penable(_zy_simnet_kme_apb_penable_41_w$) ,
  .apb_pwrite(_zy_simnet_kme_apb_pwrite_42_w$) ,
  .apb_pwdata(_zy_simnet_kme_apb_pwdata_43_w$) ); 
import "DPI-C" function int get_config_data (output bit [7:0] operation ,output bit [31:0] address ,output bit [31:0] data );
import "DPI-C" function int ib_service_data (output bit [63:0] tdata ,output bit [31:0] tuser_string ,output bit [7:0] tstrb ,output bit [31:0] str_get );
import "DPI-C" function int ob_service_data (output bit [63:0] tdata ,output bit [31:0] tuser_string ,output bit [7:0] tstrb ,output bit [31:0] str_get );

task tb_task;
 int _gpid;
 int _lpid;
// synopsys translate_off
 _zyifsyn_tb_task_2_ipt(_gpid);
 IXC_GFIFO.OSF.OSF_wait(_gpid,_lpid);
 _zyifsyn_tb_task_2_ipt_p2(_gpid);
// synopsys translate_on
endtask


task do_kme_config;
 config_ready = 1'b1;
 @(posedge clk)
  begin
  end
 $display("APB_INFO:  @time:%-d Exiting APB engine config ...",$time);
endtask


task service_ib_interface;
 static int stop_loop = 1000;
 saw_mega = 1'b0;
 saw_guid_tlv = 1'b0;
 mega_tlv_word_count = 0;
 have_guid_tlv = 1'b0;
 ready_ib = 1'b1;
 kme_ib_tvalid <= 1'b0;
 kme_ib_tlast <= 1'b0;
 @(posedge clk)
  begin
  end
 $display("INBOUND_INFO:  @time:%-d Exiting INBOUND thread...",$time);
endtask


task service_ob_interface;
 saw_cqe = 1'b0;
 saw_stats = 1'b0;
 watchdog_timer = 0;
 ready_ob = 1'b1;
 @(posedge clk)
  begin
  end
 $display("OUTBOUND_INFO:  @time:%-d Exiting OUTBOUND thread...",$time);
endtask


function  [24:0] reverse_translate_tuser;
 input bit [31:0] tuser ;
 if ((tuser == 32'b01011))
  // F1, L518
  begin
   // F1, L519
   $display("am i translating\n");
   return 25'b010100110110111101010100;
  end
 else
  if ((tuser == 32'b01010))
   // F1, L521
   begin
    // F1, L522
    $display("am i translating\n");
    return 25'b010001010110111101010100;
   end
  else
   // F1, L524
   begin
    // F1, L525
    return 25'b0;
   end
endfunction


function  [7:0] translate_tuser_t;
 input bit [24:0] tuser ;
 $display("inside translate function the tuser is : %s\n",tuser);
 if ((tuser == 25'b010100110110111101010100))
  // F1, L531
  begin
   // F1, L532
   return 8'b01;
  end
 else
  if ((tuser == 25'b010001010110111101010100))
   // F1, L533
   begin
    // F1, L534
    return 8'b010;
   end
  else
   // F1, L535
   begin
    // F1, L536
    return 8'b011;
   end
endfunction


function void get_config_data_zyackf_2_call;
 input int eos;
 _zygsfis_get_config_data_ack = (_zygsfis_get_config_data_ack + 32'b01);
 _zygsfis_get_config_data_eos = eos;
endfunction


function void get_config_data_zyputf_2_call;
 input bit [7:0] operation ;
 input bit [31:0] address ;
 input bit [31:0] data ;
 _zygsfis_get_config_data_fifo[_zygsfis_get_config_data_wptr] = {operation,address,data};
 _zygsfis_get_config_data_wptr = (_zygsfis_get_config_data_wptr + 32'b01);
endfunction

import "DPI-C"  context function void get_config_data_2_zyprefetch (input int size);

function int get_config_data_isf;
 output bit [7:0] operation ;
 output bit [31:0] address ;
 output bit [31:0] data ;
 int xr;
 xr = 0;
 if ((_zygsfis_get_config_data_rptr != _zygsfis_get_config_data_wptr))
  // F1, L206
  begin
   // F1, L206
   xr[0] = 1'b1;
   {operation,address,data} = _zygsfis_get_config_data_fifo[_zygsfis_get_config_data_rptr];
   _zygsfis_get_config_data_rptr = (_zygsfis_get_config_data_rptr + 32'b01);
   _zygsfis_get_config_data_space = (_zygsfis_get_config_data_space + 32'b01);
  end
 xr[1] = ((_zygsfis_get_config_data_rptr == _zygsfis_get_config_data_wptr) & _zygsfis_get_config_data_eos);
 if (( ~xr[1] ))
  // F1, L206
  begin
   // F1, L206
   if ((_zygsfis_get_config_data_req == _zygsfis_get_config_data_ack))
    _zygsfis_get_config_data_space = ( ~(_zygsfis_get_config_data_wptr - _zygsfis_get_config_data_rptr) );
   if ((_zygsfis_get_config_data_space >= 32'b01000))
    // F0, L0
    begin
     // F0, L0
     _zygsfis_get_config_data_req = (_zygsfis_get_config_data_req + 32'b01);
// synopsys translate_off
     get_config_data_2_zyprefetch(_zygsfis_get_config_data_space);
// synopsys translate_on
     _zygsfis_get_config_data_space = 5'b0;
    end
  end
 return xr;
endfunction


function void ib_service_data_zyackf_2_call;
 input int eos;
 _zygsfis_ib_service_data_ack = (_zygsfis_ib_service_data_ack + 32'b01);
 _zygsfis_ib_service_data_eos = eos;
endfunction


function void ib_service_data_zyputf_2_call;
 input bit [63:0] tdata ;
 input bit [31:0] tuser_string ;
 input bit [7:0] tstrb ;
 input bit [31:0] str_get ;
 _zygsfis_ib_service_data_fifo[_zygsfis_ib_service_data_wptr] = {tdata,tuser_string,tstrb,str_get};
 _zygsfis_ib_service_data_wptr = (_zygsfis_ib_service_data_wptr + 32'b01);
endfunction

import "DPI-C"  context function void ib_service_data_2_zyprefetch (input int size);

function int ib_service_data_isf;
 output bit [63:0] tdata ;
 output bit [31:0] tuser_string ;
 output bit [7:0] tstrb ;
 output bit [31:0] str_get ;
 int xr;
 xr = 0;
 if ((_zygsfis_ib_service_data_rptr != _zygsfis_ib_service_data_wptr))
  // F1, L207
  begin
   // F1, L207
   xr[0] = 1'b1;
   {tdata,tuser_string,tstrb,str_get} = _zygsfis_ib_service_data_fifo[_zygsfis_ib_service_data_rptr];
   _zygsfis_ib_service_data_rptr = (_zygsfis_ib_service_data_rptr + 32'b01);
   _zygsfis_ib_service_data_space = (_zygsfis_ib_service_data_space + 32'b01);
  end
 xr[1] = ((_zygsfis_ib_service_data_rptr == _zygsfis_ib_service_data_wptr) & _zygsfis_ib_service_data_eos);
 if (( ~xr[1] ))
  // F1, L207
  begin
   // F1, L207
   if ((_zygsfis_ib_service_data_req == _zygsfis_ib_service_data_ack))
    _zygsfis_ib_service_data_space = ( ~(_zygsfis_ib_service_data_wptr - _zygsfis_ib_service_data_rptr) );
   if ((_zygsfis_ib_service_data_space >= 32'b01000))
    // F0, L0
    begin
     // F0, L0
     _zygsfis_ib_service_data_req = (_zygsfis_ib_service_data_req + 32'b01);
// synopsys translate_off
     ib_service_data_2_zyprefetch(_zygsfis_ib_service_data_space);
// synopsys translate_on
     _zygsfis_ib_service_data_space = 5'b0;
    end
  end
 return xr;
endfunction


function void ob_service_data_zyackf_2_call;
 input int eos;
 _zygsfis_ob_service_data_ack = (_zygsfis_ob_service_data_ack + 32'b01);
 _zygsfis_ob_service_data_eos = eos;
endfunction


function void ob_service_data_zyputf_2_call;
 input bit [63:0] tdata ;
 input bit [31:0] tuser_string ;
 input bit [7:0] tstrb ;
 input bit [31:0] str_get ;
 _zygsfis_ob_service_data_fifo[_zygsfis_ob_service_data_wptr] = {tdata,tuser_string,tstrb,str_get};
 _zygsfis_ob_service_data_wptr = (_zygsfis_ob_service_data_wptr + 32'b01);
endfunction

import "DPI-C"  context function void ob_service_data_2_zyprefetch (input int size);

function int ob_service_data_isf;
 output bit [63:0] tdata ;
 output bit [31:0] tuser_string ;
 output bit [7:0] tstrb ;
 output bit [31:0] str_get ;
 int xr;
 xr = 0;
 if ((_zygsfis_ob_service_data_rptr != _zygsfis_ob_service_data_wptr))
  // F1, L209
  begin
   // F1, L209
   xr[0] = 1'b1;
   {tdata,tuser_string,tstrb,str_get} = _zygsfis_ob_service_data_fifo[_zygsfis_ob_service_data_rptr];
   _zygsfis_ob_service_data_rptr = (_zygsfis_ob_service_data_rptr + 32'b01);
   _zygsfis_ob_service_data_space = (_zygsfis_ob_service_data_space + 32'b01);
  end
 xr[1] = ((_zygsfis_ob_service_data_rptr == _zygsfis_ob_service_data_wptr) & _zygsfis_ob_service_data_eos);
 if (( ~xr[1] ))
  // F1, L209
  begin
   // F1, L209
   if ((_zygsfis_ob_service_data_req == _zygsfis_ob_service_data_ack))
    _zygsfis_ob_service_data_space = ( ~(_zygsfis_ob_service_data_wptr - _zygsfis_ob_service_data_rptr) );
   if ((_zygsfis_ob_service_data_space >= 32'b01000))
    // F0, L0
    begin
     // F0, L0
     _zygsfis_ob_service_data_req = (_zygsfis_ob_service_data_req + 32'b01);
// synopsys translate_off
     ob_service_data_2_zyprefetch(_zygsfis_ob_service_data_space);
// synopsys translate_on
     _zygsfis_ob_service_data_space = 5'b0;
    end
  end
 return xr;
endfunction


task _zyifsyn_tb_task_2_xpt;
 error_cntr = 0;
 rst_n = 1'b0;
 if ($test$plusargs("SEED"))
  // F1, L257
  begin
   // F1, L258
   _zz_58_258_2 = $value$plusargs("SEED=%d",seed);
  end
 else
  // F1, L259
  begin
   // F1, L260
   seed = 280'b0110001;
  end
 if ($test$plusargs("TESTNAME"))
  // F1, L263
  begin
   // F1, L264
   _zz_58_264_3 = $value$plusargs("TESTNAME=%s",testname);
   $display("TESTNAME=%s SEED=%s",testname,seed);
  end
 else
  // F1, L266
  begin
   // F1, L267
   testname = 280'b01110101011011100110101101101110011011110111011101101110;
   $display("TESTNAME=%s SEED=%s",testname,seed);
  end
 $display("--- \"rst_n\" is being asserted for 100ns ---");
 repeat (125)
  // F1, L273
  begin
   // F1, L274
   @(posedge clk)
    begin
    end
  end
 $display("STOP \n");
 kme_ib_tid <= 1'b0;
 kme_ib_tvalid <= 1'b0;
 kme_ib_tlast <= 1'b0;
 kme_ib_tdata <= 64'b0;
 kme_ib_tstrb <= 8'b0;
 kme_ib_tuser <= 8'b0;
 kme_ob_tready <= 1'b1;
 repeat (6.2500000000000000e+01)
  // F1, L286
  begin
   // F1, L287
   @(posedge clk)
    begin
    end
  end
 $display("--- \"rst_n\" has been DE-ASSERTED! ---");
 rst_n = 1'b1;
 repeat (125)
  // F1, L292
  begin
   // F1, L293
   @(posedge clk)
    begin
    end
  end
 @(posedge clk)
  begin
  end
 do_kme_config;
 config_done = 1'b1;
 repeat (1.2500000000000000e+01)
  // F1, L299
  begin
   // F1, L300
   @(posedge clk)
    begin
    end
  end
endtask

import "DPI-C"  context task _zyifsyn_tb_task_2_ipt (output int gpid);
import "DPI-C"  context task _zyifsyn_tb_task_2_ipt_p2 (input int gpid);

function void get_config_data_zyackf_m2p0_sim;
 input bit [31:0] iarg ;
 output bit oarg;
 // F1, L206
 begin
  // F1, L206
  get_config_data_zyackf_2_call(iarg[31:0]);
 end
endfunction

import "DPI-C"  context function void get_config_data_zyackf (input int eos);

function void get_config_data_zyputf_m2p0_sim;
 input bit [71:0] iarg ;
 output bit oarg;
 // F1, L206
 begin
  // F1, L206
  get_config_data_zyputf_2_call(iarg[7:0],iarg[39:8],iarg[71:40]);
 end
endfunction

import "DPI-C"  context function void get_config_data_zyputf (input bit [7:0] operation ,input bit [31:0] address ,input bit [31:0] data );

function void ib_service_data_zyackf_m2p0_sim;
 input bit [31:0] iarg ;
 output bit oarg;
 // F1, L207
 begin
  // F1, L207
  ib_service_data_zyackf_2_call(iarg[31:0]);
 end
endfunction

import "DPI-C"  context function void ib_service_data_zyackf (input int eos);

function void ib_service_data_zyputf_m2p0_sim;
 input bit [135:0] iarg ;
 output bit oarg;
 // F1, L207
 begin
  // F1, L207
  ib_service_data_zyputf_2_call(iarg[63:0],iarg[95:64],iarg[103:96],iarg[135:104]);
 end
endfunction

import "DPI-C"  context function void ib_service_data_zyputf (input bit [63:0] tdata ,input bit [31:0] tuser_string ,input bit [7:0] tstrb ,input bit [31:0] str_get );

function void ob_service_data_zyackf_m2p0_sim;
 input bit [31:0] iarg ;
 output bit oarg;
 // F1, L209
 begin
  // F1, L209
  ob_service_data_zyackf_2_call(iarg[31:0]);
 end
endfunction

import "DPI-C"  context function void ob_service_data_zyackf (input int eos);

function void ob_service_data_zyputf_m2p0_sim;
 input bit [135:0] iarg ;
 output bit oarg;
 // F1, L209
 begin
  // F1, L209
  ob_service_data_zyputf_2_call(iarg[63:0],iarg[95:64],iarg[103:96],iarg[135:104]);
 end
endfunction

import "DPI-C"  context function void ob_service_data_zyputf (input bit [63:0] tdata ,input bit [31:0] tuser_string ,input bit [7:0] tstrb ,input bit [31:0] str_get );

task _zzictd_finishT_L10_0;
 $finish;
endtask

import "DPI-C"  context function void xc_gfifo_sim (input int cbid,input int len,input bit [] data );
// F1, L10
initial 
 // F1, L10
 begin
  // F1, L306
  _zyL306_meState0 = 1'b0;
  _zyL312_meState2 = 1'b0;
  _zyL368_meState4 = 1'b0;
  _zyL439_meState8 = 2'b0;
 end

import "DPI-C" context function int xc_gfifo_new(string name, string cbidVar, string offVar, int needsTime, int forceLocal, int forceToSvChannel, int svContext, int argLen, int varArgs);

const bit [19:0] _zyGfifo__gfdL435_34_P0_m2_cbid_cv = xc_gfifo_new("_gfdL435_34_P0_gfifo_m2p0", "_zyGfifo__gfdL435_34_P0_m2_cbid", "_zyGfifo__gfdL435_34_P0_m2_gfOff", 1, 0, 0, 0, 0, 0);
initial _zyGfifo__gfdL435_34_P0_m2_cbid = _zyGfifo__gfdL435_34_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL513_33_P0_m2_cbid_cv = xc_gfifo_new("_gfdL513_33_P0_gfifo_m2p0", "_zyGfifo__gfdL513_33_P0_m2_cbid", "_zyGfifo__gfdL513_33_P0_m2_gfOff", 1, 0, 0, 0, 0, 0);
initial _zyGfifo__gfdL513_33_P0_m2_cbid = _zyGfifo__gfdL513_33_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL316_32_P0_m2_cbid_cv = xc_gfifo_new("_gfdL316_32_P0_gfifo_m2p0", "_zyGfifo__gfdL316_32_P0_m2_cbid", "_zyGfifo__gfdL316_32_P0_m2_gfOff", 0, 0, 0, 0, 9, 0);
initial _zyGfifo__gfdL316_32_P0_m2_cbid = _zyGfifo__gfdL316_32_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL318_31_P0_m2_cbid_cv = xc_gfifo_new("_gfdL318_31_P0_gfifo_m2p0", "_zyGfifo__gfdL318_31_P0_m2_cbid", "_zyGfifo__gfdL318_31_P0_m2_gfOff", 0, 0, 0, 0, 9, 0);
initial _zyGfifo__gfdL318_31_P0_m2_cbid = _zyGfifo__gfdL318_31_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo_get_config_data_2_zyprefetch_m2_cbid_cv = xc_gfifo_new("get_config_data_2_zyprefetch_gfifo_m2p0", "_zyGfifo_get_config_data_2_zyprefetch_m2_cbid", "_zyGfifo_get_config_data_2_zyprefetch_m2_gfOff", 0, 0, 0, 0, 1, 0);
initial _zyGfifo_get_config_data_2_zyprefetch_m2_cbid = _zyGfifo_get_config_data_2_zyprefetch_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL327_30_P0_m2_cbid_cv = xc_gfifo_new("_gfdL327_30_P0_gfifo_m2p0", "_zyGfifo__gfdL327_30_P0_m2_cbid", "_zyGfifo__gfdL327_30_P0_m2_gfOff", 0, 0, 0, 0, 1, 0);
initial _zyGfifo__gfdL327_30_P0_m2_cbid = _zyGfifo__gfdL327_30_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL330_29_P0_m2_cbid_cv = xc_gfifo_new("_gfdL330_29_P0_gfifo_m2p0", "_zyGfifo__gfdL330_29_P0_m2_cbid", "_zyGfifo__gfdL330_29_P0_m2_gfOff", 0, 0, 0, 0, 3, 0);
initial _zyGfifo__gfdL330_29_P0_m2_cbid = _zyGfifo__gfdL330_29_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL334_28_P0_m2_cbid_cv = xc_gfifo_new("_gfdL334_28_P0_gfifo_m2p0", "_zyGfifo__gfdL334_28_P0_m2_cbid", "_zyGfifo__gfdL334_28_P0_m2_gfOff", 0, 0, 0, 0, 3, 0);
initial _zyGfifo__gfdL334_28_P0_m2_cbid = _zyGfifo__gfdL334_28_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL336_27_P0_m2_cbid_cv = xc_gfifo_new("_gfdL336_27_P0_gfifo_m2p0", "_zyGfifo__gfdL336_27_P0_m2_cbid", "_zyGfifo__gfdL336_27_P0_m2_gfOff", 1, 0, 0, 0, 1, 0);
initial _zyGfifo__gfdL336_27_P0_m2_cbid = _zyGfifo__gfdL336_27_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL341_26_P0_m2_cbid_cv = xc_gfifo_new("_gfdL341_26_P0_gfifo_m2p0", "_zyGfifo__gfdL341_26_P0_m2_cbid", "_zyGfifo__gfdL341_26_P0_m2_gfOff", 1, 0, 0, 0, 2, 0);
initial _zyGfifo__gfdL341_26_P0_m2_cbid = _zyGfifo__gfdL341_26_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL351_25_P0_m2_cbid_cv = xc_gfifo_new("_gfdL351_25_P0_gfifo_m2p0", "_zyGfifo__gfdL351_25_P0_m2_cbid", "_zyGfifo__gfdL351_25_P0_m2_gfOff", 1, 0, 0, 0, 1, 0);
initial _zyGfifo__gfdL351_25_P0_m2_cbid = _zyGfifo__gfdL351_25_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo_ib_service_data_2_zyprefetch_m2_cbid_cv = xc_gfifo_new("ib_service_data_2_zyprefetch_gfifo_m2p0", "_zyGfifo_ib_service_data_2_zyprefetch_m2_cbid", "_zyGfifo_ib_service_data_2_zyprefetch_m2_gfOff", 0, 0, 0, 0, 1, 0);
initial _zyGfifo_ib_service_data_2_zyprefetch_m2_cbid = _zyGfifo_ib_service_data_2_zyprefetch_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL519_24_P0_m2_cbid_cv = xc_gfifo_new("_gfdL519_24_P0_gfifo_m2p0", "_zyGfifo__gfdL519_24_P0_m2_cbid", "_zyGfifo__gfdL519_24_P0_m2_gfOff", 0, 0, 0, 0, 0, 0);
initial _zyGfifo__gfdL519_24_P0_m2_cbid = _zyGfifo__gfdL519_24_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL522_23_P0_m2_cbid_cv = xc_gfifo_new("_gfdL522_23_P0_gfifo_m2p0", "_zyGfifo__gfdL522_23_P0_m2_cbid", "_zyGfifo__gfdL522_23_P0_m2_gfOff", 0, 0, 0, 0, 0, 0);
initial _zyGfifo__gfdL522_23_P0_m2_cbid = _zyGfifo__gfdL522_23_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL373_22_P0_m2_cbid_cv = xc_gfifo_new("_gfdL373_22_P0_gfifo_m2p0", "_zyGfifo__gfdL373_22_P0_m2_cbid", "_zyGfifo__gfdL373_22_P0_m2_gfOff", 0, 0, 0, 0, 1, 0);
initial _zyGfifo__gfdL373_22_P0_m2_cbid = _zyGfifo__gfdL373_22_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL375_21_P0_m2_cbid_cv = xc_gfifo_new("_gfdL375_21_P0_gfifo_m2p0", "_zyGfifo__gfdL375_21_P0_m2_cbid", "_zyGfifo__gfdL375_21_P0_m2_gfOff", 0, 0, 0, 0, 5, 0);
initial _zyGfifo__gfdL375_21_P0_m2_cbid = _zyGfifo__gfdL375_21_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL381_20_P0_m2_cbid_cv = xc_gfifo_new("_gfdL381_20_P0_gfifo_m2p0", "_zyGfifo__gfdL381_20_P0_m2_cbid", "_zyGfifo__gfdL381_20_P0_m2_gfOff", 0, 0, 0, 0, 0, 0);
initial _zyGfifo__gfdL381_20_P0_m2_cbid = _zyGfifo__gfdL381_20_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL390_19_P0_m2_cbid_cv = xc_gfifo_new("_gfdL390_19_P0_gfifo_m2p0", "_zyGfifo__gfdL390_19_P0_m2_cbid", "_zyGfifo__gfdL390_19_P0_m2_gfOff", 0, 0, 0, 0, 2, 0);
initial _zyGfifo__gfdL390_19_P0_m2_cbid = _zyGfifo__gfdL390_19_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL530_18_P0_m2_cbid_cv = xc_gfifo_new("_gfdL530_18_P0_gfifo_m2p0", "_zyGfifo__gfdL530_18_P0_m2_cbid", "_zyGfifo__gfdL530_18_P0_m2_gfOff", 0, 0, 0, 0, 1, 0);
initial _zyGfifo__gfdL530_18_P0_m2_cbid = _zyGfifo__gfdL530_18_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL412_17_P0_m2_cbid_cv = xc_gfifo_new("_gfdL412_17_P0_gfifo_m2p0", "_zyGfifo__gfdL412_17_P0_m2_cbid", "_zyGfifo__gfdL412_17_P0_m2_gfOff", 0, 0, 0, 0, 1, 0);
initial _zyGfifo__gfdL412_17_P0_m2_cbid = _zyGfifo__gfdL412_17_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo_ob_service_data_2_zyprefetch_m2_cbid_cv = xc_gfifo_new("ob_service_data_2_zyprefetch_gfifo_m2p0", "_zyGfifo_ob_service_data_2_zyprefetch_m2_cbid", "_zyGfifo_ob_service_data_2_zyprefetch_m2_gfOff", 0, 0, 0, 0, 1, 0);
initial _zyGfifo_ob_service_data_2_zyprefetch_m2_cbid = _zyGfifo_ob_service_data_2_zyprefetch_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL519_16_P0_m2_cbid_cv = xc_gfifo_new("_gfdL519_16_P0_gfifo_m2p0", "_zyGfifo__gfdL519_16_P0_m2_cbid", "_zyGfifo__gfdL519_16_P0_m2_gfOff", 0, 0, 0, 0, 0, 0);
initial _zyGfifo__gfdL519_16_P0_m2_cbid = _zyGfifo__gfdL519_16_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL522_15_P0_m2_cbid_cv = xc_gfifo_new("_gfdL522_15_P0_gfifo_m2p0", "_zyGfifo__gfdL522_15_P0_m2_cbid", "_zyGfifo__gfdL522_15_P0_m2_gfOff", 0, 0, 0, 0, 0, 0);
initial _zyGfifo__gfdL522_15_P0_m2_cbid = _zyGfifo__gfdL522_15_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL444_14_P0_m2_cbid_cv = xc_gfifo_new("_gfdL444_14_P0_gfifo_m2p0", "_zyGfifo__gfdL444_14_P0_m2_cbid", "_zyGfifo__gfdL444_14_P0_m2_gfOff", 0, 0, 0, 0, 1, 0);
initial _zyGfifo__gfdL444_14_P0_m2_cbid = _zyGfifo__gfdL444_14_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL446_13_P0_m2_cbid_cv = xc_gfifo_new("_gfdL446_13_P0_gfifo_m2p0", "_zyGfifo__gfdL446_13_P0_m2_cbid", "_zyGfifo__gfdL446_13_P0_m2_gfOff", 0, 0, 0, 0, 5, 0);
initial _zyGfifo__gfdL446_13_P0_m2_cbid = _zyGfifo__gfdL446_13_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL460_12_P0_m2_cbid_cv = xc_gfifo_new("_gfdL460_12_P0_gfifo_m2p0", "_zyGfifo__gfdL460_12_P0_m2_cbid", "_zyGfifo__gfdL460_12_P0_m2_gfOff", 1, 0, 0, 0, 2, 0);
initial _zyGfifo__gfdL460_12_P0_m2_cbid = _zyGfifo__gfdL460_12_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL530_11_P0_m2_cbid_cv = xc_gfifo_new("_gfdL530_11_P0_gfifo_m2p0", "_zyGfifo__gfdL530_11_P0_m2_cbid", "_zyGfifo__gfdL530_11_P0_m2_gfOff", 0, 0, 0, 0, 1, 0);
initial _zyGfifo__gfdL530_11_P0_m2_cbid = _zyGfifo__gfdL530_11_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL480_10_P0_m2_cbid_cv = xc_gfifo_new("_gfdL480_10_P0_gfifo_m2p0", "_zyGfifo__gfdL480_10_P0_m2_cbid", "_zyGfifo__gfdL480_10_P0_m2_gfOff", 0, 0, 0, 0, 1, 0);
initial _zyGfifo__gfdL480_10_P0_m2_cbid = _zyGfifo__gfdL480_10_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL482_9_P0_m2_cbid_cv = xc_gfifo_new("_gfdL482_9_P0_gfifo_m2p0", "_zyGfifo__gfdL482_9_P0_m2_cbid", "_zyGfifo__gfdL482_9_P0_m2_gfOff", 1, 0, 0, 0, 4, 0);
initial _zyGfifo__gfdL482_9_P0_m2_cbid = _zyGfifo__gfdL482_9_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL487_8_P0_m2_cbid_cv = xc_gfifo_new("_gfdL487_8_P0_gfifo_m2p0", "_zyGfifo__gfdL487_8_P0_m2_cbid", "_zyGfifo__gfdL487_8_P0_m2_gfOff", 1, 0, 0, 0, 1, 0);
initial _zyGfifo__gfdL487_8_P0_m2_cbid = _zyGfifo__gfdL487_8_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL491_7_P0_m2_cbid_cv = xc_gfifo_new("_gfdL491_7_P0_gfifo_m2p0", "_zyGfifo__gfdL491_7_P0_m2_cbid", "_zyGfifo__gfdL491_7_P0_m2_gfOff", 1, 0, 0, 0, 1, 0);
initial _zyGfifo__gfdL491_7_P0_m2_cbid = _zyGfifo__gfdL491_7_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL496_6_P0_m2_cbid_cv = xc_gfifo_new("_gfdL496_6_P0_gfifo_m2p0", "_zyGfifo__gfdL496_6_P0_m2_cbid", "_zyGfifo__gfdL496_6_P0_m2_gfOff", 1, 0, 0, 0, 1, 0);
initial _zyGfifo__gfdL496_6_P0_m2_cbid = _zyGfifo__gfdL496_6_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL265_5_P0_m2_cbid_cv = xc_gfifo_new("_gfdL265_5_P0_gfifo_m2p0", "_zyGfifo__gfdL265_5_P0_m2_cbid", "_zyGfifo__gfdL265_5_P0_m2_gfOff", 0, 0, 0, 0, 18, 0);
initial _zyGfifo__gfdL265_5_P0_m2_cbid = _zyGfifo__gfdL265_5_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL268_4_P0_m2_cbid_cv = xc_gfifo_new("_gfdL268_4_P0_gfifo_m2p0", "_zyGfifo__gfdL268_4_P0_m2_cbid", "_zyGfifo__gfdL268_4_P0_m2_gfOff", 0, 0, 0, 0, 18, 0);
initial _zyGfifo__gfdL268_4_P0_m2_cbid = _zyGfifo__gfdL268_4_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL271_3_P0_m2_cbid_cv = xc_gfifo_new("_gfdL271_3_P0_gfifo_m2p0", "_zyGfifo__gfdL271_3_P0_m2_cbid", "_zyGfifo__gfdL271_3_P0_m2_gfOff", 0, 0, 0, 0, 0, 0);
initial _zyGfifo__gfdL271_3_P0_m2_cbid = _zyGfifo__gfdL271_3_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL276_2_P0_m2_cbid_cv = xc_gfifo_new("_gfdL276_2_P0_gfifo_m2p0", "_zyGfifo__gfdL276_2_P0_m2_cbid", "_zyGfifo__gfdL276_2_P0_m2_gfOff", 0, 0, 0, 0, 0, 0);
initial _zyGfifo__gfdL276_2_P0_m2_cbid = _zyGfifo__gfdL276_2_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL289_1_P0_m2_cbid_cv = xc_gfifo_new("_gfdL289_1_P0_gfifo_m2p0", "_zyGfifo__gfdL289_1_P0_m2_cbid", "_zyGfifo__gfdL289_1_P0_m2_gfOff", 0, 0, 0, 0, 0, 0);
initial _zyGfifo__gfdL289_1_P0_m2_cbid = _zyGfifo__gfdL289_1_P0_m2_cbid_cv;

const bit [19:0] _zyGfifo__gfdL365_0_P0_m2_cbid_cv = xc_gfifo_new("_gfdL365_0_P0_gfifo_m2p0", "_zyGfifo__gfdL365_0_P0_m2_cbid", "_zyGfifo__gfdL365_0_P0_m2_gfOff", 1, 0, 0, 0, 0, 0);
initial _zyGfifo__gfdL365_0_P0_m2_cbid = _zyGfifo__gfdL365_0_P0_m2_cbid_cv;

// F1, L306
always 
 // F1, L306
 begin
  // F1, L433
  @(posedge clk)
   begin
   end
  // F1, L306
  begin:_zyL306_meSwitch0
   int _zystop_loop_L422_tfiV0_meV0;
   reg _zyL306_meEn1;
   // F1, L306
   _zyL306_meEn1 = 1'b1;
   case (_zyL306_meState0)
    1'b0:
     // F1, L306
     begin
      // F1, L306
      // F1, L306
      begin
       // F1, L307
       if ((config_done == 32'b01))
        // F1, L307
        begin
         // F1, L421
         // F1, L421
         begin:_zz_gfdinlCscp0_L308_service_ib_interface_meScp1
          // F1, L422
          _zystop_loop_L422_tfiV0_meV0 = 1000;
          saw_mega = 1'b0;
          saw_guid_tlv = 1'b0;
          mega_tlv_word_count = 0;
          have_guid_tlv = 1'b0;
          ready_ib = 1'b1;
          kme_ib_tvalid <= 1'b0;
          kme_ib_tlast <= 1'b0;
          _zyL306_meState0 = 1'b1;
          _zyL306_meEn1 = 1'b0;
         end
        end
      end
      if (_zyL306_meEn1)
       // F1, L306
       begin
        // F1, L306
        // F1, L306
        begin
         // F1, L306
         _zyL306_meState0 = 1'b0;
        end
       end
     end
    1'b1:
     // F1, L435
     begin
      // F1, L435
      _zyGfifoF0_L435_req_0 = (_zyGfifo__gfdL435_34_P0_m2_gfOff == _zyGfifoF0_L435_req_0);
// synopsys translate_off
      xc_gfifo_sim(_zyGfifo__gfdL435_34_P0_m2_cbid,32'b0,_zyGfifo_mod2_simData);
// synopsys translate_on
      // F1, L306
      begin
       // F1, L306
       _zyL306_meState0 = 1'b0;
      end
     end
   endcase
  end
 end
// F1, L312
always 
 // F1, L312
 begin
  // F1, L511
  @(posedge clk)
   begin
   end
  // F1, L312
  begin:_zyL312_meSwitch2
   reg _zyL312_meEn2;
   // F1, L312
   _zyL312_meEn2 = 1'b1;
   case (_zyL312_meState2)
    1'b0:
     // F1, L312
     begin
      // F1, L312
      // F1, L312
      begin
       // F1, L313
       if ((config_done == 32'b01))
        // F1, L313
        begin
         // F1, L505
         // F1, L505
         begin:_zz_gfdinlCscp1_L314_service_ob_interface_meScp3
          // F1, L506
          saw_cqe = 1'b0;
          saw_stats = 1'b0;
          watchdog_timer = 0;
          ready_ob = 1'b1;
          _zyL312_meState2 = 1'b1;
          _zyL312_meEn2 = 1'b0;
         end
        end
      end
      if (_zyL312_meEn2)
       // F1, L312
       begin
        // F1, L312
        // F1, L312
        begin
         // F1, L312
         _zyL312_meState2 = 1'b0;
        end
       end
     end
    1'b1:
     // F1, L513
     begin
      // F1, L513
      _zyGfifoF1_L513_req_0 = (_zyGfifo__gfdL513_33_P0_m2_gfOff == _zyGfifoF1_L513_req_0);
// synopsys translate_off
      xc_gfifo_sim(_zyGfifo__gfdL513_33_P0_m2_cbid,32'b0,_zyGfifo_mod2_simData);
// synopsys translate_on
      if (error_cntr)
       // F1, L315
       begin
        // F1, L316
        _zyGfifoF0_L312_s2_cbid_0 = _zyGfifo__gfdL316_32_P0_m2_cbid;
        _zyGfifoF0_L312_s2_data_0[279:0] = {280{1'b0}};
        _zyGfifoF0_L312_s2_data_0[279:0] = testname;
        _zyGfifoF0_L312_s2_req_0 = (_zyGfifo__gfdL316_32_P0_m2_gfOff == _zyGfifoF0_L312_s2_req_0);
// synopsys translate_off
        xc_gfifo_sim(_zyGfifo__gfdL316_32_P0_m2_cbid,32'b01001,_zyGfifoF0_L312_s2_data_0);
// synopsys translate_on
       end
      else
       // F1, L317
       begin
        // F1, L318
        _zyGfifoF0_L312_s2_cbid_0 = _zyGfifo__gfdL318_31_P0_m2_cbid;
        _zyGfifoF0_L312_s2_data_0[279:0] = {280{1'b0}};
        _zyGfifoF0_L312_s2_data_0[279:0] = testname;
        _zyGfifoF0_L312_s2_req_0 = (_zyGfifo__gfdL318_31_P0_m2_gfOff == _zyGfifoF0_L312_s2_req_0);
// synopsys translate_off
        xc_gfifo_sim(_zyGfifo__gfdL318_31_P0_m2_cbid,32'b01001,_zyGfifoF0_L312_s2_data_0);
// synopsys translate_on
       end
      _zyictd_finish_L320_0 = 1'b1;
      // F1, L312
      begin
       // F1, L312
       _zyL312_meState2 = 1'b0;
      end
     end
   endcase
  end
 end
// F1, L324
always 
 // F1, L324
 begin
  // F1, L324
  @(posedge _zyM2L324_pbcMevClk4)
   begin
   end
  // F1, L324
  begin:_zyM2L324_pbcFsm0
   // F1, L324
   case (_zyM2L324_pbcFsm0_s)
    3'b0:
     // F1, L324
     begin
      // F1, L324
      _zyM2L324_pbcEn13 = 1'b1;
      _zyM2L324_pbcCapEn0 = 1'b0;
      if ((config_ready == 32'b01))
       // F1, L325
       begin
        // F1, L206
        // F1, L206
        begin:_zygfifotfiCscp0_L326_get_config_data_isf_M2_pbcScp1
         // F0, L0
         _zyxr_L206_tfiV3_M2_pbcG3 = 0;
         if ((_zygsfis_get_config_data_rptr != _zygsfis_get_config_data_wptr))
          // F1, L206
          begin
          // F1, L206
          _zyxr_L206_tfiV3_M2_pbcG3[0] = 1'b1;
          {_zyoperation_L206_tfiV0_M2_pbcG0,_zyaddress_L206_tfiV1_M2_pbcG1,_zydata_L206_tfiV2_M2_pbcG2} = _zygsfis_get_config_data_fifo[_zygsfis_get_config_data_rptr];
          _zygsfis_get_config_data_rptr = (_zygsfis_get_config_data_rptr + 32'b01);
          _zygsfis_get_config_data_space = (_zygsfis_get_config_data_space + 32'b01);
          end
         _zyxr_L206_tfiV3_M2_pbcG3[1] = ((_zygsfis_get_config_data_rptr == _zygsfis_get_config_data_wptr) & _zygsfis_get_config_data_eos);
         if (( ~_zyxr_L206_tfiV3_M2_pbcG3[1] ))
          // F1, L206
          begin
          // F1, L206
          if ((_zygsfis_get_config_data_req == _zygsfis_get_config_data_ack))
          _zygsfis_get_config_data_space = ( ~(_zygsfis_get_config_data_wptr - _zygsfis_get_config_data_rptr) );
          if ((_zygsfis_get_config_data_space >= 32'b01000))
          // F0, L0
          begin
          // F0, L0
          _zygsfis_get_config_data_req = (_zygsfis_get_config_data_req + 32'b01);
          _zyGfifoF0_L324_s3_cbid_1 = _zyGfifo_get_config_data_2_zyprefetch_m2_cbid;
          _zyGfifoF0_L324_s3_len_1 = 12'b01;
          _zyGfifoF0_L324_s3_data_1[95:0] = 96'b0;
          _zyGfifoF0_L324_s3_data_1[31:0] = _zygsfis_get_config_data_space;
          _zyGfifoF0_L324_s3_req_1 = (_zyGfifo_get_config_data_2_zyprefetch_m2_gfOff == _zyGfifoF0_L324_s3_req_1);
// synopsys translate_off
          xc_gfifo_sim(_zyGfifo_get_config_data_2_zyprefetch_m2_cbid,32'b01,_zyGfifoF0_L324_s3_data_1);
// synopsys translate_on
          _zygsfis_get_config_data_space = 5'b0;
          end
          end
         _zyL326_tfiRv17 = _zyxr_L206_tfiV3_M2_pbcG3;
         operation = _zyoperation_L206_tfiV0_M2_pbcG0;
         address = _zyaddress_L206_tfiV1_M2_pbcG1;
         data = _zydata_L206_tfiV2_M2_pbcG2;
        end
        retval = _zyL326_tfiRv17;
        _zyGfifoF1_L324_s2_cbid_2 = _zyGfifo__gfdL327_30_P0_m2_cbid;
        _zyGfifoF1_L324_s2_data_2[31:0] = 32'b0;
        _zyGfifoF1_L324_s2_data_2[31:0] = retval;
        _zyGfifoF1_L324_s2_req_2 = (_zyGfifo__gfdL327_30_P0_m2_gfOff == _zyGfifoF1_L324_s2_req_2);
// synopsys translate_off
        xc_gfifo_sim(_zyGfifo__gfdL327_30_P0_m2_cbid,32'b01,_zyGfifoF1_L324_s2_data_2);
// synopsys translate_on
        if ((retval == 1))
         // F1, L328
         begin
          // F1, L330
          _zyGfifoF2_L324_s2_cbid_3 = _zyGfifo__gfdL330_29_P0_m2_cbid;
          _zyGfifoF2_L324_s2_len_3 = 12'b011;
          _zyGfifoF2_L324_s2_data_3[71:0] = 72'b0;
          _zyGfifoF2_L324_s2_data_3[71:64] = operation;
          _zyGfifoF2_L324_s2_data_3[63:32] = address;
          _zyGfifoF2_L324_s2_data_3[31:0] = data;
          _zyGfifoF2_L324_s2_req_3 = (_zyGfifo__gfdL330_29_P0_m2_gfOff == _zyGfifoF2_L324_s2_req_3);
// synopsys translate_off
          xc_gfifo_sim(_zyGfifo__gfdL330_29_P0_m2_cbid,32'b011,_zyGfifoF2_L324_s2_data_3);
// synopsys translate_on
          if (((((operation == 8'b01110010) || (operation == 8'b01010010)) || (operation == 8'b01110111)) || (operation == 8'b01010111)))
          // F1, L331
          begin
          // F1, L332
          if (((operation == 8'b01110010) || (operation == 8'b01010010)))
          // F1, L332
          begin
          // F1, L333
          _zyL94_iscX1c0_i0 = address;
          _zyL94_iscX1c0_s = _zyL94_iscX1c0_n;
          _zyL94_iscX1c0_n = ( ~_zyL94_iscX1c0_n );
          _zyM2L333_pbcCapEn1 = 1'b1;
          _zyM2L324_pbcFsm0_s = 3'b01;
          _zyM2L324_pbcEn13 = 1'b0;
          end
          else
          if (((operation == 8'b01110111) || (operation == 8'b01010111)))
          // F1, L348
          begin
          // F1, L349
          _zyL61_iscX2c0_i0 = address;
          _zyL61_iscX2c0_i1 = data;
          _zyL61_iscX2c0_s = _zyL61_iscX2c0_n;
          _zyL61_iscX2c0_n = ( ~_zyL61_iscX2c0_n );
          _zyM2L349_pbcCapEn2 = 1'b1;
          _zyM2L324_pbcFsm0_s = 3'b010;
          _zyM2L324_pbcEn13 = 1'b0;
          end
          if (_zyM2L324_pbcEn13)
          // F1, L355
          begin
          // F1, L355
          _zyM2L355_pbcCapEn3 = 1'b1;
          _zyM2L324_pbcFsm0_s = 3'b011;
          _zyM2L324_pbcEn13 = 1'b0;
          end
          end
         end
       end
      if (_zyM2L324_pbcEn13)
       // F1, L324
       begin
        // F1, L324
        _zyM2L324_pbcCapEn0 = 1'b1;
        _zyM2L324_pbcFsm0_s = 3'b0;
       end
     end
    3'b01:
     // F1, L333
     begin
      // F1, L333
      _zyM2L333_pbcCapEn1 = 1'b0;
      returned_data = _zyL94_iscX1c0_o1;
      response = _zyL94_iscX1c0_o2;
      _zyGfifoF0_L324_s3_cbid_1 = _zyGfifo__gfdL334_28_P0_m2_cbid;
      _zyGfifoF0_L324_s3_len_1 = 12'b011;
      _zyGfifoF0_L324_s3_data_1[95:0] = 96'b0;
      _zyGfifoF0_L324_s3_data_1[95:64] = address;
      _zyGfifoF0_L324_s3_data_1[63:32] = data;
      _zyGfifoF0_L324_s3_data_1[31:0] = returned_data;
      _zyGfifoF0_L324_s3_req_1 = (_zyGfifo__gfdL334_28_P0_m2_gfOff == _zyGfifoF0_L324_s3_req_1);
// synopsys translate_off
      xc_gfifo_sim(_zyGfifo__gfdL334_28_P0_m2_cbid,32'b011,_zyGfifoF0_L324_s3_data_1);
// synopsys translate_on
      if ((response !== 32'b0))
       // F1, L335
       begin
        // F1, L336
        _zyGfifoF1_L324_s2_cbid_2 = _zyGfifo__gfdL336_27_P0_m2_cbid;
        _zyGfifoF1_L324_s2_data_2[31:0] = 32'b0;
        _zyGfifoF1_L324_s2_data_2[31:0] = address;
        _zyGfifoF1_L324_s2_req_2 = (_zyGfifo__gfdL336_27_P0_m2_gfOff == _zyGfifoF1_L324_s2_req_2);
// synopsys translate_off
        xc_gfifo_sim(_zyGfifo__gfdL336_27_P0_m2_cbid,32'b01,_zyGfifoF1_L324_s2_data_2);
// synopsys translate_on
        _zyictd_finish_L338_1 = 1'b1;
       end
      if ((returned_data !== data))
       // F1, L340
       begin
        // F1, L341
        _zyGfifoF2_L324_s2_cbid_3 = _zyGfifo__gfdL341_26_P0_m2_cbid;
        _zyGfifoF2_L324_s2_len_3 = 12'b010;
        _zyGfifoF2_L324_s2_data_3[71:0] = 72'b0;
        _zyGfifoF2_L324_s2_data_3[63:32] = returned_data;
        _zyGfifoF2_L324_s2_data_3[31:0] = data;
        _zyGfifoF2_L324_s2_req_3 = (_zyGfifo__gfdL341_26_P0_m2_gfOff == _zyGfifoF2_L324_s2_req_3);
// synopsys translate_off
        xc_gfifo_sim(_zyGfifo__gfdL341_26_P0_m2_cbid,32'b010,_zyGfifoF2_L324_s2_data_3);
// synopsys translate_on
        error_cntr = (error_cntr + 1);
        if ((error_cntr > 10))
         // F1, L343
         begin
          // F1, L344
          _zyictd_finish_L338_1 = 1'b1;
         end
       end
      _zyM2L355_pbcCapEn3 = 1'b1;
      _zyM2L324_pbcFsm0_s = 3'b011;
     end
    3'b010:
     // F1, L349
     begin
      // F1, L349
      _zyM2L349_pbcCapEn2 = 1'b0;
      response = _zyL61_iscX2c0_o2;
      if ((response !== 32'b0))
       // F1, L350
       begin
        // F1, L351
        _zyGfifoF0_L324_s3_cbid_1 = _zyGfifo__gfdL351_25_P0_m2_cbid;
        _zyGfifoF0_L324_s3_len_1 = 12'b01;
        _zyGfifoF0_L324_s3_data_1[95:0] = 96'b0;
        _zyGfifoF0_L324_s3_data_1[31:0] = address;
        _zyGfifoF0_L324_s3_req_1 = (_zyGfifo__gfdL351_25_P0_m2_gfOff == _zyGfifoF0_L324_s3_req_1);
// synopsys translate_off
        xc_gfifo_sim(_zyGfifo__gfdL351_25_P0_m2_cbid,32'b01,_zyGfifoF0_L324_s3_data_1);
// synopsys translate_on
        _zyictd_finish_L338_1 = 1'b1;
       end
      _zyM2L355_pbcCapEn3 = 1'b1;
      _zyM2L324_pbcFsm0_s = 3'b011;
     end
    3'b011:
     // F1, L355
     begin
      // F1, L355
      _zyM2L355_pbcCapEn3 = 1'b0;
      _zyM2L324_pbcCapEn0 = 1'b1;
      _zyM2L324_pbcFsm0_s = 3'b0;
     end
   endcase
  end
 end
// F1, L368
always 
 // F1, L368
 begin
  // F1, L416
  @(posedge clk)
   begin
   end
  // F1, L368
  begin:_zyL368_meSwitch4
   reg _zyL368_meEn3;
   // F1, L368
   _zyL368_meEn3 = 1'b1;
   case (_zyL368_meState4)
    1'b0:
     // F1, L368
     begin
      // F1, L368
      // F1, L368
      begin
       // F1, L369
       if ((ready_ib == 32'b01))
        // F1, L369
        begin
         // F1, L207
         // F1, L207
         begin:_zygfifotfiCscp1_L370_ib_service_data_isf_meScp5
          bit [63:0] _zytdata_L207_tfiV5 ;
          bit [31:0] _zytuser_string_L207_tfiV6 ;
          bit [7:0] _zytstrb_L207_tfiV7 ;
          bit [31:0] _zystr_get_L207_tfiV8 ;
          int _zyxr_L207_tfiV9;
          // F0, L0
          _zyxr_L207_tfiV9 = 0;
          if ((_zygsfis_ib_service_data_rptr != _zygsfis_ib_service_data_wptr))
          // F1, L207
          begin
          // F1, L207
          _zyxr_L207_tfiV9[0] = 1'b1;
          {_zytdata_L207_tfiV5,_zytuser_string_L207_tfiV6,_zytstrb_L207_tfiV7,_zystr_get_L207_tfiV8} = _zygsfis_ib_service_data_fifo[_zygsfis_ib_service_data_rptr];
          _zygsfis_ib_service_data_rptr = (_zygsfis_ib_service_data_rptr + 32'b01);
          _zygsfis_ib_service_data_space = (_zygsfis_ib_service_data_space + 32'b01);
          end
          _zyxr_L207_tfiV9[1] = ((_zygsfis_ib_service_data_rptr == _zygsfis_ib_service_data_wptr) & _zygsfis_ib_service_data_eos);
          if (( ~_zyxr_L207_tfiV9[1] ))
          // F1, L207
          begin
          // F1, L207
          if ((_zygsfis_ib_service_data_req == _zygsfis_ib_service_data_ack))
          _zygsfis_ib_service_data_space = ( ~(_zygsfis_ib_service_data_wptr - _zygsfis_ib_service_data_rptr) );
          if ((_zygsfis_ib_service_data_space >= 32'b01000))
          // F0, L0
          begin
          // F0, L0
          _zygsfis_ib_service_data_req = (_zygsfis_ib_service_data_req + 32'b01);
          _zyGfifoF11_L207_data_0 = _zygsfis_ib_service_data_space;
          _zyGfifoF11_L207_req_0 = (_zyGfifo_ib_service_data_2_zyprefetch_m2_gfOff == _zyGfifoF11_L207_req_0);
// synopsys translate_off
          xc_gfifo_sim(_zyGfifo_ib_service_data_2_zyprefetch_m2_cbid,32'b01,_zyGfifoF11_L207_data_0);
// synopsys translate_on
          _zygsfis_ib_service_data_space = 5'b0;
          end
          end
          _zyL370_tfiRv18 = _zyxr_L207_tfiV9;
          tdata_ib = _zytdata_L207_tfiV5;
          tuser_string_ib = _zytuser_string_L207_tfiV6;
          tstrb_ib = _zytstrb_L207_tfiV7;
          str_get_ib = _zystr_get_L207_tfiV8;
         end
         retval_ib = _zyL370_tfiRv18;
         // F1, L517
         begin:_zz_gfdinlCscp2_L372_reverse_translate_tuser_meScp6
          bit [31:0] _zytuser_L517_tfiV1 ;
          // F1, L372
          _zytuser_L517_tfiV1 = tuser_string_ib;
          if ((_zytuser_L517_tfiV1 == 32'b01011))
          // F1, L518
          begin
          // F1, L519
          _zyGfifoF0_L368_s2_cbid_4 = _zyGfifo__gfdL519_24_P0_m2_cbid;
          _zyGfifoF0_L368_s2_req_4 = (_zyGfifo__gfdL519_24_P0_m2_gfOff == _zyGfifoF0_L368_s2_req_4);
// synopsys translate_off
          xc_gfifo_sim(_zyGfifo__gfdL519_24_P0_m2_cbid,32'b0,_zyGfifo_mod2_simData);
// synopsys translate_on
          _zyL372_tfiRv5 = 25'b010100110110111101010100;
          end
          else
          if ((_zytuser_L517_tfiV1 == 32'b01010))
          // F1, L521
          begin
          // F1, L522
          _zyGfifoF0_L368_s2_cbid_4 = _zyGfifo__gfdL522_23_P0_m2_cbid;
          _zyGfifoF0_L368_s2_req_4 = (_zyGfifo__gfdL522_23_P0_m2_gfOff == _zyGfifoF0_L368_s2_req_4);
// synopsys translate_off
          xc_gfifo_sim(_zyGfifo__gfdL522_23_P0_m2_cbid,32'b0,_zyGfifo_mod2_simData);
// synopsys translate_on
          _zyL372_tfiRv5 = 25'b010001010110111101010100;
          end
          else
          // F1, L524
          begin
          // F1, L525
          _zyL372_tfiRv5 = 25'b0;
          end
         end
         user_string_ib = _zyL372_tfiRv5;
         _zyGfifoF14_L373_data_0 = user_string_ib;
         _zyGfifoF14_L373_req_0 = (_zyGfifo__gfdL373_22_P0_m2_gfOff == _zyGfifoF14_L373_req_0);
// synopsys translate_off
         xc_gfifo_sim(_zyGfifo__gfdL373_22_P0_m2_cbid,32'b01,_zyGfifoF14_L373_data_0);
// synopsys translate_on
         if ((retval_ib == 1))
          // F1, L374
          begin
          // F1, L375
          _zyGfifoF15_L375_data_0[135:72] = tdata_ib;
          _zyGfifoF15_L375_data_0[71:40] = tuser_string_ib;
          _zyGfifoF15_L375_data_0[39:32] = tstrb_ib;
          _zyGfifoF15_L375_data_0[31:0] = str_get_ib;
          _zyGfifoF15_L375_req_0 = (_zyGfifo__gfdL375_21_P0_m2_gfOff == _zyGfifoF15_L375_req_0);
// synopsys translate_off
          xc_gfifo_sim(_zyGfifo__gfdL375_21_P0_m2_cbid,32'b0101,_zyGfifoF15_L375_data_0);
// synopsys translate_on
          if ((kme_ib_tready === 1'b1))
          // F1, L376
          begin
          // F1, L377
          kme_ib_tlast <= 1'b0;
          kme_ib_tvalid <= 1'b0;
          if ((str_get_ib == 32'b011))
          // F1, L379
          begin
          // F1, L380
          if (((user_string_ib == 25'b010100110110111101010100) && (tdata_ib[7:0] >= 8'b010101)))
          // F1, L380
          begin
          // F1, L381
          _zyGfifoF16_L381_req_0 = (_zyGfifo__gfdL381_20_P0_m2_gfOff == _zyGfifoF16_L381_req_0);
// synopsys translate_off
          xc_gfifo_sim(_zyGfifo__gfdL381_20_P0_m2_cbid,32'b0,_zyGfifo_mod2_simData);
// synopsys translate_on
          saw_mega = 1'b1;
          end
          else
          if ((tdata_ib[7:0] == 8'b01010))
          // F1, L384
          begin
          // F1, L385
          saw_guid_tlv = 1'b1;
          end
          if ((saw_mega == 32'b01))
          // F1, L387
          begin
          // F1, L388
          mega_tlv_word_count = (mega_tlv_word_count + 1);
          if ((mega_tlv_word_count == 2))
          // F1, L389
          begin
          // F1, L390
          _zyGfifoF17_L390_data_0 = tdata_ib;
          _zyGfifoF17_L390_req_0 = (_zyGfifo__gfdL390_19_P0_m2_gfOff == _zyGfifoF17_L390_req_0);
// synopsys translate_off
          xc_gfifo_sim(_zyGfifo__gfdL390_19_P0_m2_cbid,32'b010,_zyGfifoF17_L390_data_0);
// synopsys translate_on
          if ((tdata_ib[4] == 32'b01))
          // F1, L391
          begin
          // F1, L392
          have_guid_tlv = 1'b1;
          end
          end
          end
          if (((user_string_ib == 25'b010001010110111101010100) && (saw_mega == 32'b01)))
          // F1, L396
          begin
          // F1, L397
          if ((have_guid_tlv == 32'b0))
          // F1, L397
          begin
          // F1, L398
          kme_ib_tlast <= 1'b1;
          end
          saw_mega = 1'b0;
          end
          else
          if (((user_string_ib == 25'b010001010110111101010100) && (saw_guid_tlv == 32'b01)))
          // F1, L402
          begin
          // F1, L403
          kme_ib_tlast <= 1'b1;
          saw_guid_tlv = 1'b0;
          end
          // F1, L529
          begin:_zz_gfdinlCscp3_L406_translate_tuser_t_meScp7
          bit [24:0] _zytuser_L529_tfiV3 ;
          // F1, L406
          _zytuser_L529_tfiV3 = user_string_ib;
          _zyGfifoF18_L530_data_0 = _zytuser_L529_tfiV3;
          _zyGfifoF18_L530_req_0 = (_zyGfifo__gfdL530_18_P0_m2_gfOff == _zyGfifoF18_L530_req_0);
// synopsys translate_off
          xc_gfifo_sim(_zyGfifo__gfdL530_18_P0_m2_cbid,32'b01,_zyGfifoF18_L530_data_0);
// synopsys translate_on
          if ((_zytuser_L529_tfiV3 == 25'b010100110110111101010100))
          // F1, L531
          begin
          // F1, L532
          _zyL406_tfiRv6 = 8'b01;
          end
          else
          if ((_zytuser_L529_tfiV3 == 25'b010001010110111101010100))
          // F1, L533
          begin
          // F1, L534
          _zyL406_tfiRv6 = 8'b010;
          end
          else
          // F1, L535
          begin
          // F1, L536
          _zyL406_tfiRv6 = 8'b011;
          end
          end
          kme_ib_tuser <= _zyL406_tfiRv6;
          end
          else
          // F1, L407
          begin
          // F1, L408
          kme_ib_tuser <= 8'b0;
          end
          kme_ib_tvalid <= 1'b1;
          kme_ib_tdata <= tdata_ib;
          _zyGfifoF19_L412_data_0 = tstrb_ib;
          _zyGfifoF19_L412_req_0 = (_zyGfifo__gfdL412_17_P0_m2_gfOff == _zyGfifoF19_L412_req_0);
// synopsys translate_off
          xc_gfifo_sim(_zyGfifo__gfdL412_17_P0_m2_cbid,32'b01,_zyGfifoF19_L412_data_0);
// synopsys translate_on
          kme_ib_tstrb <= tstrb_ib;
          end
          _zyL368_meState4 = 1'b1;
          _zyL368_meEn3 = 1'b0;
          end
        end
      end
      if (_zyL368_meEn3)
       // F1, L368
       begin
        // F1, L368
        // F1, L368
        begin
         // F1, L368
         _zyL368_meState4 = 1'b0;
        end
       end
     end
    1'b1:
     // F1, L368
     begin
      // F1, L368
      _zyL368_meState4 = 1'b0;
     end
   endcase
  end
 end
// F1, L439
always 
 // F1, L439
 begin
  // F1, L500
  @(posedge clk)
   begin
   end
  // F1, L439
  begin:_zyL439_meSwitch8
   reg _zyL439_meEn4;
   // F1, L439
   _zyL439_meEn4 = 1'b1;
   case (_zyL439_meState8)
    2'b0:
     // F1, L439
     begin
      // F1, L439
      // F1, L439
      begin
       // F1, L440
       if ((ready_ob == 32'b01))
        // F1, L440
        begin
         // F1, L209
         // F1, L209
         begin:_zygfifotfiCscp2_L441_ob_service_data_isf_meScp9
          bit [63:0] _zytdata_L209_tfiV11 ;
          bit [31:0] _zytuser_string_L209_tfiV12 ;
          bit [7:0] _zytstrb_L209_tfiV13 ;
          bit [31:0] _zystr_get_L209_tfiV14 ;
          int _zyxr_L209_tfiV15;
          // F0, L0
          _zyxr_L209_tfiV15 = 0;
          if ((_zygsfis_ob_service_data_rptr != _zygsfis_ob_service_data_wptr))
          // F1, L209
          begin
          // F1, L209
          _zyxr_L209_tfiV15[0] = 1'b1;
          {_zytdata_L209_tfiV11,_zytuser_string_L209_tfiV12,_zytstrb_L209_tfiV13,_zystr_get_L209_tfiV14} = _zygsfis_ob_service_data_fifo[_zygsfis_ob_service_data_rptr];
          _zygsfis_ob_service_data_rptr = (_zygsfis_ob_service_data_rptr + 32'b01);
          _zygsfis_ob_service_data_space = (_zygsfis_ob_service_data_space + 32'b01);
          end
          _zyxr_L209_tfiV15[1] = ((_zygsfis_ob_service_data_rptr == _zygsfis_ob_service_data_wptr) & _zygsfis_ob_service_data_eos);
          if (( ~_zyxr_L209_tfiV15[1] ))
          // F1, L209
          begin
          // F1, L209
          if ((_zygsfis_ob_service_data_req == _zygsfis_ob_service_data_ack))
          _zygsfis_ob_service_data_space = ( ~(_zygsfis_ob_service_data_wptr - _zygsfis_ob_service_data_rptr) );
          if ((_zygsfis_ob_service_data_space >= 32'b01000))
          // F0, L0
          begin
          // F0, L0
          _zygsfis_ob_service_data_req = (_zygsfis_ob_service_data_req + 32'b01);
          _zyGfifoF20_L209_data_0 = _zygsfis_ob_service_data_space;
          _zyGfifoF20_L209_req_0 = (_zyGfifo_ob_service_data_2_zyprefetch_m2_gfOff == _zyGfifoF20_L209_req_0);
// synopsys translate_off
          xc_gfifo_sim(_zyGfifo_ob_service_data_2_zyprefetch_m2_cbid,32'b01,_zyGfifoF20_L209_data_0);
// synopsys translate_on
          _zygsfis_ob_service_data_space = 5'b0;
          end
          end
          _zyL441_tfiRv19 = _zyxr_L209_tfiV15;
          tdata_ob = _zytdata_L209_tfiV11;
          tuser_string_ob = _zytuser_string_L209_tfiV12;
          tstrb_ob = _zytstrb_L209_tfiV13;
          str_get_ob = _zystr_get_L209_tfiV14;
         end
         retval_ob = _zyL441_tfiRv19;
         // F1, L517
         begin:_zz_gfdinlCscp4_L443_reverse_translate_tuser_meScp10
          bit [31:0] _zytuser_L517_tfiV1 ;
          // F1, L443
          _zytuser_L517_tfiV1 = tuser_string_ob;
          if ((_zytuser_L517_tfiV1 == 32'b01011))
          // F1, L518
          begin
          // F1, L519
          _zyGfifoF0_L439_s2_cbid_5 = _zyGfifo__gfdL519_16_P0_m2_cbid;
          _zyGfifoF0_L439_s2_req_5 = (_zyGfifo__gfdL519_16_P0_m2_gfOff == _zyGfifoF0_L439_s2_req_5);
// synopsys translate_off
          xc_gfifo_sim(_zyGfifo__gfdL519_16_P0_m2_cbid,32'b0,_zyGfifo_mod2_simData);
// synopsys translate_on
          _zyL443_tfiRv7 = 25'b010100110110111101010100;
          end
          else
          if ((_zytuser_L517_tfiV1 == 32'b01010))
          // F1, L521
          begin
          // F1, L522
          _zyGfifoF0_L439_s2_cbid_5 = _zyGfifo__gfdL522_15_P0_m2_cbid;
          _zyGfifoF0_L439_s2_req_5 = (_zyGfifo__gfdL522_15_P0_m2_gfOff == _zyGfifoF0_L439_s2_req_5);
// synopsys translate_off
          xc_gfifo_sim(_zyGfifo__gfdL522_15_P0_m2_cbid,32'b0,_zyGfifo_mod2_simData);
// synopsys translate_on
          _zyL443_tfiRv7 = 25'b010001010110111101010100;
          end
          else
          // F1, L524
          begin
          // F1, L525
          _zyL443_tfiRv7 = 25'b0;
          end
         end
         user_string_ob = _zyL443_tfiRv7;
         _zyGfifoF23_L444_data_0 = user_string_ob;
         _zyGfifoF23_L444_req_0 = (_zyGfifo__gfdL444_14_P0_m2_gfOff == _zyGfifoF23_L444_req_0);
// synopsys translate_off
         xc_gfifo_sim(_zyGfifo__gfdL444_14_P0_m2_cbid,32'b01,_zyGfifoF23_L444_data_0);
// synopsys translate_on
         if ((retval_ob == 1))
          // F1, L445
          begin
          // F1, L446
          _zyGfifoF24_L446_data_0[135:72] = tdata_ob;
          _zyGfifoF24_L446_data_0[71:40] = tuser_string_ob;
          _zyGfifoF24_L446_data_0[39:32] = tstrb_ob;
          _zyGfifoF24_L446_data_0[31:0] = str_get_ob;
          _zyGfifoF24_L446_req_0 = (_zyGfifo__gfdL446_13_P0_m2_gfOff == _zyGfifoF24_L446_req_0);
// synopsys translate_off
          xc_gfifo_sim(_zyGfifo__gfdL446_13_P0_m2_cbid,32'b0101,_zyGfifoF24_L446_data_0);
// synopsys translate_on
          if ((kme_ob_tvalid === 1'b0))
          // F1, L448
          begin
          // F1, L449
          _zyL439_meState8 = 2'b01;
          _zyL439_meEn4 = 1'b0;
          end
          if (_zyL439_meEn4)
          // F1, L457
          begin
          // F1, L457
          watchdog_timer = 0;
          tlast = 1'b0;
          ignore_compare_result = 1'b0;
          _zyGfifoF25_L460_data_0 = kme_ob_tdata;
          _zyGfifoF25_L460_req_0 = (_zyGfifo__gfdL460_12_P0_m2_gfOff == _zyGfifoF25_L460_req_0);
// synopsys translate_off
          xc_gfifo_sim(_zyGfifo__gfdL460_12_P0_m2_cbid,32'b010,_zyGfifoF25_L460_data_0);
// synopsys translate_on
          if ((str_get_ob == 32'b011))
          // F1, L461
          begin
          // F1, L529
          // F1, L529
          begin:_zz_gfdinlCscp5_L462_translate_tuser_t_meScp11
          bit [24:0] _zytuser_L529_tfiV3 ;
          // F1, L462
          _zytuser_L529_tfiV3 = user_string_ob;
          _zyGfifoF26_L530_data_0 = _zytuser_L529_tfiV3;
          _zyGfifoF26_L530_req_0 = (_zyGfifo__gfdL530_11_P0_m2_gfOff == _zyGfifoF26_L530_req_0);
// synopsys translate_off
          xc_gfifo_sim(_zyGfifo__gfdL530_11_P0_m2_cbid,32'b01,_zyGfifoF26_L530_data_0);
// synopsys translate_on
          if ((_zytuser_L529_tfiV3 == 25'b010100110110111101010100))
          // F1, L531
          begin
          // F1, L532
          _zyL462_tfiRv8 = 8'b01;
          end
          else
          if ((_zytuser_L529_tfiV3 == 25'b010001010110111101010100))
          // F1, L533
          begin
          // F1, L534
          _zyL462_tfiRv8 = 8'b010;
          end
          else
          // F1, L535
          begin
          // F1, L536
          _zyL462_tfiRv8 = 8'b011;
          end
          end
          tuser = _zyL462_tfiRv8;
          if (((user_string_ob == 25'b010100110110111101010100) && (tdata_ob[7:0] == 8'b01001)))
          // F1, L463
          begin
          // F1, L464
          saw_cqe = 1'b1;
          end
          if ((user_string_ob == 25'b010001010110111101010100))
          // F1, L466
          begin
          // F1, L467
          tlast = 1'b1;
          saw_cqe = 1'b0;
          end
          if (((user_string_ob == 25'b010100110110111101010100) && (tdata_ob[7:0] == 8'b01000)))
          // F1, L470
          begin
          // F1, L471
          saw_stats = 1'b1;
          end
          if (((user_string_ob == 25'b010001010110111101010100) && (saw_stats == 32'b01)))
          // F1, L473
          begin
          // F1, L474
          ignore_compare_result = 1'b1;
          saw_stats = 1'b0;
          end
          end
          else
          // F1, L477
          begin
          // F1, L478
          tuser = 8'b0;
          end
          _zyGfifoF27_L480_data_0 = tuser;
          _zyGfifoF27_L480_req_0 = (_zyGfifo__gfdL480_10_P0_m2_gfOff == _zyGfifoF27_L480_req_0);
// synopsys translate_off
          xc_gfifo_sim(_zyGfifo__gfdL480_10_P0_m2_cbid,32'b01,_zyGfifoF27_L480_data_0);
// synopsys translate_on
          if (((kme_ob_tdata !== tdata_ob) && (ignore_compare_result == 32'b0)))
          // F1, L481
          begin
          // F1, L482
          _zyGfifoF28_L482_data_0[127:64] = kme_ob_tdata;
          _zyGfifoF28_L482_data_0[63:0] = tdata_ob;
          _zyGfifoF28_L482_req_0 = (_zyGfifo__gfdL482_9_P0_m2_gfOff == _zyGfifoF28_L482_req_0);
// synopsys translate_off
          xc_gfifo_sim(_zyGfifo__gfdL482_9_P0_m2_cbid,32'b0100,_zyGfifoF28_L482_data_0);
// synopsys translate_on
          error_cntr = (error_cntr + 1);
          end
          if ((kme_ob_tuser !== tuser))
          // F1, L486
          begin
          // F1, L487
          _zyGfifoF29_L487_data_0[15:8] = kme_ob_tuser;
          _zyGfifoF29_L487_data_0[7:0] = tuser;
          _zyGfifoF29_L487_req_0 = (_zyGfifo__gfdL487_8_P0_m2_gfOff == _zyGfifoF29_L487_req_0);
// synopsys translate_off
          xc_gfifo_sim(_zyGfifo__gfdL487_8_P0_m2_cbid,32'b01,_zyGfifoF29_L487_data_0);
// synopsys translate_on
          error_cntr = (error_cntr + 1);
          end
          if ((kme_ob_tstrb !== tstrb_ob))
          // F1, L490
          begin
          // F1, L491
          _zyGfifoF30_L491_data_0[15:8] = kme_ob_tstrb;
          _zyGfifoF30_L491_data_0[7:0] = tstrb_ob;
          _zyGfifoF30_L491_req_0 = (_zyGfifo__gfdL491_7_P0_m2_gfOff == _zyGfifoF30_L491_req_0);
// synopsys translate_off
          xc_gfifo_sim(_zyGfifo__gfdL491_7_P0_m2_cbid,32'b01,_zyGfifoF30_L491_data_0);
// synopsys translate_on
          error_cntr = (error_cntr + 1);
          end
          if ((kme_ob_tlast !== tlast))
          // F1, L495
          begin
          // F1, L496
          _zyGfifoF31_L496_data_0[8] = kme_ob_tlast;
          _zyGfifoF31_L496_data_0[0] = tlast;
          _zyGfifoF31_L496_req_0 = (_zyGfifo__gfdL496_6_P0_m2_gfOff == _zyGfifoF31_L496_req_0);
// synopsys translate_off
          xc_gfifo_sim(_zyGfifo__gfdL496_6_P0_m2_cbid,32'b01,_zyGfifoF31_L496_data_0);
// synopsys translate_on
          error_cntr = (error_cntr + 1);
          end
          end
          end
         if (_zyL439_meEn4)
          // F1, L500
          begin
          // F1, L500
          _zyL439_meState8 = 2'b10;
          _zyL439_meEn4 = 1'b0;
          end
        end
      end
      if (_zyL439_meEn4)
       // F1, L439
       begin
        // F1, L439
        // F1, L439
        begin
         // F1, L439
         _zyL439_meState8 = 2'b0;
        end
       end
     end
    2'b01:
     // F1, L450
     begin
      // F1, L450
      watchdog_timer = (watchdog_timer + 1);
      if ((watchdog_timer > 10000))
       // F1, L451
       begin
        // F1, L452
        error_cntr = (error_cntr + 1);
        $display("\nOUTBOUND_ERROR:  @time:%-d  Watchdog timer EXPIRED!\n",$time);
        _zyictd_finish_L454_2 = 1'b1;
       end
      if ((kme_ob_tvalid === 1'b0))
       // F1, L448
       begin
        // F1, L449
        _zyL439_meState8 = 2'b01;
        _zyL439_meEn4 = 1'b0;
       end
      if (_zyL439_meEn4)
       // F1, L457
       begin
        // F1, L457
        watchdog_timer = 0;
        tlast = 1'b0;
        ignore_compare_result = 1'b0;
        _zyGfifoF25_L460_data_0 = kme_ob_tdata;
        _zyGfifoF25_L460_req_0 = (_zyGfifo__gfdL460_12_P0_m2_gfOff == _zyGfifoF25_L460_req_0);
// synopsys translate_off
        xc_gfifo_sim(_zyGfifo__gfdL460_12_P0_m2_cbid,32'b010,_zyGfifoF25_L460_data_0);
// synopsys translate_on
        if ((str_get_ob == 32'b011))
         // F1, L461
         begin
          // F1, L529
          // F1, L529
          begin:_zz_gfdinlCscp5_L462_translate_tuser_t_meScp12
          bit [24:0] _zytuser_L529_tfiV3 ;
          // F1, L462
          _zytuser_L529_tfiV3 = user_string_ob;
          _zyGfifoF26_L530_data_0 = _zytuser_L529_tfiV3;
          _zyGfifoF26_L530_req_0 = (_zyGfifo__gfdL530_11_P0_m2_gfOff == _zyGfifoF26_L530_req_0);
// synopsys translate_off
          xc_gfifo_sim(_zyGfifo__gfdL530_11_P0_m2_cbid,32'b01,_zyGfifoF26_L530_data_0);
// synopsys translate_on
          if ((_zytuser_L529_tfiV3 == 25'b010100110110111101010100))
          // F1, L531
          begin
          // F1, L532
          _zyL462_tfiRv8 = 8'b01;
          end
          else
          if ((_zytuser_L529_tfiV3 == 25'b010001010110111101010100))
          // F1, L533
          begin
          // F1, L534
          _zyL462_tfiRv8 = 8'b010;
          end
          else
          // F1, L535
          begin
          // F1, L536
          _zyL462_tfiRv8 = 8'b011;
          end
          end
          tuser = _zyL462_tfiRv8;
          if (((user_string_ob == 25'b010100110110111101010100) && (tdata_ob[7:0] == 8'b01001)))
          // F1, L463
          begin
          // F1, L464
          saw_cqe = 1'b1;
          end
          if ((user_string_ob == 25'b010001010110111101010100))
          // F1, L466
          begin
          // F1, L467
          tlast = 1'b1;
          saw_cqe = 1'b0;
          end
          if (((user_string_ob == 25'b010100110110111101010100) && (tdata_ob[7:0] == 8'b01000)))
          // F1, L470
          begin
          // F1, L471
          saw_stats = 1'b1;
          end
          if (((user_string_ob == 25'b010001010110111101010100) && (saw_stats == 32'b01)))
          // F1, L473
          begin
          // F1, L474
          ignore_compare_result = 1'b1;
          saw_stats = 1'b0;
          end
         end
        else
         // F1, L477
         begin
          // F1, L478
          tuser = 8'b0;
         end
        _zyGfifoF27_L480_data_0 = tuser;
        _zyGfifoF27_L480_req_0 = (_zyGfifo__gfdL480_10_P0_m2_gfOff == _zyGfifoF27_L480_req_0);
// synopsys translate_off
        xc_gfifo_sim(_zyGfifo__gfdL480_10_P0_m2_cbid,32'b01,_zyGfifoF27_L480_data_0);
// synopsys translate_on
        if (((kme_ob_tdata !== tdata_ob) && (ignore_compare_result == 32'b0)))
         // F1, L481
         begin
          // F1, L482
          _zyGfifoF28_L482_data_0[127:64] = kme_ob_tdata;
          _zyGfifoF28_L482_data_0[63:0] = tdata_ob;
          _zyGfifoF28_L482_req_0 = (_zyGfifo__gfdL482_9_P0_m2_gfOff == _zyGfifoF28_L482_req_0);
// synopsys translate_off
          xc_gfifo_sim(_zyGfifo__gfdL482_9_P0_m2_cbid,32'b0100,_zyGfifoF28_L482_data_0);
// synopsys translate_on
          error_cntr = (error_cntr + 1);
         end
        if ((kme_ob_tuser !== tuser))
         // F1, L486
         begin
          // F1, L487
          _zyGfifoF29_L487_data_0[15:8] = kme_ob_tuser;
          _zyGfifoF29_L487_data_0[7:0] = tuser;
          _zyGfifoF29_L487_req_0 = (_zyGfifo__gfdL487_8_P0_m2_gfOff == _zyGfifoF29_L487_req_0);
// synopsys translate_off
          xc_gfifo_sim(_zyGfifo__gfdL487_8_P0_m2_cbid,32'b01,_zyGfifoF29_L487_data_0);
// synopsys translate_on
          error_cntr = (error_cntr + 1);
         end
        if ((kme_ob_tstrb !== tstrb_ob))
         // F1, L490
         begin
          // F1, L491
          _zyGfifoF30_L491_data_0[15:8] = kme_ob_tstrb;
          _zyGfifoF30_L491_data_0[7:0] = tstrb_ob;
          _zyGfifoF30_L491_req_0 = (_zyGfifo__gfdL491_7_P0_m2_gfOff == _zyGfifoF30_L491_req_0);
// synopsys translate_off
          xc_gfifo_sim(_zyGfifo__gfdL491_7_P0_m2_cbid,32'b01,_zyGfifoF30_L491_data_0);
// synopsys translate_on
          error_cntr = (error_cntr + 1);
         end
        if ((kme_ob_tlast !== tlast))
         // F1, L495
         begin
          // F1, L496
          _zyGfifoF31_L496_data_0[8] = kme_ob_tlast;
          _zyGfifoF31_L496_data_0[0] = tlast;
          _zyGfifoF31_L496_req_0 = (_zyGfifo__gfdL496_6_P0_m2_gfOff == _zyGfifoF31_L496_req_0);
// synopsys translate_off
          xc_gfifo_sim(_zyGfifo__gfdL496_6_P0_m2_cbid,32'b01,_zyGfifoF31_L496_data_0);
// synopsys translate_on
          error_cntr = (error_cntr + 1);
         end
        _zyL439_meState8 = 2'b10;
       end
     end
    2'b10:
     // F1, L439
     begin
      // F1, L439
      _zyL439_meState8 = 2'b0;
     end
   endcase
  end
 end
// F1, L10
initial 
 begin
 end
// F1, L253
always 
 // F1, L253
 begin
  // F1, L253
  @(posedge _zyM2L253_pbcMevClk12)
   begin
   end
  // F1, L253
  begin:_zyM2L253_pbcFsm2
   // F1, L253
   case (_zyM2L253_pbcFsm2_s)
    3'b0:
     // F1, L253
     begin
      // F1, L253
      _zyM2L253_pbcCapEn5 = 1'b0;
      // F1, L253
      begin:_zy_zzblk_0_0_M2L253_pbcScp3
       // F1, L253
       // F1, L253
       begin:_zyifsyneCscp1_L253_M2_pbcScp4
        // F1, L254
        error_cntr = 0;
        rst_n = 1'b0;
        if (_zyictd_sysfunc_11_L257_2)
         // F1, L257
         begin
          // F1, L258
          seed = _zyictd_sysfunc_36_L258_0;
          _zz_58_258_2 = _zyictd_sysfunc_36_L258_1;
         end
        else
         // F1, L259
         begin
          // F1, L260
          seed = 280'b0110001;
         end
        if (_zyictd_sysfunc_11_L263_5)
         // F1, L263
         begin
          // F1, L264
          testname = _zyictd_sysfunc_36_L264_3;
          _zz_58_264_3 = _zyictd_sysfunc_36_L264_4;
          _zyGfifoF0_L253_s4_cbid_6 = _zyGfifo__gfdL265_5_P0_m2_cbid;
          _zyGfifoF0_L253_s4_len_6 = 12'b010010;
          _zyGfifoF0_L253_s4_data_6[559:0] = {560{1'b0}};
          _zyGfifoF0_L253_s4_data_6[559:280] = testname;
          _zyGfifoF0_L253_s4_data_6[279:0] = seed;
          _zyGfifoF0_L253_s4_req_6 = (_zyGfifo__gfdL265_5_P0_m2_gfOff == _zyGfifoF0_L253_s4_req_6);
// synopsys translate_off
          xc_gfifo_sim(_zyGfifo__gfdL265_5_P0_m2_cbid,32'b010010,_zyGfifoF0_L253_s4_data_6);
// synopsys translate_on
         end
        else
         // F1, L266
         begin
          // F1, L267
          testname = 280'b01110101011011100110101101101110011011110111011101101110;
          _zyGfifoF0_L253_s4_cbid_6 = _zyGfifo__gfdL268_4_P0_m2_cbid;
          _zyGfifoF0_L253_s4_len_6 = 12'b010010;
          _zyGfifoF0_L253_s4_data_6[559:0] = {560{1'b0}};
          _zyGfifoF0_L253_s4_data_6[559:280] = 280'b01110101011011100110101101101110011011110111011101101110;
          _zyGfifoF0_L253_s4_data_6[279:0] = seed;
          _zyGfifoF0_L253_s4_req_6 = (_zyGfifo__gfdL268_4_P0_m2_gfOff == _zyGfifoF0_L253_s4_req_6);
// synopsys translate_off
          xc_gfifo_sim(_zyGfifo__gfdL268_4_P0_m2_cbid,32'b010010,_zyGfifoF0_L253_s4_data_6);
// synopsys translate_on
         end
        _zyGfifoF1_L253_s2_cbid_7 = _zyGfifo__gfdL271_3_P0_m2_cbid;
        _zyGfifoF1_L253_s2_req_7 = (_zyGfifo__gfdL271_3_P0_m2_gfOff == _zyGfifoF1_L253_s2_req_7);
// synopsys translate_off
        xc_gfifo_sim(_zyGfifo__gfdL271_3_P0_m2_cbid,32'b0,_zyGfifo_mod2_simData);
// synopsys translate_on
        _zyM2L273_pbcT0 = 125;
        _zyM2L274_pbcCapEn6 = 1'b1;
        _zyM2L253_pbcFsm2_s = 3'b01;
       end
      end
     end
    3'b01:
     // F1, L274
     begin
      // F1, L253
      _zyM2L253_pbcEn14 = 1'b1;
      _zyM2L274_pbcCapEn6 = 1'b0;
      _zyM2L273_pbcT0 = (_zyM2L273_pbcT0 - 32'b01);
      if ((_zyM2L273_pbcT0 > 32'b0))
       // F1, L273
       begin
        // F1, L274
        _zyM2L274_pbcCapEn6 = 1'b1;
        _zyM2L253_pbcFsm2_s = 3'b01;
        _zyM2L253_pbcEn14 = 1'b0;
       end
      if (_zyM2L253_pbcEn14)
       // F1, L276
       begin
        // F1, L276
        _zyGfifoF0_L253_s4_cbid_6 = _zyGfifo__gfdL276_2_P0_m2_cbid;
        _zyGfifoF0_L253_s4_len_6 = 12'b0;
        _zyGfifoF0_L253_s4_data_6[559:0] = {560{1'b0}};
        _zyGfifoF0_L253_s4_req_6 = (_zyGfifo__gfdL276_2_P0_m2_gfOff == _zyGfifoF0_L253_s4_req_6);
// synopsys translate_off
        xc_gfifo_sim(_zyGfifo__gfdL276_2_P0_m2_cbid,32'b0,_zyGfifo_mod2_simData);
// synopsys translate_on
        kme_ib_tid <= 1'b0;
        kme_ib_tvalid <= 1'b0;
        kme_ib_tlast <= 1'b0;
        kme_ib_tdata <= 64'b0;
        kme_ib_tstrb <= 8'b0;
        kme_ib_tuser <= 8'b0;
        kme_ob_tready <= 1'b1;
        _zyM2L286_pbcT1 = 63;
        _zyM2L287_pbcCapEn7 = 1'b1;
        _zyM2L253_pbcFsm2_s = 3'b010;
       end
     end
    3'b010:
     // F1, L287
     begin
      // F1, L253
      _zyM2L253_pbcEn14 = 1'b1;
      _zyM2L287_pbcCapEn7 = 1'b0;
      _zyM2L286_pbcT1 = (_zyM2L286_pbcT1 - 32'b01);
      if ((_zyM2L286_pbcT1 > 32'b0))
       // F1, L286
       begin
        // F1, L287
        _zyM2L287_pbcCapEn7 = 1'b1;
        _zyM2L253_pbcFsm2_s = 3'b010;
        _zyM2L253_pbcEn14 = 1'b0;
       end
      if (_zyM2L253_pbcEn14)
       // F1, L289
       begin
        // F1, L289
        _zyGfifoF1_L253_s2_cbid_7 = _zyGfifo__gfdL289_1_P0_m2_cbid;
        _zyGfifoF1_L253_s2_req_7 = (_zyGfifo__gfdL289_1_P0_m2_gfOff == _zyGfifoF1_L253_s2_req_7);
// synopsys translate_off
        xc_gfifo_sim(_zyGfifo__gfdL289_1_P0_m2_cbid,32'b0,_zyGfifo_mod2_simData);
// synopsys translate_on
        rst_n = 1'b1;
        _zyM2L292_pbcT2 = 125;
        _zyM2L293_pbcCapEn8 = 1'b1;
        _zyM2L253_pbcFsm2_s = 3'b011;
       end
     end
    3'b011:
     // F1, L293
     begin
      // F1, L253
      _zyM2L253_pbcEn14 = 1'b1;
      _zyM2L293_pbcCapEn8 = 1'b0;
      _zyM2L292_pbcT2 = (_zyM2L292_pbcT2 - 32'b01);
      if ((_zyM2L292_pbcT2 > 32'b0))
       // F1, L292
       begin
        // F1, L293
        _zyM2L293_pbcCapEn8 = 1'b1;
        _zyM2L253_pbcFsm2_s = 3'b011;
        _zyM2L253_pbcEn14 = 1'b0;
       end
      if (_zyM2L253_pbcEn14)
       // F1, L295
       begin
        // F1, L295
        _zyM2L295_pbcCapEn9 = 1'b1;
        _zyM2L253_pbcFsm2_s = 3'b100;
       end
     end
    3'b100:
     // F1, L295
     begin
      // F1, L295
      _zyM2L295_pbcCapEn9 = 1'b0;
      // F1, L362
      begin:_zyifsyneCscp0_L296_do_kme_config_M2_pbcScp5
       // F1, L363
       config_ready = 1'b1;
       _zyM2L364_pbcCapEn10 = 1'b1;
       _zyM2L253_pbcFsm2_s = 3'b101;
      end
     end
    3'b101:
     // F1, L364
     begin
      // F1, L364
      _zyM2L364_pbcCapEn10 = 1'b0;
      _zyGfifoF0_L253_s4_cbid_6 = _zyGfifo__gfdL365_0_P0_m2_cbid;
      _zyGfifoF0_L253_s4_len_6 = 12'b0;
      _zyGfifoF0_L253_s4_data_6[559:0] = {560{1'b0}};
      _zyGfifoF0_L253_s4_req_6 = (_zyGfifo__gfdL365_0_P0_m2_gfOff == _zyGfifoF0_L253_s4_req_6);
// synopsys translate_off
      xc_gfifo_sim(_zyGfifo__gfdL365_0_P0_m2_cbid,32'b0,_zyGfifo_mod2_simData);
// synopsys translate_on
      config_done = 1'b1;
      _zyM2L299_pbcT3 = 13;
      _zyM2L300_pbcCapEn11 = 1'b1;
      _zyM2L253_pbcFsm2_s = 3'b110;
     end
    3'b110:
     // F1, L300
     begin
      // F1, L253
      _zyM2L253_pbcEn14 = 1'b1;
      _zyM2L300_pbcCapEn11 = 1'b0;
      _zyM2L299_pbcT3 = (_zyM2L299_pbcT3 - 32'b01);
      if ((_zyM2L299_pbcT3 > 32'b0))
       // F1, L299
       begin
        // F1, L300
        _zyM2L300_pbcCapEn11 = 1'b1;
        _zyM2L253_pbcFsm2_s = 3'b110;
        _zyM2L253_pbcEn14 = 1'b0;
       end
      if (_zyM2L253_pbcEn14)
       // F0, L0
       begin
        // F0, L0
        _zyixc_port_0_0_ack = ( ~_zyixc_port_0_0_ack );
        _zyM2L253_pbcCapEn5 = 1'b1;
        _zyM2L253_pbcFsm2_s = 3'b0;
       end
     end
   endcase
  end
 end

  import "DPI-C" context function int xctf_register_task(input int channel, input string name, input int exportTF, int isFunc, int openarr, input int partitionId, input int mid, input int iwidth, input int owidth, input string file, input int line);
  import "DPI-C" context function void xctf_register_port_task(input int channel, input int lpid, input int ltid, input int gtid);
  import "DPI-C" context function void xctf_register_port_marg(input int channel, input int lpid, input int lmargid, input string memspec);
  import "DPI-C" context function int xctf_define_port_task_n_marg_reg_call(input int channel, input int lpid, input int piomem, input int s2hwidth, input int h2swidth, input int lmargCnt, input int ltidwidth, input int ltid, input int gtid, input int lmargid, input string memspec);

  function bit do_sf_init;
    static bit [15:0] _zyifsyn_tb_task_2_xpt_gtid = xctf_register_task(0, "_zyifsyn_tb_task_2_xpt", 1, 0, 0, 0, 2, 0, 0, "/home/ibarry/Project-Zipline-master/dv/KME/run/kme_tb.sv", 253);
    integer _zyport_0_0_gpid;
    begin
      _zyport_0_0_gpid = xctf_define_port_task_n_marg_reg_call(0, 0, 1, 0, 0, 0, 0, 0, _zyifsyn_tb_task_2_xpt_gtid, 0, "");
      IXC_GFIFO.OSF.OSF_create_wait_event(_zyport_0_0_gpid);
      return 0;
    end
  endfunction

  const bit _zydummy_do_init = do_sf_init();

// F1, L206
always 
 @(posedge _zySfifoF0_call)
  // F1, L206
  begin
   // F1, L206
   // F1, L206
   begin:_zypbctfiCscp0_L206_get_config_data_zyackf_2_call
    int _zyeos_L206_tfiV0;
    // F1, L206
    _zyeos_L206_tfiV0 = _zySfifoF0_iarg[31:0];
    _zygsfis_get_config_data_ack = (_zygsfis_get_config_data_ack + 32'b01);
    _zygsfis_get_config_data_eos = _zyeos_L206_tfiV0;
   end
  end
// F1, L206
always 
 @(posedge _zySfifoF1_call)
  // F1, L206
  begin
   // F1, L206
   // F1, L206
   begin:_zypbctfiCscp1_L206_get_config_data_zyputf_2_call
    bit [7:0] _zyoperation_L206_tfiV2 ;
    bit [31:0] _zyaddress_L206_tfiV3 ;
    bit [31:0] _zydata_L206_tfiV4 ;
    // F1, L206
    _zyoperation_L206_tfiV2 = _zySfifoF1_iarg[7:0];
    _zyaddress_L206_tfiV3 = _zySfifoF1_iarg[39:8];
    _zydata_L206_tfiV4 = _zySfifoF1_iarg[71:40];
    _zygsfis_get_config_data_fifo[_zygsfis_get_config_data_wptr] = {_zyoperation_L206_tfiV2,_zyaddress_L206_tfiV3,_zydata_L206_tfiV4};
    _zygsfis_get_config_data_wptr = (_zygsfis_get_config_data_wptr + 32'b01);
   end
  end
// F1, L207
always 
 @(posedge _zySfifoF2_call)
  // F1, L207
  begin
   // F1, L207
   // F1, L207
   begin:_zypbctfiCscp2_L207_ib_service_data_zyackf_2_call
    int _zyeos_L207_tfiV6;
    // F1, L207
    _zyeos_L207_tfiV6 = _zySfifoF2_iarg[31:0];
    _zygsfis_ib_service_data_ack = (_zygsfis_ib_service_data_ack + 32'b01);
    _zygsfis_ib_service_data_eos = _zyeos_L207_tfiV6;
   end
  end
// F1, L207
always 
 @(posedge _zySfifoF3_call)
  // F1, L207
  begin
   // F1, L207
   // F1, L207
   begin:_zypbctfiCscp3_L207_ib_service_data_zyputf_2_call
    bit [63:0] _zytdata_L207_tfiV8 ;
    bit [31:0] _zytuser_string_L207_tfiV9 ;
    bit [7:0] _zytstrb_L207_tfiV10 ;
    bit [31:0] _zystr_get_L207_tfiV11 ;
    // F1, L207
    _zytdata_L207_tfiV8 = _zySfifoF3_iarg[63:0];
    _zytuser_string_L207_tfiV9 = _zySfifoF3_iarg[95:64];
    _zytstrb_L207_tfiV10 = _zySfifoF3_iarg[103:96];
    _zystr_get_L207_tfiV11 = _zySfifoF3_iarg[135:104];
    _zygsfis_ib_service_data_fifo[_zygsfis_ib_service_data_wptr] = {_zytdata_L207_tfiV8,_zytuser_string_L207_tfiV9,_zytstrb_L207_tfiV10,_zystr_get_L207_tfiV11};
    _zygsfis_ib_service_data_wptr = (_zygsfis_ib_service_data_wptr + 32'b01);
   end
  end
// F1, L209
always 
 @(posedge _zySfifoF4_call)
  // F1, L209
  begin
   // F1, L209
   // F1, L209
   begin:_zypbctfiCscp4_L209_ob_service_data_zyackf_2_call
    int _zyeos_L209_tfiV13;
    // F1, L209
    _zyeos_L209_tfiV13 = _zySfifoF4_iarg[31:0];
    _zygsfis_ob_service_data_ack = (_zygsfis_ob_service_data_ack + 32'b01);
    _zygsfis_ob_service_data_eos = _zyeos_L209_tfiV13;
   end
  end
// F1, L209
always 
 @(posedge _zySfifoF5_call)
  // F1, L209
  begin
   // F1, L209
   // F1, L209
   begin:_zypbctfiCscp5_L209_ob_service_data_zyputf_2_call
    bit [63:0] _zytdata_L209_tfiV15 ;
    bit [31:0] _zytuser_string_L209_tfiV16 ;
    bit [7:0] _zytstrb_L209_tfiV17 ;
    bit [31:0] _zystr_get_L209_tfiV18 ;
    // F1, L209
    _zytdata_L209_tfiV15 = _zySfifoF5_iarg[63:0];
    _zytuser_string_L209_tfiV16 = _zySfifoF5_iarg[95:64];
    _zytstrb_L209_tfiV17 = _zySfifoF5_iarg[103:96];
    _zystr_get_L209_tfiV18 = _zySfifoF5_iarg[135:104];
    _zygsfis_ob_service_data_fifo[_zygsfis_ob_service_data_wptr] = {_zytdata_L209_tfiV15,_zytuser_string_L209_tfiV16,_zytstrb_L209_tfiV17,_zystr_get_L209_tfiV18};
    _zygsfis_ob_service_data_wptr = (_zygsfis_ob_service_data_wptr + 32'b01);
   end
  end

import "DPI-C" context function
  int xc_sfifo_new(input string fn, input string portName, int umodId, int partitionId, int iargL, int oargL, int oargC, int noflush, int gargL, int forceToSvChannel);

export "DPI-C" function xc_sfifo_mod_id;
function int xc_sfifo_mod_id; return 2; endfunction

export "DPI-C" function xc_sfifo_partition_id;
function int xc_sfifo_partition_id; return 0; endfunction

export "DPI-C" function get_config_data_zyackf_m2p0_sim;
const int _zySfifoF0_get_config_data_zyackf_tid_sz = 0;
const bit [21:0] _zySfifoF0_get_config_data_zyackf_tid_cv = xc_sfifo_new("get_config_data_zyackf", "_zzSfifoF0_L206_p", 2, 0, 1, 0, 0, 1, _zySfifoF0_get_config_data_zyackf_tid_sz, 0);
initial _zySfifoF0_get_config_data_zyackf_tid = _zySfifoF0_get_config_data_zyackf_tid_cv;

export "DPI-C" function get_config_data_zyputf_m2p0_sim;
const int _zySfifoF1_get_config_data_zyputf_tid_sz = 0;
const bit [21:0] _zySfifoF1_get_config_data_zyputf_tid_cv = xc_sfifo_new("get_config_data_zyputf", "_zzSfifoF1_L206_p", 2, 0, 3, 0, 0, 1, _zySfifoF1_get_config_data_zyputf_tid_sz, 0);
initial _zySfifoF1_get_config_data_zyputf_tid = _zySfifoF1_get_config_data_zyputf_tid_cv;

export "DPI-C" function ib_service_data_zyackf_m2p0_sim;
const int _zySfifoF2_ib_service_data_zyackf_tid_sz = 0;
const bit [21:0] _zySfifoF2_ib_service_data_zyackf_tid_cv = xc_sfifo_new("ib_service_data_zyackf", "_zzSfifoF2_L207_p", 2, 0, 1, 0, 0, 1, _zySfifoF2_ib_service_data_zyackf_tid_sz, 0);
initial _zySfifoF2_ib_service_data_zyackf_tid = _zySfifoF2_ib_service_data_zyackf_tid_cv;

export "DPI-C" function ib_service_data_zyputf_m2p0_sim;
const int _zySfifoF3_ib_service_data_zyputf_tid_sz = 0;
const bit [21:0] _zySfifoF3_ib_service_data_zyputf_tid_cv = xc_sfifo_new("ib_service_data_zyputf", "_zzSfifoF3_L207_p", 2, 0, 5, 0, 0, 1, _zySfifoF3_ib_service_data_zyputf_tid_sz, 0);
initial _zySfifoF3_ib_service_data_zyputf_tid = _zySfifoF3_ib_service_data_zyputf_tid_cv;

export "DPI-C" function ob_service_data_zyackf_m2p0_sim;
const int _zySfifoF4_ob_service_data_zyackf_tid_sz = 0;
const bit [21:0] _zySfifoF4_ob_service_data_zyackf_tid_cv = xc_sfifo_new("ob_service_data_zyackf", "_zzSfifoF4_L209_p", 2, 0, 1, 0, 0, 1, _zySfifoF4_ob_service_data_zyackf_tid_sz, 0);
initial _zySfifoF4_ob_service_data_zyackf_tid = _zySfifoF4_ob_service_data_zyackf_tid_cv;

export "DPI-C" function ob_service_data_zyputf_m2p0_sim;
const int _zySfifoF5_ob_service_data_zyputf_tid_sz = 0;
const bit [21:0] _zySfifoF5_ob_service_data_zyputf_tid_cv = xc_sfifo_new("ob_service_data_zyputf", "_zzSfifoF5_L209_p", 2, 0, 5, 0, 0, 1, _zySfifoF5_ob_service_data_zyputf_tid_sz, 0);
initial _zySfifoF5_ob_service_data_zyputf_tid = _zySfifoF5_ob_service_data_zyputf_tid_cv;

// F1, L10
initial 
 // F1, L10
 begin
  // F2, L94
  _zyL94_iscX1c0_s = 1'b0;
  _zyL94_iscX1c0_n = 1'b1;
  _zyL61_iscX2c0_s = 1'b0;
  _zyL61_iscX2c0_n = 1'b1;
 end
// F1, L10
initial 
 // F1, L10
 begin
  // F1, L324
  _zyM2L324_pbcCapEn0 = 1'b1;
  _zyM2L333_pbcCapEn1 = 1'b0;
  _zyM2L349_pbcCapEn2 = 1'b0;
  _zyM2L355_pbcCapEn3 = 1'b0;
  _zyM2L253_pbcCapEn5 = 1'b1;
  _zyM2L274_pbcCapEn6 = 1'b0;
  _zyM2L287_pbcCapEn7 = 1'b0;
  _zyM2L293_pbcCapEn8 = 1'b0;
  _zyM2L295_pbcCapEn9 = 1'b0;
  _zyM2L364_pbcCapEn10 = 1'b0;
  _zyM2L300_pbcCapEn11 = 1'b0;
  _zyM2L324_pbcFsm0_s = 3'b0;
  _zyM2L253_pbcFsm2_s = 3'b0;
  begin
  end
 end
endmodule

