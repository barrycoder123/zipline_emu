
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module cr_kme_key_tlv_compare_split ( set_key_tlv_miscmp_int, 
	cceip_encrypt_ob_full, cceip_encrypt_ob_afull, 
	cceip_validate_ob_full, cceip_validate_ob_afull, cceip_ob_wr, 
	.cceip_ob_tlv( {\cceip_ob_tlv[3].insert , 
	\cceip_ob_tlv[3].ordern[12] , \cceip_ob_tlv[3].ordern[11] , 
	\cceip_ob_tlv[3].ordern[10] , \cceip_ob_tlv[3].ordern[9] , 
	\cceip_ob_tlv[3].ordern[8] , \cceip_ob_tlv[3].ordern[7] , 
	\cceip_ob_tlv[3].ordern[6] , \cceip_ob_tlv[3].ordern[5] , 
	\cceip_ob_tlv[3].ordern[4] , \cceip_ob_tlv[3].ordern[3] , 
	\cceip_ob_tlv[3].ordern[2] , \cceip_ob_tlv[3].ordern[1] , 
	\cceip_ob_tlv[3].ordern[0] , \cceip_ob_tlv[3].typen[7] , 
	\cceip_ob_tlv[3].typen[6] , \cceip_ob_tlv[3].typen[5] , 
	\cceip_ob_tlv[3].typen[4] , \cceip_ob_tlv[3].typen[3] , 
	\cceip_ob_tlv[3].typen[2] , \cceip_ob_tlv[3].typen[1] , 
	\cceip_ob_tlv[3].typen[0] , \cceip_ob_tlv[3].sot , 
	\cceip_ob_tlv[3].eot , \cceip_ob_tlv[3].tlast , 
	\cceip_ob_tlv[3].tid[0] , \cceip_ob_tlv[3].tstrb[7] , 
	\cceip_ob_tlv[3].tstrb[6] , \cceip_ob_tlv[3].tstrb[5] , 
	\cceip_ob_tlv[3].tstrb[4] , \cceip_ob_tlv[3].tstrb[3] , 
	\cceip_ob_tlv[3].tstrb[2] , \cceip_ob_tlv[3].tstrb[1] , 
	\cceip_ob_tlv[3].tstrb[0] , \cceip_ob_tlv[3].tuser[7] , 
	\cceip_ob_tlv[3].tuser[6] , \cceip_ob_tlv[3].tuser[5] , 
	\cceip_ob_tlv[3].tuser[4] , \cceip_ob_tlv[3].tuser[3] , 
	\cceip_ob_tlv[3].tuser[2] , \cceip_ob_tlv[3].tuser[1] , 
	\cceip_ob_tlv[3].tuser[0] , \cceip_ob_tlv[3].tdata[63] , 
	\cceip_ob_tlv[3].tdata[62] , \cceip_ob_tlv[3].tdata[61] , 
	\cceip_ob_tlv[3].tdata[60] , \cceip_ob_tlv[3].tdata[59] , 
	\cceip_ob_tlv[3].tdata[58] , \cceip_ob_tlv[3].tdata[57] , 
	\cceip_ob_tlv[3].tdata[56] , \cceip_ob_tlv[3].tdata[55] , 
	\cceip_ob_tlv[3].tdata[54] , \cceip_ob_tlv[3].tdata[53] , 
	\cceip_ob_tlv[3].tdata[52] , \cceip_ob_tlv[3].tdata[51] , 
	\cceip_ob_tlv[3].tdata[50] , \cceip_ob_tlv[3].tdata[49] , 
	\cceip_ob_tlv[3].tdata[48] , \cceip_ob_tlv[3].tdata[47] , 
	\cceip_ob_tlv[3].tdata[46] , \cceip_ob_tlv[3].tdata[45] , 
	\cceip_ob_tlv[3].tdata[44] , \cceip_ob_tlv[3].tdata[43] , 
	\cceip_ob_tlv[3].tdata[42] , \cceip_ob_tlv[3].tdata[41] , 
	\cceip_ob_tlv[3].tdata[40] , \cceip_ob_tlv[3].tdata[39] , 
	\cceip_ob_tlv[3].tdata[38] , \cceip_ob_tlv[3].tdata[37] , 
	\cceip_ob_tlv[3].tdata[36] , \cceip_ob_tlv[3].tdata[35] , 
	\cceip_ob_tlv[3].tdata[34] , \cceip_ob_tlv[3].tdata[33] , 
	\cceip_ob_tlv[3].tdata[32] , \cceip_ob_tlv[3].tdata[31] , 
	\cceip_ob_tlv[3].tdata[30] , \cceip_ob_tlv[3].tdata[29] , 
	\cceip_ob_tlv[3].tdata[28] , \cceip_ob_tlv[3].tdata[27] , 
	\cceip_ob_tlv[3].tdata[26] , \cceip_ob_tlv[3].tdata[25] , 
	\cceip_ob_tlv[3].tdata[24] , \cceip_ob_tlv[3].tdata[23] , 
	\cceip_ob_tlv[3].tdata[22] , \cceip_ob_tlv[3].tdata[21] , 
	\cceip_ob_tlv[3].tdata[20] , \cceip_ob_tlv[3].tdata[19] , 
	\cceip_ob_tlv[3].tdata[18] , \cceip_ob_tlv[3].tdata[17] , 
	\cceip_ob_tlv[3].tdata[16] , \cceip_ob_tlv[3].tdata[15] , 
	\cceip_ob_tlv[3].tdata[14] , \cceip_ob_tlv[3].tdata[13] , 
	\cceip_ob_tlv[3].tdata[12] , \cceip_ob_tlv[3].tdata[11] , 
	\cceip_ob_tlv[3].tdata[10] , \cceip_ob_tlv[3].tdata[9] , 
	\cceip_ob_tlv[3].tdata[8] , \cceip_ob_tlv[3].tdata[7] , 
	\cceip_ob_tlv[3].tdata[6] , \cceip_ob_tlv[3].tdata[5] , 
	\cceip_ob_tlv[3].tdata[4] , \cceip_ob_tlv[3].tdata[3] , 
	\cceip_ob_tlv[3].tdata[2] , \cceip_ob_tlv[3].tdata[1] , 
	\cceip_ob_tlv[3].tdata[0] , \cceip_ob_tlv[2].insert , 
	\cceip_ob_tlv[2].ordern[12] , \cceip_ob_tlv[2].ordern[11] , 
	\cceip_ob_tlv[2].ordern[10] , \cceip_ob_tlv[2].ordern[9] , 
	\cceip_ob_tlv[2].ordern[8] , \cceip_ob_tlv[2].ordern[7] , 
	\cceip_ob_tlv[2].ordern[6] , \cceip_ob_tlv[2].ordern[5] , 
	\cceip_ob_tlv[2].ordern[4] , \cceip_ob_tlv[2].ordern[3] , 
	\cceip_ob_tlv[2].ordern[2] , \cceip_ob_tlv[2].ordern[1] , 
	\cceip_ob_tlv[2].ordern[0] , \cceip_ob_tlv[2].typen[7] , 
	\cceip_ob_tlv[2].typen[6] , \cceip_ob_tlv[2].typen[5] , 
	\cceip_ob_tlv[2].typen[4] , \cceip_ob_tlv[2].typen[3] , 
	\cceip_ob_tlv[2].typen[2] , \cceip_ob_tlv[2].typen[1] , 
	\cceip_ob_tlv[2].typen[0] , \cceip_ob_tlv[2].sot , 
	\cceip_ob_tlv[2].eot , \cceip_ob_tlv[2].tlast , 
	\cceip_ob_tlv[2].tid[0] , \cceip_ob_tlv[2].tstrb[7] , 
	\cceip_ob_tlv[2].tstrb[6] , \cceip_ob_tlv[2].tstrb[5] , 
	\cceip_ob_tlv[2].tstrb[4] , \cceip_ob_tlv[2].tstrb[3] , 
	\cceip_ob_tlv[2].tstrb[2] , \cceip_ob_tlv[2].tstrb[1] , 
	\cceip_ob_tlv[2].tstrb[0] , \cceip_ob_tlv[2].tuser[7] , 
	\cceip_ob_tlv[2].tuser[6] , \cceip_ob_tlv[2].tuser[5] , 
	\cceip_ob_tlv[2].tuser[4] , \cceip_ob_tlv[2].tuser[3] , 
	\cceip_ob_tlv[2].tuser[2] , \cceip_ob_tlv[2].tuser[1] , 
	\cceip_ob_tlv[2].tuser[0] , \cceip_ob_tlv[2].tdata[63] , 
	\cceip_ob_tlv[2].tdata[62] , \cceip_ob_tlv[2].tdata[61] , 
	\cceip_ob_tlv[2].tdata[60] , \cceip_ob_tlv[2].tdata[59] , 
	\cceip_ob_tlv[2].tdata[58] , \cceip_ob_tlv[2].tdata[57] , 
	\cceip_ob_tlv[2].tdata[56] , \cceip_ob_tlv[2].tdata[55] , 
	\cceip_ob_tlv[2].tdata[54] , \cceip_ob_tlv[2].tdata[53] , 
	\cceip_ob_tlv[2].tdata[52] , \cceip_ob_tlv[2].tdata[51] , 
	\cceip_ob_tlv[2].tdata[50] , \cceip_ob_tlv[2].tdata[49] , 
	\cceip_ob_tlv[2].tdata[48] , \cceip_ob_tlv[2].tdata[47] , 
	\cceip_ob_tlv[2].tdata[46] , \cceip_ob_tlv[2].tdata[45] , 
	\cceip_ob_tlv[2].tdata[44] , \cceip_ob_tlv[2].tdata[43] , 
	\cceip_ob_tlv[2].tdata[42] , \cceip_ob_tlv[2].tdata[41] , 
	\cceip_ob_tlv[2].tdata[40] , \cceip_ob_tlv[2].tdata[39] , 
	\cceip_ob_tlv[2].tdata[38] , \cceip_ob_tlv[2].tdata[37] , 
	\cceip_ob_tlv[2].tdata[36] , \cceip_ob_tlv[2].tdata[35] , 
	\cceip_ob_tlv[2].tdata[34] , \cceip_ob_tlv[2].tdata[33] , 
	\cceip_ob_tlv[2].tdata[32] , \cceip_ob_tlv[2].tdata[31] , 
	\cceip_ob_tlv[2].tdata[30] , \cceip_ob_tlv[2].tdata[29] , 
	\cceip_ob_tlv[2].tdata[28] , \cceip_ob_tlv[2].tdata[27] , 
	\cceip_ob_tlv[2].tdata[26] , \cceip_ob_tlv[2].tdata[25] , 
	\cceip_ob_tlv[2].tdata[24] , \cceip_ob_tlv[2].tdata[23] , 
	\cceip_ob_tlv[2].tdata[22] , \cceip_ob_tlv[2].tdata[21] , 
	\cceip_ob_tlv[2].tdata[20] , \cceip_ob_tlv[2].tdata[19] , 
	\cceip_ob_tlv[2].tdata[18] , \cceip_ob_tlv[2].tdata[17] , 
	\cceip_ob_tlv[2].tdata[16] , \cceip_ob_tlv[2].tdata[15] , 
	\cceip_ob_tlv[2].tdata[14] , \cceip_ob_tlv[2].tdata[13] , 
	\cceip_ob_tlv[2].tdata[12] , \cceip_ob_tlv[2].tdata[11] , 
	\cceip_ob_tlv[2].tdata[10] , \cceip_ob_tlv[2].tdata[9] , 
	\cceip_ob_tlv[2].tdata[8] , \cceip_ob_tlv[2].tdata[7] , 
	\cceip_ob_tlv[2].tdata[6] , \cceip_ob_tlv[2].tdata[5] , 
	\cceip_ob_tlv[2].tdata[4] , \cceip_ob_tlv[2].tdata[3] , 
	\cceip_ob_tlv[2].tdata[2] , \cceip_ob_tlv[2].tdata[1] , 
	\cceip_ob_tlv[2].tdata[0] , \cceip_ob_tlv[1].insert , 
	\cceip_ob_tlv[1].ordern[12] , \cceip_ob_tlv[1].ordern[11] , 
	\cceip_ob_tlv[1].ordern[10] , \cceip_ob_tlv[1].ordern[9] , 
	\cceip_ob_tlv[1].ordern[8] , \cceip_ob_tlv[1].ordern[7] , 
	\cceip_ob_tlv[1].ordern[6] , \cceip_ob_tlv[1].ordern[5] , 
	\cceip_ob_tlv[1].ordern[4] , \cceip_ob_tlv[1].ordern[3] , 
	\cceip_ob_tlv[1].ordern[2] , \cceip_ob_tlv[1].ordern[1] , 
	\cceip_ob_tlv[1].ordern[0] , \cceip_ob_tlv[1].typen[7] , 
	\cceip_ob_tlv[1].typen[6] , \cceip_ob_tlv[1].typen[5] , 
	\cceip_ob_tlv[1].typen[4] , \cceip_ob_tlv[1].typen[3] , 
	\cceip_ob_tlv[1].typen[2] , \cceip_ob_tlv[1].typen[1] , 
	\cceip_ob_tlv[1].typen[0] , \cceip_ob_tlv[1].sot , 
	\cceip_ob_tlv[1].eot , \cceip_ob_tlv[1].tlast , 
	\cceip_ob_tlv[1].tid[0] , \cceip_ob_tlv[1].tstrb[7] , 
	\cceip_ob_tlv[1].tstrb[6] , \cceip_ob_tlv[1].tstrb[5] , 
	\cceip_ob_tlv[1].tstrb[4] , \cceip_ob_tlv[1].tstrb[3] , 
	\cceip_ob_tlv[1].tstrb[2] , \cceip_ob_tlv[1].tstrb[1] , 
	\cceip_ob_tlv[1].tstrb[0] , \cceip_ob_tlv[1].tuser[7] , 
	\cceip_ob_tlv[1].tuser[6] , \cceip_ob_tlv[1].tuser[5] , 
	\cceip_ob_tlv[1].tuser[4] , \cceip_ob_tlv[1].tuser[3] , 
	\cceip_ob_tlv[1].tuser[2] , \cceip_ob_tlv[1].tuser[1] , 
	\cceip_ob_tlv[1].tuser[0] , \cceip_ob_tlv[1].tdata[63] , 
	\cceip_ob_tlv[1].tdata[62] , \cceip_ob_tlv[1].tdata[61] , 
	\cceip_ob_tlv[1].tdata[60] , \cceip_ob_tlv[1].tdata[59] , 
	\cceip_ob_tlv[1].tdata[58] , \cceip_ob_tlv[1].tdata[57] , 
	\cceip_ob_tlv[1].tdata[56] , \cceip_ob_tlv[1].tdata[55] , 
	\cceip_ob_tlv[1].tdata[54] , \cceip_ob_tlv[1].tdata[53] , 
	\cceip_ob_tlv[1].tdata[52] , \cceip_ob_tlv[1].tdata[51] , 
	\cceip_ob_tlv[1].tdata[50] , \cceip_ob_tlv[1].tdata[49] , 
	\cceip_ob_tlv[1].tdata[48] , \cceip_ob_tlv[1].tdata[47] , 
	\cceip_ob_tlv[1].tdata[46] , \cceip_ob_tlv[1].tdata[45] , 
	\cceip_ob_tlv[1].tdata[44] , \cceip_ob_tlv[1].tdata[43] , 
	\cceip_ob_tlv[1].tdata[42] , \cceip_ob_tlv[1].tdata[41] , 
	\cceip_ob_tlv[1].tdata[40] , \cceip_ob_tlv[1].tdata[39] , 
	\cceip_ob_tlv[1].tdata[38] , \cceip_ob_tlv[1].tdata[37] , 
	\cceip_ob_tlv[1].tdata[36] , \cceip_ob_tlv[1].tdata[35] , 
	\cceip_ob_tlv[1].tdata[34] , \cceip_ob_tlv[1].tdata[33] , 
	\cceip_ob_tlv[1].tdata[32] , \cceip_ob_tlv[1].tdata[31] , 
	\cceip_ob_tlv[1].tdata[30] , \cceip_ob_tlv[1].tdata[29] , 
	\cceip_ob_tlv[1].tdata[28] , \cceip_ob_tlv[1].tdata[27] , 
	\cceip_ob_tlv[1].tdata[26] , \cceip_ob_tlv[1].tdata[25] , 
	\cceip_ob_tlv[1].tdata[24] , \cceip_ob_tlv[1].tdata[23] , 
	\cceip_ob_tlv[1].tdata[22] , \cceip_ob_tlv[1].tdata[21] , 
	\cceip_ob_tlv[1].tdata[20] , \cceip_ob_tlv[1].tdata[19] , 
	\cceip_ob_tlv[1].tdata[18] , \cceip_ob_tlv[1].tdata[17] , 
	\cceip_ob_tlv[1].tdata[16] , \cceip_ob_tlv[1].tdata[15] , 
	\cceip_ob_tlv[1].tdata[14] , \cceip_ob_tlv[1].tdata[13] , 
	\cceip_ob_tlv[1].tdata[12] , \cceip_ob_tlv[1].tdata[11] , 
	\cceip_ob_tlv[1].tdata[10] , \cceip_ob_tlv[1].tdata[9] , 
	\cceip_ob_tlv[1].tdata[8] , \cceip_ob_tlv[1].tdata[7] , 
	\cceip_ob_tlv[1].tdata[6] , \cceip_ob_tlv[1].tdata[5] , 
	\cceip_ob_tlv[1].tdata[4] , \cceip_ob_tlv[1].tdata[3] , 
	\cceip_ob_tlv[1].tdata[2] , \cceip_ob_tlv[1].tdata[1] , 
	\cceip_ob_tlv[1].tdata[0] , \cceip_ob_tlv[0].insert , 
	\cceip_ob_tlv[0].ordern[12] , \cceip_ob_tlv[0].ordern[11] , 
	\cceip_ob_tlv[0].ordern[10] , \cceip_ob_tlv[0].ordern[9] , 
	\cceip_ob_tlv[0].ordern[8] , \cceip_ob_tlv[0].ordern[7] , 
	\cceip_ob_tlv[0].ordern[6] , \cceip_ob_tlv[0].ordern[5] , 
	\cceip_ob_tlv[0].ordern[4] , \cceip_ob_tlv[0].ordern[3] , 
	\cceip_ob_tlv[0].ordern[2] , \cceip_ob_tlv[0].ordern[1] , 
	\cceip_ob_tlv[0].ordern[0] , \cceip_ob_tlv[0].typen[7] , 
	\cceip_ob_tlv[0].typen[6] , \cceip_ob_tlv[0].typen[5] , 
	\cceip_ob_tlv[0].typen[4] , \cceip_ob_tlv[0].typen[3] , 
	\cceip_ob_tlv[0].typen[2] , \cceip_ob_tlv[0].typen[1] , 
	\cceip_ob_tlv[0].typen[0] , \cceip_ob_tlv[0].sot , 
	\cceip_ob_tlv[0].eot , \cceip_ob_tlv[0].tlast , 
	\cceip_ob_tlv[0].tid[0] , \cceip_ob_tlv[0].tstrb[7] , 
	\cceip_ob_tlv[0].tstrb[6] , \cceip_ob_tlv[0].tstrb[5] , 
	\cceip_ob_tlv[0].tstrb[4] , \cceip_ob_tlv[0].tstrb[3] , 
	\cceip_ob_tlv[0].tstrb[2] , \cceip_ob_tlv[0].tstrb[1] , 
	\cceip_ob_tlv[0].tstrb[0] , \cceip_ob_tlv[0].tuser[7] , 
	\cceip_ob_tlv[0].tuser[6] , \cceip_ob_tlv[0].tuser[5] , 
	\cceip_ob_tlv[0].tuser[4] , \cceip_ob_tlv[0].tuser[3] , 
	\cceip_ob_tlv[0].tuser[2] , \cceip_ob_tlv[0].tuser[1] , 
	\cceip_ob_tlv[0].tuser[0] , \cceip_ob_tlv[0].tdata[63] , 
	\cceip_ob_tlv[0].tdata[62] , \cceip_ob_tlv[0].tdata[61] , 
	\cceip_ob_tlv[0].tdata[60] , \cceip_ob_tlv[0].tdata[59] , 
	\cceip_ob_tlv[0].tdata[58] , \cceip_ob_tlv[0].tdata[57] , 
	\cceip_ob_tlv[0].tdata[56] , \cceip_ob_tlv[0].tdata[55] , 
	\cceip_ob_tlv[0].tdata[54] , \cceip_ob_tlv[0].tdata[53] , 
	\cceip_ob_tlv[0].tdata[52] , \cceip_ob_tlv[0].tdata[51] , 
	\cceip_ob_tlv[0].tdata[50] , \cceip_ob_tlv[0].tdata[49] , 
	\cceip_ob_tlv[0].tdata[48] , \cceip_ob_tlv[0].tdata[47] , 
	\cceip_ob_tlv[0].tdata[46] , \cceip_ob_tlv[0].tdata[45] , 
	\cceip_ob_tlv[0].tdata[44] , \cceip_ob_tlv[0].tdata[43] , 
	\cceip_ob_tlv[0].tdata[42] , \cceip_ob_tlv[0].tdata[41] , 
	\cceip_ob_tlv[0].tdata[40] , \cceip_ob_tlv[0].tdata[39] , 
	\cceip_ob_tlv[0].tdata[38] , \cceip_ob_tlv[0].tdata[37] , 
	\cceip_ob_tlv[0].tdata[36] , \cceip_ob_tlv[0].tdata[35] , 
	\cceip_ob_tlv[0].tdata[34] , \cceip_ob_tlv[0].tdata[33] , 
	\cceip_ob_tlv[0].tdata[32] , \cceip_ob_tlv[0].tdata[31] , 
	\cceip_ob_tlv[0].tdata[30] , \cceip_ob_tlv[0].tdata[29] , 
	\cceip_ob_tlv[0].tdata[28] , \cceip_ob_tlv[0].tdata[27] , 
	\cceip_ob_tlv[0].tdata[26] , \cceip_ob_tlv[0].tdata[25] , 
	\cceip_ob_tlv[0].tdata[24] , \cceip_ob_tlv[0].tdata[23] , 
	\cceip_ob_tlv[0].tdata[22] , \cceip_ob_tlv[0].tdata[21] , 
	\cceip_ob_tlv[0].tdata[20] , \cceip_ob_tlv[0].tdata[19] , 
	\cceip_ob_tlv[0].tdata[18] , \cceip_ob_tlv[0].tdata[17] , 
	\cceip_ob_tlv[0].tdata[16] , \cceip_ob_tlv[0].tdata[15] , 
	\cceip_ob_tlv[0].tdata[14] , \cceip_ob_tlv[0].tdata[13] , 
	\cceip_ob_tlv[0].tdata[12] , \cceip_ob_tlv[0].tdata[11] , 
	\cceip_ob_tlv[0].tdata[10] , \cceip_ob_tlv[0].tdata[9] , 
	\cceip_ob_tlv[0].tdata[8] , \cceip_ob_tlv[0].tdata[7] , 
	\cceip_ob_tlv[0].tdata[6] , \cceip_ob_tlv[0].tdata[5] , 
	\cceip_ob_tlv[0].tdata[4] , \cceip_ob_tlv[0].tdata[3] , 
	\cceip_ob_tlv[0].tdata[2] , \cceip_ob_tlv[0].tdata[1] , 
	\cceip_ob_tlv[0].tdata[0] } ), clk, rst_n, suppress_key_tlvs, 
	cceip_encrypt_ob_wr, .cceip_encrypt_ob_tlv( {
	\cceip_encrypt_ob_tlv.insert , \cceip_encrypt_ob_tlv.ordern [12], 
	\cceip_encrypt_ob_tlv.ordern [11], \cceip_encrypt_ob_tlv.ordern [10], 
	\cceip_encrypt_ob_tlv.ordern [9], \cceip_encrypt_ob_tlv.ordern [8], 
	\cceip_encrypt_ob_tlv.ordern [7], \cceip_encrypt_ob_tlv.ordern [6], 
	\cceip_encrypt_ob_tlv.ordern [5], \cceip_encrypt_ob_tlv.ordern [4], 
	\cceip_encrypt_ob_tlv.ordern [3], \cceip_encrypt_ob_tlv.ordern [2], 
	\cceip_encrypt_ob_tlv.ordern [1], \cceip_encrypt_ob_tlv.ordern [0], 
	\cceip_encrypt_ob_tlv.typen [7], \cceip_encrypt_ob_tlv.typen [6], 
	\cceip_encrypt_ob_tlv.typen [5], \cceip_encrypt_ob_tlv.typen [4], 
	\cceip_encrypt_ob_tlv.typen [3], \cceip_encrypt_ob_tlv.typen [2], 
	\cceip_encrypt_ob_tlv.typen [1], \cceip_encrypt_ob_tlv.typen [0], 
	\cceip_encrypt_ob_tlv.sot , \cceip_encrypt_ob_tlv.eot , 
	\cceip_encrypt_ob_tlv.tlast , \cceip_encrypt_ob_tlv.tid [0], 
	\cceip_encrypt_ob_tlv.tstrb [7], \cceip_encrypt_ob_tlv.tstrb [6], 
	\cceip_encrypt_ob_tlv.tstrb [5], \cceip_encrypt_ob_tlv.tstrb [4], 
	\cceip_encrypt_ob_tlv.tstrb [3], \cceip_encrypt_ob_tlv.tstrb [2], 
	\cceip_encrypt_ob_tlv.tstrb [1], \cceip_encrypt_ob_tlv.tstrb [0], 
	\cceip_encrypt_ob_tlv.tuser [7], \cceip_encrypt_ob_tlv.tuser [6], 
	\cceip_encrypt_ob_tlv.tuser [5], \cceip_encrypt_ob_tlv.tuser [4], 
	\cceip_encrypt_ob_tlv.tuser [3], \cceip_encrypt_ob_tlv.tuser [2], 
	\cceip_encrypt_ob_tlv.tuser [1], \cceip_encrypt_ob_tlv.tuser [0], 
	\cceip_encrypt_ob_tlv.tdata [63], \cceip_encrypt_ob_tlv.tdata [62], 
	\cceip_encrypt_ob_tlv.tdata [61], \cceip_encrypt_ob_tlv.tdata [60], 
	\cceip_encrypt_ob_tlv.tdata [59], \cceip_encrypt_ob_tlv.tdata [58], 
	\cceip_encrypt_ob_tlv.tdata [57], \cceip_encrypt_ob_tlv.tdata [56], 
	\cceip_encrypt_ob_tlv.tdata [55], \cceip_encrypt_ob_tlv.tdata [54], 
	\cceip_encrypt_ob_tlv.tdata [53], \cceip_encrypt_ob_tlv.tdata [52], 
	\cceip_encrypt_ob_tlv.tdata [51], \cceip_encrypt_ob_tlv.tdata [50], 
	\cceip_encrypt_ob_tlv.tdata [49], \cceip_encrypt_ob_tlv.tdata [48], 
	\cceip_encrypt_ob_tlv.tdata [47], \cceip_encrypt_ob_tlv.tdata [46], 
	\cceip_encrypt_ob_tlv.tdata [45], \cceip_encrypt_ob_tlv.tdata [44], 
	\cceip_encrypt_ob_tlv.tdata [43], \cceip_encrypt_ob_tlv.tdata [42], 
	\cceip_encrypt_ob_tlv.tdata [41], \cceip_encrypt_ob_tlv.tdata [40], 
	\cceip_encrypt_ob_tlv.tdata [39], \cceip_encrypt_ob_tlv.tdata [38], 
	\cceip_encrypt_ob_tlv.tdata [37], \cceip_encrypt_ob_tlv.tdata [36], 
	\cceip_encrypt_ob_tlv.tdata [35], \cceip_encrypt_ob_tlv.tdata [34], 
	\cceip_encrypt_ob_tlv.tdata [33], \cceip_encrypt_ob_tlv.tdata [32], 
	\cceip_encrypt_ob_tlv.tdata [31], \cceip_encrypt_ob_tlv.tdata [30], 
	\cceip_encrypt_ob_tlv.tdata [29], \cceip_encrypt_ob_tlv.tdata [28], 
	\cceip_encrypt_ob_tlv.tdata [27], \cceip_encrypt_ob_tlv.tdata [26], 
	\cceip_encrypt_ob_tlv.tdata [25], \cceip_encrypt_ob_tlv.tdata [24], 
	\cceip_encrypt_ob_tlv.tdata [23], \cceip_encrypt_ob_tlv.tdata [22], 
	\cceip_encrypt_ob_tlv.tdata [21], \cceip_encrypt_ob_tlv.tdata [20], 
	\cceip_encrypt_ob_tlv.tdata [19], \cceip_encrypt_ob_tlv.tdata [18], 
	\cceip_encrypt_ob_tlv.tdata [17], \cceip_encrypt_ob_tlv.tdata [16], 
	\cceip_encrypt_ob_tlv.tdata [15], \cceip_encrypt_ob_tlv.tdata [14], 
	\cceip_encrypt_ob_tlv.tdata [13], \cceip_encrypt_ob_tlv.tdata [12], 
	\cceip_encrypt_ob_tlv.tdata [11], \cceip_encrypt_ob_tlv.tdata [10], 
	\cceip_encrypt_ob_tlv.tdata [9], \cceip_encrypt_ob_tlv.tdata [8], 
	\cceip_encrypt_ob_tlv.tdata [7], \cceip_encrypt_ob_tlv.tdata [6], 
	\cceip_encrypt_ob_tlv.tdata [5], \cceip_encrypt_ob_tlv.tdata [4], 
	\cceip_encrypt_ob_tlv.tdata [3], \cceip_encrypt_ob_tlv.tdata [2], 
	\cceip_encrypt_ob_tlv.tdata [1], \cceip_encrypt_ob_tlv.tdata [0]} ), 
	cceip_validate_ob_wr, .cceip_validate_ob_tlv( {
	\cceip_validate_ob_tlv.insert , \cceip_validate_ob_tlv.ordern [12], 
	\cceip_validate_ob_tlv.ordern [11], 
	\cceip_validate_ob_tlv.ordern [10], 
	\cceip_validate_ob_tlv.ordern [9], \cceip_validate_ob_tlv.ordern [8], 
	\cceip_validate_ob_tlv.ordern [7], \cceip_validate_ob_tlv.ordern [6], 
	\cceip_validate_ob_tlv.ordern [5], \cceip_validate_ob_tlv.ordern [4], 
	\cceip_validate_ob_tlv.ordern [3], \cceip_validate_ob_tlv.ordern [2], 
	\cceip_validate_ob_tlv.ordern [1], \cceip_validate_ob_tlv.ordern [0], 
	\cceip_validate_ob_tlv.typen [7], \cceip_validate_ob_tlv.typen [6], 
	\cceip_validate_ob_tlv.typen [5], \cceip_validate_ob_tlv.typen [4], 
	\cceip_validate_ob_tlv.typen [3], \cceip_validate_ob_tlv.typen [2], 
	\cceip_validate_ob_tlv.typen [1], \cceip_validate_ob_tlv.typen [0], 
	\cceip_validate_ob_tlv.sot , \cceip_validate_ob_tlv.eot , 
	\cceip_validate_ob_tlv.tlast , \cceip_validate_ob_tlv.tid [0], 
	\cceip_validate_ob_tlv.tstrb [7], \cceip_validate_ob_tlv.tstrb [6], 
	\cceip_validate_ob_tlv.tstrb [5], \cceip_validate_ob_tlv.tstrb [4], 
	\cceip_validate_ob_tlv.tstrb [3], \cceip_validate_ob_tlv.tstrb [2], 
	\cceip_validate_ob_tlv.tstrb [1], \cceip_validate_ob_tlv.tstrb [0], 
	\cceip_validate_ob_tlv.tuser [7], \cceip_validate_ob_tlv.tuser [6], 
	\cceip_validate_ob_tlv.tuser [5], \cceip_validate_ob_tlv.tuser [4], 
	\cceip_validate_ob_tlv.tuser [3], \cceip_validate_ob_tlv.tuser [2], 
	\cceip_validate_ob_tlv.tuser [1], \cceip_validate_ob_tlv.tuser [0], 
	\cceip_validate_ob_tlv.tdata [63], \cceip_validate_ob_tlv.tdata [62], 
	\cceip_validate_ob_tlv.tdata [61], \cceip_validate_ob_tlv.tdata [60], 
	\cceip_validate_ob_tlv.tdata [59], \cceip_validate_ob_tlv.tdata [58], 
	\cceip_validate_ob_tlv.tdata [57], \cceip_validate_ob_tlv.tdata [56], 
	\cceip_validate_ob_tlv.tdata [55], \cceip_validate_ob_tlv.tdata [54], 
	\cceip_validate_ob_tlv.tdata [53], \cceip_validate_ob_tlv.tdata [52], 
	\cceip_validate_ob_tlv.tdata [51], \cceip_validate_ob_tlv.tdata [50], 
	\cceip_validate_ob_tlv.tdata [49], \cceip_validate_ob_tlv.tdata [48], 
	\cceip_validate_ob_tlv.tdata [47], \cceip_validate_ob_tlv.tdata [46], 
	\cceip_validate_ob_tlv.tdata [45], \cceip_validate_ob_tlv.tdata [44], 
	\cceip_validate_ob_tlv.tdata [43], \cceip_validate_ob_tlv.tdata [42], 
	\cceip_validate_ob_tlv.tdata [41], \cceip_validate_ob_tlv.tdata [40], 
	\cceip_validate_ob_tlv.tdata [39], \cceip_validate_ob_tlv.tdata [38], 
	\cceip_validate_ob_tlv.tdata [37], \cceip_validate_ob_tlv.tdata [36], 
	\cceip_validate_ob_tlv.tdata [35], \cceip_validate_ob_tlv.tdata [34], 
	\cceip_validate_ob_tlv.tdata [33], \cceip_validate_ob_tlv.tdata [32], 
	\cceip_validate_ob_tlv.tdata [31], \cceip_validate_ob_tlv.tdata [30], 
	\cceip_validate_ob_tlv.tdata [29], \cceip_validate_ob_tlv.tdata [28], 
	\cceip_validate_ob_tlv.tdata [27], \cceip_validate_ob_tlv.tdata [26], 
	\cceip_validate_ob_tlv.tdata [25], \cceip_validate_ob_tlv.tdata [24], 
	\cceip_validate_ob_tlv.tdata [23], \cceip_validate_ob_tlv.tdata [22], 
	\cceip_validate_ob_tlv.tdata [21], \cceip_validate_ob_tlv.tdata [20], 
	\cceip_validate_ob_tlv.tdata [19], \cceip_validate_ob_tlv.tdata [18], 
	\cceip_validate_ob_tlv.tdata [17], \cceip_validate_ob_tlv.tdata [16], 
	\cceip_validate_ob_tlv.tdata [15], \cceip_validate_ob_tlv.tdata [14], 
	\cceip_validate_ob_tlv.tdata [13], \cceip_validate_ob_tlv.tdata [12], 
	\cceip_validate_ob_tlv.tdata [11], \cceip_validate_ob_tlv.tdata [10], 
	\cceip_validate_ob_tlv.tdata [9], \cceip_validate_ob_tlv.tdata [8], 
	\cceip_validate_ob_tlv.tdata [7], \cceip_validate_ob_tlv.tdata [6], 
	\cceip_validate_ob_tlv.tdata [5], \cceip_validate_ob_tlv.tdata [4], 
	\cceip_validate_ob_tlv.tdata [3], \cceip_validate_ob_tlv.tdata [2], 
	\cceip_validate_ob_tlv.tdata [1], \cceip_validate_ob_tlv.tdata [0]} ), 
	cceip_ob_full, cceip_ob_afull);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output set_key_tlv_miscmp_int;
output cceip_encrypt_ob_full;
output cceip_encrypt_ob_afull;
output cceip_validate_ob_full;
output cceip_validate_ob_afull;
output [3:0] cceip_ob_wr;
output \cceip_ob_tlv[3].insert ,\cceip_ob_tlv[3].ordern[12] 
	,\cceip_ob_tlv[3].ordern[11] ,\cceip_ob_tlv[3].ordern[10] 
	,\cceip_ob_tlv[3].ordern[9] ,\cceip_ob_tlv[3].ordern[8] 
	,\cceip_ob_tlv[3].ordern[7] ,\cceip_ob_tlv[3].ordern[6] 
	,\cceip_ob_tlv[3].ordern[5] ,\cceip_ob_tlv[3].ordern[4] 
	,\cceip_ob_tlv[3].ordern[3] ,\cceip_ob_tlv[3].ordern[2] 
	,\cceip_ob_tlv[3].ordern[1] ,\cceip_ob_tlv[3].ordern[0] 
	,\cceip_ob_tlv[3].typen[7] ,\cceip_ob_tlv[3].typen[6] 
	,\cceip_ob_tlv[3].typen[5] ,\cceip_ob_tlv[3].typen[4] 
	,\cceip_ob_tlv[3].typen[3] ,\cceip_ob_tlv[3].typen[2] 
	,\cceip_ob_tlv[3].typen[1] ,\cceip_ob_tlv[3].typen[0] 
	,\cceip_ob_tlv[3].sot ,\cceip_ob_tlv[3].eot ,\cceip_ob_tlv[3].tlast 
	,\cceip_ob_tlv[3].tid[0] ,\cceip_ob_tlv[3].tstrb[7] 
	,\cceip_ob_tlv[3].tstrb[6] ,\cceip_ob_tlv[3].tstrb[5] 
	,\cceip_ob_tlv[3].tstrb[4] ,\cceip_ob_tlv[3].tstrb[3] 
	,\cceip_ob_tlv[3].tstrb[2] ,\cceip_ob_tlv[3].tstrb[1] 
	,\cceip_ob_tlv[3].tstrb[0] ,\cceip_ob_tlv[3].tuser[7] 
	,\cceip_ob_tlv[3].tuser[6] ,\cceip_ob_tlv[3].tuser[5] 
	,\cceip_ob_tlv[3].tuser[4] ,\cceip_ob_tlv[3].tuser[3] 
	,\cceip_ob_tlv[3].tuser[2] ,\cceip_ob_tlv[3].tuser[1] 
	,\cceip_ob_tlv[3].tuser[0] ,\cceip_ob_tlv[3].tdata[63] 
	,\cceip_ob_tlv[3].tdata[62] ,\cceip_ob_tlv[3].tdata[61] 
	,\cceip_ob_tlv[3].tdata[60] ,\cceip_ob_tlv[3].tdata[59] 
	,\cceip_ob_tlv[3].tdata[58] ,\cceip_ob_tlv[3].tdata[57] 
	,\cceip_ob_tlv[3].tdata[56] ,\cceip_ob_tlv[3].tdata[55] 
	,\cceip_ob_tlv[3].tdata[54] ,\cceip_ob_tlv[3].tdata[53] 
	,\cceip_ob_tlv[3].tdata[52] ,\cceip_ob_tlv[3].tdata[51] 
	,\cceip_ob_tlv[3].tdata[50] ,\cceip_ob_tlv[3].tdata[49] 
	,\cceip_ob_tlv[3].tdata[48] ,\cceip_ob_tlv[3].tdata[47] 
	,\cceip_ob_tlv[3].tdata[46] ,\cceip_ob_tlv[3].tdata[45] 
	,\cceip_ob_tlv[3].tdata[44] ,\cceip_ob_tlv[3].tdata[43] 
	,\cceip_ob_tlv[3].tdata[42] ,\cceip_ob_tlv[3].tdata[41] 
	,\cceip_ob_tlv[3].tdata[40] ,\cceip_ob_tlv[3].tdata[39] 
	,\cceip_ob_tlv[3].tdata[38] ,\cceip_ob_tlv[3].tdata[37] 
	,\cceip_ob_tlv[3].tdata[36] ,\cceip_ob_tlv[3].tdata[35] 
	,\cceip_ob_tlv[3].tdata[34] ,\cceip_ob_tlv[3].tdata[33] 
	,\cceip_ob_tlv[3].tdata[32] ,\cceip_ob_tlv[3].tdata[31] 
	,\cceip_ob_tlv[3].tdata[30] ,\cceip_ob_tlv[3].tdata[29] 
	,\cceip_ob_tlv[3].tdata[28] ,\cceip_ob_tlv[3].tdata[27] 
	,\cceip_ob_tlv[3].tdata[26] ,\cceip_ob_tlv[3].tdata[25] 
	,\cceip_ob_tlv[3].tdata[24] ,\cceip_ob_tlv[3].tdata[23] 
	,\cceip_ob_tlv[3].tdata[22] ,\cceip_ob_tlv[3].tdata[21] 
	,\cceip_ob_tlv[3].tdata[20] ,\cceip_ob_tlv[3].tdata[19] 
	,\cceip_ob_tlv[3].tdata[18] ,\cceip_ob_tlv[3].tdata[17] 
	,\cceip_ob_tlv[3].tdata[16] ,\cceip_ob_tlv[3].tdata[15] 
	,\cceip_ob_tlv[3].tdata[14] ,\cceip_ob_tlv[3].tdata[13] 
	,\cceip_ob_tlv[3].tdata[12] ,\cceip_ob_tlv[3].tdata[11] 
	,\cceip_ob_tlv[3].tdata[10] ,\cceip_ob_tlv[3].tdata[9] 
	,\cceip_ob_tlv[3].tdata[8] ,\cceip_ob_tlv[3].tdata[7] 
	,\cceip_ob_tlv[3].tdata[6] ,\cceip_ob_tlv[3].tdata[5] 
	,\cceip_ob_tlv[3].tdata[4] ,\cceip_ob_tlv[3].tdata[3] 
	,\cceip_ob_tlv[3].tdata[2] ,\cceip_ob_tlv[3].tdata[1] 
	,\cceip_ob_tlv[3].tdata[0] ,\cceip_ob_tlv[2].insert 
	,\cceip_ob_tlv[2].ordern[12] ,\cceip_ob_tlv[2].ordern[11] 
	,\cceip_ob_tlv[2].ordern[10] ,\cceip_ob_tlv[2].ordern[9] 
	,\cceip_ob_tlv[2].ordern[8] ,\cceip_ob_tlv[2].ordern[7] 
	,\cceip_ob_tlv[2].ordern[6] ,\cceip_ob_tlv[2].ordern[5] 
	,\cceip_ob_tlv[2].ordern[4] ,\cceip_ob_tlv[2].ordern[3] 
	,\cceip_ob_tlv[2].ordern[2] ,\cceip_ob_tlv[2].ordern[1] 
	,\cceip_ob_tlv[2].ordern[0] ,\cceip_ob_tlv[2].typen[7] 
	,\cceip_ob_tlv[2].typen[6] ,\cceip_ob_tlv[2].typen[5] 
	,\cceip_ob_tlv[2].typen[4] ,\cceip_ob_tlv[2].typen[3] 
	,\cceip_ob_tlv[2].typen[2] ,\cceip_ob_tlv[2].typen[1] 
	,\cceip_ob_tlv[2].typen[0] ,\cceip_ob_tlv[2].sot 
	,\cceip_ob_tlv[2].eot ,\cceip_ob_tlv[2].tlast 
	,\cceip_ob_tlv[2].tid[0] ,\cceip_ob_tlv[2].tstrb[7] 
	,\cceip_ob_tlv[2].tstrb[6] ,\cceip_ob_tlv[2].tstrb[5] 
	,\cceip_ob_tlv[2].tstrb[4] ,\cceip_ob_tlv[2].tstrb[3] 
	,\cceip_ob_tlv[2].tstrb[2] ,\cceip_ob_tlv[2].tstrb[1] 
	,\cceip_ob_tlv[2].tstrb[0] ,\cceip_ob_tlv[2].tuser[7] 
	,\cceip_ob_tlv[2].tuser[6] ,\cceip_ob_tlv[2].tuser[5] 
	,\cceip_ob_tlv[2].tuser[4] ,\cceip_ob_tlv[2].tuser[3] 
	,\cceip_ob_tlv[2].tuser[2] ,\cceip_ob_tlv[2].tuser[1] 
	,\cceip_ob_tlv[2].tuser[0] ,\cceip_ob_tlv[2].tdata[63] 
	,\cceip_ob_tlv[2].tdata[62] ,\cceip_ob_tlv[2].tdata[61] 
	,\cceip_ob_tlv[2].tdata[60] ,\cceip_ob_tlv[2].tdata[59] 
	,\cceip_ob_tlv[2].tdata[58] ,\cceip_ob_tlv[2].tdata[57] 
	,\cceip_ob_tlv[2].tdata[56] ,\cceip_ob_tlv[2].tdata[55] 
	,\cceip_ob_tlv[2].tdata[54] ,\cceip_ob_tlv[2].tdata[53] 
	,\cceip_ob_tlv[2].tdata[52] ,\cceip_ob_tlv[2].tdata[51] 
	,\cceip_ob_tlv[2].tdata[50] ,\cceip_ob_tlv[2].tdata[49] 
	,\cceip_ob_tlv[2].tdata[48] ,\cceip_ob_tlv[2].tdata[47] 
	,\cceip_ob_tlv[2].tdata[46] ,\cceip_ob_tlv[2].tdata[45] 
	,\cceip_ob_tlv[2].tdata[44] ,\cceip_ob_tlv[2].tdata[43] 
	,\cceip_ob_tlv[2].tdata[42] ,\cceip_ob_tlv[2].tdata[41] 
	,\cceip_ob_tlv[2].tdata[40] ,\cceip_ob_tlv[2].tdata[39] 
	,\cceip_ob_tlv[2].tdata[38] ,\cceip_ob_tlv[2].tdata[37] 
	,\cceip_ob_tlv[2].tdata[36] ,\cceip_ob_tlv[2].tdata[35] 
	,\cceip_ob_tlv[2].tdata[34] ,\cceip_ob_tlv[2].tdata[33] 
	,\cceip_ob_tlv[2].tdata[32] ,\cceip_ob_tlv[2].tdata[31] 
	,\cceip_ob_tlv[2].tdata[30] ,\cceip_ob_tlv[2].tdata[29] 
	,\cceip_ob_tlv[2].tdata[28] ,\cceip_ob_tlv[2].tdata[27] 
	,\cceip_ob_tlv[2].tdata[26] ,\cceip_ob_tlv[2].tdata[25] 
	,\cceip_ob_tlv[2].tdata[24] ,\cceip_ob_tlv[2].tdata[23] 
	,\cceip_ob_tlv[2].tdata[22] ,\cceip_ob_tlv[2].tdata[21] 
	,\cceip_ob_tlv[2].tdata[20] ,\cceip_ob_tlv[2].tdata[19] 
	,\cceip_ob_tlv[2].tdata[18] ,\cceip_ob_tlv[2].tdata[17] 
	,\cceip_ob_tlv[2].tdata[16] ,\cceip_ob_tlv[2].tdata[15] 
	,\cceip_ob_tlv[2].tdata[14] ,\cceip_ob_tlv[2].tdata[13] 
	,\cceip_ob_tlv[2].tdata[12] ,\cceip_ob_tlv[2].tdata[11] 
	,\cceip_ob_tlv[2].tdata[10] ,\cceip_ob_tlv[2].tdata[9] 
	,\cceip_ob_tlv[2].tdata[8] ,\cceip_ob_tlv[2].tdata[7] 
	,\cceip_ob_tlv[2].tdata[6] ,\cceip_ob_tlv[2].tdata[5] 
	,\cceip_ob_tlv[2].tdata[4] ,\cceip_ob_tlv[2].tdata[3] 
	,\cceip_ob_tlv[2].tdata[2] ,\cceip_ob_tlv[2].tdata[1] 
	,\cceip_ob_tlv[2].tdata[0] ,\cceip_ob_tlv[1].insert 
	,\cceip_ob_tlv[1].ordern[12] ,\cceip_ob_tlv[1].ordern[11] 
	,\cceip_ob_tlv[1].ordern[10] ,\cceip_ob_tlv[1].ordern[9] 
	,\cceip_ob_tlv[1].ordern[8] ,\cceip_ob_tlv[1].ordern[7] 
	,\cceip_ob_tlv[1].ordern[6] ,\cceip_ob_tlv[1].ordern[5] 
	,\cceip_ob_tlv[1].ordern[4] ,\cceip_ob_tlv[1].ordern[3] 
	,\cceip_ob_tlv[1].ordern[2] ,\cceip_ob_tlv[1].ordern[1] 
	,\cceip_ob_tlv[1].ordern[0] ,\cceip_ob_tlv[1].typen[7] 
	,\cceip_ob_tlv[1].typen[6] ,\cceip_ob_tlv[1].typen[5] 
	,\cceip_ob_tlv[1].typen[4] ,\cceip_ob_tlv[1].typen[3] 
	,\cceip_ob_tlv[1].typen[2] ,\cceip_ob_tlv[1].typen[1] 
	,\cceip_ob_tlv[1].typen[0] ,\cceip_ob_tlv[1].sot 
	,\cceip_ob_tlv[1].eot ,\cceip_ob_tlv[1].tlast 
	,\cceip_ob_tlv[1].tid[0] ,\cceip_ob_tlv[1].tstrb[7] 
	,\cceip_ob_tlv[1].tstrb[6] ,\cceip_ob_tlv[1].tstrb[5] 
	,\cceip_ob_tlv[1].tstrb[4] ,\cceip_ob_tlv[1].tstrb[3] 
	,\cceip_ob_tlv[1].tstrb[2] ,\cceip_ob_tlv[1].tstrb[1] 
	,\cceip_ob_tlv[1].tstrb[0] ,\cceip_ob_tlv[1].tuser[7] 
	,\cceip_ob_tlv[1].tuser[6] ,\cceip_ob_tlv[1].tuser[5] 
	,\cceip_ob_tlv[1].tuser[4] ,\cceip_ob_tlv[1].tuser[3] 
	,\cceip_ob_tlv[1].tuser[2] ,\cceip_ob_tlv[1].tuser[1] 
	,\cceip_ob_tlv[1].tuser[0] ,\cceip_ob_tlv[1].tdata[63] 
	,\cceip_ob_tlv[1].tdata[62] ,\cceip_ob_tlv[1].tdata[61] 
	,\cceip_ob_tlv[1].tdata[60] ,\cceip_ob_tlv[1].tdata[59] 
	,\cceip_ob_tlv[1].tdata[58] ,\cceip_ob_tlv[1].tdata[57] 
	,\cceip_ob_tlv[1].tdata[56] ,\cceip_ob_tlv[1].tdata[55] 
	,\cceip_ob_tlv[1].tdata[54] ,\cceip_ob_tlv[1].tdata[53] 
	,\cceip_ob_tlv[1].tdata[52] ,\cceip_ob_tlv[1].tdata[51] 
	,\cceip_ob_tlv[1].tdata[50] ,\cceip_ob_tlv[1].tdata[49] 
	,\cceip_ob_tlv[1].tdata[48] ,\cceip_ob_tlv[1].tdata[47] 
	,\cceip_ob_tlv[1].tdata[46] ,\cceip_ob_tlv[1].tdata[45] 
	,\cceip_ob_tlv[1].tdata[44] ,\cceip_ob_tlv[1].tdata[43] 
	,\cceip_ob_tlv[1].tdata[42] ,\cceip_ob_tlv[1].tdata[41] 
	,\cceip_ob_tlv[1].tdata[40] ,\cceip_ob_tlv[1].tdata[39] 
	,\cceip_ob_tlv[1].tdata[38] ,\cceip_ob_tlv[1].tdata[37] 
	,\cceip_ob_tlv[1].tdata[36] ,\cceip_ob_tlv[1].tdata[35] 
	,\cceip_ob_tlv[1].tdata[34] ,\cceip_ob_tlv[1].tdata[33] 
	,\cceip_ob_tlv[1].tdata[32] ,\cceip_ob_tlv[1].tdata[31] 
	,\cceip_ob_tlv[1].tdata[30] ,\cceip_ob_tlv[1].tdata[29] 
	,\cceip_ob_tlv[1].tdata[28] ,\cceip_ob_tlv[1].tdata[27] 
	,\cceip_ob_tlv[1].tdata[26] ,\cceip_ob_tlv[1].tdata[25] 
	,\cceip_ob_tlv[1].tdata[24] ,\cceip_ob_tlv[1].tdata[23] 
	,\cceip_ob_tlv[1].tdata[22] ,\cceip_ob_tlv[1].tdata[21] 
	,\cceip_ob_tlv[1].tdata[20] ,\cceip_ob_tlv[1].tdata[19] 
	,\cceip_ob_tlv[1].tdata[18] ,\cceip_ob_tlv[1].tdata[17] 
	,\cceip_ob_tlv[1].tdata[16] ,\cceip_ob_tlv[1].tdata[15] 
	,\cceip_ob_tlv[1].tdata[14] ,\cceip_ob_tlv[1].tdata[13] 
	,\cceip_ob_tlv[1].tdata[12] ,\cceip_ob_tlv[1].tdata[11] 
	,\cceip_ob_tlv[1].tdata[10] ,\cceip_ob_tlv[1].tdata[9] 
	,\cceip_ob_tlv[1].tdata[8] ,\cceip_ob_tlv[1].tdata[7] 
	,\cceip_ob_tlv[1].tdata[6] ,\cceip_ob_tlv[1].tdata[5] 
	,\cceip_ob_tlv[1].tdata[4] ,\cceip_ob_tlv[1].tdata[3] 
	,\cceip_ob_tlv[1].tdata[2] ,\cceip_ob_tlv[1].tdata[1] 
	,\cceip_ob_tlv[1].tdata[0] ,\cceip_ob_tlv[0].insert 
	,\cceip_ob_tlv[0].ordern[12] ,\cceip_ob_tlv[0].ordern[11] 
	,\cceip_ob_tlv[0].ordern[10] ,\cceip_ob_tlv[0].ordern[9] 
	,\cceip_ob_tlv[0].ordern[8] ,\cceip_ob_tlv[0].ordern[7] 
	,\cceip_ob_tlv[0].ordern[6] ,\cceip_ob_tlv[0].ordern[5] 
	,\cceip_ob_tlv[0].ordern[4] ,\cceip_ob_tlv[0].ordern[3] 
	,\cceip_ob_tlv[0].ordern[2] ,\cceip_ob_tlv[0].ordern[1] 
	,\cceip_ob_tlv[0].ordern[0] ,\cceip_ob_tlv[0].typen[7] 
	,\cceip_ob_tlv[0].typen[6] ,\cceip_ob_tlv[0].typen[5] 
	,\cceip_ob_tlv[0].typen[4] ,\cceip_ob_tlv[0].typen[3] 
	,\cceip_ob_tlv[0].typen[2] ,\cceip_ob_tlv[0].typen[1] 
	,\cceip_ob_tlv[0].typen[0] ,\cceip_ob_tlv[0].sot 
	,\cceip_ob_tlv[0].eot ,\cceip_ob_tlv[0].tlast 
	,\cceip_ob_tlv[0].tid[0] ,\cceip_ob_tlv[0].tstrb[7] 
	,\cceip_ob_tlv[0].tstrb[6] ,\cceip_ob_tlv[0].tstrb[5] 
	,\cceip_ob_tlv[0].tstrb[4] ,\cceip_ob_tlv[0].tstrb[3] 
	,\cceip_ob_tlv[0].tstrb[2] ,\cceip_ob_tlv[0].tstrb[1] 
	,\cceip_ob_tlv[0].tstrb[0] ,\cceip_ob_tlv[0].tuser[7] 
	,\cceip_ob_tlv[0].tuser[6] ,\cceip_ob_tlv[0].tuser[5] 
	,\cceip_ob_tlv[0].tuser[4] ,\cceip_ob_tlv[0].tuser[3] 
	,\cceip_ob_tlv[0].tuser[2] ,\cceip_ob_tlv[0].tuser[1] 
	,\cceip_ob_tlv[0].tuser[0] ,\cceip_ob_tlv[0].tdata[63] 
	,\cceip_ob_tlv[0].tdata[62] ,\cceip_ob_tlv[0].tdata[61] 
	,\cceip_ob_tlv[0].tdata[60] ,\cceip_ob_tlv[0].tdata[59] 
	,\cceip_ob_tlv[0].tdata[58] ,\cceip_ob_tlv[0].tdata[57] 
	,\cceip_ob_tlv[0].tdata[56] ,\cceip_ob_tlv[0].tdata[55] 
	,\cceip_ob_tlv[0].tdata[54] ,\cceip_ob_tlv[0].tdata[53] 
	,\cceip_ob_tlv[0].tdata[52] ,\cceip_ob_tlv[0].tdata[51] 
	,\cceip_ob_tlv[0].tdata[50] ,\cceip_ob_tlv[0].tdata[49] 
	,\cceip_ob_tlv[0].tdata[48] ,\cceip_ob_tlv[0].tdata[47] 
	,\cceip_ob_tlv[0].tdata[46] ,\cceip_ob_tlv[0].tdata[45] 
	,\cceip_ob_tlv[0].tdata[44] ,\cceip_ob_tlv[0].tdata[43] 
	,\cceip_ob_tlv[0].tdata[42] ,\cceip_ob_tlv[0].tdata[41] 
	,\cceip_ob_tlv[0].tdata[40] ,\cceip_ob_tlv[0].tdata[39] 
	,\cceip_ob_tlv[0].tdata[38] ,\cceip_ob_tlv[0].tdata[37] 
	,\cceip_ob_tlv[0].tdata[36] ,\cceip_ob_tlv[0].tdata[35] 
	,\cceip_ob_tlv[0].tdata[34] ,\cceip_ob_tlv[0].tdata[33] 
	,\cceip_ob_tlv[0].tdata[32] ,\cceip_ob_tlv[0].tdata[31] 
	,\cceip_ob_tlv[0].tdata[30] ,\cceip_ob_tlv[0].tdata[29] 
	,\cceip_ob_tlv[0].tdata[28] ,\cceip_ob_tlv[0].tdata[27] 
	,\cceip_ob_tlv[0].tdata[26] ,\cceip_ob_tlv[0].tdata[25] 
	,\cceip_ob_tlv[0].tdata[24] ,\cceip_ob_tlv[0].tdata[23] 
	,\cceip_ob_tlv[0].tdata[22] ,\cceip_ob_tlv[0].tdata[21] 
	,\cceip_ob_tlv[0].tdata[20] ,\cceip_ob_tlv[0].tdata[19] 
	,\cceip_ob_tlv[0].tdata[18] ,\cceip_ob_tlv[0].tdata[17] 
	,\cceip_ob_tlv[0].tdata[16] ,\cceip_ob_tlv[0].tdata[15] 
	,\cceip_ob_tlv[0].tdata[14] ,\cceip_ob_tlv[0].tdata[13] 
	,\cceip_ob_tlv[0].tdata[12] ,\cceip_ob_tlv[0].tdata[11] 
	,\cceip_ob_tlv[0].tdata[10] ,\cceip_ob_tlv[0].tdata[9] 
	,\cceip_ob_tlv[0].tdata[8] ,\cceip_ob_tlv[0].tdata[7] 
	,\cceip_ob_tlv[0].tdata[6] ,\cceip_ob_tlv[0].tdata[5] 
	,\cceip_ob_tlv[0].tdata[4] ,\cceip_ob_tlv[0].tdata[3] 
	,\cceip_ob_tlv[0].tdata[2] ,\cceip_ob_tlv[0].tdata[1] 
	,\cceip_ob_tlv[0].tdata[0] ;
input clk;
input rst_n;
input suppress_key_tlvs;
input cceip_encrypt_ob_wr;
input \cceip_encrypt_ob_tlv.insert ;
input [12:0] \cceip_encrypt_ob_tlv.ordern ;
input [7:0] \cceip_encrypt_ob_tlv.typen ;
input \cceip_encrypt_ob_tlv.sot ;
input \cceip_encrypt_ob_tlv.eot ;
input \cceip_encrypt_ob_tlv.tlast ;
input [0:0] \cceip_encrypt_ob_tlv.tid ;
input [7:0] \cceip_encrypt_ob_tlv.tstrb ;
input [7:0] \cceip_encrypt_ob_tlv.tuser ;
input [63:0] \cceip_encrypt_ob_tlv.tdata ;
wire [105:0] cceip_encrypt_ob_tlv;
input cceip_validate_ob_wr;
input \cceip_validate_ob_tlv.insert ;
input [12:0] \cceip_validate_ob_tlv.ordern ;
input [7:0] \cceip_validate_ob_tlv.typen ;
input \cceip_validate_ob_tlv.sot ;
input \cceip_validate_ob_tlv.eot ;
input \cceip_validate_ob_tlv.tlast ;
input [0:0] \cceip_validate_ob_tlv.tid ;
input [7:0] \cceip_validate_ob_tlv.tstrb ;
input [7:0] \cceip_validate_ob_tlv.tuser ;
input [63:0] \cceip_validate_ob_tlv.tdata ;
wire [105:0] cceip_validate_ob_tlv;
input [3:0] cceip_ob_full;
input [3:0] cceip_ob_afull;
wire encrypt_out_valid;
wire validate_out_valid;
wire [0:3] _zy_simnet_cceip_ob_wr_0_w$;
wire [0:423] _zy_simnet_cceip_ob_tlv_1_w$;
wire [0:105] _zy_simnet_encrypt_out_2_w$;
wire _zy_simnet_dio_3;
wire _zy_simnet_dio_4;
wire _zy_simnet_encrypt_out_ack_5_w$;
wire _zy_simnet_cio_6;
wire [0:105] _zy_simnet_validate_out_7_w$;
wire _zy_simnet_dio_8;
wire _zy_simnet_dio_9;
wire _zy_simnet_validate_out_ack_10_w$;
wire _zy_simnet_cio_11;
wire _zy_sva_brcm_cceip_1_reset_or;
wire _zy_sva_brcm_cceip_2_reset_or;
wire _zy_sva_brcm_cceip_3_reset_or;
wire _zy_sva_brcm_cceip_4_reset_or;
wire _zy_sva_b0_t;
wire _zy_sva_b1_t;
wire _zy_sva_b2_t;
wire _zy_sva_b3_t;
wire [0:0] cur_state;
wire [0:0] nxt_state;
wire [1:0] engine_select;
wire [1:0] nxt_engine_select;
wire [105:0] encrypt_out;
wire encrypt_out_ack;
wire [105:0] validate_out;
wire validate_out_ack;
wire [63:0] key_tlv_w0;
wire tlv_miscmp;
wire set_tlv_miscmp;
wire clr_tlv_miscmp;
wire [31:0] i;
`_2_ wire [0:0] _zy_sva_brcm_cceip_1_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_cceip_1_cpass;
`_2_ wire _zy_sva_b0;
`_2_ wire [0:0] _zy_sva_brcm_cceip_2_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_cceip_2_cpass;
`_2_ wire _zy_sva_b1;
`_2_ wire [0:0] _zy_sva_brcm_cceip_3_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_cceip_3_cpass;
`_2_ wire _zy_sva_b2;
`_2_ wire [0:0] _zy_sva_brcm_cceip_4_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_cceip_4_cpass;
`_2_ wire _zy_sva_b3;
supply0 n324;
supply1 n517;
wire \encrypt_out.insert ;
wire [12:0] \encrypt_out.ordern ;
wire [7:0] \encrypt_out.typen ;
wire \encrypt_out.sot ;
wire \encrypt_out.eot ;
wire \encrypt_out.tlast ;
wire [0:0] \encrypt_out.tid ;
wire [7:0] \encrypt_out.tstrb ;
wire [7:0] \encrypt_out.tuser ;
wire [63:0] \encrypt_out.tdata ;
wire \validate_out.insert ;
wire [12:0] \validate_out.ordern ;
wire [7:0] \validate_out.typen ;
wire \validate_out.sot ;
wire \validate_out.eot ;
wire \validate_out.tlast ;
wire [0:0] \validate_out.tid ;
wire [7:0] \validate_out.tstrb ;
wire [7:0] \validate_out.tuser ;
wire [63:0] \validate_out.tdata ;
wire [1:0] \key_tlv_w0.tlv_bip2 ;
wire [18:0] \key_tlv_w0.resv0 ;
wire [10:0] \key_tlv_w0.tlv_frame_num ;
wire [3:0] \key_tlv_w0.resv1 ;
wire [3:0] \key_tlv_w0.tlv_eng_id ;
wire [7:0] \key_tlv_w0.tlv_seq_num ;
wire [7:0] \key_tlv_w0.tlv_len ;
wire [7:0] \key_tlv_w0.tlv_type ;
tran (\cceip_ob_tlv[0][0] , \cceip_ob_tlv[0].tdata[0] );
tran (\cceip_ob_tlv[0][1] , \cceip_ob_tlv[0].tdata[1] );
tran (\cceip_ob_tlv[0][2] , \cceip_ob_tlv[0].tdata[2] );
tran (\cceip_ob_tlv[0][3] , \cceip_ob_tlv[0].tdata[3] );
tran (\cceip_ob_tlv[0][4] , \cceip_ob_tlv[0].tdata[4] );
tran (\cceip_ob_tlv[0][5] , \cceip_ob_tlv[0].tdata[5] );
tran (\cceip_ob_tlv[0][6] , \cceip_ob_tlv[0].tdata[6] );
tran (\cceip_ob_tlv[0][7] , \cceip_ob_tlv[0].tdata[7] );
tran (\cceip_ob_tlv[0][8] , \cceip_ob_tlv[0].tdata[8] );
tran (\cceip_ob_tlv[0][9] , \cceip_ob_tlv[0].tdata[9] );
tran (\cceip_ob_tlv[0][10] , \cceip_ob_tlv[0].tdata[10] );
tran (\cceip_ob_tlv[0][11] , \cceip_ob_tlv[0].tdata[11] );
tran (\cceip_ob_tlv[0][12] , \cceip_ob_tlv[0].tdata[12] );
tran (\cceip_ob_tlv[0][13] , \cceip_ob_tlv[0].tdata[13] );
tran (\cceip_ob_tlv[0][14] , \cceip_ob_tlv[0].tdata[14] );
tran (\cceip_ob_tlv[0][15] , \cceip_ob_tlv[0].tdata[15] );
tran (\cceip_ob_tlv[0][16] , \cceip_ob_tlv[0].tdata[16] );
tran (\cceip_ob_tlv[0][17] , \cceip_ob_tlv[0].tdata[17] );
tran (\cceip_ob_tlv[0][18] , \cceip_ob_tlv[0].tdata[18] );
tran (\cceip_ob_tlv[0][19] , \cceip_ob_tlv[0].tdata[19] );
tran (\cceip_ob_tlv[0][20] , \cceip_ob_tlv[0].tdata[20] );
tran (\cceip_ob_tlv[0][21] , \cceip_ob_tlv[0].tdata[21] );
tran (\cceip_ob_tlv[0][22] , \cceip_ob_tlv[0].tdata[22] );
tran (\cceip_ob_tlv[0][23] , \cceip_ob_tlv[0].tdata[23] );
tran (\cceip_ob_tlv[0][24] , \cceip_ob_tlv[0].tdata[24] );
tran (\cceip_ob_tlv[0][25] , \cceip_ob_tlv[0].tdata[25] );
tran (\cceip_ob_tlv[0][26] , \cceip_ob_tlv[0].tdata[26] );
tran (\cceip_ob_tlv[0][27] , \cceip_ob_tlv[0].tdata[27] );
tran (\cceip_ob_tlv[0][28] , \cceip_ob_tlv[0].tdata[28] );
tran (\cceip_ob_tlv[0][29] , \cceip_ob_tlv[0].tdata[29] );
tran (\cceip_ob_tlv[0][30] , \cceip_ob_tlv[0].tdata[30] );
tran (\cceip_ob_tlv[0][31] , \cceip_ob_tlv[0].tdata[31] );
tran (\cceip_ob_tlv[0][32] , \cceip_ob_tlv[0].tdata[32] );
tran (\cceip_ob_tlv[0][33] , \cceip_ob_tlv[0].tdata[33] );
tran (\cceip_ob_tlv[0][34] , \cceip_ob_tlv[0].tdata[34] );
tran (\cceip_ob_tlv[0][35] , \cceip_ob_tlv[0].tdata[35] );
tran (\cceip_ob_tlv[0][36] , \cceip_ob_tlv[0].tdata[36] );
tran (\cceip_ob_tlv[0][37] , \cceip_ob_tlv[0].tdata[37] );
tran (\cceip_ob_tlv[0][38] , \cceip_ob_tlv[0].tdata[38] );
tran (\cceip_ob_tlv[0][39] , \cceip_ob_tlv[0].tdata[39] );
tran (\cceip_ob_tlv[0][40] , \cceip_ob_tlv[0].tdata[40] );
tran (\cceip_ob_tlv[0][41] , \cceip_ob_tlv[0].tdata[41] );
tran (\cceip_ob_tlv[0][42] , \cceip_ob_tlv[0].tdata[42] );
tran (\cceip_ob_tlv[0][43] , \cceip_ob_tlv[0].tdata[43] );
tran (\cceip_ob_tlv[0][44] , \cceip_ob_tlv[0].tdata[44] );
tran (\cceip_ob_tlv[0][45] , \cceip_ob_tlv[0].tdata[45] );
tran (\cceip_ob_tlv[0][46] , \cceip_ob_tlv[0].tdata[46] );
tran (\cceip_ob_tlv[0][47] , \cceip_ob_tlv[0].tdata[47] );
tran (\cceip_ob_tlv[0][48] , \cceip_ob_tlv[0].tdata[48] );
tran (\cceip_ob_tlv[0][49] , \cceip_ob_tlv[0].tdata[49] );
tran (\cceip_ob_tlv[0][50] , \cceip_ob_tlv[0].tdata[50] );
tran (\cceip_ob_tlv[0][51] , \cceip_ob_tlv[0].tdata[51] );
tran (\cceip_ob_tlv[0][52] , \cceip_ob_tlv[0].tdata[52] );
tran (\cceip_ob_tlv[0][53] , \cceip_ob_tlv[0].tdata[53] );
tran (\cceip_ob_tlv[0][54] , \cceip_ob_tlv[0].tdata[54] );
tran (\cceip_ob_tlv[0][55] , \cceip_ob_tlv[0].tdata[55] );
tran (\cceip_ob_tlv[0][56] , \cceip_ob_tlv[0].tdata[56] );
tran (\cceip_ob_tlv[0][57] , \cceip_ob_tlv[0].tdata[57] );
tran (\cceip_ob_tlv[0][58] , \cceip_ob_tlv[0].tdata[58] );
tran (\cceip_ob_tlv[0][59] , \cceip_ob_tlv[0].tdata[59] );
tran (\cceip_ob_tlv[0][60] , \cceip_ob_tlv[0].tdata[60] );
tran (\cceip_ob_tlv[0][61] , \cceip_ob_tlv[0].tdata[61] );
tran (\cceip_ob_tlv[0][62] , \cceip_ob_tlv[0].tdata[62] );
tran (\cceip_ob_tlv[0][63] , \cceip_ob_tlv[0].tdata[63] );
tran (\cceip_ob_tlv[0][64] , \cceip_ob_tlv[0].tuser[0] );
tran (\cceip_ob_tlv[0][65] , \cceip_ob_tlv[0].tuser[1] );
tran (\cceip_ob_tlv[0][66] , \cceip_ob_tlv[0].tuser[2] );
tran (\cceip_ob_tlv[0][67] , \cceip_ob_tlv[0].tuser[3] );
tran (\cceip_ob_tlv[0][68] , \cceip_ob_tlv[0].tuser[4] );
tran (\cceip_ob_tlv[0][69] , \cceip_ob_tlv[0].tuser[5] );
tran (\cceip_ob_tlv[0][70] , \cceip_ob_tlv[0].tuser[6] );
tran (\cceip_ob_tlv[0][71] , \cceip_ob_tlv[0].tuser[7] );
tran (\cceip_ob_tlv[0][72] , \cceip_ob_tlv[0].tstrb[0] );
tran (\cceip_ob_tlv[0][73] , \cceip_ob_tlv[0].tstrb[1] );
tran (\cceip_ob_tlv[0][74] , \cceip_ob_tlv[0].tstrb[2] );
tran (\cceip_ob_tlv[0][75] , \cceip_ob_tlv[0].tstrb[3] );
tran (\cceip_ob_tlv[0][76] , \cceip_ob_tlv[0].tstrb[4] );
tran (\cceip_ob_tlv[0][77] , \cceip_ob_tlv[0].tstrb[5] );
tran (\cceip_ob_tlv[0][78] , \cceip_ob_tlv[0].tstrb[6] );
tran (\cceip_ob_tlv[0][79] , \cceip_ob_tlv[0].tstrb[7] );
tran (\cceip_ob_tlv[0][80] , \cceip_ob_tlv[0].tid[0] );
tran (\cceip_ob_tlv[0][81] , \cceip_ob_tlv[0].tlast );
tran (\cceip_ob_tlv[0][82] , \cceip_ob_tlv[0].eot );
tran (\cceip_ob_tlv[0][83] , \cceip_ob_tlv[0].sot );
tran (\cceip_ob_tlv[0][84] , \cceip_ob_tlv[0].typen[0] );
tran (\cceip_ob_tlv[0][85] , \cceip_ob_tlv[0].typen[1] );
tran (\cceip_ob_tlv[0][86] , \cceip_ob_tlv[0].typen[2] );
tran (\cceip_ob_tlv[0][87] , \cceip_ob_tlv[0].typen[3] );
tran (\cceip_ob_tlv[0][88] , \cceip_ob_tlv[0].typen[4] );
tran (\cceip_ob_tlv[0][89] , \cceip_ob_tlv[0].typen[5] );
tran (\cceip_ob_tlv[0][90] , \cceip_ob_tlv[0].typen[6] );
tran (\cceip_ob_tlv[0][91] , \cceip_ob_tlv[0].typen[7] );
tran (\cceip_ob_tlv[0][92] , \cceip_ob_tlv[0].ordern[0] );
tran (\cceip_ob_tlv[0][93] , \cceip_ob_tlv[0].ordern[1] );
tran (\cceip_ob_tlv[0][94] , \cceip_ob_tlv[0].ordern[2] );
tran (\cceip_ob_tlv[0][95] , \cceip_ob_tlv[0].ordern[3] );
tran (\cceip_ob_tlv[0][96] , \cceip_ob_tlv[0].ordern[4] );
tran (\cceip_ob_tlv[0][97] , \cceip_ob_tlv[0].ordern[5] );
tran (\cceip_ob_tlv[0][98] , \cceip_ob_tlv[0].ordern[6] );
tran (\cceip_ob_tlv[0][99] , \cceip_ob_tlv[0].ordern[7] );
tran (\cceip_ob_tlv[0][100] , \cceip_ob_tlv[0].ordern[8] );
tran (\cceip_ob_tlv[0][101] , \cceip_ob_tlv[0].ordern[9] );
tran (\cceip_ob_tlv[0][102] , \cceip_ob_tlv[0].ordern[10] );
tran (\cceip_ob_tlv[0][103] , \cceip_ob_tlv[0].ordern[11] );
tran (\cceip_ob_tlv[0][104] , \cceip_ob_tlv[0].ordern[12] );
tran (\cceip_ob_tlv[0][105] , \cceip_ob_tlv[0].insert );
tran (\cceip_ob_tlv[1][0] , \cceip_ob_tlv[1].tdata[0] );
tran (\cceip_ob_tlv[1][1] , \cceip_ob_tlv[1].tdata[1] );
tran (\cceip_ob_tlv[1][2] , \cceip_ob_tlv[1].tdata[2] );
tran (\cceip_ob_tlv[1][3] , \cceip_ob_tlv[1].tdata[3] );
tran (\cceip_ob_tlv[1][4] , \cceip_ob_tlv[1].tdata[4] );
tran (\cceip_ob_tlv[1][5] , \cceip_ob_tlv[1].tdata[5] );
tran (\cceip_ob_tlv[1][6] , \cceip_ob_tlv[1].tdata[6] );
tran (\cceip_ob_tlv[1][7] , \cceip_ob_tlv[1].tdata[7] );
tran (\cceip_ob_tlv[1][8] , \cceip_ob_tlv[1].tdata[8] );
tran (\cceip_ob_tlv[1][9] , \cceip_ob_tlv[1].tdata[9] );
tran (\cceip_ob_tlv[1][10] , \cceip_ob_tlv[1].tdata[10] );
tran (\cceip_ob_tlv[1][11] , \cceip_ob_tlv[1].tdata[11] );
tran (\cceip_ob_tlv[1][12] , \cceip_ob_tlv[1].tdata[12] );
tran (\cceip_ob_tlv[1][13] , \cceip_ob_tlv[1].tdata[13] );
tran (\cceip_ob_tlv[1][14] , \cceip_ob_tlv[1].tdata[14] );
tran (\cceip_ob_tlv[1][15] , \cceip_ob_tlv[1].tdata[15] );
tran (\cceip_ob_tlv[1][16] , \cceip_ob_tlv[1].tdata[16] );
tran (\cceip_ob_tlv[1][17] , \cceip_ob_tlv[1].tdata[17] );
tran (\cceip_ob_tlv[1][18] , \cceip_ob_tlv[1].tdata[18] );
tran (\cceip_ob_tlv[1][19] , \cceip_ob_tlv[1].tdata[19] );
tran (\cceip_ob_tlv[1][20] , \cceip_ob_tlv[1].tdata[20] );
tran (\cceip_ob_tlv[1][21] , \cceip_ob_tlv[1].tdata[21] );
tran (\cceip_ob_tlv[1][22] , \cceip_ob_tlv[1].tdata[22] );
tran (\cceip_ob_tlv[1][23] , \cceip_ob_tlv[1].tdata[23] );
tran (\cceip_ob_tlv[1][24] , \cceip_ob_tlv[1].tdata[24] );
tran (\cceip_ob_tlv[1][25] , \cceip_ob_tlv[1].tdata[25] );
tran (\cceip_ob_tlv[1][26] , \cceip_ob_tlv[1].tdata[26] );
tran (\cceip_ob_tlv[1][27] , \cceip_ob_tlv[1].tdata[27] );
tran (\cceip_ob_tlv[1][28] , \cceip_ob_tlv[1].tdata[28] );
tran (\cceip_ob_tlv[1][29] , \cceip_ob_tlv[1].tdata[29] );
tran (\cceip_ob_tlv[1][30] , \cceip_ob_tlv[1].tdata[30] );
tran (\cceip_ob_tlv[1][31] , \cceip_ob_tlv[1].tdata[31] );
tran (\cceip_ob_tlv[1][32] , \cceip_ob_tlv[1].tdata[32] );
tran (\cceip_ob_tlv[1][33] , \cceip_ob_tlv[1].tdata[33] );
tran (\cceip_ob_tlv[1][34] , \cceip_ob_tlv[1].tdata[34] );
tran (\cceip_ob_tlv[1][35] , \cceip_ob_tlv[1].tdata[35] );
tran (\cceip_ob_tlv[1][36] , \cceip_ob_tlv[1].tdata[36] );
tran (\cceip_ob_tlv[1][37] , \cceip_ob_tlv[1].tdata[37] );
tran (\cceip_ob_tlv[1][38] , \cceip_ob_tlv[1].tdata[38] );
tran (\cceip_ob_tlv[1][39] , \cceip_ob_tlv[1].tdata[39] );
tran (\cceip_ob_tlv[1][40] , \cceip_ob_tlv[1].tdata[40] );
tran (\cceip_ob_tlv[1][41] , \cceip_ob_tlv[1].tdata[41] );
tran (\cceip_ob_tlv[1][42] , \cceip_ob_tlv[1].tdata[42] );
tran (\cceip_ob_tlv[1][43] , \cceip_ob_tlv[1].tdata[43] );
tran (\cceip_ob_tlv[1][44] , \cceip_ob_tlv[1].tdata[44] );
tran (\cceip_ob_tlv[1][45] , \cceip_ob_tlv[1].tdata[45] );
tran (\cceip_ob_tlv[1][46] , \cceip_ob_tlv[1].tdata[46] );
tran (\cceip_ob_tlv[1][47] , \cceip_ob_tlv[1].tdata[47] );
tran (\cceip_ob_tlv[1][48] , \cceip_ob_tlv[1].tdata[48] );
tran (\cceip_ob_tlv[1][49] , \cceip_ob_tlv[1].tdata[49] );
tran (\cceip_ob_tlv[1][50] , \cceip_ob_tlv[1].tdata[50] );
tran (\cceip_ob_tlv[1][51] , \cceip_ob_tlv[1].tdata[51] );
tran (\cceip_ob_tlv[1][52] , \cceip_ob_tlv[1].tdata[52] );
tran (\cceip_ob_tlv[1][53] , \cceip_ob_tlv[1].tdata[53] );
tran (\cceip_ob_tlv[1][54] , \cceip_ob_tlv[1].tdata[54] );
tran (\cceip_ob_tlv[1][55] , \cceip_ob_tlv[1].tdata[55] );
tran (\cceip_ob_tlv[1][56] , \cceip_ob_tlv[1].tdata[56] );
tran (\cceip_ob_tlv[1][57] , \cceip_ob_tlv[1].tdata[57] );
tran (\cceip_ob_tlv[1][58] , \cceip_ob_tlv[1].tdata[58] );
tran (\cceip_ob_tlv[1][59] , \cceip_ob_tlv[1].tdata[59] );
tran (\cceip_ob_tlv[1][60] , \cceip_ob_tlv[1].tdata[60] );
tran (\cceip_ob_tlv[1][61] , \cceip_ob_tlv[1].tdata[61] );
tran (\cceip_ob_tlv[1][62] , \cceip_ob_tlv[1].tdata[62] );
tran (\cceip_ob_tlv[1][63] , \cceip_ob_tlv[1].tdata[63] );
tran (\cceip_ob_tlv[1][64] , \cceip_ob_tlv[1].tuser[0] );
tran (\cceip_ob_tlv[1][65] , \cceip_ob_tlv[1].tuser[1] );
tran (\cceip_ob_tlv[1][66] , \cceip_ob_tlv[1].tuser[2] );
tran (\cceip_ob_tlv[1][67] , \cceip_ob_tlv[1].tuser[3] );
tran (\cceip_ob_tlv[1][68] , \cceip_ob_tlv[1].tuser[4] );
tran (\cceip_ob_tlv[1][69] , \cceip_ob_tlv[1].tuser[5] );
tran (\cceip_ob_tlv[1][70] , \cceip_ob_tlv[1].tuser[6] );
tran (\cceip_ob_tlv[1][71] , \cceip_ob_tlv[1].tuser[7] );
tran (\cceip_ob_tlv[1][72] , \cceip_ob_tlv[1].tstrb[0] );
tran (\cceip_ob_tlv[1][73] , \cceip_ob_tlv[1].tstrb[1] );
tran (\cceip_ob_tlv[1][74] , \cceip_ob_tlv[1].tstrb[2] );
tran (\cceip_ob_tlv[1][75] , \cceip_ob_tlv[1].tstrb[3] );
tran (\cceip_ob_tlv[1][76] , \cceip_ob_tlv[1].tstrb[4] );
tran (\cceip_ob_tlv[1][77] , \cceip_ob_tlv[1].tstrb[5] );
tran (\cceip_ob_tlv[1][78] , \cceip_ob_tlv[1].tstrb[6] );
tran (\cceip_ob_tlv[1][79] , \cceip_ob_tlv[1].tstrb[7] );
tran (\cceip_ob_tlv[1][80] , \cceip_ob_tlv[1].tid[0] );
tran (\cceip_ob_tlv[1][81] , \cceip_ob_tlv[1].tlast );
tran (\cceip_ob_tlv[1][82] , \cceip_ob_tlv[1].eot );
tran (\cceip_ob_tlv[1][83] , \cceip_ob_tlv[1].sot );
tran (\cceip_ob_tlv[1][84] , \cceip_ob_tlv[1].typen[0] );
tran (\cceip_ob_tlv[1][85] , \cceip_ob_tlv[1].typen[1] );
tran (\cceip_ob_tlv[1][86] , \cceip_ob_tlv[1].typen[2] );
tran (\cceip_ob_tlv[1][87] , \cceip_ob_tlv[1].typen[3] );
tran (\cceip_ob_tlv[1][88] , \cceip_ob_tlv[1].typen[4] );
tran (\cceip_ob_tlv[1][89] , \cceip_ob_tlv[1].typen[5] );
tran (\cceip_ob_tlv[1][90] , \cceip_ob_tlv[1].typen[6] );
tran (\cceip_ob_tlv[1][91] , \cceip_ob_tlv[1].typen[7] );
tran (\cceip_ob_tlv[1][92] , \cceip_ob_tlv[1].ordern[0] );
tran (\cceip_ob_tlv[1][93] , \cceip_ob_tlv[1].ordern[1] );
tran (\cceip_ob_tlv[1][94] , \cceip_ob_tlv[1].ordern[2] );
tran (\cceip_ob_tlv[1][95] , \cceip_ob_tlv[1].ordern[3] );
tran (\cceip_ob_tlv[1][96] , \cceip_ob_tlv[1].ordern[4] );
tran (\cceip_ob_tlv[1][97] , \cceip_ob_tlv[1].ordern[5] );
tran (\cceip_ob_tlv[1][98] , \cceip_ob_tlv[1].ordern[6] );
tran (\cceip_ob_tlv[1][99] , \cceip_ob_tlv[1].ordern[7] );
tran (\cceip_ob_tlv[1][100] , \cceip_ob_tlv[1].ordern[8] );
tran (\cceip_ob_tlv[1][101] , \cceip_ob_tlv[1].ordern[9] );
tran (\cceip_ob_tlv[1][102] , \cceip_ob_tlv[1].ordern[10] );
tran (\cceip_ob_tlv[1][103] , \cceip_ob_tlv[1].ordern[11] );
tran (\cceip_ob_tlv[1][104] , \cceip_ob_tlv[1].ordern[12] );
tran (\cceip_ob_tlv[1][105] , \cceip_ob_tlv[1].insert );
tran (\cceip_ob_tlv[2][0] , \cceip_ob_tlv[2].tdata[0] );
tran (\cceip_ob_tlv[2][1] , \cceip_ob_tlv[2].tdata[1] );
tran (\cceip_ob_tlv[2][2] , \cceip_ob_tlv[2].tdata[2] );
tran (\cceip_ob_tlv[2][3] , \cceip_ob_tlv[2].tdata[3] );
tran (\cceip_ob_tlv[2][4] , \cceip_ob_tlv[2].tdata[4] );
tran (\cceip_ob_tlv[2][5] , \cceip_ob_tlv[2].tdata[5] );
tran (\cceip_ob_tlv[2][6] , \cceip_ob_tlv[2].tdata[6] );
tran (\cceip_ob_tlv[2][7] , \cceip_ob_tlv[2].tdata[7] );
tran (\cceip_ob_tlv[2][8] , \cceip_ob_tlv[2].tdata[8] );
tran (\cceip_ob_tlv[2][9] , \cceip_ob_tlv[2].tdata[9] );
tran (\cceip_ob_tlv[2][10] , \cceip_ob_tlv[2].tdata[10] );
tran (\cceip_ob_tlv[2][11] , \cceip_ob_tlv[2].tdata[11] );
tran (\cceip_ob_tlv[2][12] , \cceip_ob_tlv[2].tdata[12] );
tran (\cceip_ob_tlv[2][13] , \cceip_ob_tlv[2].tdata[13] );
tran (\cceip_ob_tlv[2][14] , \cceip_ob_tlv[2].tdata[14] );
tran (\cceip_ob_tlv[2][15] , \cceip_ob_tlv[2].tdata[15] );
tran (\cceip_ob_tlv[2][16] , \cceip_ob_tlv[2].tdata[16] );
tran (\cceip_ob_tlv[2][17] , \cceip_ob_tlv[2].tdata[17] );
tran (\cceip_ob_tlv[2][18] , \cceip_ob_tlv[2].tdata[18] );
tran (\cceip_ob_tlv[2][19] , \cceip_ob_tlv[2].tdata[19] );
tran (\cceip_ob_tlv[2][20] , \cceip_ob_tlv[2].tdata[20] );
tran (\cceip_ob_tlv[2][21] , \cceip_ob_tlv[2].tdata[21] );
tran (\cceip_ob_tlv[2][22] , \cceip_ob_tlv[2].tdata[22] );
tran (\cceip_ob_tlv[2][23] , \cceip_ob_tlv[2].tdata[23] );
tran (\cceip_ob_tlv[2][24] , \cceip_ob_tlv[2].tdata[24] );
tran (\cceip_ob_tlv[2][25] , \cceip_ob_tlv[2].tdata[25] );
tran (\cceip_ob_tlv[2][26] , \cceip_ob_tlv[2].tdata[26] );
tran (\cceip_ob_tlv[2][27] , \cceip_ob_tlv[2].tdata[27] );
tran (\cceip_ob_tlv[2][28] , \cceip_ob_tlv[2].tdata[28] );
tran (\cceip_ob_tlv[2][29] , \cceip_ob_tlv[2].tdata[29] );
tran (\cceip_ob_tlv[2][30] , \cceip_ob_tlv[2].tdata[30] );
tran (\cceip_ob_tlv[2][31] , \cceip_ob_tlv[2].tdata[31] );
tran (\cceip_ob_tlv[2][32] , \cceip_ob_tlv[2].tdata[32] );
tran (\cceip_ob_tlv[2][33] , \cceip_ob_tlv[2].tdata[33] );
tran (\cceip_ob_tlv[2][34] , \cceip_ob_tlv[2].tdata[34] );
tran (\cceip_ob_tlv[2][35] , \cceip_ob_tlv[2].tdata[35] );
tran (\cceip_ob_tlv[2][36] , \cceip_ob_tlv[2].tdata[36] );
tran (\cceip_ob_tlv[2][37] , \cceip_ob_tlv[2].tdata[37] );
tran (\cceip_ob_tlv[2][38] , \cceip_ob_tlv[2].tdata[38] );
tran (\cceip_ob_tlv[2][39] , \cceip_ob_tlv[2].tdata[39] );
tran (\cceip_ob_tlv[2][40] , \cceip_ob_tlv[2].tdata[40] );
tran (\cceip_ob_tlv[2][41] , \cceip_ob_tlv[2].tdata[41] );
tran (\cceip_ob_tlv[2][42] , \cceip_ob_tlv[2].tdata[42] );
tran (\cceip_ob_tlv[2][43] , \cceip_ob_tlv[2].tdata[43] );
tran (\cceip_ob_tlv[2][44] , \cceip_ob_tlv[2].tdata[44] );
tran (\cceip_ob_tlv[2][45] , \cceip_ob_tlv[2].tdata[45] );
tran (\cceip_ob_tlv[2][46] , \cceip_ob_tlv[2].tdata[46] );
tran (\cceip_ob_tlv[2][47] , \cceip_ob_tlv[2].tdata[47] );
tran (\cceip_ob_tlv[2][48] , \cceip_ob_tlv[2].tdata[48] );
tran (\cceip_ob_tlv[2][49] , \cceip_ob_tlv[2].tdata[49] );
tran (\cceip_ob_tlv[2][50] , \cceip_ob_tlv[2].tdata[50] );
tran (\cceip_ob_tlv[2][51] , \cceip_ob_tlv[2].tdata[51] );
tran (\cceip_ob_tlv[2][52] , \cceip_ob_tlv[2].tdata[52] );
tran (\cceip_ob_tlv[2][53] , \cceip_ob_tlv[2].tdata[53] );
tran (\cceip_ob_tlv[2][54] , \cceip_ob_tlv[2].tdata[54] );
tran (\cceip_ob_tlv[2][55] , \cceip_ob_tlv[2].tdata[55] );
tran (\cceip_ob_tlv[2][56] , \cceip_ob_tlv[2].tdata[56] );
tran (\cceip_ob_tlv[2][57] , \cceip_ob_tlv[2].tdata[57] );
tran (\cceip_ob_tlv[2][58] , \cceip_ob_tlv[2].tdata[58] );
tran (\cceip_ob_tlv[2][59] , \cceip_ob_tlv[2].tdata[59] );
tran (\cceip_ob_tlv[2][60] , \cceip_ob_tlv[2].tdata[60] );
tran (\cceip_ob_tlv[2][61] , \cceip_ob_tlv[2].tdata[61] );
tran (\cceip_ob_tlv[2][62] , \cceip_ob_tlv[2].tdata[62] );
tran (\cceip_ob_tlv[2][63] , \cceip_ob_tlv[2].tdata[63] );
tran (\cceip_ob_tlv[2][64] , \cceip_ob_tlv[2].tuser[0] );
tran (\cceip_ob_tlv[2][65] , \cceip_ob_tlv[2].tuser[1] );
tran (\cceip_ob_tlv[2][66] , \cceip_ob_tlv[2].tuser[2] );
tran (\cceip_ob_tlv[2][67] , \cceip_ob_tlv[2].tuser[3] );
tran (\cceip_ob_tlv[2][68] , \cceip_ob_tlv[2].tuser[4] );
tran (\cceip_ob_tlv[2][69] , \cceip_ob_tlv[2].tuser[5] );
tran (\cceip_ob_tlv[2][70] , \cceip_ob_tlv[2].tuser[6] );
tran (\cceip_ob_tlv[2][71] , \cceip_ob_tlv[2].tuser[7] );
tran (\cceip_ob_tlv[2][72] , \cceip_ob_tlv[2].tstrb[0] );
tran (\cceip_ob_tlv[2][73] , \cceip_ob_tlv[2].tstrb[1] );
tran (\cceip_ob_tlv[2][74] , \cceip_ob_tlv[2].tstrb[2] );
tran (\cceip_ob_tlv[2][75] , \cceip_ob_tlv[2].tstrb[3] );
tran (\cceip_ob_tlv[2][76] , \cceip_ob_tlv[2].tstrb[4] );
tran (\cceip_ob_tlv[2][77] , \cceip_ob_tlv[2].tstrb[5] );
tran (\cceip_ob_tlv[2][78] , \cceip_ob_tlv[2].tstrb[6] );
tran (\cceip_ob_tlv[2][79] , \cceip_ob_tlv[2].tstrb[7] );
tran (\cceip_ob_tlv[2][80] , \cceip_ob_tlv[2].tid[0] );
tran (\cceip_ob_tlv[2][81] , \cceip_ob_tlv[2].tlast );
tran (\cceip_ob_tlv[2][82] , \cceip_ob_tlv[2].eot );
tran (\cceip_ob_tlv[2][83] , \cceip_ob_tlv[2].sot );
tran (\cceip_ob_tlv[2][84] , \cceip_ob_tlv[2].typen[0] );
tran (\cceip_ob_tlv[2][85] , \cceip_ob_tlv[2].typen[1] );
tran (\cceip_ob_tlv[2][86] , \cceip_ob_tlv[2].typen[2] );
tran (\cceip_ob_tlv[2][87] , \cceip_ob_tlv[2].typen[3] );
tran (\cceip_ob_tlv[2][88] , \cceip_ob_tlv[2].typen[4] );
tran (\cceip_ob_tlv[2][89] , \cceip_ob_tlv[2].typen[5] );
tran (\cceip_ob_tlv[2][90] , \cceip_ob_tlv[2].typen[6] );
tran (\cceip_ob_tlv[2][91] , \cceip_ob_tlv[2].typen[7] );
tran (\cceip_ob_tlv[2][92] , \cceip_ob_tlv[2].ordern[0] );
tran (\cceip_ob_tlv[2][93] , \cceip_ob_tlv[2].ordern[1] );
tran (\cceip_ob_tlv[2][94] , \cceip_ob_tlv[2].ordern[2] );
tran (\cceip_ob_tlv[2][95] , \cceip_ob_tlv[2].ordern[3] );
tran (\cceip_ob_tlv[2][96] , \cceip_ob_tlv[2].ordern[4] );
tran (\cceip_ob_tlv[2][97] , \cceip_ob_tlv[2].ordern[5] );
tran (\cceip_ob_tlv[2][98] , \cceip_ob_tlv[2].ordern[6] );
tran (\cceip_ob_tlv[2][99] , \cceip_ob_tlv[2].ordern[7] );
tran (\cceip_ob_tlv[2][100] , \cceip_ob_tlv[2].ordern[8] );
tran (\cceip_ob_tlv[2][101] , \cceip_ob_tlv[2].ordern[9] );
tran (\cceip_ob_tlv[2][102] , \cceip_ob_tlv[2].ordern[10] );
tran (\cceip_ob_tlv[2][103] , \cceip_ob_tlv[2].ordern[11] );
tran (\cceip_ob_tlv[2][104] , \cceip_ob_tlv[2].ordern[12] );
tran (\cceip_ob_tlv[2][105] , \cceip_ob_tlv[2].insert );
tran (\cceip_ob_tlv[3][0] , \cceip_ob_tlv[3].tdata[0] );
tran (\cceip_ob_tlv[3][1] , \cceip_ob_tlv[3].tdata[1] );
tran (\cceip_ob_tlv[3][2] , \cceip_ob_tlv[3].tdata[2] );
tran (\cceip_ob_tlv[3][3] , \cceip_ob_tlv[3].tdata[3] );
tran (\cceip_ob_tlv[3][4] , \cceip_ob_tlv[3].tdata[4] );
tran (\cceip_ob_tlv[3][5] , \cceip_ob_tlv[3].tdata[5] );
tran (\cceip_ob_tlv[3][6] , \cceip_ob_tlv[3].tdata[6] );
tran (\cceip_ob_tlv[3][7] , \cceip_ob_tlv[3].tdata[7] );
tran (\cceip_ob_tlv[3][8] , \cceip_ob_tlv[3].tdata[8] );
tran (\cceip_ob_tlv[3][9] , \cceip_ob_tlv[3].tdata[9] );
tran (\cceip_ob_tlv[3][10] , \cceip_ob_tlv[3].tdata[10] );
tran (\cceip_ob_tlv[3][11] , \cceip_ob_tlv[3].tdata[11] );
tran (\cceip_ob_tlv[3][12] , \cceip_ob_tlv[3].tdata[12] );
tran (\cceip_ob_tlv[3][13] , \cceip_ob_tlv[3].tdata[13] );
tran (\cceip_ob_tlv[3][14] , \cceip_ob_tlv[3].tdata[14] );
tran (\cceip_ob_tlv[3][15] , \cceip_ob_tlv[3].tdata[15] );
tran (\cceip_ob_tlv[3][16] , \cceip_ob_tlv[3].tdata[16] );
tran (\cceip_ob_tlv[3][17] , \cceip_ob_tlv[3].tdata[17] );
tran (\cceip_ob_tlv[3][18] , \cceip_ob_tlv[3].tdata[18] );
tran (\cceip_ob_tlv[3][19] , \cceip_ob_tlv[3].tdata[19] );
tran (\cceip_ob_tlv[3][20] , \cceip_ob_tlv[3].tdata[20] );
tran (\cceip_ob_tlv[3][21] , \cceip_ob_tlv[3].tdata[21] );
tran (\cceip_ob_tlv[3][22] , \cceip_ob_tlv[3].tdata[22] );
tran (\cceip_ob_tlv[3][23] , \cceip_ob_tlv[3].tdata[23] );
tran (\cceip_ob_tlv[3][24] , \cceip_ob_tlv[3].tdata[24] );
tran (\cceip_ob_tlv[3][25] , \cceip_ob_tlv[3].tdata[25] );
tran (\cceip_ob_tlv[3][26] , \cceip_ob_tlv[3].tdata[26] );
tran (\cceip_ob_tlv[3][27] , \cceip_ob_tlv[3].tdata[27] );
tran (\cceip_ob_tlv[3][28] , \cceip_ob_tlv[3].tdata[28] );
tran (\cceip_ob_tlv[3][29] , \cceip_ob_tlv[3].tdata[29] );
tran (\cceip_ob_tlv[3][30] , \cceip_ob_tlv[3].tdata[30] );
tran (\cceip_ob_tlv[3][31] , \cceip_ob_tlv[3].tdata[31] );
tran (\cceip_ob_tlv[3][32] , \cceip_ob_tlv[3].tdata[32] );
tran (\cceip_ob_tlv[3][33] , \cceip_ob_tlv[3].tdata[33] );
tran (\cceip_ob_tlv[3][34] , \cceip_ob_tlv[3].tdata[34] );
tran (\cceip_ob_tlv[3][35] , \cceip_ob_tlv[3].tdata[35] );
tran (\cceip_ob_tlv[3][36] , \cceip_ob_tlv[3].tdata[36] );
tran (\cceip_ob_tlv[3][37] , \cceip_ob_tlv[3].tdata[37] );
tran (\cceip_ob_tlv[3][38] , \cceip_ob_tlv[3].tdata[38] );
tran (\cceip_ob_tlv[3][39] , \cceip_ob_tlv[3].tdata[39] );
tran (\cceip_ob_tlv[3][40] , \cceip_ob_tlv[3].tdata[40] );
tran (\cceip_ob_tlv[3][41] , \cceip_ob_tlv[3].tdata[41] );
tran (\cceip_ob_tlv[3][42] , \cceip_ob_tlv[3].tdata[42] );
tran (\cceip_ob_tlv[3][43] , \cceip_ob_tlv[3].tdata[43] );
tran (\cceip_ob_tlv[3][44] , \cceip_ob_tlv[3].tdata[44] );
tran (\cceip_ob_tlv[3][45] , \cceip_ob_tlv[3].tdata[45] );
tran (\cceip_ob_tlv[3][46] , \cceip_ob_tlv[3].tdata[46] );
tran (\cceip_ob_tlv[3][47] , \cceip_ob_tlv[3].tdata[47] );
tran (\cceip_ob_tlv[3][48] , \cceip_ob_tlv[3].tdata[48] );
tran (\cceip_ob_tlv[3][49] , \cceip_ob_tlv[3].tdata[49] );
tran (\cceip_ob_tlv[3][50] , \cceip_ob_tlv[3].tdata[50] );
tran (\cceip_ob_tlv[3][51] , \cceip_ob_tlv[3].tdata[51] );
tran (\cceip_ob_tlv[3][52] , \cceip_ob_tlv[3].tdata[52] );
tran (\cceip_ob_tlv[3][53] , \cceip_ob_tlv[3].tdata[53] );
tran (\cceip_ob_tlv[3][54] , \cceip_ob_tlv[3].tdata[54] );
tran (\cceip_ob_tlv[3][55] , \cceip_ob_tlv[3].tdata[55] );
tran (\cceip_ob_tlv[3][56] , \cceip_ob_tlv[3].tdata[56] );
tran (\cceip_ob_tlv[3][57] , \cceip_ob_tlv[3].tdata[57] );
tran (\cceip_ob_tlv[3][58] , \cceip_ob_tlv[3].tdata[58] );
tran (\cceip_ob_tlv[3][59] , \cceip_ob_tlv[3].tdata[59] );
tran (\cceip_ob_tlv[3][60] , \cceip_ob_tlv[3].tdata[60] );
tran (\cceip_ob_tlv[3][61] , \cceip_ob_tlv[3].tdata[61] );
tran (\cceip_ob_tlv[3][62] , \cceip_ob_tlv[3].tdata[62] );
tran (\cceip_ob_tlv[3][63] , \cceip_ob_tlv[3].tdata[63] );
tran (\cceip_ob_tlv[3][64] , \cceip_ob_tlv[3].tuser[0] );
tran (\cceip_ob_tlv[3][65] , \cceip_ob_tlv[3].tuser[1] );
tran (\cceip_ob_tlv[3][66] , \cceip_ob_tlv[3].tuser[2] );
tran (\cceip_ob_tlv[3][67] , \cceip_ob_tlv[3].tuser[3] );
tran (\cceip_ob_tlv[3][68] , \cceip_ob_tlv[3].tuser[4] );
tran (\cceip_ob_tlv[3][69] , \cceip_ob_tlv[3].tuser[5] );
tran (\cceip_ob_tlv[3][70] , \cceip_ob_tlv[3].tuser[6] );
tran (\cceip_ob_tlv[3][71] , \cceip_ob_tlv[3].tuser[7] );
tran (\cceip_ob_tlv[3][72] , \cceip_ob_tlv[3].tstrb[0] );
tran (\cceip_ob_tlv[3][73] , \cceip_ob_tlv[3].tstrb[1] );
tran (\cceip_ob_tlv[3][74] , \cceip_ob_tlv[3].tstrb[2] );
tran (\cceip_ob_tlv[3][75] , \cceip_ob_tlv[3].tstrb[3] );
tran (\cceip_ob_tlv[3][76] , \cceip_ob_tlv[3].tstrb[4] );
tran (\cceip_ob_tlv[3][77] , \cceip_ob_tlv[3].tstrb[5] );
tran (\cceip_ob_tlv[3][78] , \cceip_ob_tlv[3].tstrb[6] );
tran (\cceip_ob_tlv[3][79] , \cceip_ob_tlv[3].tstrb[7] );
tran (\cceip_ob_tlv[3][80] , \cceip_ob_tlv[3].tid[0] );
tran (\cceip_ob_tlv[3][81] , \cceip_ob_tlv[3].tlast );
tran (\cceip_ob_tlv[3][82] , \cceip_ob_tlv[3].eot );
tran (\cceip_ob_tlv[3][83] , \cceip_ob_tlv[3].sot );
tran (\cceip_ob_tlv[3][84] , \cceip_ob_tlv[3].typen[0] );
tran (\cceip_ob_tlv[3][85] , \cceip_ob_tlv[3].typen[1] );
tran (\cceip_ob_tlv[3][86] , \cceip_ob_tlv[3].typen[2] );
tran (\cceip_ob_tlv[3][87] , \cceip_ob_tlv[3].typen[3] );
tran (\cceip_ob_tlv[3][88] , \cceip_ob_tlv[3].typen[4] );
tran (\cceip_ob_tlv[3][89] , \cceip_ob_tlv[3].typen[5] );
tran (\cceip_ob_tlv[3][90] , \cceip_ob_tlv[3].typen[6] );
tran (\cceip_ob_tlv[3][91] , \cceip_ob_tlv[3].typen[7] );
tran (\cceip_ob_tlv[3][92] , \cceip_ob_tlv[3].ordern[0] );
tran (\cceip_ob_tlv[3][93] , \cceip_ob_tlv[3].ordern[1] );
tran (\cceip_ob_tlv[3][94] , \cceip_ob_tlv[3].ordern[2] );
tran (\cceip_ob_tlv[3][95] , \cceip_ob_tlv[3].ordern[3] );
tran (\cceip_ob_tlv[3][96] , \cceip_ob_tlv[3].ordern[4] );
tran (\cceip_ob_tlv[3][97] , \cceip_ob_tlv[3].ordern[5] );
tran (\cceip_ob_tlv[3][98] , \cceip_ob_tlv[3].ordern[6] );
tran (\cceip_ob_tlv[3][99] , \cceip_ob_tlv[3].ordern[7] );
tran (\cceip_ob_tlv[3][100] , \cceip_ob_tlv[3].ordern[8] );
tran (\cceip_ob_tlv[3][101] , \cceip_ob_tlv[3].ordern[9] );
tran (\cceip_ob_tlv[3][102] , \cceip_ob_tlv[3].ordern[10] );
tran (\cceip_ob_tlv[3][103] , \cceip_ob_tlv[3].ordern[11] );
tran (\cceip_ob_tlv[3][104] , \cceip_ob_tlv[3].ordern[12] );
tran (\cceip_ob_tlv[3][105] , \cceip_ob_tlv[3].insert );
tran (cceip_encrypt_ob_tlv[105], \cceip_encrypt_ob_tlv.insert );
tran (cceip_encrypt_ob_tlv[104], \cceip_encrypt_ob_tlv.ordern [12]);
tran (cceip_encrypt_ob_tlv[103], \cceip_encrypt_ob_tlv.ordern [11]);
tran (cceip_encrypt_ob_tlv[102], \cceip_encrypt_ob_tlv.ordern [10]);
tran (cceip_encrypt_ob_tlv[101], \cceip_encrypt_ob_tlv.ordern [9]);
tran (cceip_encrypt_ob_tlv[100], \cceip_encrypt_ob_tlv.ordern [8]);
tran (cceip_encrypt_ob_tlv[99], \cceip_encrypt_ob_tlv.ordern [7]);
tran (cceip_encrypt_ob_tlv[98], \cceip_encrypt_ob_tlv.ordern [6]);
tran (cceip_encrypt_ob_tlv[97], \cceip_encrypt_ob_tlv.ordern [5]);
tran (cceip_encrypt_ob_tlv[96], \cceip_encrypt_ob_tlv.ordern [4]);
tran (cceip_encrypt_ob_tlv[95], \cceip_encrypt_ob_tlv.ordern [3]);
tran (cceip_encrypt_ob_tlv[94], \cceip_encrypt_ob_tlv.ordern [2]);
tran (cceip_encrypt_ob_tlv[93], \cceip_encrypt_ob_tlv.ordern [1]);
tran (cceip_encrypt_ob_tlv[92], \cceip_encrypt_ob_tlv.ordern [0]);
tran (cceip_encrypt_ob_tlv[91], \cceip_encrypt_ob_tlv.typen [7]);
tran (cceip_encrypt_ob_tlv[90], \cceip_encrypt_ob_tlv.typen [6]);
tran (cceip_encrypt_ob_tlv[89], \cceip_encrypt_ob_tlv.typen [5]);
tran (cceip_encrypt_ob_tlv[88], \cceip_encrypt_ob_tlv.typen [4]);
tran (cceip_encrypt_ob_tlv[87], \cceip_encrypt_ob_tlv.typen [3]);
tran (cceip_encrypt_ob_tlv[86], \cceip_encrypt_ob_tlv.typen [2]);
tran (cceip_encrypt_ob_tlv[85], \cceip_encrypt_ob_tlv.typen [1]);
tran (cceip_encrypt_ob_tlv[84], \cceip_encrypt_ob_tlv.typen [0]);
tran (cceip_encrypt_ob_tlv[83], \cceip_encrypt_ob_tlv.sot );
tran (cceip_encrypt_ob_tlv[82], \cceip_encrypt_ob_tlv.eot );
tran (cceip_encrypt_ob_tlv[81], \cceip_encrypt_ob_tlv.tlast );
tran (cceip_encrypt_ob_tlv[80], \cceip_encrypt_ob_tlv.tid [0]);
tran (cceip_encrypt_ob_tlv[79], \cceip_encrypt_ob_tlv.tstrb [7]);
tran (cceip_encrypt_ob_tlv[78], \cceip_encrypt_ob_tlv.tstrb [6]);
tran (cceip_encrypt_ob_tlv[77], \cceip_encrypt_ob_tlv.tstrb [5]);
tran (cceip_encrypt_ob_tlv[76], \cceip_encrypt_ob_tlv.tstrb [4]);
tran (cceip_encrypt_ob_tlv[75], \cceip_encrypt_ob_tlv.tstrb [3]);
tran (cceip_encrypt_ob_tlv[74], \cceip_encrypt_ob_tlv.tstrb [2]);
tran (cceip_encrypt_ob_tlv[73], \cceip_encrypt_ob_tlv.tstrb [1]);
tran (cceip_encrypt_ob_tlv[72], \cceip_encrypt_ob_tlv.tstrb [0]);
tran (cceip_encrypt_ob_tlv[71], \cceip_encrypt_ob_tlv.tuser [7]);
tran (cceip_encrypt_ob_tlv[70], \cceip_encrypt_ob_tlv.tuser [6]);
tran (cceip_encrypt_ob_tlv[69], \cceip_encrypt_ob_tlv.tuser [5]);
tran (cceip_encrypt_ob_tlv[68], \cceip_encrypt_ob_tlv.tuser [4]);
tran (cceip_encrypt_ob_tlv[67], \cceip_encrypt_ob_tlv.tuser [3]);
tran (cceip_encrypt_ob_tlv[66], \cceip_encrypt_ob_tlv.tuser [2]);
tran (cceip_encrypt_ob_tlv[65], \cceip_encrypt_ob_tlv.tuser [1]);
tran (cceip_encrypt_ob_tlv[64], \cceip_encrypt_ob_tlv.tuser [0]);
tran (cceip_encrypt_ob_tlv[63], \cceip_encrypt_ob_tlv.tdata [63]);
tran (cceip_encrypt_ob_tlv[62], \cceip_encrypt_ob_tlv.tdata [62]);
tran (cceip_encrypt_ob_tlv[61], \cceip_encrypt_ob_tlv.tdata [61]);
tran (cceip_encrypt_ob_tlv[60], \cceip_encrypt_ob_tlv.tdata [60]);
tran (cceip_encrypt_ob_tlv[59], \cceip_encrypt_ob_tlv.tdata [59]);
tran (cceip_encrypt_ob_tlv[58], \cceip_encrypt_ob_tlv.tdata [58]);
tran (cceip_encrypt_ob_tlv[57], \cceip_encrypt_ob_tlv.tdata [57]);
tran (cceip_encrypt_ob_tlv[56], \cceip_encrypt_ob_tlv.tdata [56]);
tran (cceip_encrypt_ob_tlv[55], \cceip_encrypt_ob_tlv.tdata [55]);
tran (cceip_encrypt_ob_tlv[54], \cceip_encrypt_ob_tlv.tdata [54]);
tran (cceip_encrypt_ob_tlv[53], \cceip_encrypt_ob_tlv.tdata [53]);
tran (cceip_encrypt_ob_tlv[52], \cceip_encrypt_ob_tlv.tdata [52]);
tran (cceip_encrypt_ob_tlv[51], \cceip_encrypt_ob_tlv.tdata [51]);
tran (cceip_encrypt_ob_tlv[50], \cceip_encrypt_ob_tlv.tdata [50]);
tran (cceip_encrypt_ob_tlv[49], \cceip_encrypt_ob_tlv.tdata [49]);
tran (cceip_encrypt_ob_tlv[48], \cceip_encrypt_ob_tlv.tdata [48]);
tran (cceip_encrypt_ob_tlv[47], \cceip_encrypt_ob_tlv.tdata [47]);
tran (cceip_encrypt_ob_tlv[46], \cceip_encrypt_ob_tlv.tdata [46]);
tran (cceip_encrypt_ob_tlv[45], \cceip_encrypt_ob_tlv.tdata [45]);
tran (cceip_encrypt_ob_tlv[44], \cceip_encrypt_ob_tlv.tdata [44]);
tran (cceip_encrypt_ob_tlv[43], \cceip_encrypt_ob_tlv.tdata [43]);
tran (cceip_encrypt_ob_tlv[42], \cceip_encrypt_ob_tlv.tdata [42]);
tran (cceip_encrypt_ob_tlv[41], \cceip_encrypt_ob_tlv.tdata [41]);
tran (cceip_encrypt_ob_tlv[40], \cceip_encrypt_ob_tlv.tdata [40]);
tran (cceip_encrypt_ob_tlv[39], \cceip_encrypt_ob_tlv.tdata [39]);
tran (cceip_encrypt_ob_tlv[38], \cceip_encrypt_ob_tlv.tdata [38]);
tran (cceip_encrypt_ob_tlv[37], \cceip_encrypt_ob_tlv.tdata [37]);
tran (cceip_encrypt_ob_tlv[36], \cceip_encrypt_ob_tlv.tdata [36]);
tran (cceip_encrypt_ob_tlv[35], \cceip_encrypt_ob_tlv.tdata [35]);
tran (cceip_encrypt_ob_tlv[34], \cceip_encrypt_ob_tlv.tdata [34]);
tran (cceip_encrypt_ob_tlv[33], \cceip_encrypt_ob_tlv.tdata [33]);
tran (cceip_encrypt_ob_tlv[32], \cceip_encrypt_ob_tlv.tdata [32]);
tran (cceip_encrypt_ob_tlv[31], \cceip_encrypt_ob_tlv.tdata [31]);
tran (cceip_encrypt_ob_tlv[30], \cceip_encrypt_ob_tlv.tdata [30]);
tran (cceip_encrypt_ob_tlv[29], \cceip_encrypt_ob_tlv.tdata [29]);
tran (cceip_encrypt_ob_tlv[28], \cceip_encrypt_ob_tlv.tdata [28]);
tran (cceip_encrypt_ob_tlv[27], \cceip_encrypt_ob_tlv.tdata [27]);
tran (cceip_encrypt_ob_tlv[26], \cceip_encrypt_ob_tlv.tdata [26]);
tran (cceip_encrypt_ob_tlv[25], \cceip_encrypt_ob_tlv.tdata [25]);
tran (cceip_encrypt_ob_tlv[24], \cceip_encrypt_ob_tlv.tdata [24]);
tran (cceip_encrypt_ob_tlv[23], \cceip_encrypt_ob_tlv.tdata [23]);
tran (cceip_encrypt_ob_tlv[22], \cceip_encrypt_ob_tlv.tdata [22]);
tran (cceip_encrypt_ob_tlv[21], \cceip_encrypt_ob_tlv.tdata [21]);
tran (cceip_encrypt_ob_tlv[20], \cceip_encrypt_ob_tlv.tdata [20]);
tran (cceip_encrypt_ob_tlv[19], \cceip_encrypt_ob_tlv.tdata [19]);
tran (cceip_encrypt_ob_tlv[18], \cceip_encrypt_ob_tlv.tdata [18]);
tran (cceip_encrypt_ob_tlv[17], \cceip_encrypt_ob_tlv.tdata [17]);
tran (cceip_encrypt_ob_tlv[16], \cceip_encrypt_ob_tlv.tdata [16]);
tran (cceip_encrypt_ob_tlv[15], \cceip_encrypt_ob_tlv.tdata [15]);
tran (cceip_encrypt_ob_tlv[14], \cceip_encrypt_ob_tlv.tdata [14]);
tran (cceip_encrypt_ob_tlv[13], \cceip_encrypt_ob_tlv.tdata [13]);
tran (cceip_encrypt_ob_tlv[12], \cceip_encrypt_ob_tlv.tdata [12]);
tran (cceip_encrypt_ob_tlv[11], \cceip_encrypt_ob_tlv.tdata [11]);
tran (cceip_encrypt_ob_tlv[10], \cceip_encrypt_ob_tlv.tdata [10]);
tran (cceip_encrypt_ob_tlv[9], \cceip_encrypt_ob_tlv.tdata [9]);
tran (cceip_encrypt_ob_tlv[8], \cceip_encrypt_ob_tlv.tdata [8]);
tran (cceip_encrypt_ob_tlv[7], \cceip_encrypt_ob_tlv.tdata [7]);
tran (cceip_encrypt_ob_tlv[6], \cceip_encrypt_ob_tlv.tdata [6]);
tran (cceip_encrypt_ob_tlv[5], \cceip_encrypt_ob_tlv.tdata [5]);
tran (cceip_encrypt_ob_tlv[4], \cceip_encrypt_ob_tlv.tdata [4]);
tran (cceip_encrypt_ob_tlv[3], \cceip_encrypt_ob_tlv.tdata [3]);
tran (cceip_encrypt_ob_tlv[2], \cceip_encrypt_ob_tlv.tdata [2]);
tran (cceip_encrypt_ob_tlv[1], \cceip_encrypt_ob_tlv.tdata [1]);
tran (cceip_encrypt_ob_tlv[0], \cceip_encrypt_ob_tlv.tdata [0]);
tran (cceip_validate_ob_tlv[105], \cceip_validate_ob_tlv.insert );
tran (cceip_validate_ob_tlv[104], \cceip_validate_ob_tlv.ordern [12]);
tran (cceip_validate_ob_tlv[103], \cceip_validate_ob_tlv.ordern [11]);
tran (cceip_validate_ob_tlv[102], \cceip_validate_ob_tlv.ordern [10]);
tran (cceip_validate_ob_tlv[101], \cceip_validate_ob_tlv.ordern [9]);
tran (cceip_validate_ob_tlv[100], \cceip_validate_ob_tlv.ordern [8]);
tran (cceip_validate_ob_tlv[99], \cceip_validate_ob_tlv.ordern [7]);
tran (cceip_validate_ob_tlv[98], \cceip_validate_ob_tlv.ordern [6]);
tran (cceip_validate_ob_tlv[97], \cceip_validate_ob_tlv.ordern [5]);
tran (cceip_validate_ob_tlv[96], \cceip_validate_ob_tlv.ordern [4]);
tran (cceip_validate_ob_tlv[95], \cceip_validate_ob_tlv.ordern [3]);
tran (cceip_validate_ob_tlv[94], \cceip_validate_ob_tlv.ordern [2]);
tran (cceip_validate_ob_tlv[93], \cceip_validate_ob_tlv.ordern [1]);
tran (cceip_validate_ob_tlv[92], \cceip_validate_ob_tlv.ordern [0]);
tran (cceip_validate_ob_tlv[91], \cceip_validate_ob_tlv.typen [7]);
tran (cceip_validate_ob_tlv[90], \cceip_validate_ob_tlv.typen [6]);
tran (cceip_validate_ob_tlv[89], \cceip_validate_ob_tlv.typen [5]);
tran (cceip_validate_ob_tlv[88], \cceip_validate_ob_tlv.typen [4]);
tran (cceip_validate_ob_tlv[87], \cceip_validate_ob_tlv.typen [3]);
tran (cceip_validate_ob_tlv[86], \cceip_validate_ob_tlv.typen [2]);
tran (cceip_validate_ob_tlv[85], \cceip_validate_ob_tlv.typen [1]);
tran (cceip_validate_ob_tlv[84], \cceip_validate_ob_tlv.typen [0]);
tran (cceip_validate_ob_tlv[83], \cceip_validate_ob_tlv.sot );
tran (cceip_validate_ob_tlv[82], \cceip_validate_ob_tlv.eot );
tran (cceip_validate_ob_tlv[81], \cceip_validate_ob_tlv.tlast );
tran (cceip_validate_ob_tlv[80], \cceip_validate_ob_tlv.tid [0]);
tran (cceip_validate_ob_tlv[79], \cceip_validate_ob_tlv.tstrb [7]);
tran (cceip_validate_ob_tlv[78], \cceip_validate_ob_tlv.tstrb [6]);
tran (cceip_validate_ob_tlv[77], \cceip_validate_ob_tlv.tstrb [5]);
tran (cceip_validate_ob_tlv[76], \cceip_validate_ob_tlv.tstrb [4]);
tran (cceip_validate_ob_tlv[75], \cceip_validate_ob_tlv.tstrb [3]);
tran (cceip_validate_ob_tlv[74], \cceip_validate_ob_tlv.tstrb [2]);
tran (cceip_validate_ob_tlv[73], \cceip_validate_ob_tlv.tstrb [1]);
tran (cceip_validate_ob_tlv[72], \cceip_validate_ob_tlv.tstrb [0]);
tran (cceip_validate_ob_tlv[71], \cceip_validate_ob_tlv.tuser [7]);
tran (cceip_validate_ob_tlv[70], \cceip_validate_ob_tlv.tuser [6]);
tran (cceip_validate_ob_tlv[69], \cceip_validate_ob_tlv.tuser [5]);
tran (cceip_validate_ob_tlv[68], \cceip_validate_ob_tlv.tuser [4]);
tran (cceip_validate_ob_tlv[67], \cceip_validate_ob_tlv.tuser [3]);
tran (cceip_validate_ob_tlv[66], \cceip_validate_ob_tlv.tuser [2]);
tran (cceip_validate_ob_tlv[65], \cceip_validate_ob_tlv.tuser [1]);
tran (cceip_validate_ob_tlv[64], \cceip_validate_ob_tlv.tuser [0]);
tran (cceip_validate_ob_tlv[63], \cceip_validate_ob_tlv.tdata [63]);
tran (cceip_validate_ob_tlv[62], \cceip_validate_ob_tlv.tdata [62]);
tran (cceip_validate_ob_tlv[61], \cceip_validate_ob_tlv.tdata [61]);
tran (cceip_validate_ob_tlv[60], \cceip_validate_ob_tlv.tdata [60]);
tran (cceip_validate_ob_tlv[59], \cceip_validate_ob_tlv.tdata [59]);
tran (cceip_validate_ob_tlv[58], \cceip_validate_ob_tlv.tdata [58]);
tran (cceip_validate_ob_tlv[57], \cceip_validate_ob_tlv.tdata [57]);
tran (cceip_validate_ob_tlv[56], \cceip_validate_ob_tlv.tdata [56]);
tran (cceip_validate_ob_tlv[55], \cceip_validate_ob_tlv.tdata [55]);
tran (cceip_validate_ob_tlv[54], \cceip_validate_ob_tlv.tdata [54]);
tran (cceip_validate_ob_tlv[53], \cceip_validate_ob_tlv.tdata [53]);
tran (cceip_validate_ob_tlv[52], \cceip_validate_ob_tlv.tdata [52]);
tran (cceip_validate_ob_tlv[51], \cceip_validate_ob_tlv.tdata [51]);
tran (cceip_validate_ob_tlv[50], \cceip_validate_ob_tlv.tdata [50]);
tran (cceip_validate_ob_tlv[49], \cceip_validate_ob_tlv.tdata [49]);
tran (cceip_validate_ob_tlv[48], \cceip_validate_ob_tlv.tdata [48]);
tran (cceip_validate_ob_tlv[47], \cceip_validate_ob_tlv.tdata [47]);
tran (cceip_validate_ob_tlv[46], \cceip_validate_ob_tlv.tdata [46]);
tran (cceip_validate_ob_tlv[45], \cceip_validate_ob_tlv.tdata [45]);
tran (cceip_validate_ob_tlv[44], \cceip_validate_ob_tlv.tdata [44]);
tran (cceip_validate_ob_tlv[43], \cceip_validate_ob_tlv.tdata [43]);
tran (cceip_validate_ob_tlv[42], \cceip_validate_ob_tlv.tdata [42]);
tran (cceip_validate_ob_tlv[41], \cceip_validate_ob_tlv.tdata [41]);
tran (cceip_validate_ob_tlv[40], \cceip_validate_ob_tlv.tdata [40]);
tran (cceip_validate_ob_tlv[39], \cceip_validate_ob_tlv.tdata [39]);
tran (cceip_validate_ob_tlv[38], \cceip_validate_ob_tlv.tdata [38]);
tran (cceip_validate_ob_tlv[37], \cceip_validate_ob_tlv.tdata [37]);
tran (cceip_validate_ob_tlv[36], \cceip_validate_ob_tlv.tdata [36]);
tran (cceip_validate_ob_tlv[35], \cceip_validate_ob_tlv.tdata [35]);
tran (cceip_validate_ob_tlv[34], \cceip_validate_ob_tlv.tdata [34]);
tran (cceip_validate_ob_tlv[33], \cceip_validate_ob_tlv.tdata [33]);
tran (cceip_validate_ob_tlv[32], \cceip_validate_ob_tlv.tdata [32]);
tran (cceip_validate_ob_tlv[31], \cceip_validate_ob_tlv.tdata [31]);
tran (cceip_validate_ob_tlv[30], \cceip_validate_ob_tlv.tdata [30]);
tran (cceip_validate_ob_tlv[29], \cceip_validate_ob_tlv.tdata [29]);
tran (cceip_validate_ob_tlv[28], \cceip_validate_ob_tlv.tdata [28]);
tran (cceip_validate_ob_tlv[27], \cceip_validate_ob_tlv.tdata [27]);
tran (cceip_validate_ob_tlv[26], \cceip_validate_ob_tlv.tdata [26]);
tran (cceip_validate_ob_tlv[25], \cceip_validate_ob_tlv.tdata [25]);
tran (cceip_validate_ob_tlv[24], \cceip_validate_ob_tlv.tdata [24]);
tran (cceip_validate_ob_tlv[23], \cceip_validate_ob_tlv.tdata [23]);
tran (cceip_validate_ob_tlv[22], \cceip_validate_ob_tlv.tdata [22]);
tran (cceip_validate_ob_tlv[21], \cceip_validate_ob_tlv.tdata [21]);
tran (cceip_validate_ob_tlv[20], \cceip_validate_ob_tlv.tdata [20]);
tran (cceip_validate_ob_tlv[19], \cceip_validate_ob_tlv.tdata [19]);
tran (cceip_validate_ob_tlv[18], \cceip_validate_ob_tlv.tdata [18]);
tran (cceip_validate_ob_tlv[17], \cceip_validate_ob_tlv.tdata [17]);
tran (cceip_validate_ob_tlv[16], \cceip_validate_ob_tlv.tdata [16]);
tran (cceip_validate_ob_tlv[15], \cceip_validate_ob_tlv.tdata [15]);
tran (cceip_validate_ob_tlv[14], \cceip_validate_ob_tlv.tdata [14]);
tran (cceip_validate_ob_tlv[13], \cceip_validate_ob_tlv.tdata [13]);
tran (cceip_validate_ob_tlv[12], \cceip_validate_ob_tlv.tdata [12]);
tran (cceip_validate_ob_tlv[11], \cceip_validate_ob_tlv.tdata [11]);
tran (cceip_validate_ob_tlv[10], \cceip_validate_ob_tlv.tdata [10]);
tran (cceip_validate_ob_tlv[9], \cceip_validate_ob_tlv.tdata [9]);
tran (cceip_validate_ob_tlv[8], \cceip_validate_ob_tlv.tdata [8]);
tran (cceip_validate_ob_tlv[7], \cceip_validate_ob_tlv.tdata [7]);
tran (cceip_validate_ob_tlv[6], \cceip_validate_ob_tlv.tdata [6]);
tran (cceip_validate_ob_tlv[5], \cceip_validate_ob_tlv.tdata [5]);
tran (cceip_validate_ob_tlv[4], \cceip_validate_ob_tlv.tdata [4]);
tran (cceip_validate_ob_tlv[3], \cceip_validate_ob_tlv.tdata [3]);
tran (cceip_validate_ob_tlv[2], \cceip_validate_ob_tlv.tdata [2]);
tran (cceip_validate_ob_tlv[1], \cceip_validate_ob_tlv.tdata [1]);
tran (cceip_validate_ob_tlv[0], \cceip_validate_ob_tlv.tdata [0]);
tran (key_tlv_w0[0], \key_tlv_w0.tlv_type [0]);
tran (key_tlv_w0[1], \key_tlv_w0.tlv_type [1]);
tran (key_tlv_w0[2], \key_tlv_w0.tlv_type [2]);
tran (key_tlv_w0[3], \key_tlv_w0.tlv_type [3]);
tran (key_tlv_w0[4], \key_tlv_w0.tlv_type [4]);
tran (key_tlv_w0[5], \key_tlv_w0.tlv_type [5]);
tran (key_tlv_w0[6], \key_tlv_w0.tlv_type [6]);
tran (key_tlv_w0[7], \key_tlv_w0.tlv_type [7]);
tran (key_tlv_w0[8], \key_tlv_w0.tlv_len [0]);
tran (key_tlv_w0[9], \key_tlv_w0.tlv_len [1]);
tran (key_tlv_w0[10], \key_tlv_w0.tlv_len [2]);
tran (key_tlv_w0[11], \key_tlv_w0.tlv_len [3]);
tran (key_tlv_w0[12], \key_tlv_w0.tlv_len [4]);
tran (key_tlv_w0[13], \key_tlv_w0.tlv_len [5]);
tran (key_tlv_w0[14], \key_tlv_w0.tlv_len [6]);
tran (key_tlv_w0[15], \key_tlv_w0.tlv_len [7]);
tran (key_tlv_w0[16], \key_tlv_w0.tlv_seq_num [0]);
tran (key_tlv_w0[17], \key_tlv_w0.tlv_seq_num [1]);
tran (key_tlv_w0[18], \key_tlv_w0.tlv_seq_num [2]);
tran (key_tlv_w0[19], \key_tlv_w0.tlv_seq_num [3]);
tran (key_tlv_w0[20], \key_tlv_w0.tlv_seq_num [4]);
tran (key_tlv_w0[21], \key_tlv_w0.tlv_seq_num [5]);
tran (key_tlv_w0[22], \key_tlv_w0.tlv_seq_num [6]);
tran (key_tlv_w0[23], \key_tlv_w0.tlv_seq_num [7]);
tran (key_tlv_w0[24], \key_tlv_w0.tlv_eng_id [0]);
tran (key_tlv_w0[25], \key_tlv_w0.tlv_eng_id [1]);
tran (key_tlv_w0[26], \key_tlv_w0.tlv_eng_id [2]);
tran (key_tlv_w0[27], \key_tlv_w0.tlv_eng_id [3]);
tran (key_tlv_w0[28], \key_tlv_w0.resv1 [0]);
tran (key_tlv_w0[29], \key_tlv_w0.resv1 [1]);
tran (key_tlv_w0[30], \key_tlv_w0.resv1 [2]);
tran (key_tlv_w0[31], \key_tlv_w0.resv1 [3]);
tran (key_tlv_w0[32], \key_tlv_w0.tlv_frame_num [0]);
tran (key_tlv_w0[33], \key_tlv_w0.tlv_frame_num [1]);
tran (key_tlv_w0[34], \key_tlv_w0.tlv_frame_num [2]);
tran (key_tlv_w0[35], \key_tlv_w0.tlv_frame_num [3]);
tran (key_tlv_w0[36], \key_tlv_w0.tlv_frame_num [4]);
tran (key_tlv_w0[37], \key_tlv_w0.tlv_frame_num [5]);
tran (key_tlv_w0[38], \key_tlv_w0.tlv_frame_num [6]);
tran (key_tlv_w0[39], \key_tlv_w0.tlv_frame_num [7]);
tran (key_tlv_w0[40], \key_tlv_w0.tlv_frame_num [8]);
tran (key_tlv_w0[41], \key_tlv_w0.tlv_frame_num [9]);
tran (key_tlv_w0[42], \key_tlv_w0.tlv_frame_num [10]);
tran (key_tlv_w0[43], \key_tlv_w0.resv0 [0]);
tran (key_tlv_w0[44], \key_tlv_w0.resv0 [1]);
tran (key_tlv_w0[45], \key_tlv_w0.resv0 [2]);
tran (key_tlv_w0[46], \key_tlv_w0.resv0 [3]);
tran (key_tlv_w0[47], \key_tlv_w0.resv0 [4]);
tran (key_tlv_w0[48], \key_tlv_w0.resv0 [5]);
tran (key_tlv_w0[49], \key_tlv_w0.resv0 [6]);
tran (key_tlv_w0[50], \key_tlv_w0.resv0 [7]);
tran (key_tlv_w0[51], \key_tlv_w0.resv0 [8]);
tran (key_tlv_w0[52], \key_tlv_w0.resv0 [9]);
tran (key_tlv_w0[53], \key_tlv_w0.resv0 [10]);
tran (key_tlv_w0[54], \key_tlv_w0.resv0 [11]);
tran (key_tlv_w0[55], \key_tlv_w0.resv0 [12]);
tran (key_tlv_w0[56], \key_tlv_w0.resv0 [13]);
tran (key_tlv_w0[57], \key_tlv_w0.resv0 [14]);
tran (key_tlv_w0[58], \key_tlv_w0.resv0 [15]);
tran (key_tlv_w0[59], \key_tlv_w0.resv0 [16]);
tran (key_tlv_w0[60], \key_tlv_w0.resv0 [17]);
tran (key_tlv_w0[61], \key_tlv_w0.resv0 [18]);
tran (key_tlv_w0[62], \key_tlv_w0.tlv_bip2 [0]);
tran (key_tlv_w0[63], \key_tlv_w0.tlv_bip2 [1]);
tran (encrypt_out[105], \encrypt_out.insert );
tran (encrypt_out[104], \encrypt_out.ordern [12]);
tran (encrypt_out[103], \encrypt_out.ordern [11]);
tran (encrypt_out[102], \encrypt_out.ordern [10]);
tran (encrypt_out[101], \encrypt_out.ordern [9]);
tran (encrypt_out[100], \encrypt_out.ordern [8]);
tran (encrypt_out[99], \encrypt_out.ordern [7]);
tran (encrypt_out[98], \encrypt_out.ordern [6]);
tran (encrypt_out[97], \encrypt_out.ordern [5]);
tran (encrypt_out[96], \encrypt_out.ordern [4]);
tran (encrypt_out[95], \encrypt_out.ordern [3]);
tran (encrypt_out[94], \encrypt_out.ordern [2]);
tran (encrypt_out[93], \encrypt_out.ordern [1]);
tran (encrypt_out[92], \encrypt_out.ordern [0]);
tran (encrypt_out[91], \encrypt_out.typen [7]);
tran (encrypt_out[90], \encrypt_out.typen [6]);
tran (encrypt_out[89], \encrypt_out.typen [5]);
tran (encrypt_out[88], \encrypt_out.typen [4]);
tran (encrypt_out[87], \encrypt_out.typen [3]);
tran (encrypt_out[86], \encrypt_out.typen [2]);
tran (encrypt_out[85], \encrypt_out.typen [1]);
tran (encrypt_out[84], \encrypt_out.typen [0]);
tran (encrypt_out[83], \encrypt_out.sot );
tran (encrypt_out[82], \encrypt_out.eot );
tran (encrypt_out[81], \encrypt_out.tlast );
tran (encrypt_out[80], \encrypt_out.tid [0]);
tran (encrypt_out[79], \encrypt_out.tstrb [7]);
tran (encrypt_out[78], \encrypt_out.tstrb [6]);
tran (encrypt_out[77], \encrypt_out.tstrb [5]);
tran (encrypt_out[76], \encrypt_out.tstrb [4]);
tran (encrypt_out[75], \encrypt_out.tstrb [3]);
tran (encrypt_out[74], \encrypt_out.tstrb [2]);
tran (encrypt_out[73], \encrypt_out.tstrb [1]);
tran (encrypt_out[72], \encrypt_out.tstrb [0]);
tran (encrypt_out[71], \encrypt_out.tuser [7]);
tran (encrypt_out[70], \encrypt_out.tuser [6]);
tran (encrypt_out[69], \encrypt_out.tuser [5]);
tran (encrypt_out[68], \encrypt_out.tuser [4]);
tran (encrypt_out[67], \encrypt_out.tuser [3]);
tran (encrypt_out[66], \encrypt_out.tuser [2]);
tran (encrypt_out[65], \encrypt_out.tuser [1]);
tran (encrypt_out[64], \encrypt_out.tuser [0]);
tran (validate_out[105], \validate_out.insert );
tran (validate_out[104], \validate_out.ordern [12]);
tran (validate_out[103], \validate_out.ordern [11]);
tran (validate_out[102], \validate_out.ordern [10]);
tran (validate_out[101], \validate_out.ordern [9]);
tran (validate_out[100], \validate_out.ordern [8]);
tran (validate_out[99], \validate_out.ordern [7]);
tran (validate_out[98], \validate_out.ordern [6]);
tran (validate_out[97], \validate_out.ordern [5]);
tran (validate_out[96], \validate_out.ordern [4]);
tran (validate_out[95], \validate_out.ordern [3]);
tran (validate_out[94], \validate_out.ordern [2]);
tran (validate_out[93], \validate_out.ordern [1]);
tran (validate_out[92], \validate_out.ordern [0]);
tran (validate_out[91], \validate_out.typen [7]);
tran (validate_out[90], \validate_out.typen [6]);
tran (validate_out[89], \validate_out.typen [5]);
tran (validate_out[88], \validate_out.typen [4]);
tran (validate_out[87], \validate_out.typen [3]);
tran (validate_out[86], \validate_out.typen [2]);
tran (validate_out[85], \validate_out.typen [1]);
tran (validate_out[84], \validate_out.typen [0]);
tran (validate_out[83], \validate_out.sot );
tran (validate_out[82], \validate_out.eot );
tran (validate_out[81], \validate_out.tlast );
tran (validate_out[80], \validate_out.tid [0]);
tran (validate_out[79], \validate_out.tstrb [7]);
tran (validate_out[78], \validate_out.tstrb [6]);
tran (validate_out[77], \validate_out.tstrb [5]);
tran (validate_out[76], \validate_out.tstrb [4]);
tran (validate_out[75], \validate_out.tstrb [3]);
tran (validate_out[74], \validate_out.tstrb [2]);
tran (validate_out[73], \validate_out.tstrb [1]);
tran (validate_out[72], \validate_out.tstrb [0]);
tran (validate_out[71], \validate_out.tuser [7]);
tran (validate_out[70], \validate_out.tuser [6]);
tran (validate_out[69], \validate_out.tuser [5]);
tran (validate_out[68], \validate_out.tuser [4]);
tran (validate_out[67], \validate_out.tuser [3]);
tran (validate_out[66], \validate_out.tuser [2]);
tran (validate_out[65], \validate_out.tuser [1]);
tran (validate_out[64], \validate_out.tuser [0]);
tran (validate_out[63], \validate_out.tdata [63]);
tran (validate_out[62], \validate_out.tdata [62]);
tran (validate_out[61], \validate_out.tdata [61]);
tran (validate_out[60], \validate_out.tdata [60]);
tran (validate_out[59], \validate_out.tdata [59]);
tran (validate_out[58], \validate_out.tdata [58]);
tran (validate_out[57], \validate_out.tdata [57]);
tran (validate_out[56], \validate_out.tdata [56]);
tran (validate_out[55], \validate_out.tdata [55]);
tran (validate_out[54], \validate_out.tdata [54]);
tran (validate_out[53], \validate_out.tdata [53]);
tran (validate_out[52], \validate_out.tdata [52]);
tran (validate_out[51], \validate_out.tdata [51]);
tran (validate_out[50], \validate_out.tdata [50]);
tran (validate_out[49], \validate_out.tdata [49]);
tran (validate_out[48], \validate_out.tdata [48]);
tran (validate_out[47], \validate_out.tdata [47]);
tran (validate_out[46], \validate_out.tdata [46]);
tran (validate_out[45], \validate_out.tdata [45]);
tran (validate_out[44], \validate_out.tdata [44]);
tran (validate_out[43], \validate_out.tdata [43]);
tran (validate_out[42], \validate_out.tdata [42]);
tran (validate_out[41], \validate_out.tdata [41]);
tran (validate_out[40], \validate_out.tdata [40]);
tran (validate_out[39], \validate_out.tdata [39]);
tran (validate_out[38], \validate_out.tdata [38]);
tran (validate_out[37], \validate_out.tdata [37]);
tran (validate_out[36], \validate_out.tdata [36]);
tran (validate_out[35], \validate_out.tdata [35]);
tran (validate_out[34], \validate_out.tdata [34]);
tran (validate_out[33], \validate_out.tdata [33]);
tran (validate_out[32], \validate_out.tdata [32]);
tran (validate_out[31], \validate_out.tdata [31]);
tran (validate_out[30], \validate_out.tdata [30]);
tran (validate_out[29], \validate_out.tdata [29]);
tran (validate_out[28], \validate_out.tdata [28]);
tran (validate_out[27], \validate_out.tdata [27]);
tran (validate_out[26], \validate_out.tdata [26]);
tran (validate_out[25], \validate_out.tdata [25]);
tran (validate_out[24], \validate_out.tdata [24]);
tran (validate_out[23], \validate_out.tdata [23]);
tran (validate_out[22], \validate_out.tdata [22]);
tran (validate_out[21], \validate_out.tdata [21]);
tran (validate_out[20], \validate_out.tdata [20]);
tran (validate_out[19], \validate_out.tdata [19]);
tran (validate_out[18], \validate_out.tdata [18]);
tran (validate_out[17], \validate_out.tdata [17]);
tran (validate_out[16], \validate_out.tdata [16]);
tran (validate_out[15], \validate_out.tdata [15]);
tran (validate_out[14], \validate_out.tdata [14]);
tran (validate_out[13], \validate_out.tdata [13]);
tran (validate_out[12], \validate_out.tdata [12]);
tran (validate_out[11], \validate_out.tdata [11]);
tran (validate_out[10], \validate_out.tdata [10]);
tran (validate_out[9], \validate_out.tdata [9]);
tran (validate_out[8], \validate_out.tdata [8]);
tran (validate_out[7], \validate_out.tdata [7]);
tran (validate_out[6], \validate_out.tdata [6]);
tran (validate_out[5], \validate_out.tdata [5]);
tran (validate_out[4], \validate_out.tdata [4]);
tran (validate_out[3], \validate_out.tdata [3]);
tran (validate_out[2], \validate_out.tdata [2]);
tran (validate_out[1], \validate_out.tdata [1]);
tran (validate_out[0], \validate_out.tdata [0]);
tran (encrypt_out[63], \encrypt_out.tdata [63]);
tran (encrypt_out[62], \encrypt_out.tdata [62]);
tran (encrypt_out[61], \encrypt_out.tdata [61]);
tran (encrypt_out[60], \encrypt_out.tdata [60]);
tran (encrypt_out[59], \encrypt_out.tdata [59]);
tran (encrypt_out[58], \encrypt_out.tdata [58]);
tran (encrypt_out[57], \encrypt_out.tdata [57]);
tran (encrypt_out[56], \encrypt_out.tdata [56]);
tran (encrypt_out[55], \encrypt_out.tdata [55]);
tran (encrypt_out[54], \encrypt_out.tdata [54]);
tran (encrypt_out[53], \encrypt_out.tdata [53]);
tran (encrypt_out[52], \encrypt_out.tdata [52]);
tran (encrypt_out[51], \encrypt_out.tdata [51]);
tran (encrypt_out[50], \encrypt_out.tdata [50]);
tran (encrypt_out[49], \encrypt_out.tdata [49]);
tran (encrypt_out[48], \encrypt_out.tdata [48]);
tran (encrypt_out[47], \encrypt_out.tdata [47]);
tran (encrypt_out[46], \encrypt_out.tdata [46]);
tran (encrypt_out[45], \encrypt_out.tdata [45]);
tran (encrypt_out[44], \encrypt_out.tdata [44]);
tran (encrypt_out[43], \encrypt_out.tdata [43]);
tran (encrypt_out[42], \encrypt_out.tdata [42]);
tran (encrypt_out[41], \encrypt_out.tdata [41]);
tran (encrypt_out[40], \encrypt_out.tdata [40]);
tran (encrypt_out[39], \encrypt_out.tdata [39]);
tran (encrypt_out[38], \encrypt_out.tdata [38]);
tran (encrypt_out[37], \encrypt_out.tdata [37]);
tran (encrypt_out[36], \encrypt_out.tdata [36]);
tran (encrypt_out[35], \encrypt_out.tdata [35]);
tran (encrypt_out[34], \encrypt_out.tdata [34]);
tran (encrypt_out[33], \encrypt_out.tdata [33]);
tran (encrypt_out[32], \encrypt_out.tdata [32]);
tran (encrypt_out[31], \encrypt_out.tdata [31]);
tran (encrypt_out[30], \encrypt_out.tdata [30]);
tran (encrypt_out[29], \encrypt_out.tdata [29]);
tran (encrypt_out[28], \encrypt_out.tdata [28]);
tran (encrypt_out[27], \encrypt_out.tdata [27]);
tran (encrypt_out[26], \encrypt_out.tdata [26]);
tran (encrypt_out[25], \encrypt_out.tdata [25]);
tran (encrypt_out[24], \encrypt_out.tdata [24]);
tran (encrypt_out[23], \encrypt_out.tdata [23]);
tran (encrypt_out[22], \encrypt_out.tdata [22]);
tran (encrypt_out[21], \encrypt_out.tdata [21]);
tran (encrypt_out[20], \encrypt_out.tdata [20]);
tran (encrypt_out[19], \encrypt_out.tdata [19]);
tran (encrypt_out[18], \encrypt_out.tdata [18]);
tran (encrypt_out[17], \encrypt_out.tdata [17]);
tran (encrypt_out[16], \encrypt_out.tdata [16]);
tran (encrypt_out[15], \encrypt_out.tdata [15]);
tran (encrypt_out[14], \encrypt_out.tdata [14]);
tran (encrypt_out[13], \encrypt_out.tdata [13]);
tran (encrypt_out[12], \encrypt_out.tdata [12]);
tran (encrypt_out[11], \encrypt_out.tdata [11]);
tran (encrypt_out[10], \encrypt_out.tdata [10]);
tran (encrypt_out[9], \encrypt_out.tdata [9]);
tran (encrypt_out[8], \encrypt_out.tdata [8]);
tran (encrypt_out[7], \encrypt_out.tdata [7]);
tran (encrypt_out[6], \encrypt_out.tdata [6]);
tran (encrypt_out[5], \encrypt_out.tdata [5]);
tran (encrypt_out[4], \encrypt_out.tdata [4]);
tran (encrypt_out[3], \encrypt_out.tdata [3]);
tran (encrypt_out[2], \encrypt_out.tdata [2]);
tran (encrypt_out[1], \encrypt_out.tdata [1]);
tran (encrypt_out[0], \encrypt_out.tdata [0]);
Q_BUF U0 ( .A(n324), .Z(cceip_validate_ob_afull));
Q_BUF U1 ( .A(n324), .Z(cceip_encrypt_ob_afull));
Q_BUF U2 ( .A(n324), .Z(_zy_simnet_cio_11));
Q_BUF U3 ( .A(n324), .Z(_zy_simnet_cio_6));
Q_BUF U4 ( .A(_zy_sva_brcm_cceip_3_reset_or), .Z(_zy_sva_brcm_cceip_2_reset_or));
Q_BUF U5 ( .A(_zy_sva_brcm_cceip_4_reset_or), .Z(_zy_sva_brcm_cceip_3_reset_or));
Q_BUF U6 ( .A(_zy_sva_brcm_cceip_1_reset_or), .Z(_zy_sva_brcm_cceip_4_reset_or));
Q_ASSIGN U7 ( .B(encrypt_out[0]), .A(key_tlv_w0[0]));
Q_ASSIGN U8 ( .B(encrypt_out[1]), .A(key_tlv_w0[1]));
Q_ASSIGN U9 ( .B(encrypt_out[2]), .A(key_tlv_w0[2]));
Q_ASSIGN U10 ( .B(encrypt_out[3]), .A(key_tlv_w0[3]));
Q_ASSIGN U11 ( .B(encrypt_out[4]), .A(key_tlv_w0[4]));
Q_ASSIGN U12 ( .B(encrypt_out[5]), .A(key_tlv_w0[5]));
Q_ASSIGN U13 ( .B(encrypt_out[6]), .A(key_tlv_w0[6]));
Q_ASSIGN U14 ( .B(encrypt_out[7]), .A(key_tlv_w0[7]));
Q_ASSIGN U15 ( .B(encrypt_out[8]), .A(key_tlv_w0[8]));
Q_ASSIGN U16 ( .B(encrypt_out[9]), .A(key_tlv_w0[9]));
Q_ASSIGN U17 ( .B(encrypt_out[10]), .A(key_tlv_w0[10]));
Q_ASSIGN U18 ( .B(encrypt_out[11]), .A(key_tlv_w0[11]));
Q_ASSIGN U19 ( .B(encrypt_out[12]), .A(key_tlv_w0[12]));
Q_ASSIGN U20 ( .B(encrypt_out[13]), .A(key_tlv_w0[13]));
Q_ASSIGN U21 ( .B(encrypt_out[14]), .A(key_tlv_w0[14]));
Q_ASSIGN U22 ( .B(encrypt_out[15]), .A(key_tlv_w0[15]));
Q_ASSIGN U23 ( .B(encrypt_out[16]), .A(key_tlv_w0[16]));
Q_ASSIGN U24 ( .B(encrypt_out[17]), .A(key_tlv_w0[17]));
Q_ASSIGN U25 ( .B(encrypt_out[18]), .A(key_tlv_w0[18]));
Q_ASSIGN U26 ( .B(encrypt_out[19]), .A(key_tlv_w0[19]));
Q_ASSIGN U27 ( .B(encrypt_out[20]), .A(key_tlv_w0[20]));
Q_ASSIGN U28 ( .B(encrypt_out[21]), .A(key_tlv_w0[21]));
Q_ASSIGN U29 ( .B(encrypt_out[22]), .A(key_tlv_w0[22]));
Q_ASSIGN U30 ( .B(encrypt_out[23]), .A(key_tlv_w0[23]));
Q_ASSIGN U31 ( .B(encrypt_out[24]), .A(key_tlv_w0[24]));
Q_ASSIGN U32 ( .B(encrypt_out[25]), .A(key_tlv_w0[25]));
Q_ASSIGN U33 ( .B(encrypt_out[26]), .A(key_tlv_w0[26]));
Q_ASSIGN U34 ( .B(encrypt_out[27]), .A(key_tlv_w0[27]));
Q_ASSIGN U35 ( .B(encrypt_out[28]), .A(key_tlv_w0[28]));
Q_ASSIGN U36 ( .B(encrypt_out[29]), .A(key_tlv_w0[29]));
Q_ASSIGN U37 ( .B(encrypt_out[30]), .A(key_tlv_w0[30]));
Q_ASSIGN U38 ( .B(encrypt_out[31]), .A(key_tlv_w0[31]));
Q_ASSIGN U39 ( .B(encrypt_out[32]), .A(key_tlv_w0[32]));
Q_ASSIGN U40 ( .B(encrypt_out[33]), .A(key_tlv_w0[33]));
Q_ASSIGN U41 ( .B(encrypt_out[34]), .A(key_tlv_w0[34]));
Q_ASSIGN U42 ( .B(encrypt_out[35]), .A(key_tlv_w0[35]));
Q_ASSIGN U43 ( .B(encrypt_out[36]), .A(key_tlv_w0[36]));
Q_ASSIGN U44 ( .B(encrypt_out[37]), .A(key_tlv_w0[37]));
Q_ASSIGN U45 ( .B(encrypt_out[38]), .A(key_tlv_w0[38]));
Q_ASSIGN U46 ( .B(encrypt_out[39]), .A(key_tlv_w0[39]));
Q_ASSIGN U47 ( .B(encrypt_out[40]), .A(key_tlv_w0[40]));
Q_ASSIGN U48 ( .B(encrypt_out[41]), .A(key_tlv_w0[41]));
Q_ASSIGN U49 ( .B(encrypt_out[42]), .A(key_tlv_w0[42]));
Q_ASSIGN U50 ( .B(encrypt_out[43]), .A(key_tlv_w0[43]));
Q_ASSIGN U51 ( .B(encrypt_out[44]), .A(key_tlv_w0[44]));
Q_ASSIGN U52 ( .B(encrypt_out[45]), .A(key_tlv_w0[45]));
Q_ASSIGN U53 ( .B(encrypt_out[46]), .A(key_tlv_w0[46]));
Q_ASSIGN U54 ( .B(encrypt_out[47]), .A(key_tlv_w0[47]));
Q_ASSIGN U55 ( .B(encrypt_out[48]), .A(key_tlv_w0[48]));
Q_ASSIGN U56 ( .B(encrypt_out[49]), .A(key_tlv_w0[49]));
Q_ASSIGN U57 ( .B(encrypt_out[50]), .A(key_tlv_w0[50]));
Q_ASSIGN U58 ( .B(encrypt_out[51]), .A(key_tlv_w0[51]));
Q_ASSIGN U59 ( .B(encrypt_out[52]), .A(key_tlv_w0[52]));
Q_ASSIGN U60 ( .B(encrypt_out[53]), .A(key_tlv_w0[53]));
Q_ASSIGN U61 ( .B(encrypt_out[54]), .A(key_tlv_w0[54]));
Q_ASSIGN U62 ( .B(encrypt_out[55]), .A(key_tlv_w0[55]));
Q_ASSIGN U63 ( .B(encrypt_out[56]), .A(key_tlv_w0[56]));
Q_ASSIGN U64 ( .B(encrypt_out[57]), .A(key_tlv_w0[57]));
Q_ASSIGN U65 ( .B(encrypt_out[58]), .A(key_tlv_w0[58]));
Q_ASSIGN U66 ( .B(encrypt_out[59]), .A(key_tlv_w0[59]));
Q_ASSIGN U67 ( .B(encrypt_out[60]), .A(key_tlv_w0[60]));
Q_ASSIGN U68 ( .B(encrypt_out[61]), .A(key_tlv_w0[61]));
Q_ASSIGN U69 ( .B(encrypt_out[62]), .A(key_tlv_w0[62]));
Q_ASSIGN U70 ( .B(encrypt_out[63]), .A(key_tlv_w0[63]));
Q_BUF U71 ( .A(validate_out_ack), .Z(encrypt_out_ack));
Q_BUF U72 ( .A(n324), .Z(\cceip_ob_tlv[3][104] ));
Q_BUF U73 ( .A(n324), .Z(\cceip_ob_tlv[3][103] ));
Q_BUF U74 ( .A(n324), .Z(\cceip_ob_tlv[3][102] ));
Q_BUF U75 ( .A(n324), .Z(\cceip_ob_tlv[3][101] ));
Q_BUF U76 ( .A(n324), .Z(\cceip_ob_tlv[3][100] ));
Q_BUF U77 ( .A(n324), .Z(\cceip_ob_tlv[3][99] ));
Q_BUF U78 ( .A(n324), .Z(\cceip_ob_tlv[3][98] ));
Q_BUF U79 ( .A(n324), .Z(\cceip_ob_tlv[3][97] ));
Q_BUF U80 ( .A(n324), .Z(\cceip_ob_tlv[3][96] ));
Q_BUF U81 ( .A(n324), .Z(\cceip_ob_tlv[3][95] ));
Q_BUF U82 ( .A(n324), .Z(\cceip_ob_tlv[3][94] ));
Q_BUF U83 ( .A(n324), .Z(\cceip_ob_tlv[3][93] ));
Q_BUF U84 ( .A(\cceip_ob_tlv[3][81] ), .Z(\cceip_ob_tlv[3][82] ));
Q_BUF U85 ( .A(n324), .Z(\cceip_ob_tlv[2][104] ));
Q_BUF U86 ( .A(n324), .Z(\cceip_ob_tlv[2][103] ));
Q_BUF U87 ( .A(n324), .Z(\cceip_ob_tlv[2][102] ));
Q_BUF U88 ( .A(n324), .Z(\cceip_ob_tlv[2][101] ));
Q_BUF U89 ( .A(n324), .Z(\cceip_ob_tlv[2][100] ));
Q_BUF U90 ( .A(n324), .Z(\cceip_ob_tlv[2][99] ));
Q_BUF U91 ( .A(n324), .Z(\cceip_ob_tlv[2][98] ));
Q_BUF U92 ( .A(n324), .Z(\cceip_ob_tlv[2][97] ));
Q_BUF U93 ( .A(n324), .Z(\cceip_ob_tlv[2][96] ));
Q_BUF U94 ( .A(n324), .Z(\cceip_ob_tlv[2][95] ));
Q_BUF U95 ( .A(n324), .Z(\cceip_ob_tlv[2][94] ));
Q_BUF U96 ( .A(n324), .Z(\cceip_ob_tlv[2][93] ));
Q_BUF U97 ( .A(\cceip_ob_tlv[2][81] ), .Z(\cceip_ob_tlv[2][82] ));
Q_BUF U98 ( .A(n324), .Z(\cceip_ob_tlv[1][104] ));
Q_BUF U99 ( .A(n324), .Z(\cceip_ob_tlv[1][103] ));
Q_BUF U100 ( .A(n324), .Z(\cceip_ob_tlv[1][102] ));
Q_BUF U101 ( .A(n324), .Z(\cceip_ob_tlv[1][101] ));
Q_BUF U102 ( .A(n324), .Z(\cceip_ob_tlv[1][100] ));
Q_BUF U103 ( .A(n324), .Z(\cceip_ob_tlv[1][99] ));
Q_BUF U104 ( .A(n324), .Z(\cceip_ob_tlv[1][98] ));
Q_BUF U105 ( .A(n324), .Z(\cceip_ob_tlv[1][97] ));
Q_BUF U106 ( .A(n324), .Z(\cceip_ob_tlv[1][96] ));
Q_BUF U107 ( .A(n324), .Z(\cceip_ob_tlv[1][95] ));
Q_BUF U108 ( .A(n324), .Z(\cceip_ob_tlv[1][94] ));
Q_BUF U109 ( .A(n324), .Z(\cceip_ob_tlv[1][93] ));
Q_BUF U110 ( .A(\cceip_ob_tlv[1][81] ), .Z(\cceip_ob_tlv[1][82] ));
Q_BUF U111 ( .A(n324), .Z(\cceip_ob_tlv[0][104] ));
Q_BUF U112 ( .A(n324), .Z(\cceip_ob_tlv[0][103] ));
Q_BUF U113 ( .A(n324), .Z(\cceip_ob_tlv[0][102] ));
Q_BUF U114 ( .A(n324), .Z(\cceip_ob_tlv[0][101] ));
Q_BUF U115 ( .A(n324), .Z(\cceip_ob_tlv[0][100] ));
Q_BUF U116 ( .A(n324), .Z(\cceip_ob_tlv[0][99] ));
Q_BUF U117 ( .A(n324), .Z(\cceip_ob_tlv[0][98] ));
Q_BUF U118 ( .A(n324), .Z(\cceip_ob_tlv[0][97] ));
Q_BUF U119 ( .A(n324), .Z(\cceip_ob_tlv[0][96] ));
Q_BUF U120 ( .A(n324), .Z(\cceip_ob_tlv[0][95] ));
Q_BUF U121 ( .A(n324), .Z(\cceip_ob_tlv[0][94] ));
Q_BUF U122 ( .A(n324), .Z(\cceip_ob_tlv[0][93] ));
Q_BUF U123 ( .A(\cceip_ob_tlv[0][81] ), .Z(\cceip_ob_tlv[0][82] ));
wire [2:0] n519 = 3'b000;
Q_ASSERT \engine_3_.brcm_cceip  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_cceip_4_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_cceip_4_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n519[0]));
// pragma CVASTRPROP INSTANCE "\engine_3_.brcm_cceip " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\engine_3_.brcm_cceip " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_key_tlv_compare_split.v"
//pragma CVAINTPROP INSTANCE "\engine_3_.brcm_cceip " ASSERT_LINE 265
wire [2:0] n520 = 3'b000;
Q_ASSERT \engine_2_.brcm_cceip  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_cceip_3_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_cceip_3_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n520[0]));
// pragma CVASTRPROP INSTANCE "\engine_2_.brcm_cceip " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\engine_2_.brcm_cceip " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_key_tlv_compare_split.v"
//pragma CVAINTPROP INSTANCE "\engine_2_.brcm_cceip " ASSERT_LINE 265
wire [2:0] n521 = 3'b000;
Q_ASSERT \engine_1_.brcm_cceip  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_cceip_2_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_cceip_2_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n521[0]));
// pragma CVASTRPROP INSTANCE "\engine_1_.brcm_cceip " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\engine_1_.brcm_cceip " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_key_tlv_compare_split.v"
//pragma CVAINTPROP INSTANCE "\engine_1_.brcm_cceip " ASSERT_LINE 265
wire [2:0] n522 = 3'b000;
Q_ASSERT \engine_0_.brcm_cceip  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_cceip_1_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_cceip_1_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n522[0]));
// pragma CVASTRPROP INSTANCE "\engine_0_.brcm_cceip " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\engine_0_.brcm_cceip " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_key_tlv_compare_split.v"
//pragma CVAINTPROP INSTANCE "\engine_0_.brcm_cceip " ASSERT_LINE 265
cr_kme_fifo_xcm44 validate_fifo ( .fifo_in_stall( cceip_validate_ob_full), 
	.fifo_out( _zy_simnet_validate_out_7_w$[0:105]), .fifo_out_valid( 
	validate_out_valid), .fifo_overflow( _zy_simnet_dio_8), 
	.fifo_underflow( _zy_simnet_dio_9), .clk( clk), .rst_n( rst_n), 
	.fifo_in( cceip_validate_ob_tlv[105:0]), .fifo_in_valid( 
	cceip_validate_ob_wr), .fifo_out_ack( 
	_zy_simnet_validate_out_ack_10_w$), .fifo_in_stall_override( 
	_zy_simnet_cio_11));
cr_kme_fifo_xcm44 encrypt_fifo ( .fifo_in_stall( cceip_encrypt_ob_full), 
	.fifo_out( _zy_simnet_encrypt_out_2_w$[0:105]), .fifo_out_valid( 
	encrypt_out_valid), .fifo_overflow( _zy_simnet_dio_3), 
	.fifo_underflow( _zy_simnet_dio_4), .clk( clk), .rst_n( rst_n), 
	.fifo_in( cceip_encrypt_ob_tlv[105:0]), .fifo_in_valid( 
	cceip_encrypt_ob_wr), .fifo_out_ack( 
	_zy_simnet_encrypt_out_ack_5_w$), .fifo_in_stall_override( 
	_zy_simnet_cio_6));
ixc_sample_logic_1_3 _zz_zy_sva_b3 ( _zy_sva_b3, _zy_sva_b3_t);
ixc_sample_logic_1_3 _zz_zy_sva_b2 ( _zy_sva_b2, _zy_sva_b2_t);
ixc_sample_logic_1_3 _zz_zy_sva_b1 ( _zy_sva_b1, _zy_sva_b1_t);
ixc_sample_logic_1_3 _zz_zy_sva_b0 ( _zy_sva_b0, _zy_sva_b0_t);
Q_AN03 U134 ( .A0(encrypt_out_ack), .A1(encrypt_out[82]), .A2(n6), .Z(_zy_sva_b3_t));
Q_AN02 U135 ( .A0(engine_select[0]), .A1(engine_select[1]), .Z(n6));
Q_AN03 U136 ( .A0(encrypt_out_ack), .A1(encrypt_out[82]), .A2(n5), .Z(_zy_sva_b2_t));
Q_AN02 U137 ( .A0(n4), .A1(engine_select[1]), .Z(n5));
Q_AN03 U138 ( .A0(encrypt_out_ack), .A1(encrypt_out[82]), .A2(n3), .Z(_zy_sva_b1_t));
Q_AN02 U139 ( .A0(engine_select[0]), .A1(n2), .Z(n3));
Q_AN03 U140 ( .A0(encrypt_out_ack), .A1(encrypt_out[82]), .A2(n1), .Z(_zy_sva_b0_t));
Q_NR02 U141 ( .A0(engine_select[0]), .A1(engine_select[1]), .Z(n1));
Q_INV U142 ( .A(rst_n), .Z(_zy_sva_brcm_cceip_1_reset_or));
ixc_assign _zz_strnp_6 ( _zy_simnet_validate_out_ack_10_w$, encrypt_out_ack);
ixc_assign_106 _zz_strnp_5 ( validate_out[105:0], 
	_zy_simnet_validate_out_7_w$[0:105]);
ixc_assign _zz_strnp_4 ( _zy_simnet_encrypt_out_ack_5_w$, encrypt_out_ack);
ixc_assign_106 _zz_strnp_3 ( encrypt_out[105:0], 
	_zy_simnet_encrypt_out_2_w$[0:105]);
ixc_assign_424 _zz_strnp_2 ( _zy_simnet_cceip_ob_tlv_1_w$[0:423], { 
	\cceip_ob_tlv[3][105] , n324, n324, n324, n324, n324, n324, n324, 
	n324, n324, n324, n324, n324, \cceip_ob_tlv[3][92] , 
	\cceip_ob_tlv[3][91] , \cceip_ob_tlv[3][90] , \cceip_ob_tlv[3][89] , 
	\cceip_ob_tlv[3][88] , \cceip_ob_tlv[3][87] , \cceip_ob_tlv[3][86] , 
	\cceip_ob_tlv[3][85] , \cceip_ob_tlv[3][84] , \cceip_ob_tlv[3][83] , 
	\cceip_ob_tlv[3][81] , \cceip_ob_tlv[3][81] , \cceip_ob_tlv[3][80] , 
	\cceip_ob_tlv[3][79] , \cceip_ob_tlv[3][78] , \cceip_ob_tlv[3][77] , 
	\cceip_ob_tlv[3][76] , \cceip_ob_tlv[3][75] , \cceip_ob_tlv[3][74] , 
	\cceip_ob_tlv[3][73] , \cceip_ob_tlv[3][72] , \cceip_ob_tlv[3][71] , 
	\cceip_ob_tlv[3][70] , \cceip_ob_tlv[3][69] , \cceip_ob_tlv[3][68] , 
	\cceip_ob_tlv[3][67] , \cceip_ob_tlv[3][66] , \cceip_ob_tlv[3][65] , 
	\cceip_ob_tlv[3][64] , \cceip_ob_tlv[3][63] , \cceip_ob_tlv[3][62] , 
	\cceip_ob_tlv[3][61] , \cceip_ob_tlv[3][60] , \cceip_ob_tlv[3][59] , 
	\cceip_ob_tlv[3][58] , \cceip_ob_tlv[3][57] , \cceip_ob_tlv[3][56] , 
	\cceip_ob_tlv[3][55] , \cceip_ob_tlv[3][54] , \cceip_ob_tlv[3][53] , 
	\cceip_ob_tlv[3][52] , \cceip_ob_tlv[3][51] , \cceip_ob_tlv[3][50] , 
	\cceip_ob_tlv[3][49] , \cceip_ob_tlv[3][48] , \cceip_ob_tlv[3][47] , 
	\cceip_ob_tlv[3][46] , \cceip_ob_tlv[3][45] , \cceip_ob_tlv[3][44] , 
	\cceip_ob_tlv[3][43] , \cceip_ob_tlv[3][42] , \cceip_ob_tlv[3][41] , 
	\cceip_ob_tlv[3][40] , \cceip_ob_tlv[3][39] , \cceip_ob_tlv[3][38] , 
	\cceip_ob_tlv[3][37] , \cceip_ob_tlv[3][36] , \cceip_ob_tlv[3][35] , 
	\cceip_ob_tlv[3][34] , \cceip_ob_tlv[3][33] , \cceip_ob_tlv[3][32] , 
	\cceip_ob_tlv[3][31] , \cceip_ob_tlv[3][30] , \cceip_ob_tlv[3][29] , 
	\cceip_ob_tlv[3][28] , \cceip_ob_tlv[3][27] , \cceip_ob_tlv[3][26] , 
	\cceip_ob_tlv[3][25] , \cceip_ob_tlv[3][24] , \cceip_ob_tlv[3][23] , 
	\cceip_ob_tlv[3][22] , \cceip_ob_tlv[3][21] , \cceip_ob_tlv[3][20] , 
	\cceip_ob_tlv[3][19] , \cceip_ob_tlv[3][18] , \cceip_ob_tlv[3][17] , 
	\cceip_ob_tlv[3][16] , \cceip_ob_tlv[3][15] , \cceip_ob_tlv[3][14] , 
	\cceip_ob_tlv[3][13] , \cceip_ob_tlv[3][12] , \cceip_ob_tlv[3][11] , 
	\cceip_ob_tlv[3][10] , \cceip_ob_tlv[3][9] , \cceip_ob_tlv[3][8] , 
	\cceip_ob_tlv[3][7] , \cceip_ob_tlv[3][6] , \cceip_ob_tlv[3][5] , 
	\cceip_ob_tlv[3][4] , \cceip_ob_tlv[3][3] , \cceip_ob_tlv[3][2] , 
	\cceip_ob_tlv[3][1] , \cceip_ob_tlv[3][0] , \cceip_ob_tlv[2][105] , 
	n324, n324, n324, n324, n324, n324, n324, n324, n324, n324, n324, 
	n324, \cceip_ob_tlv[2][92] , \cceip_ob_tlv[2][91] , 
	\cceip_ob_tlv[2][90] , \cceip_ob_tlv[2][89] , \cceip_ob_tlv[2][88] , 
	\cceip_ob_tlv[2][87] , \cceip_ob_tlv[2][86] , \cceip_ob_tlv[2][85] , 
	\cceip_ob_tlv[2][84] , \cceip_ob_tlv[2][83] , \cceip_ob_tlv[2][81] , 
	\cceip_ob_tlv[2][81] , \cceip_ob_tlv[2][80] , \cceip_ob_tlv[2][79] , 
	\cceip_ob_tlv[2][78] , \cceip_ob_tlv[2][77] , \cceip_ob_tlv[2][76] , 
	\cceip_ob_tlv[2][75] , \cceip_ob_tlv[2][74] , \cceip_ob_tlv[2][73] , 
	\cceip_ob_tlv[2][72] , \cceip_ob_tlv[2][71] , \cceip_ob_tlv[2][70] , 
	\cceip_ob_tlv[2][69] , \cceip_ob_tlv[2][68] , \cceip_ob_tlv[2][67] , 
	\cceip_ob_tlv[2][66] , \cceip_ob_tlv[2][65] , \cceip_ob_tlv[2][64] , 
	\cceip_ob_tlv[2][63] , \cceip_ob_tlv[2][62] , \cceip_ob_tlv[2][61] , 
	\cceip_ob_tlv[2][60] , \cceip_ob_tlv[2][59] , \cceip_ob_tlv[2][58] , 
	\cceip_ob_tlv[2][57] , \cceip_ob_tlv[2][56] , \cceip_ob_tlv[2][55] , 
	\cceip_ob_tlv[2][54] , \cceip_ob_tlv[2][53] , \cceip_ob_tlv[2][52] , 
	\cceip_ob_tlv[2][51] , \cceip_ob_tlv[2][50] , \cceip_ob_tlv[2][49] , 
	\cceip_ob_tlv[2][48] , \cceip_ob_tlv[2][47] , \cceip_ob_tlv[2][46] , 
	\cceip_ob_tlv[2][45] , \cceip_ob_tlv[2][44] , \cceip_ob_tlv[2][43] , 
	\cceip_ob_tlv[2][42] , \cceip_ob_tlv[2][41] , \cceip_ob_tlv[2][40] , 
	\cceip_ob_tlv[2][39] , \cceip_ob_tlv[2][38] , \cceip_ob_tlv[2][37] , 
	\cceip_ob_tlv[2][36] , \cceip_ob_tlv[2][35] , \cceip_ob_tlv[2][34] , 
	\cceip_ob_tlv[2][33] , \cceip_ob_tlv[2][32] , \cceip_ob_tlv[2][31] , 
	\cceip_ob_tlv[2][30] , \cceip_ob_tlv[2][29] , \cceip_ob_tlv[2][28] , 
	\cceip_ob_tlv[2][27] , \cceip_ob_tlv[2][26] , \cceip_ob_tlv[2][25] , 
	\cceip_ob_tlv[2][24] , \cceip_ob_tlv[2][23] , \cceip_ob_tlv[2][22] , 
	\cceip_ob_tlv[2][21] , \cceip_ob_tlv[2][20] , \cceip_ob_tlv[2][19] , 
	\cceip_ob_tlv[2][18] , \cceip_ob_tlv[2][17] , \cceip_ob_tlv[2][16] , 
	\cceip_ob_tlv[2][15] , \cceip_ob_tlv[2][14] , \cceip_ob_tlv[2][13] , 
	\cceip_ob_tlv[2][12] , \cceip_ob_tlv[2][11] , \cceip_ob_tlv[2][10] , 
	\cceip_ob_tlv[2][9] , \cceip_ob_tlv[2][8] , \cceip_ob_tlv[2][7] , 
	\cceip_ob_tlv[2][6] , \cceip_ob_tlv[2][5] , \cceip_ob_tlv[2][4] , 
	\cceip_ob_tlv[2][3] , \cceip_ob_tlv[2][2] , \cceip_ob_tlv[2][1] , 
	\cceip_ob_tlv[2][0] , \cceip_ob_tlv[1][105] , n324, n324, n324, n324, 
	n324, n324, n324, n324, n324, n324, n324, n324, 
	\cceip_ob_tlv[1][92] , \cceip_ob_tlv[1][91] , \cceip_ob_tlv[1][90] , 
	\cceip_ob_tlv[1][89] , \cceip_ob_tlv[1][88] , \cceip_ob_tlv[1][87] , 
	\cceip_ob_tlv[1][86] , \cceip_ob_tlv[1][85] , \cceip_ob_tlv[1][84] , 
	\cceip_ob_tlv[1][83] , \cceip_ob_tlv[1][81] , \cceip_ob_tlv[1][81] , 
	\cceip_ob_tlv[1][80] , \cceip_ob_tlv[1][79] , \cceip_ob_tlv[1][78] , 
	\cceip_ob_tlv[1][77] , \cceip_ob_tlv[1][76] , \cceip_ob_tlv[1][75] , 
	\cceip_ob_tlv[1][74] , \cceip_ob_tlv[1][73] , \cceip_ob_tlv[1][72] , 
	\cceip_ob_tlv[1][71] , \cceip_ob_tlv[1][70] , \cceip_ob_tlv[1][69] , 
	\cceip_ob_tlv[1][68] , \cceip_ob_tlv[1][67] , \cceip_ob_tlv[1][66] , 
	\cceip_ob_tlv[1][65] , \cceip_ob_tlv[1][64] , \cceip_ob_tlv[1][63] , 
	\cceip_ob_tlv[1][62] , \cceip_ob_tlv[1][61] , \cceip_ob_tlv[1][60] , 
	\cceip_ob_tlv[1][59] , \cceip_ob_tlv[1][58] , \cceip_ob_tlv[1][57] , 
	\cceip_ob_tlv[1][56] , \cceip_ob_tlv[1][55] , \cceip_ob_tlv[1][54] , 
	\cceip_ob_tlv[1][53] , \cceip_ob_tlv[1][52] , \cceip_ob_tlv[1][51] , 
	\cceip_ob_tlv[1][50] , \cceip_ob_tlv[1][49] , \cceip_ob_tlv[1][48] , 
	\cceip_ob_tlv[1][47] , \cceip_ob_tlv[1][46] , \cceip_ob_tlv[1][45] , 
	\cceip_ob_tlv[1][44] , \cceip_ob_tlv[1][43] , \cceip_ob_tlv[1][42] , 
	\cceip_ob_tlv[1][41] , \cceip_ob_tlv[1][40] , \cceip_ob_tlv[1][39] , 
	\cceip_ob_tlv[1][38] , \cceip_ob_tlv[1][37] , \cceip_ob_tlv[1][36] , 
	\cceip_ob_tlv[1][35] , \cceip_ob_tlv[1][34] , \cceip_ob_tlv[1][33] , 
	\cceip_ob_tlv[1][32] , \cceip_ob_tlv[1][31] , \cceip_ob_tlv[1][30] , 
	\cceip_ob_tlv[1][29] , \cceip_ob_tlv[1][28] , \cceip_ob_tlv[1][27] , 
	\cceip_ob_tlv[1][26] , \cceip_ob_tlv[1][25] , \cceip_ob_tlv[1][24] , 
	\cceip_ob_tlv[1][23] , \cceip_ob_tlv[1][22] , \cceip_ob_tlv[1][21] , 
	\cceip_ob_tlv[1][20] , \cceip_ob_tlv[1][19] , \cceip_ob_tlv[1][18] , 
	\cceip_ob_tlv[1][17] , \cceip_ob_tlv[1][16] , \cceip_ob_tlv[1][15] , 
	\cceip_ob_tlv[1][14] , \cceip_ob_tlv[1][13] , \cceip_ob_tlv[1][12] , 
	\cceip_ob_tlv[1][11] , \cceip_ob_tlv[1][10] , \cceip_ob_tlv[1][9] , 
	\cceip_ob_tlv[1][8] , \cceip_ob_tlv[1][7] , \cceip_ob_tlv[1][6] , 
	\cceip_ob_tlv[1][5] , \cceip_ob_tlv[1][4] , \cceip_ob_tlv[1][3] , 
	\cceip_ob_tlv[1][2] , \cceip_ob_tlv[1][1] , \cceip_ob_tlv[1][0] , 
	\cceip_ob_tlv[0][105] , n324, n324, n324, n324, n324, n324, n324, 
	n324, n324, n324, n324, n324, \cceip_ob_tlv[0][92] , 
	\cceip_ob_tlv[0][91] , \cceip_ob_tlv[0][90] , \cceip_ob_tlv[0][89] , 
	\cceip_ob_tlv[0][88] , \cceip_ob_tlv[0][87] , \cceip_ob_tlv[0][86] , 
	\cceip_ob_tlv[0][85] , \cceip_ob_tlv[0][84] , \cceip_ob_tlv[0][83] , 
	\cceip_ob_tlv[0][81] , \cceip_ob_tlv[0][81] , \cceip_ob_tlv[0][80] , 
	\cceip_ob_tlv[0][79] , \cceip_ob_tlv[0][78] , \cceip_ob_tlv[0][77] , 
	\cceip_ob_tlv[0][76] , \cceip_ob_tlv[0][75] , \cceip_ob_tlv[0][74] , 
	\cceip_ob_tlv[0][73] , \cceip_ob_tlv[0][72] , \cceip_ob_tlv[0][71] , 
	\cceip_ob_tlv[0][70] , \cceip_ob_tlv[0][69] , \cceip_ob_tlv[0][68] , 
	\cceip_ob_tlv[0][67] , \cceip_ob_tlv[0][66] , \cceip_ob_tlv[0][65] , 
	\cceip_ob_tlv[0][64] , \cceip_ob_tlv[0][63] , \cceip_ob_tlv[0][62] , 
	\cceip_ob_tlv[0][61] , \cceip_ob_tlv[0][60] , \cceip_ob_tlv[0][59] , 
	\cceip_ob_tlv[0][58] , \cceip_ob_tlv[0][57] , \cceip_ob_tlv[0][56] , 
	\cceip_ob_tlv[0][55] , \cceip_ob_tlv[0][54] , \cceip_ob_tlv[0][53] , 
	\cceip_ob_tlv[0][52] , \cceip_ob_tlv[0][51] , \cceip_ob_tlv[0][50] , 
	\cceip_ob_tlv[0][49] , \cceip_ob_tlv[0][48] , \cceip_ob_tlv[0][47] , 
	\cceip_ob_tlv[0][46] , \cceip_ob_tlv[0][45] , \cceip_ob_tlv[0][44] , 
	\cceip_ob_tlv[0][43] , \cceip_ob_tlv[0][42] , \cceip_ob_tlv[0][41] , 
	\cceip_ob_tlv[0][40] , \cceip_ob_tlv[0][39] , \cceip_ob_tlv[0][38] , 
	\cceip_ob_tlv[0][37] , \cceip_ob_tlv[0][36] , \cceip_ob_tlv[0][35] , 
	\cceip_ob_tlv[0][34] , \cceip_ob_tlv[0][33] , \cceip_ob_tlv[0][32] , 
	\cceip_ob_tlv[0][31] , \cceip_ob_tlv[0][30] , \cceip_ob_tlv[0][29] , 
	\cceip_ob_tlv[0][28] , \cceip_ob_tlv[0][27] , \cceip_ob_tlv[0][26] , 
	\cceip_ob_tlv[0][25] , \cceip_ob_tlv[0][24] , \cceip_ob_tlv[0][23] , 
	\cceip_ob_tlv[0][22] , \cceip_ob_tlv[0][21] , \cceip_ob_tlv[0][20] , 
	\cceip_ob_tlv[0][19] , \cceip_ob_tlv[0][18] , \cceip_ob_tlv[0][17] , 
	\cceip_ob_tlv[0][16] , \cceip_ob_tlv[0][15] , \cceip_ob_tlv[0][14] , 
	\cceip_ob_tlv[0][13] , \cceip_ob_tlv[0][12] , \cceip_ob_tlv[0][11] , 
	\cceip_ob_tlv[0][10] , \cceip_ob_tlv[0][9] , \cceip_ob_tlv[0][8] , 
	\cceip_ob_tlv[0][7] , \cceip_ob_tlv[0][6] , \cceip_ob_tlv[0][5] , 
	\cceip_ob_tlv[0][4] , \cceip_ob_tlv[0][3] , \cceip_ob_tlv[0][2] , 
	\cceip_ob_tlv[0][1] , \cceip_ob_tlv[0][0] });
ixc_assign_4 _zz_strnp_1 ( _zy_simnet_cceip_ob_wr_0_w$[0:3], cceip_ob_wr[3:0]);
ixc_assign _zz_strnp_0 ( set_key_tlv_miscmp_int, set_tlv_miscmp);
Q_AN02 U150 ( .A0(rst_n), .A1(_zy_sva_b0), .Z(n7));
Q_AN02 U151 ( .A0(rst_n), .A1(_zy_sva_b1), .Z(n8));
Q_AN02 U152 ( .A0(rst_n), .A1(_zy_sva_b2), .Z(n9));
Q_AN02 U153 ( .A0(rst_n), .A1(_zy_sva_b3), .Z(n10));
Q_FDP1 \engine_select_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_engine_select[0]), .Q(engine_select[0]), .QN(n4));
Q_FDP1 \engine_select_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_engine_select[1]), .Q(engine_select[1]), .QN(n2));
Q_FDP1 \cur_state_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_state[0]), .Q(cur_state[0]), .QN( ));
Q_AN02 U157 ( .A0(encrypt_out_ack), .A1(encrypt_out[82]), .Z(clr_tlv_miscmp));
Q_MX02 U158 ( .S(cur_state[0]), .A0(encrypt_out_valid), .A1(n11), .Z(nxt_state[0]));
Q_INV U159 ( .A(clr_tlv_miscmp), .Z(n11));
Q_INV U160 ( .A(suppress_key_tlvs), .Z(n12));
Q_INV U161 ( .A(encrypt_out[0]), .Z(n13));
Q_INV U162 ( .A(encrypt_out[1]), .Z(n14));
Q_INV U163 ( .A(encrypt_out[2]), .Z(n15));
Q_INV U164 ( .A(encrypt_out[3]), .Z(n16));
Q_INV U165 ( .A(encrypt_out[4]), .Z(n17));
Q_INV U166 ( .A(encrypt_out[5]), .Z(n18));
Q_INV U167 ( .A(encrypt_out[6]), .Z(n19));
Q_INV U168 ( .A(encrypt_out[7]), .Z(n20));
Q_INV U169 ( .A(encrypt_out[8]), .Z(n21));
Q_INV U170 ( .A(encrypt_out[9]), .Z(n22));
Q_INV U171 ( .A(encrypt_out[10]), .Z(n23));
Q_INV U172 ( .A(encrypt_out[11]), .Z(n24));
Q_INV U173 ( .A(encrypt_out[12]), .Z(n25));
Q_INV U174 ( .A(encrypt_out[13]), .Z(n26));
Q_INV U175 ( .A(encrypt_out[14]), .Z(n27));
Q_INV U176 ( .A(encrypt_out[15]), .Z(n28));
Q_INV U177 ( .A(encrypt_out[16]), .Z(n29));
Q_INV U178 ( .A(encrypt_out[17]), .Z(n30));
Q_INV U179 ( .A(encrypt_out[18]), .Z(n31));
Q_INV U180 ( .A(encrypt_out[19]), .Z(n32));
Q_INV U181 ( .A(encrypt_out[20]), .Z(n33));
Q_INV U182 ( .A(encrypt_out[21]), .Z(n34));
Q_INV U183 ( .A(encrypt_out[22]), .Z(n35));
Q_INV U184 ( .A(encrypt_out[23]), .Z(n36));
Q_INV U185 ( .A(encrypt_out[24]), .Z(n37));
Q_INV U186 ( .A(encrypt_out[25]), .Z(n38));
Q_INV U187 ( .A(encrypt_out[26]), .Z(n39));
Q_INV U188 ( .A(encrypt_out[27]), .Z(n40));
Q_INV U189 ( .A(encrypt_out[28]), .Z(n41));
Q_INV U190 ( .A(encrypt_out[29]), .Z(n42));
Q_INV U191 ( .A(encrypt_out[30]), .Z(n43));
Q_INV U192 ( .A(encrypt_out[31]), .Z(n44));
Q_INV U193 ( .A(encrypt_out[32]), .Z(n45));
Q_INV U194 ( .A(encrypt_out[33]), .Z(n46));
Q_INV U195 ( .A(encrypt_out[34]), .Z(n47));
Q_INV U196 ( .A(encrypt_out[35]), .Z(n48));
Q_INV U197 ( .A(encrypt_out[36]), .Z(n49));
Q_INV U198 ( .A(encrypt_out[37]), .Z(n50));
Q_INV U199 ( .A(encrypt_out[38]), .Z(n51));
Q_INV U200 ( .A(encrypt_out[39]), .Z(n52));
Q_INV U201 ( .A(encrypt_out[40]), .Z(n53));
Q_INV U202 ( .A(encrypt_out[41]), .Z(n54));
Q_INV U203 ( .A(encrypt_out[42]), .Z(n55));
Q_INV U204 ( .A(encrypt_out[43]), .Z(n56));
Q_INV U205 ( .A(encrypt_out[44]), .Z(n57));
Q_INV U206 ( .A(encrypt_out[45]), .Z(n58));
Q_INV U207 ( .A(encrypt_out[46]), .Z(n59));
Q_INV U208 ( .A(encrypt_out[47]), .Z(n60));
Q_INV U209 ( .A(encrypt_out[48]), .Z(n61));
Q_INV U210 ( .A(encrypt_out[49]), .Z(n62));
Q_INV U211 ( .A(encrypt_out[50]), .Z(n63));
Q_INV U212 ( .A(encrypt_out[51]), .Z(n64));
Q_INV U213 ( .A(encrypt_out[52]), .Z(n65));
Q_INV U214 ( .A(encrypt_out[53]), .Z(n66));
Q_INV U215 ( .A(encrypt_out[54]), .Z(n67));
Q_INV U216 ( .A(encrypt_out[55]), .Z(n68));
Q_INV U217 ( .A(encrypt_out[56]), .Z(n69));
Q_INV U218 ( .A(encrypt_out[57]), .Z(n70));
Q_INV U219 ( .A(encrypt_out[58]), .Z(n71));
Q_INV U220 ( .A(encrypt_out[59]), .Z(n72));
Q_INV U221 ( .A(encrypt_out[60]), .Z(n73));
Q_INV U222 ( .A(encrypt_out[61]), .Z(n74));
Q_INV U223 ( .A(encrypt_out[62]), .Z(n75));
Q_INV U224 ( .A(encrypt_out[63]), .Z(n76));
Q_AN03 U225 ( .A0(tlv_miscmp), .A1(encrypt_out[82]), .A2(encrypt_out_ack), .Z(n245));
Q_XNR2 U226 ( .A0(encrypt_out[0]), .A1(validate_out[0]), .Z(n77));
Q_XNR2 U227 ( .A0(encrypt_out[1]), .A1(validate_out[1]), .Z(n78));
Q_XNR2 U228 ( .A0(encrypt_out[2]), .A1(validate_out[2]), .Z(n79));
Q_XNR2 U229 ( .A0(encrypt_out[3]), .A1(validate_out[3]), .Z(n80));
Q_XNR2 U230 ( .A0(encrypt_out[4]), .A1(validate_out[4]), .Z(n81));
Q_XNR2 U231 ( .A0(encrypt_out[5]), .A1(validate_out[5]), .Z(n82));
Q_XNR2 U232 ( .A0(encrypt_out[6]), .A1(validate_out[6]), .Z(n83));
Q_XNR2 U233 ( .A0(encrypt_out[7]), .A1(validate_out[7]), .Z(n84));
Q_XNR2 U234 ( .A0(encrypt_out[8]), .A1(validate_out[8]), .Z(n85));
Q_XNR2 U235 ( .A0(encrypt_out[9]), .A1(validate_out[9]), .Z(n86));
Q_XNR2 U236 ( .A0(encrypt_out[10]), .A1(validate_out[10]), .Z(n87));
Q_XNR2 U237 ( .A0(encrypt_out[11]), .A1(validate_out[11]), .Z(n88));
Q_XNR2 U238 ( .A0(encrypt_out[12]), .A1(validate_out[12]), .Z(n89));
Q_XNR2 U239 ( .A0(encrypt_out[13]), .A1(validate_out[13]), .Z(n90));
Q_XNR2 U240 ( .A0(encrypt_out[14]), .A1(validate_out[14]), .Z(n91));
Q_XNR2 U241 ( .A0(encrypt_out[15]), .A1(validate_out[15]), .Z(n92));
Q_XNR2 U242 ( .A0(encrypt_out[16]), .A1(validate_out[16]), .Z(n93));
Q_XNR2 U243 ( .A0(encrypt_out[17]), .A1(validate_out[17]), .Z(n94));
Q_XNR2 U244 ( .A0(encrypt_out[18]), .A1(validate_out[18]), .Z(n95));
Q_XNR2 U245 ( .A0(encrypt_out[19]), .A1(validate_out[19]), .Z(n96));
Q_XNR2 U246 ( .A0(encrypt_out[20]), .A1(validate_out[20]), .Z(n97));
Q_XNR2 U247 ( .A0(encrypt_out[21]), .A1(validate_out[21]), .Z(n98));
Q_XNR2 U248 ( .A0(encrypt_out[22]), .A1(validate_out[22]), .Z(n99));
Q_XNR2 U249 ( .A0(encrypt_out[23]), .A1(validate_out[23]), .Z(n100));
Q_XNR2 U250 ( .A0(encrypt_out[24]), .A1(validate_out[24]), .Z(n101));
Q_XNR2 U251 ( .A0(encrypt_out[25]), .A1(validate_out[25]), .Z(n102));
Q_XNR2 U252 ( .A0(encrypt_out[26]), .A1(validate_out[26]), .Z(n103));
Q_XNR2 U253 ( .A0(encrypt_out[27]), .A1(validate_out[27]), .Z(n104));
Q_XNR2 U254 ( .A0(encrypt_out[28]), .A1(validate_out[28]), .Z(n105));
Q_XNR2 U255 ( .A0(encrypt_out[29]), .A1(validate_out[29]), .Z(n106));
Q_XNR2 U256 ( .A0(encrypt_out[30]), .A1(validate_out[30]), .Z(n107));
Q_XNR2 U257 ( .A0(encrypt_out[31]), .A1(validate_out[31]), .Z(n108));
Q_XNR2 U258 ( .A0(encrypt_out[32]), .A1(validate_out[32]), .Z(n109));
Q_XNR2 U259 ( .A0(encrypt_out[33]), .A1(validate_out[33]), .Z(n110));
Q_XNR2 U260 ( .A0(encrypt_out[34]), .A1(validate_out[34]), .Z(n111));
Q_XNR2 U261 ( .A0(encrypt_out[35]), .A1(validate_out[35]), .Z(n112));
Q_XNR2 U262 ( .A0(encrypt_out[36]), .A1(validate_out[36]), .Z(n113));
Q_XNR2 U263 ( .A0(encrypt_out[37]), .A1(validate_out[37]), .Z(n114));
Q_XNR2 U264 ( .A0(encrypt_out[38]), .A1(validate_out[38]), .Z(n115));
Q_XNR2 U265 ( .A0(encrypt_out[39]), .A1(validate_out[39]), .Z(n116));
Q_XNR2 U266 ( .A0(encrypt_out[40]), .A1(validate_out[40]), .Z(n117));
Q_XNR2 U267 ( .A0(encrypt_out[41]), .A1(validate_out[41]), .Z(n118));
Q_XNR2 U268 ( .A0(encrypt_out[42]), .A1(validate_out[42]), .Z(n119));
Q_XNR2 U269 ( .A0(encrypt_out[43]), .A1(validate_out[43]), .Z(n120));
Q_XNR2 U270 ( .A0(encrypt_out[44]), .A1(validate_out[44]), .Z(n121));
Q_XNR2 U271 ( .A0(encrypt_out[45]), .A1(validate_out[45]), .Z(n122));
Q_XNR2 U272 ( .A0(encrypt_out[46]), .A1(validate_out[46]), .Z(n123));
Q_XNR2 U273 ( .A0(encrypt_out[47]), .A1(validate_out[47]), .Z(n124));
Q_XNR2 U274 ( .A0(encrypt_out[48]), .A1(validate_out[48]), .Z(n125));
Q_XNR2 U275 ( .A0(encrypt_out[49]), .A1(validate_out[49]), .Z(n126));
Q_XNR2 U276 ( .A0(encrypt_out[50]), .A1(validate_out[50]), .Z(n127));
Q_XNR2 U277 ( .A0(encrypt_out[51]), .A1(validate_out[51]), .Z(n128));
Q_XNR2 U278 ( .A0(encrypt_out[52]), .A1(validate_out[52]), .Z(n129));
Q_XNR2 U279 ( .A0(encrypt_out[53]), .A1(validate_out[53]), .Z(n130));
Q_XNR2 U280 ( .A0(encrypt_out[54]), .A1(validate_out[54]), .Z(n131));
Q_XNR2 U281 ( .A0(encrypt_out[55]), .A1(validate_out[55]), .Z(n132));
Q_XNR2 U282 ( .A0(encrypt_out[56]), .A1(validate_out[56]), .Z(n133));
Q_XNR2 U283 ( .A0(encrypt_out[57]), .A1(validate_out[57]), .Z(n134));
Q_XNR2 U284 ( .A0(encrypt_out[58]), .A1(validate_out[58]), .Z(n135));
Q_XNR2 U285 ( .A0(encrypt_out[59]), .A1(validate_out[59]), .Z(n136));
Q_XNR2 U286 ( .A0(encrypt_out[60]), .A1(validate_out[60]), .Z(n137));
Q_XNR2 U287 ( .A0(encrypt_out[61]), .A1(validate_out[61]), .Z(n138));
Q_XNR2 U288 ( .A0(encrypt_out[62]), .A1(validate_out[62]), .Z(n139));
Q_XNR2 U289 ( .A0(encrypt_out[63]), .A1(validate_out[63]), .Z(n140));
Q_XNR2 U290 ( .A0(encrypt_out[64]), .A1(validate_out[64]), .Z(n141));
Q_XNR2 U291 ( .A0(encrypt_out[65]), .A1(validate_out[65]), .Z(n142));
Q_XNR2 U292 ( .A0(encrypt_out[66]), .A1(validate_out[66]), .Z(n143));
Q_XNR2 U293 ( .A0(encrypt_out[67]), .A1(validate_out[67]), .Z(n144));
Q_XNR2 U294 ( .A0(encrypt_out[68]), .A1(validate_out[68]), .Z(n145));
Q_XNR2 U295 ( .A0(encrypt_out[69]), .A1(validate_out[69]), .Z(n146));
Q_XNR2 U296 ( .A0(encrypt_out[70]), .A1(validate_out[70]), .Z(n147));
Q_XNR2 U297 ( .A0(encrypt_out[71]), .A1(validate_out[71]), .Z(n148));
Q_XNR2 U298 ( .A0(encrypt_out[72]), .A1(validate_out[72]), .Z(n149));
Q_XNR2 U299 ( .A0(encrypt_out[73]), .A1(validate_out[73]), .Z(n150));
Q_XNR2 U300 ( .A0(encrypt_out[74]), .A1(validate_out[74]), .Z(n151));
Q_XNR2 U301 ( .A0(encrypt_out[75]), .A1(validate_out[75]), .Z(n152));
Q_XNR2 U302 ( .A0(encrypt_out[76]), .A1(validate_out[76]), .Z(n153));
Q_XNR2 U303 ( .A0(encrypt_out[77]), .A1(validate_out[77]), .Z(n154));
Q_XNR2 U304 ( .A0(encrypt_out[78]), .A1(validate_out[78]), .Z(n155));
Q_XNR2 U305 ( .A0(encrypt_out[79]), .A1(validate_out[79]), .Z(n156));
Q_XNR2 U306 ( .A0(encrypt_out[80]), .A1(validate_out[80]), .Z(n157));
Q_XNR2 U307 ( .A0(encrypt_out[81]), .A1(validate_out[81]), .Z(n158));
Q_XNR2 U308 ( .A0(encrypt_out[82]), .A1(validate_out[82]), .Z(n159));
Q_XNR2 U309 ( .A0(encrypt_out[83]), .A1(validate_out[83]), .Z(n160));
Q_XNR2 U310 ( .A0(encrypt_out[84]), .A1(validate_out[84]), .Z(n161));
Q_XNR2 U311 ( .A0(encrypt_out[85]), .A1(validate_out[85]), .Z(n162));
Q_XNR2 U312 ( .A0(encrypt_out[86]), .A1(validate_out[86]), .Z(n163));
Q_XNR2 U313 ( .A0(encrypt_out[87]), .A1(validate_out[87]), .Z(n164));
Q_XNR2 U314 ( .A0(encrypt_out[88]), .A1(validate_out[88]), .Z(n165));
Q_XNR2 U315 ( .A0(encrypt_out[89]), .A1(validate_out[89]), .Z(n166));
Q_XNR2 U316 ( .A0(encrypt_out[90]), .A1(validate_out[90]), .Z(n167));
Q_XNR2 U317 ( .A0(encrypt_out[91]), .A1(validate_out[91]), .Z(n168));
Q_XNR2 U318 ( .A0(encrypt_out[92]), .A1(validate_out[92]), .Z(n169));
Q_XNR2 U319 ( .A0(encrypt_out[93]), .A1(validate_out[93]), .Z(n170));
Q_XNR2 U320 ( .A0(encrypt_out[94]), .A1(validate_out[94]), .Z(n171));
Q_XNR2 U321 ( .A0(encrypt_out[95]), .A1(validate_out[95]), .Z(n172));
Q_XNR2 U322 ( .A0(encrypt_out[96]), .A1(validate_out[96]), .Z(n173));
Q_XNR2 U323 ( .A0(encrypt_out[97]), .A1(validate_out[97]), .Z(n174));
Q_XNR2 U324 ( .A0(encrypt_out[98]), .A1(validate_out[98]), .Z(n175));
Q_XNR2 U325 ( .A0(encrypt_out[99]), .A1(validate_out[99]), .Z(n176));
Q_XNR2 U326 ( .A0(encrypt_out[100]), .A1(validate_out[100]), .Z(n177));
Q_XNR2 U327 ( .A0(encrypt_out[101]), .A1(validate_out[101]), .Z(n178));
Q_XNR2 U328 ( .A0(encrypt_out[102]), .A1(validate_out[102]), .Z(n179));
Q_XNR2 U329 ( .A0(encrypt_out[103]), .A1(validate_out[103]), .Z(n180));
Q_XNR2 U330 ( .A0(encrypt_out[104]), .A1(validate_out[104]), .Z(n181));
Q_XNR2 U331 ( .A0(encrypt_out[105]), .A1(validate_out[105]), .Z(n182));
Q_AN03 U332 ( .A0(n182), .A1(n181), .A2(n180), .Z(n183));
Q_AN03 U333 ( .A0(n179), .A1(n178), .A2(n177), .Z(n184));
Q_AN03 U334 ( .A0(n176), .A1(n175), .A2(n174), .Z(n185));
Q_AN03 U335 ( .A0(n173), .A1(n172), .A2(n171), .Z(n186));
Q_AN03 U336 ( .A0(n170), .A1(n169), .A2(n168), .Z(n187));
Q_AN03 U337 ( .A0(n167), .A1(n166), .A2(n165), .Z(n188));
Q_AN03 U338 ( .A0(n164), .A1(n163), .A2(n162), .Z(n189));
Q_AN03 U339 ( .A0(n161), .A1(n160), .A2(n159), .Z(n190));
Q_AN03 U340 ( .A0(n158), .A1(n157), .A2(n156), .Z(n191));
Q_AN03 U341 ( .A0(n155), .A1(n154), .A2(n153), .Z(n192));
Q_AN03 U342 ( .A0(n152), .A1(n151), .A2(n150), .Z(n193));
Q_AN03 U343 ( .A0(n149), .A1(n148), .A2(n147), .Z(n194));
Q_AN03 U344 ( .A0(n146), .A1(n145), .A2(n144), .Z(n195));
Q_AN03 U345 ( .A0(n143), .A1(n142), .A2(n141), .Z(n196));
Q_AN03 U346 ( .A0(n140), .A1(n139), .A2(n138), .Z(n197));
Q_AN03 U347 ( .A0(n137), .A1(n136), .A2(n135), .Z(n198));
Q_AN03 U348 ( .A0(n134), .A1(n133), .A2(n132), .Z(n199));
Q_AN03 U349 ( .A0(n131), .A1(n130), .A2(n129), .Z(n200));
Q_AN03 U350 ( .A0(n128), .A1(n127), .A2(n126), .Z(n201));
Q_AN03 U351 ( .A0(n125), .A1(n124), .A2(n123), .Z(n202));
Q_AN03 U352 ( .A0(n122), .A1(n121), .A2(n120), .Z(n203));
Q_AN03 U353 ( .A0(n119), .A1(n118), .A2(n117), .Z(n204));
Q_AN03 U354 ( .A0(n116), .A1(n115), .A2(n114), .Z(n205));
Q_AN03 U355 ( .A0(n113), .A1(n112), .A2(n111), .Z(n206));
Q_AN03 U356 ( .A0(n110), .A1(n109), .A2(n108), .Z(n207));
Q_AN03 U357 ( .A0(n107), .A1(n106), .A2(n105), .Z(n208));
Q_AN03 U358 ( .A0(n104), .A1(n103), .A2(n102), .Z(n209));
Q_AN03 U359 ( .A0(n101), .A1(n100), .A2(n99), .Z(n210));
Q_AN03 U360 ( .A0(n98), .A1(n97), .A2(n96), .Z(n211));
Q_AN03 U361 ( .A0(n95), .A1(n94), .A2(n93), .Z(n212));
Q_AN03 U362 ( .A0(n92), .A1(n91), .A2(n90), .Z(n213));
Q_AN03 U363 ( .A0(n89), .A1(n88), .A2(n87), .Z(n214));
Q_AN03 U364 ( .A0(n86), .A1(n85), .A2(n84), .Z(n215));
Q_AN03 U365 ( .A0(n83), .A1(n82), .A2(n81), .Z(n216));
Q_AN03 U366 ( .A0(n80), .A1(n79), .A2(n78), .Z(n217));
Q_AN03 U367 ( .A0(n77), .A1(n183), .A2(n184), .Z(n218));
Q_AN03 U368 ( .A0(n185), .A1(n186), .A2(n187), .Z(n219));
Q_AN03 U369 ( .A0(n188), .A1(n189), .A2(n190), .Z(n220));
Q_AN03 U370 ( .A0(n191), .A1(n192), .A2(n193), .Z(n221));
Q_AN03 U371 ( .A0(n194), .A1(n195), .A2(n196), .Z(n222));
Q_AN03 U372 ( .A0(n197), .A1(n198), .A2(n199), .Z(n223));
Q_AN03 U373 ( .A0(n200), .A1(n201), .A2(n202), .Z(n224));
Q_AN03 U374 ( .A0(n203), .A1(n204), .A2(n205), .Z(n225));
Q_AN03 U375 ( .A0(n206), .A1(n207), .A2(n208), .Z(n226));
Q_AN03 U376 ( .A0(n209), .A1(n210), .A2(n211), .Z(n227));
Q_AN03 U377 ( .A0(n212), .A1(n213), .A2(n214), .Z(n228));
Q_AN03 U378 ( .A0(n215), .A1(n216), .A2(n217), .Z(n229));
Q_AN03 U379 ( .A0(n218), .A1(n219), .A2(n220), .Z(n230));
Q_AN03 U380 ( .A0(n221), .A1(n222), .A2(n223), .Z(n231));
Q_AN03 U381 ( .A0(n224), .A1(n225), .A2(n226), .Z(n232));
Q_AN03 U382 ( .A0(n227), .A1(n228), .A2(n229), .Z(n233));
Q_AN03 U383 ( .A0(n230), .A1(n231), .A2(n232), .Z(n234));
Q_ND02 U384 ( .A0(n233), .A1(n234), .Z(n235));
Q_MX04 U385 ( .S0(engine_select[0]), .S1(engine_select[1]), .A0(cceip_ob_full[0]), .A1(cceip_ob_full[1]), .A2(cceip_ob_full[2]), .A3(cceip_ob_full[3]), .Z(n236));
Q_INV U386 ( .A(n236), .Z(n237));
Q_AN03 U387 ( .A0(n237), .A1(encrypt_out_valid), .A2(validate_out_valid), .Z(n246));
Q_AN02 U388 ( .A0(encrypt_out_ack), .A1(n235), .Z(set_tlv_miscmp));
Q_AN02 U389 ( .A0(cur_state[0]), .A1(engine_select[0]), .Z(nxt_engine_select[0]));
Q_AN02 U390 ( .A0(cur_state[0]), .A1(engine_select[1]), .Z(nxt_engine_select[1]));
Q_NR02 U391 ( .A0(n238), .A1(suppress_key_tlvs), .Z(cceip_ob_wr[0]));
Q_NR02 U392 ( .A0(n240), .A1(suppress_key_tlvs), .Z(cceip_ob_wr[1]));
Q_NR02 U393 ( .A0(n242), .A1(suppress_key_tlvs), .Z(cceip_ob_wr[2]));
Q_OR02 U394 ( .A0(engine_select[0]), .A1(n239), .Z(n238));
Q_OR02 U395 ( .A0(n4), .A1(n239), .Z(n240));
Q_OR02 U396 ( .A0(engine_select[1]), .A1(n241), .Z(n239));
Q_INV U397 ( .A(encrypt_out_ack), .Z(n241));
Q_OR02 U398 ( .A0(engine_select[0]), .A1(n243), .Z(n242));
Q_INV U399 ( .A(n244), .Z(n243));
Q_AN03 U400 ( .A0(engine_select[0]), .A1(n244), .A2(n12), .Z(cceip_ob_wr[3]));
Q_AN02 U401 ( .A0(engine_select[1]), .A1(encrypt_out_ack), .Z(n244));
Q_AN02 U402 ( .A0(n246), .A1(cur_state[0]), .Z(validate_out_ack));
Q_OR02 U403 ( .A0(clr_tlv_miscmp), .A1(set_tlv_miscmp), .Z(n247));
Q_AN02 U404 ( .A0(engine_select[0]), .A1(encrypt_out_ack), .Z(n248));
Q_INV U405 ( .A(n248), .Z(n249));
Q_NR02 U406 ( .A0(n244), .A1(n248), .Z(n250));
Q_AN02 U407 ( .A0(engine_select[0]), .A1(n245), .Z(n251));
Q_AN02 U408 ( .A0(engine_select[1]), .A1(n245), .Z(n252));
Q_INV U409 ( .A(n251), .Z(n253));
Q_INV U410 ( .A(n252), .Z(n254));
Q_NR02 U411 ( .A0(n252), .A1(n251), .Z(n255));
Q_AN02 U412 ( .A0(n254), .A1(n251), .Z(n256));
Q_AN02 U413 ( .A0(n252), .A1(n253), .Z(n257));
Q_AN02 U414 ( .A0(n252), .A1(n251), .Z(n258));
Q_AN02 U415 ( .A0(n255), .A1(n245), .Z(n259));
Q_AN02 U416 ( .A0(n243), .A1(n248), .Z(\cceip_ob_tlv[1][92] ));
Q_AN02 U417 ( .A0(n244), .A1(n249), .Z(\cceip_ob_tlv[2][92] ));
Q_AN02 U418 ( .A0(n244), .A1(n248), .Z(\cceip_ob_tlv[3][92] ));
Q_AN02 U419 ( .A0(n250), .A1(encrypt_out_ack), .Z(\cceip_ob_tlv[0][92] ));
Q_AN02 U420 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[0]), .Z(n260));
Q_MX02 U421 ( .S(n259), .A0(n260), .A1(n13), .Z(\cceip_ob_tlv[0][0] ));
Q_AN02 U422 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[1]), .Z(n261));
Q_MX02 U423 ( .S(n259), .A0(n261), .A1(n14), .Z(\cceip_ob_tlv[0][1] ));
Q_AN02 U424 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[2]), .Z(n262));
Q_MX02 U425 ( .S(n259), .A0(n262), .A1(n15), .Z(\cceip_ob_tlv[0][2] ));
Q_AN02 U426 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[3]), .Z(n263));
Q_MX02 U427 ( .S(n259), .A0(n263), .A1(n16), .Z(\cceip_ob_tlv[0][3] ));
Q_AN02 U428 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[4]), .Z(n264));
Q_MX02 U429 ( .S(n259), .A0(n264), .A1(n17), .Z(\cceip_ob_tlv[0][4] ));
Q_AN02 U430 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[5]), .Z(n265));
Q_MX02 U431 ( .S(n259), .A0(n265), .A1(n18), .Z(\cceip_ob_tlv[0][5] ));
Q_AN02 U432 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[6]), .Z(n266));
Q_MX02 U433 ( .S(n259), .A0(n266), .A1(n19), .Z(\cceip_ob_tlv[0][6] ));
Q_AN02 U434 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[7]), .Z(n267));
Q_MX02 U435 ( .S(n259), .A0(n267), .A1(n20), .Z(\cceip_ob_tlv[0][7] ));
Q_AN02 U436 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[8]), .Z(n268));
Q_MX02 U437 ( .S(n259), .A0(n268), .A1(n21), .Z(\cceip_ob_tlv[0][8] ));
Q_AN02 U438 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[9]), .Z(n269));
Q_MX02 U439 ( .S(n259), .A0(n269), .A1(n22), .Z(\cceip_ob_tlv[0][9] ));
Q_AN02 U440 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[10]), .Z(n270));
Q_MX02 U441 ( .S(n259), .A0(n270), .A1(n23), .Z(\cceip_ob_tlv[0][10] ));
Q_AN02 U442 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[11]), .Z(n271));
Q_MX02 U443 ( .S(n259), .A0(n271), .A1(n24), .Z(\cceip_ob_tlv[0][11] ));
Q_AN02 U444 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[12]), .Z(n272));
Q_MX02 U445 ( .S(n259), .A0(n272), .A1(n25), .Z(\cceip_ob_tlv[0][12] ));
Q_AN02 U446 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[13]), .Z(n273));
Q_MX02 U447 ( .S(n259), .A0(n273), .A1(n26), .Z(\cceip_ob_tlv[0][13] ));
Q_AN02 U448 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[14]), .Z(n274));
Q_MX02 U449 ( .S(n259), .A0(n274), .A1(n27), .Z(\cceip_ob_tlv[0][14] ));
Q_AN02 U450 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[15]), .Z(n275));
Q_MX02 U451 ( .S(n259), .A0(n275), .A1(n28), .Z(\cceip_ob_tlv[0][15] ));
Q_AN02 U452 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[16]), .Z(n276));
Q_MX02 U453 ( .S(n259), .A0(n276), .A1(n29), .Z(\cceip_ob_tlv[0][16] ));
Q_AN02 U454 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[17]), .Z(n277));
Q_MX02 U455 ( .S(n259), .A0(n277), .A1(n30), .Z(\cceip_ob_tlv[0][17] ));
Q_AN02 U456 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[18]), .Z(n278));
Q_MX02 U457 ( .S(n259), .A0(n278), .A1(n31), .Z(\cceip_ob_tlv[0][18] ));
Q_AN02 U458 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[19]), .Z(n279));
Q_MX02 U459 ( .S(n259), .A0(n279), .A1(n32), .Z(\cceip_ob_tlv[0][19] ));
Q_AN02 U460 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[20]), .Z(n280));
Q_MX02 U461 ( .S(n259), .A0(n280), .A1(n33), .Z(\cceip_ob_tlv[0][20] ));
Q_AN02 U462 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[21]), .Z(n281));
Q_MX02 U463 ( .S(n259), .A0(n281), .A1(n34), .Z(\cceip_ob_tlv[0][21] ));
Q_AN02 U464 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[22]), .Z(n282));
Q_MX02 U465 ( .S(n259), .A0(n282), .A1(n35), .Z(\cceip_ob_tlv[0][22] ));
Q_AN02 U466 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[23]), .Z(n283));
Q_MX02 U467 ( .S(n259), .A0(n283), .A1(n36), .Z(\cceip_ob_tlv[0][23] ));
Q_AN02 U468 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[24]), .Z(n284));
Q_MX02 U469 ( .S(n259), .A0(n284), .A1(n37), .Z(\cceip_ob_tlv[0][24] ));
Q_AN02 U470 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[25]), .Z(n285));
Q_MX02 U471 ( .S(n259), .A0(n285), .A1(n38), .Z(\cceip_ob_tlv[0][25] ));
Q_AN02 U472 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[26]), .Z(n286));
Q_MX02 U473 ( .S(n259), .A0(n286), .A1(n39), .Z(\cceip_ob_tlv[0][26] ));
Q_AN02 U474 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[27]), .Z(n287));
Q_MX02 U475 ( .S(n259), .A0(n287), .A1(n40), .Z(\cceip_ob_tlv[0][27] ));
Q_AN02 U476 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[28]), .Z(n288));
Q_MX02 U477 ( .S(n259), .A0(n288), .A1(n41), .Z(\cceip_ob_tlv[0][28] ));
Q_AN02 U478 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[29]), .Z(n289));
Q_MX02 U479 ( .S(n259), .A0(n289), .A1(n42), .Z(\cceip_ob_tlv[0][29] ));
Q_AN02 U480 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[30]), .Z(n290));
Q_MX02 U481 ( .S(n259), .A0(n290), .A1(n43), .Z(\cceip_ob_tlv[0][30] ));
Q_AN02 U482 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[31]), .Z(n291));
Q_MX02 U483 ( .S(n259), .A0(n291), .A1(n44), .Z(\cceip_ob_tlv[0][31] ));
Q_AN02 U484 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[32]), .Z(n292));
Q_MX02 U485 ( .S(n259), .A0(n292), .A1(n45), .Z(\cceip_ob_tlv[0][32] ));
Q_AN02 U486 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[33]), .Z(n293));
Q_MX02 U487 ( .S(n259), .A0(n293), .A1(n46), .Z(\cceip_ob_tlv[0][33] ));
Q_AN02 U488 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[34]), .Z(n294));
Q_MX02 U489 ( .S(n259), .A0(n294), .A1(n47), .Z(\cceip_ob_tlv[0][34] ));
Q_AN02 U490 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[35]), .Z(n295));
Q_MX02 U491 ( .S(n259), .A0(n295), .A1(n48), .Z(\cceip_ob_tlv[0][35] ));
Q_AN02 U492 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[36]), .Z(n296));
Q_MX02 U493 ( .S(n259), .A0(n296), .A1(n49), .Z(\cceip_ob_tlv[0][36] ));
Q_AN02 U494 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[37]), .Z(n297));
Q_MX02 U495 ( .S(n259), .A0(n297), .A1(n50), .Z(\cceip_ob_tlv[0][37] ));
Q_AN02 U496 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[38]), .Z(n298));
Q_MX02 U497 ( .S(n259), .A0(n298), .A1(n51), .Z(\cceip_ob_tlv[0][38] ));
Q_AN02 U498 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[39]), .Z(n299));
Q_MX02 U499 ( .S(n259), .A0(n299), .A1(n52), .Z(\cceip_ob_tlv[0][39] ));
Q_AN02 U500 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[40]), .Z(n300));
Q_MX02 U501 ( .S(n259), .A0(n300), .A1(n53), .Z(\cceip_ob_tlv[0][40] ));
Q_AN02 U502 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[41]), .Z(n301));
Q_MX02 U503 ( .S(n259), .A0(n301), .A1(n54), .Z(\cceip_ob_tlv[0][41] ));
Q_AN02 U504 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[42]), .Z(n302));
Q_MX02 U505 ( .S(n259), .A0(n302), .A1(n55), .Z(\cceip_ob_tlv[0][42] ));
Q_AN02 U506 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[43]), .Z(n303));
Q_MX02 U507 ( .S(n259), .A0(n303), .A1(n56), .Z(\cceip_ob_tlv[0][43] ));
Q_AN02 U508 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[44]), .Z(n304));
Q_MX02 U509 ( .S(n259), .A0(n304), .A1(n57), .Z(\cceip_ob_tlv[0][44] ));
Q_AN02 U510 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[45]), .Z(n305));
Q_MX02 U511 ( .S(n259), .A0(n305), .A1(n58), .Z(\cceip_ob_tlv[0][45] ));
Q_AN02 U512 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[46]), .Z(n306));
Q_MX02 U513 ( .S(n259), .A0(n306), .A1(n59), .Z(\cceip_ob_tlv[0][46] ));
Q_AN02 U514 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[47]), .Z(n307));
Q_MX02 U515 ( .S(n259), .A0(n307), .A1(n60), .Z(\cceip_ob_tlv[0][47] ));
Q_AN02 U516 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[48]), .Z(n308));
Q_MX02 U517 ( .S(n259), .A0(n308), .A1(n61), .Z(\cceip_ob_tlv[0][48] ));
Q_AN02 U518 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[49]), .Z(n309));
Q_MX02 U519 ( .S(n259), .A0(n309), .A1(n62), .Z(\cceip_ob_tlv[0][49] ));
Q_AN02 U520 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[50]), .Z(n310));
Q_MX02 U521 ( .S(n259), .A0(n310), .A1(n63), .Z(\cceip_ob_tlv[0][50] ));
Q_AN02 U522 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[51]), .Z(n311));
Q_MX02 U523 ( .S(n259), .A0(n311), .A1(n64), .Z(\cceip_ob_tlv[0][51] ));
Q_AN02 U524 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[52]), .Z(n312));
Q_MX02 U525 ( .S(n259), .A0(n312), .A1(n65), .Z(\cceip_ob_tlv[0][52] ));
Q_AN02 U526 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[53]), .Z(n313));
Q_MX02 U527 ( .S(n259), .A0(n313), .A1(n66), .Z(\cceip_ob_tlv[0][53] ));
Q_AN02 U528 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[54]), .Z(n314));
Q_MX02 U529 ( .S(n259), .A0(n314), .A1(n67), .Z(\cceip_ob_tlv[0][54] ));
Q_AN02 U530 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[55]), .Z(n315));
Q_MX02 U531 ( .S(n259), .A0(n315), .A1(n68), .Z(\cceip_ob_tlv[0][55] ));
Q_AN02 U532 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[56]), .Z(n316));
Q_MX02 U533 ( .S(n259), .A0(n316), .A1(n69), .Z(\cceip_ob_tlv[0][56] ));
Q_AN02 U534 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[57]), .Z(n317));
Q_MX02 U535 ( .S(n259), .A0(n317), .A1(n70), .Z(\cceip_ob_tlv[0][57] ));
Q_AN02 U536 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[58]), .Z(n318));
Q_MX02 U537 ( .S(n259), .A0(n318), .A1(n71), .Z(\cceip_ob_tlv[0][58] ));
Q_AN02 U538 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[59]), .Z(n319));
Q_MX02 U539 ( .S(n259), .A0(n319), .A1(n72), .Z(\cceip_ob_tlv[0][59] ));
Q_AN02 U540 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[60]), .Z(n320));
Q_MX02 U541 ( .S(n259), .A0(n320), .A1(n73), .Z(\cceip_ob_tlv[0][60] ));
Q_AN02 U542 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[61]), .Z(n321));
Q_MX02 U543 ( .S(n259), .A0(n321), .A1(n74), .Z(\cceip_ob_tlv[0][61] ));
Q_AN02 U544 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[62]), .Z(n322));
Q_MX02 U545 ( .S(n259), .A0(n322), .A1(n75), .Z(\cceip_ob_tlv[0][62] ));
Q_AN02 U546 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[63]), .Z(n323));
Q_MX02 U547 ( .S(n259), .A0(n323), .A1(n76), .Z(\cceip_ob_tlv[0][63] ));
Q_AN02 U548 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[64]), .Z(\cceip_ob_tlv[0][64] ));
Q_AN02 U549 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[65]), .Z(\cceip_ob_tlv[0][65] ));
Q_AN02 U550 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[66]), .Z(\cceip_ob_tlv[0][66] ));
Q_AN02 U551 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[67]), .Z(\cceip_ob_tlv[0][67] ));
Q_AN02 U552 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[68]), .Z(\cceip_ob_tlv[0][68] ));
Q_AN02 U553 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[69]), .Z(\cceip_ob_tlv[0][69] ));
Q_AN02 U554 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[70]), .Z(\cceip_ob_tlv[0][70] ));
Q_AN02 U555 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[71]), .Z(\cceip_ob_tlv[0][71] ));
Q_AN02 U556 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[72]), .Z(\cceip_ob_tlv[0][72] ));
Q_AN02 U557 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[73]), .Z(\cceip_ob_tlv[0][73] ));
Q_AN02 U558 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[74]), .Z(\cceip_ob_tlv[0][74] ));
Q_AN02 U559 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[75]), .Z(\cceip_ob_tlv[0][75] ));
Q_AN02 U560 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[76]), .Z(\cceip_ob_tlv[0][76] ));
Q_AN02 U561 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[77]), .Z(\cceip_ob_tlv[0][77] ));
Q_AN02 U562 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[78]), .Z(\cceip_ob_tlv[0][78] ));
Q_AN02 U563 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[79]), .Z(\cceip_ob_tlv[0][79] ));
Q_AN02 U564 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[80]), .Z(\cceip_ob_tlv[0][80] ));
Q_AN02 U565 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[82]), .Z(\cceip_ob_tlv[0][81] ));
Q_AN02 U566 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[83]), .Z(\cceip_ob_tlv[0][83] ));
Q_AN02 U567 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[84]), .Z(\cceip_ob_tlv[0][84] ));
Q_AN02 U568 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[85]), .Z(\cceip_ob_tlv[0][85] ));
Q_AN02 U569 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[86]), .Z(\cceip_ob_tlv[0][86] ));
Q_AN02 U570 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[87]), .Z(\cceip_ob_tlv[0][87] ));
Q_AN02 U571 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[88]), .Z(\cceip_ob_tlv[0][88] ));
Q_AN02 U572 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[89]), .Z(\cceip_ob_tlv[0][89] ));
Q_AN02 U573 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[90]), .Z(\cceip_ob_tlv[0][90] ));
Q_AN02 U574 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[91]), .Z(\cceip_ob_tlv[0][91] ));
Q_AN02 U575 ( .A0(\cceip_ob_tlv[0][92] ), .A1(encrypt_out[105]), .Z(\cceip_ob_tlv[0][105] ));
Q_AN02 U576 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[0]), .Z(n325));
Q_MX02 U577 ( .S(n256), .A0(n325), .A1(n13), .Z(\cceip_ob_tlv[1][0] ));
Q_AN02 U578 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[1]), .Z(n326));
Q_MX02 U579 ( .S(n256), .A0(n326), .A1(n14), .Z(\cceip_ob_tlv[1][1] ));
Q_AN02 U580 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[2]), .Z(n327));
Q_MX02 U581 ( .S(n256), .A0(n327), .A1(n15), .Z(\cceip_ob_tlv[1][2] ));
Q_AN02 U582 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[3]), .Z(n328));
Q_MX02 U583 ( .S(n256), .A0(n328), .A1(n16), .Z(\cceip_ob_tlv[1][3] ));
Q_AN02 U584 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[4]), .Z(n329));
Q_MX02 U585 ( .S(n256), .A0(n329), .A1(n17), .Z(\cceip_ob_tlv[1][4] ));
Q_AN02 U586 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[5]), .Z(n330));
Q_MX02 U587 ( .S(n256), .A0(n330), .A1(n18), .Z(\cceip_ob_tlv[1][5] ));
Q_AN02 U588 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[6]), .Z(n331));
Q_MX02 U589 ( .S(n256), .A0(n331), .A1(n19), .Z(\cceip_ob_tlv[1][6] ));
Q_AN02 U590 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[7]), .Z(n332));
Q_MX02 U591 ( .S(n256), .A0(n332), .A1(n20), .Z(\cceip_ob_tlv[1][7] ));
Q_AN02 U592 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[8]), .Z(n333));
Q_MX02 U593 ( .S(n256), .A0(n333), .A1(n21), .Z(\cceip_ob_tlv[1][8] ));
Q_AN02 U594 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[9]), .Z(n334));
Q_MX02 U595 ( .S(n256), .A0(n334), .A1(n22), .Z(\cceip_ob_tlv[1][9] ));
Q_AN02 U596 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[10]), .Z(n335));
Q_MX02 U597 ( .S(n256), .A0(n335), .A1(n23), .Z(\cceip_ob_tlv[1][10] ));
Q_AN02 U598 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[11]), .Z(n336));
Q_MX02 U599 ( .S(n256), .A0(n336), .A1(n24), .Z(\cceip_ob_tlv[1][11] ));
Q_AN02 U600 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[12]), .Z(n337));
Q_MX02 U601 ( .S(n256), .A0(n337), .A1(n25), .Z(\cceip_ob_tlv[1][12] ));
Q_AN02 U602 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[13]), .Z(n338));
Q_MX02 U603 ( .S(n256), .A0(n338), .A1(n26), .Z(\cceip_ob_tlv[1][13] ));
Q_AN02 U604 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[14]), .Z(n339));
Q_MX02 U605 ( .S(n256), .A0(n339), .A1(n27), .Z(\cceip_ob_tlv[1][14] ));
Q_AN02 U606 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[15]), .Z(n340));
Q_MX02 U607 ( .S(n256), .A0(n340), .A1(n28), .Z(\cceip_ob_tlv[1][15] ));
Q_AN02 U608 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[16]), .Z(n341));
Q_MX02 U609 ( .S(n256), .A0(n341), .A1(n29), .Z(\cceip_ob_tlv[1][16] ));
Q_AN02 U610 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[17]), .Z(n342));
Q_MX02 U611 ( .S(n256), .A0(n342), .A1(n30), .Z(\cceip_ob_tlv[1][17] ));
Q_AN02 U612 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[18]), .Z(n343));
Q_MX02 U613 ( .S(n256), .A0(n343), .A1(n31), .Z(\cceip_ob_tlv[1][18] ));
Q_AN02 U614 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[19]), .Z(n344));
Q_MX02 U615 ( .S(n256), .A0(n344), .A1(n32), .Z(\cceip_ob_tlv[1][19] ));
Q_AN02 U616 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[20]), .Z(n345));
Q_MX02 U617 ( .S(n256), .A0(n345), .A1(n33), .Z(\cceip_ob_tlv[1][20] ));
Q_AN02 U618 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[21]), .Z(n346));
Q_MX02 U619 ( .S(n256), .A0(n346), .A1(n34), .Z(\cceip_ob_tlv[1][21] ));
Q_AN02 U620 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[22]), .Z(n347));
Q_MX02 U621 ( .S(n256), .A0(n347), .A1(n35), .Z(\cceip_ob_tlv[1][22] ));
Q_AN02 U622 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[23]), .Z(n348));
Q_MX02 U623 ( .S(n256), .A0(n348), .A1(n36), .Z(\cceip_ob_tlv[1][23] ));
Q_AN02 U624 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[24]), .Z(n349));
Q_MX02 U625 ( .S(n256), .A0(n349), .A1(n37), .Z(\cceip_ob_tlv[1][24] ));
Q_AN02 U626 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[25]), .Z(n350));
Q_MX02 U627 ( .S(n256), .A0(n350), .A1(n38), .Z(\cceip_ob_tlv[1][25] ));
Q_AN02 U628 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[26]), .Z(n351));
Q_MX02 U629 ( .S(n256), .A0(n351), .A1(n39), .Z(\cceip_ob_tlv[1][26] ));
Q_AN02 U630 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[27]), .Z(n352));
Q_MX02 U631 ( .S(n256), .A0(n352), .A1(n40), .Z(\cceip_ob_tlv[1][27] ));
Q_AN02 U632 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[28]), .Z(n353));
Q_MX02 U633 ( .S(n256), .A0(n353), .A1(n41), .Z(\cceip_ob_tlv[1][28] ));
Q_AN02 U634 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[29]), .Z(n354));
Q_MX02 U635 ( .S(n256), .A0(n354), .A1(n42), .Z(\cceip_ob_tlv[1][29] ));
Q_AN02 U636 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[30]), .Z(n355));
Q_MX02 U637 ( .S(n256), .A0(n355), .A1(n43), .Z(\cceip_ob_tlv[1][30] ));
Q_AN02 U638 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[31]), .Z(n356));
Q_MX02 U639 ( .S(n256), .A0(n356), .A1(n44), .Z(\cceip_ob_tlv[1][31] ));
Q_AN02 U640 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[32]), .Z(n357));
Q_MX02 U641 ( .S(n256), .A0(n357), .A1(n45), .Z(\cceip_ob_tlv[1][32] ));
Q_AN02 U642 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[33]), .Z(n358));
Q_MX02 U643 ( .S(n256), .A0(n358), .A1(n46), .Z(\cceip_ob_tlv[1][33] ));
Q_AN02 U644 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[34]), .Z(n359));
Q_MX02 U645 ( .S(n256), .A0(n359), .A1(n47), .Z(\cceip_ob_tlv[1][34] ));
Q_AN02 U646 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[35]), .Z(n360));
Q_MX02 U647 ( .S(n256), .A0(n360), .A1(n48), .Z(\cceip_ob_tlv[1][35] ));
Q_AN02 U648 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[36]), .Z(n361));
Q_MX02 U649 ( .S(n256), .A0(n361), .A1(n49), .Z(\cceip_ob_tlv[1][36] ));
Q_AN02 U650 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[37]), .Z(n362));
Q_MX02 U651 ( .S(n256), .A0(n362), .A1(n50), .Z(\cceip_ob_tlv[1][37] ));
Q_AN02 U652 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[38]), .Z(n363));
Q_MX02 U653 ( .S(n256), .A0(n363), .A1(n51), .Z(\cceip_ob_tlv[1][38] ));
Q_AN02 U654 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[39]), .Z(n364));
Q_MX02 U655 ( .S(n256), .A0(n364), .A1(n52), .Z(\cceip_ob_tlv[1][39] ));
Q_AN02 U656 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[40]), .Z(n365));
Q_MX02 U657 ( .S(n256), .A0(n365), .A1(n53), .Z(\cceip_ob_tlv[1][40] ));
Q_AN02 U658 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[41]), .Z(n366));
Q_MX02 U659 ( .S(n256), .A0(n366), .A1(n54), .Z(\cceip_ob_tlv[1][41] ));
Q_AN02 U660 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[42]), .Z(n367));
Q_MX02 U661 ( .S(n256), .A0(n367), .A1(n55), .Z(\cceip_ob_tlv[1][42] ));
Q_AN02 U662 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[43]), .Z(n368));
Q_MX02 U663 ( .S(n256), .A0(n368), .A1(n56), .Z(\cceip_ob_tlv[1][43] ));
Q_AN02 U664 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[44]), .Z(n369));
Q_MX02 U665 ( .S(n256), .A0(n369), .A1(n57), .Z(\cceip_ob_tlv[1][44] ));
Q_AN02 U666 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[45]), .Z(n370));
Q_MX02 U667 ( .S(n256), .A0(n370), .A1(n58), .Z(\cceip_ob_tlv[1][45] ));
Q_AN02 U668 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[46]), .Z(n371));
Q_MX02 U669 ( .S(n256), .A0(n371), .A1(n59), .Z(\cceip_ob_tlv[1][46] ));
Q_AN02 U670 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[47]), .Z(n372));
Q_MX02 U671 ( .S(n256), .A0(n372), .A1(n60), .Z(\cceip_ob_tlv[1][47] ));
Q_AN02 U672 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[48]), .Z(n373));
Q_MX02 U673 ( .S(n256), .A0(n373), .A1(n61), .Z(\cceip_ob_tlv[1][48] ));
Q_AN02 U674 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[49]), .Z(n374));
Q_MX02 U675 ( .S(n256), .A0(n374), .A1(n62), .Z(\cceip_ob_tlv[1][49] ));
Q_AN02 U676 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[50]), .Z(n375));
Q_MX02 U677 ( .S(n256), .A0(n375), .A1(n63), .Z(\cceip_ob_tlv[1][50] ));
Q_AN02 U678 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[51]), .Z(n376));
Q_MX02 U679 ( .S(n256), .A0(n376), .A1(n64), .Z(\cceip_ob_tlv[1][51] ));
Q_AN02 U680 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[52]), .Z(n377));
Q_MX02 U681 ( .S(n256), .A0(n377), .A1(n65), .Z(\cceip_ob_tlv[1][52] ));
Q_AN02 U682 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[53]), .Z(n378));
Q_MX02 U683 ( .S(n256), .A0(n378), .A1(n66), .Z(\cceip_ob_tlv[1][53] ));
Q_AN02 U684 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[54]), .Z(n379));
Q_MX02 U685 ( .S(n256), .A0(n379), .A1(n67), .Z(\cceip_ob_tlv[1][54] ));
Q_AN02 U686 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[55]), .Z(n380));
Q_MX02 U687 ( .S(n256), .A0(n380), .A1(n68), .Z(\cceip_ob_tlv[1][55] ));
Q_AN02 U688 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[56]), .Z(n381));
Q_MX02 U689 ( .S(n256), .A0(n381), .A1(n69), .Z(\cceip_ob_tlv[1][56] ));
Q_AN02 U690 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[57]), .Z(n382));
Q_MX02 U691 ( .S(n256), .A0(n382), .A1(n70), .Z(\cceip_ob_tlv[1][57] ));
Q_AN02 U692 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[58]), .Z(n383));
Q_MX02 U693 ( .S(n256), .A0(n383), .A1(n71), .Z(\cceip_ob_tlv[1][58] ));
Q_AN02 U694 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[59]), .Z(n384));
Q_MX02 U695 ( .S(n256), .A0(n384), .A1(n72), .Z(\cceip_ob_tlv[1][59] ));
Q_AN02 U696 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[60]), .Z(n385));
Q_MX02 U697 ( .S(n256), .A0(n385), .A1(n73), .Z(\cceip_ob_tlv[1][60] ));
Q_AN02 U698 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[61]), .Z(n386));
Q_MX02 U699 ( .S(n256), .A0(n386), .A1(n74), .Z(\cceip_ob_tlv[1][61] ));
Q_AN02 U700 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[62]), .Z(n387));
Q_MX02 U701 ( .S(n256), .A0(n387), .A1(n75), .Z(\cceip_ob_tlv[1][62] ));
Q_AN02 U702 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[63]), .Z(n388));
Q_MX02 U703 ( .S(n256), .A0(n388), .A1(n76), .Z(\cceip_ob_tlv[1][63] ));
Q_AN02 U704 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[64]), .Z(\cceip_ob_tlv[1][64] ));
Q_AN02 U705 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[65]), .Z(\cceip_ob_tlv[1][65] ));
Q_AN02 U706 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[66]), .Z(\cceip_ob_tlv[1][66] ));
Q_AN02 U707 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[67]), .Z(\cceip_ob_tlv[1][67] ));
Q_AN02 U708 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[68]), .Z(\cceip_ob_tlv[1][68] ));
Q_AN02 U709 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[69]), .Z(\cceip_ob_tlv[1][69] ));
Q_AN02 U710 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[70]), .Z(\cceip_ob_tlv[1][70] ));
Q_AN02 U711 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[71]), .Z(\cceip_ob_tlv[1][71] ));
Q_AN02 U712 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[72]), .Z(\cceip_ob_tlv[1][72] ));
Q_AN02 U713 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[73]), .Z(\cceip_ob_tlv[1][73] ));
Q_AN02 U714 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[74]), .Z(\cceip_ob_tlv[1][74] ));
Q_AN02 U715 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[75]), .Z(\cceip_ob_tlv[1][75] ));
Q_AN02 U716 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[76]), .Z(\cceip_ob_tlv[1][76] ));
Q_AN02 U717 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[77]), .Z(\cceip_ob_tlv[1][77] ));
Q_AN02 U718 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[78]), .Z(\cceip_ob_tlv[1][78] ));
Q_AN02 U719 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[79]), .Z(\cceip_ob_tlv[1][79] ));
Q_AN02 U720 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[80]), .Z(\cceip_ob_tlv[1][80] ));
Q_AN02 U721 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[82]), .Z(\cceip_ob_tlv[1][81] ));
Q_AN02 U722 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[83]), .Z(\cceip_ob_tlv[1][83] ));
Q_AN02 U723 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[84]), .Z(\cceip_ob_tlv[1][84] ));
Q_AN02 U724 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[85]), .Z(\cceip_ob_tlv[1][85] ));
Q_AN02 U725 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[86]), .Z(\cceip_ob_tlv[1][86] ));
Q_AN02 U726 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[87]), .Z(\cceip_ob_tlv[1][87] ));
Q_AN02 U727 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[88]), .Z(\cceip_ob_tlv[1][88] ));
Q_AN02 U728 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[89]), .Z(\cceip_ob_tlv[1][89] ));
Q_AN02 U729 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[90]), .Z(\cceip_ob_tlv[1][90] ));
Q_AN02 U730 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[91]), .Z(\cceip_ob_tlv[1][91] ));
Q_AN02 U731 ( .A0(\cceip_ob_tlv[1][92] ), .A1(encrypt_out[105]), .Z(\cceip_ob_tlv[1][105] ));
Q_AN02 U732 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[0]), .Z(n389));
Q_MX02 U733 ( .S(n257), .A0(n389), .A1(n13), .Z(\cceip_ob_tlv[2][0] ));
Q_AN02 U734 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[1]), .Z(n390));
Q_MX02 U735 ( .S(n257), .A0(n390), .A1(n14), .Z(\cceip_ob_tlv[2][1] ));
Q_AN02 U736 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[2]), .Z(n391));
Q_MX02 U737 ( .S(n257), .A0(n391), .A1(n15), .Z(\cceip_ob_tlv[2][2] ));
Q_AN02 U738 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[3]), .Z(n392));
Q_MX02 U739 ( .S(n257), .A0(n392), .A1(n16), .Z(\cceip_ob_tlv[2][3] ));
Q_AN02 U740 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[4]), .Z(n393));
Q_MX02 U741 ( .S(n257), .A0(n393), .A1(n17), .Z(\cceip_ob_tlv[2][4] ));
Q_AN02 U742 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[5]), .Z(n394));
Q_MX02 U743 ( .S(n257), .A0(n394), .A1(n18), .Z(\cceip_ob_tlv[2][5] ));
Q_AN02 U744 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[6]), .Z(n395));
Q_MX02 U745 ( .S(n257), .A0(n395), .A1(n19), .Z(\cceip_ob_tlv[2][6] ));
Q_AN02 U746 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[7]), .Z(n396));
Q_MX02 U747 ( .S(n257), .A0(n396), .A1(n20), .Z(\cceip_ob_tlv[2][7] ));
Q_AN02 U748 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[8]), .Z(n397));
Q_MX02 U749 ( .S(n257), .A0(n397), .A1(n21), .Z(\cceip_ob_tlv[2][8] ));
Q_AN02 U750 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[9]), .Z(n398));
Q_MX02 U751 ( .S(n257), .A0(n398), .A1(n22), .Z(\cceip_ob_tlv[2][9] ));
Q_AN02 U752 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[10]), .Z(n399));
Q_MX02 U753 ( .S(n257), .A0(n399), .A1(n23), .Z(\cceip_ob_tlv[2][10] ));
Q_AN02 U754 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[11]), .Z(n400));
Q_MX02 U755 ( .S(n257), .A0(n400), .A1(n24), .Z(\cceip_ob_tlv[2][11] ));
Q_AN02 U756 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[12]), .Z(n401));
Q_MX02 U757 ( .S(n257), .A0(n401), .A1(n25), .Z(\cceip_ob_tlv[2][12] ));
Q_AN02 U758 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[13]), .Z(n402));
Q_MX02 U759 ( .S(n257), .A0(n402), .A1(n26), .Z(\cceip_ob_tlv[2][13] ));
Q_AN02 U760 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[14]), .Z(n403));
Q_MX02 U761 ( .S(n257), .A0(n403), .A1(n27), .Z(\cceip_ob_tlv[2][14] ));
Q_AN02 U762 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[15]), .Z(n404));
Q_MX02 U763 ( .S(n257), .A0(n404), .A1(n28), .Z(\cceip_ob_tlv[2][15] ));
Q_AN02 U764 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[16]), .Z(n405));
Q_MX02 U765 ( .S(n257), .A0(n405), .A1(n29), .Z(\cceip_ob_tlv[2][16] ));
Q_AN02 U766 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[17]), .Z(n406));
Q_MX02 U767 ( .S(n257), .A0(n406), .A1(n30), .Z(\cceip_ob_tlv[2][17] ));
Q_AN02 U768 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[18]), .Z(n407));
Q_MX02 U769 ( .S(n257), .A0(n407), .A1(n31), .Z(\cceip_ob_tlv[2][18] ));
Q_AN02 U770 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[19]), .Z(n408));
Q_MX02 U771 ( .S(n257), .A0(n408), .A1(n32), .Z(\cceip_ob_tlv[2][19] ));
Q_AN02 U772 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[20]), .Z(n409));
Q_MX02 U773 ( .S(n257), .A0(n409), .A1(n33), .Z(\cceip_ob_tlv[2][20] ));
Q_AN02 U774 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[21]), .Z(n410));
Q_MX02 U775 ( .S(n257), .A0(n410), .A1(n34), .Z(\cceip_ob_tlv[2][21] ));
Q_AN02 U776 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[22]), .Z(n411));
Q_MX02 U777 ( .S(n257), .A0(n411), .A1(n35), .Z(\cceip_ob_tlv[2][22] ));
Q_AN02 U778 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[23]), .Z(n412));
Q_MX02 U779 ( .S(n257), .A0(n412), .A1(n36), .Z(\cceip_ob_tlv[2][23] ));
Q_AN02 U780 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[24]), .Z(n413));
Q_MX02 U781 ( .S(n257), .A0(n413), .A1(n37), .Z(\cceip_ob_tlv[2][24] ));
Q_AN02 U782 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[25]), .Z(n414));
Q_MX02 U783 ( .S(n257), .A0(n414), .A1(n38), .Z(\cceip_ob_tlv[2][25] ));
Q_AN02 U784 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[26]), .Z(n415));
Q_MX02 U785 ( .S(n257), .A0(n415), .A1(n39), .Z(\cceip_ob_tlv[2][26] ));
Q_AN02 U786 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[27]), .Z(n416));
Q_MX02 U787 ( .S(n257), .A0(n416), .A1(n40), .Z(\cceip_ob_tlv[2][27] ));
Q_AN02 U788 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[28]), .Z(n417));
Q_MX02 U789 ( .S(n257), .A0(n417), .A1(n41), .Z(\cceip_ob_tlv[2][28] ));
Q_AN02 U790 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[29]), .Z(n418));
Q_MX02 U791 ( .S(n257), .A0(n418), .A1(n42), .Z(\cceip_ob_tlv[2][29] ));
Q_AN02 U792 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[30]), .Z(n419));
Q_MX02 U793 ( .S(n257), .A0(n419), .A1(n43), .Z(\cceip_ob_tlv[2][30] ));
Q_AN02 U794 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[31]), .Z(n420));
Q_MX02 U795 ( .S(n257), .A0(n420), .A1(n44), .Z(\cceip_ob_tlv[2][31] ));
Q_AN02 U796 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[32]), .Z(n421));
Q_MX02 U797 ( .S(n257), .A0(n421), .A1(n45), .Z(\cceip_ob_tlv[2][32] ));
Q_AN02 U798 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[33]), .Z(n422));
Q_MX02 U799 ( .S(n257), .A0(n422), .A1(n46), .Z(\cceip_ob_tlv[2][33] ));
Q_AN02 U800 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[34]), .Z(n423));
Q_MX02 U801 ( .S(n257), .A0(n423), .A1(n47), .Z(\cceip_ob_tlv[2][34] ));
Q_AN02 U802 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[35]), .Z(n424));
Q_MX02 U803 ( .S(n257), .A0(n424), .A1(n48), .Z(\cceip_ob_tlv[2][35] ));
Q_AN02 U804 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[36]), .Z(n425));
Q_MX02 U805 ( .S(n257), .A0(n425), .A1(n49), .Z(\cceip_ob_tlv[2][36] ));
Q_AN02 U806 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[37]), .Z(n426));
Q_MX02 U807 ( .S(n257), .A0(n426), .A1(n50), .Z(\cceip_ob_tlv[2][37] ));
Q_AN02 U808 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[38]), .Z(n427));
Q_MX02 U809 ( .S(n257), .A0(n427), .A1(n51), .Z(\cceip_ob_tlv[2][38] ));
Q_AN02 U810 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[39]), .Z(n428));
Q_MX02 U811 ( .S(n257), .A0(n428), .A1(n52), .Z(\cceip_ob_tlv[2][39] ));
Q_AN02 U812 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[40]), .Z(n429));
Q_MX02 U813 ( .S(n257), .A0(n429), .A1(n53), .Z(\cceip_ob_tlv[2][40] ));
Q_AN02 U814 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[41]), .Z(n430));
Q_MX02 U815 ( .S(n257), .A0(n430), .A1(n54), .Z(\cceip_ob_tlv[2][41] ));
Q_AN02 U816 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[42]), .Z(n431));
Q_MX02 U817 ( .S(n257), .A0(n431), .A1(n55), .Z(\cceip_ob_tlv[2][42] ));
Q_AN02 U818 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[43]), .Z(n432));
Q_MX02 U819 ( .S(n257), .A0(n432), .A1(n56), .Z(\cceip_ob_tlv[2][43] ));
Q_AN02 U820 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[44]), .Z(n433));
Q_MX02 U821 ( .S(n257), .A0(n433), .A1(n57), .Z(\cceip_ob_tlv[2][44] ));
Q_AN02 U822 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[45]), .Z(n434));
Q_MX02 U823 ( .S(n257), .A0(n434), .A1(n58), .Z(\cceip_ob_tlv[2][45] ));
Q_AN02 U824 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[46]), .Z(n435));
Q_MX02 U825 ( .S(n257), .A0(n435), .A1(n59), .Z(\cceip_ob_tlv[2][46] ));
Q_AN02 U826 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[47]), .Z(n436));
Q_MX02 U827 ( .S(n257), .A0(n436), .A1(n60), .Z(\cceip_ob_tlv[2][47] ));
Q_AN02 U828 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[48]), .Z(n437));
Q_MX02 U829 ( .S(n257), .A0(n437), .A1(n61), .Z(\cceip_ob_tlv[2][48] ));
Q_AN02 U830 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[49]), .Z(n438));
Q_MX02 U831 ( .S(n257), .A0(n438), .A1(n62), .Z(\cceip_ob_tlv[2][49] ));
Q_AN02 U832 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[50]), .Z(n439));
Q_MX02 U833 ( .S(n257), .A0(n439), .A1(n63), .Z(\cceip_ob_tlv[2][50] ));
Q_AN02 U834 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[51]), .Z(n440));
Q_MX02 U835 ( .S(n257), .A0(n440), .A1(n64), .Z(\cceip_ob_tlv[2][51] ));
Q_AN02 U836 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[52]), .Z(n441));
Q_MX02 U837 ( .S(n257), .A0(n441), .A1(n65), .Z(\cceip_ob_tlv[2][52] ));
Q_AN02 U838 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[53]), .Z(n442));
Q_MX02 U839 ( .S(n257), .A0(n442), .A1(n66), .Z(\cceip_ob_tlv[2][53] ));
Q_AN02 U840 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[54]), .Z(n443));
Q_MX02 U841 ( .S(n257), .A0(n443), .A1(n67), .Z(\cceip_ob_tlv[2][54] ));
Q_AN02 U842 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[55]), .Z(n444));
Q_MX02 U843 ( .S(n257), .A0(n444), .A1(n68), .Z(\cceip_ob_tlv[2][55] ));
Q_AN02 U844 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[56]), .Z(n445));
Q_MX02 U845 ( .S(n257), .A0(n445), .A1(n69), .Z(\cceip_ob_tlv[2][56] ));
Q_AN02 U846 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[57]), .Z(n446));
Q_MX02 U847 ( .S(n257), .A0(n446), .A1(n70), .Z(\cceip_ob_tlv[2][57] ));
Q_AN02 U848 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[58]), .Z(n447));
Q_MX02 U849 ( .S(n257), .A0(n447), .A1(n71), .Z(\cceip_ob_tlv[2][58] ));
Q_AN02 U850 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[59]), .Z(n448));
Q_MX02 U851 ( .S(n257), .A0(n448), .A1(n72), .Z(\cceip_ob_tlv[2][59] ));
Q_AN02 U852 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[60]), .Z(n449));
Q_MX02 U853 ( .S(n257), .A0(n449), .A1(n73), .Z(\cceip_ob_tlv[2][60] ));
Q_AN02 U854 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[61]), .Z(n450));
Q_MX02 U855 ( .S(n257), .A0(n450), .A1(n74), .Z(\cceip_ob_tlv[2][61] ));
Q_AN02 U856 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[62]), .Z(n451));
Q_MX02 U857 ( .S(n257), .A0(n451), .A1(n75), .Z(\cceip_ob_tlv[2][62] ));
Q_AN02 U858 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[63]), .Z(n452));
Q_MX02 U859 ( .S(n257), .A0(n452), .A1(n76), .Z(\cceip_ob_tlv[2][63] ));
Q_AN02 U860 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[64]), .Z(\cceip_ob_tlv[2][64] ));
Q_AN02 U861 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[65]), .Z(\cceip_ob_tlv[2][65] ));
Q_AN02 U862 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[66]), .Z(\cceip_ob_tlv[2][66] ));
Q_AN02 U863 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[67]), .Z(\cceip_ob_tlv[2][67] ));
Q_AN02 U864 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[68]), .Z(\cceip_ob_tlv[2][68] ));
Q_AN02 U865 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[69]), .Z(\cceip_ob_tlv[2][69] ));
Q_AN02 U866 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[70]), .Z(\cceip_ob_tlv[2][70] ));
Q_AN02 U867 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[71]), .Z(\cceip_ob_tlv[2][71] ));
Q_AN02 U868 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[72]), .Z(\cceip_ob_tlv[2][72] ));
Q_AN02 U869 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[73]), .Z(\cceip_ob_tlv[2][73] ));
Q_AN02 U870 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[74]), .Z(\cceip_ob_tlv[2][74] ));
Q_AN02 U871 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[75]), .Z(\cceip_ob_tlv[2][75] ));
Q_AN02 U872 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[76]), .Z(\cceip_ob_tlv[2][76] ));
Q_AN02 U873 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[77]), .Z(\cceip_ob_tlv[2][77] ));
Q_AN02 U874 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[78]), .Z(\cceip_ob_tlv[2][78] ));
Q_AN02 U875 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[79]), .Z(\cceip_ob_tlv[2][79] ));
Q_AN02 U876 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[80]), .Z(\cceip_ob_tlv[2][80] ));
Q_AN02 U877 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[82]), .Z(\cceip_ob_tlv[2][81] ));
Q_AN02 U878 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[83]), .Z(\cceip_ob_tlv[2][83] ));
Q_AN02 U879 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[84]), .Z(\cceip_ob_tlv[2][84] ));
Q_AN02 U880 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[85]), .Z(\cceip_ob_tlv[2][85] ));
Q_AN02 U881 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[86]), .Z(\cceip_ob_tlv[2][86] ));
Q_AN02 U882 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[87]), .Z(\cceip_ob_tlv[2][87] ));
Q_AN02 U883 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[88]), .Z(\cceip_ob_tlv[2][88] ));
Q_AN02 U884 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[89]), .Z(\cceip_ob_tlv[2][89] ));
Q_AN02 U885 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[90]), .Z(\cceip_ob_tlv[2][90] ));
Q_AN02 U886 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[91]), .Z(\cceip_ob_tlv[2][91] ));
Q_AN02 U887 ( .A0(\cceip_ob_tlv[2][92] ), .A1(encrypt_out[105]), .Z(\cceip_ob_tlv[2][105] ));
Q_AN02 U888 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[0]), .Z(n453));
Q_MX02 U889 ( .S(n258), .A0(n453), .A1(n13), .Z(\cceip_ob_tlv[3][0] ));
Q_AN02 U890 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[1]), .Z(n454));
Q_MX02 U891 ( .S(n258), .A0(n454), .A1(n14), .Z(\cceip_ob_tlv[3][1] ));
Q_AN02 U892 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[2]), .Z(n455));
Q_MX02 U893 ( .S(n258), .A0(n455), .A1(n15), .Z(\cceip_ob_tlv[3][2] ));
Q_AN02 U894 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[3]), .Z(n456));
Q_MX02 U895 ( .S(n258), .A0(n456), .A1(n16), .Z(\cceip_ob_tlv[3][3] ));
Q_AN02 U896 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[4]), .Z(n457));
Q_MX02 U897 ( .S(n258), .A0(n457), .A1(n17), .Z(\cceip_ob_tlv[3][4] ));
Q_AN02 U898 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[5]), .Z(n458));
Q_MX02 U899 ( .S(n258), .A0(n458), .A1(n18), .Z(\cceip_ob_tlv[3][5] ));
Q_AN02 U900 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[6]), .Z(n459));
Q_MX02 U901 ( .S(n258), .A0(n459), .A1(n19), .Z(\cceip_ob_tlv[3][6] ));
Q_AN02 U902 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[7]), .Z(n460));
Q_MX02 U903 ( .S(n258), .A0(n460), .A1(n20), .Z(\cceip_ob_tlv[3][7] ));
Q_AN02 U904 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[8]), .Z(n461));
Q_MX02 U905 ( .S(n258), .A0(n461), .A1(n21), .Z(\cceip_ob_tlv[3][8] ));
Q_AN02 U906 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[9]), .Z(n462));
Q_MX02 U907 ( .S(n258), .A0(n462), .A1(n22), .Z(\cceip_ob_tlv[3][9] ));
Q_AN02 U908 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[10]), .Z(n463));
Q_MX02 U909 ( .S(n258), .A0(n463), .A1(n23), .Z(\cceip_ob_tlv[3][10] ));
Q_AN02 U910 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[11]), .Z(n464));
Q_MX02 U911 ( .S(n258), .A0(n464), .A1(n24), .Z(\cceip_ob_tlv[3][11] ));
Q_AN02 U912 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[12]), .Z(n465));
Q_MX02 U913 ( .S(n258), .A0(n465), .A1(n25), .Z(\cceip_ob_tlv[3][12] ));
Q_AN02 U914 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[13]), .Z(n466));
Q_MX02 U915 ( .S(n258), .A0(n466), .A1(n26), .Z(\cceip_ob_tlv[3][13] ));
Q_AN02 U916 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[14]), .Z(n467));
Q_MX02 U917 ( .S(n258), .A0(n467), .A1(n27), .Z(\cceip_ob_tlv[3][14] ));
Q_AN02 U918 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[15]), .Z(n468));
Q_MX02 U919 ( .S(n258), .A0(n468), .A1(n28), .Z(\cceip_ob_tlv[3][15] ));
Q_AN02 U920 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[16]), .Z(n469));
Q_MX02 U921 ( .S(n258), .A0(n469), .A1(n29), .Z(\cceip_ob_tlv[3][16] ));
Q_AN02 U922 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[17]), .Z(n470));
Q_MX02 U923 ( .S(n258), .A0(n470), .A1(n30), .Z(\cceip_ob_tlv[3][17] ));
Q_AN02 U924 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[18]), .Z(n471));
Q_MX02 U925 ( .S(n258), .A0(n471), .A1(n31), .Z(\cceip_ob_tlv[3][18] ));
Q_AN02 U926 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[19]), .Z(n472));
Q_MX02 U927 ( .S(n258), .A0(n472), .A1(n32), .Z(\cceip_ob_tlv[3][19] ));
Q_AN02 U928 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[20]), .Z(n473));
Q_MX02 U929 ( .S(n258), .A0(n473), .A1(n33), .Z(\cceip_ob_tlv[3][20] ));
Q_AN02 U930 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[21]), .Z(n474));
Q_MX02 U931 ( .S(n258), .A0(n474), .A1(n34), .Z(\cceip_ob_tlv[3][21] ));
Q_AN02 U932 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[22]), .Z(n475));
Q_MX02 U933 ( .S(n258), .A0(n475), .A1(n35), .Z(\cceip_ob_tlv[3][22] ));
Q_AN02 U934 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[23]), .Z(n476));
Q_MX02 U935 ( .S(n258), .A0(n476), .A1(n36), .Z(\cceip_ob_tlv[3][23] ));
Q_AN02 U936 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[24]), .Z(n477));
Q_MX02 U937 ( .S(n258), .A0(n477), .A1(n37), .Z(\cceip_ob_tlv[3][24] ));
Q_AN02 U938 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[25]), .Z(n478));
Q_MX02 U939 ( .S(n258), .A0(n478), .A1(n38), .Z(\cceip_ob_tlv[3][25] ));
Q_AN02 U940 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[26]), .Z(n479));
Q_MX02 U941 ( .S(n258), .A0(n479), .A1(n39), .Z(\cceip_ob_tlv[3][26] ));
Q_AN02 U942 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[27]), .Z(n480));
Q_MX02 U943 ( .S(n258), .A0(n480), .A1(n40), .Z(\cceip_ob_tlv[3][27] ));
Q_AN02 U944 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[28]), .Z(n481));
Q_MX02 U945 ( .S(n258), .A0(n481), .A1(n41), .Z(\cceip_ob_tlv[3][28] ));
Q_AN02 U946 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[29]), .Z(n482));
Q_MX02 U947 ( .S(n258), .A0(n482), .A1(n42), .Z(\cceip_ob_tlv[3][29] ));
Q_AN02 U948 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[30]), .Z(n483));
Q_MX02 U949 ( .S(n258), .A0(n483), .A1(n43), .Z(\cceip_ob_tlv[3][30] ));
Q_AN02 U950 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[31]), .Z(n484));
Q_MX02 U951 ( .S(n258), .A0(n484), .A1(n44), .Z(\cceip_ob_tlv[3][31] ));
Q_AN02 U952 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[32]), .Z(n485));
Q_MX02 U953 ( .S(n258), .A0(n485), .A1(n45), .Z(\cceip_ob_tlv[3][32] ));
Q_AN02 U954 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[33]), .Z(n486));
Q_MX02 U955 ( .S(n258), .A0(n486), .A1(n46), .Z(\cceip_ob_tlv[3][33] ));
Q_AN02 U956 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[34]), .Z(n487));
Q_MX02 U957 ( .S(n258), .A0(n487), .A1(n47), .Z(\cceip_ob_tlv[3][34] ));
Q_AN02 U958 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[35]), .Z(n488));
Q_MX02 U959 ( .S(n258), .A0(n488), .A1(n48), .Z(\cceip_ob_tlv[3][35] ));
Q_AN02 U960 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[36]), .Z(n489));
Q_MX02 U961 ( .S(n258), .A0(n489), .A1(n49), .Z(\cceip_ob_tlv[3][36] ));
Q_AN02 U962 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[37]), .Z(n490));
Q_MX02 U963 ( .S(n258), .A0(n490), .A1(n50), .Z(\cceip_ob_tlv[3][37] ));
Q_AN02 U964 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[38]), .Z(n491));
Q_MX02 U965 ( .S(n258), .A0(n491), .A1(n51), .Z(\cceip_ob_tlv[3][38] ));
Q_AN02 U966 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[39]), .Z(n492));
Q_MX02 U967 ( .S(n258), .A0(n492), .A1(n52), .Z(\cceip_ob_tlv[3][39] ));
Q_AN02 U968 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[40]), .Z(n493));
Q_MX02 U969 ( .S(n258), .A0(n493), .A1(n53), .Z(\cceip_ob_tlv[3][40] ));
Q_AN02 U970 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[41]), .Z(n494));
Q_MX02 U971 ( .S(n258), .A0(n494), .A1(n54), .Z(\cceip_ob_tlv[3][41] ));
Q_AN02 U972 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[42]), .Z(n495));
Q_MX02 U973 ( .S(n258), .A0(n495), .A1(n55), .Z(\cceip_ob_tlv[3][42] ));
Q_AN02 U974 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[43]), .Z(n496));
Q_MX02 U975 ( .S(n258), .A0(n496), .A1(n56), .Z(\cceip_ob_tlv[3][43] ));
Q_AN02 U976 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[44]), .Z(n497));
Q_MX02 U977 ( .S(n258), .A0(n497), .A1(n57), .Z(\cceip_ob_tlv[3][44] ));
Q_AN02 U978 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[45]), .Z(n498));
Q_MX02 U979 ( .S(n258), .A0(n498), .A1(n58), .Z(\cceip_ob_tlv[3][45] ));
Q_AN02 U980 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[46]), .Z(n499));
Q_MX02 U981 ( .S(n258), .A0(n499), .A1(n59), .Z(\cceip_ob_tlv[3][46] ));
Q_AN02 U982 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[47]), .Z(n500));
Q_MX02 U983 ( .S(n258), .A0(n500), .A1(n60), .Z(\cceip_ob_tlv[3][47] ));
Q_AN02 U984 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[48]), .Z(n501));
Q_MX02 U985 ( .S(n258), .A0(n501), .A1(n61), .Z(\cceip_ob_tlv[3][48] ));
Q_AN02 U986 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[49]), .Z(n502));
Q_MX02 U987 ( .S(n258), .A0(n502), .A1(n62), .Z(\cceip_ob_tlv[3][49] ));
Q_AN02 U988 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[50]), .Z(n503));
Q_MX02 U989 ( .S(n258), .A0(n503), .A1(n63), .Z(\cceip_ob_tlv[3][50] ));
Q_AN02 U990 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[51]), .Z(n504));
Q_MX02 U991 ( .S(n258), .A0(n504), .A1(n64), .Z(\cceip_ob_tlv[3][51] ));
Q_AN02 U992 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[52]), .Z(n505));
Q_MX02 U993 ( .S(n258), .A0(n505), .A1(n65), .Z(\cceip_ob_tlv[3][52] ));
Q_AN02 U994 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[53]), .Z(n506));
Q_MX02 U995 ( .S(n258), .A0(n506), .A1(n66), .Z(\cceip_ob_tlv[3][53] ));
Q_AN02 U996 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[54]), .Z(n507));
Q_MX02 U997 ( .S(n258), .A0(n507), .A1(n67), .Z(\cceip_ob_tlv[3][54] ));
Q_AN02 U998 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[55]), .Z(n508));
Q_MX02 U999 ( .S(n258), .A0(n508), .A1(n68), .Z(\cceip_ob_tlv[3][55] ));
Q_AN02 U1000 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[56]), .Z(n509));
Q_MX02 U1001 ( .S(n258), .A0(n509), .A1(n69), .Z(\cceip_ob_tlv[3][56] ));
Q_AN02 U1002 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[57]), .Z(n510));
Q_MX02 U1003 ( .S(n258), .A0(n510), .A1(n70), .Z(\cceip_ob_tlv[3][57] ));
Q_AN02 U1004 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[58]), .Z(n511));
Q_MX02 U1005 ( .S(n258), .A0(n511), .A1(n71), .Z(\cceip_ob_tlv[3][58] ));
Q_AN02 U1006 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[59]), .Z(n512));
Q_MX02 U1007 ( .S(n258), .A0(n512), .A1(n72), .Z(\cceip_ob_tlv[3][59] ));
Q_AN02 U1008 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[60]), .Z(n513));
Q_MX02 U1009 ( .S(n258), .A0(n513), .A1(n73), .Z(\cceip_ob_tlv[3][60] ));
Q_AN02 U1010 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[61]), .Z(n514));
Q_MX02 U1011 ( .S(n258), .A0(n514), .A1(n74), .Z(\cceip_ob_tlv[3][61] ));
Q_AN02 U1012 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[62]), .Z(n515));
Q_MX02 U1013 ( .S(n258), .A0(n515), .A1(n75), .Z(\cceip_ob_tlv[3][62] ));
Q_AN02 U1014 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[63]), .Z(n516));
Q_MX02 U1015 ( .S(n258), .A0(n516), .A1(n76), .Z(\cceip_ob_tlv[3][63] ));
Q_AN02 U1016 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[64]), .Z(\cceip_ob_tlv[3][64] ));
Q_AN02 U1017 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[65]), .Z(\cceip_ob_tlv[3][65] ));
Q_AN02 U1018 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[66]), .Z(\cceip_ob_tlv[3][66] ));
Q_AN02 U1019 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[67]), .Z(\cceip_ob_tlv[3][67] ));
Q_AN02 U1020 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[68]), .Z(\cceip_ob_tlv[3][68] ));
Q_AN02 U1021 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[69]), .Z(\cceip_ob_tlv[3][69] ));
Q_AN02 U1022 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[70]), .Z(\cceip_ob_tlv[3][70] ));
Q_AN02 U1023 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[71]), .Z(\cceip_ob_tlv[3][71] ));
Q_AN02 U1024 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[72]), .Z(\cceip_ob_tlv[3][72] ));
Q_AN02 U1025 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[73]), .Z(\cceip_ob_tlv[3][73] ));
Q_AN02 U1026 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[74]), .Z(\cceip_ob_tlv[3][74] ));
Q_AN02 U1027 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[75]), .Z(\cceip_ob_tlv[3][75] ));
Q_AN02 U1028 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[76]), .Z(\cceip_ob_tlv[3][76] ));
Q_AN02 U1029 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[77]), .Z(\cceip_ob_tlv[3][77] ));
Q_AN02 U1030 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[78]), .Z(\cceip_ob_tlv[3][78] ));
Q_AN02 U1031 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[79]), .Z(\cceip_ob_tlv[3][79] ));
Q_AN02 U1032 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[80]), .Z(\cceip_ob_tlv[3][80] ));
Q_AN02 U1033 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[82]), .Z(\cceip_ob_tlv[3][81] ));
Q_AN02 U1034 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[83]), .Z(\cceip_ob_tlv[3][83] ));
Q_AN02 U1035 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[84]), .Z(\cceip_ob_tlv[3][84] ));
Q_AN02 U1036 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[85]), .Z(\cceip_ob_tlv[3][85] ));
Q_AN02 U1037 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[86]), .Z(\cceip_ob_tlv[3][86] ));
Q_AN02 U1038 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[87]), .Z(\cceip_ob_tlv[3][87] ));
Q_AN02 U1039 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[88]), .Z(\cceip_ob_tlv[3][88] ));
Q_AN02 U1040 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[89]), .Z(\cceip_ob_tlv[3][89] ));
Q_AN02 U1041 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[90]), .Z(\cceip_ob_tlv[3][90] ));
Q_AN02 U1042 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[91]), .Z(\cceip_ob_tlv[3][91] ));
Q_AN02 U1043 ( .A0(\cceip_ob_tlv[3][92] ), .A1(encrypt_out[105]), .Z(\cceip_ob_tlv[3][105] ));
Q_FDP4EP tlv_miscmp_REG  ( .CK(clk), .CE(n247), .R(n518), .D(n11), .Q(tlv_miscmp));
Q_INV U1045 ( .A(rst_n), .Z(n518));
Q_FDP4EP \_zy_sva_brcm_cceip_4_cpass_REG[0] ( .CK(clk), .CE(n10), .R(n324), .D(n517), .Q(_zy_sva_brcm_cceip_4_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_cceip_4_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n324), .D(n517), .Q(_zy_sva_brcm_cceip_4_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_cceip_3_cpass_REG[0] ( .CK(clk), .CE(n9), .R(n324), .D(n517), .Q(_zy_sva_brcm_cceip_3_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_cceip_3_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n324), .D(n517), .Q(_zy_sva_brcm_cceip_3_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_cceip_2_cpass_REG[0] ( .CK(clk), .CE(n8), .R(n324), .D(n517), .Q(_zy_sva_brcm_cceip_2_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_cceip_2_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n324), .D(n517), .Q(_zy_sva_brcm_cceip_2_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_cceip_1_cpass_REG[0] ( .CK(clk), .CE(n7), .R(n324), .D(n517), .Q(_zy_sva_brcm_cceip_1_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_cceip_1_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n324), .D(n517), .Q(_zy_sva_brcm_cceip_1_ccheck[0]));
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m1 "cceip_ob_tlv (2,0) 1 105 0 3 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_NON_CMM "1"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "\cceip_ob_tlv%s.ordern  1 12 0 3 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m2 "\cceip_ob_tlv%s.typen  1 7 0 3 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m3 "\cceip_ob_tlv%s.tid  1 0 0 3 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m4 "\cceip_ob_tlv%s.tstrb  1 7 0 3 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m5 "\cceip_ob_tlv%s.tuser  1 7 0 3 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m6 "\cceip_ob_tlv%s.tdata  1 63 0 3 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m7 "\cceip_encrypt_ob_tlv.ordern  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m8 "\cceip_encrypt_ob_tlv.typen  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m9 "\cceip_encrypt_ob_tlv.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m10 "\cceip_encrypt_ob_tlv.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m11 "\cceip_encrypt_ob_tlv.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m12 "\cceip_encrypt_ob_tlv.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m13 "\cceip_validate_ob_tlv.ordern  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m14 "\cceip_validate_ob_tlv.typen  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m15 "\cceip_validate_ob_tlv.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m16 "\cceip_validate_ob_tlv.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m17 "\cceip_validate_ob_tlv.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m18 "\cceip_validate_ob_tlv.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m19 "\encrypt_out.ordern  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m20 "\encrypt_out.typen  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m21 "\encrypt_out.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m22 "\encrypt_out.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m23 "\encrypt_out.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m24 "\encrypt_out.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m25 "\validate_out.ordern  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m26 "\validate_out.typen  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m27 "\validate_out.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m28 "\validate_out.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m29 "\validate_out.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m30 "\validate_out.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m31 "\key_tlv_w0.tlv_bip2  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m32 "\key_tlv_w0.resv0  (1,0) 1 18 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m33 "\key_tlv_w0.tlv_frame_num  (1,0) 1 10 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m34 "\key_tlv_w0.resv1  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m35 "\key_tlv_w0.tlv_eng_id  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m36 "\key_tlv_w0.tlv_seq_num  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m37 "\key_tlv_w0.tlv_len  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m38 "\key_tlv_w0.tlv_type  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "38"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r1 "cceip_ob_tlv%s 10 \cceip_ob_tlv%s.insert  \cceip_ob_tlv%s.ordern  \cceip_ob_tlv%s.typen  \cceip_ob_tlv%s.sot  \cceip_ob_tlv%s.eot  \cceip_ob_tlv%s.tlast  \cceip_ob_tlv%s.tid  \cceip_ob_tlv%s.tstrb  \cceip_ob_tlv%s.tuser  \cceip_ob_tlv%s.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r2 "cceip_encrypt_ob_tlv 10 \cceip_encrypt_ob_tlv.insert  \cceip_encrypt_ob_tlv.ordern  \cceip_encrypt_ob_tlv.typen  \cceip_encrypt_ob_tlv.sot  \cceip_encrypt_ob_tlv.eot  \cceip_encrypt_ob_tlv.tlast  \cceip_encrypt_ob_tlv.tid  \cceip_encrypt_ob_tlv.tstrb  \cceip_encrypt_ob_tlv.tuser  \cceip_encrypt_ob_tlv.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r3 "cceip_validate_ob_tlv 10 \cceip_validate_ob_tlv.insert  \cceip_validate_ob_tlv.ordern  \cceip_validate_ob_tlv.typen  \cceip_validate_ob_tlv.sot  \cceip_validate_ob_tlv.eot  \cceip_validate_ob_tlv.tlast  \cceip_validate_ob_tlv.tid  \cceip_validate_ob_tlv.tstrb  \cceip_validate_ob_tlv.tuser  \cceip_validate_ob_tlv.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r4 "encrypt_out 10 \encrypt_out.insert  \encrypt_out.ordern  \encrypt_out.typen  \encrypt_out.sot  \encrypt_out.eot  \encrypt_out.tlast  \encrypt_out.tid  \encrypt_out.tstrb  \encrypt_out.tuser  \encrypt_out.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r5 "validate_out 10 \validate_out.insert  \validate_out.ordern  \validate_out.typen  \validate_out.sot  \validate_out.eot  \validate_out.tlast  \validate_out.tid  \validate_out.tstrb  \validate_out.tuser  \validate_out.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r6 "key_tlv_w0 8 \key_tlv_w0.tlv_bip2  \key_tlv_w0.resv0  \key_tlv_w0.tlv_frame_num  \key_tlv_w0.resv1  \key_tlv_w0.tlv_eng_id  \key_tlv_w0.tlv_seq_num  \key_tlv_w0.tlv_len  \key_tlv_w0.tlv_type "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_NUM "6"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_0 "-1 engine 0 3 "
// pragma CVASTRPROP MODULE HDLICE PROP_RANOFF TRUE
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "engine[3]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "engine[2]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "engine[1]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "engine[0]"
endmodule
