library ieee, quickturn ;
use ieee.std_logic_1164.all ;
use quickturn.verilog.all ;
entity ixcEcmHoldOtb is
  attribute _2_state_: integer;
  attribute upf_always_on : integer;
  attribute upf_always_on of ixcEcmHoldOtb: entity is 1 ;
  attribute _2_state_ of ixcEcmHoldOtb: entity is 1 ;
end ixcEcmHoldOtb ;
