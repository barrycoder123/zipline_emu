architecture module of ixc_gfifo_bind_12_2 is

begin
end module;
