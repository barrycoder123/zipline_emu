architecture module of cr_kme_tlv_parser is
  -- quickturn multiple_driver_resolution
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "key_type[0]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "key_type[1]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "key_type[2]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "key_type[3]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "key_type[4]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "key_type[5]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "key_type[6]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "key_type[7]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "key_type[8]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "key_type[9]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "key_type[10]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "key_type[11]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "key_type[12]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "key_type[13]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[0]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[0].dek_op[0]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[0].dek_op[0].dak_op[0]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[0].dek_op[0].dak_op[1]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[0].dek_op[1]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[0].dek_op[1].dak_op[0]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[0].dek_op[1].dak_op[1]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[1]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[1].dek_op[0]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[1].dek_op[0].dak_op[0]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[1].dek_op[0].dak_op[1]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[1].dek_op[1]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[1].dek_op[1].dak_op[0]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[1].dek_op[1].dak_op[1]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[2]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[2].dek_op[0]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[2].dek_op[0].dak_op[0]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[2].dek_op[0].dak_op[1]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[2].dek_op[1]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[2].dek_op[1].dak_op[0]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[2].dek_op[1].dak_op[1]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[3]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[3].dek_op[0]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[3].dek_op[0].dak_op[0]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[3].dek_op[0].dak_op[1]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[3].dek_op[1]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[3].dek_op[1].dak_op[0]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[3].dek_op[1].dak_op[1]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "key_type_enc_dek[7]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "key_type_enc_dek[8]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "key_type_enc_dek_dak[10]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "key_type_enc_dek_dak[11]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "key_type_enc_dek_dak[12]"
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate "key_type_enc_dek_dak[13]"
  -- quickturn CVASTRPROP MODULE HDLICE PROP_RANOFF TRUE
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate_0 "-1 key_type 0 13 "
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate_1 "-1 kdf_mode 0 3 "
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate_2 "1 dek_op 0 1 "
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate_3 "2 dak_op 0 1 "
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate_4 "-1 key_type_enc_dek 7 8 "
  -- quickturn CVASTRPROP MODULE HDLICE cva_for_generate_5 "-1 key_type_enc_dek_dak 10 13 "
  component ixc_assign
    generic (
      W : integer := 1
    ) ;
    port (
      L : out std_logic_vector((W - 1) downto 0) ;
    R : in std_logic_vector((W - 1) downto 0) := (others => 'X') ) ;
  end component ;

  component cr_kme_fifo_xcm58
    generic (
      DATA_SIZE : integer := 71 ;
      FIFO_DEPTH : integer := 2 ;
      OVERRIDE_EN : integer := 0 ;
      STALL_AT : integer := 0
    ) ;
    port (
      fifo_in_stall : out std_logic ;
      fifo_out : out std_logic_vector(70 downto 0) ;
      fifo_out_valid : out std_logic ;
      fifo_overflow : out std_logic ;
      fifo_underflow : out std_logic ;
      clk : in std_logic := 'X' ;
      rst_n : in std_logic := 'X' ;
      fifo_in : in std_logic_vector(70 downto 0) := (others => 'X') ;
      fifo_in_valid : in std_logic := 'X' ;
      fifo_out_ack : in std_logic := 'X' ;
    fifo_in_stall_override : in std_logic := 'X' ) ;
  end component ;

  component ixc_sample_logic
    generic (
      WIDTH : integer := 1 ;
      RD_TYPE : integer := 0 ;
      subtype StateType is std_logic ;
      type DUMMY2 is array(integer range <>) of std_logic
    ) ;
    port (
      sv : out DUMMY2((WIDTH - 1) downto 0) ;
    v : in DUMMY2((WIDTH - 1) downto 0) ) ;
  end component ;

  type $_axi4s_dp_rdy_t is
  record
    tready : std_logic ;
  end record ;
  subtype axi4s_dp_rdy_t is $_axi4s_dp_rdy_t std_logic_vector(0 downto 0) ;
  type $_rbus_in_t is
  record
    addr : std_logic_vector(19 downto 0) ;
    wr_strb : std_logic ;
    wr_data : std_logic_vector(31 downto 0) ;
    rd_strb : std_logic ;
  end record ;
  subtype rbus_in_t is $_rbus_in_t std_logic_vector(53 downto 0) ;
  type $_rbus_out_t is
  record
    rd_data : std_logic_vector(31 downto 0) ;
    ack : std_logic ;
    err_ack : std_logic ;
  end record ;
  subtype rbus_out_t is $_rbus_out_t std_logic_vector(33 downto 0) ;
  type $_rbus_ring_t is
  record
    addr : std_logic_vector(19 downto 0) ;
    wr_strb : std_logic ;
    wr_data : std_logic_vector(31 downto 0) ;
    rd_strb : std_logic ;
    rd_data : std_logic_vector(31 downto 0) ;
    ack : std_logic ;
    err_ack : std_logic ;
  end record ;
  subtype rbus_ring_t is $_rbus_ring_t std_logic_vector(87 downto 0) ;
  type $_kme_rbus_ring_t is
  record
    addr : std_logic_vector(15 downto 0) ;
    wr_strb : std_logic ;
    wr_data : std_logic_vector(31 downto 0) ;
    rd_strb : std_logic ;
    rd_data : std_logic_vector(31 downto 0) ;
    ack : std_logic ;
    err_ack : std_logic ;
  end record ;
  subtype kme_rbus_ring_t is $_kme_rbus_ring_t std_logic_vector(83 downto 0) ;
  type $_im_desc_t is
  record
    eob : std_logic ;
    bytes_vld : std_logic_vector(7 downto 0) ;
    im_meta : std_logic_vector(22 downto 0) ;
  end record ;
  subtype im_desc_t is $_im_desc_t std_logic_vector(31 downto 0) ;
  type $_im_data_t is
  record
    data : std_logic_vector(63 downto 0) ;
  end record ;
  subtype im_data_t is $_im_data_t std_logic_vector(63 downto 0) ;
  type $_im_din_t is
  record
    data : im_data_t ;
    desc : im_desc_t ;
  end record ;
  subtype im_din_t is $_im_din_t std_logic_vector(95 downto 0) ;
  type $_im_available_t is
  record
    bank_hi : std_logic ;
    bank_lo : std_logic ;
  end record ;
  subtype im_available_t is $_im_available_t std_logic_vector(1 downto 0) ;
  type $_im_consumed_t is
  record
    bank_hi : std_logic ;
    bank_lo : std_logic ;
  end record ;
  subtype im_consumed_t is $_im_consumed_t std_logic_vector(1 downto 0) ;
  type $_frame_latency_if_bus_t is
  record
    valid : std_logic ;
    seq_num : std_logic_vector(7 downto 0) ;
  end record ;
  subtype frame_latency_if_bus_t is $_frame_latency_if_bus_t std_logic_vector(8
   downto 0) ;
  type $_sched_update_if_bus_t is
  record
    valid : std_logic ;
    rqe_sched_handle : std_logic_vector(15 downto 0) ;
    last : std_logic ;
    tlv_frame_num : std_logic_vector(10 downto 0) ;
    tlv_eng_id : std_logic_vector(3 downto 0) ;
    tlv_seq_num : std_logic_vector(7 downto 0) ;
    bytes_in : std_logic_vector(23 downto 0) ;
    bytes_out : std_logic_vector(23 downto 0) ;
    basis : std_logic_vector(23 downto 0) ;
  end record ;
  subtype sched_update_if_bus_t is $_sched_update_if_bus_t std_logic_vector(112
   downto 0) ;
  type $_tlvp_if_bus_t is
  record
    insert : std_logic ;
    ordern : std_logic_vector(12 downto 0) ;
    typen : tlv_types_e ;
    sot : std_logic ;
    eot : std_logic ;
    tlast : std_logic ;
    tid : std_logic_vector(0 downto 0) ;
    tstrb : std_logic_vector(7 downto 0) ;
    tuser : std_logic_vector(7 downto 0) ;
    tdata : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlvp_if_bus_t is $_tlvp_if_bus_t std_logic_vector(105 downto 0) ;
  type $_lz_symbol_bus_t is
  record
    framing : std_logic_vector(3 downto 0) ;
    data0 : std_logic_vector(7 downto 0) ;
    data1 : std_logic_vector(7 downto 0) ;
    data2 : std_logic_vector(7 downto 0) ;
    data3 : std_logic_vector(7 downto 0) ;
    backref : std_logic ;
    backref_type : std_logic ;
    backref_lane : std_logic_vector(1 downto 0) ;
    offset_msb : std_logic_vector(7 downto 0) ;
    length : std_logic_vector(15 downto 0) ;
  end record ;
  subtype lz_symbol_bus_t is $_lz_symbol_bus_t std_logic_vector(63 downto 0) ;
  type $_tlv_word_0_t is
  record
    tlv_bip2 : std_logic_vector(1 downto 0) ;
    resv0 : std_logic_vector(18 downto 0) ;
    tlv_frame_num : std_logic_vector(10 downto 0) ;
    resv1 : std_logic_vector(3 downto 0) ;
    tlv_eng_id : std_logic_vector(3 downto 0) ;
    tlv_seq_num : std_logic_vector(7 downto 0) ;
    tlv_len : std_logic_vector(7 downto 0) ;
    tlv_type : tlv_types_e ;
  end record ;
  subtype tlv_word_0_t is $_tlv_word_0_t std_logic_vector(63 downto 0) ;
  type $_tlv_rqe_word_0_t is
  record
    tlv_bip2 : std_logic_vector(1 downto 0) ;
    no_data : std_logic ;
    aux_frmd_crc : std_logic ;
    frame_size : rqe_frame_size_e ;
    vf_valid : std_logic ;
    trace : rqe_trace_e ;
    unused : std_logic_vector(10 downto 0) ;
    tlv_frame_num : std_logic_vector(10 downto 0) ;
    resv0 : std_logic_vector(3 downto 0) ;
    tlv_eng_id : std_logic_vector(3 downto 0) ;
    tlv_seq_num : std_logic_vector(7 downto 0) ;
    tlv_len : std_logic_vector(7 downto 0) ;
    tlv_type : tlv_types_e ;
  end record ;
  subtype tlv_rqe_word_0_t is $_tlv_rqe_word_0_t std_logic_vector(63 downto 0) ;
  type $_tlv_data_word_0_t is
  record
    tlv_bip2 : std_logic_vector(1 downto 0) ;
    last_of_command : std_logic ;
    resv0 : std_logic_vector(15 downto 0) ;
    coding : frmd_coding_e ;
    tlv_frame_num : std_logic_vector(10 downto 0) ;
    resv1 : std_logic_vector(3 downto 0) ;
    tlv_eng_id : std_logic_vector(3 downto 0) ;
    tlv_seq_num : std_logic_vector(7 downto 0) ;
    tlv_len : std_logic_vector(7 downto 0) ;
    tlv_type : tlv_types_e ;
  end record ;
  subtype tlv_data_word_0_t is $_tlv_data_word_0_t std_logic_vector(63 downto 0)
   ;
  type $_tlv_rqe_word_1_t is
  record
    pf_number : std_logic_vector(3 downto 0) ;
    vf_number : std_logic_vector(11 downto 0) ;
    scheduler_handle : std_logic_vector(15 downto 0) ;
    src_data_len : std_logic_vector(31 downto 0) ;
  end record ;
  subtype tlv_rqe_word_1_t is $_tlv_rqe_word_1_t std_logic_vector(63 downto 0) ;
  type $_cmd_debug_t is
  record
    tlvp_corrupt : tlvp_corrupt_e ;
    cmd_mode : cmd_mode_e ;
    module_id : std_logic_vector(4 downto 0) ;
    cmd_type : cmd_type_e ;
    tlv_num : std_logic_vector(4 downto 0) ;
    byte_num : std_logic_vector(9 downto 0) ;
    byte_msk : std_logic_vector(7 downto 0) ;
  end record ;
  subtype cmd_debug_t is $_cmd_debug_t std_logic_vector(31 downto 0) ;
  type $_bp_debug_t is
  record
    rsvd : std_logic_vector(0 downto 0) ;
    on_count : std_logic_vector(10 downto 0) ;
    off_count : std_logic_vector(10 downto 0) ;
  end record ;
  subtype bp_debug_t is $_bp_debug_t std_logic_vector(22 downto 0) ;
  type $_tlv_cmd_word_1_t is
  record
    debug : cmd_debug_t ;
    trace : std_logic ;
    dst_guid_present : std_logic ;
    frmd_out_type : std_logic_vector(6 downto 0) ;
    md_op : cmd_md_op_e ;
    md_type : cmd_md_type_e ;
    frmd_in_type : std_logic_vector(6 downto 0) ;
    frmd_in_aux : std_logic_vector(5 downto 0) ;
    frmd_crc_in : cmd_frmd_crc_in_e ;
    src_guid_present : cmd_guid_present_e ;
    compound_cmd_frm_size : cmd_compound_cmd_frm_size_e ;
  end record ;
  subtype tlv_cmd_word_1_t is $_tlv_cmd_word_1_t std_logic_vector(63 downto 0) ;
  type $_tlv_cmd_word_2_t is
  record
    rsvd2 : std_logic ;
    key_type : aux_key_type_e ;
    rsvd1 : std_logic_vector(1 downto 0) ;
    cipher_pad : cmd_cipher_pad_e ;
    iv_op : cmd_iv_op_e ;
    aad_len : std_logic_vector(7 downto 0) ;
    cipher_op : cmd_cipher_op_e ;
    auth_op : cmd_auth_op_e ;
    raw_auth_op : cmd_auth_op_e ;
    rsvd0 : std_logic_vector(7 downto 0) ;
    chu_comp_thrsh : cmd_chu_comp_thrsh_e ;
    xp10_crc_mode : cmd_xp10_crc_mode_e ;
    xp10_user_prefix_size : std_logic_vector(5 downto 0) ;
    xp10_prefix_mode : cmd_xp10_prefix_mode_e ;
    lz77_max_symb_len : cmd_lz77_max_symb_len_e ;
    lz77_min_match_len : cmd_lz77_min_match_len_e ;
    lz77_dly_match_win : cmd_lz77_dly_match_win_e ;
    lz77_win_size : cmd_lz77_win_size_e ;
    comp_mode : cmd_comp_mode_e ;
  end record ;
  subtype tlv_cmd_word_2_t is $_tlv_cmd_word_2_t std_logic_vector(63 downto 0) ;
  type $_tlv_key_word1_t is
  record
    guid : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_key_word1_t is $_tlv_key_word1_t std_logic_vector(63 downto 0) ;
  type $_tlv_key_word2_t is
  record
    guid : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_key_word2_t is $_tlv_key_word2_t std_logic_vector(63 downto 0) ;
  type $_tlv_key_word3_t is
  record
    guid : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_key_word3_t is $_tlv_key_word3_t std_logic_vector(63 downto 0) ;
  type $_tlv_key_word4_t is
  record
    guid : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_key_word4_t is $_tlv_key_word4_t std_logic_vector(63 downto 0) ;
  type $_tlv_key_word5_t is
  record
    ivtweak : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_key_word5_t is $_tlv_key_word5_t std_logic_vector(63 downto 0) ;
  type $_tlv_key_word6_t is
  record
    ivtweak : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_key_word6_t is $_tlv_key_word6_t std_logic_vector(63 downto 0) ;
  type $_tlv_key_word7_t is
  record
    dek : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_key_word7_t is $_tlv_key_word7_t std_logic_vector(63 downto 0) ;
  type $_tlv_key_word8_t is
  record
    dek : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_key_word8_t is $_tlv_key_word8_t std_logic_vector(63 downto 0) ;
  type $_tlv_key_word9_t is
  record
    dek : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_key_word9_t is $_tlv_key_word9_t std_logic_vector(63 downto 0) ;
  type $_tlv_key_word10_t is
  record
    dek : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_key_word10_t is $_tlv_key_word10_t std_logic_vector(63 downto 0) ;
  type $_tlv_key_word11_t is
  record
    dek : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_key_word11_t is $_tlv_key_word11_t std_logic_vector(63 downto 0) ;
  type $_tlv_key_word12_t is
  record
    dek : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_key_word12_t is $_tlv_key_word12_t std_logic_vector(63 downto 0) ;
  type $_tlv_key_word13_t is
  record
    dek : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_key_word13_t is $_tlv_key_word13_t std_logic_vector(63 downto 0) ;
  type $_tlv_key_word14_t is
  record
    dek : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_key_word14_t is $_tlv_key_word14_t std_logic_vector(63 downto 0) ;
  type $_tlv_key_word15_t is
  record
    dak : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_key_word15_t is $_tlv_key_word15_t std_logic_vector(63 downto 0) ;
  type $_tlv_key_word16_t is
  record
    dak : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_key_word16_t is $_tlv_key_word16_t std_logic_vector(63 downto 0) ;
  type $_tlv_key_word17_t is
  record
    dak : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_key_word17_t is $_tlv_key_word17_t std_logic_vector(63 downto 0) ;
  type $_tlv_key_word18_t is
  record
    dak : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_key_word18_t is $_tlv_key_word18_t std_logic_vector(63 downto 0) ;
  type $_tlv_key_word19_t is
  record
    rsvd : std_logic_vector(55 downto 0) ;
    kme_errors : zipline_error_e ;
  end record ;
  subtype tlv_key_word19_t is $_tlv_key_word19_t std_logic_vector(63 downto 0) ;
  type $_tlv_key_word20_t is
  record
    rsvd : std_logic_vector(31 downto 0) ;
    crc32 : std_logic_vector(31 downto 0) ;
  end record ;
  subtype tlv_key_word20_t is $_tlv_key_word20_t std_logic_vector(63 downto 0) ;
  type $_tlv_phd_word1_t is
  record
    rsvd : std_logic_vector(63 downto 6) ;
    xp10_prefix_sel : std_logic_vector(5 downto 0) ;
  end record ;
  subtype tlv_phd_word1_t is $_tlv_phd_word1_t std_logic_vector(63 downto 0) ;
  type $_tlv_pfd_word0_t is
  record
    tlv_bip2 : std_logic_vector(1 downto 0) ;
    resv0 : std_logic_vector(11 downto 0) ;
    prefix_src : std_logic ;
    xp10_prefix_sel : std_logic_vector(5 downto 0) ;
    tlv_frame_num : std_logic_vector(10 downto 0) ;
    resv1 : std_logic_vector(3 downto 0) ;
    tlv_eng_id : std_logic_vector(3 downto 0) ;
    tlv_seq_num : std_logic_vector(7 downto 0) ;
    tlv_len : std_logic_vector(7 downto 0) ;
    tlv_type : tlv_types_e ;
  end record ;
  subtype tlv_pfd_word0_t is $_tlv_pfd_word0_t std_logic_vector(63 downto 0) ;
  type $_tlv_pfd_word1_t is
  record
    rsvd : std_logic_vector(63 downto 6) ;
    xp10_prefix_sel : std_logic_vector(5 downto 0) ;
  end record ;
  subtype tlv_pfd_word1_t is $_tlv_pfd_word1_t std_logic_vector(63 downto 0) ;
  type $_tlv_guid_word1_t is
  record
    guid : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_guid_word1_t is $_tlv_guid_word1_t std_logic_vector(63 downto 0) ;
  type $_tlv_guid_word2_t is
  record
    guid : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_guid_word2_t is $_tlv_guid_word2_t std_logic_vector(63 downto 0) ;
  type $_tlv_guid_word3_t is
  record
    guid : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_guid_word3_t is $_tlv_guid_word3_t std_logic_vector(63 downto 0) ;
  type $_tlv_guid_word4_t is
  record
    guid : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_guid_word4_t is $_tlv_guid_word4_t std_logic_vector(63 downto 0) ;
  type $_tlv_ftr_word0_t is
  record
    tlv_bip2 : std_logic_vector(1 downto 0) ;
    rsvd3 : std_logic_vector(1 downto 0) ;
    gen_frmd_out_type : std_logic_vector(7 downto 0) ;
    rsvd2 : std_logic_vector(1 downto 0) ;
    raw_data_mac_size : frmd_mac_size_e ;
    enc_cmp_data_mac_size : frmd_mac_size_e ;
    coding : frmd_coding_e ;
    rsvd1 : std_logic ;
    tlv_frame_num : std_logic_vector(10 downto 0) ;
    rsvd0 : std_logic_vector(3 downto 0) ;
    tlv_eng_id : std_logic_vector(3 downto 0) ;
    tlv_seq_num : std_logic_vector(7 downto 0) ;
    tlv_len : std_logic_vector(7 downto 0) ;
    tlv_type : tlv_types_e ;
  end record ;
  subtype tlv_ftr_word0_t is $_tlv_ftr_word0_t std_logic_vector(63 downto 0) ;
  type $_tlv_ftr_word1_t is
  record
    raw_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_ftr_word1_t is $_tlv_ftr_word1_t std_logic_vector(63 downto 0) ;
  type $_tlv_ftr_word2_t is
  record
    raw_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_ftr_word2_t is $_tlv_ftr_word2_t std_logic_vector(63 downto 0) ;
  type $_tlv_ftr_word3_t is
  record
    raw_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_ftr_word3_t is $_tlv_ftr_word3_t std_logic_vector(63 downto 0) ;
  type $_tlv_ftr_word4_t is
  record
    raw_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_ftr_word4_t is $_tlv_ftr_word4_t std_logic_vector(63 downto 0) ;
  type $_tlv_ftr_word5_t is
  record
    raw_data_cksum : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_ftr_word5_t is $_tlv_ftr_word5_t std_logic_vector(63 downto 0) ;
  type $_tlv_ftr_word6_t is
  record
    raw_data_cksum_protocol : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_ftr_word6_t is $_tlv_ftr_word6_t std_logic_vector(63 downto 0) ;
  type $_tlv_ftr_word7_t is
  record
    enc_cmp_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_ftr_word7_t is $_tlv_ftr_word7_t std_logic_vector(63 downto 0) ;
  type $_tlv_ftr_word8_t is
  record
    enc_cmp_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_ftr_word8_t is $_tlv_ftr_word8_t std_logic_vector(63 downto 0) ;
  type $_tlv_ftr_word9_t is
  record
    enc_cmp_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_ftr_word9_t is $_tlv_ftr_word9_t std_logic_vector(63 downto 0) ;
  type $_tlv_ftr_word10_t is
  record
    enc_cmp_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_ftr_word10_t is $_tlv_ftr_word10_t std_logic_vector(63 downto 0) ;
  type $_tlv_ftr_word11_t is
  record
    enc_cmp_data_cksum : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_ftr_word11_t is $_tlv_ftr_word11_t std_logic_vector(63 downto 0) ;
  type $_tlv_ftr_word12_t is
  record
    nvme_raw_cksum_crc16t : std_logic_vector(15 downto 0) ;
    bytes_in : std_logic_vector(23 downto 0) ;
    bytes_out : std_logic_vector(23 downto 0) ;
  end record ;
  subtype tlv_ftr_word12_t is $_tlv_ftr_word12_t std_logic_vector(63 downto 0) ;
  type $_tlv_ftr_word13_t is
  record
    rsvd1 : std_logic_vector(19 downto 0) ;
    compressed_length : std_logic_vector(23 downto 0) ;
    error_code : zipline_error_e ;
    rsvd0 : std_logic ;
    errored_frame_number : std_logic_vector(10 downto 0) ;
  end record ;
  subtype tlv_ftr_word13_t is $_tlv_ftr_word13_t std_logic_vector(63 downto 0) ;
  type $_tlv_ftr_guid_word0_t is
  record
    guid : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_ftr_guid_word0_t is $_tlv_ftr_guid_word0_t std_logic_vector(63
   downto 0) ;
  type $_tlv_ftr_guid_word1_t is
  record
    guid : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_ftr_guid_word1_t is $_tlv_ftr_guid_word1_t std_logic_vector(63
   downto 0) ;
  type $_tlv_ftr_guid_word2_t is
  record
    guid : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_ftr_guid_word2_t is $_tlv_ftr_guid_word2_t std_logic_vector(63
   downto 0) ;
  type $_tlv_ftr_guid_word3_t is
  record
    guid : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_ftr_guid_word3_t is $_tlv_ftr_guid_word3_t std_logic_vector(63
   downto 0) ;
  type $_tlv_ftr_iv_word0_t is
  record
    rsvd : std_logic_vector(31 downto 0) ;
    iv : std_logic_vector(31 downto 0) ;
  end record ;
  subtype tlv_ftr_iv_word0_t is $_tlv_ftr_iv_word0_t std_logic_vector(63 downto
   0) ;
  type $_tlv_ftr_iv_word1_t is
  record
    iv : std_logic_vector(63 downto 0) ;
  end record ;
  subtype tlv_ftr_iv_word1_t is $_tlv_ftr_iv_word1_t std_logic_vector(63 downto
   0) ;
  type $_tlv_stats_word1_t is
  record
    rsvd1 : std_logic_vector(7 downto 0) ;
    bytes_in : std_logic_vector(23 downto 0) ;
    rsvd0 : std_logic_vector(7 downto 0) ;
    bytes_out : std_logic_vector(23 downto 0) ;
  end record ;
  subtype tlv_stats_word1_t is $_tlv_stats_word1_t std_logic_vector(63 downto 0)
   ;
  type $_tlv_stats_word2_t is
  record
    rsvd1 : std_logic_vector(30 downto 0) ;
    frame_error : std_logic ;
    rsvd0 : std_logic_vector(7 downto 0) ;
    latency : std_logic_vector(23 downto 0) ;
  end record ;
  subtype tlv_stats_word2_t is $_tlv_stats_word2_t std_logic_vector(63 downto 0)
   ;
  type $_tlv_cqe_word1_t is
  record
    status_code : std_logic_vector(7 downto 0) ;
    do_not_resend : std_logic ;
    vf_valid : std_logic ;
    rsvd0 : std_logic_vector(1 downto 0) ;
    error_code : std_logic_vector(7 downto 0) ;
    errored_frame_number : std_logic_vector(11 downto 0) ;
    status_code_type : std_logic_vector(2 downto 0) ;
    stat_cts : std_logic_vector(12 downto 0) ;
    pf_number : std_logic_vector(3 downto 0) ;
    vf_number : std_logic_vector(11 downto 0) ;
  end record ;
  subtype tlv_cqe_word1_t is $_tlv_cqe_word1_t std_logic_vector(63 downto 0) ;
  type $_fmd_user_pi16_word1_t is
  record
    rsvd : std_logic_vector(47 downto 0) ;
    nvme_raw_cksum_crc16t : std_logic_vector(15 downto 0) ;
  end record ;
  subtype fmd_user_pi16_word1_t is $_fmd_user_pi16_word1_t std_logic_vector(63
   downto 0) ;
  type $_fmd_user_pi64_word1_t is
  record
    raw_data_cksum : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_user_pi64_word1_t is $_fmd_user_pi64_word1_t std_logic_vector(63
   downto 0) ;
  type $_fmd_user_vm_word1_t is
  record
    ivtweak : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_user_vm_word1_t is $_fmd_user_vm_word1_t std_logic_vector(63
   downto 0) ;
  type $_fmd_user_vm_word2_t is
  record
    ivtweak : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_user_vm_word2_t is $_fmd_user_vm_word2_t std_logic_vector(63
   downto 0) ;
  type $_fmd_user_vm_word3_t is
  record
    raw_data_cksum : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_user_vm_word3_t is $_fmd_user_vm_word3_t std_logic_vector(63
   downto 0) ;
  type $_fmd_user_vm_word4_t is
  record
    raw_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_user_vm_word4_t is $_fmd_user_vm_word4_t std_logic_vector(63
   downto 0) ;
  type $_fmd_user_vm_word5_t is
  record
    raw_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_user_vm_word5_t is $_fmd_user_vm_word5_t std_logic_vector(63
   downto 0) ;
  type $_fmd_user_vm_word6_t is
  record
    raw_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_user_vm_word6_t is $_fmd_user_vm_word6_t std_logic_vector(63
   downto 0) ;
  type $_fmd_user_vm_word7_t is
  record
    raw_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_user_vm_word7_t is $_fmd_user_vm_word7_t std_logic_vector(63
   downto 0) ;
  type $_fmd_int_app_word6_t is
  record
    rsvd : std_logic_vector(31 downto 0) ;
    rsvd0 : std_logic_vector(5 downto 0) ;
    coding : frmd_coding_e ;
    compressed_length : std_logic_vector(23 downto 0) ;
  end record ;
  subtype fmd_int_app_word6_t is $_fmd_int_app_word6_t std_logic_vector(63
   downto 0) ;
  type $_fmd_int_app_word1_t is
  record
    enc_cmp_data_cksum : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_app_word1_t is $_fmd_int_app_word1_t std_logic_vector(63
   downto 0) ;
  type $_fmd_int_app_word2_t is
  record
    enc_cmp_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_app_word2_t is $_fmd_int_app_word2_t std_logic_vector(63
   downto 0) ;
  type $_fmd_int_app_word3_t is
  record
    enc_cmp_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_app_word3_t is $_fmd_int_app_word3_t std_logic_vector(63
   downto 0) ;
  type $_fmd_int_app_word4_t is
  record
    ivtweak : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_app_word4_t is $_fmd_int_app_word4_t std_logic_vector(63
   downto 0) ;
  type $_fmd_int_app_word5_t is
  record
    rsvd : std_logic_vector(31 downto 0) ;
    ivtweak : std_logic_vector(31 downto 0) ;
  end record ;
  subtype fmd_int_app_word5_t is $_fmd_int_app_word5_t std_logic_vector(63
   downto 0) ;
  type $_fmd_int_sip_word3_t is
  record
    rsvd : std_logic_vector(31 downto 0) ;
    rsvd0 : std_logic_vector(5 downto 0) ;
    coding : frmd_coding_e ;
    compressed_length : std_logic_vector(23 downto 0) ;
  end record ;
  subtype fmd_int_sip_word3_t is $_fmd_int_sip_word3_t std_logic_vector(63
   downto 0) ;
  type $_fmd_int_sip_word1_t is
  record
    enc_cmp_data_cksum : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_sip_word1_t is $_fmd_int_sip_word1_t std_logic_vector(63
   downto 0) ;
  type $_fmd_int_sip_word2_t is
  record
    raw_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_sip_word2_t is $_fmd_int_sip_word2_t std_logic_vector(63
   downto 0) ;
  type $_fmd_int_lip_word6_t is
  record
    rsvd : std_logic_vector(31 downto 0) ;
    rsvd0 : std_logic_vector(5 downto 0) ;
    coding : frmd_coding_e ;
    compressed_length : std_logic_vector(23 downto 0) ;
  end record ;
  subtype fmd_int_lip_word6_t is $_fmd_int_lip_word6_t std_logic_vector(63
   downto 0) ;
  type $_fmd_int_lip_word1_t is
  record
    enc_cmp_data_cksum : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_lip_word1_t is $_fmd_int_lip_word1_t std_logic_vector(63
   downto 0) ;
  type $_fmd_int_lip_word2_t is
  record
    raw_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_lip_word2_t is $_fmd_int_lip_word2_t std_logic_vector(63
   downto 0) ;
  type $_fmd_int_lip_word3_t is
  record
    raw_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_lip_word3_t is $_fmd_int_lip_word3_t std_logic_vector(63
   downto 0) ;
  type $_fmd_int_lip_word4_t is
  record
    raw_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_lip_word4_t is $_fmd_int_lip_word4_t std_logic_vector(63
   downto 0) ;
  type $_fmd_int_lip_word5_t is
  record
    raw_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_lip_word5_t is $_fmd_int_lip_word5_t std_logic_vector(63
   downto 0) ;
  type $_fmd_int_vm_word12_t is
  record
    rsvd : std_logic_vector(31 downto 0) ;
    rsvd0 : std_logic_vector(5 downto 0) ;
    coding : frmd_coding_e ;
    compressed_length : std_logic_vector(23 downto 0) ;
  end record ;
  subtype fmd_int_vm_word12_t is $_fmd_int_vm_word12_t std_logic_vector(63
   downto 0) ;
  type $_fmd_int_vm_word1_t is
  record
    enc_cmp_data_cksum : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_vm_word1_t is $_fmd_int_vm_word1_t std_logic_vector(63 downto
   0) ;
  type $_fmd_int_vm_word2_t is
  record
    enc_cmp_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_vm_word2_t is $_fmd_int_vm_word2_t std_logic_vector(63 downto
   0) ;
  type $_fmd_int_vm_word3_t is
  record
    enc_cmp_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_vm_word3_t is $_fmd_int_vm_word3_t std_logic_vector(63 downto
   0) ;
  type $_fmd_int_vm_word4_t is
  record
    enc_cmp_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_vm_word4_t is $_fmd_int_vm_word4_t std_logic_vector(63 downto
   0) ;
  type $_fmd_int_vm_word5_t is
  record
    enc_cmp_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_vm_word5_t is $_fmd_int_vm_word5_t std_logic_vector(63 downto
   0) ;
  type $_fmd_int_vm_word6_t is
  record
    raw_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_vm_word6_t is $_fmd_int_vm_word6_t std_logic_vector(63 downto
   0) ;
  type $_fmd_int_vm_word7_t is
  record
    raw_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_vm_word7_t is $_fmd_int_vm_word7_t std_logic_vector(63 downto
   0) ;
  type $_fmd_int_vm_word8_t is
  record
    raw_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_vm_word8_t is $_fmd_int_vm_word8_t std_logic_vector(63 downto
   0) ;
  type $_fmd_int_vm_word9_t is
  record
    raw_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_vm_word9_t is $_fmd_int_vm_word9_t std_logic_vector(63 downto
   0) ;
  type $_fmd_int_vm_word10_t is
  record
    ivtweak : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_vm_word10_t is $_fmd_int_vm_word10_t std_logic_vector(63
   downto 0) ;
  type $_fmd_int_vm_word11_t is
  record
    ivtweak : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_vm_word11_t is $_fmd_int_vm_word11_t std_logic_vector(63
   downto 0) ;
  type $_fmd_int_vm_short_word9_t is
  record
    rsvd : std_logic_vector(31 downto 0) ;
    rsvd0 : std_logic_vector(5 downto 0) ;
    coding : frmd_coding_e ;
    compressed_length : std_logic_vector(23 downto 0) ;
  end record ;
  subtype fmd_int_vm_short_word9_t is $_fmd_int_vm_short_word9_t
   std_logic_vector(63 downto 0) ;
  type $_fmd_int_vm_short_word1_t is
  record
    enc_cmp_data_cksum : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_vm_short_word1_t is $_fmd_int_vm_short_word1_t
   std_logic_vector(63 downto 0) ;
  type $_fmd_int_vm_short_word2_t is
  record
    enc_cmp_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_vm_short_word2_t is $_fmd_int_vm_short_word2_t
   std_logic_vector(63 downto 0) ;
  type $_fmd_int_vm_short_word3_t is
  record
    enc_cmp_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_vm_short_word3_t is $_fmd_int_vm_short_word3_t
   std_logic_vector(63 downto 0) ;
  type $_fmd_int_vm_short_word4_t is
  record
    enc_cmp_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_vm_short_word4_t is $_fmd_int_vm_short_word4_t
   std_logic_vector(63 downto 0) ;
  type $_fmd_int_vm_short_word5_t is
  record
    enc_cmp_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_vm_short_word5_t is $_fmd_int_vm_short_word5_t
   std_logic_vector(63 downto 0) ;
  type $_fmd_int_vm_short_word6_t is
  record
    raw_data_mac : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_vm_short_word6_t is $_fmd_int_vm_short_word6_t
   std_logic_vector(63 downto 0) ;
  type $_fmd_int_vm_short_word7_t is
  record
    ivtweak : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_vm_short_word7_t is $_fmd_int_vm_short_word7_t
   std_logic_vector(63 downto 0) ;
  type $_fmd_int_vm_short_word8_t is
  record
    ivtweak : std_logic_vector(63 downto 0) ;
  end record ;
  subtype fmd_int_vm_short_word8_t is $_fmd_int_vm_short_word8_t
   std_logic_vector(63 downto 0) ;
  type $_s_sm_seq_id_intf is
  record
    predet_mem_mask : std_logic ;
    predet_mem_id : std_logic_vector(3 downto 0) ;
    comp_mode : cmd_comp_mode_e ;
    lz77_win_size : cmd_lz77_win_size_e ;
    lz77_min_match_len : cmd_lz77_min_match_len_e ;
    xp10_prefix_mode : cmd_xp10_prefix_mode_e ;
    xp10_user_prefix_size : std_logic_vector(5 downto 0) ;
    xp10_crc_mode : cmd_xp10_crc_mode_e ;
    chu_comp_thrsh : cmd_chu_comp_thrsh_e ;
    tid : std_logic_vector(0 downto 0) ;
    tuser : std_logic_vector(7 downto 0) ;
    raw_byte_count : std_logic_vector(23 downto 0) ;
    extra_bit_count : std_logic_vector(17 downto 0) ;
    blk_count : std_logic_vector(10 downto 0) ;
    blk_last : std_logic ;
    pdh_crc_err : std_logic ;
    raw_crc : std_logic_vector(63 downto 0) ;
  end record ;
  subtype s_sm_seq_id_intf is $_s_sm_seq_id_intf std_logic_vector(152 downto 0)
   ;
  type $_s_seq_id_type_intf is
  record
    comp_mode : cmd_comp_mode_e ;
    lz77_win_size : cmd_lz77_win_size_e ;
    xp10_prefix_mode : cmd_xp10_prefix_mode_e ;
  end record ;
  subtype s_seq_id_type_intf is $_s_seq_id_type_intf std_logic_vector(9 downto 0
  ) ;
  type $_counter_50_t is
  record
    count_part1 : std_logic_vector(17 downto 0) ;
    count_part0 : std_logic_vector(31 downto 0) ;
  end record ;
  subtype counter_50_t is $_counter_50_t std_logic_vector(49 downto 0) ;
  type $_cg_stats_t is
  record
    cqe_out : std_logic ;
    cqe_sys_err : std_logic ;
    cqe_err_sel : std_logic ;
    cqe_eng_err : std_logic ;
  end record ;
  subtype cg_stats_t is $_cg_stats_t std_logic_vector(3 downto 0) ;
  type $_osf_stats_t is
  record
    rsvd : std_logic_vector(59 downto 0) ;
    ob_stall : std_logic ;
    ob_sys_bp : std_logic ;
    pdt_fifo_stall : std_logic ;
    dat_fifo_stall : std_logic ;
  end record ;
  subtype osf_stats_t is $_osf_stats_t std_logic_vector(63 downto 0) ;
  type $_isf_stats_t is
  record
    rsvd : std_logic_vector(54 downto 0) ;
    aux_cmd_match3 : std_logic ;
    aux_cmd_match2 : std_logic ;
    aux_cmd_match1 : std_logic ;
    aux_cmd_match0 : std_logic ;
    ob_sys_bp : std_logic ;
    ib_sys_stall : std_logic ;
    ib_stall : std_logic ;
    ib_frame : std_logic ;
    ib_cmd : std_logic ;
  end record ;
  subtype isf_stats_t is $_isf_stats_t std_logic_vector(63 downto 0) ;
  type $_huf_comp_stats_t is
  record
    huff_comp_rsvd : std_logic_vector(9 downto 0) ;
    lz77_stall_stb : std_logic ;
    encrypt_stall_stb : std_logic ;
    byte_7_stb : std_logic ;
    byte_6_stb : std_logic ;
    byte_5_stb : std_logic ;
    byte_4_stb : std_logic ;
    byte_3_stb : std_logic ;
    byte_2_stb : std_logic ;
    byte_1_stb : std_logic ;
    byte_0_stb : std_logic ;
    pass_thru_frm_stb : std_logic ;
    df_frm_stb : std_logic ;
    df_blk_long_ret_stb : std_logic ;
    df_blk_shrt_ret_stb : std_logic ;
    df_blk_long_sim_stb : std_logic ;
    df_blk_shrt_sim_stb : std_logic ;
    df_blk_raw_stb : std_logic ;
    df_blk_enc_stb : std_logic ;
    chu4_cmd_stb : std_logic ;
    chu4_frm_long_pre_stb : std_logic ;
    chu4_frm_shrt_pre_stb : std_logic ;
    chu4_frm_long_ret_stb : std_logic ;
    chu4_frm_shrt_ret_stb : std_logic ;
    chu4_frm_long_sim_stb : std_logic ;
    chu4_frm_shrt_sim_stb : std_logic ;
    chu4_frm_enc_stb : std_logic ;
    chu4_frm_raw_stb : std_logic ;
    chu8_cmd_stb : std_logic ;
    chu8_frm_long_pre_stb : std_logic ;
    chu8_frm_shrt_pre_stb : std_logic ;
    chu8_frm_long_ret_stb : std_logic ;
    chu8_frm_shrt_ret_stb : std_logic ;
    chu8_frm_long_sim_stb : std_logic ;
    chu8_frm_shrt_sim_stb : std_logic ;
    chu8_frm_enc_stb : std_logic ;
    chu8_frm_raw_stb : std_logic ;
    xp10_frm_stb : std_logic ;
    xp10_blk_long_pre_stb : std_logic ;
    xp10_blk_shrt_pre_stb : std_logic ;
    xp10_blk_long_ret_stb : std_logic ;
    xp10_blk_shrt_ret_stb : std_logic ;
    xp10_blk_long_sim_stb : std_logic ;
    xp10_blk_shrt_sim_stb : std_logic ;
    xp10_blk_raw_stb : std_logic ;
    xp10_blk_enc_stb : std_logic ;
    xp9_blk_long_ret_stb : std_logic ;
    xp9_blk_shrt_ret_stb : std_logic ;
    xp9_blk_long_sim_stb : std_logic ;
    xp9_blk_shrt_sim_stb : std_logic ;
    xp9_frm_stb : std_logic ;
    xp9_frm_raw_stb : std_logic ;
    xp9_blk_enc_stb : std_logic ;
    long_map_err_stb : std_logic ;
    shrt_map_err_stb : std_logic ;
  end record ;
  subtype huf_comp_stats_t is $_huf_comp_stats_t std_logic_vector(63 downto 0) ;
  type $_crypto_stats_t is
  record
    unused : std_logic_vector(48 downto 0) ;
    cipher_aes_gcm : std_logic_vector(0 downto 0) ;
    cipher_aes_xts : std_logic_vector(0 downto 0) ;
    cipher_aes_xex : std_logic_vector(0 downto 0) ;
    cipher_nop : std_logic_vector(0 downto 0) ;
    auth_aes_gmac : std_logic_vector(0 downto 0) ;
    auth_sha256 : std_logic_vector(0 downto 0) ;
    auth_sha256_hmac : std_logic_vector(0 downto 0) ;
    auth_nop : std_logic_vector(0 downto 0) ;
    gcm_tag_fail : std_logic_vector(0 downto 0) ;
    gmac_tag_fail : std_logic_vector(0 downto 0) ;
    sha256_tag_fail : std_logic_vector(0 downto 0) ;
    hmac_sha256_tag_fail : std_logic_vector(0 downto 0) ;
    seq_id_mismatch : std_logic_vector(0 downto 0) ;
    eng_id_mismatch : std_logic_vector(0 downto 0) ;
    reserved : std_logic_vector(0 downto 0) ;
  end record ;
  subtype crypto_stats_t is $_crypto_stats_t std_logic_vector(63 downto 0) ;
  type $_aux_key_ctrl_t is
  record
    dak_key_op : aux_key_op_e ;
    dak_key_ref : std_logic_vector(13 downto 0) ;
    kdf_mode : aux_kdf_mode_e ;
    dek_key_op : aux_key_op_e ;
    dek_key_ref : std_logic_vector(13 downto 0) ;
  end record ;
  subtype aux_key_ctrl_t is $_aux_key_ctrl_t std_logic_vector(31 downto 0) ;
  type $_axi4s_su_dp_bus_t is
  record
    tvalid : std_logic ;
    tlast : std_logic ;
    tuser : std_logic_vector(1 downto 0) ;
    tdata : std_logic_vector(7 downto 0) ;
  end record ;
  subtype axi4s_su_dp_bus_t is $_axi4s_su_dp_bus_t std_logic_vector(11 downto 0)
   ;
  type $_generic_int_t is
  record
    tlvp_err : std_logic ;
    uncor_ecc_err : std_logic ;
    bimc_int : std_logic ;
  end record ;
  subtype generic_int_t is $_generic_int_t std_logic_vector(2 downto 0) ;
  type $_ecc_int_t is
  record
    uncor_ecc_err : std_logic ;
  end record ;
  subtype ecc_int_t is $_ecc_int_t std_logic_vector(0 downto 0) ;
  type $_tlvp_int_t is
  record
    tlvp_err : std_logic ;
  end record ;
  subtype tlvp_int_t is $_tlvp_int_t std_logic_vector(0 downto 0) ;
  type $_bimc_int_t is
  record
    bimc_err : std_logic ;
  end record ;
  subtype bimc_int_t is $_bimc_int_t std_logic_vector(0 downto 0) ;
  type $_crypto_int_t is
  record
    seed_expire : std_logic ;
    id_mismatch : std_logic ;
    tlvp_err : std_logic ;
    uncor_ecc_err : std_logic ;
  end record ;
  subtype crypto_int_t is $_crypto_int_t std_logic_vector(3 downto 0) ;
  type $_crypto_ckmic_int_t is
  record
    id_mismatch : std_logic ;
    tlvp_err : std_logic ;
  end record ;
  subtype crypto_ckmic_int_t is $_crypto_ckmic_int_t std_logic_vector(1 downto 0
  ) ;
  type $_osf_int_t is
  record
    tlvp_err : std_logic ;
    uncor_ecc_err : std_logic ;
  end record ;
  subtype osf_int_t is $_osf_int_t std_logic_vector(1 downto 0) ;
  type $_isf_int_t is
  record
    sys_stall : std_logic ;
    ovfl : std_logic ;
    prot_err : std_logic ;
    tlvp_int : std_logic ;
    uncor_ecc_err : std_logic ;
  end record ;
  subtype isf_int_t is $_isf_int_t std_logic_vector(4 downto 0) ;
  type $_prefix_attach_int_t is
  record
    tlvp_err : std_logic ;
    uncor_ecc_err : std_logic ;
  end record ;
  subtype prefix_attach_int_t is $_prefix_attach_int_t std_logic_vector(1 downto
   0) ;
  type $_ftr_error_t is
  record
    error_code : zipline_error_e ;
    errored_frame_number : std_logic_vector(10 downto 0) ;
  end record ;
  subtype ftr_error_t is $_ftr_error_t std_logic_vector(18 downto 0) ;
  type $_kim_entry_t is
  record
    valid : std_logic_vector(0 downto 0) ;
    label_index : std_logic_vector(2 downto 0) ;
    ckv_length : std_logic_vector(1 downto 0) ;
    ckv_pointer : std_logic_vector(14 downto 0) ;
    pf_num : std_logic_vector(3 downto 0) ;
    vf_num : std_logic_vector(11 downto 0) ;
    vf_valid : std_logic_vector(0 downto 0) ;
  end record ;
  subtype kim_entry_t is $_kim_entry_t std_logic_vector(37 downto 0) ;
  type $_label_t is
  record
    guid_size : std_logic_vector(0 downto 0) ;
    label_size : std_logic_vector(5 downto 0) ;
    DUMMY1 : std_logic_vector(255 downto 0) ;
    delimiter_valid : std_logic_vector(0 downto 0) ;
    delimiter : std_logic_vector(7 downto 0) ;
  end record ;
  subtype label_t is $_label_t std_logic_vector(271 downto 0) ;
  type $_kim_ckv_resp_t is
  record
    valid : std_logic_vector(0 downto 0) ;
    label_index : std_logic_vector(2 downto 0) ;
    pf_num : std_logic_vector(0 downto 0) ;
    vf_valid : std_logic_vector(0 downto 0) ;
    vf_num : std_logic_vector(8 downto 0) ;
    ckv_key : std_logic_vector(511 downto 0) ;
  end record ;
  subtype kim_ckv_resp_t is $_kim_ckv_resp_t std_logic_vector(526 downto 0) ;
  type $_kme_internal_word_0_t is
  record
    tlv_bip2 : std_logic_vector(1 downto 0) ;
    resv0 : std_logic_vector(12 downto 0) ;
    kdf_dek_iter : std_logic_vector(0 downto 0) ;
    keyless_algos : std_logic_vector(0 downto 0) ;
    needs_dek : std_logic_vector(0 downto 0) ;
    needs_dak : std_logic_vector(0 downto 0) ;
    key_type : aux_key_type_e ;
    tlv_frame_num : std_logic_vector(10 downto 0) ;
    tlv_eng_id : std_logic_vector(3 downto 0) ;
    tlv_seq_num : std_logic_vector(7 downto 0) ;
    tlv_len : std_logic_vector(7 downto 0) ;
    tlv_type : tlv_types_e ;
  end record ;
  subtype kme_internal_word_0_t is $_kme_internal_word_0_t std_logic_vector(63
   downto 0) ;
  type $_kme_internal_word_8_t is
  record
    dek_kim_entry : kim_entry_t ;
    unused : std_logic_vector(5 downto 0) ;
    missing_iv : std_logic_vector(0 downto 0) ;
    missing_guid : std_logic_vector(0 downto 0) ;
    validate_dek : std_logic_vector(0 downto 0) ;
    vf_valid : std_logic_vector(0 downto 0) ;
    pf_num : std_logic_vector(3 downto 0) ;
    vf_num : std_logic_vector(11 downto 0) ;
  end record ;
  subtype kme_internal_word_8_t is $_kme_internal_word_8_t std_logic_vector(63
   downto 0) ;
  type $_kme_internal_word_9_t is
  record
    dak_kim_entry : kim_entry_t ;
    unused : std_logic_vector(7 downto 0) ;
    validate_dak : std_logic_vector(0 downto 0) ;
    vf_valid : std_logic_vector(0 downto 0) ;
    pf_num : std_logic_vector(3 downto 0) ;
    vf_num : std_logic_vector(11 downto 0) ;
  end record ;
  subtype kme_internal_word_9_t is $_kme_internal_word_9_t std_logic_vector(63
   downto 0) ;
  type $_kme_internal_word_42_t is
  record
    corrupt_crc32 : std_logic_vector(0 downto 0) ;
    unused : std_logic_vector(46 downto 0) ;
    error_code : zipline_error_e ;
  end record ;
  subtype kme_internal_word_42_t is $_kme_internal_word_42_t std_logic_vector(55
   downto 0) ;
  type $_gcm_cmd_t is
  record
    key0 : std_logic_vector(255 downto 0) ;
    key1 : std_logic_vector(255 downto 0) ;
    iv : std_logic_vector(95 downto 0) ;
    op : gcm_op_e ;
  end record ;
  subtype gcm_cmd_t is $_gcm_cmd_t std_logic_vector(610 downto 0) ;
  type $_gcm_status_t is
  record
    tag_mismatch : std_logic_vector(0 downto 0) ;
  end record ;
  subtype gcm_status_t is $_gcm_status_t std_logic_vector(0 downto 0) ;
  type $_keyfilter_cmd_t is
  record
    combo_mode : std_logic_vector(0 downto 0) ;
  end record ;
  subtype keyfilter_cmd_t is $_keyfilter_cmd_t std_logic_vector(0 downto 0) ;
  type $_kdf_cmd_t is
  record
    kdf_dek_iter : std_logic_vector(0 downto 0) ;
    combo_mode : std_logic_vector(0 downto 0) ;
    dek_key_op : aux_key_op_e ;
    dak_key_op : aux_key_op_e ;
  end record ;
  subtype kdf_cmd_t is $_kdf_cmd_t std_logic_vector(3 downto 0) ;
  type $_kdfstream_cmd_t is
  record
    combo_mode : std_logic_vector(0 downto 0) ;
    skip : std_logic_vector(0 downto 0) ;
    guid : std_logic_vector(255 downto 0) ;
    label_index : std_logic_vector(2 downto 0) ;
    num_iter : std_logic_vector(1 downto 0) ;
  end record ;
  subtype kdfstream_cmd_t is $_kdfstream_cmd_t std_logic_vector(262 downto 0) ;
  type $_skip_control is
  record
    start : std_logic_vector(0 downto 0) ;
    partial : std_logic_vector(0 downto 0) ;
    endian_swap : std_logic_vector(0 downto 0) ;
    till : kme_internal_id ;
  end record ;
  subtype skip_control is $_skip_control std_logic_vector(6 downto 0) ;
  signal fifo_in_stall : std_logic ;
  signal stitcher_sot : std_logic ;
  signal stitcher_eot : std_logic ;
  signal DUMMY2 : std_logic ;
  signal DUMMY3 : std_logic_vector(0 to 70) ;
  signal DUMMY4 : std_logic_vector(0 to 70) ;
  signal _zy_simnet_dio_3 : std_logic ;
  signal _zy_simnet_dio_4 : std_logic ;
  signal DUMMY5 : std_logic_vector(0 to 70) ;
  signal DUMMY6 : std_logic ;
  signal _zy_simnet_cio_7 : std_logic ;
  signal _zy_sva_key_type0_line4_1_reset_or : std_logic ;
  signal _zy_sva_key_type0_line5a_2_reset_or : std_logic ;
  signal _zy_sva_key_type0_line5b_3_reset_or : std_logic ;
  signal _zy_sva_key_type1_line7a_4_reset_or : std_logic ;
  signal _zy_sva_key_type1_line7b_5_reset_or : std_logic ;
  signal _zy_sva_key_type1_line8a_6_reset_or : std_logic ;
  signal _zy_sva_key_type1_line8b_7_reset_or : std_logic ;
  signal _zy_sva_key_type1_line9_8_reset_or : std_logic ;
  signal _zy_sva_key_type1_line10_9_reset_or : std_logic ;
  signal _zy_sva_key_type1_line11a_10_reset_or : std_logic ;
  signal _zy_sva_key_type1_line11b_11_reset_or : std_logic ;
  signal _zy_sva_key_type1_line11c_12_reset_or : std_logic ;
  signal _zy_sva_key_type1_line11d_13_reset_or : std_logic ;
  signal _zy_sva_key_type1_line12a_14_reset_or : std_logic ;
  signal _zy_sva_key_type1_line12b_15_reset_or : std_logic ;
  signal _zy_sva_key_type9_line14_16_reset_or : std_logic ;
  signal _zy_sva_key_type9_line15_17_reset_or : std_logic ;
  signal _zy_sva_key_type9_line16a_18_reset_or : std_logic ;
  signal _zy_sva_key_type9_line16b_19_reset_or : std_logic ;
  signal _zy_sva_key_type9_line17a_20_reset_or : std_logic ;
  signal _zy_sva_key_type9_line17b_21_reset_or : std_logic ;
  signal _zy_sva_key_type9_line18a_22_reset_or : std_logic ;
  signal _zy_sva_key_type9_line18b_23_reset_or : std_logic ;
  signal _zy_sva_key_type9_line19a_24_reset_or : std_logic ;
  signal _zy_sva_key_type9_line19b_25_reset_or : std_logic ;
  signal _zy_sva_key_type9_line19c_26_reset_or : std_logic ;
  signal _zy_sva_key_type9_line19d_27_reset_or : std_logic ;
  signal _zy_sva_guid_miss_aux_cmd_0_28_reset_or : std_logic ;
  signal _zy_sva_guid_miss_aux_cmd_1_29_reset_or : std_logic ;
  signal _zy_sva_guid_miss_aux_cmd_2_30_reset_or : std_logic ;
  signal _zy_sva_guid_miss_aux_cmd_3_31_reset_or : std_logic ;
  signal _zy_sva_guid_miss_aux_cmd_iv_0_32_reset_or : std_logic ;
  signal _zy_sva_guid_miss_aux_cmd_iv_1_33_reset_or : std_logic ;
  signal _zy_sva_guid_miss_aux_cmd_iv_2_34_reset_or : std_logic ;
  signal _zy_sva_guid_miss_aux_cmd_iv_3_35_reset_or : std_logic ;
  signal _zy_sva_iv_miss_aux_cmd_0_36_reset_or : std_logic ;
  signal _zy_sva_iv_miss_aux_cmd_1_37_reset_or : std_logic ;
  signal _zy_sva_iv_miss_aux_cmd_guid_38_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_39_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_iv_40_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_guid_41_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_42_reset_or : std_logic ;
  signal _zy_sva_brcm_key_type_43_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_44_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_iv_45_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_guid_46_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_47_reset_or : std_logic ;
  signal _zy_sva_brcm_key_type_48_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_49_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_iv_50_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_guid_51_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_52_reset_or : std_logic ;
  signal _zy_sva_brcm_key_type_53_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_54_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_iv_55_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_guid_56_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_57_reset_or : std_logic ;
  signal _zy_sva_brcm_key_type_58_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_59_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_iv_60_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_guid_61_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_62_reset_or : std_logic ;
  signal _zy_sva_brcm_key_type_63_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_64_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_iv_65_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_guid_66_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_67_reset_or : std_logic ;
  signal _zy_sva_brcm_key_type_68_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_69_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_iv_70_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_guid_71_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_72_reset_or : std_logic ;
  signal _zy_sva_brcm_key_type_73_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_74_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_iv_75_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_guid_76_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_77_reset_or : std_logic ;
  signal _zy_sva_brcm_key_type_78_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_79_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_iv_80_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_guid_81_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_82_reset_or : std_logic ;
  signal _zy_sva_brcm_key_type_83_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_84_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_iv_85_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_guid_86_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_87_reset_or : std_logic ;
  signal _zy_sva_brcm_key_type_88_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_89_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_iv_90_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_guid_91_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_92_reset_or : std_logic ;
  signal _zy_sva_brcm_key_type_93_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_94_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_iv_95_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_guid_96_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_97_reset_or : std_logic ;
  signal _zy_sva_brcm_key_type_98_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_99_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_iv_100_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_guid_101_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_102_reset_or : std_logic ;
  signal _zy_sva_brcm_key_type_103_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_104_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_iv_105_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_guid_106_reset_or : std_logic ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_107_reset_or : std_logic ;
  signal _zy_sva_brcm_key_type_108_reset_or : std_logic ;
  signal _zy_sva_brcm_kdf_ops_109_reset_or : std_logic ;
  signal _zy_sva_brcm_kdf_ops_110_reset_or : std_logic ;
  signal _zy_sva_brcm_kdf_ops_111_reset_or : std_logic ;
  signal _zy_sva_brcm_kdf_ops_112_reset_or : std_logic ;
  signal _zy_sva_brcm_kdf_ops_113_reset_or : std_logic ;
  signal _zy_sva_brcm_kdf_ops_114_reset_or : std_logic ;
  signal _zy_sva_brcm_kdf_ops_115_reset_or : std_logic ;
  signal _zy_sva_brcm_kdf_ops_116_reset_or : std_logic ;
  signal _zy_sva_brcm_kdf_ops_117_reset_or : std_logic ;
  signal _zy_sva_brcm_kdf_ops_118_reset_or : std_logic ;
  signal _zy_sva_brcm_kdf_ops_119_reset_or : std_logic ;
  signal _zy_sva_brcm_kdf_ops_120_reset_or : std_logic ;
  signal _zy_sva_brcm_kdf_ops_121_reset_or : std_logic ;
  signal _zy_sva_brcm_kdf_ops_122_reset_or : std_logic ;
  signal _zy_sva_brcm_kdf_ops_123_reset_or : std_logic ;
  signal _zy_sva_brcm_kdf_ops_124_reset_or : std_logic ;
  signal _zy_sva_null_gcm_125_reset_or : std_logic ;
  signal _zy_sva_sha_gcm_126_reset_or : std_logic ;
  signal _zy_sva_null_xts_127_reset_or : std_logic ;
  signal _zy_sva_sha_xts_128_reset_or : std_logic ;
  signal _zy_sva_null_null_129_reset_or : std_logic ;
  signal _zy_sva_sha_null_130_reset_or : std_logic ;
  signal _zy_sva_hmac_gcm_131_reset_or : std_logic ;
  signal _zy_sva_hmac_xts_132_reset_or : std_logic ;
  signal _zy_sva_hmac_null_133_reset_or : std_logic ;
  signal _zy_sva_null_gcm_134_reset_or : std_logic ;
  signal _zy_sva_sha_gcm_135_reset_or : std_logic ;
  signal _zy_sva_null_xts_136_reset_or : std_logic ;
  signal _zy_sva_sha_xts_137_reset_or : std_logic ;
  signal _zy_sva_null_null_138_reset_or : std_logic ;
  signal _zy_sva_sha_null_139_reset_or : std_logic ;
  signal _zy_sva_hmac_gcm_140_reset_or : std_logic ;
  signal _zy_sva_hmac_xts_141_reset_or : std_logic ;
  signal _zy_sva_hmac_null_142_reset_or : std_logic ;
  signal _zy_sva_null_gcm_143_reset_or : std_logic ;
  signal _zy_sva_sha_gcm_144_reset_or : std_logic ;
  signal _zy_sva_null_xts_145_reset_or : std_logic ;
  signal _zy_sva_sha_xts_146_reset_or : std_logic ;
  signal _zy_sva_null_null_147_reset_or : std_logic ;
  signal _zy_sva_sha_null_148_reset_or : std_logic ;
  signal _zy_sva_hmac_gcm_149_reset_or : std_logic ;
  signal _zy_sva_hmac_xts_150_reset_or : std_logic ;
  signal _zy_sva_hmac_null_151_reset_or : std_logic ;
  signal _zy_sva_null_gcm_152_reset_or : std_logic ;
  signal _zy_sva_sha_gcm_153_reset_or : std_logic ;
  signal _zy_sva_null_xts_154_reset_or : std_logic ;
  signal _zy_sva_sha_xts_155_reset_or : std_logic ;
  signal _zy_sva_null_null_156_reset_or : std_logic ;
  signal _zy_sva_sha_null_157_reset_or : std_logic ;
  signal _zy_sva_hmac_gcm_158_reset_or : std_logic ;
  signal _zy_sva_hmac_xts_159_reset_or : std_logic ;
  signal _zy_sva_hmac_null_160_reset_or : std_logic ;
  signal _zy_sva_null_gcm_161_reset_or : std_logic ;
  signal _zy_sva_sha_gcm_162_reset_or : std_logic ;
  signal _zy_sva_null_xts_163_reset_or : std_logic ;
  signal _zy_sva_sha_xts_164_reset_or : std_logic ;
  signal _zy_sva_null_null_165_reset_or : std_logic ;
  signal _zy_sva_sha_null_166_reset_or : std_logic ;
  signal _zy_sva_hmac_gcm_167_reset_or : std_logic ;
  signal _zy_sva_hmac_xts_168_reset_or : std_logic ;
  signal _zy_sva_hmac_null_169_reset_or : std_logic ;
  signal _zy_sva_null_gcm_170_reset_or : std_logic ;
  signal _zy_sva_sha_gcm_171_reset_or : std_logic ;
  signal _zy_sva_null_xts_172_reset_or : std_logic ;
  signal _zy_sva_sha_xts_173_reset_or : std_logic ;
  signal _zy_sva_null_null_174_reset_or : std_logic ;
  signal _zy_sva_sha_null_175_reset_or : std_logic ;
  signal _zy_sva_hmac_gcm_176_reset_or : std_logic ;
  signal _zy_sva_hmac_xts_177_reset_or : std_logic ;
  signal _zy_sva_hmac_null_178_reset_or : std_logic ;
  signal _zy_sva_b0_t : std_logic ;
  signal _zy_sva_b1_t : std_logic ;
  signal _zy_sva_b2_t : std_logic ;
  signal _zy_sva_b3_t : std_logic ;
  signal _zy_sva_b4_t : std_logic ;
  signal _zy_sva_b5_t : std_logic ;
  signal _zy_sva_b6_t : std_logic ;
  signal _zy_sva_b7_t : std_logic ;
  signal _zy_sva_b8_t : std_logic ;
  signal _zy_sva_b9_t : std_logic ;
  signal _zy_sva_b10_t : std_logic ;
  signal _zy_sva_b11_t : std_logic ;
  signal _zy_sva_b12_t : std_logic ;
  signal _zy_sva_b13_t : std_logic ;
  signal _zy_sva_b14_t : std_logic ;
  signal _zy_sva_b15_t : std_logic ;
  signal _zy_sva_b16_t : std_logic ;
  signal _zy_sva_b17_t : std_logic ;
  signal _zy_sva_b18_t : std_logic ;
  signal _zy_sva_b19_t : std_logic ;
  signal _zy_sva_b20_t : std_logic ;
  signal _zy_sva_b21_t : std_logic ;
  signal _zy_sva_b22_t : std_logic ;
  signal _zy_sva_b23_t : std_logic ;
  signal _zy_sva_b24_t : std_logic ;
  signal _zy_sva_b25_t : std_logic ;
  signal _zy_sva_b26_t : std_logic ;
  signal _zy_sva_b27_t : std_logic ;
  signal _zy_sva_b28_t : std_logic ;
  signal _zy_sva_b29_t : std_logic ;
  signal _zy_sva_b30_t : std_logic ;
  signal _zy_sva_b31_t : std_logic ;
  signal _zy_sva_b32_t : std_logic ;
  signal _zy_sva_b33_t : std_logic ;
  signal _zy_sva_b34_t : std_logic ;
  signal _zy_sva_b35_t : std_logic ;
  signal _zy_sva_b36_t : std_logic ;
  signal _zy_sva_b37_t : std_logic ;
  signal _zy_sva_b38_t : std_logic ;
  signal _zy_sva_b39_t : std_logic ;
  signal _zy_sva_b40_t : std_logic ;
  signal _zy_sva_b41_t : std_logic ;
  signal _zy_sva_b42_t : std_logic ;
  signal _zy_sva_b43_t : std_logic ;
  signal _zy_sva_b44_t : std_logic ;
  signal _zy_sva_b45_t : std_logic ;
  signal _zy_sva_b46_t : std_logic ;
  signal _zy_sva_b47_t : std_logic ;
  signal _zy_sva_b48_t : std_logic ;
  signal _zy_sva_b49_t : std_logic ;
  signal _zy_sva_b50_t : std_logic ;
  signal _zy_sva_b51_t : std_logic ;
  signal _zy_sva_b52_t : std_logic ;
  signal _zy_sva_b53_t : std_logic ;
  signal _zy_sva_b54_t : std_logic ;
  signal _zy_sva_b55_t : std_logic ;
  signal _zy_sva_b56_t : std_logic ;
  signal _zy_sva_b57_t : std_logic ;
  signal _zy_sva_b58_t : std_logic ;
  signal _zy_sva_b59_t : std_logic ;
  signal _zy_sva_b60_t : std_logic ;
  signal _zy_sva_b61_t : std_logic ;
  signal _zy_sva_b62_t : std_logic ;
  signal _zy_sva_b63_t : std_logic ;
  signal _zy_sva_b64_t : std_logic ;
  signal _zy_sva_b65_t : std_logic ;
  signal _zy_sva_b66_t : std_logic ;
  signal _zy_sva_b67_t : std_logic ;
  signal _zy_sva_b68_t : std_logic ;
  signal _zy_sva_b69_t : std_logic ;
  signal _zy_sva_b70_t : std_logic ;
  signal _zy_sva_b71_t : std_logic ;
  signal _zy_sva_b72_t : std_logic ;
  signal _zy_sva_b73_t : std_logic ;
  signal _zy_sva_b74_t : std_logic ;
  signal _zy_sva_b75_t : std_logic ;
  signal _zy_sva_b76_t : std_logic ;
  signal _zy_sva_b77_t : std_logic ;
  signal _zy_sva_b78_t : std_logic ;
  signal _zy_sva_b79_t : std_logic ;
  signal _zy_sva_b80_t : std_logic ;
  signal _zy_sva_b81_t : std_logic ;
  signal _zy_sva_b82_t : std_logic ;
  signal _zy_sva_b83_t : std_logic ;
  signal _zy_sva_b84_t : std_logic ;
  signal _zy_sva_b85_t : std_logic ;
  signal _zy_sva_b86_t : std_logic ;
  signal _zy_sva_b87_t : std_logic ;
  signal _zy_sva_b88_t : std_logic ;
  signal _zy_sva_b89_t : std_logic ;
  signal _zy_sva_b90_t : std_logic ;
  signal _zy_sva_b91_t : std_logic ;
  signal _zy_sva_b92_t : std_logic ;
  signal _zy_sva_b93_t : std_logic ;
  signal _zy_sva_b94_t : std_logic ;
  signal _zy_sva_b95_t : std_logic ;
  signal _zy_sva_b96_t : std_logic ;
  signal _zy_sva_b97_t : std_logic ;
  signal _zy_sva_b98_t : std_logic ;
  signal _zy_sva_b99_t : std_logic ;
  signal _zy_sva_b100_t : std_logic ;
  signal _zy_sva_b101_t : std_logic ;
  signal _zy_sva_b102_t : std_logic ;
  signal _zy_sva_b103_t : std_logic ;
  signal _zy_sva_b104_t : std_logic ;
  signal _zy_sva_b105_t : std_logic ;
  signal _zy_sva_b106_t : std_logic ;
  signal _zy_sva_b107_t : std_logic ;
  signal _zy_sva_b108_t : std_logic ;
  signal _zy_sva_b109_t : std_logic ;
  signal _zy_sva_b110_t : std_logic ;
  signal _zy_sva_b111_t : std_logic ;
  signal _zy_sva_b112_t : std_logic ;
  signal _zy_sva_b113_t : std_logic ;
  signal _zy_sva_b114_t : std_logic ;
  signal _zy_sva_b115_t : std_logic ;
  signal _zy_sva_b116_t : std_logic ;
  signal _zy_sva_b117_t : std_logic ;
  signal _zy_sva_b118_t : std_logic ;
  signal _zy_sva_b119_t : std_logic ;
  signal _zy_sva_b120_t : std_logic ;
  signal _zy_sva_b121_t : std_logic ;
  signal _zy_sva_b122_t : std_logic ;
  signal _zy_sva_b123_t : std_logic ;
  signal _zy_sva_b124_t : std_logic ;
  signal _zy_sva_b125_t : std_logic ;
  signal _zy_sva_b126_t : std_logic ;
  signal _zy_sva_b127_t : std_logic ;
  signal _zy_sva_b128_t : std_logic ;
  signal _zy_sva_b129_t : std_logic ;
  signal _zy_sva_b130_t : std_logic ;
  signal _zy_sva_b131_t : std_logic ;
  signal _zy_sva_b132_t : std_logic ;
  signal _zy_sva_b133_t : std_logic ;
  signal _zy_sva_b134_t : std_logic ;
  signal _zy_sva_b135_t : std_logic ;
  signal _zy_sva_b136_t : std_logic ;
  signal _zy_sva_b137_t : std_logic ;
  signal _zy_sva_b138_t : std_logic ;
  signal _zy_sva_b139_t : std_logic ;
  signal _zy_sva_b140_t : std_logic ;
  signal _zy_sva_b141_t : std_logic ;
  signal _zy_sva_b142_t : std_logic ;
  signal _zy_sva_b143_t : std_logic ;
  signal _zy_sva_b144_t : std_logic ;
  signal _zy_sva_b145_t : std_logic ;
  signal _zy_sva_b146_t : std_logic ;
  signal _zy_sva_b147_t : std_logic ;
  signal _zy_sva_b148_t : std_logic ;
  signal _zy_sva_b149_t : std_logic ;
  signal _zy_sva_b150_t : std_logic ;
  signal _zy_sva_b151_t : std_logic ;
  signal _zy_sva_b152_t : std_logic ;
  signal _zy_sva_b153_t : std_logic ;
  signal _zy_sva_b154_t : std_logic ;
  signal _zy_sva_b155_t : std_logic ;
  signal _zy_sva_b156_t : std_logic ;
  signal _zy_sva_b157_t : std_logic ;
  signal _zy_sva_b158_t : std_logic ;
  signal _zy_sva_b159_t : std_logic ;
  signal _zy_sva_b160_t : std_logic ;
  signal _zy_sva_b161_t : std_logic ;
  signal _zy_sva_b162_t : std_logic ;
  signal _zy_sva_b163_t : std_logic ;
  signal _zy_sva_b164_t : std_logic ;
  signal _zy_sva_b165_t : std_logic ;
  signal _zy_sva_b166_t : std_logic ;
  signal _zy_sva_b167_t : std_logic ;
  signal _zy_sva_b168_t : std_logic ;
  signal _zy_sva_b169_t : std_logic ;
  signal _zy_sva_b170_t : std_logic ;
  signal _zy_sva_b171_t : std_logic ;
  signal _zy_sva_b172_t : std_logic ;
  signal _zy_sva_b173_t : std_logic ;
  signal _zy_sva_b174_t : std_logic ;
  signal _zy_sva_b175_t : std_logic ;
  signal _zy_sva_b176_t : std_logic ;
  signal _zy_sva_b177_t : std_logic ;
  signal fifo_in : kme_internal_t ;
  signal fifo_in_valid : std_logic ;
  signal key_blob_region : std_logic ;
  signal int_tlv_counter : std_logic_vector(5 downto 0) ;
  signal tlv_counter : std_logic_vector(4 downto 0) ;
  signal tlv_word0 : tlv_rqe_word_0_t ;
  signal tlv_word1 : tlv_rqe_word_1_t ;
  signal tlv_word2 : tlv_cmd_word_2_t ;
  signal nxt_fifo_in_id : kme_internal_id ;
  signal frame_word : tlv_cmd_word_1_t ;
  signal kme_internal_word0 : kme_internal_word_0_t ;
  signal nxt_kme_internal_word0 : kme_internal_word_0_t ;
  signal kme_internal_dek_kim_word : kme_internal_word_8_t ;
  signal nxt_kme_internal_dek_kim_word : kme_internal_word_8_t ;
  signal kme_internal_dak_kim_word : kme_internal_word_9_t ;
  signal nxt_kme_internal_dak_kim_word : kme_internal_word_9_t ;
  signal tlv_type : tlv_types_e ;
  signal nxt_tlv_type : tlv_types_e ;
  signal aux_key_type : aux_key_type_e ;
  signal nxt_aux_key_type : aux_key_type_e ;
  signal aux_iv_op : cmd_iv_op_e ;
  signal nxt_aux_iv_op : cmd_iv_op_e ;
  signal aux_cipher_op : cmd_cipher_op_e ;
  signal nxt_aux_cipher_op : cmd_cipher_op_e ;
  signal aux_auth_op : cmd_auth_op_e ;
  signal nxt_aux_auth_op : cmd_auth_op_e ;
  signal aux_raw_auth_op : cmd_auth_op_e ;
  signal nxt_aux_raw_auth_op : cmd_auth_op_e ;
  signal debug_cmd : cmd_debug_t ;
  signal nxt_debug_cmd : cmd_debug_t ;
  signal aux_key_header : aux_key_ctrl_t ;
  signal nxt_aux_key_header : aux_key_ctrl_t ;
  signal skip : skip_control ;
  signal nxt_skip : skip_control ;
  signal guid0 : std_logic_vector(63 downto 0) ;
  signal nxt_guid0 : std_logic_vector(63 downto 0) ;
  signal guid1 : std_logic_vector(63 downto 0) ;
  signal nxt_guid1 : std_logic_vector(63 downto 0) ;
  signal guid2 : std_logic_vector(63 downto 0) ;
  signal nxt_guid2 : std_logic_vector(63 downto 0) ;
  signal guid3 : std_logic_vector(63 downto 0) ;
  signal nxt_guid3 : std_logic_vector(63 downto 0) ;
  signal iv0 : std_logic_vector(63 downto 0) ;
  signal nxt_iv0 : std_logic_vector(63 downto 0) ;
  signal iv1 : std_logic_vector(63 downto 0) ;
  signal nxt_iv1 : std_logic_vector(63 downto 0) ;
  signal DUMMY7 : std_logic_vector(31 downto 0) ;
  signal nxt_buffer : std_logic_vector(31 downto 0) ;
  signal _zy_sva_key_type0_line4_1_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type0_line4_1_ccheck: signal is 1 ;
  signal _zy_sva_key_type0_line4_1_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type0_line4_1_cpass: signal is 1 ;
  signal _zy_sva_b0 : std_logic ;
  attribute _2_state_ of _zy_sva_b0: signal is 1 ;
  signal _zy_sva_key_type0_line5a_2_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type0_line5a_2_ccheck: signal is 1 ;
  signal _zy_sva_key_type0_line5a_2_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type0_line5a_2_cpass: signal is 1 ;
  signal _zy_sva_b1 : std_logic ;
  attribute _2_state_ of _zy_sva_b1: signal is 1 ;
  signal _zy_sva_key_type0_line5b_3_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type0_line5b_3_ccheck: signal is 1 ;
  signal _zy_sva_key_type0_line5b_3_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type0_line5b_3_cpass: signal is 1 ;
  signal _zy_sva_b2 : std_logic ;
  attribute _2_state_ of _zy_sva_b2: signal is 1 ;
  signal _zy_sva_key_type1_line7a_4_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type1_line7a_4_ccheck: signal is 1 ;
  signal _zy_sva_key_type1_line7a_4_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type1_line7a_4_cpass: signal is 1 ;
  signal _zy_sva_b3 : std_logic ;
  attribute _2_state_ of _zy_sva_b3: signal is 1 ;
  signal _zy_sva_key_type1_line7b_5_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type1_line7b_5_ccheck: signal is 1 ;
  signal _zy_sva_key_type1_line7b_5_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type1_line7b_5_cpass: signal is 1 ;
  signal _zy_sva_b4 : std_logic ;
  attribute _2_state_ of _zy_sva_b4: signal is 1 ;
  signal _zy_sva_key_type1_line8a_6_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type1_line8a_6_ccheck: signal is 1 ;
  signal _zy_sva_key_type1_line8a_6_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type1_line8a_6_cpass: signal is 1 ;
  signal _zy_sva_b5 : std_logic ;
  attribute _2_state_ of _zy_sva_b5: signal is 1 ;
  signal _zy_sva_key_type1_line8b_7_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type1_line8b_7_ccheck: signal is 1 ;
  signal _zy_sva_key_type1_line8b_7_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type1_line8b_7_cpass: signal is 1 ;
  signal _zy_sva_b6 : std_logic ;
  attribute _2_state_ of _zy_sva_b6: signal is 1 ;
  signal _zy_sva_key_type1_line9_8_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type1_line9_8_ccheck: signal is 1 ;
  signal _zy_sva_key_type1_line9_8_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type1_line9_8_cpass: signal is 1 ;
  signal _zy_sva_b7 : std_logic ;
  attribute _2_state_ of _zy_sva_b7: signal is 1 ;
  signal _zy_sva_key_type1_line10_9_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type1_line10_9_ccheck: signal is 1 ;
  signal _zy_sva_key_type1_line10_9_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type1_line10_9_cpass: signal is 1 ;
  signal _zy_sva_b8 : std_logic ;
  attribute _2_state_ of _zy_sva_b8: signal is 1 ;
  signal _zy_sva_key_type1_line11a_10_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type1_line11a_10_ccheck: signal is 1 ;
  signal _zy_sva_key_type1_line11a_10_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type1_line11a_10_cpass: signal is 1 ;
  signal _zy_sva_b9 : std_logic ;
  attribute _2_state_ of _zy_sva_b9: signal is 1 ;
  signal _zy_sva_key_type1_line11b_11_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type1_line11b_11_ccheck: signal is 1 ;
  signal _zy_sva_key_type1_line11b_11_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type1_line11b_11_cpass: signal is 1 ;
  signal _zy_sva_b10 : std_logic ;
  attribute _2_state_ of _zy_sva_b10: signal is 1 ;
  signal _zy_sva_key_type1_line11c_12_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type1_line11c_12_ccheck: signal is 1 ;
  signal _zy_sva_key_type1_line11c_12_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type1_line11c_12_cpass: signal is 1 ;
  signal _zy_sva_b11 : std_logic ;
  attribute _2_state_ of _zy_sva_b11: signal is 1 ;
  signal _zy_sva_key_type1_line11d_13_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type1_line11d_13_ccheck: signal is 1 ;
  signal _zy_sva_key_type1_line11d_13_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type1_line11d_13_cpass: signal is 1 ;
  signal _zy_sva_b12 : std_logic ;
  attribute _2_state_ of _zy_sva_b12: signal is 1 ;
  signal _zy_sva_key_type1_line12a_14_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type1_line12a_14_ccheck: signal is 1 ;
  signal _zy_sva_key_type1_line12a_14_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type1_line12a_14_cpass: signal is 1 ;
  signal _zy_sva_b13 : std_logic ;
  attribute _2_state_ of _zy_sva_b13: signal is 1 ;
  signal _zy_sva_key_type1_line12b_15_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type1_line12b_15_ccheck: signal is 1 ;
  signal _zy_sva_key_type1_line12b_15_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type1_line12b_15_cpass: signal is 1 ;
  signal _zy_sva_b14 : std_logic ;
  attribute _2_state_ of _zy_sva_b14: signal is 1 ;
  signal _zy_sva_key_type9_line14_16_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type9_line14_16_ccheck: signal is 1 ;
  signal _zy_sva_key_type9_line14_16_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type9_line14_16_cpass: signal is 1 ;
  signal _zy_sva_b15 : std_logic ;
  attribute _2_state_ of _zy_sva_b15: signal is 1 ;
  signal _zy_sva_key_type9_line15_17_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type9_line15_17_ccheck: signal is 1 ;
  signal _zy_sva_key_type9_line15_17_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type9_line15_17_cpass: signal is 1 ;
  signal _zy_sva_b16 : std_logic ;
  attribute _2_state_ of _zy_sva_b16: signal is 1 ;
  signal _zy_sva_key_type9_line16a_18_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type9_line16a_18_ccheck: signal is 1 ;
  signal _zy_sva_key_type9_line16a_18_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type9_line16a_18_cpass: signal is 1 ;
  signal _zy_sva_b17 : std_logic ;
  attribute _2_state_ of _zy_sva_b17: signal is 1 ;
  signal _zy_sva_key_type9_line16b_19_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type9_line16b_19_ccheck: signal is 1 ;
  signal _zy_sva_key_type9_line16b_19_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type9_line16b_19_cpass: signal is 1 ;
  signal _zy_sva_b18 : std_logic ;
  attribute _2_state_ of _zy_sva_b18: signal is 1 ;
  signal _zy_sva_key_type9_line17a_20_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type9_line17a_20_ccheck: signal is 1 ;
  signal _zy_sva_key_type9_line17a_20_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type9_line17a_20_cpass: signal is 1 ;
  signal _zy_sva_b19 : std_logic ;
  attribute _2_state_ of _zy_sva_b19: signal is 1 ;
  signal _zy_sva_key_type9_line17b_21_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type9_line17b_21_ccheck: signal is 1 ;
  signal _zy_sva_key_type9_line17b_21_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type9_line17b_21_cpass: signal is 1 ;
  signal _zy_sva_b20 : std_logic ;
  attribute _2_state_ of _zy_sva_b20: signal is 1 ;
  signal _zy_sva_key_type9_line18a_22_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type9_line18a_22_ccheck: signal is 1 ;
  signal _zy_sva_key_type9_line18a_22_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type9_line18a_22_cpass: signal is 1 ;
  signal _zy_sva_b21 : std_logic ;
  attribute _2_state_ of _zy_sva_b21: signal is 1 ;
  signal _zy_sva_key_type9_line18b_23_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type9_line18b_23_ccheck: signal is 1 ;
  signal _zy_sva_key_type9_line18b_23_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type9_line18b_23_cpass: signal is 1 ;
  signal _zy_sva_b22 : std_logic ;
  attribute _2_state_ of _zy_sva_b22: signal is 1 ;
  signal _zy_sva_key_type9_line19a_24_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type9_line19a_24_ccheck: signal is 1 ;
  signal _zy_sva_key_type9_line19a_24_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type9_line19a_24_cpass: signal is 1 ;
  signal _zy_sva_b23 : std_logic ;
  attribute _2_state_ of _zy_sva_b23: signal is 1 ;
  signal _zy_sva_key_type9_line19b_25_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type9_line19b_25_ccheck: signal is 1 ;
  signal _zy_sva_key_type9_line19b_25_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type9_line19b_25_cpass: signal is 1 ;
  signal _zy_sva_b24 : std_logic ;
  attribute _2_state_ of _zy_sva_b24: signal is 1 ;
  signal _zy_sva_key_type9_line19c_26_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type9_line19c_26_ccheck: signal is 1 ;
  signal _zy_sva_key_type9_line19c_26_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type9_line19c_26_cpass: signal is 1 ;
  signal _zy_sva_b25 : std_logic ;
  attribute _2_state_ of _zy_sva_b25: signal is 1 ;
  signal _zy_sva_key_type9_line19d_27_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type9_line19d_27_ccheck: signal is 1 ;
  signal _zy_sva_key_type9_line19d_27_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_key_type9_line19d_27_cpass: signal is 1 ;
  signal _zy_sva_b26 : std_logic ;
  attribute _2_state_ of _zy_sva_b26: signal is 1 ;
  signal _zy_sva_guid_miss_aux_cmd_0_28_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_guid_miss_aux_cmd_0_28_ccheck: signal is 1 ;
  signal _zy_sva_guid_miss_aux_cmd_0_28_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_guid_miss_aux_cmd_0_28_cpass: signal is 1 ;
  signal _zy_sva_b27 : std_logic ;
  attribute _2_state_ of _zy_sva_b27: signal is 1 ;
  signal _zy_sva_guid_miss_aux_cmd_1_29_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_guid_miss_aux_cmd_1_29_ccheck: signal is 1 ;
  signal _zy_sva_guid_miss_aux_cmd_1_29_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_guid_miss_aux_cmd_1_29_cpass: signal is 1 ;
  signal _zy_sva_b28 : std_logic ;
  attribute _2_state_ of _zy_sva_b28: signal is 1 ;
  signal _zy_sva_guid_miss_aux_cmd_2_30_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_guid_miss_aux_cmd_2_30_ccheck: signal is 1 ;
  signal _zy_sva_guid_miss_aux_cmd_2_30_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_guid_miss_aux_cmd_2_30_cpass: signal is 1 ;
  signal _zy_sva_b29 : std_logic ;
  attribute _2_state_ of _zy_sva_b29: signal is 1 ;
  signal _zy_sva_guid_miss_aux_cmd_3_31_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_guid_miss_aux_cmd_3_31_ccheck: signal is 1 ;
  signal _zy_sva_guid_miss_aux_cmd_3_31_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_guid_miss_aux_cmd_3_31_cpass: signal is 1 ;
  signal _zy_sva_b30 : std_logic ;
  attribute _2_state_ of _zy_sva_b30: signal is 1 ;
  signal _zy_sva_guid_miss_aux_cmd_iv_0_32_ccheck : std_logic_vector(0 downto 0)
   := std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_guid_miss_aux_cmd_iv_0_32_ccheck: signal is 1 ;
  signal _zy_sva_guid_miss_aux_cmd_iv_0_32_cpass : std_logic_vector(0 downto 0)
   := std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_guid_miss_aux_cmd_iv_0_32_cpass: signal is 1 ;
  signal _zy_sva_b31 : std_logic ;
  attribute _2_state_ of _zy_sva_b31: signal is 1 ;
  signal _zy_sva_guid_miss_aux_cmd_iv_1_33_ccheck : std_logic_vector(0 downto 0)
   := std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_guid_miss_aux_cmd_iv_1_33_ccheck: signal is 1 ;
  signal _zy_sva_guid_miss_aux_cmd_iv_1_33_cpass : std_logic_vector(0 downto 0)
   := std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_guid_miss_aux_cmd_iv_1_33_cpass: signal is 1 ;
  signal _zy_sva_b32 : std_logic ;
  attribute _2_state_ of _zy_sva_b32: signal is 1 ;
  signal _zy_sva_guid_miss_aux_cmd_iv_2_34_ccheck : std_logic_vector(0 downto 0)
   := std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_guid_miss_aux_cmd_iv_2_34_ccheck: signal is 1 ;
  signal _zy_sva_guid_miss_aux_cmd_iv_2_34_cpass : std_logic_vector(0 downto 0)
   := std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_guid_miss_aux_cmd_iv_2_34_cpass: signal is 1 ;
  signal _zy_sva_b33 : std_logic ;
  attribute _2_state_ of _zy_sva_b33: signal is 1 ;
  signal _zy_sva_guid_miss_aux_cmd_iv_3_35_ccheck : std_logic_vector(0 downto 0)
   := std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_guid_miss_aux_cmd_iv_3_35_ccheck: signal is 1 ;
  signal _zy_sva_guid_miss_aux_cmd_iv_3_35_cpass : std_logic_vector(0 downto 0)
   := std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_guid_miss_aux_cmd_iv_3_35_cpass: signal is 1 ;
  signal _zy_sva_b34 : std_logic ;
  attribute _2_state_ of _zy_sva_b34: signal is 1 ;
  signal _zy_sva_iv_miss_aux_cmd_0_36_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_iv_miss_aux_cmd_0_36_ccheck: signal is 1 ;
  signal _zy_sva_iv_miss_aux_cmd_0_36_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_iv_miss_aux_cmd_0_36_cpass: signal is 1 ;
  signal _zy_sva_b35 : std_logic ;
  attribute _2_state_ of _zy_sva_b35: signal is 1 ;
  signal _zy_sva_iv_miss_aux_cmd_1_37_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_iv_miss_aux_cmd_1_37_ccheck: signal is 1 ;
  signal _zy_sva_iv_miss_aux_cmd_1_37_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_iv_miss_aux_cmd_1_37_cpass: signal is 1 ;
  signal _zy_sva_b36 : std_logic ;
  attribute _2_state_ of _zy_sva_b36: signal is 1 ;
  signal _zy_sva_iv_miss_aux_cmd_guid_38_ccheck : std_logic_vector(0 downto 0)
   := std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_iv_miss_aux_cmd_guid_38_ccheck: signal is 1 ;
  signal _zy_sva_iv_miss_aux_cmd_guid_38_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_iv_miss_aux_cmd_guid_38_cpass: signal is 1 ;
  signal _zy_sva_b37 : std_logic ;
  attribute _2_state_ of _zy_sva_b37: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_39_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_39_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_39_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_39_cpass: signal is 1 ;
  signal _zy_sva_b38 : std_logic ;
  attribute _2_state_ of _zy_sva_b38: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_iv_40_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_iv_40_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_iv_40_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_iv_40_cpass: signal is 1 ;
  signal _zy_sva_b39 : std_logic ;
  attribute _2_state_ of _zy_sva_b39: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_41_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_41_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_41_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_41_cpass: signal is 1 ;
  signal _zy_sva_b40 : std_logic ;
  attribute _2_state_ of _zy_sva_b40: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_42_ccheck : std_logic_vector(0 downto 0)
   := std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_iv_42_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_42_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_iv_42_cpass: signal is 1 ;
  signal _zy_sva_b41 : std_logic ;
  attribute _2_state_ of _zy_sva_b41: signal is 1 ;
  signal _zy_sva_brcm_key_type_43_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_key_type_43_ccheck: signal is 1 ;
  signal _zy_sva_brcm_key_type_43_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_key_type_43_cpass: signal is 1 ;
  signal _zy_sva_b42 : std_logic ;
  attribute _2_state_ of _zy_sva_b42: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_44_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_44_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_44_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_44_cpass: signal is 1 ;
  signal _zy_sva_b43 : std_logic ;
  attribute _2_state_ of _zy_sva_b43: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_iv_45_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_iv_45_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_iv_45_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_iv_45_cpass: signal is 1 ;
  signal _zy_sva_b44 : std_logic ;
  attribute _2_state_ of _zy_sva_b44: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_46_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_46_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_46_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_46_cpass: signal is 1 ;
  signal _zy_sva_b45 : std_logic ;
  attribute _2_state_ of _zy_sva_b45: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_47_ccheck : std_logic_vector(0 downto 0)
   := std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_iv_47_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_47_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_iv_47_cpass: signal is 1 ;
  signal _zy_sva_b46 : std_logic ;
  attribute _2_state_ of _zy_sva_b46: signal is 1 ;
  signal _zy_sva_brcm_key_type_48_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_key_type_48_ccheck: signal is 1 ;
  signal _zy_sva_brcm_key_type_48_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_key_type_48_cpass: signal is 1 ;
  signal _zy_sva_b47 : std_logic ;
  attribute _2_state_ of _zy_sva_b47: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_49_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_49_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_49_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_49_cpass: signal is 1 ;
  signal _zy_sva_b48 : std_logic ;
  attribute _2_state_ of _zy_sva_b48: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_iv_50_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_iv_50_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_iv_50_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_iv_50_cpass: signal is 1 ;
  signal _zy_sva_b49 : std_logic ;
  attribute _2_state_ of _zy_sva_b49: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_51_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_51_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_51_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_51_cpass: signal is 1 ;
  signal _zy_sva_b50 : std_logic ;
  attribute _2_state_ of _zy_sva_b50: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_52_ccheck : std_logic_vector(0 downto 0)
   := std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_iv_52_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_52_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_iv_52_cpass: signal is 1 ;
  signal _zy_sva_b51 : std_logic ;
  attribute _2_state_ of _zy_sva_b51: signal is 1 ;
  signal _zy_sva_brcm_key_type_53_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_key_type_53_ccheck: signal is 1 ;
  signal _zy_sva_brcm_key_type_53_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_key_type_53_cpass: signal is 1 ;
  signal _zy_sva_b52 : std_logic ;
  attribute _2_state_ of _zy_sva_b52: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_54_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_54_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_54_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_54_cpass: signal is 1 ;
  signal _zy_sva_b53 : std_logic ;
  attribute _2_state_ of _zy_sva_b53: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_iv_55_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_iv_55_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_iv_55_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_iv_55_cpass: signal is 1 ;
  signal _zy_sva_b54 : std_logic ;
  attribute _2_state_ of _zy_sva_b54: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_56_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_56_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_56_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_56_cpass: signal is 1 ;
  signal _zy_sva_b55 : std_logic ;
  attribute _2_state_ of _zy_sva_b55: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_57_ccheck : std_logic_vector(0 downto 0)
   := std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_iv_57_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_57_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_iv_57_cpass: signal is 1 ;
  signal _zy_sva_b56 : std_logic ;
  attribute _2_state_ of _zy_sva_b56: signal is 1 ;
  signal _zy_sva_brcm_key_type_58_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_key_type_58_ccheck: signal is 1 ;
  signal _zy_sva_brcm_key_type_58_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_key_type_58_cpass: signal is 1 ;
  signal _zy_sva_b57 : std_logic ;
  attribute _2_state_ of _zy_sva_b57: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_59_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_59_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_59_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_59_cpass: signal is 1 ;
  signal _zy_sva_b58 : std_logic ;
  attribute _2_state_ of _zy_sva_b58: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_iv_60_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_iv_60_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_iv_60_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_iv_60_cpass: signal is 1 ;
  signal _zy_sva_b59 : std_logic ;
  attribute _2_state_ of _zy_sva_b59: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_61_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_61_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_61_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_61_cpass: signal is 1 ;
  signal _zy_sva_b60 : std_logic ;
  attribute _2_state_ of _zy_sva_b60: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_62_ccheck : std_logic_vector(0 downto 0)
   := std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_iv_62_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_62_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_iv_62_cpass: signal is 1 ;
  signal _zy_sva_b61 : std_logic ;
  attribute _2_state_ of _zy_sva_b61: signal is 1 ;
  signal _zy_sva_brcm_key_type_63_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_key_type_63_ccheck: signal is 1 ;
  signal _zy_sva_brcm_key_type_63_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_key_type_63_cpass: signal is 1 ;
  signal _zy_sva_b62 : std_logic ;
  attribute _2_state_ of _zy_sva_b62: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_64_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_64_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_64_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_64_cpass: signal is 1 ;
  signal _zy_sva_b63 : std_logic ;
  attribute _2_state_ of _zy_sva_b63: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_iv_65_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_iv_65_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_iv_65_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_iv_65_cpass: signal is 1 ;
  signal _zy_sva_b64 : std_logic ;
  attribute _2_state_ of _zy_sva_b64: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_66_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_66_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_66_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_66_cpass: signal is 1 ;
  signal _zy_sva_b65 : std_logic ;
  attribute _2_state_ of _zy_sva_b65: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_67_ccheck : std_logic_vector(0 downto 0)
   := std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_iv_67_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_67_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_iv_67_cpass: signal is 1 ;
  signal _zy_sva_b66 : std_logic ;
  attribute _2_state_ of _zy_sva_b66: signal is 1 ;
  signal _zy_sva_brcm_key_type_68_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_key_type_68_ccheck: signal is 1 ;
  signal _zy_sva_brcm_key_type_68_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_key_type_68_cpass: signal is 1 ;
  signal _zy_sva_b67 : std_logic ;
  attribute _2_state_ of _zy_sva_b67: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_69_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_69_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_69_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_69_cpass: signal is 1 ;
  signal _zy_sva_b68 : std_logic ;
  attribute _2_state_ of _zy_sva_b68: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_iv_70_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_iv_70_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_iv_70_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_iv_70_cpass: signal is 1 ;
  signal _zy_sva_b69 : std_logic ;
  attribute _2_state_ of _zy_sva_b69: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_71_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_71_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_71_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_71_cpass: signal is 1 ;
  signal _zy_sva_b70 : std_logic ;
  attribute _2_state_ of _zy_sva_b70: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_72_ccheck : std_logic_vector(0 downto 0)
   := std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_iv_72_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_72_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_iv_72_cpass: signal is 1 ;
  signal _zy_sva_b71 : std_logic ;
  attribute _2_state_ of _zy_sva_b71: signal is 1 ;
  signal _zy_sva_brcm_key_type_73_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_key_type_73_ccheck: signal is 1 ;
  signal _zy_sva_brcm_key_type_73_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_key_type_73_cpass: signal is 1 ;
  signal _zy_sva_b72 : std_logic ;
  attribute _2_state_ of _zy_sva_b72: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_74_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_74_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_74_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_74_cpass: signal is 1 ;
  signal _zy_sva_b73 : std_logic ;
  attribute _2_state_ of _zy_sva_b73: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_iv_75_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_iv_75_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_iv_75_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_iv_75_cpass: signal is 1 ;
  signal _zy_sva_b74 : std_logic ;
  attribute _2_state_ of _zy_sva_b74: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_76_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_76_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_76_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_76_cpass: signal is 1 ;
  signal _zy_sva_b75 : std_logic ;
  attribute _2_state_ of _zy_sva_b75: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_77_ccheck : std_logic_vector(0 downto 0)
   := std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_iv_77_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_77_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_iv_77_cpass: signal is 1 ;
  signal _zy_sva_b76 : std_logic ;
  attribute _2_state_ of _zy_sva_b76: signal is 1 ;
  signal _zy_sva_brcm_key_type_78_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_key_type_78_ccheck: signal is 1 ;
  signal _zy_sva_brcm_key_type_78_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_key_type_78_cpass: signal is 1 ;
  signal _zy_sva_b77 : std_logic ;
  attribute _2_state_ of _zy_sva_b77: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_79_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_79_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_79_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_79_cpass: signal is 1 ;
  signal _zy_sva_b78 : std_logic ;
  attribute _2_state_ of _zy_sva_b78: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_iv_80_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_iv_80_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_iv_80_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_iv_80_cpass: signal is 1 ;
  signal _zy_sva_b79 : std_logic ;
  attribute _2_state_ of _zy_sva_b79: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_81_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_81_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_81_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_81_cpass: signal is 1 ;
  signal _zy_sva_b80 : std_logic ;
  attribute _2_state_ of _zy_sva_b80: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_82_ccheck : std_logic_vector(0 downto 0)
   := std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_iv_82_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_82_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_iv_82_cpass: signal is 1 ;
  signal _zy_sva_b81 : std_logic ;
  attribute _2_state_ of _zy_sva_b81: signal is 1 ;
  signal _zy_sva_brcm_key_type_83_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_key_type_83_ccheck: signal is 1 ;
  signal _zy_sva_brcm_key_type_83_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_key_type_83_cpass: signal is 1 ;
  signal _zy_sva_b82 : std_logic ;
  attribute _2_state_ of _zy_sva_b82: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_84_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_84_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_84_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_84_cpass: signal is 1 ;
  signal _zy_sva_b83 : std_logic ;
  attribute _2_state_ of _zy_sva_b83: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_iv_85_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_iv_85_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_iv_85_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_iv_85_cpass: signal is 1 ;
  signal _zy_sva_b84 : std_logic ;
  attribute _2_state_ of _zy_sva_b84: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_86_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_86_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_86_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_86_cpass: signal is 1 ;
  signal _zy_sva_b85 : std_logic ;
  attribute _2_state_ of _zy_sva_b85: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_87_ccheck : std_logic_vector(0 downto 0)
   := std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_iv_87_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_87_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_iv_87_cpass: signal is 1 ;
  signal _zy_sva_b86 : std_logic ;
  attribute _2_state_ of _zy_sva_b86: signal is 1 ;
  signal _zy_sva_brcm_key_type_88_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_key_type_88_ccheck: signal is 1 ;
  signal _zy_sva_brcm_key_type_88_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_key_type_88_cpass: signal is 1 ;
  signal _zy_sva_b87 : std_logic ;
  attribute _2_state_ of _zy_sva_b87: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_89_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_89_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_89_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_89_cpass: signal is 1 ;
  signal _zy_sva_b88 : std_logic ;
  attribute _2_state_ of _zy_sva_b88: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_iv_90_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_iv_90_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_iv_90_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_iv_90_cpass: signal is 1 ;
  signal _zy_sva_b89 : std_logic ;
  attribute _2_state_ of _zy_sva_b89: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_91_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_91_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_91_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_91_cpass: signal is 1 ;
  signal _zy_sva_b90 : std_logic ;
  attribute _2_state_ of _zy_sva_b90: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_92_ccheck : std_logic_vector(0 downto 0)
   := std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_iv_92_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_92_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_iv_92_cpass: signal is 1 ;
  signal _zy_sva_b91 : std_logic ;
  attribute _2_state_ of _zy_sva_b91: signal is 1 ;
  signal _zy_sva_brcm_key_type_93_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_key_type_93_ccheck: signal is 1 ;
  signal _zy_sva_brcm_key_type_93_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_key_type_93_cpass: signal is 1 ;
  signal _zy_sva_b92 : std_logic ;
  attribute _2_state_ of _zy_sva_b92: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_94_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_94_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_94_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_94_cpass: signal is 1 ;
  signal _zy_sva_b93 : std_logic ;
  attribute _2_state_ of _zy_sva_b93: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_iv_95_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_iv_95_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_iv_95_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_iv_95_cpass: signal is 1 ;
  signal _zy_sva_b94 : std_logic ;
  attribute _2_state_ of _zy_sva_b94: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_96_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_96_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_96_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_96_cpass: signal is 1 ;
  signal _zy_sva_b95 : std_logic ;
  attribute _2_state_ of _zy_sva_b95: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_97_ccheck : std_logic_vector(0 downto 0)
   := std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_iv_97_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_97_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_iv_97_cpass: signal is 1 ;
  signal _zy_sva_b96 : std_logic ;
  attribute _2_state_ of _zy_sva_b96: signal is 1 ;
  signal _zy_sva_brcm_key_type_98_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_key_type_98_ccheck: signal is 1 ;
  signal _zy_sva_brcm_key_type_98_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_key_type_98_cpass: signal is 1 ;
  signal _zy_sva_b97 : std_logic ;
  attribute _2_state_ of _zy_sva_b97: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_99_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_99_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_99_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_99_cpass: signal is 1 ;
  signal _zy_sva_b98 : std_logic ;
  attribute _2_state_ of _zy_sva_b98: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_iv_100_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_iv_100_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_iv_100_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_iv_100_cpass: signal is 1 ;
  signal _zy_sva_b99 : std_logic ;
  attribute _2_state_ of _zy_sva_b99: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_101_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_101_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_101_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_101_cpass: signal is 1 ;
  signal _zy_sva_b100 : std_logic ;
  attribute _2_state_ of _zy_sva_b100: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_102_ccheck : std_logic_vector(0 downto 0)
   := std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_iv_102_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_102_cpass : std_logic_vector(0 downto 0)
   := std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_iv_102_cpass: signal is 1 ;
  signal _zy_sva_b101 : std_logic ;
  attribute _2_state_ of _zy_sva_b101: signal is 1 ;
  signal _zy_sva_brcm_key_type_103_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_key_type_103_ccheck: signal is 1 ;
  signal _zy_sva_brcm_key_type_103_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_key_type_103_cpass: signal is 1 ;
  signal _zy_sva_b102 : std_logic ;
  attribute _2_state_ of _zy_sva_b102: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_104_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_104_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_104_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_104_cpass: signal is 1 ;
  signal _zy_sva_b103 : std_logic ;
  attribute _2_state_ of _zy_sva_b103: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_iv_105_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_iv_105_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_iv_105_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_iv_105_cpass: signal is 1 ;
  signal _zy_sva_b104 : std_logic ;
  attribute _2_state_ of _zy_sva_b104: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_106_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_106_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_106_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_106_cpass: signal is 1 ;
  signal _zy_sva_b105 : std_logic ;
  attribute _2_state_ of _zy_sva_b105: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_107_ccheck : std_logic_vector(0 downto 0)
   := std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_iv_107_ccheck: signal is 1 ;
  signal _zy_sva_brcm_aux_cmd_guid_iv_107_cpass : std_logic_vector(0 downto 0)
   := std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_aux_cmd_guid_iv_107_cpass: signal is 1 ;
  signal _zy_sva_b106 : std_logic ;
  attribute _2_state_ of _zy_sva_b106: signal is 1 ;
  signal _zy_sva_brcm_key_type_108_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_key_type_108_ccheck: signal is 1 ;
  signal _zy_sva_brcm_key_type_108_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_key_type_108_cpass: signal is 1 ;
  signal _zy_sva_b107 : std_logic ;
  attribute _2_state_ of _zy_sva_b107: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_109_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_109_ccheck: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_109_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_109_cpass: signal is 1 ;
  signal _zy_sva_b108 : std_logic ;
  attribute _2_state_ of _zy_sva_b108: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_110_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_110_ccheck: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_110_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_110_cpass: signal is 1 ;
  signal _zy_sva_b109 : std_logic ;
  attribute _2_state_ of _zy_sva_b109: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_111_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_111_ccheck: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_111_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_111_cpass: signal is 1 ;
  signal _zy_sva_b110 : std_logic ;
  attribute _2_state_ of _zy_sva_b110: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_112_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_112_ccheck: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_112_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_112_cpass: signal is 1 ;
  signal _zy_sva_b111 : std_logic ;
  attribute _2_state_ of _zy_sva_b111: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_113_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_113_ccheck: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_113_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_113_cpass: signal is 1 ;
  signal _zy_sva_b112 : std_logic ;
  attribute _2_state_ of _zy_sva_b112: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_114_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_114_ccheck: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_114_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_114_cpass: signal is 1 ;
  signal _zy_sva_b113 : std_logic ;
  attribute _2_state_ of _zy_sva_b113: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_115_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_115_ccheck: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_115_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_115_cpass: signal is 1 ;
  signal _zy_sva_b114 : std_logic ;
  attribute _2_state_ of _zy_sva_b114: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_116_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_116_ccheck: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_116_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_116_cpass: signal is 1 ;
  signal _zy_sva_b115 : std_logic ;
  attribute _2_state_ of _zy_sva_b115: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_117_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_117_ccheck: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_117_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_117_cpass: signal is 1 ;
  signal _zy_sva_b116 : std_logic ;
  attribute _2_state_ of _zy_sva_b116: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_118_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_118_ccheck: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_118_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_118_cpass: signal is 1 ;
  signal _zy_sva_b117 : std_logic ;
  attribute _2_state_ of _zy_sva_b117: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_119_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_119_ccheck: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_119_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_119_cpass: signal is 1 ;
  signal _zy_sva_b118 : std_logic ;
  attribute _2_state_ of _zy_sva_b118: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_120_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_120_ccheck: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_120_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_120_cpass: signal is 1 ;
  signal _zy_sva_b119 : std_logic ;
  attribute _2_state_ of _zy_sva_b119: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_121_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_121_ccheck: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_121_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_121_cpass: signal is 1 ;
  signal _zy_sva_b120 : std_logic ;
  attribute _2_state_ of _zy_sva_b120: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_122_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_122_ccheck: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_122_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_122_cpass: signal is 1 ;
  signal _zy_sva_b121 : std_logic ;
  attribute _2_state_ of _zy_sva_b121: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_123_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_123_ccheck: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_123_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_123_cpass: signal is 1 ;
  signal _zy_sva_b122 : std_logic ;
  attribute _2_state_ of _zy_sva_b122: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_124_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_124_ccheck: signal is 1 ;
  signal _zy_sva_brcm_kdf_ops_124_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_brcm_kdf_ops_124_cpass: signal is 1 ;
  signal _zy_sva_b123 : std_logic ;
  attribute _2_state_ of _zy_sva_b123: signal is 1 ;
  signal _zy_sva_null_gcm_125_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_gcm_125_ccheck: signal is 1 ;
  signal _zy_sva_null_gcm_125_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_gcm_125_cpass: signal is 1 ;
  signal _zy_sva_b124 : std_logic ;
  attribute _2_state_ of _zy_sva_b124: signal is 1 ;
  signal _zy_sva_sha_gcm_126_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_gcm_126_ccheck: signal is 1 ;
  signal _zy_sva_sha_gcm_126_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_gcm_126_cpass: signal is 1 ;
  signal _zy_sva_b125 : std_logic ;
  attribute _2_state_ of _zy_sva_b125: signal is 1 ;
  signal _zy_sva_null_xts_127_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_xts_127_ccheck: signal is 1 ;
  signal _zy_sva_null_xts_127_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_xts_127_cpass: signal is 1 ;
  signal _zy_sva_b126 : std_logic ;
  attribute _2_state_ of _zy_sva_b126: signal is 1 ;
  signal _zy_sva_sha_xts_128_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_xts_128_ccheck: signal is 1 ;
  signal _zy_sva_sha_xts_128_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_xts_128_cpass: signal is 1 ;
  signal _zy_sva_b127 : std_logic ;
  attribute _2_state_ of _zy_sva_b127: signal is 1 ;
  signal _zy_sva_null_null_129_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_null_129_ccheck: signal is 1 ;
  signal _zy_sva_null_null_129_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_null_129_cpass: signal is 1 ;
  signal _zy_sva_b128 : std_logic ;
  attribute _2_state_ of _zy_sva_b128: signal is 1 ;
  signal _zy_sva_sha_null_130_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_null_130_ccheck: signal is 1 ;
  signal _zy_sva_sha_null_130_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_null_130_cpass: signal is 1 ;
  signal _zy_sva_b129 : std_logic ;
  attribute _2_state_ of _zy_sva_b129: signal is 1 ;
  signal _zy_sva_hmac_gcm_131_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_gcm_131_ccheck: signal is 1 ;
  signal _zy_sva_hmac_gcm_131_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_gcm_131_cpass: signal is 1 ;
  signal _zy_sva_b130 : std_logic ;
  attribute _2_state_ of _zy_sva_b130: signal is 1 ;
  signal _zy_sva_hmac_xts_132_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_xts_132_ccheck: signal is 1 ;
  signal _zy_sva_hmac_xts_132_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_xts_132_cpass: signal is 1 ;
  signal _zy_sva_b131 : std_logic ;
  attribute _2_state_ of _zy_sva_b131: signal is 1 ;
  signal _zy_sva_hmac_null_133_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_null_133_ccheck: signal is 1 ;
  signal _zy_sva_hmac_null_133_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_null_133_cpass: signal is 1 ;
  signal _zy_sva_b132 : std_logic ;
  attribute _2_state_ of _zy_sva_b132: signal is 1 ;
  signal _zy_sva_null_gcm_134_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_gcm_134_ccheck: signal is 1 ;
  signal _zy_sva_null_gcm_134_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_gcm_134_cpass: signal is 1 ;
  signal _zy_sva_b133 : std_logic ;
  attribute _2_state_ of _zy_sva_b133: signal is 1 ;
  signal _zy_sva_sha_gcm_135_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_gcm_135_ccheck: signal is 1 ;
  signal _zy_sva_sha_gcm_135_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_gcm_135_cpass: signal is 1 ;
  signal _zy_sva_b134 : std_logic ;
  attribute _2_state_ of _zy_sva_b134: signal is 1 ;
  signal _zy_sva_null_xts_136_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_xts_136_ccheck: signal is 1 ;
  signal _zy_sva_null_xts_136_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_xts_136_cpass: signal is 1 ;
  signal _zy_sva_b135 : std_logic ;
  attribute _2_state_ of _zy_sva_b135: signal is 1 ;
  signal _zy_sva_sha_xts_137_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_xts_137_ccheck: signal is 1 ;
  signal _zy_sva_sha_xts_137_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_xts_137_cpass: signal is 1 ;
  signal _zy_sva_b136 : std_logic ;
  attribute _2_state_ of _zy_sva_b136: signal is 1 ;
  signal _zy_sva_null_null_138_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_null_138_ccheck: signal is 1 ;
  signal _zy_sva_null_null_138_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_null_138_cpass: signal is 1 ;
  signal _zy_sva_b137 : std_logic ;
  attribute _2_state_ of _zy_sva_b137: signal is 1 ;
  signal _zy_sva_sha_null_139_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_null_139_ccheck: signal is 1 ;
  signal _zy_sva_sha_null_139_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_null_139_cpass: signal is 1 ;
  signal _zy_sva_b138 : std_logic ;
  attribute _2_state_ of _zy_sva_b138: signal is 1 ;
  signal _zy_sva_hmac_gcm_140_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_gcm_140_ccheck: signal is 1 ;
  signal _zy_sva_hmac_gcm_140_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_gcm_140_cpass: signal is 1 ;
  signal _zy_sva_b139 : std_logic ;
  attribute _2_state_ of _zy_sva_b139: signal is 1 ;
  signal _zy_sva_hmac_xts_141_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_xts_141_ccheck: signal is 1 ;
  signal _zy_sva_hmac_xts_141_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_xts_141_cpass: signal is 1 ;
  signal _zy_sva_b140 : std_logic ;
  attribute _2_state_ of _zy_sva_b140: signal is 1 ;
  signal _zy_sva_hmac_null_142_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_null_142_ccheck: signal is 1 ;
  signal _zy_sva_hmac_null_142_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_null_142_cpass: signal is 1 ;
  signal _zy_sva_b141 : std_logic ;
  attribute _2_state_ of _zy_sva_b141: signal is 1 ;
  signal _zy_sva_null_gcm_143_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_gcm_143_ccheck: signal is 1 ;
  signal _zy_sva_null_gcm_143_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_gcm_143_cpass: signal is 1 ;
  signal _zy_sva_b142 : std_logic ;
  attribute _2_state_ of _zy_sva_b142: signal is 1 ;
  signal _zy_sva_sha_gcm_144_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_gcm_144_ccheck: signal is 1 ;
  signal _zy_sva_sha_gcm_144_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_gcm_144_cpass: signal is 1 ;
  signal _zy_sva_b143 : std_logic ;
  attribute _2_state_ of _zy_sva_b143: signal is 1 ;
  signal _zy_sva_null_xts_145_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_xts_145_ccheck: signal is 1 ;
  signal _zy_sva_null_xts_145_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_xts_145_cpass: signal is 1 ;
  signal _zy_sva_b144 : std_logic ;
  attribute _2_state_ of _zy_sva_b144: signal is 1 ;
  signal _zy_sva_sha_xts_146_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_xts_146_ccheck: signal is 1 ;
  signal _zy_sva_sha_xts_146_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_xts_146_cpass: signal is 1 ;
  signal _zy_sva_b145 : std_logic ;
  attribute _2_state_ of _zy_sva_b145: signal is 1 ;
  signal _zy_sva_null_null_147_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_null_147_ccheck: signal is 1 ;
  signal _zy_sva_null_null_147_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_null_147_cpass: signal is 1 ;
  signal _zy_sva_b146 : std_logic ;
  attribute _2_state_ of _zy_sva_b146: signal is 1 ;
  signal _zy_sva_sha_null_148_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_null_148_ccheck: signal is 1 ;
  signal _zy_sva_sha_null_148_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_null_148_cpass: signal is 1 ;
  signal _zy_sva_b147 : std_logic ;
  attribute _2_state_ of _zy_sva_b147: signal is 1 ;
  signal _zy_sva_hmac_gcm_149_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_gcm_149_ccheck: signal is 1 ;
  signal _zy_sva_hmac_gcm_149_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_gcm_149_cpass: signal is 1 ;
  signal _zy_sva_b148 : std_logic ;
  attribute _2_state_ of _zy_sva_b148: signal is 1 ;
  signal _zy_sva_hmac_xts_150_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_xts_150_ccheck: signal is 1 ;
  signal _zy_sva_hmac_xts_150_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_xts_150_cpass: signal is 1 ;
  signal _zy_sva_b149 : std_logic ;
  attribute _2_state_ of _zy_sva_b149: signal is 1 ;
  signal _zy_sva_hmac_null_151_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_null_151_ccheck: signal is 1 ;
  signal _zy_sva_hmac_null_151_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_null_151_cpass: signal is 1 ;
  signal _zy_sva_b150 : std_logic ;
  attribute _2_state_ of _zy_sva_b150: signal is 1 ;
  signal _zy_sva_null_gcm_152_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_gcm_152_ccheck: signal is 1 ;
  signal _zy_sva_null_gcm_152_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_gcm_152_cpass: signal is 1 ;
  signal _zy_sva_b151 : std_logic ;
  attribute _2_state_ of _zy_sva_b151: signal is 1 ;
  signal _zy_sva_sha_gcm_153_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_gcm_153_ccheck: signal is 1 ;
  signal _zy_sva_sha_gcm_153_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_gcm_153_cpass: signal is 1 ;
  signal _zy_sva_b152 : std_logic ;
  attribute _2_state_ of _zy_sva_b152: signal is 1 ;
  signal _zy_sva_null_xts_154_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_xts_154_ccheck: signal is 1 ;
  signal _zy_sva_null_xts_154_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_xts_154_cpass: signal is 1 ;
  signal _zy_sva_b153 : std_logic ;
  attribute _2_state_ of _zy_sva_b153: signal is 1 ;
  signal _zy_sva_sha_xts_155_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_xts_155_ccheck: signal is 1 ;
  signal _zy_sva_sha_xts_155_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_xts_155_cpass: signal is 1 ;
  signal _zy_sva_b154 : std_logic ;
  attribute _2_state_ of _zy_sva_b154: signal is 1 ;
  signal _zy_sva_null_null_156_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_null_156_ccheck: signal is 1 ;
  signal _zy_sva_null_null_156_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_null_156_cpass: signal is 1 ;
  signal _zy_sva_b155 : std_logic ;
  attribute _2_state_ of _zy_sva_b155: signal is 1 ;
  signal _zy_sva_sha_null_157_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_null_157_ccheck: signal is 1 ;
  signal _zy_sva_sha_null_157_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_null_157_cpass: signal is 1 ;
  signal _zy_sva_b156 : std_logic ;
  attribute _2_state_ of _zy_sva_b156: signal is 1 ;
  signal _zy_sva_hmac_gcm_158_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_gcm_158_ccheck: signal is 1 ;
  signal _zy_sva_hmac_gcm_158_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_gcm_158_cpass: signal is 1 ;
  signal _zy_sva_b157 : std_logic ;
  attribute _2_state_ of _zy_sva_b157: signal is 1 ;
  signal _zy_sva_hmac_xts_159_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_xts_159_ccheck: signal is 1 ;
  signal _zy_sva_hmac_xts_159_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_xts_159_cpass: signal is 1 ;
  signal _zy_sva_b158 : std_logic ;
  attribute _2_state_ of _zy_sva_b158: signal is 1 ;
  signal _zy_sva_hmac_null_160_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_null_160_ccheck: signal is 1 ;
  signal _zy_sva_hmac_null_160_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_null_160_cpass: signal is 1 ;
  signal _zy_sva_b159 : std_logic ;
  attribute _2_state_ of _zy_sva_b159: signal is 1 ;
  signal _zy_sva_null_gcm_161_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_gcm_161_ccheck: signal is 1 ;
  signal _zy_sva_null_gcm_161_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_gcm_161_cpass: signal is 1 ;
  signal _zy_sva_b160 : std_logic ;
  attribute _2_state_ of _zy_sva_b160: signal is 1 ;
  signal _zy_sva_sha_gcm_162_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_gcm_162_ccheck: signal is 1 ;
  signal _zy_sva_sha_gcm_162_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_gcm_162_cpass: signal is 1 ;
  signal _zy_sva_b161 : std_logic ;
  attribute _2_state_ of _zy_sva_b161: signal is 1 ;
  signal _zy_sva_null_xts_163_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_xts_163_ccheck: signal is 1 ;
  signal _zy_sva_null_xts_163_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_xts_163_cpass: signal is 1 ;
  signal _zy_sva_b162 : std_logic ;
  attribute _2_state_ of _zy_sva_b162: signal is 1 ;
  signal _zy_sva_sha_xts_164_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_xts_164_ccheck: signal is 1 ;
  signal _zy_sva_sha_xts_164_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_xts_164_cpass: signal is 1 ;
  signal _zy_sva_b163 : std_logic ;
  attribute _2_state_ of _zy_sva_b163: signal is 1 ;
  signal _zy_sva_null_null_165_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_null_165_ccheck: signal is 1 ;
  signal _zy_sva_null_null_165_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_null_165_cpass: signal is 1 ;
  signal _zy_sva_b164 : std_logic ;
  attribute _2_state_ of _zy_sva_b164: signal is 1 ;
  signal _zy_sva_sha_null_166_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_null_166_ccheck: signal is 1 ;
  signal _zy_sva_sha_null_166_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_null_166_cpass: signal is 1 ;
  signal _zy_sva_b165 : std_logic ;
  attribute _2_state_ of _zy_sva_b165: signal is 1 ;
  signal _zy_sva_hmac_gcm_167_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_gcm_167_ccheck: signal is 1 ;
  signal _zy_sva_hmac_gcm_167_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_gcm_167_cpass: signal is 1 ;
  signal _zy_sva_b166 : std_logic ;
  attribute _2_state_ of _zy_sva_b166: signal is 1 ;
  signal _zy_sva_hmac_xts_168_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_xts_168_ccheck: signal is 1 ;
  signal _zy_sva_hmac_xts_168_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_xts_168_cpass: signal is 1 ;
  signal _zy_sva_b167 : std_logic ;
  attribute _2_state_ of _zy_sva_b167: signal is 1 ;
  signal _zy_sva_hmac_null_169_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_null_169_ccheck: signal is 1 ;
  signal _zy_sva_hmac_null_169_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_null_169_cpass: signal is 1 ;
  signal _zy_sva_b168 : std_logic ;
  attribute _2_state_ of _zy_sva_b168: signal is 1 ;
  signal _zy_sva_null_gcm_170_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_gcm_170_ccheck: signal is 1 ;
  signal _zy_sva_null_gcm_170_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_gcm_170_cpass: signal is 1 ;
  signal _zy_sva_b169 : std_logic ;
  attribute _2_state_ of _zy_sva_b169: signal is 1 ;
  signal _zy_sva_sha_gcm_171_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_gcm_171_ccheck: signal is 1 ;
  signal _zy_sva_sha_gcm_171_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_gcm_171_cpass: signal is 1 ;
  signal _zy_sva_b170 : std_logic ;
  attribute _2_state_ of _zy_sva_b170: signal is 1 ;
  signal _zy_sva_null_xts_172_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_xts_172_ccheck: signal is 1 ;
  signal _zy_sva_null_xts_172_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_xts_172_cpass: signal is 1 ;
  signal _zy_sva_b171 : std_logic ;
  attribute _2_state_ of _zy_sva_b171: signal is 1 ;
  signal _zy_sva_sha_xts_173_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_xts_173_ccheck: signal is 1 ;
  signal _zy_sva_sha_xts_173_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_xts_173_cpass: signal is 1 ;
  signal _zy_sva_b172 : std_logic ;
  attribute _2_state_ of _zy_sva_b172: signal is 1 ;
  signal _zy_sva_null_null_174_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_null_174_ccheck: signal is 1 ;
  signal _zy_sva_null_null_174_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_null_null_174_cpass: signal is 1 ;
  signal _zy_sva_b173 : std_logic ;
  attribute _2_state_ of _zy_sva_b173: signal is 1 ;
  signal _zy_sva_sha_null_175_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_null_175_ccheck: signal is 1 ;
  signal _zy_sva_sha_null_175_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_sha_null_175_cpass: signal is 1 ;
  signal _zy_sva_b174 : std_logic ;
  attribute _2_state_ of _zy_sva_b174: signal is 1 ;
  signal _zy_sva_hmac_gcm_176_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_gcm_176_ccheck: signal is 1 ;
  signal _zy_sva_hmac_gcm_176_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_gcm_176_cpass: signal is 1 ;
  signal _zy_sva_b175 : std_logic ;
  attribute _2_state_ of _zy_sva_b175: signal is 1 ;
  signal _zy_sva_hmac_xts_177_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_xts_177_ccheck: signal is 1 ;
  signal _zy_sva_hmac_xts_177_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_xts_177_cpass: signal is 1 ;
  signal _zy_sva_b176 : std_logic ;
  attribute _2_state_ of _zy_sva_b176: signal is 1 ;
  signal _zy_sva_hmac_null_178_ccheck : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_null_178_ccheck: signal is 1 ;
  signal _zy_sva_hmac_null_178_cpass : std_logic_vector(0 downto 0) :=
   std_logic_vector'("0") ;
  attribute _2_state_ of _zy_sva_hmac_null_178_cpass: signal is 1 ;
  signal _zy_sva_b177 : std_logic ;
  attribute _2_state_ of _zy_sva_b177: signal is 1 ;
  signal _zyL234_tfiRv52 : std_logic_vector(63 downto 0) ;
  signal _zyL252_tfiRv53 : std_logic ;
  signal _zyL253_tfiRv54 : std_logic ;
  signal _zyL254_tfiRv55 : std_logic ;
  signal _zyL255_tfiRv56 : std_logic ;
  signal _zyL288_tfiRv57 : std_logic_vector(63 downto 0) ;
  signal _zyL293_tfiRv58 : std_logic_vector(63 downto 0) ;
  signal _zyL301_tfiRv59 : std_logic_vector(63 downto 0) ;
  signal _zyL306_tfiRv60 : std_logic_vector(63 downto 0) ;
  signal _zyL313_tfiRv61 : std_logic_vector(63 downto 0) ;
  signal _zyL321_tfiRv62 : std_logic_vector(63 downto 0) ;
  signal _zyL327_tfiRv63 : std_logic_vector(63 downto 0) ;
  signal _zyL337_tfiRv64 : std_logic_vector(63 downto 0) ;
  signal _zyL346_tfiRv65 : std_logic_vector(63 downto 0) ;
  signal _zyL354_tfiRv66 : std_logic_vector(63 downto 0) ;
  signal _zyL359_tfiRv67 : std_logic_vector(63 downto 0) ;
  signal _zyL368_tfiRv68 : std_logic_vector(63 downto 0) ;
  signal _zyL373_tfiRv69 : std_logic_vector(63 downto 0) ;
  signal _zyL382_tfiRv70 : std_logic_vector(63 downto 0) ;
  signal _zyL390_tfiRv71 : std_logic_vector(63 downto 0) ;
  signal _zyL395_tfiRv72 : std_logic_vector(63 downto 0) ;
  signal _zyL410_tfiRv73 : std_logic_vector(63 downto 0) ;
  signal _zyL485_tfiRv74 : std_logic ;
  signal _zyL486_tfiRv75 : std_logic ;
  signal _zyL489_tfiRv76 : std_logic ;
  signal _zyL489_tfiRv77 : std_logic ;
  signal _zyL492_tfiRv78 : std_logic ;
  signal _zyL526_tfiRv79 : std_logic_vector(63 downto 0) ;
  signal _zyL527_tfiRv80 : std_logic_vector(63 downto 0) ;
  signal _zyL541_tfiRv81 : std_logic_vector(63 downto 0) ;
  signal _zyL542_tfiRv82 : std_logic_vector(63 downto 0) ;
  signal _zyL555_tfiRv83 : std_logic_vector(63 downto 0) ;
  signal _zyL556_tfiRv84 : std_logic_vector(63 downto 0) ;
  signal _zyL569_tfiRv85 : std_logic_vector(63 downto 0) ;
  signal _zyL570_tfiRv86 : std_logic_vector(63 downto 0) ;
  -- quickturn keep_net _zy_sva_key_type0_line4_1_ccheck
  -- quickturn keep_net _zy_sva_key_type0_line4_1_cpass
  -- quickturn keep_net _zy_sva_key_type0_line5a_2_ccheck
  -- quickturn keep_net _zy_sva_key_type0_line5a_2_cpass
  -- quickturn keep_net _zy_sva_key_type0_line5b_3_ccheck
  -- quickturn keep_net _zy_sva_key_type0_line5b_3_cpass
  -- quickturn keep_net _zy_sva_key_type1_line7a_4_ccheck
  -- quickturn keep_net _zy_sva_key_type1_line7a_4_cpass
  -- quickturn keep_net _zy_sva_key_type1_line7b_5_ccheck
  -- quickturn keep_net _zy_sva_key_type1_line7b_5_cpass
  -- quickturn keep_net _zy_sva_key_type1_line8a_6_ccheck
  -- quickturn keep_net _zy_sva_key_type1_line8a_6_cpass
  -- quickturn keep_net _zy_sva_key_type1_line8b_7_ccheck
  -- quickturn keep_net _zy_sva_key_type1_line8b_7_cpass
  -- quickturn keep_net _zy_sva_key_type1_line9_8_ccheck
  -- quickturn keep_net _zy_sva_key_type1_line9_8_cpass
  -- quickturn keep_net _zy_sva_key_type1_line10_9_ccheck
  -- quickturn keep_net _zy_sva_key_type1_line10_9_cpass
  -- quickturn keep_net _zy_sva_key_type1_line11a_10_ccheck
  -- quickturn keep_net _zy_sva_key_type1_line11a_10_cpass
  -- quickturn keep_net _zy_sva_key_type1_line11b_11_ccheck
  -- quickturn keep_net _zy_sva_key_type1_line11b_11_cpass
  -- quickturn keep_net _zy_sva_key_type1_line11c_12_ccheck
  -- quickturn keep_net _zy_sva_key_type1_line11c_12_cpass
  -- quickturn keep_net _zy_sva_key_type1_line11d_13_ccheck
  -- quickturn keep_net _zy_sva_key_type1_line11d_13_cpass
  -- quickturn keep_net _zy_sva_key_type1_line12a_14_ccheck
  -- quickturn keep_net _zy_sva_key_type1_line12a_14_cpass
  -- quickturn keep_net _zy_sva_key_type1_line12b_15_ccheck
  -- quickturn keep_net _zy_sva_key_type1_line12b_15_cpass
  -- quickturn keep_net _zy_sva_key_type9_line14_16_ccheck
  -- quickturn keep_net _zy_sva_key_type9_line14_16_cpass
  -- quickturn keep_net _zy_sva_key_type9_line15_17_ccheck
  -- quickturn keep_net _zy_sva_key_type9_line15_17_cpass
  -- quickturn keep_net _zy_sva_key_type9_line16a_18_ccheck
  -- quickturn keep_net _zy_sva_key_type9_line16a_18_cpass
  -- quickturn keep_net _zy_sva_key_type9_line16b_19_ccheck
  -- quickturn keep_net _zy_sva_key_type9_line16b_19_cpass
  -- quickturn keep_net _zy_sva_key_type9_line17a_20_ccheck
  -- quickturn keep_net _zy_sva_key_type9_line17a_20_cpass
  -- quickturn keep_net _zy_sva_key_type9_line17b_21_ccheck
  -- quickturn keep_net _zy_sva_key_type9_line17b_21_cpass
  -- quickturn keep_net _zy_sva_key_type9_line18a_22_ccheck
  -- quickturn keep_net _zy_sva_key_type9_line18a_22_cpass
  -- quickturn keep_net _zy_sva_key_type9_line18b_23_ccheck
  -- quickturn keep_net _zy_sva_key_type9_line18b_23_cpass
  -- quickturn keep_net _zy_sva_key_type9_line19a_24_ccheck
  -- quickturn keep_net _zy_sva_key_type9_line19a_24_cpass
  -- quickturn keep_net _zy_sva_key_type9_line19b_25_ccheck
  -- quickturn keep_net _zy_sva_key_type9_line19b_25_cpass
  -- quickturn keep_net _zy_sva_key_type9_line19c_26_ccheck
  -- quickturn keep_net _zy_sva_key_type9_line19c_26_cpass
  -- quickturn keep_net _zy_sva_key_type9_line19d_27_ccheck
  -- quickturn keep_net _zy_sva_key_type9_line19d_27_cpass
  -- quickturn keep_net _zy_sva_guid_miss_aux_cmd_0_28_ccheck
  -- quickturn keep_net _zy_sva_guid_miss_aux_cmd_0_28_cpass
  -- quickturn keep_net _zy_sva_guid_miss_aux_cmd_1_29_ccheck
  -- quickturn keep_net _zy_sva_guid_miss_aux_cmd_1_29_cpass
  -- quickturn keep_net _zy_sva_guid_miss_aux_cmd_2_30_ccheck
  -- quickturn keep_net _zy_sva_guid_miss_aux_cmd_2_30_cpass
  -- quickturn keep_net _zy_sva_guid_miss_aux_cmd_3_31_ccheck
  -- quickturn keep_net _zy_sva_guid_miss_aux_cmd_3_31_cpass
  -- quickturn keep_net _zy_sva_guid_miss_aux_cmd_iv_0_32_ccheck
  -- quickturn keep_net _zy_sva_guid_miss_aux_cmd_iv_0_32_cpass
  -- quickturn keep_net _zy_sva_guid_miss_aux_cmd_iv_1_33_ccheck
  -- quickturn keep_net _zy_sva_guid_miss_aux_cmd_iv_1_33_cpass
  -- quickturn keep_net _zy_sva_guid_miss_aux_cmd_iv_2_34_ccheck
  -- quickturn keep_net _zy_sva_guid_miss_aux_cmd_iv_2_34_cpass
  -- quickturn keep_net _zy_sva_guid_miss_aux_cmd_iv_3_35_ccheck
  -- quickturn keep_net _zy_sva_guid_miss_aux_cmd_iv_3_35_cpass
  -- quickturn keep_net _zy_sva_iv_miss_aux_cmd_0_36_ccheck
  -- quickturn keep_net _zy_sva_iv_miss_aux_cmd_0_36_cpass
  -- quickturn keep_net _zy_sva_iv_miss_aux_cmd_1_37_ccheck
  -- quickturn keep_net _zy_sva_iv_miss_aux_cmd_1_37_cpass
  -- quickturn keep_net _zy_sva_iv_miss_aux_cmd_guid_38_ccheck
  -- quickturn keep_net _zy_sva_iv_miss_aux_cmd_guid_38_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_39_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_39_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_iv_40_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_iv_40_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_41_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_41_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_42_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_42_cpass
  -- quickturn keep_net _zy_sva_brcm_key_type_43_ccheck
  -- quickturn keep_net _zy_sva_brcm_key_type_43_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_44_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_44_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_iv_45_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_iv_45_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_46_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_46_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_47_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_47_cpass
  -- quickturn keep_net _zy_sva_brcm_key_type_48_ccheck
  -- quickturn keep_net _zy_sva_brcm_key_type_48_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_49_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_49_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_iv_50_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_iv_50_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_51_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_51_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_52_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_52_cpass
  -- quickturn keep_net _zy_sva_brcm_key_type_53_ccheck
  -- quickturn keep_net _zy_sva_brcm_key_type_53_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_54_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_54_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_iv_55_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_iv_55_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_56_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_56_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_57_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_57_cpass
  -- quickturn keep_net _zy_sva_brcm_key_type_58_ccheck
  -- quickturn keep_net _zy_sva_brcm_key_type_58_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_59_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_59_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_iv_60_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_iv_60_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_61_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_61_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_62_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_62_cpass
  -- quickturn keep_net _zy_sva_brcm_key_type_63_ccheck
  -- quickturn keep_net _zy_sva_brcm_key_type_63_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_64_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_64_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_iv_65_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_iv_65_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_66_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_66_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_67_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_67_cpass
  -- quickturn keep_net _zy_sva_brcm_key_type_68_ccheck
  -- quickturn keep_net _zy_sva_brcm_key_type_68_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_69_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_69_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_iv_70_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_iv_70_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_71_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_71_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_72_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_72_cpass
  -- quickturn keep_net _zy_sva_brcm_key_type_73_ccheck
  -- quickturn keep_net _zy_sva_brcm_key_type_73_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_74_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_74_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_iv_75_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_iv_75_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_76_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_76_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_77_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_77_cpass
  -- quickturn keep_net _zy_sva_brcm_key_type_78_ccheck
  -- quickturn keep_net _zy_sva_brcm_key_type_78_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_79_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_79_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_iv_80_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_iv_80_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_81_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_81_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_82_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_82_cpass
  -- quickturn keep_net _zy_sva_brcm_key_type_83_ccheck
  -- quickturn keep_net _zy_sva_brcm_key_type_83_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_84_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_84_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_iv_85_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_iv_85_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_86_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_86_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_87_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_87_cpass
  -- quickturn keep_net _zy_sva_brcm_key_type_88_ccheck
  -- quickturn keep_net _zy_sva_brcm_key_type_88_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_89_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_89_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_iv_90_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_iv_90_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_91_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_91_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_92_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_92_cpass
  -- quickturn keep_net _zy_sva_brcm_key_type_93_ccheck
  -- quickturn keep_net _zy_sva_brcm_key_type_93_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_94_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_94_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_iv_95_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_iv_95_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_96_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_96_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_97_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_97_cpass
  -- quickturn keep_net _zy_sva_brcm_key_type_98_ccheck
  -- quickturn keep_net _zy_sva_brcm_key_type_98_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_99_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_99_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_iv_100_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_iv_100_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_101_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_101_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_102_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_102_cpass
  -- quickturn keep_net _zy_sva_brcm_key_type_103_ccheck
  -- quickturn keep_net _zy_sva_brcm_key_type_103_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_104_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_104_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_iv_105_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_iv_105_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_106_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_106_cpass
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_107_ccheck
  -- quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_107_cpass
  -- quickturn keep_net _zy_sva_brcm_key_type_108_ccheck
  -- quickturn keep_net _zy_sva_brcm_key_type_108_cpass
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_109_ccheck
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_109_cpass
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_110_ccheck
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_110_cpass
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_111_ccheck
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_111_cpass
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_112_ccheck
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_112_cpass
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_113_ccheck
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_113_cpass
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_114_ccheck
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_114_cpass
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_115_ccheck
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_115_cpass
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_116_ccheck
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_116_cpass
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_117_ccheck
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_117_cpass
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_118_ccheck
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_118_cpass
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_119_ccheck
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_119_cpass
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_120_ccheck
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_120_cpass
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_121_ccheck
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_121_cpass
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_122_ccheck
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_122_cpass
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_123_ccheck
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_123_cpass
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_124_ccheck
  -- quickturn keep_net _zy_sva_brcm_kdf_ops_124_cpass
  -- quickturn keep_net _zy_sva_null_gcm_125_ccheck
  -- quickturn keep_net _zy_sva_null_gcm_125_cpass
  -- quickturn keep_net _zy_sva_sha_gcm_126_ccheck
  -- quickturn keep_net _zy_sva_sha_gcm_126_cpass
  -- quickturn keep_net _zy_sva_null_xts_127_ccheck
  -- quickturn keep_net _zy_sva_null_xts_127_cpass
  -- quickturn keep_net _zy_sva_sha_xts_128_ccheck
  -- quickturn keep_net _zy_sva_sha_xts_128_cpass
  -- quickturn keep_net _zy_sva_null_null_129_ccheck
  -- quickturn keep_net _zy_sva_null_null_129_cpass
  -- quickturn keep_net _zy_sva_sha_null_130_ccheck
  -- quickturn keep_net _zy_sva_sha_null_130_cpass
  -- quickturn keep_net _zy_sva_hmac_gcm_131_ccheck
  -- quickturn keep_net _zy_sva_hmac_gcm_131_cpass
  -- quickturn keep_net _zy_sva_hmac_xts_132_ccheck
  -- quickturn keep_net _zy_sva_hmac_xts_132_cpass
  -- quickturn keep_net _zy_sva_hmac_null_133_ccheck
  -- quickturn keep_net _zy_sva_hmac_null_133_cpass
  -- quickturn keep_net _zy_sva_null_gcm_134_ccheck
  -- quickturn keep_net _zy_sva_null_gcm_134_cpass
  -- quickturn keep_net _zy_sva_sha_gcm_135_ccheck
  -- quickturn keep_net _zy_sva_sha_gcm_135_cpass
  -- quickturn keep_net _zy_sva_null_xts_136_ccheck
  -- quickturn keep_net _zy_sva_null_xts_136_cpass
  -- quickturn keep_net _zy_sva_sha_xts_137_ccheck
  -- quickturn keep_net _zy_sva_sha_xts_137_cpass
  -- quickturn keep_net _zy_sva_null_null_138_ccheck
  -- quickturn keep_net _zy_sva_null_null_138_cpass
  -- quickturn keep_net _zy_sva_sha_null_139_ccheck
  -- quickturn keep_net _zy_sva_sha_null_139_cpass
  -- quickturn keep_net _zy_sva_hmac_gcm_140_ccheck
  -- quickturn keep_net _zy_sva_hmac_gcm_140_cpass
  -- quickturn keep_net _zy_sva_hmac_xts_141_ccheck
  -- quickturn keep_net _zy_sva_hmac_xts_141_cpass
  -- quickturn keep_net _zy_sva_hmac_null_142_ccheck
  -- quickturn keep_net _zy_sva_hmac_null_142_cpass
  -- quickturn keep_net _zy_sva_null_gcm_143_ccheck
  -- quickturn keep_net _zy_sva_null_gcm_143_cpass
  -- quickturn keep_net _zy_sva_sha_gcm_144_ccheck
  -- quickturn keep_net _zy_sva_sha_gcm_144_cpass
  -- quickturn keep_net _zy_sva_null_xts_145_ccheck
  -- quickturn keep_net _zy_sva_null_xts_145_cpass
  -- quickturn keep_net _zy_sva_sha_xts_146_ccheck
  -- quickturn keep_net _zy_sva_sha_xts_146_cpass
  -- quickturn keep_net _zy_sva_null_null_147_ccheck
  -- quickturn keep_net _zy_sva_null_null_147_cpass
  -- quickturn keep_net _zy_sva_sha_null_148_ccheck
  -- quickturn keep_net _zy_sva_sha_null_148_cpass
  -- quickturn keep_net _zy_sva_hmac_gcm_149_ccheck
  -- quickturn keep_net _zy_sva_hmac_gcm_149_cpass
  -- quickturn keep_net _zy_sva_hmac_xts_150_ccheck
  -- quickturn keep_net _zy_sva_hmac_xts_150_cpass
  -- quickturn keep_net _zy_sva_hmac_null_151_ccheck
  -- quickturn keep_net _zy_sva_hmac_null_151_cpass
  -- quickturn keep_net _zy_sva_null_gcm_152_ccheck
  -- quickturn keep_net _zy_sva_null_gcm_152_cpass
  -- quickturn keep_net _zy_sva_sha_gcm_153_ccheck
  -- quickturn keep_net _zy_sva_sha_gcm_153_cpass
  -- quickturn keep_net _zy_sva_null_xts_154_ccheck
  -- quickturn keep_net _zy_sva_null_xts_154_cpass
  -- quickturn keep_net _zy_sva_sha_xts_155_ccheck
  -- quickturn keep_net _zy_sva_sha_xts_155_cpass
  -- quickturn keep_net _zy_sva_null_null_156_ccheck
  -- quickturn keep_net _zy_sva_null_null_156_cpass
  -- quickturn keep_net _zy_sva_sha_null_157_ccheck
  -- quickturn keep_net _zy_sva_sha_null_157_cpass
  -- quickturn keep_net _zy_sva_hmac_gcm_158_ccheck
  -- quickturn keep_net _zy_sva_hmac_gcm_158_cpass
  -- quickturn keep_net _zy_sva_hmac_xts_159_ccheck
  -- quickturn keep_net _zy_sva_hmac_xts_159_cpass
  -- quickturn keep_net _zy_sva_hmac_null_160_ccheck
  -- quickturn keep_net _zy_sva_hmac_null_160_cpass
  -- quickturn keep_net _zy_sva_null_gcm_161_ccheck
  -- quickturn keep_net _zy_sva_null_gcm_161_cpass
  -- quickturn keep_net _zy_sva_sha_gcm_162_ccheck
  -- quickturn keep_net _zy_sva_sha_gcm_162_cpass
  -- quickturn keep_net _zy_sva_null_xts_163_ccheck
  -- quickturn keep_net _zy_sva_null_xts_163_cpass
  -- quickturn keep_net _zy_sva_sha_xts_164_ccheck
  -- quickturn keep_net _zy_sva_sha_xts_164_cpass
  -- quickturn keep_net _zy_sva_null_null_165_ccheck
  -- quickturn keep_net _zy_sva_null_null_165_cpass
  -- quickturn keep_net _zy_sva_sha_null_166_ccheck
  -- quickturn keep_net _zy_sva_sha_null_166_cpass
  -- quickturn keep_net _zy_sva_hmac_gcm_167_ccheck
  -- quickturn keep_net _zy_sva_hmac_gcm_167_cpass
  -- quickturn keep_net _zy_sva_hmac_xts_168_ccheck
  -- quickturn keep_net _zy_sva_hmac_xts_168_cpass
  -- quickturn keep_net _zy_sva_hmac_null_169_ccheck
  -- quickturn keep_net _zy_sva_hmac_null_169_cpass
  -- quickturn keep_net _zy_sva_null_gcm_170_ccheck
  -- quickturn keep_net _zy_sva_null_gcm_170_cpass
  -- quickturn keep_net _zy_sva_sha_gcm_171_ccheck
  -- quickturn keep_net _zy_sva_sha_gcm_171_cpass
  -- quickturn keep_net _zy_sva_null_xts_172_ccheck
  -- quickturn keep_net _zy_sva_null_xts_172_cpass
  -- quickturn keep_net _zy_sva_sha_xts_173_ccheck
  -- quickturn keep_net _zy_sva_sha_xts_173_cpass
  -- quickturn keep_net _zy_sva_null_null_174_ccheck
  -- quickturn keep_net _zy_sva_null_null_174_cpass
  -- quickturn keep_net _zy_sva_sha_null_175_ccheck
  -- quickturn keep_net _zy_sva_sha_null_175_cpass
  -- quickturn keep_net _zy_sva_hmac_gcm_176_ccheck
  -- quickturn keep_net _zy_sva_hmac_gcm_176_cpass
  -- quickturn keep_net _zy_sva_hmac_xts_177_ccheck
  -- quickturn keep_net _zy_sva_hmac_xts_177_cpass
  -- quickturn keep_net _zy_sva_hmac_null_178_ccheck
  -- quickturn keep_net _zy_sva_hmac_null_178_cpass

begin
  stitcher_sot <= boolean_to_std(stitcher_out(64+7 downto 64) =
   std_logic_vector'("00000001")) ;
  stitcher_eot <= boolean_to_std(stitcher_out(64+7 downto 64) =
   std_logic_vector'("00000010")) ;
  tlv_parser_idle <= (stitcher_empty and boolean_to_std(tlv_counter =
   std_logic_vector'("00000"))) ;
  tlv_parser_int_tlv_start_pulse <= (fifo_in_valid and it_conv_std_logic(fifo_in
  (70 downto 70))) ;
  _zz_strnp_0 : ixc_assign
    generic map(W => 1)
    port map (
       DUMMY2
      ,stitcher_rd
    ) ;
  _zz_strnp_1 : ixc_assign
    generic map(W => 71)
    port map (
       DUMMY3
      ,parser_kimreader_data
    ) ;
  _zz_strnp_2 : ixc_assign
    generic map(W => 71)
    port map (
       parser_kimreader_data
      ,DUMMY4
    ) ;
  _zz_strnp_3 : ixc_assign
    generic map(W => 71)
    port map (
       DUMMY5
      ,fifo_in
    ) ;
  _zz_strnp_4 : ixc_assign
    generic map(W => 1)
    port map (
       DUMMY6
      ,fifo_in_valid
    ) ;
  _zy_simnet_cio_7 <= '0' ;
  _zy_sva_key_type0_line4_1_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_key_type0_line5a_2_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_key_type0_line5b_3_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_key_type1_line7a_4_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_key_type1_line7b_5_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_key_type1_line8a_6_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_key_type1_line8b_7_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_key_type1_line9_8_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_key_type1_line10_9_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_key_type1_line11a_10_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_key_type1_line11b_11_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_key_type1_line11c_12_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_key_type1_line11d_13_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_key_type1_line12a_14_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_key_type1_line12b_15_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_key_type9_line14_16_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_key_type9_line15_17_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_key_type9_line16a_18_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_key_type9_line16b_19_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_key_type9_line17a_20_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_key_type9_line17b_21_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_key_type9_line18a_22_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_key_type9_line18b_23_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_key_type9_line19a_24_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_key_type9_line19b_25_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_key_type9_line19c_26_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_key_type9_line19d_27_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_guid_miss_aux_cmd_0_28_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_guid_miss_aux_cmd_1_29_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_guid_miss_aux_cmd_2_30_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_guid_miss_aux_cmd_3_31_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_guid_miss_aux_cmd_iv_0_32_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_guid_miss_aux_cmd_iv_1_33_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_guid_miss_aux_cmd_iv_2_34_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_guid_miss_aux_cmd_iv_3_35_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_iv_miss_aux_cmd_0_36_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_iv_miss_aux_cmd_1_37_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_iv_miss_aux_cmd_guid_38_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_39_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_iv_40_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_guid_41_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_guid_iv_42_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_key_type_43_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_44_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_iv_45_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_guid_46_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_guid_iv_47_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_key_type_48_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_49_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_iv_50_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_guid_51_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_guid_iv_52_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_key_type_53_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_54_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_iv_55_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_guid_56_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_guid_iv_57_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_key_type_58_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_59_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_iv_60_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_guid_61_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_guid_iv_62_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_key_type_63_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_64_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_iv_65_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_guid_66_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_guid_iv_67_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_key_type_68_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_69_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_iv_70_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_guid_71_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_guid_iv_72_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_key_type_73_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_74_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_iv_75_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_guid_76_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_guid_iv_77_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_key_type_78_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_79_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_iv_80_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_guid_81_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_guid_iv_82_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_key_type_83_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_84_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_iv_85_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_guid_86_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_guid_iv_87_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_key_type_88_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_89_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_iv_90_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_guid_91_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_guid_iv_92_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_key_type_93_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_94_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_iv_95_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_guid_96_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_guid_iv_97_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_key_type_98_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_99_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_iv_100_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_guid_101_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_guid_iv_102_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_key_type_103_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_104_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_iv_105_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_guid_106_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_aux_cmd_guid_iv_107_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_key_type_108_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_kdf_ops_109_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_kdf_ops_110_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_kdf_ops_111_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_kdf_ops_112_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_kdf_ops_113_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_kdf_ops_114_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_kdf_ops_115_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_kdf_ops_116_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_kdf_ops_117_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_kdf_ops_118_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_kdf_ops_119_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_kdf_ops_120_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_kdf_ops_121_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_kdf_ops_122_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_kdf_ops_123_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_brcm_kdf_ops_124_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_null_gcm_125_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_sha_gcm_126_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_null_xts_127_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_sha_xts_128_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_null_null_129_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_sha_null_130_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_hmac_gcm_131_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_hmac_xts_132_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_hmac_null_133_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_null_gcm_134_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_sha_gcm_135_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_null_xts_136_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_sha_xts_137_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_null_null_138_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_sha_null_139_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_hmac_gcm_140_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_hmac_xts_141_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_hmac_null_142_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_null_gcm_143_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_sha_gcm_144_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_null_xts_145_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_sha_xts_146_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_null_null_147_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_sha_null_148_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_hmac_gcm_149_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_hmac_xts_150_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_hmac_null_151_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_null_gcm_152_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_sha_gcm_153_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_null_xts_154_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_sha_xts_155_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_null_null_156_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_sha_null_157_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_hmac_gcm_158_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_hmac_xts_159_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_hmac_null_160_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_null_gcm_161_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_sha_gcm_162_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_null_xts_163_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_sha_xts_164_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_null_null_165_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_sha_null_166_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_hmac_gcm_167_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_hmac_xts_168_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_hmac_null_169_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_null_gcm_170_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_sha_gcm_171_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_null_xts_172_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_sha_xts_173_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_null_null_174_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_sha_null_175_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_hmac_gcm_176_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_hmac_xts_177_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_hmac_null_178_reset_or <= boolean_to_std(ext(rst_n,32) /=
   std_logic_vector'("00000000000000000000000000000001")) ;
  _zy_sva_b0_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and 
  (aux_auth_op = HMAC_SHA2 or aux_raw_auth_op = HMAC_SHA2) and aux_cipher_op =
   CPH_NULL and aux_key_type = NO_AUX_KEY)) ;
  _zy_sva_b1_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op /= HMAC_SHA2 and aux_raw_auth_op /= HMAC_SHA2 and aux_cipher_op =
   AES_XTS_XEX and aux_key_type = NO_AUX_KEY)) ;
  _zy_sva_b2_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op /= HMAC_SHA2 and aux_raw_auth_op /= HMAC_SHA2 and aux_cipher_op =
   AES_GCM and aux_key_type = NO_AUX_KEY)) ;
  _zy_sva_b3_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = AUTH_NULL and aux_raw_auth_op = AUTH_NULL and aux_cipher_op =
   CPH_NULL and aux_key_type = AUX_KEY_ONLY and aux_key_header(15+1 downto 15)
   /= KDF_MODE_COMB_GUID and aux_key_header(15+1 downto 15) /=
   KDF_MODE_COMB_RGUID)) ;
  _zy_sva_b4_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = SHA2 and aux_raw_auth_op = SHA2 and aux_cipher_op = CPH_NULL
   and aux_key_type = AUX_KEY_ONLY and aux_key_header(15+1 downto 15) /=
   KDF_MODE_COMB_GUID and aux_key_header(15+1 downto 15) /= KDF_MODE_COMB_RGUID)
  ) ;
  _zy_sva_b5_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = AUTH_NULL and aux_raw_auth_op = AUTH_NULL and aux_cipher_op =
   CPH_NULL and aux_key_type = AUX_KEY_ONLY and (aux_key_header(15+1 downto 15)
   = KDF_MODE_COMB_GUID or aux_key_header(15+1 downto 15) = KDF_MODE_COMB_RGUID)
  )) ;
  _zy_sva_b6_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = SHA2 and aux_raw_auth_op = SHA2 and aux_cipher_op = CPH_NULL
   and aux_key_type = AUX_KEY_ONLY and (aux_key_header(15+1 downto 15) =
   KDF_MODE_COMB_GUID or aux_key_header(15+1 downto 15) = KDF_MODE_COMB_RGUID)))
   ;
  _zy_sva_b7_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = HMAC_SHA2 and aux_raw_auth_op = HMAC_SHA2 and aux_cipher_op =
   CPH_NULL and aux_key_type = AUX_KEY_ONLY and aux_key_header(15+1 downto 15)
   /= KDF_MODE_COMB_GUID and aux_key_header(15+1 downto 15) /=
   KDF_MODE_COMB_RGUID)) ;
  _zy_sva_b8_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = HMAC_SHA2 and aux_raw_auth_op = HMAC_SHA2 and aux_cipher_op =
   CPH_NULL and aux_key_type = AUX_KEY_ONLY and (aux_key_header(15+1 downto 15)
   = KDF_MODE_COMB_GUID or aux_key_header(15+1 downto 15) = KDF_MODE_COMB_RGUID)
  )) ;
  _zy_sva_b9_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = AUTH_NULL and aux_raw_auth_op = AUTH_NULL and aux_cipher_op =
   AES_GCM and aux_key_type = AUX_KEY_ONLY)) ;
  _zy_sva_b10_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = AUTH_NULL and aux_raw_auth_op = AUTH_NULL and aux_cipher_op =
   AES_XTS_XEX and aux_key_type = AUX_KEY_ONLY)) ;
  _zy_sva_b11_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = SHA2 and aux_raw_auth_op = SHA2 and aux_cipher_op = AES_GCM and
   aux_key_type = AUX_KEY_ONLY)) ;
  _zy_sva_b12_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = SHA2 and aux_raw_auth_op = SHA2 and aux_cipher_op = AES_XTS_XEX
   and aux_key_type = AUX_KEY_ONLY)) ;
  _zy_sva_b13_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = HMAC_SHA2 and aux_raw_auth_op = HMAC_SHA2 and aux_cipher_op =
   AES_GCM and aux_key_type = AUX_KEY_ONLY)) ;
  _zy_sva_b14_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = HMAC_SHA2 and aux_raw_auth_op = HMAC_SHA2 and aux_cipher_op =
   AES_XTS_XEX and aux_key_type = AUX_KEY_ONLY)) ;
  _zy_sva_b15_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = HMAC_SHA2 and aux_raw_auth_op = HMAC_SHA2 and aux_cipher_op =
   CPH_NULL and aux_key_type = ENC_DAK and aux_key_header(15+1 downto 15) /=
   KDF_MODE_COMB_GUID and aux_key_header(15+1 downto 15) /= KDF_MODE_COMB_RGUID)
  ) ;
  _zy_sva_b16_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = HMAC_SHA2 and aux_raw_auth_op = HMAC_SHA2 and aux_cipher_op =
   CPH_NULL and aux_key_type = ENC_DAK and (aux_key_header(15+1 downto 15) =
   KDF_MODE_COMB_GUID or aux_key_header(15+1 downto 15) = KDF_MODE_COMB_RGUID)))
   ;
  _zy_sva_b17_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = HMAC_SHA2 and aux_raw_auth_op = HMAC_SHA2 and aux_cipher_op =
   AES_GCM and aux_key_type = ENC_DAK)) ;
  _zy_sva_b18_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = HMAC_SHA2 and aux_raw_auth_op = HMAC_SHA2 and aux_cipher_op =
   AES_XTS_XEX and aux_key_type = ENC_DAK)) ;
  _zy_sva_b19_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = AUTH_NULL and aux_raw_auth_op = AUTH_NULL and aux_cipher_op =
   CPH_NULL and aux_key_type = ENC_DAK and aux_key_header(15+1 downto 15) /=
   KDF_MODE_COMB_GUID and aux_key_header(15+1 downto 15) /= KDF_MODE_COMB_RGUID)
  ) ;
  _zy_sva_b20_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = SHA2 and aux_raw_auth_op = SHA2 and aux_cipher_op = CPH_NULL
   and aux_key_type = ENC_DAK and aux_key_header(15+1 downto 15) /=
   KDF_MODE_COMB_GUID and aux_key_header(15+1 downto 15) /= KDF_MODE_COMB_RGUID)
  ) ;
  _zy_sva_b21_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = AUTH_NULL and aux_raw_auth_op = AUTH_NULL and aux_cipher_op =
   CPH_NULL and aux_key_type = ENC_DAK and (aux_key_header(15+1 downto 15) =
   KDF_MODE_COMB_GUID or aux_key_header(15+1 downto 15) = KDF_MODE_COMB_RGUID)))
   ;
  _zy_sva_b22_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = SHA2 and aux_raw_auth_op = SHA2 and aux_cipher_op = CPH_NULL
   and aux_key_type = ENC_DAK and (aux_key_header(15+1 downto 15) =
   KDF_MODE_COMB_GUID or aux_key_header(15+1 downto 15) = KDF_MODE_COMB_RGUID)))
   ;
  _zy_sva_b23_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = AUTH_NULL and aux_raw_auth_op = AUTH_NULL and aux_cipher_op =
   AES_GCM and aux_key_type = ENC_DAK)) ;
  _zy_sva_b24_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = SHA2 and aux_raw_auth_op = SHA2 and aux_cipher_op = AES_GCM and
   aux_key_type = ENC_DAK)) ;
  _zy_sva_b25_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = AUTH_NULL and aux_raw_auth_op = AUTH_NULL and aux_cipher_op =
   AES_XTS_XEX and aux_key_type = ENC_DAK)) ;
  _zy_sva_b26_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = SHA2 and aux_raw_auth_op = SHA2 and aux_cipher_op = AES_XTS_XEX
   and aux_key_type = ENC_DAK)) ;
  _zy_sva_b27_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   tlv_type = AUX_CMD and aux_key_header(15+1 downto 15) = KDF_MODE_GUID and
   aux_key_header(14 downto 14) = KDF and aux_key_header(31 downto 31) = NOOP))
   ;
  _zy_sva_b28_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   tlv_type = AUX_CMD and aux_key_header(15+1 downto 15) = KDF_MODE_GUID and
   aux_key_header(14 downto 14) = NOOP and aux_key_header(31 downto 31) = KDF))
   ;
  _zy_sva_b29_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   tlv_type = AUX_CMD and aux_key_header(15+1 downto 15) = KDF_MODE_COMB_GUID
   and aux_key_header(14 downto 14) = KDF and aux_key_header(31 downto 31) =
   NOOP)) ;
  _zy_sva_b30_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   tlv_type = AUX_CMD and aux_key_header(15+1 downto 15) = KDF_MODE_COMB_GUID
   and aux_key_header(14 downto 14) = NOOP and aux_key_header(31 downto 31) =
   KDF)) ;
  _zy_sva_b31_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   tlv_type = AUX_CMD_IV and aux_key_header(15+1 downto 15) = KDF_MODE_GUID and
   aux_key_header(14 downto 14) = KDF and aux_key_header(31 downto 31) = NOOP))
   ;
  _zy_sva_b32_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   tlv_type = AUX_CMD_IV and aux_key_header(15+1 downto 15) = KDF_MODE_GUID and
   aux_key_header(14 downto 14) = NOOP and aux_key_header(31 downto 31) = KDF))
   ;
  _zy_sva_b33_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   tlv_type = AUX_CMD_IV and aux_key_header(15+1 downto 15) = KDF_MODE_COMB_GUID
   and aux_key_header(14 downto 14) = KDF and aux_key_header(31 downto 31) =
   NOOP)) ;
  _zy_sva_b34_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   tlv_type = AUX_CMD_IV and aux_key_header(15+1 downto 15) = KDF_MODE_COMB_GUID
   and aux_key_header(14 downto 14) = NOOP and aux_key_header(31 downto 31) =
   KDF)) ;
  _zy_sva_b35_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   tlv_type = AUX_CMD and aux_iv_op = IV_INC and aux_cipher_op = AES_GCM)) ;
  _zy_sva_b36_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   tlv_type = AUX_CMD and aux_iv_op = IV_INC and aux_cipher_op = AES_XTS_XEX)) ;
  _zy_sva_b37_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   tlv_type = AUX_CMD_GUID and aux_iv_op = IV_INC and aux_cipher_op =
   AES_XTS_XEX)) ;
  _zy_sva_b38_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000010101"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000000"))) ;
  _zy_sva_b39_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000010111"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000000"))) ;
  _zy_sva_b40_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000011000"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000000"))) ;
  _zy_sva_b41_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000011001"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000000"))) ;
  _zy_sva_b42_t <= ((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_word2(57+5 downto 57),32) =
   std_logic_vector'("00000000000000000000000000000000"))) ;
  _zy_sva_b43_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000010101"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000001"))) ;
  _zy_sva_b44_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000010111"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000001"))) ;
  _zy_sva_b45_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000011000"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000001"))) ;
  _zy_sva_b46_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000011001"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000001"))) ;
  _zy_sva_b47_t <= ((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_word2(57+5 downto 57),32) =
   std_logic_vector'("00000000000000000000000000000001"))) ;
  _zy_sva_b48_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000010101"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000010"))) ;
  _zy_sva_b49_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000010111"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000010"))) ;
  _zy_sva_b50_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000011000"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000010"))) ;
  _zy_sva_b51_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000011001"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000010"))) ;
  _zy_sva_b52_t <= ((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_word2(57+5 downto 57),32) =
   std_logic_vector'("00000000000000000000000000000010"))) ;
  _zy_sva_b53_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000010101"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000011"))) ;
  _zy_sva_b54_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000010111"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000011"))) ;
  _zy_sva_b55_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000011000"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000011"))) ;
  _zy_sva_b56_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000011001"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000011"))) ;
  _zy_sva_b57_t <= ((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_word2(57+5 downto 57),32) =
   std_logic_vector'("00000000000000000000000000000011"))) ;
  _zy_sva_b58_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000010101"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000100"))) ;
  _zy_sva_b59_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000010111"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000100"))) ;
  _zy_sva_b60_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000011000"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000100"))) ;
  _zy_sva_b61_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000011001"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000100"))) ;
  _zy_sva_b62_t <= ((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_word2(57+5 downto 57),32) =
   std_logic_vector'("00000000000000000000000000000100"))) ;
  _zy_sva_b63_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000010101"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000101"))) ;
  _zy_sva_b64_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000010111"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000101"))) ;
  _zy_sva_b65_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000011000"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000101"))) ;
  _zy_sva_b66_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000011001"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000101"))) ;
  _zy_sva_b67_t <= ((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_word2(57+5 downto 57),32) =
   std_logic_vector'("00000000000000000000000000000101"))) ;
  _zy_sva_b68_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000010101"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000110"))) ;
  _zy_sva_b69_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000010111"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000110"))) ;
  _zy_sva_b70_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000011000"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000110"))) ;
  _zy_sva_b71_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000011001"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000110"))) ;
  _zy_sva_b72_t <= ((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_word2(57+5 downto 57),32) =
   std_logic_vector'("00000000000000000000000000000110"))) ;
  _zy_sva_b73_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000010101"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000111"))) ;
  _zy_sva_b74_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000010111"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000111"))) ;
  _zy_sva_b75_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000011000"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000111"))) ;
  _zy_sva_b76_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000011001"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000000111"))) ;
  _zy_sva_b77_t <= ((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_word2(57+5 downto 57),32) =
   std_logic_vector'("00000000000000000000000000000111"))) ;
  _zy_sva_b78_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000010101"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000001000"))) ;
  _zy_sva_b79_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000010111"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000001000"))) ;
  _zy_sva_b80_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000011000"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000001000"))) ;
  _zy_sva_b81_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000011001"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000001000"))) ;
  _zy_sva_b82_t <= ((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_word2(57+5 downto 57),32) =
   std_logic_vector'("00000000000000000000000000001000"))) ;
  _zy_sva_b83_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000010101"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000001001"))) ;
  _zy_sva_b84_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000010111"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000001001"))) ;
  _zy_sva_b85_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000011000"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000001001"))) ;
  _zy_sva_b86_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000011001"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000001001"))) ;
  _zy_sva_b87_t <= ((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_word2(57+5 downto 57),32) =
   std_logic_vector'("00000000000000000000000000001001"))) ;
  _zy_sva_b88_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000010101"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000001010"))) ;
  _zy_sva_b89_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000010111"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000001010"))) ;
  _zy_sva_b90_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000011000"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000001010"))) ;
  _zy_sva_b91_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000011001"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000001010"))) ;
  _zy_sva_b92_t <= ((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_word2(57+5 downto 57),32) =
   std_logic_vector'("00000000000000000000000000001010"))) ;
  _zy_sva_b93_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000010101"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000001011"))) ;
  _zy_sva_b94_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000010111"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000001011"))) ;
  _zy_sva_b95_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000011000"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000001011"))) ;
  _zy_sva_b96_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000011001"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000001011"))) ;
  _zy_sva_b97_t <= ((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_word2(57+5 downto 57),32) =
   std_logic_vector'("00000000000000000000000000001011"))) ;
  _zy_sva_b98_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000010101"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000001100"))) ;
  _zy_sva_b99_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000010111"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000001100"))) ;
  _zy_sva_b100_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64)
   = KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000011000"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000001100"))) ;
  _zy_sva_b101_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64)
   = KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000011001"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000001100"))) ;
  _zy_sva_b102_t <= ((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_word2(57+5 downto 57),32) =
   std_logic_vector'("00000000000000000000000000001100"))) ;
  _zy_sva_b103_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64)
   = KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000010101"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000001101"))) ;
  _zy_sva_b104_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64)
   = KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000010111"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000001101"))) ;
  _zy_sva_b105_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64)
   = KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000011000"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000001101"))) ;
  _zy_sva_b106_t <= (((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64)
   = KME_WORD0)) and boolean_to_std(ext(tlv_type,32) = std_logic_vector'
  ("00000000000000000000000000011001"))) and boolean_to_std(ext(tlv_word2(57+5
   downto 57),32) = std_logic_vector'("00000000000000000000000000001101"))) ;
  _zy_sva_b107_t <= ((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64) =
   KME_WORD0)) and boolean_to_std(ext(tlv_word2(57+5 downto 57),32) =
   std_logic_vector'("00000000000000000000000000001101"))) ;
  _zy_sva_b108_t <= ((((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64)
   = KME_ERROR)) and boolean_to_std(ext(aux_key_header(15+1 downto 15),32) =
   std_logic_vector'("00000000000000000000000000000000"))) and boolean_to_std
  (ext(aux_key_header(14 downto 14),32) = std_logic_vector'
  ("00000000000000000000000000000000"))) and boolean_to_std(ext(aux_key_header
  (31 downto 31),32) = std_logic_vector'("00000000000000000000000000000000"))) ;
  _zy_sva_b109_t <= ((((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64)
   = KME_ERROR)) and boolean_to_std(ext(aux_key_header(15+1 downto 15),32) =
   std_logic_vector'("00000000000000000000000000000000"))) and boolean_to_std
  (ext(aux_key_header(14 downto 14),32) = std_logic_vector'
  ("00000000000000000000000000000000"))) and boolean_to_std(ext(aux_key_header
  (31 downto 31),32) = std_logic_vector'("00000000000000000000000000000001"))) ;
  _zy_sva_b110_t <= ((((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64)
   = KME_ERROR)) and boolean_to_std(ext(aux_key_header(15+1 downto 15),32) =
   std_logic_vector'("00000000000000000000000000000000"))) and boolean_to_std
  (ext(aux_key_header(14 downto 14),32) = std_logic_vector'
  ("00000000000000000000000000000001"))) and boolean_to_std(ext(aux_key_header
  (31 downto 31),32) = std_logic_vector'("00000000000000000000000000000000"))) ;
  _zy_sva_b111_t <= ((((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64)
   = KME_ERROR)) and boolean_to_std(ext(aux_key_header(15+1 downto 15),32) =
   std_logic_vector'("00000000000000000000000000000000"))) and boolean_to_std
  (ext(aux_key_header(14 downto 14),32) = std_logic_vector'
  ("00000000000000000000000000000001"))) and boolean_to_std(ext(aux_key_header
  (31 downto 31),32) = std_logic_vector'("00000000000000000000000000000001"))) ;
  _zy_sva_b112_t <= ((((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64)
   = KME_ERROR)) and boolean_to_std(ext(aux_key_header(15+1 downto 15),32) =
   std_logic_vector'("00000000000000000000000000000001"))) and boolean_to_std
  (ext(aux_key_header(14 downto 14),32) = std_logic_vector'
  ("00000000000000000000000000000000"))) and boolean_to_std(ext(aux_key_header
  (31 downto 31),32) = std_logic_vector'("00000000000000000000000000000000"))) ;
  _zy_sva_b113_t <= ((((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64)
   = KME_ERROR)) and boolean_to_std(ext(aux_key_header(15+1 downto 15),32) =
   std_logic_vector'("00000000000000000000000000000001"))) and boolean_to_std
  (ext(aux_key_header(14 downto 14),32) = std_logic_vector'
  ("00000000000000000000000000000000"))) and boolean_to_std(ext(aux_key_header
  (31 downto 31),32) = std_logic_vector'("00000000000000000000000000000001"))) ;
  _zy_sva_b114_t <= ((((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64)
   = KME_ERROR)) and boolean_to_std(ext(aux_key_header(15+1 downto 15),32) =
   std_logic_vector'("00000000000000000000000000000001"))) and boolean_to_std
  (ext(aux_key_header(14 downto 14),32) = std_logic_vector'
  ("00000000000000000000000000000001"))) and boolean_to_std(ext(aux_key_header
  (31 downto 31),32) = std_logic_vector'("00000000000000000000000000000000"))) ;
  _zy_sva_b115_t <= ((((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64)
   = KME_ERROR)) and boolean_to_std(ext(aux_key_header(15+1 downto 15),32) =
   std_logic_vector'("00000000000000000000000000000001"))) and boolean_to_std
  (ext(aux_key_header(14 downto 14),32) = std_logic_vector'
  ("00000000000000000000000000000001"))) and boolean_to_std(ext(aux_key_header
  (31 downto 31),32) = std_logic_vector'("00000000000000000000000000000001"))) ;
  _zy_sva_b116_t <= ((((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64)
   = KME_ERROR)) and boolean_to_std(ext(aux_key_header(15+1 downto 15),32) =
   std_logic_vector'("00000000000000000000000000000010"))) and boolean_to_std
  (ext(aux_key_header(14 downto 14),32) = std_logic_vector'
  ("00000000000000000000000000000000"))) and boolean_to_std(ext(aux_key_header
  (31 downto 31),32) = std_logic_vector'("00000000000000000000000000000000"))) ;
  _zy_sva_b117_t <= ((((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64)
   = KME_ERROR)) and boolean_to_std(ext(aux_key_header(15+1 downto 15),32) =
   std_logic_vector'("00000000000000000000000000000010"))) and boolean_to_std
  (ext(aux_key_header(14 downto 14),32) = std_logic_vector'
  ("00000000000000000000000000000000"))) and boolean_to_std(ext(aux_key_header
  (31 downto 31),32) = std_logic_vector'("00000000000000000000000000000001"))) ;
  _zy_sva_b118_t <= ((((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64)
   = KME_ERROR)) and boolean_to_std(ext(aux_key_header(15+1 downto 15),32) =
   std_logic_vector'("00000000000000000000000000000010"))) and boolean_to_std
  (ext(aux_key_header(14 downto 14),32) = std_logic_vector'
  ("00000000000000000000000000000001"))) and boolean_to_std(ext(aux_key_header
  (31 downto 31),32) = std_logic_vector'("00000000000000000000000000000000"))) ;
  _zy_sva_b119_t <= ((((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64)
   = KME_ERROR)) and boolean_to_std(ext(aux_key_header(15+1 downto 15),32) =
   std_logic_vector'("00000000000000000000000000000010"))) and boolean_to_std
  (ext(aux_key_header(14 downto 14),32) = std_logic_vector'
  ("00000000000000000000000000000001"))) and boolean_to_std(ext(aux_key_header
  (31 downto 31),32) = std_logic_vector'("00000000000000000000000000000001"))) ;
  _zy_sva_b120_t <= ((((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64)
   = KME_ERROR)) and boolean_to_std(ext(aux_key_header(15+1 downto 15),32) =
   std_logic_vector'("00000000000000000000000000000011"))) and boolean_to_std
  (ext(aux_key_header(14 downto 14),32) = std_logic_vector'
  ("00000000000000000000000000000000"))) and boolean_to_std(ext(aux_key_header
  (31 downto 31),32) = std_logic_vector'("00000000000000000000000000000000"))) ;
  _zy_sva_b121_t <= ((((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64)
   = KME_ERROR)) and boolean_to_std(ext(aux_key_header(15+1 downto 15),32) =
   std_logic_vector'("00000000000000000000000000000011"))) and boolean_to_std
  (ext(aux_key_header(14 downto 14),32) = std_logic_vector'
  ("00000000000000000000000000000000"))) and boolean_to_std(ext(aux_key_header
  (31 downto 31),32) = std_logic_vector'("00000000000000000000000000000001"))) ;
  _zy_sva_b122_t <= ((((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64)
   = KME_ERROR)) and boolean_to_std(ext(aux_key_header(15+1 downto 15),32) =
   std_logic_vector'("00000000000000000000000000000011"))) and boolean_to_std
  (ext(aux_key_header(14 downto 14),32) = std_logic_vector'
  ("00000000000000000000000000000001"))) and boolean_to_std(ext(aux_key_header
  (31 downto 31),32) = std_logic_vector'("00000000000000000000000000000000"))) ;
  _zy_sva_b123_t <= ((((fifo_in_valid and boolean_to_std(fifo_in(64+3 downto 64)
   = KME_ERROR)) and boolean_to_std(ext(aux_key_header(15+1 downto 15),32) =
   std_logic_vector'("00000000000000000000000000000011"))) and boolean_to_std
  (ext(aux_key_header(14 downto 14),32) = std_logic_vector'
  ("00000000000000000000000000000001"))) and boolean_to_std(ext(aux_key_header
  (31 downto 31),32) = std_logic_vector'("00000000000000000000000000000001"))) ;
  _zy_sva_b124_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = AUTH_NULL and aux_raw_auth_op = AUTH_NULL and aux_cipher_op =
   AES_GCM and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000000111"))) ;
  _zy_sva_b125_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = SHA2 and aux_raw_auth_op = SHA2 and aux_cipher_op = AES_GCM and
   ext(aux_key_type,32) = std_logic_vector'("00000000000000000000000000000111"))
  ) ;
  _zy_sva_b126_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = AUTH_NULL and aux_raw_auth_op = AUTH_NULL and aux_cipher_op =
   AES_XTS_XEX and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000000111"))) ;
  _zy_sva_b127_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = SHA2 and aux_raw_auth_op = SHA2 and aux_cipher_op = AES_XTS_XEX
   and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000000111"))) ;
  _zy_sva_b128_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = AUTH_NULL and aux_raw_auth_op = AUTH_NULL and aux_cipher_op =
   CPH_NULL and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000000111"))) ;
  _zy_sva_b129_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = SHA2 and aux_raw_auth_op = SHA2 and aux_cipher_op = CPH_NULL
   and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000000111"))) ;
  _zy_sva_b130_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = HMAC_SHA2 and aux_raw_auth_op = HMAC_SHA2 and aux_cipher_op =
   AES_GCM and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000000111"))) ;
  _zy_sva_b131_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = HMAC_SHA2 and aux_raw_auth_op = HMAC_SHA2 and aux_cipher_op =
   AES_XTS_XEX and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000000111"))) ;
  _zy_sva_b132_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = HMAC_SHA2 and aux_raw_auth_op = HMAC_SHA2 and aux_cipher_op =
   CPH_NULL and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000000111"))) ;
  _zy_sva_b133_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = AUTH_NULL and aux_raw_auth_op = AUTH_NULL and aux_cipher_op =
   AES_GCM and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001000"))) ;
  _zy_sva_b134_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = SHA2 and aux_raw_auth_op = SHA2 and aux_cipher_op = AES_GCM and
   ext(aux_key_type,32) = std_logic_vector'("00000000000000000000000000001000"))
  ) ;
  _zy_sva_b135_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = AUTH_NULL and aux_raw_auth_op = AUTH_NULL and aux_cipher_op =
   AES_XTS_XEX and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001000"))) ;
  _zy_sva_b136_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = SHA2 and aux_raw_auth_op = SHA2 and aux_cipher_op = AES_XTS_XEX
   and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001000"))) ;
  _zy_sva_b137_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = AUTH_NULL and aux_raw_auth_op = AUTH_NULL and aux_cipher_op =
   CPH_NULL and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001000"))) ;
  _zy_sva_b138_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = SHA2 and aux_raw_auth_op = SHA2 and aux_cipher_op = CPH_NULL
   and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001000"))) ;
  _zy_sva_b139_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = HMAC_SHA2 and aux_raw_auth_op = HMAC_SHA2 and aux_cipher_op =
   AES_GCM and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001000"))) ;
  _zy_sva_b140_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = HMAC_SHA2 and aux_raw_auth_op = HMAC_SHA2 and aux_cipher_op =
   AES_XTS_XEX and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001000"))) ;
  _zy_sva_b141_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = HMAC_SHA2 and aux_raw_auth_op = HMAC_SHA2 and aux_cipher_op =
   CPH_NULL and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001000"))) ;
  _zy_sva_b142_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = AUTH_NULL and aux_raw_auth_op = AUTH_NULL and aux_cipher_op =
   AES_GCM and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001010"))) ;
  _zy_sva_b143_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = SHA2 and aux_raw_auth_op = SHA2 and aux_cipher_op = AES_GCM and
   ext(aux_key_type,32) = std_logic_vector'("00000000000000000000000000001010"))
  ) ;
  _zy_sva_b144_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = AUTH_NULL and aux_raw_auth_op = AUTH_NULL and aux_cipher_op =
   AES_XTS_XEX and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001010"))) ;
  _zy_sva_b145_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = SHA2 and aux_raw_auth_op = SHA2 and aux_cipher_op = AES_XTS_XEX
   and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001010"))) ;
  _zy_sva_b146_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = AUTH_NULL and aux_raw_auth_op = AUTH_NULL and aux_cipher_op =
   CPH_NULL and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001010"))) ;
  _zy_sva_b147_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = SHA2 and aux_raw_auth_op = SHA2 and aux_cipher_op = CPH_NULL
   and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001010"))) ;
  _zy_sva_b148_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = HMAC_SHA2 and aux_raw_auth_op = HMAC_SHA2 and aux_cipher_op =
   AES_GCM and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001010"))) ;
  _zy_sva_b149_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = HMAC_SHA2 and aux_raw_auth_op = HMAC_SHA2 and aux_cipher_op =
   AES_XTS_XEX and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001010"))) ;
  _zy_sva_b150_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = HMAC_SHA2 and aux_raw_auth_op = HMAC_SHA2 and aux_cipher_op =
   CPH_NULL and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001010"))) ;
  _zy_sva_b151_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = AUTH_NULL and aux_raw_auth_op = AUTH_NULL and aux_cipher_op =
   AES_GCM and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001011"))) ;
  _zy_sva_b152_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = SHA2 and aux_raw_auth_op = SHA2 and aux_cipher_op = AES_GCM and
   ext(aux_key_type,32) = std_logic_vector'("00000000000000000000000000001011"))
  ) ;
  _zy_sva_b153_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = AUTH_NULL and aux_raw_auth_op = AUTH_NULL and aux_cipher_op =
   AES_XTS_XEX and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001011"))) ;
  _zy_sva_b154_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = SHA2 and aux_raw_auth_op = SHA2 and aux_cipher_op = AES_XTS_XEX
   and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001011"))) ;
  _zy_sva_b155_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = AUTH_NULL and aux_raw_auth_op = AUTH_NULL and aux_cipher_op =
   CPH_NULL and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001011"))) ;
  _zy_sva_b156_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = SHA2 and aux_raw_auth_op = SHA2 and aux_cipher_op = CPH_NULL
   and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001011"))) ;
  _zy_sva_b157_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = HMAC_SHA2 and aux_raw_auth_op = HMAC_SHA2 and aux_cipher_op =
   AES_GCM and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001011"))) ;
  _zy_sva_b158_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = HMAC_SHA2 and aux_raw_auth_op = HMAC_SHA2 and aux_cipher_op =
   AES_XTS_XEX and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001011"))) ;
  _zy_sva_b159_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = HMAC_SHA2 and aux_raw_auth_op = HMAC_SHA2 and aux_cipher_op =
   CPH_NULL and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001011"))) ;
  _zy_sva_b160_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = AUTH_NULL and aux_raw_auth_op = AUTH_NULL and aux_cipher_op =
   AES_GCM and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001100"))) ;
  _zy_sva_b161_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = SHA2 and aux_raw_auth_op = SHA2 and aux_cipher_op = AES_GCM and
   ext(aux_key_type,32) = std_logic_vector'("00000000000000000000000000001100"))
  ) ;
  _zy_sva_b162_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = AUTH_NULL and aux_raw_auth_op = AUTH_NULL and aux_cipher_op =
   AES_XTS_XEX and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001100"))) ;
  _zy_sva_b163_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = SHA2 and aux_raw_auth_op = SHA2 and aux_cipher_op = AES_XTS_XEX
   and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001100"))) ;
  _zy_sva_b164_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = AUTH_NULL and aux_raw_auth_op = AUTH_NULL and aux_cipher_op =
   CPH_NULL and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001100"))) ;
  _zy_sva_b165_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = SHA2 and aux_raw_auth_op = SHA2 and aux_cipher_op = CPH_NULL
   and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001100"))) ;
  _zy_sva_b166_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = HMAC_SHA2 and aux_raw_auth_op = HMAC_SHA2 and aux_cipher_op =
   AES_GCM and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001100"))) ;
  _zy_sva_b167_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = HMAC_SHA2 and aux_raw_auth_op = HMAC_SHA2 and aux_cipher_op =
   AES_XTS_XEX and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001100"))) ;
  _zy_sva_b168_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = HMAC_SHA2 and aux_raw_auth_op = HMAC_SHA2 and aux_cipher_op =
   CPH_NULL and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001100"))) ;
  _zy_sva_b169_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = AUTH_NULL and aux_raw_auth_op = AUTH_NULL and aux_cipher_op =
   AES_GCM and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001101"))) ;
  _zy_sva_b170_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = SHA2 and aux_raw_auth_op = SHA2 and aux_cipher_op = AES_GCM and
   ext(aux_key_type,32) = std_logic_vector'("00000000000000000000000000001101"))
  ) ;
  _zy_sva_b171_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = AUTH_NULL and aux_raw_auth_op = AUTH_NULL and aux_cipher_op =
   AES_XTS_XEX and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001101"))) ;
  _zy_sva_b172_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = SHA2 and aux_raw_auth_op = SHA2 and aux_cipher_op = AES_XTS_XEX
   and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001101"))) ;
  _zy_sva_b173_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = AUTH_NULL and aux_raw_auth_op = AUTH_NULL and aux_cipher_op =
   CPH_NULL and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001101"))) ;
  _zy_sva_b174_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = SHA2 and aux_raw_auth_op = SHA2 and aux_cipher_op = CPH_NULL
   and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001101"))) ;
  _zy_sva_b175_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = HMAC_SHA2 and aux_raw_auth_op = HMAC_SHA2 and aux_cipher_op =
   AES_GCM and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001101"))) ;
  _zy_sva_b176_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = HMAC_SHA2 and aux_raw_auth_op = HMAC_SHA2 and aux_cipher_op =
   AES_XTS_XEX and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001101"))) ;
  _zy_sva_b177_t <= boolean_to_std((int_tlv_counter = IDX_KME_IVTWEAK and
   aux_auth_op = HMAC_SHA2 and aux_raw_auth_op = HMAC_SHA2 and aux_cipher_op =
   CPH_NULL and ext(aux_key_type,32) = std_logic_vector'
  ("00000000000000000000000000001101"))) ;
  _zz_zy_sva_b0 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b0
      ,_zy_sva_b0_t
    ) ;
  _zz_zy_sva_b1 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b1
      ,_zy_sva_b1_t
    ) ;
  _zz_zy_sva_b2 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b2
      ,_zy_sva_b2_t
    ) ;
  _zz_zy_sva_b3 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b3
      ,_zy_sva_b3_t
    ) ;
  _zz_zy_sva_b4 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b4
      ,_zy_sva_b4_t
    ) ;
  _zz_zy_sva_b5 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b5
      ,_zy_sva_b5_t
    ) ;
  _zz_zy_sva_b6 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b6
      ,_zy_sva_b6_t
    ) ;
  _zz_zy_sva_b7 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b7
      ,_zy_sva_b7_t
    ) ;
  _zz_zy_sva_b8 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b8
      ,_zy_sva_b8_t
    ) ;
  _zz_zy_sva_b9 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b9
      ,_zy_sva_b9_t
    ) ;
  _zz_zy_sva_b10 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b10
      ,_zy_sva_b10_t
    ) ;
  _zz_zy_sva_b11 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b11
      ,_zy_sva_b11_t
    ) ;
  _zz_zy_sva_b12 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b12
      ,_zy_sva_b12_t
    ) ;
  _zz_zy_sva_b13 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b13
      ,_zy_sva_b13_t
    ) ;
  _zz_zy_sva_b14 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b14
      ,_zy_sva_b14_t
    ) ;
  _zz_zy_sva_b15 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b15
      ,_zy_sva_b15_t
    ) ;
  _zz_zy_sva_b16 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b16
      ,_zy_sva_b16_t
    ) ;
  _zz_zy_sva_b17 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b17
      ,_zy_sva_b17_t
    ) ;
  _zz_zy_sva_b18 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b18
      ,_zy_sva_b18_t
    ) ;
  _zz_zy_sva_b19 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b19
      ,_zy_sva_b19_t
    ) ;
  _zz_zy_sva_b20 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b20
      ,_zy_sva_b20_t
    ) ;
  _zz_zy_sva_b21 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b21
      ,_zy_sva_b21_t
    ) ;
  _zz_zy_sva_b22 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b22
      ,_zy_sva_b22_t
    ) ;
  _zz_zy_sva_b23 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b23
      ,_zy_sva_b23_t
    ) ;
  _zz_zy_sva_b24 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b24
      ,_zy_sva_b24_t
    ) ;
  _zz_zy_sva_b25 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b25
      ,_zy_sva_b25_t
    ) ;
  _zz_zy_sva_b26 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b26
      ,_zy_sva_b26_t
    ) ;
  _zz_zy_sva_b27 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b27
      ,_zy_sva_b27_t
    ) ;
  _zz_zy_sva_b28 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b28
      ,_zy_sva_b28_t
    ) ;
  _zz_zy_sva_b29 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b29
      ,_zy_sva_b29_t
    ) ;
  _zz_zy_sva_b30 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b30
      ,_zy_sva_b30_t
    ) ;
  _zz_zy_sva_b31 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b31
      ,_zy_sva_b31_t
    ) ;
  _zz_zy_sva_b32 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b32
      ,_zy_sva_b32_t
    ) ;
  _zz_zy_sva_b33 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b33
      ,_zy_sva_b33_t
    ) ;
  _zz_zy_sva_b34 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b34
      ,_zy_sva_b34_t
    ) ;
  _zz_zy_sva_b35 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b35
      ,_zy_sva_b35_t
    ) ;
  _zz_zy_sva_b36 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b36
      ,_zy_sva_b36_t
    ) ;
  _zz_zy_sva_b37 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b37
      ,_zy_sva_b37_t
    ) ;
  _zz_zy_sva_b38 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b38
      ,_zy_sva_b38_t
    ) ;
  _zz_zy_sva_b39 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b39
      ,_zy_sva_b39_t
    ) ;
  _zz_zy_sva_b40 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b40
      ,_zy_sva_b40_t
    ) ;
  _zz_zy_sva_b41 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b41
      ,_zy_sva_b41_t
    ) ;
  _zz_zy_sva_b42 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b42
      ,_zy_sva_b42_t
    ) ;
  _zz_zy_sva_b43 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b43
      ,_zy_sva_b43_t
    ) ;
  _zz_zy_sva_b44 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b44
      ,_zy_sva_b44_t
    ) ;
  _zz_zy_sva_b45 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b45
      ,_zy_sva_b45_t
    ) ;
  _zz_zy_sva_b46 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b46
      ,_zy_sva_b46_t
    ) ;
  _zz_zy_sva_b47 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b47
      ,_zy_sva_b47_t
    ) ;
  _zz_zy_sva_b48 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b48
      ,_zy_sva_b48_t
    ) ;
  _zz_zy_sva_b49 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b49
      ,_zy_sva_b49_t
    ) ;
  _zz_zy_sva_b50 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b50
      ,_zy_sva_b50_t
    ) ;
  _zz_zy_sva_b51 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b51
      ,_zy_sva_b51_t
    ) ;
  _zz_zy_sva_b52 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b52
      ,_zy_sva_b52_t
    ) ;
  _zz_zy_sva_b53 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b53
      ,_zy_sva_b53_t
    ) ;
  _zz_zy_sva_b54 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b54
      ,_zy_sva_b54_t
    ) ;
  _zz_zy_sva_b55 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b55
      ,_zy_sva_b55_t
    ) ;
  _zz_zy_sva_b56 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b56
      ,_zy_sva_b56_t
    ) ;
  _zz_zy_sva_b57 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b57
      ,_zy_sva_b57_t
    ) ;
  _zz_zy_sva_b58 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b58
      ,_zy_sva_b58_t
    ) ;
  _zz_zy_sva_b59 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b59
      ,_zy_sva_b59_t
    ) ;
  _zz_zy_sva_b60 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b60
      ,_zy_sva_b60_t
    ) ;
  _zz_zy_sva_b61 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b61
      ,_zy_sva_b61_t
    ) ;
  _zz_zy_sva_b62 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b62
      ,_zy_sva_b62_t
    ) ;
  _zz_zy_sva_b63 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b63
      ,_zy_sva_b63_t
    ) ;
  _zz_zy_sva_b64 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b64
      ,_zy_sva_b64_t
    ) ;
  _zz_zy_sva_b65 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b65
      ,_zy_sva_b65_t
    ) ;
  _zz_zy_sva_b66 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b66
      ,_zy_sva_b66_t
    ) ;
  _zz_zy_sva_b67 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b67
      ,_zy_sva_b67_t
    ) ;
  _zz_zy_sva_b68 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b68
      ,_zy_sva_b68_t
    ) ;
  _zz_zy_sva_b69 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b69
      ,_zy_sva_b69_t
    ) ;
  _zz_zy_sva_b70 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b70
      ,_zy_sva_b70_t
    ) ;
  _zz_zy_sva_b71 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b71
      ,_zy_sva_b71_t
    ) ;
  _zz_zy_sva_b72 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b72
      ,_zy_sva_b72_t
    ) ;
  _zz_zy_sva_b73 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b73
      ,_zy_sva_b73_t
    ) ;
  _zz_zy_sva_b74 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b74
      ,_zy_sva_b74_t
    ) ;
  _zz_zy_sva_b75 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b75
      ,_zy_sva_b75_t
    ) ;
  _zz_zy_sva_b76 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b76
      ,_zy_sva_b76_t
    ) ;
  _zz_zy_sva_b77 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b77
      ,_zy_sva_b77_t
    ) ;
  _zz_zy_sva_b78 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b78
      ,_zy_sva_b78_t
    ) ;
  _zz_zy_sva_b79 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b79
      ,_zy_sva_b79_t
    ) ;
  _zz_zy_sva_b80 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b80
      ,_zy_sva_b80_t
    ) ;
  _zz_zy_sva_b81 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b81
      ,_zy_sva_b81_t
    ) ;
  _zz_zy_sva_b82 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b82
      ,_zy_sva_b82_t
    ) ;
  _zz_zy_sva_b83 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b83
      ,_zy_sva_b83_t
    ) ;
  _zz_zy_sva_b84 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b84
      ,_zy_sva_b84_t
    ) ;
  _zz_zy_sva_b85 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b85
      ,_zy_sva_b85_t
    ) ;
  _zz_zy_sva_b86 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b86
      ,_zy_sva_b86_t
    ) ;
  _zz_zy_sva_b87 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b87
      ,_zy_sva_b87_t
    ) ;
  _zz_zy_sva_b88 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b88
      ,_zy_sva_b88_t
    ) ;
  _zz_zy_sva_b89 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b89
      ,_zy_sva_b89_t
    ) ;
  _zz_zy_sva_b90 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b90
      ,_zy_sva_b90_t
    ) ;
  _zz_zy_sva_b91 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b91
      ,_zy_sva_b91_t
    ) ;
  _zz_zy_sva_b92 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b92
      ,_zy_sva_b92_t
    ) ;
  _zz_zy_sva_b93 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b93
      ,_zy_sva_b93_t
    ) ;
  _zz_zy_sva_b94 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b94
      ,_zy_sva_b94_t
    ) ;
  _zz_zy_sva_b95 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b95
      ,_zy_sva_b95_t
    ) ;
  _zz_zy_sva_b96 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b96
      ,_zy_sva_b96_t
    ) ;
  _zz_zy_sva_b97 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b97
      ,_zy_sva_b97_t
    ) ;
  _zz_zy_sva_b98 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b98
      ,_zy_sva_b98_t
    ) ;
  _zz_zy_sva_b99 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b99
      ,_zy_sva_b99_t
    ) ;
  _zz_zy_sva_b100 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b100
      ,_zy_sva_b100_t
    ) ;
  _zz_zy_sva_b101 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b101
      ,_zy_sva_b101_t
    ) ;
  _zz_zy_sva_b102 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b102
      ,_zy_sva_b102_t
    ) ;
  _zz_zy_sva_b103 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b103
      ,_zy_sva_b103_t
    ) ;
  _zz_zy_sva_b104 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b104
      ,_zy_sva_b104_t
    ) ;
  _zz_zy_sva_b105 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b105
      ,_zy_sva_b105_t
    ) ;
  _zz_zy_sva_b106 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b106
      ,_zy_sva_b106_t
    ) ;
  _zz_zy_sva_b107 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b107
      ,_zy_sva_b107_t
    ) ;
  _zz_zy_sva_b108 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b108
      ,_zy_sva_b108_t
    ) ;
  _zz_zy_sva_b109 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b109
      ,_zy_sva_b109_t
    ) ;
  _zz_zy_sva_b110 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b110
      ,_zy_sva_b110_t
    ) ;
  _zz_zy_sva_b111 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b111
      ,_zy_sva_b111_t
    ) ;
  _zz_zy_sva_b112 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b112
      ,_zy_sva_b112_t
    ) ;
  _zz_zy_sva_b113 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b113
      ,_zy_sva_b113_t
    ) ;
  _zz_zy_sva_b114 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b114
      ,_zy_sva_b114_t
    ) ;
  _zz_zy_sva_b115 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b115
      ,_zy_sva_b115_t
    ) ;
  _zz_zy_sva_b116 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b116
      ,_zy_sva_b116_t
    ) ;
  _zz_zy_sva_b117 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b117
      ,_zy_sva_b117_t
    ) ;
  _zz_zy_sva_b118 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b118
      ,_zy_sva_b118_t
    ) ;
  _zz_zy_sva_b119 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b119
      ,_zy_sva_b119_t
    ) ;
  _zz_zy_sva_b120 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b120
      ,_zy_sva_b120_t
    ) ;
  _zz_zy_sva_b121 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b121
      ,_zy_sva_b121_t
    ) ;
  _zz_zy_sva_b122 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b122
      ,_zy_sva_b122_t
    ) ;
  _zz_zy_sva_b123 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b123
      ,_zy_sva_b123_t
    ) ;
  _zz_zy_sva_b124 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b124
      ,_zy_sva_b124_t
    ) ;
  _zz_zy_sva_b125 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b125
      ,_zy_sva_b125_t
    ) ;
  _zz_zy_sva_b126 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b126
      ,_zy_sva_b126_t
    ) ;
  _zz_zy_sva_b127 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b127
      ,_zy_sva_b127_t
    ) ;
  _zz_zy_sva_b128 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b128
      ,_zy_sva_b128_t
    ) ;
  _zz_zy_sva_b129 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b129
      ,_zy_sva_b129_t
    ) ;
  _zz_zy_sva_b130 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b130
      ,_zy_sva_b130_t
    ) ;
  _zz_zy_sva_b131 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b131
      ,_zy_sva_b131_t
    ) ;
  _zz_zy_sva_b132 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b132
      ,_zy_sva_b132_t
    ) ;
  _zz_zy_sva_b133 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b133
      ,_zy_sva_b133_t
    ) ;
  _zz_zy_sva_b134 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b134
      ,_zy_sva_b134_t
    ) ;
  _zz_zy_sva_b135 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b135
      ,_zy_sva_b135_t
    ) ;
  _zz_zy_sva_b136 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b136
      ,_zy_sva_b136_t
    ) ;
  _zz_zy_sva_b137 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b137
      ,_zy_sva_b137_t
    ) ;
  _zz_zy_sva_b138 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b138
      ,_zy_sva_b138_t
    ) ;
  _zz_zy_sva_b139 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b139
      ,_zy_sva_b139_t
    ) ;
  _zz_zy_sva_b140 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b140
      ,_zy_sva_b140_t
    ) ;
  _zz_zy_sva_b141 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b141
      ,_zy_sva_b141_t
    ) ;
  _zz_zy_sva_b142 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b142
      ,_zy_sva_b142_t
    ) ;
  _zz_zy_sva_b143 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b143
      ,_zy_sva_b143_t
    ) ;
  _zz_zy_sva_b144 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b144
      ,_zy_sva_b144_t
    ) ;
  _zz_zy_sva_b145 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b145
      ,_zy_sva_b145_t
    ) ;
  _zz_zy_sva_b146 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b146
      ,_zy_sva_b146_t
    ) ;
  _zz_zy_sva_b147 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b147
      ,_zy_sva_b147_t
    ) ;
  _zz_zy_sva_b148 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b148
      ,_zy_sva_b148_t
    ) ;
  _zz_zy_sva_b149 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b149
      ,_zy_sva_b149_t
    ) ;
  _zz_zy_sva_b150 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b150
      ,_zy_sva_b150_t
    ) ;
  _zz_zy_sva_b151 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b151
      ,_zy_sva_b151_t
    ) ;
  _zz_zy_sva_b152 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b152
      ,_zy_sva_b152_t
    ) ;
  _zz_zy_sva_b153 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b153
      ,_zy_sva_b153_t
    ) ;
  _zz_zy_sva_b154 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b154
      ,_zy_sva_b154_t
    ) ;
  _zz_zy_sva_b155 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b155
      ,_zy_sva_b155_t
    ) ;
  _zz_zy_sva_b156 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b156
      ,_zy_sva_b156_t
    ) ;
  _zz_zy_sva_b157 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b157
      ,_zy_sva_b157_t
    ) ;
  _zz_zy_sva_b158 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b158
      ,_zy_sva_b158_t
    ) ;
  _zz_zy_sva_b159 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b159
      ,_zy_sva_b159_t
    ) ;
  _zz_zy_sva_b160 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b160
      ,_zy_sva_b160_t
    ) ;
  _zz_zy_sva_b161 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b161
      ,_zy_sva_b161_t
    ) ;
  _zz_zy_sva_b162 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b162
      ,_zy_sva_b162_t
    ) ;
  _zz_zy_sva_b163 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b163
      ,_zy_sva_b163_t
    ) ;
  _zz_zy_sva_b164 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b164
      ,_zy_sva_b164_t
    ) ;
  _zz_zy_sva_b165 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b165
      ,_zy_sva_b165_t
    ) ;
  _zz_zy_sva_b166 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b166
      ,_zy_sva_b166_t
    ) ;
  _zz_zy_sva_b167 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b167
      ,_zy_sva_b167_t
    ) ;
  _zz_zy_sva_b168 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b168
      ,_zy_sva_b168_t
    ) ;
  _zz_zy_sva_b169 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b169
      ,_zy_sva_b169_t
    ) ;
  _zz_zy_sva_b170 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b170
      ,_zy_sva_b170_t
    ) ;
  _zz_zy_sva_b171 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b171
      ,_zy_sva_b171_t
    ) ;
  _zz_zy_sva_b172 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b172
      ,_zy_sva_b172_t
    ) ;
  _zz_zy_sva_b173 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b173
      ,_zy_sva_b173_t
    ) ;
  _zz_zy_sva_b174 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b174
      ,_zy_sva_b174_t
    ) ;
  _zz_zy_sva_b175 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b175
      ,_zy_sva_b175_t
    ) ;
  _zz_zy_sva_b176 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b176
      ,_zy_sva_b176_t
    ) ;
  _zz_zy_sva_b177 : ixc_sample_logic
    generic map(WIDTH => 1,RD_TYPE => 3)
    port map (
       _zy_sva_b177
      ,_zy_sva_b177_t
    ) ;
  parser_fifo : cr_kme_fifo_xcm58
    port map (
       fifo_in_stall => fifo_in_stall
      ,fifo_out => DUMMY4
      ,fifo_out_valid => parser_kimreader_valid
      ,fifo_overflow => _zy_simnet_dio_3
      ,fifo_underflow => _zy_simnet_dio_4
      ,clk => clk
      ,rst_n => rst_n
      ,fifo_in => DUMMY5
      ,fifo_in_valid => DUMMY6
      ,fifo_out_ack => kimreader_parser_ack
      ,fifo_in_stall_override => _zy_simnet_cio_7
    ) ;

  process --:o2835
  (clk,_zy_sva_key_type0_line4_1_reset_or)
    variable DUMMY8 : std_logic ;
  begin
    if (_zy_sva_key_type0_line4_1_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY8 := _zy_sva_b0 ;
      _zy_sva_key_type0_line4_1_ccheck <= "1" ;
      if (DUMMY8 = '1') then
        _zy_sva_key_type0_line4_1_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o2852
  (clk,_zy_sva_key_type0_line5a_2_reset_or)
    variable DUMMY9 : std_logic ;
  begin
    if (_zy_sva_key_type0_line5a_2_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY9 := _zy_sva_b1 ;
      _zy_sva_key_type0_line5a_2_ccheck <= "1" ;
      if (DUMMY9 = '1') then
        _zy_sva_key_type0_line5a_2_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o2869
  (clk,_zy_sva_key_type0_line5b_3_reset_or)
    variable DUMMY10 : std_logic ;
  begin
    if (_zy_sva_key_type0_line5b_3_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY10 := _zy_sva_b2 ;
      _zy_sva_key_type0_line5b_3_ccheck <= "1" ;
      if (DUMMY10 = '1') then
        _zy_sva_key_type0_line5b_3_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o2886
  (clk,_zy_sva_key_type1_line7a_4_reset_or)
    variable DUMMY11 : std_logic ;
  begin
    if (_zy_sva_key_type1_line7a_4_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY11 := _zy_sva_b3 ;
      _zy_sva_key_type1_line7a_4_ccheck <= "1" ;
      if (DUMMY11 = '1') then
        _zy_sva_key_type1_line7a_4_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o2903
  (clk,_zy_sva_key_type1_line7b_5_reset_or)
    variable DUMMY12 : std_logic ;
  begin
    if (_zy_sva_key_type1_line7b_5_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY12 := _zy_sva_b4 ;
      _zy_sva_key_type1_line7b_5_ccheck <= "1" ;
      if (DUMMY12 = '1') then
        _zy_sva_key_type1_line7b_5_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o2920
  (clk,_zy_sva_key_type1_line8a_6_reset_or)
    variable DUMMY13 : std_logic ;
  begin
    if (_zy_sva_key_type1_line8a_6_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY13 := _zy_sva_b5 ;
      _zy_sva_key_type1_line8a_6_ccheck <= "1" ;
      if (DUMMY13 = '1') then
        _zy_sva_key_type1_line8a_6_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o2937
  (clk,_zy_sva_key_type1_line8b_7_reset_or)
    variable DUMMY14 : std_logic ;
  begin
    if (_zy_sva_key_type1_line8b_7_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY14 := _zy_sva_b6 ;
      _zy_sva_key_type1_line8b_7_ccheck <= "1" ;
      if (DUMMY14 = '1') then
        _zy_sva_key_type1_line8b_7_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o2954
  (clk,_zy_sva_key_type1_line9_8_reset_or)
    variable DUMMY15 : std_logic ;
  begin
    if (_zy_sva_key_type1_line9_8_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY15 := _zy_sva_b7 ;
      _zy_sva_key_type1_line9_8_ccheck <= "1" ;
      if (DUMMY15 = '1') then
        _zy_sva_key_type1_line9_8_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o2971
  (clk,_zy_sva_key_type1_line10_9_reset_or)
    variable DUMMY16 : std_logic ;
  begin
    if (_zy_sva_key_type1_line10_9_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY16 := _zy_sva_b8 ;
      _zy_sva_key_type1_line10_9_ccheck <= "1" ;
      if (DUMMY16 = '1') then
        _zy_sva_key_type1_line10_9_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o2988
  (clk,_zy_sva_key_type1_line11a_10_reset_or)
    variable DUMMY17 : std_logic ;
  begin
    if (_zy_sva_key_type1_line11a_10_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY17 := _zy_sva_b9 ;
      _zy_sva_key_type1_line11a_10_ccheck <= "1" ;
      if (DUMMY17 = '1') then
        _zy_sva_key_type1_line11a_10_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3005
  (clk,_zy_sva_key_type1_line11b_11_reset_or)
    variable DUMMY18 : std_logic ;
  begin
    if (_zy_sva_key_type1_line11b_11_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY18 := _zy_sva_b10 ;
      _zy_sva_key_type1_line11b_11_ccheck <= "1" ;
      if (DUMMY18 = '1') then
        _zy_sva_key_type1_line11b_11_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3022
  (clk,_zy_sva_key_type1_line11c_12_reset_or)
    variable DUMMY19 : std_logic ;
  begin
    if (_zy_sva_key_type1_line11c_12_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY19 := _zy_sva_b11 ;
      _zy_sva_key_type1_line11c_12_ccheck <= "1" ;
      if (DUMMY19 = '1') then
        _zy_sva_key_type1_line11c_12_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3039
  (clk,_zy_sva_key_type1_line11d_13_reset_or)
    variable DUMMY20 : std_logic ;
  begin
    if (_zy_sva_key_type1_line11d_13_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY20 := _zy_sva_b12 ;
      _zy_sva_key_type1_line11d_13_ccheck <= "1" ;
      if (DUMMY20 = '1') then
        _zy_sva_key_type1_line11d_13_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3056
  (clk,_zy_sva_key_type1_line12a_14_reset_or)
    variable DUMMY21 : std_logic ;
  begin
    if (_zy_sva_key_type1_line12a_14_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY21 := _zy_sva_b13 ;
      _zy_sva_key_type1_line12a_14_ccheck <= "1" ;
      if (DUMMY21 = '1') then
        _zy_sva_key_type1_line12a_14_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3073
  (clk,_zy_sva_key_type1_line12b_15_reset_or)
    variable DUMMY22 : std_logic ;
  begin
    if (_zy_sva_key_type1_line12b_15_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY22 := _zy_sva_b14 ;
      _zy_sva_key_type1_line12b_15_ccheck <= "1" ;
      if (DUMMY22 = '1') then
        _zy_sva_key_type1_line12b_15_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3090
  (clk,_zy_sva_key_type9_line14_16_reset_or)
    variable DUMMY23 : std_logic ;
  begin
    if (_zy_sva_key_type9_line14_16_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY23 := _zy_sva_b15 ;
      _zy_sva_key_type9_line14_16_ccheck <= "1" ;
      if (DUMMY23 = '1') then
        _zy_sva_key_type9_line14_16_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3107
  (clk,_zy_sva_key_type9_line15_17_reset_or)
    variable DUMMY24 : std_logic ;
  begin
    if (_zy_sva_key_type9_line15_17_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY24 := _zy_sva_b16 ;
      _zy_sva_key_type9_line15_17_ccheck <= "1" ;
      if (DUMMY24 = '1') then
        _zy_sva_key_type9_line15_17_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3124
  (clk,_zy_sva_key_type9_line16a_18_reset_or)
    variable DUMMY25 : std_logic ;
  begin
    if (_zy_sva_key_type9_line16a_18_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY25 := _zy_sva_b17 ;
      _zy_sva_key_type9_line16a_18_ccheck <= "1" ;
      if (DUMMY25 = '1') then
        _zy_sva_key_type9_line16a_18_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3141
  (clk,_zy_sva_key_type9_line16b_19_reset_or)
    variable DUMMY26 : std_logic ;
  begin
    if (_zy_sva_key_type9_line16b_19_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY26 := _zy_sva_b18 ;
      _zy_sva_key_type9_line16b_19_ccheck <= "1" ;
      if (DUMMY26 = '1') then
        _zy_sva_key_type9_line16b_19_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3158
  (clk,_zy_sva_key_type9_line17a_20_reset_or)
    variable DUMMY27 : std_logic ;
  begin
    if (_zy_sva_key_type9_line17a_20_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY27 := _zy_sva_b19 ;
      _zy_sva_key_type9_line17a_20_ccheck <= "1" ;
      if (DUMMY27 = '1') then
        _zy_sva_key_type9_line17a_20_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3175
  (clk,_zy_sva_key_type9_line17b_21_reset_or)
    variable DUMMY28 : std_logic ;
  begin
    if (_zy_sva_key_type9_line17b_21_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY28 := _zy_sva_b20 ;
      _zy_sva_key_type9_line17b_21_ccheck <= "1" ;
      if (DUMMY28 = '1') then
        _zy_sva_key_type9_line17b_21_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3192
  (clk,_zy_sva_key_type9_line18a_22_reset_or)
    variable DUMMY29 : std_logic ;
  begin
    if (_zy_sva_key_type9_line18a_22_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY29 := _zy_sva_b21 ;
      _zy_sva_key_type9_line18a_22_ccheck <= "1" ;
      if (DUMMY29 = '1') then
        _zy_sva_key_type9_line18a_22_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3209
  (clk,_zy_sva_key_type9_line18b_23_reset_or)
    variable DUMMY30 : std_logic ;
  begin
    if (_zy_sva_key_type9_line18b_23_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY30 := _zy_sva_b22 ;
      _zy_sva_key_type9_line18b_23_ccheck <= "1" ;
      if (DUMMY30 = '1') then
        _zy_sva_key_type9_line18b_23_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3226
  (clk,_zy_sva_key_type9_line19a_24_reset_or)
    variable DUMMY31 : std_logic ;
  begin
    if (_zy_sva_key_type9_line19a_24_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY31 := _zy_sva_b23 ;
      _zy_sva_key_type9_line19a_24_ccheck <= "1" ;
      if (DUMMY31 = '1') then
        _zy_sva_key_type9_line19a_24_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3243
  (clk,_zy_sva_key_type9_line19b_25_reset_or)
    variable DUMMY32 : std_logic ;
  begin
    if (_zy_sva_key_type9_line19b_25_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY32 := _zy_sva_b24 ;
      _zy_sva_key_type9_line19b_25_ccheck <= "1" ;
      if (DUMMY32 = '1') then
        _zy_sva_key_type9_line19b_25_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3260
  (clk,_zy_sva_key_type9_line19c_26_reset_or)
    variable DUMMY33 : std_logic ;
  begin
    if (_zy_sva_key_type9_line19c_26_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY33 := _zy_sva_b25 ;
      _zy_sva_key_type9_line19c_26_ccheck <= "1" ;
      if (DUMMY33 = '1') then
        _zy_sva_key_type9_line19c_26_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3277
  (clk,_zy_sva_key_type9_line19d_27_reset_or)
    variable DUMMY34 : std_logic ;
  begin
    if (_zy_sva_key_type9_line19d_27_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY34 := _zy_sva_b26 ;
      _zy_sva_key_type9_line19d_27_ccheck <= "1" ;
      if (DUMMY34 = '1') then
        _zy_sva_key_type9_line19d_27_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3294
  (clk,_zy_sva_guid_miss_aux_cmd_0_28_reset_or)
    variable DUMMY35 : std_logic ;
  begin
    if (_zy_sva_guid_miss_aux_cmd_0_28_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY35 := _zy_sva_b27 ;
      _zy_sva_guid_miss_aux_cmd_0_28_ccheck <= "1" ;
      if (DUMMY35 = '1') then
        _zy_sva_guid_miss_aux_cmd_0_28_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3311
  (clk,_zy_sva_guid_miss_aux_cmd_1_29_reset_or)
    variable DUMMY36 : std_logic ;
  begin
    if (_zy_sva_guid_miss_aux_cmd_1_29_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY36 := _zy_sva_b28 ;
      _zy_sva_guid_miss_aux_cmd_1_29_ccheck <= "1" ;
      if (DUMMY36 = '1') then
        _zy_sva_guid_miss_aux_cmd_1_29_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3328
  (clk,_zy_sva_guid_miss_aux_cmd_2_30_reset_or)
    variable DUMMY37 : std_logic ;
  begin
    if (_zy_sva_guid_miss_aux_cmd_2_30_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY37 := _zy_sva_b29 ;
      _zy_sva_guid_miss_aux_cmd_2_30_ccheck <= "1" ;
      if (DUMMY37 = '1') then
        _zy_sva_guid_miss_aux_cmd_2_30_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3345
  (clk,_zy_sva_guid_miss_aux_cmd_3_31_reset_or)
    variable DUMMY38 : std_logic ;
  begin
    if (_zy_sva_guid_miss_aux_cmd_3_31_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY38 := _zy_sva_b30 ;
      _zy_sva_guid_miss_aux_cmd_3_31_ccheck <= "1" ;
      if (DUMMY38 = '1') then
        _zy_sva_guid_miss_aux_cmd_3_31_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3362
  (clk,_zy_sva_guid_miss_aux_cmd_iv_0_32_reset_or)
    variable DUMMY39 : std_logic ;
  begin
    if (_zy_sva_guid_miss_aux_cmd_iv_0_32_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY39 := _zy_sva_b31 ;
      _zy_sva_guid_miss_aux_cmd_iv_0_32_ccheck <= "1" ;
      if (DUMMY39 = '1') then
        _zy_sva_guid_miss_aux_cmd_iv_0_32_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3379
  (clk,_zy_sva_guid_miss_aux_cmd_iv_1_33_reset_or)
    variable DUMMY40 : std_logic ;
  begin
    if (_zy_sva_guid_miss_aux_cmd_iv_1_33_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY40 := _zy_sva_b32 ;
      _zy_sva_guid_miss_aux_cmd_iv_1_33_ccheck <= "1" ;
      if (DUMMY40 = '1') then
        _zy_sva_guid_miss_aux_cmd_iv_1_33_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3396
  (clk,_zy_sva_guid_miss_aux_cmd_iv_2_34_reset_or)
    variable DUMMY41 : std_logic ;
  begin
    if (_zy_sva_guid_miss_aux_cmd_iv_2_34_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY41 := _zy_sva_b33 ;
      _zy_sva_guid_miss_aux_cmd_iv_2_34_ccheck <= "1" ;
      if (DUMMY41 = '1') then
        _zy_sva_guid_miss_aux_cmd_iv_2_34_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3413
  (clk,_zy_sva_guid_miss_aux_cmd_iv_3_35_reset_or)
    variable DUMMY42 : std_logic ;
  begin
    if (_zy_sva_guid_miss_aux_cmd_iv_3_35_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY42 := _zy_sva_b34 ;
      _zy_sva_guid_miss_aux_cmd_iv_3_35_ccheck <= "1" ;
      if (DUMMY42 = '1') then
        _zy_sva_guid_miss_aux_cmd_iv_3_35_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3430
  (clk,_zy_sva_iv_miss_aux_cmd_0_36_reset_or)
    variable DUMMY43 : std_logic ;
  begin
    if (_zy_sva_iv_miss_aux_cmd_0_36_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY43 := _zy_sva_b35 ;
      _zy_sva_iv_miss_aux_cmd_0_36_ccheck <= "1" ;
      if (DUMMY43 = '1') then
        _zy_sva_iv_miss_aux_cmd_0_36_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3447
  (clk,_zy_sva_iv_miss_aux_cmd_1_37_reset_or)
    variable DUMMY44 : std_logic ;
  begin
    if (_zy_sva_iv_miss_aux_cmd_1_37_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY44 := _zy_sva_b36 ;
      _zy_sva_iv_miss_aux_cmd_1_37_ccheck <= "1" ;
      if (DUMMY44 = '1') then
        _zy_sva_iv_miss_aux_cmd_1_37_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3464
  (clk,_zy_sva_iv_miss_aux_cmd_guid_38_reset_or)
    variable DUMMY45 : std_logic ;
  begin
    if (_zy_sva_iv_miss_aux_cmd_guid_38_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY45 := _zy_sva_b37 ;
      _zy_sva_iv_miss_aux_cmd_guid_38_ccheck <= "1" ;
      if (DUMMY45 = '1') then
        _zy_sva_iv_miss_aux_cmd_guid_38_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3481
  (clk,_zy_sva_brcm_aux_cmd_39_reset_or)
    variable DUMMY46 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_39_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY46 := _zy_sva_b38 ;
      _zy_sva_brcm_aux_cmd_39_ccheck <= "1" ;
      if (DUMMY46 = '1') then
        _zy_sva_brcm_aux_cmd_39_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3498
  (clk,_zy_sva_brcm_aux_cmd_iv_40_reset_or)
    variable DUMMY47 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_iv_40_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY47 := _zy_sva_b39 ;
      _zy_sva_brcm_aux_cmd_iv_40_ccheck <= "1" ;
      if (DUMMY47 = '1') then
        _zy_sva_brcm_aux_cmd_iv_40_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3515
  (clk,_zy_sva_brcm_aux_cmd_guid_41_reset_or)
    variable DUMMY48 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_guid_41_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY48 := _zy_sva_b40 ;
      _zy_sva_brcm_aux_cmd_guid_41_ccheck <= "1" ;
      if (DUMMY48 = '1') then
        _zy_sva_brcm_aux_cmd_guid_41_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3532
  (clk,_zy_sva_brcm_aux_cmd_guid_iv_42_reset_or)
    variable DUMMY49 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_guid_iv_42_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY49 := _zy_sva_b41 ;
      _zy_sva_brcm_aux_cmd_guid_iv_42_ccheck <= "1" ;
      if (DUMMY49 = '1') then
        _zy_sva_brcm_aux_cmd_guid_iv_42_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3549
  (clk,_zy_sva_brcm_key_type_43_reset_or)
    variable DUMMY50 : std_logic ;
  begin
    if (_zy_sva_brcm_key_type_43_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY50 := _zy_sva_b42 ;
      _zy_sva_brcm_key_type_43_ccheck <= "1" ;
      if (DUMMY50 = '1') then
        _zy_sva_brcm_key_type_43_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3566
  (clk,_zy_sva_brcm_aux_cmd_44_reset_or)
    variable DUMMY51 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_44_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY51 := _zy_sva_b43 ;
      _zy_sva_brcm_aux_cmd_44_ccheck <= "1" ;
      if (DUMMY51 = '1') then
        _zy_sva_brcm_aux_cmd_44_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3583
  (clk,_zy_sva_brcm_aux_cmd_iv_45_reset_or)
    variable DUMMY52 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_iv_45_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY52 := _zy_sva_b44 ;
      _zy_sva_brcm_aux_cmd_iv_45_ccheck <= "1" ;
      if (DUMMY52 = '1') then
        _zy_sva_brcm_aux_cmd_iv_45_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3600
  (clk,_zy_sva_brcm_aux_cmd_guid_46_reset_or)
    variable DUMMY53 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_guid_46_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY53 := _zy_sva_b45 ;
      _zy_sva_brcm_aux_cmd_guid_46_ccheck <= "1" ;
      if (DUMMY53 = '1') then
        _zy_sva_brcm_aux_cmd_guid_46_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3617
  (clk,_zy_sva_brcm_aux_cmd_guid_iv_47_reset_or)
    variable DUMMY54 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_guid_iv_47_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY54 := _zy_sva_b46 ;
      _zy_sva_brcm_aux_cmd_guid_iv_47_ccheck <= "1" ;
      if (DUMMY54 = '1') then
        _zy_sva_brcm_aux_cmd_guid_iv_47_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3634
  (clk,_zy_sva_brcm_key_type_48_reset_or)
    variable DUMMY55 : std_logic ;
  begin
    if (_zy_sva_brcm_key_type_48_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY55 := _zy_sva_b47 ;
      _zy_sva_brcm_key_type_48_ccheck <= "1" ;
      if (DUMMY55 = '1') then
        _zy_sva_brcm_key_type_48_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3651
  (clk,_zy_sva_brcm_aux_cmd_49_reset_or)
    variable DUMMY56 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_49_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY56 := _zy_sva_b48 ;
      _zy_sva_brcm_aux_cmd_49_ccheck <= "1" ;
      if (DUMMY56 = '1') then
        _zy_sva_brcm_aux_cmd_49_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3668
  (clk,_zy_sva_brcm_aux_cmd_iv_50_reset_or)
    variable DUMMY57 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_iv_50_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY57 := _zy_sva_b49 ;
      _zy_sva_brcm_aux_cmd_iv_50_ccheck <= "1" ;
      if (DUMMY57 = '1') then
        _zy_sva_brcm_aux_cmd_iv_50_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3685
  (clk,_zy_sva_brcm_aux_cmd_guid_51_reset_or)
    variable DUMMY58 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_guid_51_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY58 := _zy_sva_b50 ;
      _zy_sva_brcm_aux_cmd_guid_51_ccheck <= "1" ;
      if (DUMMY58 = '1') then
        _zy_sva_brcm_aux_cmd_guid_51_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3702
  (clk,_zy_sva_brcm_aux_cmd_guid_iv_52_reset_or)
    variable DUMMY59 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_guid_iv_52_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY59 := _zy_sva_b51 ;
      _zy_sva_brcm_aux_cmd_guid_iv_52_ccheck <= "1" ;
      if (DUMMY59 = '1') then
        _zy_sva_brcm_aux_cmd_guid_iv_52_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3719
  (clk,_zy_sva_brcm_key_type_53_reset_or)
    variable DUMMY60 : std_logic ;
  begin
    if (_zy_sva_brcm_key_type_53_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY60 := _zy_sva_b52 ;
      _zy_sva_brcm_key_type_53_ccheck <= "1" ;
      if (DUMMY60 = '1') then
        _zy_sva_brcm_key_type_53_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3736
  (clk,_zy_sva_brcm_aux_cmd_54_reset_or)
    variable DUMMY61 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_54_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY61 := _zy_sva_b53 ;
      _zy_sva_brcm_aux_cmd_54_ccheck <= "1" ;
      if (DUMMY61 = '1') then
        _zy_sva_brcm_aux_cmd_54_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3753
  (clk,_zy_sva_brcm_aux_cmd_iv_55_reset_or)
    variable DUMMY62 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_iv_55_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY62 := _zy_sva_b54 ;
      _zy_sva_brcm_aux_cmd_iv_55_ccheck <= "1" ;
      if (DUMMY62 = '1') then
        _zy_sva_brcm_aux_cmd_iv_55_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3770
  (clk,_zy_sva_brcm_aux_cmd_guid_56_reset_or)
    variable DUMMY63 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_guid_56_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY63 := _zy_sva_b55 ;
      _zy_sva_brcm_aux_cmd_guid_56_ccheck <= "1" ;
      if (DUMMY63 = '1') then
        _zy_sva_brcm_aux_cmd_guid_56_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3787
  (clk,_zy_sva_brcm_aux_cmd_guid_iv_57_reset_or)
    variable DUMMY64 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_guid_iv_57_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY64 := _zy_sva_b56 ;
      _zy_sva_brcm_aux_cmd_guid_iv_57_ccheck <= "1" ;
      if (DUMMY64 = '1') then
        _zy_sva_brcm_aux_cmd_guid_iv_57_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3804
  (clk,_zy_sva_brcm_key_type_58_reset_or)
    variable DUMMY65 : std_logic ;
  begin
    if (_zy_sva_brcm_key_type_58_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY65 := _zy_sva_b57 ;
      _zy_sva_brcm_key_type_58_ccheck <= "1" ;
      if (DUMMY65 = '1') then
        _zy_sva_brcm_key_type_58_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3821
  (clk,_zy_sva_brcm_aux_cmd_59_reset_or)
    variable DUMMY66 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_59_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY66 := _zy_sva_b58 ;
      _zy_sva_brcm_aux_cmd_59_ccheck <= "1" ;
      if (DUMMY66 = '1') then
        _zy_sva_brcm_aux_cmd_59_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3838
  (clk,_zy_sva_brcm_aux_cmd_iv_60_reset_or)
    variable DUMMY67 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_iv_60_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY67 := _zy_sva_b59 ;
      _zy_sva_brcm_aux_cmd_iv_60_ccheck <= "1" ;
      if (DUMMY67 = '1') then
        _zy_sva_brcm_aux_cmd_iv_60_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3855
  (clk,_zy_sva_brcm_aux_cmd_guid_61_reset_or)
    variable DUMMY68 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_guid_61_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY68 := _zy_sva_b60 ;
      _zy_sva_brcm_aux_cmd_guid_61_ccheck <= "1" ;
      if (DUMMY68 = '1') then
        _zy_sva_brcm_aux_cmd_guid_61_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3872
  (clk,_zy_sva_brcm_aux_cmd_guid_iv_62_reset_or)
    variable DUMMY69 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_guid_iv_62_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY69 := _zy_sva_b61 ;
      _zy_sva_brcm_aux_cmd_guid_iv_62_ccheck <= "1" ;
      if (DUMMY69 = '1') then
        _zy_sva_brcm_aux_cmd_guid_iv_62_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3889
  (clk,_zy_sva_brcm_key_type_63_reset_or)
    variable DUMMY70 : std_logic ;
  begin
    if (_zy_sva_brcm_key_type_63_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY70 := _zy_sva_b62 ;
      _zy_sva_brcm_key_type_63_ccheck <= "1" ;
      if (DUMMY70 = '1') then
        _zy_sva_brcm_key_type_63_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3906
  (clk,_zy_sva_brcm_aux_cmd_64_reset_or)
    variable DUMMY71 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_64_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY71 := _zy_sva_b63 ;
      _zy_sva_brcm_aux_cmd_64_ccheck <= "1" ;
      if (DUMMY71 = '1') then
        _zy_sva_brcm_aux_cmd_64_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3923
  (clk,_zy_sva_brcm_aux_cmd_iv_65_reset_or)
    variable DUMMY72 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_iv_65_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY72 := _zy_sva_b64 ;
      _zy_sva_brcm_aux_cmd_iv_65_ccheck <= "1" ;
      if (DUMMY72 = '1') then
        _zy_sva_brcm_aux_cmd_iv_65_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3940
  (clk,_zy_sva_brcm_aux_cmd_guid_66_reset_or)
    variable DUMMY73 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_guid_66_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY73 := _zy_sva_b65 ;
      _zy_sva_brcm_aux_cmd_guid_66_ccheck <= "1" ;
      if (DUMMY73 = '1') then
        _zy_sva_brcm_aux_cmd_guid_66_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3957
  (clk,_zy_sva_brcm_aux_cmd_guid_iv_67_reset_or)
    variable DUMMY74 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_guid_iv_67_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY74 := _zy_sva_b66 ;
      _zy_sva_brcm_aux_cmd_guid_iv_67_ccheck <= "1" ;
      if (DUMMY74 = '1') then
        _zy_sva_brcm_aux_cmd_guid_iv_67_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3974
  (clk,_zy_sva_brcm_key_type_68_reset_or)
    variable DUMMY75 : std_logic ;
  begin
    if (_zy_sva_brcm_key_type_68_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY75 := _zy_sva_b67 ;
      _zy_sva_brcm_key_type_68_ccheck <= "1" ;
      if (DUMMY75 = '1') then
        _zy_sva_brcm_key_type_68_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o3991
  (clk,_zy_sva_brcm_aux_cmd_69_reset_or)
    variable DUMMY76 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_69_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY76 := _zy_sva_b68 ;
      _zy_sva_brcm_aux_cmd_69_ccheck <= "1" ;
      if (DUMMY76 = '1') then
        _zy_sva_brcm_aux_cmd_69_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4008
  (clk,_zy_sva_brcm_aux_cmd_iv_70_reset_or)
    variable DUMMY77 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_iv_70_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY77 := _zy_sva_b69 ;
      _zy_sva_brcm_aux_cmd_iv_70_ccheck <= "1" ;
      if (DUMMY77 = '1') then
        _zy_sva_brcm_aux_cmd_iv_70_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4025
  (clk,_zy_sva_brcm_aux_cmd_guid_71_reset_or)
    variable DUMMY78 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_guid_71_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY78 := _zy_sva_b70 ;
      _zy_sva_brcm_aux_cmd_guid_71_ccheck <= "1" ;
      if (DUMMY78 = '1') then
        _zy_sva_brcm_aux_cmd_guid_71_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4042
  (clk,_zy_sva_brcm_aux_cmd_guid_iv_72_reset_or)
    variable DUMMY79 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_guid_iv_72_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY79 := _zy_sva_b71 ;
      _zy_sva_brcm_aux_cmd_guid_iv_72_ccheck <= "1" ;
      if (DUMMY79 = '1') then
        _zy_sva_brcm_aux_cmd_guid_iv_72_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4059
  (clk,_zy_sva_brcm_key_type_73_reset_or)
    variable DUMMY80 : std_logic ;
  begin
    if (_zy_sva_brcm_key_type_73_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY80 := _zy_sva_b72 ;
      _zy_sva_brcm_key_type_73_ccheck <= "1" ;
      if (DUMMY80 = '1') then
        _zy_sva_brcm_key_type_73_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4076
  (clk,_zy_sva_brcm_aux_cmd_74_reset_or)
    variable DUMMY81 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_74_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY81 := _zy_sva_b73 ;
      _zy_sva_brcm_aux_cmd_74_ccheck <= "1" ;
      if (DUMMY81 = '1') then
        _zy_sva_brcm_aux_cmd_74_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4093
  (clk,_zy_sva_brcm_aux_cmd_iv_75_reset_or)
    variable DUMMY82 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_iv_75_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY82 := _zy_sva_b74 ;
      _zy_sva_brcm_aux_cmd_iv_75_ccheck <= "1" ;
      if (DUMMY82 = '1') then
        _zy_sva_brcm_aux_cmd_iv_75_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4110
  (clk,_zy_sva_brcm_aux_cmd_guid_76_reset_or)
    variable DUMMY83 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_guid_76_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY83 := _zy_sva_b75 ;
      _zy_sva_brcm_aux_cmd_guid_76_ccheck <= "1" ;
      if (DUMMY83 = '1') then
        _zy_sva_brcm_aux_cmd_guid_76_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4127
  (clk,_zy_sva_brcm_aux_cmd_guid_iv_77_reset_or)
    variable DUMMY84 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_guid_iv_77_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY84 := _zy_sva_b76 ;
      _zy_sva_brcm_aux_cmd_guid_iv_77_ccheck <= "1" ;
      if (DUMMY84 = '1') then
        _zy_sva_brcm_aux_cmd_guid_iv_77_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4144
  (clk,_zy_sva_brcm_key_type_78_reset_or)
    variable DUMMY85 : std_logic ;
  begin
    if (_zy_sva_brcm_key_type_78_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY85 := _zy_sva_b77 ;
      _zy_sva_brcm_key_type_78_ccheck <= "1" ;
      if (DUMMY85 = '1') then
        _zy_sva_brcm_key_type_78_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4161
  (clk,_zy_sva_brcm_aux_cmd_79_reset_or)
    variable DUMMY86 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_79_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY86 := _zy_sva_b78 ;
      _zy_sva_brcm_aux_cmd_79_ccheck <= "1" ;
      if (DUMMY86 = '1') then
        _zy_sva_brcm_aux_cmd_79_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4178
  (clk,_zy_sva_brcm_aux_cmd_iv_80_reset_or)
    variable DUMMY87 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_iv_80_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY87 := _zy_sva_b79 ;
      _zy_sva_brcm_aux_cmd_iv_80_ccheck <= "1" ;
      if (DUMMY87 = '1') then
        _zy_sva_brcm_aux_cmd_iv_80_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4195
  (clk,_zy_sva_brcm_aux_cmd_guid_81_reset_or)
    variable DUMMY88 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_guid_81_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY88 := _zy_sva_b80 ;
      _zy_sva_brcm_aux_cmd_guid_81_ccheck <= "1" ;
      if (DUMMY88 = '1') then
        _zy_sva_brcm_aux_cmd_guid_81_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4212
  (clk,_zy_sva_brcm_aux_cmd_guid_iv_82_reset_or)
    variable DUMMY89 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_guid_iv_82_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY89 := _zy_sva_b81 ;
      _zy_sva_brcm_aux_cmd_guid_iv_82_ccheck <= "1" ;
      if (DUMMY89 = '1') then
        _zy_sva_brcm_aux_cmd_guid_iv_82_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4229
  (clk,_zy_sva_brcm_key_type_83_reset_or)
    variable DUMMY90 : std_logic ;
  begin
    if (_zy_sva_brcm_key_type_83_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY90 := _zy_sva_b82 ;
      _zy_sva_brcm_key_type_83_ccheck <= "1" ;
      if (DUMMY90 = '1') then
        _zy_sva_brcm_key_type_83_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4246
  (clk,_zy_sva_brcm_aux_cmd_84_reset_or)
    variable DUMMY91 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_84_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY91 := _zy_sva_b83 ;
      _zy_sva_brcm_aux_cmd_84_ccheck <= "1" ;
      if (DUMMY91 = '1') then
        _zy_sva_brcm_aux_cmd_84_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4263
  (clk,_zy_sva_brcm_aux_cmd_iv_85_reset_or)
    variable DUMMY92 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_iv_85_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY92 := _zy_sva_b84 ;
      _zy_sva_brcm_aux_cmd_iv_85_ccheck <= "1" ;
      if (DUMMY92 = '1') then
        _zy_sva_brcm_aux_cmd_iv_85_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4280
  (clk,_zy_sva_brcm_aux_cmd_guid_86_reset_or)
    variable DUMMY93 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_guid_86_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY93 := _zy_sva_b85 ;
      _zy_sva_brcm_aux_cmd_guid_86_ccheck <= "1" ;
      if (DUMMY93 = '1') then
        _zy_sva_brcm_aux_cmd_guid_86_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4297
  (clk,_zy_sva_brcm_aux_cmd_guid_iv_87_reset_or)
    variable DUMMY94 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_guid_iv_87_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY94 := _zy_sva_b86 ;
      _zy_sva_brcm_aux_cmd_guid_iv_87_ccheck <= "1" ;
      if (DUMMY94 = '1') then
        _zy_sva_brcm_aux_cmd_guid_iv_87_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4314
  (clk,_zy_sva_brcm_key_type_88_reset_or)
    variable DUMMY95 : std_logic ;
  begin
    if (_zy_sva_brcm_key_type_88_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY95 := _zy_sva_b87 ;
      _zy_sva_brcm_key_type_88_ccheck <= "1" ;
      if (DUMMY95 = '1') then
        _zy_sva_brcm_key_type_88_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4331
  (clk,_zy_sva_brcm_aux_cmd_89_reset_or)
    variable DUMMY96 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_89_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY96 := _zy_sva_b88 ;
      _zy_sva_brcm_aux_cmd_89_ccheck <= "1" ;
      if (DUMMY96 = '1') then
        _zy_sva_brcm_aux_cmd_89_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4348
  (clk,_zy_sva_brcm_aux_cmd_iv_90_reset_or)
    variable DUMMY97 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_iv_90_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY97 := _zy_sva_b89 ;
      _zy_sva_brcm_aux_cmd_iv_90_ccheck <= "1" ;
      if (DUMMY97 = '1') then
        _zy_sva_brcm_aux_cmd_iv_90_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4365
  (clk,_zy_sva_brcm_aux_cmd_guid_91_reset_or)
    variable DUMMY98 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_guid_91_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY98 := _zy_sva_b90 ;
      _zy_sva_brcm_aux_cmd_guid_91_ccheck <= "1" ;
      if (DUMMY98 = '1') then
        _zy_sva_brcm_aux_cmd_guid_91_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4382
  (clk,_zy_sva_brcm_aux_cmd_guid_iv_92_reset_or)
    variable DUMMY99 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_guid_iv_92_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY99 := _zy_sva_b91 ;
      _zy_sva_brcm_aux_cmd_guid_iv_92_ccheck <= "1" ;
      if (DUMMY99 = '1') then
        _zy_sva_brcm_aux_cmd_guid_iv_92_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4399
  (clk,_zy_sva_brcm_key_type_93_reset_or)
    variable DUMMY100 : std_logic ;
  begin
    if (_zy_sva_brcm_key_type_93_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY100 := _zy_sva_b92 ;
      _zy_sva_brcm_key_type_93_ccheck <= "1" ;
      if (DUMMY100 = '1') then
        _zy_sva_brcm_key_type_93_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4416
  (clk,_zy_sva_brcm_aux_cmd_94_reset_or)
    variable DUMMY101 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_94_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY101 := _zy_sva_b93 ;
      _zy_sva_brcm_aux_cmd_94_ccheck <= "1" ;
      if (DUMMY101 = '1') then
        _zy_sva_brcm_aux_cmd_94_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4433
  (clk,_zy_sva_brcm_aux_cmd_iv_95_reset_or)
    variable DUMMY102 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_iv_95_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY102 := _zy_sva_b94 ;
      _zy_sva_brcm_aux_cmd_iv_95_ccheck <= "1" ;
      if (DUMMY102 = '1') then
        _zy_sva_brcm_aux_cmd_iv_95_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4450
  (clk,_zy_sva_brcm_aux_cmd_guid_96_reset_or)
    variable DUMMY103 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_guid_96_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY103 := _zy_sva_b95 ;
      _zy_sva_brcm_aux_cmd_guid_96_ccheck <= "1" ;
      if (DUMMY103 = '1') then
        _zy_sva_brcm_aux_cmd_guid_96_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4467
  (clk,_zy_sva_brcm_aux_cmd_guid_iv_97_reset_or)
    variable DUMMY104 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_guid_iv_97_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY104 := _zy_sva_b96 ;
      _zy_sva_brcm_aux_cmd_guid_iv_97_ccheck <= "1" ;
      if (DUMMY104 = '1') then
        _zy_sva_brcm_aux_cmd_guid_iv_97_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4484
  (clk,_zy_sva_brcm_key_type_98_reset_or)
    variable DUMMY105 : std_logic ;
  begin
    if (_zy_sva_brcm_key_type_98_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY105 := _zy_sva_b97 ;
      _zy_sva_brcm_key_type_98_ccheck <= "1" ;
      if (DUMMY105 = '1') then
        _zy_sva_brcm_key_type_98_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4501
  (clk,_zy_sva_brcm_aux_cmd_99_reset_or)
    variable DUMMY106 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_99_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY106 := _zy_sva_b98 ;
      _zy_sva_brcm_aux_cmd_99_ccheck <= "1" ;
      if (DUMMY106 = '1') then
        _zy_sva_brcm_aux_cmd_99_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4518
  (clk,_zy_sva_brcm_aux_cmd_iv_100_reset_or)
    variable DUMMY107 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_iv_100_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY107 := _zy_sva_b99 ;
      _zy_sva_brcm_aux_cmd_iv_100_ccheck <= "1" ;
      if (DUMMY107 = '1') then
        _zy_sva_brcm_aux_cmd_iv_100_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4535
  (clk,_zy_sva_brcm_aux_cmd_guid_101_reset_or)
    variable DUMMY108 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_guid_101_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY108 := _zy_sva_b100 ;
      _zy_sva_brcm_aux_cmd_guid_101_ccheck <= "1" ;
      if (DUMMY108 = '1') then
        _zy_sva_brcm_aux_cmd_guid_101_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4552
  (clk,_zy_sva_brcm_aux_cmd_guid_iv_102_reset_or)
    variable DUMMY109 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_guid_iv_102_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY109 := _zy_sva_b101 ;
      _zy_sva_brcm_aux_cmd_guid_iv_102_ccheck <= "1" ;
      if (DUMMY109 = '1') then
        _zy_sva_brcm_aux_cmd_guid_iv_102_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4569
  (clk,_zy_sva_brcm_key_type_103_reset_or)
    variable DUMMY110 : std_logic ;
  begin
    if (_zy_sva_brcm_key_type_103_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY110 := _zy_sva_b102 ;
      _zy_sva_brcm_key_type_103_ccheck <= "1" ;
      if (DUMMY110 = '1') then
        _zy_sva_brcm_key_type_103_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4586
  (clk,_zy_sva_brcm_aux_cmd_104_reset_or)
    variable DUMMY111 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_104_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY111 := _zy_sva_b103 ;
      _zy_sva_brcm_aux_cmd_104_ccheck <= "1" ;
      if (DUMMY111 = '1') then
        _zy_sva_brcm_aux_cmd_104_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4603
  (clk,_zy_sva_brcm_aux_cmd_iv_105_reset_or)
    variable DUMMY112 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_iv_105_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY112 := _zy_sva_b104 ;
      _zy_sva_brcm_aux_cmd_iv_105_ccheck <= "1" ;
      if (DUMMY112 = '1') then
        _zy_sva_brcm_aux_cmd_iv_105_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4620
  (clk,_zy_sva_brcm_aux_cmd_guid_106_reset_or)
    variable DUMMY113 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_guid_106_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY113 := _zy_sva_b105 ;
      _zy_sva_brcm_aux_cmd_guid_106_ccheck <= "1" ;
      if (DUMMY113 = '1') then
        _zy_sva_brcm_aux_cmd_guid_106_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4637
  (clk,_zy_sva_brcm_aux_cmd_guid_iv_107_reset_or)
    variable DUMMY114 : std_logic ;
  begin
    if (_zy_sva_brcm_aux_cmd_guid_iv_107_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY114 := _zy_sva_b106 ;
      _zy_sva_brcm_aux_cmd_guid_iv_107_ccheck <= "1" ;
      if (DUMMY114 = '1') then
        _zy_sva_brcm_aux_cmd_guid_iv_107_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4654
  (clk,_zy_sva_brcm_key_type_108_reset_or)
    variable DUMMY115 : std_logic ;
  begin
    if (_zy_sva_brcm_key_type_108_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY115 := _zy_sva_b107 ;
      _zy_sva_brcm_key_type_108_ccheck <= "1" ;
      if (DUMMY115 = '1') then
        _zy_sva_brcm_key_type_108_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4671
  (clk,_zy_sva_brcm_kdf_ops_109_reset_or)
    variable DUMMY116 : std_logic ;
  begin
    if (_zy_sva_brcm_kdf_ops_109_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY116 := _zy_sva_b108 ;
      _zy_sva_brcm_kdf_ops_109_ccheck <= "1" ;
      if (DUMMY116 = '1') then
        _zy_sva_brcm_kdf_ops_109_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4688
  (clk,_zy_sva_brcm_kdf_ops_110_reset_or)
    variable DUMMY117 : std_logic ;
  begin
    if (_zy_sva_brcm_kdf_ops_110_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY117 := _zy_sva_b109 ;
      _zy_sva_brcm_kdf_ops_110_ccheck <= "1" ;
      if (DUMMY117 = '1') then
        _zy_sva_brcm_kdf_ops_110_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4705
  (clk,_zy_sva_brcm_kdf_ops_111_reset_or)
    variable DUMMY118 : std_logic ;
  begin
    if (_zy_sva_brcm_kdf_ops_111_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY118 := _zy_sva_b110 ;
      _zy_sva_brcm_kdf_ops_111_ccheck <= "1" ;
      if (DUMMY118 = '1') then
        _zy_sva_brcm_kdf_ops_111_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4722
  (clk,_zy_sva_brcm_kdf_ops_112_reset_or)
    variable DUMMY119 : std_logic ;
  begin
    if (_zy_sva_brcm_kdf_ops_112_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY119 := _zy_sva_b111 ;
      _zy_sva_brcm_kdf_ops_112_ccheck <= "1" ;
      if (DUMMY119 = '1') then
        _zy_sva_brcm_kdf_ops_112_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4739
  (clk,_zy_sva_brcm_kdf_ops_113_reset_or)
    variable DUMMY120 : std_logic ;
  begin
    if (_zy_sva_brcm_kdf_ops_113_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY120 := _zy_sva_b112 ;
      _zy_sva_brcm_kdf_ops_113_ccheck <= "1" ;
      if (DUMMY120 = '1') then
        _zy_sva_brcm_kdf_ops_113_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4756
  (clk,_zy_sva_brcm_kdf_ops_114_reset_or)
    variable DUMMY121 : std_logic ;
  begin
    if (_zy_sva_brcm_kdf_ops_114_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY121 := _zy_sva_b113 ;
      _zy_sva_brcm_kdf_ops_114_ccheck <= "1" ;
      if (DUMMY121 = '1') then
        _zy_sva_brcm_kdf_ops_114_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4773
  (clk,_zy_sva_brcm_kdf_ops_115_reset_or)
    variable DUMMY122 : std_logic ;
  begin
    if (_zy_sva_brcm_kdf_ops_115_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY122 := _zy_sva_b114 ;
      _zy_sva_brcm_kdf_ops_115_ccheck <= "1" ;
      if (DUMMY122 = '1') then
        _zy_sva_brcm_kdf_ops_115_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4790
  (clk,_zy_sva_brcm_kdf_ops_116_reset_or)
    variable DUMMY123 : std_logic ;
  begin
    if (_zy_sva_brcm_kdf_ops_116_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY123 := _zy_sva_b115 ;
      _zy_sva_brcm_kdf_ops_116_ccheck <= "1" ;
      if (DUMMY123 = '1') then
        _zy_sva_brcm_kdf_ops_116_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4807
  (clk,_zy_sva_brcm_kdf_ops_117_reset_or)
    variable DUMMY124 : std_logic ;
  begin
    if (_zy_sva_brcm_kdf_ops_117_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY124 := _zy_sva_b116 ;
      _zy_sva_brcm_kdf_ops_117_ccheck <= "1" ;
      if (DUMMY124 = '1') then
        _zy_sva_brcm_kdf_ops_117_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4824
  (clk,_zy_sva_brcm_kdf_ops_118_reset_or)
    variable DUMMY125 : std_logic ;
  begin
    if (_zy_sva_brcm_kdf_ops_118_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY125 := _zy_sva_b117 ;
      _zy_sva_brcm_kdf_ops_118_ccheck <= "1" ;
      if (DUMMY125 = '1') then
        _zy_sva_brcm_kdf_ops_118_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4841
  (clk,_zy_sva_brcm_kdf_ops_119_reset_or)
    variable DUMMY126 : std_logic ;
  begin
    if (_zy_sva_brcm_kdf_ops_119_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY126 := _zy_sva_b118 ;
      _zy_sva_brcm_kdf_ops_119_ccheck <= "1" ;
      if (DUMMY126 = '1') then
        _zy_sva_brcm_kdf_ops_119_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4858
  (clk,_zy_sva_brcm_kdf_ops_120_reset_or)
    variable DUMMY127 : std_logic ;
  begin
    if (_zy_sva_brcm_kdf_ops_120_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY127 := _zy_sva_b119 ;
      _zy_sva_brcm_kdf_ops_120_ccheck <= "1" ;
      if (DUMMY127 = '1') then
        _zy_sva_brcm_kdf_ops_120_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4875
  (clk,_zy_sva_brcm_kdf_ops_121_reset_or)
    variable DUMMY128 : std_logic ;
  begin
    if (_zy_sva_brcm_kdf_ops_121_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY128 := _zy_sva_b120 ;
      _zy_sva_brcm_kdf_ops_121_ccheck <= "1" ;
      if (DUMMY128 = '1') then
        _zy_sva_brcm_kdf_ops_121_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4892
  (clk,_zy_sva_brcm_kdf_ops_122_reset_or)
    variable DUMMY129 : std_logic ;
  begin
    if (_zy_sva_brcm_kdf_ops_122_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY129 := _zy_sva_b121 ;
      _zy_sva_brcm_kdf_ops_122_ccheck <= "1" ;
      if (DUMMY129 = '1') then
        _zy_sva_brcm_kdf_ops_122_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4909
  (clk,_zy_sva_brcm_kdf_ops_123_reset_or)
    variable DUMMY130 : std_logic ;
  begin
    if (_zy_sva_brcm_kdf_ops_123_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY130 := _zy_sva_b122 ;
      _zy_sva_brcm_kdf_ops_123_ccheck <= "1" ;
      if (DUMMY130 = '1') then
        _zy_sva_brcm_kdf_ops_123_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4926
  (clk,_zy_sva_brcm_kdf_ops_124_reset_or)
    variable DUMMY131 : std_logic ;
  begin
    if (_zy_sva_brcm_kdf_ops_124_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY131 := _zy_sva_b123 ;
      _zy_sva_brcm_kdf_ops_124_ccheck <= "1" ;
      if (DUMMY131 = '1') then
        _zy_sva_brcm_kdf_ops_124_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4943
  (clk,_zy_sva_null_gcm_125_reset_or)
    variable DUMMY132 : std_logic ;
  begin
    if (_zy_sva_null_gcm_125_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY132 := _zy_sva_b124 ;
      _zy_sva_null_gcm_125_ccheck <= "1" ;
      if (DUMMY132 = '1') then
        _zy_sva_null_gcm_125_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4960
  (clk,_zy_sva_sha_gcm_126_reset_or)
    variable DUMMY133 : std_logic ;
  begin
    if (_zy_sva_sha_gcm_126_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY133 := _zy_sva_b125 ;
      _zy_sva_sha_gcm_126_ccheck <= "1" ;
      if (DUMMY133 = '1') then
        _zy_sva_sha_gcm_126_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4977
  (clk,_zy_sva_null_xts_127_reset_or)
    variable DUMMY134 : std_logic ;
  begin
    if (_zy_sva_null_xts_127_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY134 := _zy_sva_b126 ;
      _zy_sva_null_xts_127_ccheck <= "1" ;
      if (DUMMY134 = '1') then
        _zy_sva_null_xts_127_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o4994
  (clk,_zy_sva_sha_xts_128_reset_or)
    variable DUMMY135 : std_logic ;
  begin
    if (_zy_sva_sha_xts_128_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY135 := _zy_sva_b127 ;
      _zy_sva_sha_xts_128_ccheck <= "1" ;
      if (DUMMY135 = '1') then
        _zy_sva_sha_xts_128_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5011
  (clk,_zy_sva_null_null_129_reset_or)
    variable DUMMY136 : std_logic ;
  begin
    if (_zy_sva_null_null_129_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY136 := _zy_sva_b128 ;
      _zy_sva_null_null_129_ccheck <= "1" ;
      if (DUMMY136 = '1') then
        _zy_sva_null_null_129_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5028
  (clk,_zy_sva_sha_null_130_reset_or)
    variable DUMMY137 : std_logic ;
  begin
    if (_zy_sva_sha_null_130_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY137 := _zy_sva_b129 ;
      _zy_sva_sha_null_130_ccheck <= "1" ;
      if (DUMMY137 = '1') then
        _zy_sva_sha_null_130_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5045
  (clk,_zy_sva_hmac_gcm_131_reset_or)
    variable DUMMY138 : std_logic ;
  begin
    if (_zy_sva_hmac_gcm_131_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY138 := _zy_sva_b130 ;
      _zy_sva_hmac_gcm_131_ccheck <= "1" ;
      if (DUMMY138 = '1') then
        _zy_sva_hmac_gcm_131_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5062
  (clk,_zy_sva_hmac_xts_132_reset_or)
    variable DUMMY139 : std_logic ;
  begin
    if (_zy_sva_hmac_xts_132_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY139 := _zy_sva_b131 ;
      _zy_sva_hmac_xts_132_ccheck <= "1" ;
      if (DUMMY139 = '1') then
        _zy_sva_hmac_xts_132_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5079
  (clk,_zy_sva_hmac_null_133_reset_or)
    variable DUMMY140 : std_logic ;
  begin
    if (_zy_sva_hmac_null_133_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY140 := _zy_sva_b132 ;
      _zy_sva_hmac_null_133_ccheck <= "1" ;
      if (DUMMY140 = '1') then
        _zy_sva_hmac_null_133_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5096
  (clk,_zy_sva_null_gcm_134_reset_or)
    variable DUMMY141 : std_logic ;
  begin
    if (_zy_sva_null_gcm_134_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY141 := _zy_sva_b133 ;
      _zy_sva_null_gcm_134_ccheck <= "1" ;
      if (DUMMY141 = '1') then
        _zy_sva_null_gcm_134_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5113
  (clk,_zy_sva_sha_gcm_135_reset_or)
    variable DUMMY142 : std_logic ;
  begin
    if (_zy_sva_sha_gcm_135_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY142 := _zy_sva_b134 ;
      _zy_sva_sha_gcm_135_ccheck <= "1" ;
      if (DUMMY142 = '1') then
        _zy_sva_sha_gcm_135_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5130
  (clk,_zy_sva_null_xts_136_reset_or)
    variable DUMMY143 : std_logic ;
  begin
    if (_zy_sva_null_xts_136_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY143 := _zy_sva_b135 ;
      _zy_sva_null_xts_136_ccheck <= "1" ;
      if (DUMMY143 = '1') then
        _zy_sva_null_xts_136_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5147
  (clk,_zy_sva_sha_xts_137_reset_or)
    variable DUMMY144 : std_logic ;
  begin
    if (_zy_sva_sha_xts_137_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY144 := _zy_sva_b136 ;
      _zy_sva_sha_xts_137_ccheck <= "1" ;
      if (DUMMY144 = '1') then
        _zy_sva_sha_xts_137_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5164
  (clk,_zy_sva_null_null_138_reset_or)
    variable DUMMY145 : std_logic ;
  begin
    if (_zy_sva_null_null_138_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY145 := _zy_sva_b137 ;
      _zy_sva_null_null_138_ccheck <= "1" ;
      if (DUMMY145 = '1') then
        _zy_sva_null_null_138_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5181
  (clk,_zy_sva_sha_null_139_reset_or)
    variable DUMMY146 : std_logic ;
  begin
    if (_zy_sva_sha_null_139_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY146 := _zy_sva_b138 ;
      _zy_sva_sha_null_139_ccheck <= "1" ;
      if (DUMMY146 = '1') then
        _zy_sva_sha_null_139_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5198
  (clk,_zy_sva_hmac_gcm_140_reset_or)
    variable DUMMY147 : std_logic ;
  begin
    if (_zy_sva_hmac_gcm_140_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY147 := _zy_sva_b139 ;
      _zy_sva_hmac_gcm_140_ccheck <= "1" ;
      if (DUMMY147 = '1') then
        _zy_sva_hmac_gcm_140_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5215
  (clk,_zy_sva_hmac_xts_141_reset_or)
    variable DUMMY148 : std_logic ;
  begin
    if (_zy_sva_hmac_xts_141_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY148 := _zy_sva_b140 ;
      _zy_sva_hmac_xts_141_ccheck <= "1" ;
      if (DUMMY148 = '1') then
        _zy_sva_hmac_xts_141_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5232
  (clk,_zy_sva_hmac_null_142_reset_or)
    variable DUMMY149 : std_logic ;
  begin
    if (_zy_sva_hmac_null_142_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY149 := _zy_sva_b141 ;
      _zy_sva_hmac_null_142_ccheck <= "1" ;
      if (DUMMY149 = '1') then
        _zy_sva_hmac_null_142_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5249
  (clk,_zy_sva_null_gcm_143_reset_or)
    variable DUMMY150 : std_logic ;
  begin
    if (_zy_sva_null_gcm_143_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY150 := _zy_sva_b142 ;
      _zy_sva_null_gcm_143_ccheck <= "1" ;
      if (DUMMY150 = '1') then
        _zy_sva_null_gcm_143_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5266
  (clk,_zy_sva_sha_gcm_144_reset_or)
    variable DUMMY151 : std_logic ;
  begin
    if (_zy_sva_sha_gcm_144_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY151 := _zy_sva_b143 ;
      _zy_sva_sha_gcm_144_ccheck <= "1" ;
      if (DUMMY151 = '1') then
        _zy_sva_sha_gcm_144_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5283
  (clk,_zy_sva_null_xts_145_reset_or)
    variable DUMMY152 : std_logic ;
  begin
    if (_zy_sva_null_xts_145_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY152 := _zy_sva_b144 ;
      _zy_sva_null_xts_145_ccheck <= "1" ;
      if (DUMMY152 = '1') then
        _zy_sva_null_xts_145_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5300
  (clk,_zy_sva_sha_xts_146_reset_or)
    variable DUMMY153 : std_logic ;
  begin
    if (_zy_sva_sha_xts_146_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY153 := _zy_sva_b145 ;
      _zy_sva_sha_xts_146_ccheck <= "1" ;
      if (DUMMY153 = '1') then
        _zy_sva_sha_xts_146_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5317
  (clk,_zy_sva_null_null_147_reset_or)
    variable DUMMY154 : std_logic ;
  begin
    if (_zy_sva_null_null_147_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY154 := _zy_sva_b146 ;
      _zy_sva_null_null_147_ccheck <= "1" ;
      if (DUMMY154 = '1') then
        _zy_sva_null_null_147_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5334
  (clk,_zy_sva_sha_null_148_reset_or)
    variable DUMMY155 : std_logic ;
  begin
    if (_zy_sva_sha_null_148_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY155 := _zy_sva_b147 ;
      _zy_sva_sha_null_148_ccheck <= "1" ;
      if (DUMMY155 = '1') then
        _zy_sva_sha_null_148_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5351
  (clk,_zy_sva_hmac_gcm_149_reset_or)
    variable DUMMY156 : std_logic ;
  begin
    if (_zy_sva_hmac_gcm_149_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY156 := _zy_sva_b148 ;
      _zy_sva_hmac_gcm_149_ccheck <= "1" ;
      if (DUMMY156 = '1') then
        _zy_sva_hmac_gcm_149_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5368
  (clk,_zy_sva_hmac_xts_150_reset_or)
    variable DUMMY157 : std_logic ;
  begin
    if (_zy_sva_hmac_xts_150_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY157 := _zy_sva_b149 ;
      _zy_sva_hmac_xts_150_ccheck <= "1" ;
      if (DUMMY157 = '1') then
        _zy_sva_hmac_xts_150_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5385
  (clk,_zy_sva_hmac_null_151_reset_or)
    variable DUMMY158 : std_logic ;
  begin
    if (_zy_sva_hmac_null_151_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY158 := _zy_sva_b150 ;
      _zy_sva_hmac_null_151_ccheck <= "1" ;
      if (DUMMY158 = '1') then
        _zy_sva_hmac_null_151_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5402
  (clk,_zy_sva_null_gcm_152_reset_or)
    variable DUMMY159 : std_logic ;
  begin
    if (_zy_sva_null_gcm_152_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY159 := _zy_sva_b151 ;
      _zy_sva_null_gcm_152_ccheck <= "1" ;
      if (DUMMY159 = '1') then
        _zy_sva_null_gcm_152_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5419
  (clk,_zy_sva_sha_gcm_153_reset_or)
    variable DUMMY160 : std_logic ;
  begin
    if (_zy_sva_sha_gcm_153_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY160 := _zy_sva_b152 ;
      _zy_sva_sha_gcm_153_ccheck <= "1" ;
      if (DUMMY160 = '1') then
        _zy_sva_sha_gcm_153_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5436
  (clk,_zy_sva_null_xts_154_reset_or)
    variable DUMMY161 : std_logic ;
  begin
    if (_zy_sva_null_xts_154_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY161 := _zy_sva_b153 ;
      _zy_sva_null_xts_154_ccheck <= "1" ;
      if (DUMMY161 = '1') then
        _zy_sva_null_xts_154_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5453
  (clk,_zy_sva_sha_xts_155_reset_or)
    variable DUMMY162 : std_logic ;
  begin
    if (_zy_sva_sha_xts_155_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY162 := _zy_sva_b154 ;
      _zy_sva_sha_xts_155_ccheck <= "1" ;
      if (DUMMY162 = '1') then
        _zy_sva_sha_xts_155_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5470
  (clk,_zy_sva_null_null_156_reset_or)
    variable DUMMY163 : std_logic ;
  begin
    if (_zy_sva_null_null_156_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY163 := _zy_sva_b155 ;
      _zy_sva_null_null_156_ccheck <= "1" ;
      if (DUMMY163 = '1') then
        _zy_sva_null_null_156_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5487
  (clk,_zy_sva_sha_null_157_reset_or)
    variable DUMMY164 : std_logic ;
  begin
    if (_zy_sva_sha_null_157_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY164 := _zy_sva_b156 ;
      _zy_sva_sha_null_157_ccheck <= "1" ;
      if (DUMMY164 = '1') then
        _zy_sva_sha_null_157_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5504
  (clk,_zy_sva_hmac_gcm_158_reset_or)
    variable DUMMY165 : std_logic ;
  begin
    if (_zy_sva_hmac_gcm_158_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY165 := _zy_sva_b157 ;
      _zy_sva_hmac_gcm_158_ccheck <= "1" ;
      if (DUMMY165 = '1') then
        _zy_sva_hmac_gcm_158_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5521
  (clk,_zy_sva_hmac_xts_159_reset_or)
    variable DUMMY166 : std_logic ;
  begin
    if (_zy_sva_hmac_xts_159_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY166 := _zy_sva_b158 ;
      _zy_sva_hmac_xts_159_ccheck <= "1" ;
      if (DUMMY166 = '1') then
        _zy_sva_hmac_xts_159_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5538
  (clk,_zy_sva_hmac_null_160_reset_or)
    variable DUMMY167 : std_logic ;
  begin
    if (_zy_sva_hmac_null_160_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY167 := _zy_sva_b159 ;
      _zy_sva_hmac_null_160_ccheck <= "1" ;
      if (DUMMY167 = '1') then
        _zy_sva_hmac_null_160_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5555
  (clk,_zy_sva_null_gcm_161_reset_or)
    variable DUMMY168 : std_logic ;
  begin
    if (_zy_sva_null_gcm_161_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY168 := _zy_sva_b160 ;
      _zy_sva_null_gcm_161_ccheck <= "1" ;
      if (DUMMY168 = '1') then
        _zy_sva_null_gcm_161_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5572
  (clk,_zy_sva_sha_gcm_162_reset_or)
    variable DUMMY169 : std_logic ;
  begin
    if (_zy_sva_sha_gcm_162_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY169 := _zy_sva_b161 ;
      _zy_sva_sha_gcm_162_ccheck <= "1" ;
      if (DUMMY169 = '1') then
        _zy_sva_sha_gcm_162_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5589
  (clk,_zy_sva_null_xts_163_reset_or)
    variable DUMMY170 : std_logic ;
  begin
    if (_zy_sva_null_xts_163_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY170 := _zy_sva_b162 ;
      _zy_sva_null_xts_163_ccheck <= "1" ;
      if (DUMMY170 = '1') then
        _zy_sva_null_xts_163_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5606
  (clk,_zy_sva_sha_xts_164_reset_or)
    variable DUMMY171 : std_logic ;
  begin
    if (_zy_sva_sha_xts_164_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY171 := _zy_sva_b163 ;
      _zy_sva_sha_xts_164_ccheck <= "1" ;
      if (DUMMY171 = '1') then
        _zy_sva_sha_xts_164_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5623
  (clk,_zy_sva_null_null_165_reset_or)
    variable DUMMY172 : std_logic ;
  begin
    if (_zy_sva_null_null_165_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY172 := _zy_sva_b164 ;
      _zy_sva_null_null_165_ccheck <= "1" ;
      if (DUMMY172 = '1') then
        _zy_sva_null_null_165_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5640
  (clk,_zy_sva_sha_null_166_reset_or)
    variable DUMMY173 : std_logic ;
  begin
    if (_zy_sva_sha_null_166_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY173 := _zy_sva_b165 ;
      _zy_sva_sha_null_166_ccheck <= "1" ;
      if (DUMMY173 = '1') then
        _zy_sva_sha_null_166_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5657
  (clk,_zy_sva_hmac_gcm_167_reset_or)
    variable DUMMY174 : std_logic ;
  begin
    if (_zy_sva_hmac_gcm_167_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY174 := _zy_sva_b166 ;
      _zy_sva_hmac_gcm_167_ccheck <= "1" ;
      if (DUMMY174 = '1') then
        _zy_sva_hmac_gcm_167_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5674
  (clk,_zy_sva_hmac_xts_168_reset_or)
    variable DUMMY175 : std_logic ;
  begin
    if (_zy_sva_hmac_xts_168_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY175 := _zy_sva_b167 ;
      _zy_sva_hmac_xts_168_ccheck <= "1" ;
      if (DUMMY175 = '1') then
        _zy_sva_hmac_xts_168_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5691
  (clk,_zy_sva_hmac_null_169_reset_or)
    variable DUMMY176 : std_logic ;
  begin
    if (_zy_sva_hmac_null_169_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY176 := _zy_sva_b168 ;
      _zy_sva_hmac_null_169_ccheck <= "1" ;
      if (DUMMY176 = '1') then
        _zy_sva_hmac_null_169_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5708
  (clk,_zy_sva_null_gcm_170_reset_or)
    variable DUMMY177 : std_logic ;
  begin
    if (_zy_sva_null_gcm_170_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY177 := _zy_sva_b169 ;
      _zy_sva_null_gcm_170_ccheck <= "1" ;
      if (DUMMY177 = '1') then
        _zy_sva_null_gcm_170_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5725
  (clk,_zy_sva_sha_gcm_171_reset_or)
    variable DUMMY178 : std_logic ;
  begin
    if (_zy_sva_sha_gcm_171_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY178 := _zy_sva_b170 ;
      _zy_sva_sha_gcm_171_ccheck <= "1" ;
      if (DUMMY178 = '1') then
        _zy_sva_sha_gcm_171_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5742
  (clk,_zy_sva_null_xts_172_reset_or)
    variable DUMMY179 : std_logic ;
  begin
    if (_zy_sva_null_xts_172_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY179 := _zy_sva_b171 ;
      _zy_sva_null_xts_172_ccheck <= "1" ;
      if (DUMMY179 = '1') then
        _zy_sva_null_xts_172_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5759
  (clk,_zy_sva_sha_xts_173_reset_or)
    variable DUMMY180 : std_logic ;
  begin
    if (_zy_sva_sha_xts_173_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY180 := _zy_sva_b172 ;
      _zy_sva_sha_xts_173_ccheck <= "1" ;
      if (DUMMY180 = '1') then
        _zy_sva_sha_xts_173_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5776
  (clk,_zy_sva_null_null_174_reset_or)
    variable DUMMY181 : std_logic ;
  begin
    if (_zy_sva_null_null_174_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY181 := _zy_sva_b173 ;
      _zy_sva_null_null_174_ccheck <= "1" ;
      if (DUMMY181 = '1') then
        _zy_sva_null_null_174_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5793
  (clk,_zy_sva_sha_null_175_reset_or)
    variable DUMMY182 : std_logic ;
  begin
    if (_zy_sva_sha_null_175_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY182 := _zy_sva_b174 ;
      _zy_sva_sha_null_175_ccheck <= "1" ;
      if (DUMMY182 = '1') then
        _zy_sva_sha_null_175_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5810
  (clk,_zy_sva_hmac_gcm_176_reset_or)
    variable DUMMY183 : std_logic ;
  begin
    if (_zy_sva_hmac_gcm_176_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY183 := _zy_sva_b175 ;
      _zy_sva_hmac_gcm_176_ccheck <= "1" ;
      if (DUMMY183 = '1') then
        _zy_sva_hmac_gcm_176_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5827
  (clk,_zy_sva_hmac_xts_177_reset_or)
    variable DUMMY184 : std_logic ;
  begin
    if (_zy_sva_hmac_xts_177_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY184 := _zy_sva_b176 ;
      _zy_sva_hmac_xts_177_ccheck <= "1" ;
      if (DUMMY184 = '1') then
        _zy_sva_hmac_xts_177_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5844
  (clk,_zy_sva_hmac_null_178_reset_or)
    variable DUMMY185 : std_logic ;
  begin
    if (_zy_sva_hmac_null_178_reset_or = '1') then
    elsif (clk'event and clk = '1') then
      DUMMY185 := _zy_sva_b177 ;
      _zy_sva_hmac_null_178_ccheck <= "1" ;
      if (DUMMY185 = '1') then
        _zy_sva_hmac_null_178_cpass <= "1" ;
      end if;
    end if ;
  end process ;

  process --:o5861
  (clk,rst_n)
  begin
    if (rst_n = '0') then
      tlv_counter <= "00000" ;
    elsif (clk'event and clk = '1') then
      if (stitcher_rd = '1') then
        if (stitcher_eot = '1') then
          tlv_counter <= "00000" ;
        else
          tlv_counter <= (tlv_counter + std_logic_vector'("00001")) ;
        end if;
      end if;
    end if ;
  end process ;

  process --:o5881
  (clk,rst_n)
  begin
    if (rst_n = '0') then
      tlv_type <= RQE ;
      aux_key_type <= NO_AUX_KEY ;
      aux_iv_op <= IV_SRC ;
      aux_cipher_op <= CPH_NULL ;
      aux_auth_op <= AUTH_NULL ;
      aux_raw_auth_op <= AUTH_NULL ;
      kme_internal_word0 <=
       "0000000000000000000000000000000000000000000000000000000000000000" ;
      kme_internal_dek_kim_word <=
       "0000000000000000000000000000000000000000000000000000000000000000" ;
      kme_internal_dak_kim_word <=
       "0000000000000000000000000000000000000000000000000000000000000000" ;
      debug_cmd <= "00000000000000000000000000000000" ;
      aux_key_header <= "00000000000000000000000000000000" ;
      skip <= "0000000" ;
      guid0 <=
       "0000000000000000000000000000000000000000000000000000000000000000" ;
      guid1 <=
       "0000000000000000000000000000000000000000000000000000000000000000" ;
      guid2 <=
       "0000000000000000000000000000000000000000000000000000000000000000" ;
      guid3 <=
       "0000000000000000000000000000000000000000000000000000000000000000" ;
      iv0 <= "0000000000000000000000000000000000000000000000000000000000000000"
       ;
      iv1 <= "0000000000000000000000000000000000000000000000000000000000000000"
       ;
      DUMMY7 <= "00000000000000000000000000000000" ;
      fifo_in(64+3 downto 64) <= KME_WORD0 ;
    elsif (clk'event and clk = '1') then
      tlv_type <= nxt_tlv_type ;
      aux_key_type <= nxt_aux_key_type ;
      aux_iv_op <= nxt_aux_iv_op ;
      aux_cipher_op <= nxt_aux_cipher_op ;
      aux_auth_op <= nxt_aux_auth_op ;
      aux_raw_auth_op <= nxt_aux_raw_auth_op ;
      kme_internal_word0 <= nxt_kme_internal_word0 ;
      kme_internal_dek_kim_word <= nxt_kme_internal_dek_kim_word ;
      kme_internal_dak_kim_word <= nxt_kme_internal_dak_kim_word ;
      debug_cmd <= nxt_debug_cmd ;
      aux_key_header <= nxt_aux_key_header ;
      skip <= nxt_skip ;
      guid0 <= nxt_guid0 ;
      guid1 <= nxt_guid1 ;
      guid2 <= nxt_guid2 ;
      guid3 <= nxt_guid3 ;
      iv0 <= nxt_iv0 ;
      iv1 <= nxt_iv1 ;
      DUMMY7 <= nxt_buffer ;
      fifo_in(64+3 downto 64) <= nxt_fifo_in_id ;
    end if ;
  end process ;

  process --:o5931
  (*)
    variable fifo_in_DUMMY0 : kme_internal_t ;
    variable nxt_kme_internal_word0_DUMMY1 : kme_internal_word_0_t ;
    variable nxt_aux_key_header_DUMMY2 : aux_key_ctrl_t ;
    variable nxt_buffer_DUMMY3 : std_logic_vector(31 downto 0) ;
    variable tlv_word0_DUMMY4 : tlv_rqe_word_0_t ;
    variable tlv_word1_DUMMY5 : tlv_rqe_word_1_t ;
    variable tlv_word2_DUMMY6 : tlv_cmd_word_2_t ;
    variable frame_word_DUMMY7 : tlv_cmd_word_1_t ;
    variable stitcher_rd_DUMMY8 : std_logic ;
    variable DUMMY186 : std_logic_vector(63 downto 0) ;
    variable _zyL234_tfiRv52_DUMMY9 : std_logic_vector(63 downto 0) ;
    variable DUMMY187 : std_logic ;
    variable DUMMY188 : aux_key_type_e ;
    variable DUMMY189 : cmd_cipher_op_e ;
    variable DUMMY190 : aux_kdf_mode_e ;
    variable DUMMY191 : std_logic ;
    variable DUMMY192 : std_logic ;
    variable DUMMY193 : std_logic ;
    variable DUMMY194 : std_logic ;
    variable _zyL252_tfiRv53_DUMMY10 : std_logic ;
    variable DUMMY195 : cmd_cipher_op_e ;
    variable DUMMY196 : aux_kdf_mode_e ;
    variable DUMMY197 : cmd_cipher_op_e ;
    variable DUMMY198 : aux_kdf_mode_e ;
    variable DUMMY199 : tlv_types_e ;
    variable DUMMY200 : aux_kdf_mode_e ;
    variable DUMMY201 : aux_key_op_e ;
    variable DUMMY202 : aux_key_op_e ;
    variable _zyL253_tfiRv54_DUMMY11 : std_logic ;
    variable DUMMY203 : tlv_types_e ;
    variable DUMMY204 : cmd_iv_op_e ;
    variable DUMMY205 : cmd_cipher_op_e ;
    variable DUMMY206 : std_logic ;
    variable DUMMY207 : cmd_cipher_op_e ;
    variable _zyL254_tfiRv55_DUMMY12 : std_logic ;
    variable DUMMY208 : std_logic ;
    variable DUMMY209 : aux_key_type_e ;
    variable DUMMY210 : cmd_auth_op_e ;
    variable DUMMY211 : cmd_auth_op_e ;
    variable DUMMY212 : std_logic ;
    variable DUMMY213 : std_logic ;
    variable DUMMY214 : std_logic ;
    variable _zyL255_tfiRv56_DUMMY13 : std_logic ;
    variable DUMMY215 : cmd_auth_op_e ;
    variable DUMMY216 : cmd_auth_op_e ;
    variable DUMMY217 : cmd_auth_op_e ;
    variable DUMMY218 : cmd_auth_op_e ;
    variable DUMMY219 : cmd_auth_op_e ;
    variable DUMMY220 : cmd_auth_op_e ;
    variable DUMMY221 : std_logic_vector(63 downto 0) ;
    variable _zyL288_tfiRv57_DUMMY14 : std_logic_vector(63 downto 0) ;
    variable DUMMY222 : std_logic_vector(63 downto 0) ;
    variable _zyL293_tfiRv58_DUMMY15 : std_logic_vector(63 downto 0) ;
    variable DUMMY223 : std_logic_vector(63 downto 0) ;
    variable _zyL301_tfiRv59_DUMMY16 : std_logic_vector(63 downto 0) ;
    variable DUMMY224 : std_logic_vector(63 downto 0) ;
    variable _zyL306_tfiRv60_DUMMY17 : std_logic_vector(63 downto 0) ;
    variable DUMMY225 : std_logic_vector(63 downto 0) ;
    variable _zyL313_tfiRv61_DUMMY18 : std_logic_vector(63 downto 0) ;
    variable DUMMY226 : std_logic_vector(63 downto 0) ;
    variable _zyL321_tfiRv62_DUMMY19 : std_logic_vector(63 downto 0) ;
    variable DUMMY227 : std_logic_vector(63 downto 0) ;
    variable _zyL327_tfiRv63_DUMMY20 : std_logic_vector(63 downto 0) ;
    variable DUMMY228 : std_logic_vector(63 downto 0) ;
    variable _zyL337_tfiRv64_DUMMY21 : std_logic_vector(63 downto 0) ;
    variable DUMMY229 : std_logic_vector(63 downto 0) ;
    variable _zyL346_tfiRv65_DUMMY22 : std_logic_vector(63 downto 0) ;
    variable DUMMY230 : std_logic_vector(63 downto 0) ;
    variable _zyL354_tfiRv66_DUMMY23 : std_logic_vector(63 downto 0) ;
    variable DUMMY231 : std_logic_vector(63 downto 0) ;
    variable _zyL359_tfiRv67_DUMMY24 : std_logic_vector(63 downto 0) ;
    variable DUMMY232 : std_logic_vector(63 downto 0) ;
    variable _zyL368_tfiRv68_DUMMY25 : std_logic_vector(63 downto 0) ;
    variable DUMMY233 : std_logic_vector(63 downto 0) ;
    variable _zyL373_tfiRv69_DUMMY26 : std_logic_vector(63 downto 0) ;
    variable DUMMY234 : std_logic_vector(63 downto 0) ;
    variable _zyL382_tfiRv70_DUMMY27 : std_logic_vector(63 downto 0) ;
    variable DUMMY235 : std_logic_vector(63 downto 0) ;
    variable _zyL390_tfiRv71_DUMMY28 : std_logic_vector(63 downto 0) ;
    variable DUMMY236 : std_logic_vector(63 downto 0) ;
    variable _zyL395_tfiRv72_DUMMY29 : std_logic_vector(63 downto 0) ;
    variable DUMMY237 : std_logic_vector(63 downto 0) ;
    variable _zyL410_tfiRv73_DUMMY30 : std_logic_vector(63 downto 0) ;
    variable DUMMY238 : std_logic ;
    variable DUMMY239 : aux_key_type_e ;
    variable DUMMY240 : cmd_cipher_op_e ;
    variable DUMMY241 : std_logic ;
    variable DUMMY242 : std_logic ;
    variable _zyL485_tfiRv74_DUMMY31 : std_logic ;
    variable DUMMY243 : cmd_cipher_op_e ;
    variable DUMMY244 : cmd_cipher_op_e ;
    variable DUMMY245 : std_logic ;
    variable DUMMY246 : aux_key_type_e ;
    variable DUMMY247 : cmd_auth_op_e ;
    variable DUMMY248 : cmd_auth_op_e ;
    variable DUMMY249 : std_logic ;
    variable DUMMY250 : std_logic ;
    variable DUMMY251 : std_logic ;
    variable _zyL486_tfiRv75_DUMMY32 : std_logic ;
    variable DUMMY252 : cmd_auth_op_e ;
    variable DUMMY253 : cmd_auth_op_e ;
    variable DUMMY254 : cmd_auth_op_e ;
    variable DUMMY255 : cmd_auth_op_e ;
    variable DUMMY256 : cmd_auth_op_e ;
    variable DUMMY257 : cmd_auth_op_e ;
    variable DUMMY258 : cmd_cipher_op_e ;
    variable _zyL489_tfiRv76_DUMMY33 : std_logic ;
    variable DUMMY259 : cmd_auth_op_e ;
    variable DUMMY260 : cmd_auth_op_e ;
    variable _zyL489_tfiRv77_DUMMY34 : std_logic ;
    variable DUMMY261 : cmd_cipher_op_e ;
    variable _zyL492_tfiRv78_DUMMY35 : std_logic ;
    variable DUMMY262 : std_logic_vector(63 downto 0) ;
    variable _zyL526_tfiRv79_DUMMY36 : std_logic_vector(63 downto 0) ;
    variable DUMMY263 : std_logic_vector(63 downto 0) ;
    variable _zyL527_tfiRv80_DUMMY37 : std_logic_vector(63 downto 0) ;
    variable DUMMY264 : std_logic_vector(1 to 64) ;
    variable DUMMY265 : std_logic_vector(63 downto 0) ;
    variable _zyL541_tfiRv81_DUMMY38 : std_logic_vector(63 downto 0) ;
    variable DUMMY266 : std_logic_vector(63 downto 0) ;
    variable _zyL542_tfiRv82_DUMMY39 : std_logic_vector(63 downto 0) ;
    variable DUMMY267 : std_logic_vector(63 downto 0) ;
    variable _zyL555_tfiRv83_DUMMY40 : std_logic_vector(63 downto 0) ;
    variable DUMMY268 : std_logic_vector(63 downto 0) ;
    variable _zyL556_tfiRv84_DUMMY41 : std_logic_vector(63 downto 0) ;
    variable DUMMY269 : std_logic_vector(1 to 64) ;
    variable DUMMY270 : std_logic_vector(63 downto 0) ;
    variable _zyL569_tfiRv85_DUMMY42 : std_logic_vector(63 downto 0) ;
    variable DUMMY271 : std_logic_vector(63 downto 0) ;
    variable _zyL570_tfiRv86_DUMMY43 : std_logic_vector(63 downto 0) ;
    variable DUMMY272 : std_logic_vector(1 to 64) ;
    variable DUMMY273 : std_logic_vector(1 to 64) ;
  begin
    fifo_in_DUMMY0 := fifo_in;
    nxt_kme_internal_word0_DUMMY1 := nxt_kme_internal_word0;
    nxt_aux_key_header_DUMMY2 := nxt_aux_key_header;
    nxt_buffer_DUMMY3 := nxt_buffer;
    tlv_word0_DUMMY4 := tlv_word0;
    tlv_word1_DUMMY5 := tlv_word1;
    tlv_word2_DUMMY6 := tlv_word2;
    frame_word_DUMMY7 := frame_word;
    stitcher_rd_DUMMY8 := stitcher_rd;
    _zyL234_tfiRv52_DUMMY9 := _zyL234_tfiRv52;
    _zyL252_tfiRv53_DUMMY10 := _zyL252_tfiRv53;
    _zyL253_tfiRv54_DUMMY11 := _zyL253_tfiRv54;
    _zyL254_tfiRv55_DUMMY12 := _zyL254_tfiRv55;
    _zyL255_tfiRv56_DUMMY13 := _zyL255_tfiRv56;
    _zyL288_tfiRv57_DUMMY14 := _zyL288_tfiRv57;
    _zyL293_tfiRv58_DUMMY15 := _zyL293_tfiRv58;
    _zyL301_tfiRv59_DUMMY16 := _zyL301_tfiRv59;
    _zyL306_tfiRv60_DUMMY17 := _zyL306_tfiRv60;
    _zyL313_tfiRv61_DUMMY18 := _zyL313_tfiRv61;
    _zyL321_tfiRv62_DUMMY19 := _zyL321_tfiRv62;
    _zyL327_tfiRv63_DUMMY20 := _zyL327_tfiRv63;
    _zyL337_tfiRv64_DUMMY21 := _zyL337_tfiRv64;
    _zyL346_tfiRv65_DUMMY22 := _zyL346_tfiRv65;
    _zyL354_tfiRv66_DUMMY23 := _zyL354_tfiRv66;
    _zyL359_tfiRv67_DUMMY24 := _zyL359_tfiRv67;
    _zyL368_tfiRv68_DUMMY25 := _zyL368_tfiRv68;
    _zyL373_tfiRv69_DUMMY26 := _zyL373_tfiRv69;
    _zyL382_tfiRv70_DUMMY27 := _zyL382_tfiRv70;
    _zyL390_tfiRv71_DUMMY28 := _zyL390_tfiRv71;
    _zyL395_tfiRv72_DUMMY29 := _zyL395_tfiRv72;
    _zyL410_tfiRv73_DUMMY30 := _zyL410_tfiRv73;
    _zyL485_tfiRv74_DUMMY31 := _zyL485_tfiRv74;
    _zyL486_tfiRv75_DUMMY32 := _zyL486_tfiRv75;
    _zyL489_tfiRv76_DUMMY33 := _zyL489_tfiRv76;
    _zyL489_tfiRv77_DUMMY34 := _zyL489_tfiRv77;
    _zyL492_tfiRv78_DUMMY35 := _zyL492_tfiRv78;
    _zyL526_tfiRv79_DUMMY36 := _zyL526_tfiRv79;
    _zyL527_tfiRv80_DUMMY37 := _zyL527_tfiRv80;
    _zyL541_tfiRv81_DUMMY38 := _zyL541_tfiRv81;
    _zyL542_tfiRv82_DUMMY39 := _zyL542_tfiRv82;
    _zyL555_tfiRv83_DUMMY40 := _zyL555_tfiRv83;
    _zyL556_tfiRv84_DUMMY41 := _zyL556_tfiRv84;
    _zyL569_tfiRv85_DUMMY42 := _zyL569_tfiRv85;
    _zyL570_tfiRv86_DUMMY43 := _zyL570_tfiRv86;
    fifo_in_DUMMY0(63 downto 0) :=
     "0000000000000000000000000000000000000000000000000000000000000000" ;
    fifo_in_valid <= '0' ;
    nxt_tlv_type <= tlv_type ;
    nxt_aux_key_type <= aux_key_type ;
    nxt_aux_iv_op <= aux_iv_op ;
    nxt_aux_cipher_op <= aux_cipher_op ;
    nxt_aux_auth_op <= aux_auth_op ;
    nxt_aux_raw_auth_op <= aux_raw_auth_op ;
    nxt_kme_internal_word0_DUMMY1 := kme_internal_word0 ;
    nxt_kme_internal_dek_kim_word <= kme_internal_dek_kim_word ;
    nxt_kme_internal_dak_kim_word <= kme_internal_dak_kim_word ;
    nxt_aux_key_header_DUMMY2 := aux_key_header ;
    nxt_debug_cmd <= debug_cmd ;
    nxt_skip <= skip ;
    nxt_guid0 <= guid0 ;
    nxt_guid1 <= guid1 ;
    nxt_guid2 <= guid2 ;
    nxt_guid3 <= guid3 ;
    nxt_iv0 <= iv0 ;
    nxt_iv1 <= iv1 ;
    nxt_buffer_DUMMY3 := DUMMY7 ;
    tlv_word0_DUMMY4 := stitcher_out(63 downto 0) ;
    tlv_word1_DUMMY5 := stitcher_out(63 downto 0) ;
    tlv_word2_DUMMY6 := stitcher_out(63 downto 0) ;
    frame_word_DUMMY7 := stitcher_out(63 downto 0) ;
    stitcher_rd_DUMMY8 := ((not(stitcher_empty) and not(fifo_in_stall)) and not
    (it_conv_std_logic(skip(6 downto 6)))) ;
    if ((fifo_in_stall = '0')) then
      if (skip(6 downto 6) /= "0") then
        if (fifo_in_DUMMY0(64+3 downto 64) = skip(3 downto 0)) then
          nxt_skip(6 downto 6) <= "0" ;
        else
          fifo_in_valid <= '1' ;
        end if;
        if (skip(5 downto 5) /= "0") then
          nxt_skip(5 downto 5) <= "0" ;
          nxt_skip(4 downto 4) <= "0" ;
          DUMMY186 := std_logic_vector'(std_logic_vector'
          ("00000000000000000000000000000000") & DUMMY7) ;
          _zyL234_tfiRv52_DUMMY9 := std_logic_vector'(DUMMY186(7 downto 0) &
           DUMMY186(15 downto 8) & DUMMY186(23 downto 16) & DUMMY186(31 downto
           24) & DUMMY186(39 downto 32) & DUMMY186(47 downto 40) & DUMMY186(55
           downto 48) & DUMMY186(63 downto 56)) ;
          fifo_in_DUMMY0(63 downto 0) := it_cond_op((skip(4 downto 4)
          )/="0",_zyL234_tfiRv52_DUMMY9,std_logic_vector'(DUMMY7 &
           std_logic_vector'("00000000000000000000000000000000"))) ;
        end if;

        case int_tlv_counter is
          when  "000010"  =>
            fifo_in_DUMMY0(63 downto 0) := guid0 ;
          when  "000011"  =>
            fifo_in_DUMMY0(63 downto 0) := guid1 ;
          when  "000100"  =>
            fifo_in_DUMMY0(63 downto 0) := guid2 ;
          when  "000101"  =>
            fifo_in_DUMMY0(63 downto 0) := guid3 ;
          when  "000110"  =>
            fifo_in_DUMMY0(63 downto 0) := iv0 ;
          when  "000111"  =>
            fifo_in_DUMMY0(63 downto 0) := iv1 ;
          when  "001000"  =>
            fifo_in_DUMMY0(63 downto 0) := kme_internal_dek_kim_word ;
          when  "001001"  =>
            fifo_in_DUMMY0(63 downto 0) := kme_internal_dak_kim_word ;
          when others => null ;
        end case;
        if (int_tlv_counter = IDX_KME_IVTWEAK) then
          DUMMY187 := always_validate_kim_ref ;
          DUMMY188 := aux_key_type ;
          DUMMY189 := aux_cipher_op ;
          DUMMY190 := aux_key_header(15+1 downto 15) ;
          _zyL252_tfiRv53_DUMMY10 := '1' ;
          if ((DUMMY187 = '0')) then

            case DUMMY188 is
              when  "000000"  =>
                _zyL252_tfiRv53_DUMMY10 := '0' ;
              when  "000001"  =>
                DUMMY195 := DUMMY189 ;
                DUMMY191 := not(((boolean_to_std(DUMMY195 = AES_GCM) or
                 boolean_to_std(DUMMY195 = AES_XTS_XEX)) or boolean_to_std
                (DUMMY195 = AES_GMAC))) ;
                DUMMY196 := DUMMY190 ;
                DUMMY192 := (boolean_to_std(DUMMY196 = KDF_MODE_GUID) or
                 boolean_to_std(DUMMY196 = KDF_MODE_RGUID)) ;
                if (((DUMMY191)='1' and (DUMMY192)='1')) then
                  _zyL252_tfiRv53_DUMMY10 := '0' ;
                end if;
              when  "001001"  =>
                DUMMY197 := DUMMY189 ;
                DUMMY193 := not(((boolean_to_std(DUMMY197 = AES_GCM) or
                 boolean_to_std(DUMMY197 = AES_XTS_XEX)) or boolean_to_std
                (DUMMY197 = AES_GMAC))) ;
                DUMMY198 := DUMMY190 ;
                DUMMY194 := (boolean_to_std(DUMMY198 = KDF_MODE_GUID) or
                 boolean_to_std(DUMMY198 = KDF_MODE_RGUID)) ;
                if (((DUMMY193)='1' and (DUMMY194)='1')) then
                  _zyL252_tfiRv53_DUMMY10 := '0' ;
                end if;
              when others => null ;
            end case;
          end if;
          nxt_kme_internal_dek_kim_word(17 downto 17) <= ext
          (_zyL252_tfiRv53_DUMMY10,1) ;
          DUMMY199 := tlv_type ;
          DUMMY200 := aux_key_header(15+1 downto 15) ;
          DUMMY201 := aux_key_header(14 downto 14) ;
          DUMMY202 := aux_key_header(31 downto 31) ;
          _zyL253_tfiRv54_DUMMY11 := boolean_to_std(((DUMMY199 = AUX_CMD or
           DUMMY199 = AUX_CMD_IV) and (it_conv_std_logic(DUMMY201) = '1' or
           it_conv_std_logic(DUMMY202) = '1') and (DUMMY200 = KDF_MODE_GUID or
           DUMMY200 = KDF_MODE_COMB_GUID))) ;
          nxt_kme_internal_dek_kim_word(18 downto 18) <= ext
          (_zyL253_tfiRv54_DUMMY11,1) ;
          DUMMY203 := tlv_type ;
          DUMMY204 := aux_iv_op ;
          DUMMY205 := aux_cipher_op ;
          DUMMY207 := DUMMY205 ;
          DUMMY206 := not(((boolean_to_std(DUMMY207 = AES_GCM) or boolean_to_std
          (DUMMY207 = AES_XTS_XEX)) or boolean_to_std(DUMMY207 = AES_GMAC))) ;
          _zyL254_tfiRv55_DUMMY12 := boolean_to_std(((DUMMY203 = AUX_CMD or
           DUMMY203 = AUX_CMD_GUID) and DUMMY204 = IV_INC and (not(DUMMY206)
          )='1')) ;
          nxt_kme_internal_dek_kim_word(19 downto 19) <= ext
          (_zyL254_tfiRv55_DUMMY12,1) ;
          DUMMY208 := always_validate_kim_ref ;
          DUMMY209 := aux_key_type ;
          DUMMY210 := aux_auth_op ;
          DUMMY211 := aux_raw_auth_op ;
          _zyL255_tfiRv56_DUMMY13 := '1' ;
          if ((DUMMY208 = '0')) then

            case DUMMY209 is
              when  "000000"  =>
                _zyL255_tfiRv56_DUMMY13 := '0' ;
              when  "000001"  =>
                DUMMY215 := DUMMY210 ;
                DUMMY216 := DUMMY211 ;
                DUMMY212 := (boolean_to_std(DUMMY215 /= HMAC_SHA2) and
                 boolean_to_std(DUMMY216 /= HMAC_SHA2)) ;
                if (DUMMY212 = '1') then
                  _zyL255_tfiRv56_DUMMY13 := '0' ;
                end if;
              when  "000111"  =>
                DUMMY217 := DUMMY210 ;
                DUMMY218 := DUMMY211 ;
                DUMMY213 := (boolean_to_std(DUMMY217 /= HMAC_SHA2) and
                 boolean_to_std(DUMMY218 /= HMAC_SHA2)) ;
                if (DUMMY213 = '1') then
                  _zyL255_tfiRv56_DUMMY13 := '0' ;
                end if;
              when  "001000"  =>
                DUMMY219 := DUMMY210 ;
                DUMMY220 := DUMMY211 ;
                DUMMY214 := (boolean_to_std(DUMMY219 /= HMAC_SHA2) and
                 boolean_to_std(DUMMY220 /= HMAC_SHA2)) ;
                if (DUMMY214 = '1') then
                  _zyL255_tfiRv56_DUMMY13 := '0' ;
                end if;
              when others => null ;
            end case;
          end if;
          nxt_kme_internal_dak_kim_word(17 downto 17) <= ext
          (_zyL255_tfiRv56_DUMMY13,1) ;
        end if;
      end if;
    end if;
    if (stitcher_rd_DUMMY8 = '1') then
      if (key_blob_region = '1') then

        case aux_key_type is
          when  "000010"  |  "000011"  |  "000100"  =>
            fifo_in_valid <= '1' ;
            DUMMY221 := std_logic_vector'(stitcher_out(31 downto 0) & DUMMY7) ;
            _zyL288_tfiRv57_DUMMY14 := std_logic_vector'(DUMMY221(7 downto 0) &
             DUMMY221(15 downto 8) & DUMMY221(23 downto 16) & DUMMY221(31 downto
             24) & DUMMY221(39 downto 32) & DUMMY221(47 downto 40) & DUMMY221(55
             downto 48) & DUMMY221(63 downto 56)) ;
            fifo_in_DUMMY0(63 downto 0) := _zyL288_tfiRv57_DUMMY14 ;
            nxt_buffer_DUMMY3 := stitcher_out(63 downto 32) ;
            if (stitcher_eot = '1') then
              DUMMY222 := std_logic_vector'(stitcher_out(31 downto 0) & DUMMY7)
               ;
              _zyL293_tfiRv58_DUMMY15 := std_logic_vector'(DUMMY222(7 downto 0)
               & DUMMY222(15 downto 8) & DUMMY222(23 downto 16) & DUMMY222(31
               downto 24) & DUMMY222(39 downto 32) & DUMMY222(47 downto 40) &
               DUMMY222(55 downto 48) & DUMMY222(63 downto 56)) ;
              fifo_in_DUMMY0(63 downto 0) := _zyL293_tfiRv58_DUMMY15 ;
              nxt_skip(6 downto 6) <= "1" ;
              nxt_skip(3 downto 0) <= KME_WORD0 ;
            end if;
          when  "000101"  |  "000110"  =>
            fifo_in_valid <= '1' ;
            DUMMY223 := std_logic_vector'(stitcher_out(31 downto 0) & DUMMY7) ;
            _zyL301_tfiRv59_DUMMY16 := std_logic_vector'(DUMMY223(7 downto 0) &
             DUMMY223(15 downto 8) & DUMMY223(23 downto 16) & DUMMY223(31 downto
             24) & DUMMY223(39 downto 32) & DUMMY223(47 downto 40) & DUMMY223(55
             downto 48) & DUMMY223(63 downto 56)) ;
            fifo_in_DUMMY0(63 downto 0) := _zyL301_tfiRv59_DUMMY16 ;
            nxt_buffer_DUMMY3 := stitcher_out(63 downto 32) ;
            if (ext(int_tlv_counter,32) = std_logic_vector'
            ("00000000000000000000000000011111")) then
              DUMMY224 := std_logic_vector'(stitcher_out(31 downto 0) & DUMMY7)
               ;
              _zyL306_tfiRv60_DUMMY17 := std_logic_vector'(DUMMY224(7 downto 0)
               & DUMMY224(15 downto 8) & DUMMY224(23 downto 16) & DUMMY224(31
               downto 24) & DUMMY224(39 downto 32) & DUMMY224(47 downto 40) &
               DUMMY224(55 downto 48) & DUMMY224(63 downto 56)) ;
              fifo_in_DUMMY0(63 downto 0) := _zyL306_tfiRv60_DUMMY17 ;
              nxt_skip(6 downto 6) <= "1" ;
              nxt_skip(3 downto 0) <= KME_DAK ;
            end if;
            if (stitcher_eot = '1') then
              DUMMY225 := std_logic_vector'(stitcher_out(31 downto 0) & DUMMY7)
               ;
              _zyL313_tfiRv61_DUMMY18 := std_logic_vector'(DUMMY225(7 downto 0)
               & DUMMY225(15 downto 8) & DUMMY225(23 downto 16) & DUMMY225(31
               downto 24) & DUMMY225(39 downto 32) & DUMMY225(47 downto 40) &
               DUMMY225(55 downto 48) & DUMMY225(63 downto 56)) ;
              fifo_in_DUMMY0(63 downto 0) := _zyL313_tfiRv61_DUMMY18 ;
              nxt_skip(6 downto 6) <= "1" ;
              nxt_skip(3 downto 0) <= KME_WORD0 ;
            end if;
          when  "000111"  |  "001000"  |  "001001"  =>
            fifo_in_valid <= '1' ;
            DUMMY226 := stitcher_out(63 downto 0) ;
            _zyL321_tfiRv62_DUMMY19 := std_logic_vector'(DUMMY226(7 downto 0) &
             DUMMY226(15 downto 8) & DUMMY226(23 downto 16) & DUMMY226(31 downto
             24) & DUMMY226(39 downto 32) & DUMMY226(47 downto 40) & DUMMY226(55
             downto 48) & DUMMY226(63 downto 56)) ;
            fifo_in_DUMMY0(63 downto 0) := _zyL321_tfiRv62_DUMMY19 ;
            nxt_buffer_DUMMY3 := stitcher_out(63 downto 32) ;
            if (int_tlv_counter = IDX_KME_EIV) then
              DUMMY227 := std_logic_vector'(stitcher_out(31 downto 0) & DUMMY7)
               ;
              _zyL327_tfiRv63_DUMMY20 := std_logic_vector'(DUMMY227(7 downto 0)
               & DUMMY227(15 downto 8) & DUMMY227(23 downto 16) & DUMMY227(31
               downto 24) & DUMMY227(39 downto 32) & DUMMY227(47 downto 40) &
               DUMMY227(55 downto 48) & DUMMY227(63 downto 56)) ;
              fifo_in_DUMMY0(63 downto 0) := _zyL327_tfiRv63_DUMMY20 ;
              nxt_skip(6 downto 6) <= "1" ;
              nxt_skip(5 downto 5) <= "1" ;
              nxt_skip(4 downto 4) <= "1" ;
              nxt_skip(3 downto 0) <= it_cond_op(aux_key_type =
               ENC_DEK256,KME_DEK1,KME_DEK0) ;
            end if;
            if (int_tlv_counter = IDX_KME_AIV) then
              DUMMY228 := std_logic_vector'(stitcher_out(31 downto 0) & DUMMY7)
               ;
              _zyL337_tfiRv64_DUMMY21 := std_logic_vector'(DUMMY228(7 downto 0)
               & DUMMY228(15 downto 8) & DUMMY228(23 downto 16) & DUMMY228(31
               downto 24) & DUMMY228(39 downto 32) & DUMMY228(47 downto 40) &
               DUMMY228(55 downto 48) & DUMMY228(63 downto 56)) ;
              fifo_in_DUMMY0(63 downto 0) := _zyL337_tfiRv64_DUMMY21 ;
              nxt_skip(6 downto 6) <= "1" ;
              nxt_skip(5 downto 5) <= "1" ;
              nxt_skip(4 downto 4) <= "1" ;
              nxt_skip(3 downto 0) <= KME_DAK ;
            end if;
            if (stitcher_eot = '1') then
              DUMMY229 := std_logic_vector'(std_logic_vector'
              ("00000000000000000000000000000000") & stitcher_out(31 downto 0))
               ;
              _zyL346_tfiRv65_DUMMY22 := std_logic_vector'(DUMMY229(7 downto 0)
               & DUMMY229(15 downto 8) & DUMMY229(23 downto 16) & DUMMY229(31
               downto 24) & DUMMY229(39 downto 32) & DUMMY229(47 downto 40) &
               DUMMY229(55 downto 48) & DUMMY229(63 downto 56)) ;
              fifo_in_DUMMY0(63 downto 0) := _zyL346_tfiRv65_DUMMY22 ;
              nxt_skip(6 downto 6) <= "1" ;
              nxt_skip(3 downto 0) <= KME_WORD0 ;
            end if;
          when  "001010"  |  "001011"  =>
            fifo_in_valid <= '1' ;
            DUMMY230 := stitcher_out(63 downto 0) ;
            _zyL354_tfiRv66_DUMMY23 := std_logic_vector'(DUMMY230(7 downto 0) &
             DUMMY230(15 downto 8) & DUMMY230(23 downto 16) & DUMMY230(31 downto
             24) & DUMMY230(39 downto 32) & DUMMY230(47 downto 40) & DUMMY230(55
             downto 48) & DUMMY230(63 downto 56)) ;
            fifo_in_DUMMY0(63 downto 0) := _zyL354_tfiRv66_DUMMY23 ;
            nxt_buffer_DUMMY3 := stitcher_out(63 downto 32) ;
            if (int_tlv_counter = IDX_KME_EIV) then
              DUMMY231 := std_logic_vector'(stitcher_out(31 downto 0) & DUMMY7)
               ;
              _zyL359_tfiRv67_DUMMY24 := std_logic_vector'(DUMMY231(7 downto 0)
               & DUMMY231(15 downto 8) & DUMMY231(23 downto 16) & DUMMY231(31
               downto 24) & DUMMY231(39 downto 32) & DUMMY231(47 downto 40) &
               DUMMY231(55 downto 48) & DUMMY231(63 downto 56)) ;
              fifo_in_DUMMY0(63 downto 0) := _zyL359_tfiRv67_DUMMY24 ;
              nxt_skip(6 downto 6) <= "1" ;
              nxt_skip(5 downto 5) <= "1" ;
              nxt_skip(4 downto 4) <= "1" ;
              nxt_skip(3 downto 0) <= it_cond_op(aux_key_type =
               ENC_DEK256_DAK,KME_DEK1,KME_DEK0) ;
            end if;
            if (ext(int_tlv_counter,32) = std_logic_vector'
            ("00000000000000000000000000100001")) then
              DUMMY232 := std_logic_vector'(std_logic_vector'
              ("00000000000000000000000000000000") & stitcher_out(31 downto 0))
               ;
              _zyL368_tfiRv68_DUMMY25 := std_logic_vector'(DUMMY232(7 downto 0)
               & DUMMY232(15 downto 8) & DUMMY232(23 downto 16) & DUMMY232(31
               downto 24) & DUMMY232(39 downto 32) & DUMMY232(47 downto 40) &
               DUMMY232(55 downto 48) & DUMMY232(63 downto 56)) ;
              fifo_in_DUMMY0(63 downto 0) := _zyL368_tfiRv68_DUMMY25 ;
            end if;
            if (int_tlv_counter = IDX_KME_AIV) then
              DUMMY233 := std_logic_vector'(stitcher_out(31 downto 0) & DUMMY7)
               ;
              _zyL373_tfiRv69_DUMMY26 := std_logic_vector'(DUMMY233(7 downto 0)
               & DUMMY233(15 downto 8) & DUMMY233(23 downto 16) & DUMMY233(31
               downto 24) & DUMMY233(39 downto 32) & DUMMY233(47 downto 40) &
               DUMMY233(55 downto 48) & DUMMY233(63 downto 56)) ;
              fifo_in_DUMMY0(63 downto 0) := _zyL373_tfiRv69_DUMMY26 ;
              nxt_skip(6 downto 6) <= "1" ;
              nxt_skip(5 downto 5) <= "1" ;
              nxt_skip(4 downto 4) <= "1" ;
              nxt_skip(3 downto 0) <= KME_DAK ;
            end if;
            if (stitcher_eot = '1') then
              DUMMY234 := std_logic_vector'(std_logic_vector'
              ("00000000000000000000000000000000") & stitcher_out(31 downto 0))
               ;
              _zyL382_tfiRv70_DUMMY27 := std_logic_vector'(DUMMY234(7 downto 0)
               & DUMMY234(15 downto 8) & DUMMY234(23 downto 16) & DUMMY234(31
               downto 24) & DUMMY234(39 downto 32) & DUMMY234(47 downto 40) &
               DUMMY234(55 downto 48) & DUMMY234(63 downto 56)) ;
              fifo_in_DUMMY0(63 downto 0) := _zyL382_tfiRv70_DUMMY27 ;
              nxt_skip(6 downto 6) <= "1" ;
              nxt_skip(3 downto 0) <= KME_WORD0 ;
            end if;
          when  "001100"  |  "001101"  =>
            fifo_in_valid <= '1' ;
            DUMMY235 := stitcher_out(63 downto 0) ;
            _zyL390_tfiRv71_DUMMY28 := std_logic_vector'(DUMMY235(7 downto 0) &
             DUMMY235(15 downto 8) & DUMMY235(23 downto 16) & DUMMY235(31 downto
             24) & DUMMY235(39 downto 32) & DUMMY235(47 downto 40) & DUMMY235(55
             downto 48) & DUMMY235(63 downto 56)) ;
            fifo_in_DUMMY0(63 downto 0) := _zyL390_tfiRv71_DUMMY28 ;
            nxt_buffer_DUMMY3 := stitcher_out(63 downto 32) ;
            if (int_tlv_counter = IDX_KME_EIV) then
              DUMMY236 := std_logic_vector'(stitcher_out(31 downto 0) & DUMMY7)
               ;
              _zyL395_tfiRv72_DUMMY29 := std_logic_vector'(DUMMY236(7 downto 0)
               & DUMMY236(15 downto 8) & DUMMY236(23 downto 16) & DUMMY236(31
               downto 24) & DUMMY236(39 downto 32) & DUMMY236(47 downto 40) &
               DUMMY236(55 downto 48) & DUMMY236(63 downto 56)) ;
              fifo_in_DUMMY0(63 downto 0) := _zyL395_tfiRv72_DUMMY29 ;
              nxt_skip(6 downto 6) <= "1" ;
              nxt_skip(5 downto 5) <= "1" ;
              nxt_skip(4 downto 4) <= "1" ;
              nxt_skip(3 downto 0) <= it_cond_op(aux_key_type =
               ENC_DEK256_DAK_COMB,KME_DEK1,KME_DEK0) ;
            end if;
            if (ext(int_tlv_counter,32) = std_logic_vector'
            ("00000000000000000000000000011111")) then
              nxt_skip(6 downto 6) <= "1" ;
              nxt_skip(3 downto 0) <= KME_DAK ;
            end if;
            if (stitcher_eot = '1') then
              DUMMY237 := std_logic_vector'(std_logic_vector'
              ("00000000000000000000000000000000") & stitcher_out(31 downto 0))
               ;
              _zyL410_tfiRv73_DUMMY30 := std_logic_vector'(DUMMY237(7 downto 0)
               & DUMMY237(15 downto 8) & DUMMY237(23 downto 16) & DUMMY237(31
               downto 24) & DUMMY237(39 downto 32) & DUMMY237(47 downto 40) &
               DUMMY237(55 downto 48) & DUMMY237(63 downto 56)) ;
              fifo_in_DUMMY0(63 downto 0) := _zyL410_tfiRv73_DUMMY30 ;
              nxt_skip(6 downto 6) <= "1" ;
              nxt_skip(3 downto 0) <= KME_WORD0 ;
            end if;
          when others => null ;
        end case;
      else

        case tlv_counter is
          when  "00000"  =>
            nxt_kme_internal_word0_DUMMY1 :=
             "0000000000000000000000000000000000000000000000000000000000000000"
             ;
            nxt_kme_internal_word0_DUMMY1(7 downto 0) := tlv_word0_DUMMY4(7
             downto 0) ;
            nxt_kme_internal_word0_DUMMY1(24+3 downto 24) := tlv_word0_DUMMY4
            (24+3 downto 24) ;
            nxt_kme_internal_word0_DUMMY1(16+7 downto 16) := tlv_word0_DUMMY4
            (16+7 downto 16) ;
            nxt_kme_internal_word0_DUMMY1(28+10 downto 28) := tlv_word0_DUMMY4
            (32+10 downto 32) ;
            nxt_tlv_type <= tlv_word0_DUMMY4(7 downto 0) ;
            if (tlv_word0_DUMMY4(7 downto 0) = RQE) then
              nxt_kme_internal_dek_kim_word <=
               "0000000000000000000000000000000000000000000000000000000000000000"
               ;
              nxt_kme_internal_dak_kim_word <=
               "0000000000000000000000000000000000000000000000000000000000000000"
               ;
              nxt_kme_internal_dek_kim_word(16 downto 16) <= ext
              (tlv_word0_DUMMY4(55),1) ;
              nxt_kme_internal_dak_kim_word(16 downto 16) <= ext
              (tlv_word0_DUMMY4(55),1) ;
            end if;
            nxt_aux_key_type <= NO_AUX_KEY ;
            nxt_aux_iv_op <= IV_SRC ;
            nxt_aux_cipher_op <= CPH_NULL ;
            nxt_aux_auth_op <= AUTH_NULL ;
            nxt_aux_raw_auth_op <= AUTH_NULL ;
            nxt_aux_key_header_DUMMY2 := "00000000000000000000000000000000" ;
            nxt_iv0 <=
             "0000000000000000000000000000000000000000000000000000000000000000"
             ;
            nxt_iv1 <=
             "0000000000000000000000000000000000000000000000000000000000000000"
             ;
            nxt_guid0 <=
             "0000000000000000000000000000000000000000000000000000000000000000"
             ;
            nxt_guid1 <=
             "0000000000000000000000000000000000000000000000000000000000000000"
             ;
            nxt_guid2 <=
             "0000000000000000000000000000000000000000000000000000000000000000"
             ;
            nxt_guid3 <=
             "0000000000000000000000000000000000000000000000000000000000000000"
             ;
          when  "00001"  =>
            if (tlv_type = RQE) then
              nxt_kme_internal_dek_kim_word(12+3 downto 12) <= tlv_word1_DUMMY5
              (60+3 downto 60) ;
              nxt_kme_internal_dek_kim_word(11 downto 0) <= tlv_word1_DUMMY5
              (48+11 downto 48) ;
              nxt_kme_internal_dak_kim_word(12+3 downto 12) <= tlv_word1_DUMMY5
              (60+3 downto 60) ;
              nxt_kme_internal_dak_kim_word(11 downto 0) <= tlv_word1_DUMMY5
              (48+11 downto 48) ;
            else

              case tlv_type is
                when  "00010101"  =>
                  if (frame_word_DUMMY7(4 downto 4) = GUID_PRESENT) then
                    nxt_tlv_type <= AUX_CMD_GUID ;
                  end if;
                when  "00010111"  =>
                  if (frame_word_DUMMY7(4 downto 4) = GUID_PRESENT) then
                    nxt_tlv_type <= AUX_CMD_GUID_IV ;
                  end if;
                when others => null ;
              end case;
              if (disable_debug_cmd_q = '1') then
                nxt_debug_cmd <= "00000000000000000000000000000000" ;
              else
                nxt_debug_cmd <= stitcher_out(63 downto 32) ;
              end if;
            end if;
          when  "00010"  =>
            nxt_kme_internal_word0_DUMMY1(39+5 downto 39) := tlv_word2_DUMMY6
            (57+5 downto 57) ;
            DUMMY238 := always_validate_kim_ref ;
            DUMMY239 := tlv_word2_DUMMY6(57+5 downto 57) ;
            DUMMY240 := tlv_word2_DUMMY6(40+3 downto 40) ;
            _zyL485_tfiRv74_DUMMY31 := '1' ;
            if ((DUMMY238 = '0')) then

              case DUMMY239 is
                when  "000000"  =>
                  _zyL485_tfiRv74_DUMMY31 := '0' ;
                when  "000001"  =>
                  DUMMY243 := DUMMY240 ;
                  DUMMY241 := not(((boolean_to_std(DUMMY243 = AES_GCM) or
                   boolean_to_std(DUMMY243 = AES_XTS_XEX)) or boolean_to_std
                  (DUMMY243 = AES_GMAC))) ;
                  if (DUMMY241 = '1') then
                    _zyL485_tfiRv74_DUMMY31 := '0' ;
                  end if;
                when  "001001"  =>
                  DUMMY244 := DUMMY240 ;
                  DUMMY242 := not(((boolean_to_std(DUMMY244 = AES_GCM) or
                   boolean_to_std(DUMMY244 = AES_XTS_XEX)) or boolean_to_std
                  (DUMMY244 = AES_GMAC))) ;
                  if (DUMMY242 = '1') then
                    _zyL485_tfiRv74_DUMMY31 := '0' ;
                  end if;
                when others => null ;
              end case;
            end if;
            nxt_kme_internal_word0_DUMMY1(46 downto 46) := ext
            (_zyL485_tfiRv74_DUMMY31,1) ;
            DUMMY245 := always_validate_kim_ref ;
            DUMMY246 := tlv_word2_DUMMY6(57+5 downto 57) ;
            DUMMY247 := tlv_word2_DUMMY6(36+3 downto 36) ;
            DUMMY248 := tlv_word2_DUMMY6(32+3 downto 32) ;
            _zyL486_tfiRv75_DUMMY32 := '1' ;
            if ((DUMMY245 = '0')) then

              case DUMMY246 is
                when  "000000"  =>
                  _zyL486_tfiRv75_DUMMY32 := '0' ;
                when  "000001"  =>
                  DUMMY252 := DUMMY247 ;
                  DUMMY253 := DUMMY248 ;
                  DUMMY249 := (boolean_to_std(DUMMY252 /= HMAC_SHA2) and
                   boolean_to_std(DUMMY253 /= HMAC_SHA2)) ;
                  if (DUMMY249 = '1') then
                    _zyL486_tfiRv75_DUMMY32 := '0' ;
                  end if;
                when  "000111"  =>
                  DUMMY254 := DUMMY247 ;
                  DUMMY255 := DUMMY248 ;
                  DUMMY250 := (boolean_to_std(DUMMY254 /= HMAC_SHA2) and
                   boolean_to_std(DUMMY255 /= HMAC_SHA2)) ;
                  if (DUMMY250 = '1') then
                    _zyL486_tfiRv75_DUMMY32 := '0' ;
                  end if;
                when  "001000"  =>
                  DUMMY256 := DUMMY247 ;
                  DUMMY257 := DUMMY248 ;
                  DUMMY251 := (boolean_to_std(DUMMY256 /= HMAC_SHA2) and
                   boolean_to_std(DUMMY257 /= HMAC_SHA2)) ;
                  if (DUMMY251 = '1') then
                    _zyL486_tfiRv75_DUMMY32 := '0' ;
                  end if;
                when others => null ;
              end case;
            end if;
            nxt_kme_internal_word0_DUMMY1(45 downto 45) := ext
            (_zyL486_tfiRv75_DUMMY32,1) ;
            DUMMY258 := tlv_word2_DUMMY6(40+3 downto 40) ;
            _zyL489_tfiRv76_DUMMY33 := not(((boolean_to_std(DUMMY258 = AES_GCM)
             or boolean_to_std(DUMMY258 = AES_XTS_XEX)) or boolean_to_std
            (DUMMY258 = AES_GMAC))) ;
            DUMMY259 := tlv_word2_DUMMY6(36+3 downto 36) ;
            DUMMY260 := tlv_word2_DUMMY6(32+3 downto 32) ;
            _zyL489_tfiRv77_DUMMY34 := (boolean_to_std(DUMMY259 /= HMAC_SHA2)
             and boolean_to_std(DUMMY260 /= HMAC_SHA2)) ;
            nxt_kme_internal_word0_DUMMY1(47 downto 47) := (ext
            (_zyL489_tfiRv76_DUMMY33,1) and ext(_zyL489_tfiRv77_DUMMY34,1)) ;
            DUMMY261 := tlv_word2_DUMMY6(40+3 downto 40) ;
            _zyL492_tfiRv78_DUMMY35 := it_cond_op(DUMMY261 =
             AES_XTS_XEX,std_logic'('1'),std_logic'('0')) ;
            nxt_kme_internal_word0_DUMMY1(48 downto 48) := ext
            (_zyL492_tfiRv78_DUMMY35,1) ;
            nxt_aux_key_type <= tlv_word2_DUMMY6(57+5 downto 57) ;
            nxt_aux_iv_op <= tlv_word2_DUMMY6(52+1 downto 52) ;
            nxt_aux_cipher_op <= tlv_word2_DUMMY6(40+3 downto 40) ;
            nxt_aux_auth_op <= tlv_word2_DUMMY6(36+3 downto 36) ;
            nxt_aux_raw_auth_op <= tlv_word2_DUMMY6(32+3 downto 32) ;
            fifo_in_valid <= '1' ;
            fifo_in_DUMMY0(63 downto 0) := nxt_kme_internal_word0_DUMMY1 ;
            if (stitcher_eot = '1') then
              nxt_buffer_DUMMY3 := debug_cmd ;
              nxt_skip(6 downto 6) <= "1" ;
              nxt_skip(5 downto 5) <= "1" ;
            end if;
          when  "00011"  =>

            case tlv_type is
              when  "00011000"  =>
                DUMMY262 := stitcher_out(63 downto 0) ;
                _zyL526_tfiRv79_DUMMY36 := std_logic_vector'(DUMMY262(7 downto 0
                ) & DUMMY262(15 downto 8) & DUMMY262(23 downto 16) & DUMMY262(31
                 downto 24) & DUMMY262(39 downto 32) & DUMMY262(47 downto 40) &
                 DUMMY262(55 downto 48) & DUMMY262(63 downto 56)) ;
                nxt_guid0 <= _zyL526_tfiRv79_DUMMY36 ;
              when  "00011001"  =>
                DUMMY263 := stitcher_out(63 downto 0) ;
                _zyL527_tfiRv80_DUMMY37 := std_logic_vector'(DUMMY263(7 downto 0
                ) & DUMMY263(15 downto 8) & DUMMY263(23 downto 16) & DUMMY263(31
                 downto 24) & DUMMY263(39 downto 32) & DUMMY263(47 downto 40) &
                 DUMMY263(55 downto 48) & DUMMY263(63 downto 56)) ;
                nxt_guid0 <= _zyL527_tfiRv80_DUMMY37 ;
              when  "00010111"  =>
                nxt_iv0 <= stitcher_out(63 downto 0) ;
              when others => null ;
            end case;
            if (tlv_type = AUX_CMD) then
              DUMMY264 := stitcher_out(63 downto 0) ;
              nxt_aux_key_header_DUMMY2 := DUMMY264(33 to 64) ;
              nxt_buffer_DUMMY3 := DUMMY264(1 to 32) ;
              fifo_in_valid <= '1' ;
              fifo_in_DUMMY0(63 downto 0) := std_logic_vector'(debug_cmd &
               nxt_aux_key_header_DUMMY2) ;
              nxt_skip(6 downto 6) <= "1" ;
            end if;
          when  "00100"  =>

            case tlv_type is
              when  "00011000"  =>
                DUMMY265 := stitcher_out(63 downto 0) ;
                _zyL541_tfiRv81_DUMMY38 := std_logic_vector'(DUMMY265(7 downto 0
                ) & DUMMY265(15 downto 8) & DUMMY265(23 downto 16) & DUMMY265(31
                 downto 24) & DUMMY265(39 downto 32) & DUMMY265(47 downto 40) &
                 DUMMY265(55 downto 48) & DUMMY265(63 downto 56)) ;
                nxt_guid1 <= _zyL541_tfiRv81_DUMMY38 ;
              when  "00011001"  =>
                DUMMY266 := stitcher_out(63 downto 0) ;
                _zyL542_tfiRv82_DUMMY39 := std_logic_vector'(DUMMY266(7 downto 0
                ) & DUMMY266(15 downto 8) & DUMMY266(23 downto 16) & DUMMY266(31
                 downto 24) & DUMMY266(39 downto 32) & DUMMY266(47 downto 40) &
                 DUMMY266(55 downto 48) & DUMMY266(63 downto 56)) ;
                nxt_guid1 <= _zyL542_tfiRv82_DUMMY39 ;
              when  "00010111"  =>
                nxt_iv1 <= stitcher_out(63 downto 0) ;
              when others => null ;
            end case;
            if (stitcher_eot = '1') then
              nxt_buffer_DUMMY3 := debug_cmd ;
              nxt_skip(6 downto 6) <= "1" ;
              nxt_skip(5 downto 5) <= "1" ;
            end if;
          when  "00101"  =>

            case tlv_type is
              when  "00011000"  =>
                DUMMY267 := stitcher_out(63 downto 0) ;
                _zyL555_tfiRv83_DUMMY40 := std_logic_vector'(DUMMY267(7 downto 0
                ) & DUMMY267(15 downto 8) & DUMMY267(23 downto 16) & DUMMY267(31
                 downto 24) & DUMMY267(39 downto 32) & DUMMY267(47 downto 40) &
                 DUMMY267(55 downto 48) & DUMMY267(63 downto 56)) ;
                nxt_guid2 <= _zyL555_tfiRv83_DUMMY40 ;
              when  "00011001"  =>
                DUMMY268 := stitcher_out(63 downto 0) ;
                _zyL556_tfiRv84_DUMMY41 := std_logic_vector'(DUMMY268(7 downto 0
                ) & DUMMY268(15 downto 8) & DUMMY268(23 downto 16) & DUMMY268(31
                 downto 24) & DUMMY268(39 downto 32) & DUMMY268(47 downto 40) &
                 DUMMY268(55 downto 48) & DUMMY268(63 downto 56)) ;
                nxt_guid2 <= _zyL556_tfiRv84_DUMMY41 ;
              when others => null ;
            end case;
            if (tlv_type = AUX_CMD_IV) then
              DUMMY269 := stitcher_out(63 downto 0) ;
              nxt_aux_key_header_DUMMY2 := DUMMY269(33 to 64) ;
              nxt_buffer_DUMMY3 := DUMMY269(1 to 32) ;
              fifo_in_valid <= '1' ;
              fifo_in_DUMMY0(63 downto 0) := std_logic_vector'(debug_cmd &
               nxt_aux_key_header_DUMMY2) ;
              nxt_skip(6 downto 6) <= "1" ;
            end if;
          when  "00110"  =>

            case tlv_type is
              when  "00011000"  =>
                DUMMY270 := stitcher_out(63 downto 0) ;
                _zyL569_tfiRv85_DUMMY42 := std_logic_vector'(DUMMY270(7 downto 0
                ) & DUMMY270(15 downto 8) & DUMMY270(23 downto 16) & DUMMY270(31
                 downto 24) & DUMMY270(39 downto 32) & DUMMY270(47 downto 40) &
                 DUMMY270(55 downto 48) & DUMMY270(63 downto 56)) ;
                nxt_guid3 <= _zyL569_tfiRv85_DUMMY42 ;
              when  "00011001"  =>
                DUMMY271 := stitcher_out(63 downto 0) ;
                _zyL570_tfiRv86_DUMMY43 := std_logic_vector'(DUMMY271(7 downto 0
                ) & DUMMY271(15 downto 8) & DUMMY271(23 downto 16) & DUMMY271(31
                 downto 24) & DUMMY271(39 downto 32) & DUMMY271(47 downto 40) &
                 DUMMY271(55 downto 48) & DUMMY271(63 downto 56)) ;
                nxt_guid3 <= _zyL570_tfiRv86_DUMMY43 ;
              when others => null ;
            end case;
            if (stitcher_eot = '1') then
              nxt_buffer_DUMMY3 := debug_cmd ;
              nxt_skip(6 downto 6) <= "1" ;
              nxt_skip(5 downto 5) <= "1" ;
            end if;
          when  "00111"  =>

            case tlv_type is
              when  "00011001"  =>
                nxt_iv0 <= stitcher_out(63 downto 0) ;
              when others => null ;
            end case;
            if (tlv_type = AUX_CMD_GUID) then
              DUMMY272 := stitcher_out(63 downto 0) ;
              nxt_aux_key_header_DUMMY2 := DUMMY272(33 to 64) ;
              nxt_buffer_DUMMY3 := DUMMY272(1 to 32) ;
              fifo_in_valid <= '1' ;
              fifo_in_DUMMY0(63 downto 0) := std_logic_vector'(debug_cmd &
               nxt_aux_key_header_DUMMY2) ;
              nxt_skip(6 downto 6) <= "1" ;
            end if;
          when  "01000"  =>

            case tlv_type is
              when  "00011001"  =>
                nxt_iv1 <= stitcher_out(63 downto 0) ;
              when others => null ;
            end case;
            if (stitcher_eot = '1') then
              nxt_buffer_DUMMY3 := debug_cmd ;
              nxt_skip(6 downto 6) <= "1" ;
              nxt_skip(5 downto 5) <= "1" ;
            end if;
          when  "01001"  =>
            DUMMY273 := stitcher_out(63 downto 0) ;
            nxt_aux_key_header_DUMMY2 := DUMMY273(33 to 64) ;
            nxt_buffer_DUMMY3 := DUMMY273(1 to 32) ;
            fifo_in_valid <= '1' ;
            fifo_in_DUMMY0(63 downto 0) := std_logic_vector'(debug_cmd &
             nxt_aux_key_header_DUMMY2) ;
            nxt_skip(6 downto 6) <= "1" ;
          when others => null ;
        end case;

        case aux_key_type is
          when  "000000"  =>
            nxt_skip(3 downto 0) <= KME_WORD0 ;
          when  "000001"  =>
            nxt_skip(3 downto 0) <= KME_WORD0 ;
          when  "000010"  =>
            nxt_skip(3 downto 0) <= KME_DEK1 ;
          when  "000011"  =>
            nxt_skip(3 downto 0) <= KME_DEK0 ;
          when  "000100"  =>
            nxt_skip(3 downto 0) <= KME_DAK ;
          when  "000101"  =>
            nxt_skip(3 downto 0) <= KME_DEK1 ;
          when  "000110"  =>
            nxt_skip(3 downto 0) <= KME_DEK0 ;
          when  "000111"  =>
            nxt_skip(3 downto 0) <= KME_EIV ;
          when  "001000"  =>
            nxt_skip(3 downto 0) <= KME_EIV ;
          when  "001001"  =>
            nxt_skip(3 downto 0) <= KME_AIV ;
          when  "001010"  =>
            nxt_skip(3 downto 0) <= KME_EIV ;
          when  "001011"  =>
            nxt_skip(3 downto 0) <= KME_EIV ;
          when  "001100"  =>
            nxt_skip(3 downto 0) <= KME_EIV ;
          when  "001101"  =>
            nxt_skip(3 downto 0) <= KME_EIV ;
          when others => null ;
        end case;
      end if;
    end if;
    fifo_in <= transport fifo_in_DUMMY0;
    nxt_kme_internal_word0 <= nxt_kme_internal_word0_DUMMY1;
    nxt_aux_key_header <= nxt_aux_key_header_DUMMY2;
    nxt_buffer <= nxt_buffer_DUMMY3;
    tlv_word0 <= tlv_word0_DUMMY4;
    tlv_word1 <= tlv_word1_DUMMY5;
    tlv_word2 <= tlv_word2_DUMMY6;
    frame_word <= frame_word_DUMMY7;
    stitcher_rd <= stitcher_rd_DUMMY8;
    _zyL234_tfiRv52 <= _zyL234_tfiRv52_DUMMY9;
    _zyL252_tfiRv53 <= _zyL252_tfiRv53_DUMMY10;
    _zyL253_tfiRv54 <= _zyL253_tfiRv54_DUMMY11;
    _zyL254_tfiRv55 <= _zyL254_tfiRv55_DUMMY12;
    _zyL255_tfiRv56 <= _zyL255_tfiRv56_DUMMY13;
    _zyL288_tfiRv57 <= _zyL288_tfiRv57_DUMMY14;
    _zyL293_tfiRv58 <= _zyL293_tfiRv58_DUMMY15;
    _zyL301_tfiRv59 <= _zyL301_tfiRv59_DUMMY16;
    _zyL306_tfiRv60 <= _zyL306_tfiRv60_DUMMY17;
    _zyL313_tfiRv61 <= _zyL313_tfiRv61_DUMMY18;
    _zyL321_tfiRv62 <= _zyL321_tfiRv62_DUMMY19;
    _zyL327_tfiRv63 <= _zyL327_tfiRv63_DUMMY20;
    _zyL337_tfiRv64 <= _zyL337_tfiRv64_DUMMY21;
    _zyL346_tfiRv65 <= _zyL346_tfiRv65_DUMMY22;
    _zyL354_tfiRv66 <= _zyL354_tfiRv66_DUMMY23;
    _zyL359_tfiRv67 <= _zyL359_tfiRv67_DUMMY24;
    _zyL368_tfiRv68 <= _zyL368_tfiRv68_DUMMY25;
    _zyL373_tfiRv69 <= _zyL373_tfiRv69_DUMMY26;
    _zyL382_tfiRv70 <= _zyL382_tfiRv70_DUMMY27;
    _zyL390_tfiRv71 <= _zyL390_tfiRv71_DUMMY28;
    _zyL395_tfiRv72 <= _zyL395_tfiRv72_DUMMY29;
    _zyL410_tfiRv73 <= _zyL410_tfiRv73_DUMMY30;
    _zyL485_tfiRv74 <= _zyL485_tfiRv74_DUMMY31;
    _zyL486_tfiRv75 <= _zyL486_tfiRv75_DUMMY32;
    _zyL489_tfiRv76 <= _zyL489_tfiRv76_DUMMY33;
    _zyL489_tfiRv77 <= _zyL489_tfiRv77_DUMMY34;
    _zyL492_tfiRv78 <= _zyL492_tfiRv78_DUMMY35;
    _zyL526_tfiRv79 <= _zyL526_tfiRv79_DUMMY36;
    _zyL527_tfiRv80 <= _zyL527_tfiRv80_DUMMY37;
    _zyL541_tfiRv81 <= _zyL541_tfiRv81_DUMMY38;
    _zyL542_tfiRv82 <= _zyL542_tfiRv82_DUMMY39;
    _zyL555_tfiRv83 <= _zyL555_tfiRv83_DUMMY40;
    _zyL556_tfiRv84 <= _zyL556_tfiRv84_DUMMY41;
    _zyL569_tfiRv85 <= _zyL569_tfiRv85_DUMMY42;
    _zyL570_tfiRv86 <= _zyL570_tfiRv86_DUMMY43;
  end process ;

  process --:o6732
  (clk,rst_n)
  begin
    if (rst_n = '0') then
      fifo_in(68 downto 68) <= "0" ;
      key_blob_region <= '0' ;
      int_tlv_counter <= "000000" ;
    elsif (clk'event and clk = '1') then
      if (fifo_in_valid = '1') then

        case int_tlv_counter is
          when  "101001"  =>
            fifo_in(68 downto 68) <= "1" ;
          when  "101010"  =>
            fifo_in(68 downto 68) <= "0" ;
          when others =>
            fifo_in(68 downto 68) <= fifo_in(68 downto 68) ;
        end case;

        case int_tlv_counter is
          when  "010101"  =>
            key_blob_region <= '1' ;
          when  "101010"  =>
            key_blob_region <= '0' ;
          when others =>
            key_blob_region <= key_blob_region ;
        end case;

        case int_tlv_counter is
          when  "101010"  =>
            int_tlv_counter <= "000000" ;
          when others =>
            int_tlv_counter <= (int_tlv_counter + std_logic_vector'("000001")) ;
        end case;
      end if;
    end if ;
  end process ;

  process --:o6768
  (*)
  begin
    nxt_fifo_in_id <= fifo_in(64+3 downto 64) ;
    fifo_in(70 downto 70) <= (ext(fifo_in_valid,1) and boolean_to_std(fifo_in
    (64+3 downto 64) = KME_WORD0,1)) ;
    fifo_in(69 downto 69) <= "0" ;
    if (fifo_in_valid = '1') then

      case int_tlv_counter is
        when  "000000"  =>
          nxt_fifo_in_id <= KME_DEBUG_KEYHDR ;
          fifo_in(69 downto 69) <= "1" ;
        when  "000001"  =>
          nxt_fifo_in_id <= KME_GUID ;
          fifo_in(69 downto 69) <= "1" ;
        when  "000101"  =>
          nxt_fifo_in_id <= KME_IVTWEAK ;
          fifo_in(69 downto 69) <= "1" ;
        when  "000111"  =>
          nxt_fifo_in_id <= KME_KIM ;
          fifo_in(69 downto 69) <= "1" ;
        when  "001001"  =>
          nxt_fifo_in_id <= KME_DEK_CKV0 ;
          fifo_in(69 downto 69) <= "1" ;
        when  "001101"  =>
          nxt_fifo_in_id <= KME_DEK_CKV1 ;
          fifo_in(69 downto 69) <= "1" ;
        when  "010001"  =>
          nxt_fifo_in_id <= KME_DAK_CKV ;
          fifo_in(69 downto 69) <= "1" ;
        when  "010101"  =>
          nxt_fifo_in_id <= KME_EIV ;
          fifo_in(69 downto 69) <= "1" ;
        when  "010111"  =>
          nxt_fifo_in_id <= KME_DEK0 ;
          fifo_in(69 downto 69) <= "1" ;
        when  "011011"  =>
          nxt_fifo_in_id <= KME_DEK1 ;
          fifo_in(69 downto 69) <= "1" ;
        when  "011111"  =>
          nxt_fifo_in_id <= KME_ETAG ;
          fifo_in(69 downto 69) <= "1" ;
        when  "100001"  =>
          nxt_fifo_in_id <= KME_AIV ;
          fifo_in(69 downto 69) <= "1" ;
        when  "100011"  =>
          nxt_fifo_in_id <= KME_DAK ;
          fifo_in(69 downto 69) <= "1" ;
        when  "100111"  =>
          nxt_fifo_in_id <= KME_ATAG ;
          fifo_in(69 downto 69) <= "1" ;
        when  "101001"  =>
          nxt_fifo_in_id <= KME_ERROR ;
          fifo_in(69 downto 69) <= "1" ;
        when  "101010"  =>
          nxt_fifo_in_id <= KME_WORD0 ;
          fifo_in(69 downto 69) <= "1" ;
        when others => null ;
      end case;
    end if;
  end process ;
  Generate1 : if key_type_0_ : (TRUE) generate
    constant jj : integer := 0 ;
  begin

    process --:o6864
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_39_cpass, " ",
       _zy_sva_brcm_aux_cmd_39_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       889, std_logic_vector'("000"));
    end process ;

    process --:o6865
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_iv", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_iv_40_cpass, " ",
       _zy_sva_brcm_aux_cmd_iv_40_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       890, std_logic_vector'("000"));
    end process ;

    process --:o6866
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_guid", std_logic'('0'), std_logic_vector'("10"
      ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_guid_41_cpass, " ",
       _zy_sva_brcm_aux_cmd_guid_41_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       891, std_logic_vector'("000"));
    end process ;

    process --:o6867
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_guid_iv", std_logic'('0'), std_logic_vector'
      ("10"), " ", " ", " ", " ", " ", " ",
       _zy_sva_brcm_aux_cmd_guid_iv_42_cpass, " ",
       _zy_sva_brcm_aux_cmd_guid_iv_42_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       892, std_logic_vector'("000"));
    end process ;

    process --:o6868
    (**) -- always_comb
    begin
      $axis_assert( "brcm_key_type", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_key_type_43_cpass, " ",
       _zy_sva_brcm_key_type_43_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       893, std_logic_vector'("000"));
    end process ;
  end generate ;
  Generate2 : if key_type_1_ : (TRUE) generate
    constant jj : integer := 1 ;
  begin

    process --:o6874
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_44_cpass, " ",
       _zy_sva_brcm_aux_cmd_44_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       889, std_logic_vector'("000"));
    end process ;

    process --:o6875
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_iv", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_iv_45_cpass, " ",
       _zy_sva_brcm_aux_cmd_iv_45_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       890, std_logic_vector'("000"));
    end process ;

    process --:o6876
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_guid", std_logic'('0'), std_logic_vector'("10"
      ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_guid_46_cpass, " ",
       _zy_sva_brcm_aux_cmd_guid_46_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       891, std_logic_vector'("000"));
    end process ;

    process --:o6877
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_guid_iv", std_logic'('0'), std_logic_vector'
      ("10"), " ", " ", " ", " ", " ", " ",
       _zy_sva_brcm_aux_cmd_guid_iv_47_cpass, " ",
       _zy_sva_brcm_aux_cmd_guid_iv_47_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       892, std_logic_vector'("000"));
    end process ;

    process --:o6878
    (**) -- always_comb
    begin
      $axis_assert( "brcm_key_type", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_key_type_48_cpass, " ",
       _zy_sva_brcm_key_type_48_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       893, std_logic_vector'("000"));
    end process ;
  end generate ;
  Generate3 : if key_type_2_ : (TRUE) generate
    constant jj : integer := 2 ;
  begin

    process --:o6884
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_49_cpass, " ",
       _zy_sva_brcm_aux_cmd_49_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       889, std_logic_vector'("000"));
    end process ;

    process --:o6885
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_iv", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_iv_50_cpass, " ",
       _zy_sva_brcm_aux_cmd_iv_50_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       890, std_logic_vector'("000"));
    end process ;

    process --:o6886
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_guid", std_logic'('0'), std_logic_vector'("10"
      ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_guid_51_cpass, " ",
       _zy_sva_brcm_aux_cmd_guid_51_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       891, std_logic_vector'("000"));
    end process ;

    process --:o6887
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_guid_iv", std_logic'('0'), std_logic_vector'
      ("10"), " ", " ", " ", " ", " ", " ",
       _zy_sva_brcm_aux_cmd_guid_iv_52_cpass, " ",
       _zy_sva_brcm_aux_cmd_guid_iv_52_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       892, std_logic_vector'("000"));
    end process ;

    process --:o6888
    (**) -- always_comb
    begin
      $axis_assert( "brcm_key_type", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_key_type_53_cpass, " ",
       _zy_sva_brcm_key_type_53_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       893, std_logic_vector'("000"));
    end process ;
  end generate ;
  Generate4 : if key_type_3_ : (TRUE) generate
    constant jj : integer := 3 ;
  begin

    process --:o6894
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_54_cpass, " ",
       _zy_sva_brcm_aux_cmd_54_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       889, std_logic_vector'("000"));
    end process ;

    process --:o6895
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_iv", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_iv_55_cpass, " ",
       _zy_sva_brcm_aux_cmd_iv_55_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       890, std_logic_vector'("000"));
    end process ;

    process --:o6896
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_guid", std_logic'('0'), std_logic_vector'("10"
      ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_guid_56_cpass, " ",
       _zy_sva_brcm_aux_cmd_guid_56_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       891, std_logic_vector'("000"));
    end process ;

    process --:o6897
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_guid_iv", std_logic'('0'), std_logic_vector'
      ("10"), " ", " ", " ", " ", " ", " ",
       _zy_sva_brcm_aux_cmd_guid_iv_57_cpass, " ",
       _zy_sva_brcm_aux_cmd_guid_iv_57_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       892, std_logic_vector'("000"));
    end process ;

    process --:o6898
    (**) -- always_comb
    begin
      $axis_assert( "brcm_key_type", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_key_type_58_cpass, " ",
       _zy_sva_brcm_key_type_58_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       893, std_logic_vector'("000"));
    end process ;
  end generate ;
  Generate5 : if key_type_4_ : (TRUE) generate
    constant jj : integer := 4 ;
  begin

    process --:o6904
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_59_cpass, " ",
       _zy_sva_brcm_aux_cmd_59_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       889, std_logic_vector'("000"));
    end process ;

    process --:o6905
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_iv", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_iv_60_cpass, " ",
       _zy_sva_brcm_aux_cmd_iv_60_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       890, std_logic_vector'("000"));
    end process ;

    process --:o6906
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_guid", std_logic'('0'), std_logic_vector'("10"
      ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_guid_61_cpass, " ",
       _zy_sva_brcm_aux_cmd_guid_61_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       891, std_logic_vector'("000"));
    end process ;

    process --:o6907
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_guid_iv", std_logic'('0'), std_logic_vector'
      ("10"), " ", " ", " ", " ", " ", " ",
       _zy_sva_brcm_aux_cmd_guid_iv_62_cpass, " ",
       _zy_sva_brcm_aux_cmd_guid_iv_62_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       892, std_logic_vector'("000"));
    end process ;

    process --:o6908
    (**) -- always_comb
    begin
      $axis_assert( "brcm_key_type", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_key_type_63_cpass, " ",
       _zy_sva_brcm_key_type_63_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       893, std_logic_vector'("000"));
    end process ;
  end generate ;
  Generate6 : if key_type_5_ : (TRUE) generate
    constant jj : integer := 5 ;
  begin

    process --:o6914
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_64_cpass, " ",
       _zy_sva_brcm_aux_cmd_64_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       889, std_logic_vector'("000"));
    end process ;

    process --:o6915
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_iv", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_iv_65_cpass, " ",
       _zy_sva_brcm_aux_cmd_iv_65_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       890, std_logic_vector'("000"));
    end process ;

    process --:o6916
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_guid", std_logic'('0'), std_logic_vector'("10"
      ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_guid_66_cpass, " ",
       _zy_sva_brcm_aux_cmd_guid_66_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       891, std_logic_vector'("000"));
    end process ;

    process --:o6917
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_guid_iv", std_logic'('0'), std_logic_vector'
      ("10"), " ", " ", " ", " ", " ", " ",
       _zy_sva_brcm_aux_cmd_guid_iv_67_cpass, " ",
       _zy_sva_brcm_aux_cmd_guid_iv_67_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       892, std_logic_vector'("000"));
    end process ;

    process --:o6918
    (**) -- always_comb
    begin
      $axis_assert( "brcm_key_type", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_key_type_68_cpass, " ",
       _zy_sva_brcm_key_type_68_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       893, std_logic_vector'("000"));
    end process ;
  end generate ;
  Generate7 : if key_type_6_ : (TRUE) generate
    constant jj : integer := 6 ;
  begin

    process --:o6924
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_69_cpass, " ",
       _zy_sva_brcm_aux_cmd_69_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       889, std_logic_vector'("000"));
    end process ;

    process --:o6925
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_iv", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_iv_70_cpass, " ",
       _zy_sva_brcm_aux_cmd_iv_70_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       890, std_logic_vector'("000"));
    end process ;

    process --:o6926
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_guid", std_logic'('0'), std_logic_vector'("10"
      ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_guid_71_cpass, " ",
       _zy_sva_brcm_aux_cmd_guid_71_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       891, std_logic_vector'("000"));
    end process ;

    process --:o6927
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_guid_iv", std_logic'('0'), std_logic_vector'
      ("10"), " ", " ", " ", " ", " ", " ",
       _zy_sva_brcm_aux_cmd_guid_iv_72_cpass, " ",
       _zy_sva_brcm_aux_cmd_guid_iv_72_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       892, std_logic_vector'("000"));
    end process ;

    process --:o6928
    (**) -- always_comb
    begin
      $axis_assert( "brcm_key_type", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_key_type_73_cpass, " ",
       _zy_sva_brcm_key_type_73_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       893, std_logic_vector'("000"));
    end process ;
  end generate ;
  Generate8 : if key_type_7_ : (TRUE) generate
    constant jj : integer := 7 ;
  begin

    process --:o6934
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_74_cpass, " ",
       _zy_sva_brcm_aux_cmd_74_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       889, std_logic_vector'("000"));
    end process ;

    process --:o6935
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_iv", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_iv_75_cpass, " ",
       _zy_sva_brcm_aux_cmd_iv_75_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       890, std_logic_vector'("000"));
    end process ;

    process --:o6936
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_guid", std_logic'('0'), std_logic_vector'("10"
      ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_guid_76_cpass, " ",
       _zy_sva_brcm_aux_cmd_guid_76_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       891, std_logic_vector'("000"));
    end process ;

    process --:o6937
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_guid_iv", std_logic'('0'), std_logic_vector'
      ("10"), " ", " ", " ", " ", " ", " ",
       _zy_sva_brcm_aux_cmd_guid_iv_77_cpass, " ",
       _zy_sva_brcm_aux_cmd_guid_iv_77_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       892, std_logic_vector'("000"));
    end process ;

    process --:o6938
    (**) -- always_comb
    begin
      $axis_assert( "brcm_key_type", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_key_type_78_cpass, " ",
       _zy_sva_brcm_key_type_78_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       893, std_logic_vector'("000"));
    end process ;
  end generate ;
  Generate9 : if key_type_8_ : (TRUE) generate
    constant jj : integer := 8 ;
  begin

    process --:o6944
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_79_cpass, " ",
       _zy_sva_brcm_aux_cmd_79_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       889, std_logic_vector'("000"));
    end process ;

    process --:o6945
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_iv", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_iv_80_cpass, " ",
       _zy_sva_brcm_aux_cmd_iv_80_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       890, std_logic_vector'("000"));
    end process ;

    process --:o6946
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_guid", std_logic'('0'), std_logic_vector'("10"
      ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_guid_81_cpass, " ",
       _zy_sva_brcm_aux_cmd_guid_81_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       891, std_logic_vector'("000"));
    end process ;

    process --:o6947
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_guid_iv", std_logic'('0'), std_logic_vector'
      ("10"), " ", " ", " ", " ", " ", " ",
       _zy_sva_brcm_aux_cmd_guid_iv_82_cpass, " ",
       _zy_sva_brcm_aux_cmd_guid_iv_82_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       892, std_logic_vector'("000"));
    end process ;

    process --:o6948
    (**) -- always_comb
    begin
      $axis_assert( "brcm_key_type", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_key_type_83_cpass, " ",
       _zy_sva_brcm_key_type_83_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       893, std_logic_vector'("000"));
    end process ;
  end generate ;
  Generate10 : if key_type_9_ : (TRUE) generate
    constant jj : integer := 9 ;
  begin

    process --:o6954
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_84_cpass, " ",
       _zy_sva_brcm_aux_cmd_84_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       889, std_logic_vector'("000"));
    end process ;

    process --:o6955
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_iv", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_iv_85_cpass, " ",
       _zy_sva_brcm_aux_cmd_iv_85_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       890, std_logic_vector'("000"));
    end process ;

    process --:o6956
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_guid", std_logic'('0'), std_logic_vector'("10"
      ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_guid_86_cpass, " ",
       _zy_sva_brcm_aux_cmd_guid_86_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       891, std_logic_vector'("000"));
    end process ;

    process --:o6957
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_guid_iv", std_logic'('0'), std_logic_vector'
      ("10"), " ", " ", " ", " ", " ", " ",
       _zy_sva_brcm_aux_cmd_guid_iv_87_cpass, " ",
       _zy_sva_brcm_aux_cmd_guid_iv_87_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       892, std_logic_vector'("000"));
    end process ;

    process --:o6958
    (**) -- always_comb
    begin
      $axis_assert( "brcm_key_type", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_key_type_88_cpass, " ",
       _zy_sva_brcm_key_type_88_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       893, std_logic_vector'("000"));
    end process ;
  end generate ;
  Generate11 : if key_type_10_ : (TRUE) generate
    constant jj : integer := 10 ;
  begin

    process --:o6964
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_89_cpass, " ",
       _zy_sva_brcm_aux_cmd_89_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       889, std_logic_vector'("000"));
    end process ;

    process --:o6965
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_iv", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_iv_90_cpass, " ",
       _zy_sva_brcm_aux_cmd_iv_90_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       890, std_logic_vector'("000"));
    end process ;

    process --:o6966
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_guid", std_logic'('0'), std_logic_vector'("10"
      ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_guid_91_cpass, " ",
       _zy_sva_brcm_aux_cmd_guid_91_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       891, std_logic_vector'("000"));
    end process ;

    process --:o6967
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_guid_iv", std_logic'('0'), std_logic_vector'
      ("10"), " ", " ", " ", " ", " ", " ",
       _zy_sva_brcm_aux_cmd_guid_iv_92_cpass, " ",
       _zy_sva_brcm_aux_cmd_guid_iv_92_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       892, std_logic_vector'("000"));
    end process ;

    process --:o6968
    (**) -- always_comb
    begin
      $axis_assert( "brcm_key_type", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_key_type_93_cpass, " ",
       _zy_sva_brcm_key_type_93_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       893, std_logic_vector'("000"));
    end process ;
  end generate ;
  Generate12 : if key_type_11_ : (TRUE) generate
    constant jj : integer := 11 ;
  begin

    process --:o6974
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_94_cpass, " ",
       _zy_sva_brcm_aux_cmd_94_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       889, std_logic_vector'("000"));
    end process ;

    process --:o6975
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_iv", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_iv_95_cpass, " ",
       _zy_sva_brcm_aux_cmd_iv_95_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       890, std_logic_vector'("000"));
    end process ;

    process --:o6976
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_guid", std_logic'('0'), std_logic_vector'("10"
      ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_guid_96_cpass, " ",
       _zy_sva_brcm_aux_cmd_guid_96_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       891, std_logic_vector'("000"));
    end process ;

    process --:o6977
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_guid_iv", std_logic'('0'), std_logic_vector'
      ("10"), " ", " ", " ", " ", " ", " ",
       _zy_sva_brcm_aux_cmd_guid_iv_97_cpass, " ",
       _zy_sva_brcm_aux_cmd_guid_iv_97_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       892, std_logic_vector'("000"));
    end process ;

    process --:o6978
    (**) -- always_comb
    begin
      $axis_assert( "brcm_key_type", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_key_type_98_cpass, " ",
       _zy_sva_brcm_key_type_98_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       893, std_logic_vector'("000"));
    end process ;
  end generate ;
  Generate13 : if key_type_12_ : (TRUE) generate
    constant jj : integer := 12 ;
  begin

    process --:o6984
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_99_cpass, " ",
       _zy_sva_brcm_aux_cmd_99_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       889, std_logic_vector'("000"));
    end process ;

    process --:o6985
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_iv", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_iv_100_cpass, " ",
       _zy_sva_brcm_aux_cmd_iv_100_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       890, std_logic_vector'("000"));
    end process ;

    process --:o6986
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_guid", std_logic'('0'), std_logic_vector'("10"
      ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_guid_101_cpass, " ",
       _zy_sva_brcm_aux_cmd_guid_101_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       891, std_logic_vector'("000"));
    end process ;

    process --:o6987
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_guid_iv", std_logic'('0'), std_logic_vector'
      ("10"), " ", " ", " ", " ", " ", " ",
       _zy_sva_brcm_aux_cmd_guid_iv_102_cpass, " ",
       _zy_sva_brcm_aux_cmd_guid_iv_102_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       892, std_logic_vector'("000"));
    end process ;

    process --:o6988
    (**) -- always_comb
    begin
      $axis_assert( "brcm_key_type", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_key_type_103_cpass, " ",
       _zy_sva_brcm_key_type_103_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       893, std_logic_vector'("000"));
    end process ;
  end generate ;
  Generate14 : if key_type_13_ : (TRUE) generate
    constant jj : integer := 13 ;
  begin

    process --:o6994
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_104_cpass, " ",
       _zy_sva_brcm_aux_cmd_104_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       889, std_logic_vector'("000"));
    end process ;

    process --:o6995
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_iv", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_iv_105_cpass, " ",
       _zy_sva_brcm_aux_cmd_iv_105_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       890, std_logic_vector'("000"));
    end process ;

    process --:o6996
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_guid", std_logic'('0'), std_logic_vector'("10"
      ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_aux_cmd_guid_106_cpass, " ",
       _zy_sva_brcm_aux_cmd_guid_106_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       891, std_logic_vector'("000"));
    end process ;

    process --:o6997
    (**) -- always_comb
    begin
      $axis_assert( "brcm_aux_cmd_guid_iv", std_logic'('0'), std_logic_vector'
      ("10"), " ", " ", " ", " ", " ", " ",
       _zy_sva_brcm_aux_cmd_guid_iv_107_cpass, " ",
       _zy_sva_brcm_aux_cmd_guid_iv_107_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       892, std_logic_vector'("000"));
    end process ;

    process --:o6998
    (**) -- always_comb
    begin
      $axis_assert( "brcm_key_type", std_logic'('0'), std_logic_vector'("10"),
       " ", " ", " ", " ", " ", " ", _zy_sva_brcm_key_type_108_cpass, " ",
       _zy_sva_brcm_key_type_108_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       893, std_logic_vector'("000"));
    end process ;
  end generate ;
  Generate15 : if kdf_mode_0_ : (TRUE) generate
    constant ii : integer := 0 ;
  begin
    Generate16 : if dek_op_0_ : (TRUE) generate
      constant jj : integer := 0 ;
    begin
      Generate17 : if dak_op_0_ : (TRUE) generate
        constant kk : integer := 0 ;
      begin

        process --:o7012
        (**) -- always_comb
        begin
          $axis_assert( "brcm_kdf_ops", std_logic'('0'), std_logic_vector'("10"
          ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_kdf_ops_109_cpass, " ",
           _zy_sva_brcm_kdf_ops_109_ccheck, " ",
           "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
           902, std_logic_vector'("000"));
        end process ;
      end generate ;
      Generate18 : if dak_op_1_ : (TRUE) generate
        constant kk : integer := 1 ;
      begin

        process --:o7018
        (**) -- always_comb
        begin
          $axis_assert( "brcm_kdf_ops", std_logic'('0'), std_logic_vector'("10"
          ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_kdf_ops_110_cpass, " ",
           _zy_sva_brcm_kdf_ops_110_ccheck, " ",
           "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
           902, std_logic_vector'("000"));
        end process ;
      end generate ;
    end generate ;
    Generate19 : if dek_op_1_ : (TRUE) generate
      constant jj : integer := 1 ;
    begin
      Generate20 : if dak_op_0_ : (TRUE) generate
        constant kk : integer := 0 ;
      begin

        process --:o7029
        (**) -- always_comb
        begin
          $axis_assert( "brcm_kdf_ops", std_logic'('0'), std_logic_vector'("10"
          ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_kdf_ops_111_cpass, " ",
           _zy_sva_brcm_kdf_ops_111_ccheck, " ",
           "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
           902, std_logic_vector'("000"));
        end process ;
      end generate ;
      Generate21 : if dak_op_1_ : (TRUE) generate
        constant kk : integer := 1 ;
      begin

        process --:o7035
        (**) -- always_comb
        begin
          $axis_assert( "brcm_kdf_ops", std_logic'('0'), std_logic_vector'("10"
          ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_kdf_ops_112_cpass, " ",
           _zy_sva_brcm_kdf_ops_112_ccheck, " ",
           "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
           902, std_logic_vector'("000"));
        end process ;
      end generate ;
    end generate ;
  end generate ;
  Generate22 : if kdf_mode_1_ : (TRUE) generate
    constant ii : integer := 1 ;
  begin
    Generate23 : if dek_op_0_ : (TRUE) generate
      constant jj : integer := 0 ;
    begin
      Generate24 : if dak_op_0_ : (TRUE) generate
        constant kk : integer := 0 ;
      begin

        process --:o7051
        (**) -- always_comb
        begin
          $axis_assert( "brcm_kdf_ops", std_logic'('0'), std_logic_vector'("10"
          ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_kdf_ops_113_cpass, " ",
           _zy_sva_brcm_kdf_ops_113_ccheck, " ",
           "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
           902, std_logic_vector'("000"));
        end process ;
      end generate ;
      Generate25 : if dak_op_1_ : (TRUE) generate
        constant kk : integer := 1 ;
      begin

        process --:o7057
        (**) -- always_comb
        begin
          $axis_assert( "brcm_kdf_ops", std_logic'('0'), std_logic_vector'("10"
          ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_kdf_ops_114_cpass, " ",
           _zy_sva_brcm_kdf_ops_114_ccheck, " ",
           "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
           902, std_logic_vector'("000"));
        end process ;
      end generate ;
    end generate ;
    Generate26 : if dek_op_1_ : (TRUE) generate
      constant jj : integer := 1 ;
    begin
      Generate27 : if dak_op_0_ : (TRUE) generate
        constant kk : integer := 0 ;
      begin

        process --:o7068
        (**) -- always_comb
        begin
          $axis_assert( "brcm_kdf_ops", std_logic'('0'), std_logic_vector'("10"
          ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_kdf_ops_115_cpass, " ",
           _zy_sva_brcm_kdf_ops_115_ccheck, " ",
           "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
           902, std_logic_vector'("000"));
        end process ;
      end generate ;
      Generate28 : if dak_op_1_ : (TRUE) generate
        constant kk : integer := 1 ;
      begin

        process --:o7074
        (**) -- always_comb
        begin
          $axis_assert( "brcm_kdf_ops", std_logic'('0'), std_logic_vector'("10"
          ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_kdf_ops_116_cpass, " ",
           _zy_sva_brcm_kdf_ops_116_ccheck, " ",
           "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
           902, std_logic_vector'("000"));
        end process ;
      end generate ;
    end generate ;
  end generate ;
  Generate29 : if kdf_mode_2_ : (TRUE) generate
    constant ii : integer := 2 ;
  begin
    Generate30 : if dek_op_0_ : (TRUE) generate
      constant jj : integer := 0 ;
    begin
      Generate31 : if dak_op_0_ : (TRUE) generate
        constant kk : integer := 0 ;
      begin

        process --:o7090
        (**) -- always_comb
        begin
          $axis_assert( "brcm_kdf_ops", std_logic'('0'), std_logic_vector'("10"
          ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_kdf_ops_117_cpass, " ",
           _zy_sva_brcm_kdf_ops_117_ccheck, " ",
           "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
           902, std_logic_vector'("000"));
        end process ;
      end generate ;
      Generate32 : if dak_op_1_ : (TRUE) generate
        constant kk : integer := 1 ;
      begin

        process --:o7096
        (**) -- always_comb
        begin
          $axis_assert( "brcm_kdf_ops", std_logic'('0'), std_logic_vector'("10"
          ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_kdf_ops_118_cpass, " ",
           _zy_sva_brcm_kdf_ops_118_ccheck, " ",
           "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
           902, std_logic_vector'("000"));
        end process ;
      end generate ;
    end generate ;
    Generate33 : if dek_op_1_ : (TRUE) generate
      constant jj : integer := 1 ;
    begin
      Generate34 : if dak_op_0_ : (TRUE) generate
        constant kk : integer := 0 ;
      begin

        process --:o7107
        (**) -- always_comb
        begin
          $axis_assert( "brcm_kdf_ops", std_logic'('0'), std_logic_vector'("10"
          ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_kdf_ops_119_cpass, " ",
           _zy_sva_brcm_kdf_ops_119_ccheck, " ",
           "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
           902, std_logic_vector'("000"));
        end process ;
      end generate ;
      Generate35 : if dak_op_1_ : (TRUE) generate
        constant kk : integer := 1 ;
      begin

        process --:o7113
        (**) -- always_comb
        begin
          $axis_assert( "brcm_kdf_ops", std_logic'('0'), std_logic_vector'("10"
          ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_kdf_ops_120_cpass, " ",
           _zy_sva_brcm_kdf_ops_120_ccheck, " ",
           "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
           902, std_logic_vector'("000"));
        end process ;
      end generate ;
    end generate ;
  end generate ;
  Generate36 : if kdf_mode_3_ : (TRUE) generate
    constant ii : integer := 3 ;
  begin
    Generate37 : if dek_op_0_ : (TRUE) generate
      constant jj : integer := 0 ;
    begin
      Generate38 : if dak_op_0_ : (TRUE) generate
        constant kk : integer := 0 ;
      begin

        process --:o7129
        (**) -- always_comb
        begin
          $axis_assert( "brcm_kdf_ops", std_logic'('0'), std_logic_vector'("10"
          ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_kdf_ops_121_cpass, " ",
           _zy_sva_brcm_kdf_ops_121_ccheck, " ",
           "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
           902, std_logic_vector'("000"));
        end process ;
      end generate ;
      Generate39 : if dak_op_1_ : (TRUE) generate
        constant kk : integer := 1 ;
      begin

        process --:o7135
        (**) -- always_comb
        begin
          $axis_assert( "brcm_kdf_ops", std_logic'('0'), std_logic_vector'("10"
          ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_kdf_ops_122_cpass, " ",
           _zy_sva_brcm_kdf_ops_122_ccheck, " ",
           "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
           902, std_logic_vector'("000"));
        end process ;
      end generate ;
    end generate ;
    Generate40 : if dek_op_1_ : (TRUE) generate
      constant jj : integer := 1 ;
    begin
      Generate41 : if dak_op_0_ : (TRUE) generate
        constant kk : integer := 0 ;
      begin

        process --:o7146
        (**) -- always_comb
        begin
          $axis_assert( "brcm_kdf_ops", std_logic'('0'), std_logic_vector'("10"
          ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_kdf_ops_123_cpass, " ",
           _zy_sva_brcm_kdf_ops_123_ccheck, " ",
           "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
           902, std_logic_vector'("000"));
        end process ;
      end generate ;
      Generate42 : if dak_op_1_ : (TRUE) generate
        constant kk : integer := 1 ;
      begin

        process --:o7152
        (**) -- always_comb
        begin
          $axis_assert( "brcm_kdf_ops", std_logic'('0'), std_logic_vector'("10"
          ), " ", " ", " ", " ", " ", " ", _zy_sva_brcm_kdf_ops_124_cpass, " ",
           _zy_sva_brcm_kdf_ops_124_ccheck, " ",
           "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
           902, std_logic_vector'("000"));
        end process ;
      end generate ;
    end generate ;
  end generate ;
  Generate43 : if key_type_enc_dek_7_ : (TRUE) generate
    constant nn : integer := 7 ;
  begin

    process --:o7160
    (**) -- always_comb
    begin
      $axis_assert( "null_gcm", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_null_gcm_125_cpass, " ",
       _zy_sva_null_gcm_125_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1114, std_logic_vector'("000"));
    end process ;

    process --:o7161
    (**) -- always_comb
    begin
      $axis_assert( "sha_gcm", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_sha_gcm_126_cpass, " ",
       _zy_sva_sha_gcm_126_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1121, std_logic_vector'("000"));
    end process ;

    process --:o7162
    (**) -- always_comb
    begin
      $axis_assert( "null_xts", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_null_xts_127_cpass, " ",
       _zy_sva_null_xts_127_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1127, std_logic_vector'("000"));
    end process ;

    process --:o7163
    (**) -- always_comb
    begin
      $axis_assert( "sha_xts", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_sha_xts_128_cpass, " ",
       _zy_sva_sha_xts_128_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1133, std_logic_vector'("000"));
    end process ;

    process --:o7164
    (**) -- always_comb
    begin
      $axis_assert( "null_null", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_null_null_129_cpass, " ",
       _zy_sva_null_null_129_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1139, std_logic_vector'("000"));
    end process ;

    process --:o7165
    (**) -- always_comb
    begin
      $axis_assert( "sha_null", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_sha_null_130_cpass, " ",
       _zy_sva_sha_null_130_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1145, std_logic_vector'("000"));
    end process ;

    process --:o7166
    (**) -- always_comb
    begin
      $axis_assert( "hmac_gcm", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_hmac_gcm_131_cpass, " ",
       _zy_sva_hmac_gcm_131_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1152, std_logic_vector'("000"));
    end process ;

    process --:o7167
    (**) -- always_comb
    begin
      $axis_assert( "hmac_xts", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_hmac_xts_132_cpass, " ",
       _zy_sva_hmac_xts_132_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1158, std_logic_vector'("000"));
    end process ;

    process --:o7168
    (**) -- always_comb
    begin
      $axis_assert( "hmac_null", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_hmac_null_133_cpass, " ",
       _zy_sva_hmac_null_133_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1164, std_logic_vector'("000"));
    end process ;
  end generate ;
  Generate44 : if key_type_enc_dek_8_ : (TRUE) generate
    constant nn : integer := 8 ;
  begin

    process --:o7174
    (**) -- always_comb
    begin
      $axis_assert( "null_gcm", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_null_gcm_134_cpass, " ",
       _zy_sva_null_gcm_134_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1114, std_logic_vector'("000"));
    end process ;

    process --:o7175
    (**) -- always_comb
    begin
      $axis_assert( "sha_gcm", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_sha_gcm_135_cpass, " ",
       _zy_sva_sha_gcm_135_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1121, std_logic_vector'("000"));
    end process ;

    process --:o7176
    (**) -- always_comb
    begin
      $axis_assert( "null_xts", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_null_xts_136_cpass, " ",
       _zy_sva_null_xts_136_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1127, std_logic_vector'("000"));
    end process ;

    process --:o7177
    (**) -- always_comb
    begin
      $axis_assert( "sha_xts", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_sha_xts_137_cpass, " ",
       _zy_sva_sha_xts_137_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1133, std_logic_vector'("000"));
    end process ;

    process --:o7178
    (**) -- always_comb
    begin
      $axis_assert( "null_null", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_null_null_138_cpass, " ",
       _zy_sva_null_null_138_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1139, std_logic_vector'("000"));
    end process ;

    process --:o7179
    (**) -- always_comb
    begin
      $axis_assert( "sha_null", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_sha_null_139_cpass, " ",
       _zy_sva_sha_null_139_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1145, std_logic_vector'("000"));
    end process ;

    process --:o7180
    (**) -- always_comb
    begin
      $axis_assert( "hmac_gcm", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_hmac_gcm_140_cpass, " ",
       _zy_sva_hmac_gcm_140_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1152, std_logic_vector'("000"));
    end process ;

    process --:o7181
    (**) -- always_comb
    begin
      $axis_assert( "hmac_xts", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_hmac_xts_141_cpass, " ",
       _zy_sva_hmac_xts_141_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1158, std_logic_vector'("000"));
    end process ;

    process --:o7182
    (**) -- always_comb
    begin
      $axis_assert( "hmac_null", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_hmac_null_142_cpass, " ",
       _zy_sva_hmac_null_142_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1164, std_logic_vector'("000"));
    end process ;
  end generate ;
  Generate45 : if key_type_enc_dek_dak_10_ : (TRUE) generate
    constant qq : integer := 10 ;
  begin

    process --:o7188
    (**) -- always_comb
    begin
      $axis_assert( "null_gcm", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_null_gcm_143_cpass, " ",
       _zy_sva_null_gcm_143_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1175, std_logic_vector'("000"));
    end process ;

    process --:o7189
    (**) -- always_comb
    begin
      $axis_assert( "sha_gcm", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_sha_gcm_144_cpass, " ",
       _zy_sva_sha_gcm_144_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1182, std_logic_vector'("000"));
    end process ;

    process --:o7190
    (**) -- always_comb
    begin
      $axis_assert( "null_xts", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_null_xts_145_cpass, " ",
       _zy_sva_null_xts_145_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1188, std_logic_vector'("000"));
    end process ;

    process --:o7191
    (**) -- always_comb
    begin
      $axis_assert( "sha_xts", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_sha_xts_146_cpass, " ",
       _zy_sva_sha_xts_146_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1194, std_logic_vector'("000"));
    end process ;

    process --:o7192
    (**) -- always_comb
    begin
      $axis_assert( "null_null", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_null_null_147_cpass, " ",
       _zy_sva_null_null_147_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1200, std_logic_vector'("000"));
    end process ;

    process --:o7193
    (**) -- always_comb
    begin
      $axis_assert( "sha_null", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_sha_null_148_cpass, " ",
       _zy_sva_sha_null_148_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1206, std_logic_vector'("000"));
    end process ;

    process --:o7194
    (**) -- always_comb
    begin
      $axis_assert( "hmac_gcm", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_hmac_gcm_149_cpass, " ",
       _zy_sva_hmac_gcm_149_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1213, std_logic_vector'("000"));
    end process ;

    process --:o7195
    (**) -- always_comb
    begin
      $axis_assert( "hmac_xts", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_hmac_xts_150_cpass, " ",
       _zy_sva_hmac_xts_150_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1219, std_logic_vector'("000"));
    end process ;

    process --:o7196
    (**) -- always_comb
    begin
      $axis_assert( "hmac_null", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_hmac_null_151_cpass, " ",
       _zy_sva_hmac_null_151_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1225, std_logic_vector'("000"));
    end process ;
  end generate ;
  Generate46 : if key_type_enc_dek_dak_11_ : (TRUE) generate
    constant qq : integer := 11 ;
  begin

    process --:o7202
    (**) -- always_comb
    begin
      $axis_assert( "null_gcm", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_null_gcm_152_cpass, " ",
       _zy_sva_null_gcm_152_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1175, std_logic_vector'("000"));
    end process ;

    process --:o7203
    (**) -- always_comb
    begin
      $axis_assert( "sha_gcm", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_sha_gcm_153_cpass, " ",
       _zy_sva_sha_gcm_153_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1182, std_logic_vector'("000"));
    end process ;

    process --:o7204
    (**) -- always_comb
    begin
      $axis_assert( "null_xts", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_null_xts_154_cpass, " ",
       _zy_sva_null_xts_154_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1188, std_logic_vector'("000"));
    end process ;

    process --:o7205
    (**) -- always_comb
    begin
      $axis_assert( "sha_xts", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_sha_xts_155_cpass, " ",
       _zy_sva_sha_xts_155_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1194, std_logic_vector'("000"));
    end process ;

    process --:o7206
    (**) -- always_comb
    begin
      $axis_assert( "null_null", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_null_null_156_cpass, " ",
       _zy_sva_null_null_156_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1200, std_logic_vector'("000"));
    end process ;

    process --:o7207
    (**) -- always_comb
    begin
      $axis_assert( "sha_null", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_sha_null_157_cpass, " ",
       _zy_sva_sha_null_157_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1206, std_logic_vector'("000"));
    end process ;

    process --:o7208
    (**) -- always_comb
    begin
      $axis_assert( "hmac_gcm", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_hmac_gcm_158_cpass, " ",
       _zy_sva_hmac_gcm_158_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1213, std_logic_vector'("000"));
    end process ;

    process --:o7209
    (**) -- always_comb
    begin
      $axis_assert( "hmac_xts", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_hmac_xts_159_cpass, " ",
       _zy_sva_hmac_xts_159_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1219, std_logic_vector'("000"));
    end process ;

    process --:o7210
    (**) -- always_comb
    begin
      $axis_assert( "hmac_null", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_hmac_null_160_cpass, " ",
       _zy_sva_hmac_null_160_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1225, std_logic_vector'("000"));
    end process ;
  end generate ;
  Generate47 : if key_type_enc_dek_dak_12_ : (TRUE) generate
    constant qq : integer := 12 ;
  begin

    process --:o7216
    (**) -- always_comb
    begin
      $axis_assert( "null_gcm", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_null_gcm_161_cpass, " ",
       _zy_sva_null_gcm_161_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1175, std_logic_vector'("000"));
    end process ;

    process --:o7217
    (**) -- always_comb
    begin
      $axis_assert( "sha_gcm", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_sha_gcm_162_cpass, " ",
       _zy_sva_sha_gcm_162_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1182, std_logic_vector'("000"));
    end process ;

    process --:o7218
    (**) -- always_comb
    begin
      $axis_assert( "null_xts", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_null_xts_163_cpass, " ",
       _zy_sva_null_xts_163_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1188, std_logic_vector'("000"));
    end process ;

    process --:o7219
    (**) -- always_comb
    begin
      $axis_assert( "sha_xts", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_sha_xts_164_cpass, " ",
       _zy_sva_sha_xts_164_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1194, std_logic_vector'("000"));
    end process ;

    process --:o7220
    (**) -- always_comb
    begin
      $axis_assert( "null_null", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_null_null_165_cpass, " ",
       _zy_sva_null_null_165_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1200, std_logic_vector'("000"));
    end process ;

    process --:o7221
    (**) -- always_comb
    begin
      $axis_assert( "sha_null", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_sha_null_166_cpass, " ",
       _zy_sva_sha_null_166_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1206, std_logic_vector'("000"));
    end process ;

    process --:o7222
    (**) -- always_comb
    begin
      $axis_assert( "hmac_gcm", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_hmac_gcm_167_cpass, " ",
       _zy_sva_hmac_gcm_167_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1213, std_logic_vector'("000"));
    end process ;

    process --:o7223
    (**) -- always_comb
    begin
      $axis_assert( "hmac_xts", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_hmac_xts_168_cpass, " ",
       _zy_sva_hmac_xts_168_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1219, std_logic_vector'("000"));
    end process ;

    process --:o7224
    (**) -- always_comb
    begin
      $axis_assert( "hmac_null", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_hmac_null_169_cpass, " ",
       _zy_sva_hmac_null_169_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1225, std_logic_vector'("000"));
    end process ;
  end generate ;
  Generate48 : if key_type_enc_dek_dak_13_ : (TRUE) generate
    constant qq : integer := 13 ;
  begin

    process --:o7230
    (**) -- always_comb
    begin
      $axis_assert( "null_gcm", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_null_gcm_170_cpass, " ",
       _zy_sva_null_gcm_170_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1175, std_logic_vector'("000"));
    end process ;

    process --:o7231
    (**) -- always_comb
    begin
      $axis_assert( "sha_gcm", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_sha_gcm_171_cpass, " ",
       _zy_sva_sha_gcm_171_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1182, std_logic_vector'("000"));
    end process ;

    process --:o7232
    (**) -- always_comb
    begin
      $axis_assert( "null_xts", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_null_xts_172_cpass, " ",
       _zy_sva_null_xts_172_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1188, std_logic_vector'("000"));
    end process ;

    process --:o7233
    (**) -- always_comb
    begin
      $axis_assert( "sha_xts", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_sha_xts_173_cpass, " ",
       _zy_sva_sha_xts_173_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1194, std_logic_vector'("000"));
    end process ;

    process --:o7234
    (**) -- always_comb
    begin
      $axis_assert( "null_null", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_null_null_174_cpass, " ",
       _zy_sva_null_null_174_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1200, std_logic_vector'("000"));
    end process ;

    process --:o7235
    (**) -- always_comb
    begin
      $axis_assert( "sha_null", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_sha_null_175_cpass, " ",
       _zy_sva_sha_null_175_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1206, std_logic_vector'("000"));
    end process ;

    process --:o7236
    (**) -- always_comb
    begin
      $axis_assert( "hmac_gcm", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_hmac_gcm_176_cpass, " ",
       _zy_sva_hmac_gcm_176_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1213, std_logic_vector'("000"));
    end process ;

    process --:o7237
    (**) -- always_comb
    begin
      $axis_assert( "hmac_xts", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_hmac_xts_177_cpass, " ",
       _zy_sva_hmac_xts_177_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1219, std_logic_vector'("000"));
    end process ;

    process --:o7238
    (**) -- always_comb
    begin
      $axis_assert( "hmac_null", std_logic'('0'), std_logic_vector'("10"), " ",
       " ", " ", " ", " ", " ", _zy_sva_hmac_null_178_cpass, " ",
       _zy_sva_hmac_null_178_ccheck, " ",
       "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",
       1225, std_logic_vector'("000"));
    end process ;
  end generate ;

  process --:o7240
  (**) -- always_comb
  begin
    $axis_assert( "key_type0_line4", std_logic'('0'), std_logic_vector'("10"),
     " ", " ", " ", " ", " ", " ", _zy_sva_key_type0_line4_1_cpass, " ",
     _zy_sva_key_type0_line4_1_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 914,
     std_logic_vector'("000"));
  end process ;

  process --:o7241
  (**) -- always_comb
  begin
    $axis_assert( "key_type0_line5a", std_logic'('0'), std_logic_vector'("10"),
     " ", " ", " ", " ", " ", " ", _zy_sva_key_type0_line5a_2_cpass, " ",
     _zy_sva_key_type0_line5a_2_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 920,
     std_logic_vector'("000"));
  end process ;

  process --:o7242
  (**) -- always_comb
  begin
    $axis_assert( "key_type0_line5b", std_logic'('0'), std_logic_vector'("10"),
     " ", " ", " ", " ", " ", " ", _zy_sva_key_type0_line5b_3_cpass, " ",
     _zy_sva_key_type0_line5b_3_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 926,
     std_logic_vector'("000"));
  end process ;

  process --:o7243
  (**) -- always_comb
  begin
    $axis_assert( "key_type1_line7a", std_logic'('0'), std_logic_vector'("10"),
     " ", " ", " ", " ", " ", " ", _zy_sva_key_type1_line7a_4_cpass, " ",
     _zy_sva_key_type1_line7a_4_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 936,
     std_logic_vector'("000"));
  end process ;

  process --:o7244
  (**) -- always_comb
  begin
    $axis_assert( "key_type1_line7b", std_logic'('0'), std_logic_vector'("10"),
     " ", " ", " ", " ", " ", " ", _zy_sva_key_type1_line7b_5_cpass, " ",
     _zy_sva_key_type1_line7b_5_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 944,
     std_logic_vector'("000"));
  end process ;

  process --:o7245
  (**) -- always_comb
  begin
    $axis_assert( "key_type1_line8a", std_logic'('0'), std_logic_vector'("10"),
     " ", " ", " ", " ", " ", " ", _zy_sva_key_type1_line8a_6_cpass, " ",
     _zy_sva_key_type1_line8a_6_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 952,
     std_logic_vector'("000"));
  end process ;

  process --:o7246
  (**) -- always_comb
  begin
    $axis_assert( "key_type1_line8b", std_logic'('0'), std_logic_vector'("10"),
     " ", " ", " ", " ", " ", " ", _zy_sva_key_type1_line8b_7_cpass, " ",
     _zy_sva_key_type1_line8b_7_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 960,
     std_logic_vector'("000"));
  end process ;

  process --:o7247
  (**) -- always_comb
  begin
    $axis_assert( "key_type1_line9", std_logic'('0'), std_logic_vector'("10"),
     " ", " ", " ", " ", " ", " ", _zy_sva_key_type1_line9_8_cpass, " ",
     _zy_sva_key_type1_line9_8_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 969,
     std_logic_vector'("000"));
  end process ;

  process --:o7248
  (**) -- always_comb
  begin
    $axis_assert( "key_type1_line10", std_logic'('0'), std_logic_vector'("10"),
     " ", " ", " ", " ", " ", " ", _zy_sva_key_type1_line10_9_cpass, " ",
     _zy_sva_key_type1_line10_9_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 977,
     std_logic_vector'("000"));
  end process ;

  process --:o7249
  (**) -- always_comb
  begin
    $axis_assert( "key_type1_line11a", std_logic'('0'), std_logic_vector'("10"),
     " ", " ", " ", " ", " ", " ", _zy_sva_key_type1_line11a_10_cpass, " ",
     _zy_sva_key_type1_line11a_10_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 983,
     std_logic_vector'("000"));
  end process ;

  process --:o7250
  (**) -- always_comb
  begin
    $axis_assert( "key_type1_line11b", std_logic'('0'), std_logic_vector'("10"),
     " ", " ", " ", " ", " ", " ", _zy_sva_key_type1_line11b_11_cpass, " ",
     _zy_sva_key_type1_line11b_11_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 989,
     std_logic_vector'("000"));
  end process ;

  process --:o7251
  (**) -- always_comb
  begin
    $axis_assert( "key_type1_line11c", std_logic'('0'), std_logic_vector'("10"),
     " ", " ", " ", " ", " ", " ", _zy_sva_key_type1_line11c_12_cpass, " ",
     _zy_sva_key_type1_line11c_12_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 995,
     std_logic_vector'("000"));
  end process ;

  process --:o7252
  (**) -- always_comb
  begin
    $axis_assert( "key_type1_line11d", std_logic'('0'), std_logic_vector'("10"),
     " ", " ", " ", " ", " ", " ", _zy_sva_key_type1_line11d_13_cpass, " ",
     _zy_sva_key_type1_line11d_13_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 1001,
     std_logic_vector'("000"));
  end process ;

  process --:o7253
  (**) -- always_comb
  begin
    $axis_assert( "key_type1_line12a", std_logic'('0'), std_logic_vector'("10"),
     " ", " ", " ", " ", " ", " ", _zy_sva_key_type1_line12a_14_cpass, " ",
     _zy_sva_key_type1_line12a_14_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 1007,
     std_logic_vector'("000"));
  end process ;

  process --:o7254
  (**) -- always_comb
  begin
    $axis_assert( "key_type1_line12b", std_logic'('0'), std_logic_vector'("10"),
     " ", " ", " ", " ", " ", " ", _zy_sva_key_type1_line12b_15_cpass, " ",
     _zy_sva_key_type1_line12b_15_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 1014,
     std_logic_vector'("000"));
  end process ;

  process --:o7255
  (**) -- always_comb
  begin
    $axis_assert( "key_type9_line14", std_logic'('0'), std_logic_vector'("10"),
     " ", " ", " ", " ", " ", " ", _zy_sva_key_type9_line14_16_cpass, " ",
     _zy_sva_key_type9_line14_16_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 1023,
     std_logic_vector'("000"));
  end process ;

  process --:o7256
  (**) -- always_comb
  begin
    $axis_assert( "key_type9_line15", std_logic'('0'), std_logic_vector'("10"),
     " ", " ", " ", " ", " ", " ", _zy_sva_key_type9_line15_17_cpass, " ",
     _zy_sva_key_type9_line15_17_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 1030,
     std_logic_vector'("000"));
  end process ;

  process --:o7257
  (**) -- always_comb
  begin
    $axis_assert( "key_type9_line16a", std_logic'('0'), std_logic_vector'("10"),
     " ", " ", " ", " ", " ", " ", _zy_sva_key_type9_line16a_18_cpass, " ",
     _zy_sva_key_type9_line16a_18_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 1036,
     std_logic_vector'("000"));
  end process ;

  process --:o7258
  (**) -- always_comb
  begin
    $axis_assert( "key_type9_line16b", std_logic'('0'), std_logic_vector'("10"),
     " ", " ", " ", " ", " ", " ", _zy_sva_key_type9_line16b_19_cpass, " ",
     _zy_sva_key_type9_line16b_19_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 1042,
     std_logic_vector'("000"));
  end process ;

  process --:o7259
  (**) -- always_comb
  begin
    $axis_assert( "key_type9_line17a", std_logic'('0'), std_logic_vector'("10"),
     " ", " ", " ", " ", " ", " ", _zy_sva_key_type9_line17a_20_cpass, " ",
     _zy_sva_key_type9_line17a_20_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 1050,
     std_logic_vector'("000"));
  end process ;

  process --:o7260
  (**) -- always_comb
  begin
    $axis_assert( "key_type9_line17b", std_logic'('0'), std_logic_vector'("10"),
     " ", " ", " ", " ", " ", " ", _zy_sva_key_type9_line17b_21_cpass, " ",
     _zy_sva_key_type9_line17b_21_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 1059,
     std_logic_vector'("000"));
  end process ;

  process --:o7261
  (**) -- always_comb
  begin
    $axis_assert( "key_type9_line18a", std_logic'('0'), std_logic_vector'("10"),
     " ", " ", " ", " ", " ", " ", _zy_sva_key_type9_line18a_22_cpass, " ",
     _zy_sva_key_type9_line18a_22_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 1066,
     std_logic_vector'("000"));
  end process ;

  process --:o7262
  (**) -- always_comb
  begin
    $axis_assert( "key_type9_line18b", std_logic'('0'), std_logic_vector'("10"),
     " ", " ", " ", " ", " ", " ", _zy_sva_key_type9_line18b_23_cpass, " ",
     _zy_sva_key_type9_line18b_23_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 1074,
     std_logic_vector'("000"));
  end process ;

  process --:o7263
  (**) -- always_comb
  begin
    $axis_assert( "key_type9_line19a", std_logic'('0'), std_logic_vector'("10"),
     " ", " ", " ", " ", " ", " ", _zy_sva_key_type9_line19a_24_cpass, " ",
     _zy_sva_key_type9_line19a_24_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 1081,
     std_logic_vector'("000"));
  end process ;

  process --:o7264
  (**) -- always_comb
  begin
    $axis_assert( "key_type9_line19b", std_logic'('0'), std_logic_vector'("10"),
     " ", " ", " ", " ", " ", " ", _zy_sva_key_type9_line19b_25_cpass, " ",
     _zy_sva_key_type9_line19b_25_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 1088,
     std_logic_vector'("000"));
  end process ;

  process --:o7265
  (**) -- always_comb
  begin
    $axis_assert( "key_type9_line19c", std_logic'('0'), std_logic_vector'("10"),
     " ", " ", " ", " ", " ", " ", _zy_sva_key_type9_line19c_26_cpass, " ",
     _zy_sva_key_type9_line19c_26_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 1094,
     std_logic_vector'("000"));
  end process ;

  process --:o7266
  (**) -- always_comb
  begin
    $axis_assert( "key_type9_line19d", std_logic'('0'), std_logic_vector'("10"),
     " ", " ", " ", " ", " ", " ", _zy_sva_key_type9_line19d_27_cpass, " ",
     _zy_sva_key_type9_line19d_27_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 1101,
     std_logic_vector'("000"));
  end process ;

  process --:o7267
  (**) -- always_comb
  begin
    $axis_assert( "guid_miss_aux_cmd_0", std_logic'('0'), std_logic_vector'("10"
    ), " ", " ", " ", " ", " ", " ", _zy_sva_guid_miss_aux_cmd_0_28_cpass, " ",
     _zy_sva_guid_miss_aux_cmd_0_28_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 1234,
     std_logic_vector'("000"));
  end process ;

  process --:o7268
  (**) -- always_comb
  begin
    $axis_assert( "guid_miss_aux_cmd_1", std_logic'('0'), std_logic_vector'("10"
    ), " ", " ", " ", " ", " ", " ", _zy_sva_guid_miss_aux_cmd_1_29_cpass, " ",
     _zy_sva_guid_miss_aux_cmd_1_29_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 1240,
     std_logic_vector'("000"));
  end process ;

  process --:o7269
  (**) -- always_comb
  begin
    $axis_assert( "guid_miss_aux_cmd_2", std_logic'('0'), std_logic_vector'("10"
    ), " ", " ", " ", " ", " ", " ", _zy_sva_guid_miss_aux_cmd_2_30_cpass, " ",
     _zy_sva_guid_miss_aux_cmd_2_30_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 1246,
     std_logic_vector'("000"));
  end process ;

  process --:o7270
  (**) -- always_comb
  begin
    $axis_assert( "guid_miss_aux_cmd_3", std_logic'('0'), std_logic_vector'("10"
    ), " ", " ", " ", " ", " ", " ", _zy_sva_guid_miss_aux_cmd_3_31_cpass, " ",
     _zy_sva_guid_miss_aux_cmd_3_31_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 1252,
     std_logic_vector'("000"));
  end process ;

  process --:o7271
  (**) -- always_comb
  begin
    $axis_assert( "guid_miss_aux_cmd_iv_0", std_logic'('0'), std_logic_vector'
    ("10"), " ", " ", " ", " ", " ", " ",
     _zy_sva_guid_miss_aux_cmd_iv_0_32_cpass, " ",
     _zy_sva_guid_miss_aux_cmd_iv_0_32_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 1258,
     std_logic_vector'("000"));
  end process ;

  process --:o7272
  (**) -- always_comb
  begin
    $axis_assert( "guid_miss_aux_cmd_iv_1", std_logic'('0'), std_logic_vector'
    ("10"), " ", " ", " ", " ", " ", " ",
     _zy_sva_guid_miss_aux_cmd_iv_1_33_cpass, " ",
     _zy_sva_guid_miss_aux_cmd_iv_1_33_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 1264,
     std_logic_vector'("000"));
  end process ;

  process --:o7273
  (**) -- always_comb
  begin
    $axis_assert( "guid_miss_aux_cmd_iv_2", std_logic'('0'), std_logic_vector'
    ("10"), " ", " ", " ", " ", " ", " ",
     _zy_sva_guid_miss_aux_cmd_iv_2_34_cpass, " ",
     _zy_sva_guid_miss_aux_cmd_iv_2_34_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 1270,
     std_logic_vector'("000"));
  end process ;

  process --:o7274
  (**) -- always_comb
  begin
    $axis_assert( "guid_miss_aux_cmd_iv_3", std_logic'('0'), std_logic_vector'
    ("10"), " ", " ", " ", " ", " ", " ",
     _zy_sva_guid_miss_aux_cmd_iv_3_35_cpass, " ",
     _zy_sva_guid_miss_aux_cmd_iv_3_35_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 1276,
     std_logic_vector'("000"));
  end process ;

  process --:o7275
  (**) -- always_comb
  begin
    $axis_assert( "iv_miss_aux_cmd_0", std_logic'('0'), std_logic_vector'("10"),
     " ", " ", " ", " ", " ", " ", _zy_sva_iv_miss_aux_cmd_0_36_cpass, " ",
     _zy_sva_iv_miss_aux_cmd_0_36_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 1282,
     std_logic_vector'("000"));
  end process ;

  process --:o7276
  (**) -- always_comb
  begin
    $axis_assert( "iv_miss_aux_cmd_1", std_logic'('0'), std_logic_vector'("10"),
     " ", " ", " ", " ", " ", " ", _zy_sva_iv_miss_aux_cmd_1_37_cpass, " ",
     _zy_sva_iv_miss_aux_cmd_1_37_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 1287,
     std_logic_vector'("000"));
  end process ;

  process --:o7277
  (**) -- always_comb
  begin
    $axis_assert( "iv_miss_aux_cmd_guid", std_logic'('0'), std_logic_vector'
    ("10"), " ", " ", " ", " ", " ", " ", _zy_sva_iv_miss_aux_cmd_guid_38_cpass,
     " ", _zy_sva_iv_miss_aux_cmd_guid_38_ccheck, " ",
     "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v", 1292,
     std_logic_vector'("000"));
  end process ;
end module;
