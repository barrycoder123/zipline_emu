library ieee, quickturn ;
use ieee.std_logic_1164.all ;
use quickturn.verilog.all ;
entity ifsyn_conns is
  attribute _2_state_: integer;
end ifsyn_conns ;
