library ieee, quickturn ;
use ieee.std_logic_1164.all ;
use quickturn.verilog.all ;
entity my_clks is
  attribute _2_state_: integer;
end my_clks ;
