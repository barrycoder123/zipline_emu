
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module AesSecIStub ( AesCiphOutR, AesCiphOutVldR, KeyInitStall, CiphInStall, 
	Aes128, Aes192, Aes256, CiphIn, CiphInVldR, CiphInLastR, EncryptEn, 
	KeyIn, KeyInitVldR, AesCiphOutStall, clk, rst_n);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output [127:0] AesCiphOutR;
output AesCiphOutVldR;
output KeyInitStall;
output CiphInStall;
input Aes128;
input Aes192;
input Aes256;
input [127:0] CiphIn;
input CiphInVldR;
input CiphInLastR;
input EncryptEn;
input [255:0] KeyIn;
input KeyInitVldR;
input AesCiphOutStall;
input clk;
input rst_n;
supply0 n1;
Q_BUF U0 ( .A(n1), .Z(AesCiphOutR[127]));
Q_BUF U1 ( .A(n1), .Z(AesCiphOutR[126]));
Q_BUF U2 ( .A(n1), .Z(AesCiphOutR[125]));
Q_BUF U3 ( .A(n1), .Z(AesCiphOutR[124]));
Q_BUF U4 ( .A(n1), .Z(AesCiphOutR[123]));
Q_BUF U5 ( .A(n1), .Z(AesCiphOutR[122]));
Q_BUF U6 ( .A(n1), .Z(AesCiphOutR[121]));
Q_BUF U7 ( .A(n1), .Z(AesCiphOutR[120]));
Q_BUF U8 ( .A(n1), .Z(AesCiphOutR[119]));
Q_BUF U9 ( .A(n1), .Z(AesCiphOutR[118]));
Q_BUF U10 ( .A(n1), .Z(AesCiphOutR[117]));
Q_BUF U11 ( .A(n1), .Z(AesCiphOutR[116]));
Q_BUF U12 ( .A(n1), .Z(AesCiphOutR[115]));
Q_BUF U13 ( .A(n1), .Z(AesCiphOutR[114]));
Q_BUF U14 ( .A(n1), .Z(AesCiphOutR[113]));
Q_BUF U15 ( .A(n1), .Z(AesCiphOutR[112]));
Q_BUF U16 ( .A(n1), .Z(AesCiphOutR[111]));
Q_BUF U17 ( .A(n1), .Z(AesCiphOutR[110]));
Q_BUF U18 ( .A(n1), .Z(AesCiphOutR[109]));
Q_BUF U19 ( .A(n1), .Z(AesCiphOutR[108]));
Q_BUF U20 ( .A(n1), .Z(AesCiphOutR[107]));
Q_BUF U21 ( .A(n1), .Z(AesCiphOutR[106]));
Q_BUF U22 ( .A(n1), .Z(AesCiphOutR[105]));
Q_BUF U23 ( .A(n1), .Z(AesCiphOutR[104]));
Q_BUF U24 ( .A(n1), .Z(AesCiphOutR[103]));
Q_BUF U25 ( .A(n1), .Z(AesCiphOutR[102]));
Q_BUF U26 ( .A(n1), .Z(AesCiphOutR[101]));
Q_BUF U27 ( .A(n1), .Z(AesCiphOutR[100]));
Q_BUF U28 ( .A(n1), .Z(AesCiphOutR[99]));
Q_BUF U29 ( .A(n1), .Z(AesCiphOutR[98]));
Q_BUF U30 ( .A(n1), .Z(AesCiphOutR[97]));
Q_BUF U31 ( .A(n1), .Z(AesCiphOutR[96]));
Q_BUF U32 ( .A(n1), .Z(AesCiphOutR[95]));
Q_BUF U33 ( .A(n1), .Z(AesCiphOutR[94]));
Q_BUF U34 ( .A(n1), .Z(AesCiphOutR[93]));
Q_BUF U35 ( .A(n1), .Z(AesCiphOutR[92]));
Q_BUF U36 ( .A(n1), .Z(AesCiphOutR[91]));
Q_BUF U37 ( .A(n1), .Z(AesCiphOutR[90]));
Q_BUF U38 ( .A(n1), .Z(AesCiphOutR[89]));
Q_BUF U39 ( .A(n1), .Z(AesCiphOutR[88]));
Q_BUF U40 ( .A(n1), .Z(AesCiphOutR[87]));
Q_BUF U41 ( .A(n1), .Z(AesCiphOutR[86]));
Q_BUF U42 ( .A(n1), .Z(AesCiphOutR[85]));
Q_BUF U43 ( .A(n1), .Z(AesCiphOutR[84]));
Q_BUF U44 ( .A(n1), .Z(AesCiphOutR[83]));
Q_BUF U45 ( .A(n1), .Z(AesCiphOutR[82]));
Q_BUF U46 ( .A(n1), .Z(AesCiphOutR[81]));
Q_BUF U47 ( .A(n1), .Z(AesCiphOutR[80]));
Q_BUF U48 ( .A(n1), .Z(AesCiphOutR[79]));
Q_BUF U49 ( .A(n1), .Z(AesCiphOutR[78]));
Q_BUF U50 ( .A(n1), .Z(AesCiphOutR[77]));
Q_BUF U51 ( .A(n1), .Z(AesCiphOutR[76]));
Q_BUF U52 ( .A(n1), .Z(AesCiphOutR[75]));
Q_BUF U53 ( .A(n1), .Z(AesCiphOutR[74]));
Q_BUF U54 ( .A(n1), .Z(AesCiphOutR[73]));
Q_BUF U55 ( .A(n1), .Z(AesCiphOutR[72]));
Q_BUF U56 ( .A(n1), .Z(AesCiphOutR[71]));
Q_BUF U57 ( .A(n1), .Z(AesCiphOutR[70]));
Q_BUF U58 ( .A(n1), .Z(AesCiphOutR[69]));
Q_BUF U59 ( .A(n1), .Z(AesCiphOutR[68]));
Q_BUF U60 ( .A(n1), .Z(AesCiphOutR[67]));
Q_BUF U61 ( .A(n1), .Z(AesCiphOutR[66]));
Q_BUF U62 ( .A(n1), .Z(AesCiphOutR[65]));
Q_BUF U63 ( .A(n1), .Z(AesCiphOutR[64]));
Q_BUF U64 ( .A(n1), .Z(AesCiphOutR[63]));
Q_BUF U65 ( .A(n1), .Z(AesCiphOutR[62]));
Q_BUF U66 ( .A(n1), .Z(AesCiphOutR[61]));
Q_BUF U67 ( .A(n1), .Z(AesCiphOutR[60]));
Q_BUF U68 ( .A(n1), .Z(AesCiphOutR[59]));
Q_BUF U69 ( .A(n1), .Z(AesCiphOutR[58]));
Q_BUF U70 ( .A(n1), .Z(AesCiphOutR[57]));
Q_BUF U71 ( .A(n1), .Z(AesCiphOutR[56]));
Q_BUF U72 ( .A(n1), .Z(AesCiphOutR[55]));
Q_BUF U73 ( .A(n1), .Z(AesCiphOutR[54]));
Q_BUF U74 ( .A(n1), .Z(AesCiphOutR[53]));
Q_BUF U75 ( .A(n1), .Z(AesCiphOutR[52]));
Q_BUF U76 ( .A(n1), .Z(AesCiphOutR[51]));
Q_BUF U77 ( .A(n1), .Z(AesCiphOutR[50]));
Q_BUF U78 ( .A(n1), .Z(AesCiphOutR[49]));
Q_BUF U79 ( .A(n1), .Z(AesCiphOutR[48]));
Q_BUF U80 ( .A(n1), .Z(AesCiphOutR[47]));
Q_BUF U81 ( .A(n1), .Z(AesCiphOutR[46]));
Q_BUF U82 ( .A(n1), .Z(AesCiphOutR[45]));
Q_BUF U83 ( .A(n1), .Z(AesCiphOutR[44]));
Q_BUF U84 ( .A(n1), .Z(AesCiphOutR[43]));
Q_BUF U85 ( .A(n1), .Z(AesCiphOutR[42]));
Q_BUF U86 ( .A(n1), .Z(AesCiphOutR[41]));
Q_BUF U87 ( .A(n1), .Z(AesCiphOutR[40]));
Q_BUF U88 ( .A(n1), .Z(AesCiphOutR[39]));
Q_BUF U89 ( .A(n1), .Z(AesCiphOutR[38]));
Q_BUF U90 ( .A(n1), .Z(AesCiphOutR[37]));
Q_BUF U91 ( .A(n1), .Z(AesCiphOutR[36]));
Q_BUF U92 ( .A(n1), .Z(AesCiphOutR[35]));
Q_BUF U93 ( .A(n1), .Z(AesCiphOutR[34]));
Q_BUF U94 ( .A(n1), .Z(AesCiphOutR[33]));
Q_BUF U95 ( .A(n1), .Z(AesCiphOutR[32]));
Q_BUF U96 ( .A(n1), .Z(AesCiphOutR[31]));
Q_BUF U97 ( .A(n1), .Z(AesCiphOutR[30]));
Q_BUF U98 ( .A(n1), .Z(AesCiphOutR[29]));
Q_BUF U99 ( .A(n1), .Z(AesCiphOutR[28]));
Q_BUF U100 ( .A(n1), .Z(AesCiphOutR[27]));
Q_BUF U101 ( .A(n1), .Z(AesCiphOutR[26]));
Q_BUF U102 ( .A(n1), .Z(AesCiphOutR[25]));
Q_BUF U103 ( .A(n1), .Z(AesCiphOutR[24]));
Q_BUF U104 ( .A(n1), .Z(AesCiphOutR[23]));
Q_BUF U105 ( .A(n1), .Z(AesCiphOutR[22]));
Q_BUF U106 ( .A(n1), .Z(AesCiphOutR[21]));
Q_BUF U107 ( .A(n1), .Z(AesCiphOutR[20]));
Q_BUF U108 ( .A(n1), .Z(AesCiphOutR[19]));
Q_BUF U109 ( .A(n1), .Z(AesCiphOutR[18]));
Q_BUF U110 ( .A(n1), .Z(AesCiphOutR[17]));
Q_BUF U111 ( .A(n1), .Z(AesCiphOutR[16]));
Q_BUF U112 ( .A(n1), .Z(AesCiphOutR[15]));
Q_BUF U113 ( .A(n1), .Z(AesCiphOutR[14]));
Q_BUF U114 ( .A(n1), .Z(AesCiphOutR[13]));
Q_BUF U115 ( .A(n1), .Z(AesCiphOutR[12]));
Q_BUF U116 ( .A(n1), .Z(AesCiphOutR[11]));
Q_BUF U117 ( .A(n1), .Z(AesCiphOutR[10]));
Q_BUF U118 ( .A(n1), .Z(AesCiphOutR[9]));
Q_BUF U119 ( .A(n1), .Z(AesCiphOutR[8]));
Q_BUF U120 ( .A(n1), .Z(AesCiphOutR[7]));
Q_BUF U121 ( .A(n1), .Z(AesCiphOutR[6]));
Q_BUF U122 ( .A(n1), .Z(AesCiphOutR[5]));
Q_BUF U123 ( .A(n1), .Z(AesCiphOutR[4]));
Q_BUF U124 ( .A(n1), .Z(AesCiphOutR[3]));
Q_BUF U125 ( .A(n1), .Z(AesCiphOutR[2]));
Q_BUF U126 ( .A(n1), .Z(AesCiphOutR[1]));
Q_BUF U127 ( .A(n1), .Z(AesCiphOutR[0]));
Q_BUF U128 ( .A(n1), .Z(KeyInitStall));
Q_BUF U129 ( .A(n1), .Z(CiphInStall));
Q_INV U130 ( .A(AesCiphOutStall), .Z(AesCiphOutVldR));
endmodule
