
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
(* celldefine = 1 *) 
module nx_indirect_access_cntrl_xcm113 ( clk, rst_n, wr_stb, reg_addr, cmnd_op, 
	cmnd_addr, cmnd_table_id, stat_code, stat_datawords, stat_addr, 
	stat_table_id, capability_lst, capability_type, enable, .addr_limit( {
	\addr_limit[0][8] , \addr_limit[0][7] , \addr_limit[0][6] , 
	\addr_limit[0][5] , \addr_limit[0][4] , \addr_limit[0][3] , 
	\addr_limit[0][2] , \addr_limit[0][1] , \addr_limit[0][0] } ), 
	wr_dat, rd_dat, sw_cs, sw_ce, sw_we, sw_add, sw_wdat, sw_rdat, 
	sw_match, sw_aindex, grant, yield, reset);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
input clk;
input rst_n;
input wr_stb;
input [10:0] reg_addr;
input [3:0] cmnd_op;
input [8:0] cmnd_addr;
input [0:0] cmnd_table_id;
output [2:0] stat_code;
output [4:0] stat_datawords;
output [8:0] stat_addr;
output [0:0] stat_table_id;
output [15:0] capability_lst;
output [3:0] capability_type;
output enable;
input \addr_limit[0][8] ;
input \addr_limit[0][7] ;
input \addr_limit[0][6] ;
input \addr_limit[0][5] ;
input \addr_limit[0][4] ;
input \addr_limit[0][3] ;
input \addr_limit[0][2] ;
input \addr_limit[0][1] ;
input \addr_limit[0][0] ;
input [95:0] wr_dat;
output [95:0] rd_dat;
output sw_cs;
output sw_ce;
output sw_we;
output [8:0] sw_add;
output [95:0] sw_wdat;
input [95:0] sw_rdat;
input sw_match;
input [7:0] sw_aindex;
input grant;
output yield;
output reset;
wire [0:2] _zy_simnet_stat_code_0_w$;
wire [0:4] _zy_simnet_stat_datawords_1_w$;
wire [0:8] _zy_simnet_stat_addr_2_w$;
wire _zy_simnet_stat_table_id_3_w$;
wire [0:15] _zy_simnet_capability_lst_4_w$;
wire [0:3] _zy_simnet_capability_type_5_w$;
wire _zy_simnet_enable_6_w$;
wire [0:95] _zy_simnet_rd_dat_7_w$;
wire _zy_simnet_sw_cs_8_w$;
wire _zy_simnet_sw_ce_9_w$;
wire _zy_simnet_sw_we_10_w$;
wire [0:8] _zy_simnet_sw_add_11_w$;
wire [0:95] _zy_simnet_sw_wdat_12_w$;
wire _zy_simnet_yield_13_w$;
wire _zy_simnet_reset_14_w$;
wire [3:0] cmnd;
wire init_r;
wire [0:0] inc_r;
wire init_inc_r;
wire sw_cs_r;
wire sw_ce_r;
wire rst_r;
wire rst_or_ini_r;
wire [8:0] rst_addr_r;
wire sw_we_r;
wire cmnd_rd_stb;
wire cmnd_wr_stb;
wire cmnd_ena_stb;
wire cmnd_dis_stb;
wire cmnd_rst_stb;
wire cmnd_ini_stb;
wire cmnd_inc_stb;
wire cmnd_sis_stb;
wire cmnd_tmo_stb;
wire cmnd_cmp_stb;
wire cmnd_issued;
wire ack_error;
wire unsupported_op;
wire [3:0] state_r;
wire [5:0] timer_r;
wire timeout;
wire sim_tmo_r;
wire [8:0] maxaddr;
wire badaddr;
wire igrant;
wire [2:0] stat;
supply0 n1;
supply1 n2;
Q_BUF U0 ( .A(n1), .Z(stat_datawords[0]));
Q_BUF U1 ( .A(n2), .Z(stat_datawords[1]));
Q_BUF U2 ( .A(n1), .Z(stat_datawords[2]));
Q_BUF U3 ( .A(n1), .Z(stat_datawords[3]));
Q_BUF U4 ( .A(n1), .Z(stat_datawords[4]));
Q_BUF U5 ( .A(n1), .Z(capability_type[0]));
Q_BUF U6 ( .A(n1), .Z(capability_type[1]));
Q_BUF U7 ( .A(n1), .Z(capability_type[2]));
Q_BUF U8 ( .A(n1), .Z(capability_type[3]));
Q_BUF U9 ( .A(n2), .Z(capability_lst[0]));
Q_BUF U10 ( .A(n2), .Z(capability_lst[1]));
Q_BUF U11 ( .A(n2), .Z(capability_lst[2]));
Q_BUF U12 ( .A(n2), .Z(capability_lst[3]));
Q_BUF U13 ( .A(n2), .Z(capability_lst[4]));
Q_BUF U14 ( .A(n2), .Z(capability_lst[5]));
Q_BUF U15 ( .A(n2), .Z(capability_lst[6]));
Q_BUF U16 ( .A(n1), .Z(capability_lst[7]));
Q_BUF U17 ( .A(n2), .Z(capability_lst[8]));
Q_BUF U18 ( .A(n1), .Z(capability_lst[9]));
Q_BUF U19 ( .A(n1), .Z(capability_lst[10]));
Q_BUF U20 ( .A(n1), .Z(capability_lst[11]));
Q_BUF U21 ( .A(n1), .Z(capability_lst[12]));
Q_BUF U22 ( .A(n1), .Z(capability_lst[13]));
Q_BUF U23 ( .A(n2), .Z(capability_lst[14]));
Q_BUF U24 ( .A(n2), .Z(capability_lst[15]));
Q_BUF U25 ( .A(n1), .Z(stat_table_id[0]));
ixc_assign_3 _zz_strnp_7 ( stat[2:0], stat_code[2:0]);
ixc_assign_4 _zz_strnp_1 ( cmnd[3:0], cmnd_op[3:0]);
ixc_assign \genblk1._zz_strnp_0 ( reset, rst_or_ini_r);
ixc_context_read_6 _zzixc_ctxrd_0 ( { stat_code[2], stat_code[1], 
	stat_code[0], stat[2], stat[1], stat[0]});
ixc_assign _zz_strnp_22 ( _zy_simnet_reset_14_w$, reset);
ixc_assign _zz_strnp_21 ( _zy_simnet_yield_13_w$, yield);
ixc_assign_96 _zz_strnp_20 ( _zy_simnet_sw_wdat_12_w$[0:95], sw_wdat[95:0]);
ixc_assign_9 _zz_strnp_19 ( _zy_simnet_sw_add_11_w$[0:8], sw_add[8:0]);
ixc_assign _zz_strnp_18 ( _zy_simnet_sw_we_10_w$, sw_we);
ixc_assign _zz_strnp_17 ( _zy_simnet_sw_ce_9_w$, sw_ce);
ixc_assign _zz_strnp_16 ( _zy_simnet_sw_cs_8_w$, sw_cs);
ixc_assign_96 _zz_strnp_15 ( _zy_simnet_rd_dat_7_w$[0:95], rd_dat[95:0]);
ixc_assign _zz_strnp_14 ( _zy_simnet_enable_6_w$, enable);
ixc_assign_4 _zz_strnp_13 ( _zy_simnet_capability_type_5_w$[0:3], { n1, n1, 
	n1, n1});
ixc_assign_16 _zz_strnp_12 ( _zy_simnet_capability_lst_4_w$[0:15], { n2, n2, 
	n1, n1, n1, n1, n1, n2, n1, n2, n2, n2, n2, n2, n2, n2});
ixc_assign _zz_strnp_11 ( _zy_simnet_stat_table_id_3_w$, n1);
ixc_assign_9 _zz_strnp_10 ( _zy_simnet_stat_addr_2_w$[0:8], stat_addr[8:0]);
ixc_assign_5 _zz_strnp_9 ( _zy_simnet_stat_datawords_1_w$[0:4], { n1, n1, n1, 
	n2, n1});
ixc_assign_3 _zz_strnp_8 ( _zy_simnet_stat_code_0_w$[0:2], stat_code[2:0]);
ixc_assign_9 _zz_strnp_6 ( stat_addr[8:0], maxaddr[8:0]);
Q_AN02 U46 ( .A0(n36), .A1(grant), .Z(igrant));
Q_AN02 U47 ( .A0(cmnd_issued), .A1(n35), .Z(badaddr));
Q_OR03 U48 ( .A0(n16), .A1(n34), .A2(n33), .Z(n35));
Q_AN02 U49 ( .A0(n17), .A1(n29), .Z(n34));
Q_AN02 U50 ( .A0(n17), .A1(n30), .Z(n32));
Q_AN03 U51 ( .A0(cmnd_addr[0]), .A1(n31), .A2(n32), .Z(n33));
Q_INV U52 ( .A(maxaddr[0]), .Z(n31));
Q_OR03 U53 ( .A0(n26), .A1(n25), .A2(n28), .Z(n29));
Q_OA21 U54 ( .A0(cmnd_addr[1]), .A1(n22), .B0(n24), .Z(n30));
Q_AN03 U55 ( .A0(cmnd_addr[1]), .A1(n22), .A2(n24), .Z(n25));
Q_INV U56 ( .A(maxaddr[1]), .Z(n22));
Q_OA21 U57 ( .A0(cmnd_addr[2]), .A1(n21), .B0(n23), .Z(n24));
Q_AN03 U58 ( .A0(cmnd_addr[2]), .A1(n21), .A2(n23), .Z(n26));
Q_INV U59 ( .A(maxaddr[2]), .Z(n21));
Q_OA21 U60 ( .A0(cmnd_addr[3]), .A1(n20), .B0(n19), .Z(n23));
Q_AN03 U61 ( .A0(cmnd_addr[3]), .A1(n20), .A2(n19), .Z(n27));
Q_INV U62 ( .A(maxaddr[3]), .Z(n20));
Q_OR02 U63 ( .A0(cmnd_addr[4]), .A1(n18), .Z(n19));
Q_AO21 U64 ( .A0(cmnd_addr[4]), .A1(n18), .B0(n27), .Z(n28));
Q_INV U65 ( .A(maxaddr[4]), .Z(n18));
Q_OR03 U66 ( .A0(n13), .A1(n12), .A2(n15), .Z(n16));
Q_OA21 U67 ( .A0(cmnd_addr[5]), .A1(n9), .B0(n11), .Z(n17));
Q_AN03 U68 ( .A0(cmnd_addr[5]), .A1(n9), .A2(n11), .Z(n12));
Q_INV U69 ( .A(maxaddr[5]), .Z(n9));
Q_OA21 U70 ( .A0(cmnd_addr[6]), .A1(n8), .B0(n10), .Z(n11));
Q_AN03 U71 ( .A0(cmnd_addr[6]), .A1(n8), .A2(n10), .Z(n13));
Q_INV U72 ( .A(maxaddr[6]), .Z(n8));
Q_OA21 U73 ( .A0(cmnd_addr[7]), .A1(n7), .B0(n6), .Z(n10));
Q_AN03 U74 ( .A0(cmnd_addr[7]), .A1(n7), .A2(n6), .Z(n14));
Q_INV U75 ( .A(maxaddr[7]), .Z(n7));
Q_OR02 U76 ( .A0(cmnd_addr[8]), .A1(n5), .Z(n6));
Q_AO21 U77 ( .A0(cmnd_addr[8]), .A1(n5), .B0(n14), .Z(n15));
Q_INV U78 ( .A(maxaddr[8]), .Z(n5));
Q_AN02 U79 ( .A0(n3), .A1(n4), .Z(timeout));
Q_AN03 U80 ( .A0(timer_r[2]), .A1(timer_r[1]), .A2(timer_r[0]), .Z(n4));
Q_AN03 U81 ( .A0(timer_r[5]), .A1(timer_r[4]), .A2(timer_r[3]), .Z(n3));
ixc_assign _zz_strnp_5 ( yield, timer_r[5]);
ixc_assign _zz_strnp_4 ( sw_we, sw_we_r);
ixc_assign _zz_strnp_3 ( sw_ce, sw_ce_r);
ixc_assign _zz_strnp_2 ( sw_cs, sw_cs_r);
Q_MX02 U86 ( .S(rst_or_ini_r), .A0(cmnd_addr[0]), .A1(rst_addr_r[0]), .Z(sw_add[0]));
Q_MX02 U87 ( .S(rst_or_ini_r), .A0(cmnd_addr[1]), .A1(rst_addr_r[1]), .Z(sw_add[1]));
Q_MX02 U88 ( .S(rst_or_ini_r), .A0(cmnd_addr[2]), .A1(rst_addr_r[2]), .Z(sw_add[2]));
Q_MX02 U89 ( .S(rst_or_ini_r), .A0(cmnd_addr[3]), .A1(rst_addr_r[3]), .Z(sw_add[3]));
Q_MX02 U90 ( .S(rst_or_ini_r), .A0(cmnd_addr[4]), .A1(rst_addr_r[4]), .Z(sw_add[4]));
Q_MX02 U91 ( .S(rst_or_ini_r), .A0(cmnd_addr[5]), .A1(rst_addr_r[5]), .Z(sw_add[5]));
Q_MX02 U92 ( .S(rst_or_ini_r), .A0(cmnd_addr[6]), .A1(rst_addr_r[6]), .Z(sw_add[6]));
Q_MX02 U93 ( .S(rst_or_ini_r), .A0(cmnd_addr[7]), .A1(rst_addr_r[7]), .Z(sw_add[7]));
Q_MX02 U94 ( .S(rst_or_ini_r), .A0(cmnd_addr[8]), .A1(rst_addr_r[8]), .Z(sw_add[8]));
Q_AN02 U95 ( .A0(enable), .A1(\addr_limit[0][0] ), .Z(maxaddr[0]));
Q_AN02 U96 ( .A0(enable), .A1(\addr_limit[0][1] ), .Z(maxaddr[1]));
Q_AN02 U97 ( .A0(enable), .A1(\addr_limit[0][2] ), .Z(maxaddr[2]));
Q_AN02 U98 ( .A0(enable), .A1(\addr_limit[0][3] ), .Z(maxaddr[3]));
Q_AN02 U99 ( .A0(enable), .A1(\addr_limit[0][4] ), .Z(maxaddr[4]));
Q_AN02 U100 ( .A0(enable), .A1(\addr_limit[0][5] ), .Z(maxaddr[5]));
Q_AN02 U101 ( .A0(enable), .A1(\addr_limit[0][6] ), .Z(maxaddr[6]));
Q_AN02 U102 ( .A0(enable), .A1(\addr_limit[0][7] ), .Z(maxaddr[7]));
Q_AN02 U103 ( .A0(enable), .A1(\addr_limit[0][8] ), .Z(maxaddr[8]));
Q_INV U104 ( .A(reg_addr[4]), .Z(n37));
Q_INV U105 ( .A(reg_addr[5]), .Z(n38));
Q_INV U106 ( .A(reg_addr[6]), .Z(n39));
Q_INV U107 ( .A(reg_addr[8]), .Z(n40));
Q_OR03 U108 ( .A0(reg_addr[10]), .A1(reg_addr[9]), .A2(n40), .Z(n41));
Q_OR03 U109 ( .A0(reg_addr[7]), .A1(n39), .A2(n38), .Z(n42));
Q_OR03 U110 ( .A0(n37), .A1(reg_addr[3]), .A2(reg_addr[2]), .Z(n43));
Q_OR03 U111 ( .A0(reg_addr[1]), .A1(reg_addr[0]), .A2(n41), .Z(n44));
Q_NR03 U112 ( .A0(n42), .A1(n43), .A2(n44), .Z(n45));
Q_AN02 U113 ( .A0(wr_stb), .A1(n45), .Z(n69));
Q_INV U114 ( .A(n64), .Z(cmnd_issued));
Q_INV U115 ( .A(unsupported_op), .Z(n63));
Q_OA21 U116 ( .A0(n47), .A1(n48), .B0(n46), .Z(unsupported_op));
Q_AN02 U117 ( .A0(n46), .A1(n49), .Z(ack_error));
Q_AO21 U118 ( .A0(n51), .A1(n52), .B0(n50), .Z(n64));
Q_INV U119 ( .A(n69), .Z(n50));
Q_MX02 U120 ( .S(cmnd[3]), .A0(n55), .A1(n53), .Z(n51));
Q_INV U121 ( .A(cmnd_cmp_stb), .Z(n65));
Q_AN02 U122 ( .A0(n46), .A1(n56), .Z(cmnd_cmp_stb));
Q_AN02 U123 ( .A0(n46), .A1(n57), .Z(cmnd_tmo_stb));
Q_AN03 U124 ( .A0(n46), .A1(n52), .A2(n55), .Z(cmnd_sis_stb));
Q_AN02 U125 ( .A0(n69), .A1(cmnd[3]), .Z(n46));
Q_AN02 U126 ( .A0(n58), .A1(n49), .Z(cmnd_inc_stb));
Q_AN02 U127 ( .A0(n53), .A1(cmnd[0]), .Z(n49));
Q_AN02 U128 ( .A0(n58), .A1(n57), .Z(cmnd_ini_stb));
Q_AN02 U129 ( .A0(n53), .A1(n52), .Z(n57));
Q_AN02 U130 ( .A0(cmnd[2]), .A1(cmnd[1]), .Z(n53));
Q_INV U131 ( .A(cmnd_rst_stb), .Z(n66));
Q_AN02 U132 ( .A0(n48), .A1(n59), .Z(cmnd_rst_stb));
Q_AN02 U133 ( .A0(n58), .A1(cmnd[0]), .Z(n59));
Q_AN02 U134 ( .A0(n48), .A1(n60), .Z(cmnd_dis_stb));
Q_AN02 U135 ( .A0(n58), .A1(n52), .Z(n60));
Q_AN02 U136 ( .A0(cmnd[2]), .A1(n61), .Z(n48));
Q_AN02 U137 ( .A0(n47), .A1(n59), .Z(cmnd_ena_stb));
Q_INV U138 ( .A(cmnd_wr_stb), .Z(n67));
Q_AN02 U139 ( .A0(n47), .A1(n60), .Z(cmnd_wr_stb));
Q_INV U140 ( .A(cmnd[0]), .Z(n52));
Q_AN02 U141 ( .A0(n62), .A1(cmnd[1]), .Z(n47));
Q_INV U142 ( .A(cmnd_rd_stb), .Z(n68));
Q_AN02 U143 ( .A0(n58), .A1(n56), .Z(cmnd_rd_stb));
Q_AN02 U144 ( .A0(n55), .A1(cmnd[0]), .Z(n56));
Q_NR02 U145 ( .A0(cmnd[2]), .A1(cmnd[1]), .Z(n55));
Q_INV U146 ( .A(cmnd[1]), .Z(n61));
Q_INV U147 ( .A(cmnd[2]), .Z(n62));
Q_AN02 U148 ( .A0(n69), .A1(n54), .Z(n58));
Q_INV U149 ( .A(cmnd[3]), .Z(n54));
Q_OR02 U150 ( .A0(cmnd_ini_stb), .A1(cmnd_inc_stb), .Z(n517));
Q_XNR2 U151 ( .A0(rst_addr_r[0]), .A1(maxaddr[0]), .Z(n70));
Q_XNR2 U152 ( .A0(rst_addr_r[1]), .A1(maxaddr[1]), .Z(n71));
Q_XNR2 U153 ( .A0(rst_addr_r[2]), .A1(maxaddr[2]), .Z(n72));
Q_XNR2 U154 ( .A0(rst_addr_r[3]), .A1(maxaddr[3]), .Z(n73));
Q_XNR2 U155 ( .A0(rst_addr_r[4]), .A1(maxaddr[4]), .Z(n74));
Q_XNR2 U156 ( .A0(rst_addr_r[5]), .A1(maxaddr[5]), .Z(n75));
Q_XNR2 U157 ( .A0(rst_addr_r[6]), .A1(maxaddr[6]), .Z(n76));
Q_XNR2 U158 ( .A0(rst_addr_r[7]), .A1(maxaddr[7]), .Z(n77));
Q_XNR2 U159 ( .A0(rst_addr_r[8]), .A1(maxaddr[8]), .Z(n78));
Q_AN03 U160 ( .A0(n78), .A1(n77), .A2(n76), .Z(n79));
Q_AN03 U161 ( .A0(n75), .A1(n74), .A2(n73), .Z(n80));
Q_AN03 U162 ( .A0(n72), .A1(n71), .A2(n70), .Z(n81));
Q_AN03 U163 ( .A0(n79), .A1(n80), .A2(n81), .Z(n518));
Q_XNR2 U164 ( .A0(rst_addr_r[0]), .A1(cmnd_addr[0]), .Z(n82));
Q_XNR2 U165 ( .A0(rst_addr_r[1]), .A1(cmnd_addr[1]), .Z(n83));
Q_XNR2 U166 ( .A0(rst_addr_r[2]), .A1(cmnd_addr[2]), .Z(n84));
Q_XNR2 U167 ( .A0(rst_addr_r[3]), .A1(cmnd_addr[3]), .Z(n85));
Q_XNR2 U168 ( .A0(rst_addr_r[4]), .A1(cmnd_addr[4]), .Z(n86));
Q_XNR2 U169 ( .A0(rst_addr_r[5]), .A1(cmnd_addr[5]), .Z(n87));
Q_XNR2 U170 ( .A0(rst_addr_r[6]), .A1(cmnd_addr[6]), .Z(n88));
Q_XNR2 U171 ( .A0(rst_addr_r[7]), .A1(cmnd_addr[7]), .Z(n89));
Q_XNR2 U172 ( .A0(rst_addr_r[8]), .A1(cmnd_addr[8]), .Z(n90));
Q_AN03 U173 ( .A0(n90), .A1(n89), .A2(n88), .Z(n91));
Q_AN03 U174 ( .A0(n87), .A1(n86), .A2(n85), .Z(n92));
Q_AN03 U175 ( .A0(n84), .A1(n83), .A2(n82), .Z(n93));
Q_AN03 U176 ( .A0(n91), .A1(n92), .A2(n93), .Z(n519));
Q_AN02 U177 ( .A0(init_inc_r), .A1(igrant), .Z(n94));
Q_XOR2 U178 ( .A0(inc_r[0]), .A1(n94), .Z(n95));
Q_AD01HF U179 ( .A0(rst_addr_r[0]), .B0(igrant), .S(n96), .CO(n97));
Q_AD01HF U180 ( .A0(rst_addr_r[1]), .B0(n97), .S(n98), .CO(n99));
Q_AD01HF U181 ( .A0(rst_addr_r[2]), .B0(n99), .S(n100), .CO(n101));
Q_AD01HF U182 ( .A0(rst_addr_r[3]), .B0(n101), .S(n102), .CO(n103));
Q_AD01HF U183 ( .A0(rst_addr_r[4]), .B0(n103), .S(n104), .CO(n105));
Q_AD01HF U184 ( .A0(rst_addr_r[5]), .B0(n105), .S(n106), .CO(n107));
Q_AD01HF U185 ( .A0(rst_addr_r[6]), .B0(n107), .S(n108), .CO(n109));
Q_AD01HF U186 ( .A0(rst_addr_r[7]), .B0(n109), .S(n110), .CO(n111));
Q_XOR2 U187 ( .A0(rst_addr_r[8]), .A1(n111), .Z(n112));
Q_AD01HF U188 ( .A0(timer_r[1]), .B0(timer_r[0]), .S(n114), .CO(n115));
Q_AD01HF U189 ( .A0(timer_r[2]), .B0(n115), .S(n116), .CO(n117));
Q_AD01HF U190 ( .A0(timer_r[3]), .B0(n117), .S(n118), .CO(n119));
Q_AD01HF U191 ( .A0(timer_r[4]), .B0(n119), .S(n120), .CO(n121));
Q_XOR2 U192 ( .A0(timer_r[5]), .A1(n121), .Z(n122));
Q_MX02 U193 ( .S(n436), .A0(n128), .A1(n124), .Z(n123));
Q_ND02 U194 ( .A0(n125), .A1(n126), .Z(n124));
Q_ND02 U195 ( .A0(n494), .A1(n400), .Z(n126));
Q_OR02 U196 ( .A0(n127), .A1(n400), .Z(n125));
Q_OR02 U197 ( .A0(n400), .A1(n496), .Z(n128));
Q_INV U198 ( .A(n129), .Z(n130));
Q_MX02 U199 ( .S(n436), .A0(n125), .A1(n131), .Z(n129));
Q_INV U200 ( .A(n132), .Z(n131));
Q_INV U201 ( .A(n133), .Z(n134));
Q_MX02 U202 ( .S(n436), .A0(n140), .A1(n135), .Z(n133));
Q_INV U203 ( .A(n136), .Z(n135));
Q_MX02 U204 ( .S(n400), .A0(n132), .A1(n137), .Z(n136));
Q_INV U205 ( .A(n138), .Z(n137));
Q_XOR2 U206 ( .A0(n494), .A1(n139), .Z(n132));
Q_OR02 U207 ( .A0(n495), .A1(n127), .Z(n140));
Q_OR02 U208 ( .A0(n494), .A1(n496), .Z(n127));
Q_NR02 U209 ( .A0(n497), .A1(n142), .Z(n141));
Q_MX02 U210 ( .S(n400), .A0(n138), .A1(n496), .Z(n142));
Q_OR02 U211 ( .A0(n494), .A1(n139), .Z(n138));
Q_INV U212 ( .A(n496), .Z(n139));
Q_AN03 U213 ( .A0(n495), .A1(n494), .A2(n497), .Z(n143));
Q_AO21 U214 ( .A0(n143), .A1(state_r[3]), .B0(n141), .Z(n523));
Q_AO21 U215 ( .A0(n143), .A1(state_r[2]), .B0(n134), .Z(n522));
Q_AO21 U216 ( .A0(n143), .A1(state_r[1]), .B0(n130), .Z(n521));
Q_AO21 U217 ( .A0(n143), .A1(state_r[0]), .B0(n123), .Z(n520));
Q_AN02 U218 ( .A0(n498), .A1(n113), .Z(n144));
Q_AN02 U219 ( .A0(n498), .A1(n114), .Z(n145));
Q_AN02 U220 ( .A0(n498), .A1(n116), .Z(n146));
Q_AN02 U221 ( .A0(n498), .A1(n118), .Z(n147));
Q_AN02 U222 ( .A0(n498), .A1(n120), .Z(n148));
Q_AN02 U223 ( .A0(n498), .A1(n122), .Z(n149));
Q_AN02 U224 ( .A0(n500), .A1(cmnd_addr[0]), .Z(n150));
Q_MX02 U225 ( .S(n501), .A0(n150), .A1(n96), .Z(n151));
Q_AN02 U226 ( .A0(n500), .A1(cmnd_addr[1]), .Z(n152));
Q_MX02 U227 ( .S(n501), .A0(n152), .A1(n98), .Z(n153));
Q_AN02 U228 ( .A0(n500), .A1(cmnd_addr[2]), .Z(n154));
Q_MX02 U229 ( .S(n501), .A0(n154), .A1(n100), .Z(n155));
Q_AN02 U230 ( .A0(n500), .A1(cmnd_addr[3]), .Z(n156));
Q_MX02 U231 ( .S(n501), .A0(n156), .A1(n102), .Z(n157));
Q_AN02 U232 ( .A0(n500), .A1(cmnd_addr[4]), .Z(n158));
Q_MX02 U233 ( .S(n501), .A0(n158), .A1(n104), .Z(n159));
Q_AN02 U234 ( .A0(n500), .A1(cmnd_addr[5]), .Z(n160));
Q_MX02 U235 ( .S(n501), .A0(n160), .A1(n106), .Z(n161));
Q_AN02 U236 ( .A0(n500), .A1(cmnd_addr[6]), .Z(n162));
Q_MX02 U237 ( .S(n501), .A0(n162), .A1(n108), .Z(n163));
Q_AN02 U238 ( .A0(n500), .A1(cmnd_addr[7]), .Z(n164));
Q_MX02 U239 ( .S(n501), .A0(n164), .A1(n110), .Z(n165));
Q_AN02 U240 ( .A0(n500), .A1(cmnd_addr[8]), .Z(n166));
Q_MX02 U241 ( .S(n501), .A0(n166), .A1(n112), .Z(n167));
Q_AN02 U242 ( .A0(n506), .A1(n95), .Z(n168));
Q_MX03 U243 ( .S0(n508), .S1(n509), .A0(sw_aindex[0]), .A1(wr_dat[0]), .A2(sw_rdat[0]), .Z(n169));
Q_MX03 U244 ( .S0(n508), .S1(n509), .A0(sw_aindex[1]), .A1(wr_dat[1]), .A2(sw_rdat[1]), .Z(n170));
Q_MX03 U245 ( .S0(n508), .S1(n509), .A0(sw_aindex[2]), .A1(wr_dat[2]), .A2(sw_rdat[2]), .Z(n171));
Q_MX03 U246 ( .S0(n508), .S1(n509), .A0(sw_aindex[3]), .A1(wr_dat[3]), .A2(sw_rdat[3]), .Z(n172));
Q_MX03 U247 ( .S0(n508), .S1(n509), .A0(sw_aindex[4]), .A1(wr_dat[4]), .A2(sw_rdat[4]), .Z(n173));
Q_MX03 U248 ( .S0(n508), .S1(n509), .A0(sw_aindex[5]), .A1(wr_dat[5]), .A2(sw_rdat[5]), .Z(n174));
Q_MX03 U249 ( .S0(n508), .S1(n509), .A0(sw_aindex[6]), .A1(wr_dat[6]), .A2(sw_rdat[6]), .Z(n175));
Q_MX03 U250 ( .S0(n508), .S1(n509), .A0(sw_aindex[7]), .A1(wr_dat[7]), .A2(sw_rdat[7]), .Z(n176));
Q_MX03 U251 ( .S0(n508), .S1(n509), .A0(sw_match), .A1(wr_dat[8]), .A2(sw_rdat[8]), .Z(n177));
Q_AN02 U252 ( .A0(n508), .A1(wr_dat[9]), .Z(n178));
Q_MX02 U253 ( .S(n509), .A0(n178), .A1(sw_rdat[9]), .Z(n179));
Q_AN02 U254 ( .A0(n508), .A1(wr_dat[10]), .Z(n180));
Q_MX02 U255 ( .S(n509), .A0(n180), .A1(sw_rdat[10]), .Z(n181));
Q_AN02 U256 ( .A0(n508), .A1(wr_dat[11]), .Z(n182));
Q_MX02 U257 ( .S(n509), .A0(n182), .A1(sw_rdat[11]), .Z(n183));
Q_AN02 U258 ( .A0(n508), .A1(wr_dat[12]), .Z(n184));
Q_MX02 U259 ( .S(n509), .A0(n184), .A1(sw_rdat[12]), .Z(n185));
Q_AN02 U260 ( .A0(n508), .A1(wr_dat[13]), .Z(n186));
Q_MX02 U261 ( .S(n509), .A0(n186), .A1(sw_rdat[13]), .Z(n187));
Q_AN02 U262 ( .A0(n508), .A1(wr_dat[14]), .Z(n188));
Q_MX02 U263 ( .S(n509), .A0(n188), .A1(sw_rdat[14]), .Z(n189));
Q_AN02 U264 ( .A0(n508), .A1(wr_dat[15]), .Z(n190));
Q_MX02 U265 ( .S(n509), .A0(n190), .A1(sw_rdat[15]), .Z(n191));
Q_AN02 U266 ( .A0(n508), .A1(wr_dat[16]), .Z(n192));
Q_MX02 U267 ( .S(n509), .A0(n192), .A1(sw_rdat[16]), .Z(n193));
Q_AN02 U268 ( .A0(n508), .A1(wr_dat[17]), .Z(n194));
Q_MX02 U269 ( .S(n509), .A0(n194), .A1(sw_rdat[17]), .Z(n195));
Q_AN02 U270 ( .A0(n508), .A1(wr_dat[18]), .Z(n196));
Q_MX02 U271 ( .S(n509), .A0(n196), .A1(sw_rdat[18]), .Z(n197));
Q_AN02 U272 ( .A0(n508), .A1(wr_dat[19]), .Z(n198));
Q_MX02 U273 ( .S(n509), .A0(n198), .A1(sw_rdat[19]), .Z(n199));
Q_AN02 U274 ( .A0(n508), .A1(wr_dat[20]), .Z(n200));
Q_MX02 U275 ( .S(n509), .A0(n200), .A1(sw_rdat[20]), .Z(n201));
Q_AN02 U276 ( .A0(n508), .A1(wr_dat[21]), .Z(n202));
Q_MX02 U277 ( .S(n509), .A0(n202), .A1(sw_rdat[21]), .Z(n203));
Q_AN02 U278 ( .A0(n508), .A1(wr_dat[22]), .Z(n204));
Q_MX02 U279 ( .S(n509), .A0(n204), .A1(sw_rdat[22]), .Z(n205));
Q_AN02 U280 ( .A0(n508), .A1(wr_dat[23]), .Z(n206));
Q_MX02 U281 ( .S(n509), .A0(n206), .A1(sw_rdat[23]), .Z(n207));
Q_AN02 U282 ( .A0(n508), .A1(wr_dat[24]), .Z(n208));
Q_MX02 U283 ( .S(n509), .A0(n208), .A1(sw_rdat[24]), .Z(n209));
Q_AN02 U284 ( .A0(n508), .A1(wr_dat[25]), .Z(n210));
Q_MX02 U285 ( .S(n509), .A0(n210), .A1(sw_rdat[25]), .Z(n211));
Q_AN02 U286 ( .A0(n508), .A1(wr_dat[26]), .Z(n212));
Q_MX02 U287 ( .S(n509), .A0(n212), .A1(sw_rdat[26]), .Z(n213));
Q_AN02 U288 ( .A0(n508), .A1(wr_dat[27]), .Z(n214));
Q_MX02 U289 ( .S(n509), .A0(n214), .A1(sw_rdat[27]), .Z(n215));
Q_AN02 U290 ( .A0(n508), .A1(wr_dat[28]), .Z(n216));
Q_MX02 U291 ( .S(n509), .A0(n216), .A1(sw_rdat[28]), .Z(n217));
Q_AN02 U292 ( .A0(n508), .A1(wr_dat[29]), .Z(n218));
Q_MX02 U293 ( .S(n509), .A0(n218), .A1(sw_rdat[29]), .Z(n219));
Q_AN02 U294 ( .A0(n508), .A1(wr_dat[30]), .Z(n220));
Q_MX02 U295 ( .S(n509), .A0(n220), .A1(sw_rdat[30]), .Z(n221));
Q_AN02 U296 ( .A0(n508), .A1(wr_dat[31]), .Z(n222));
Q_MX02 U297 ( .S(n509), .A0(n222), .A1(sw_rdat[31]), .Z(n223));
Q_AN02 U298 ( .A0(n508), .A1(wr_dat[32]), .Z(n224));
Q_MX02 U299 ( .S(n509), .A0(n224), .A1(sw_rdat[32]), .Z(n225));
Q_AN02 U300 ( .A0(n508), .A1(wr_dat[33]), .Z(n226));
Q_MX02 U301 ( .S(n509), .A0(n226), .A1(sw_rdat[33]), .Z(n227));
Q_AN02 U302 ( .A0(n508), .A1(wr_dat[34]), .Z(n228));
Q_MX02 U303 ( .S(n509), .A0(n228), .A1(sw_rdat[34]), .Z(n229));
Q_AN02 U304 ( .A0(n508), .A1(wr_dat[35]), .Z(n230));
Q_MX02 U305 ( .S(n509), .A0(n230), .A1(sw_rdat[35]), .Z(n231));
Q_AN02 U306 ( .A0(n508), .A1(wr_dat[36]), .Z(n232));
Q_MX02 U307 ( .S(n509), .A0(n232), .A1(sw_rdat[36]), .Z(n233));
Q_AN02 U308 ( .A0(n508), .A1(wr_dat[37]), .Z(n234));
Q_MX02 U309 ( .S(n509), .A0(n234), .A1(sw_rdat[37]), .Z(n235));
Q_AN02 U310 ( .A0(n508), .A1(wr_dat[38]), .Z(n236));
Q_MX02 U311 ( .S(n509), .A0(n236), .A1(sw_rdat[38]), .Z(n237));
Q_AN02 U312 ( .A0(n508), .A1(wr_dat[39]), .Z(n238));
Q_MX02 U313 ( .S(n509), .A0(n238), .A1(sw_rdat[39]), .Z(n239));
Q_AN02 U314 ( .A0(n508), .A1(wr_dat[40]), .Z(n240));
Q_MX02 U315 ( .S(n509), .A0(n240), .A1(sw_rdat[40]), .Z(n241));
Q_AN02 U316 ( .A0(n508), .A1(wr_dat[41]), .Z(n242));
Q_MX02 U317 ( .S(n509), .A0(n242), .A1(sw_rdat[41]), .Z(n243));
Q_AN02 U318 ( .A0(n508), .A1(wr_dat[42]), .Z(n244));
Q_MX02 U319 ( .S(n509), .A0(n244), .A1(sw_rdat[42]), .Z(n245));
Q_AN02 U320 ( .A0(n508), .A1(wr_dat[43]), .Z(n246));
Q_MX02 U321 ( .S(n509), .A0(n246), .A1(sw_rdat[43]), .Z(n247));
Q_AN02 U322 ( .A0(n508), .A1(wr_dat[44]), .Z(n248));
Q_MX02 U323 ( .S(n509), .A0(n248), .A1(sw_rdat[44]), .Z(n249));
Q_AN02 U324 ( .A0(n508), .A1(wr_dat[45]), .Z(n250));
Q_MX02 U325 ( .S(n509), .A0(n250), .A1(sw_rdat[45]), .Z(n251));
Q_AN02 U326 ( .A0(n508), .A1(wr_dat[46]), .Z(n252));
Q_MX02 U327 ( .S(n509), .A0(n252), .A1(sw_rdat[46]), .Z(n253));
Q_AN02 U328 ( .A0(n508), .A1(wr_dat[47]), .Z(n254));
Q_MX02 U329 ( .S(n509), .A0(n254), .A1(sw_rdat[47]), .Z(n255));
Q_AN02 U330 ( .A0(n508), .A1(wr_dat[48]), .Z(n256));
Q_MX02 U331 ( .S(n509), .A0(n256), .A1(sw_rdat[48]), .Z(n257));
Q_AN02 U332 ( .A0(n508), .A1(wr_dat[49]), .Z(n258));
Q_MX02 U333 ( .S(n509), .A0(n258), .A1(sw_rdat[49]), .Z(n259));
Q_AN02 U334 ( .A0(n508), .A1(wr_dat[50]), .Z(n260));
Q_MX02 U335 ( .S(n509), .A0(n260), .A1(sw_rdat[50]), .Z(n261));
Q_AN02 U336 ( .A0(n508), .A1(wr_dat[51]), .Z(n262));
Q_MX02 U337 ( .S(n509), .A0(n262), .A1(sw_rdat[51]), .Z(n263));
Q_AN02 U338 ( .A0(n508), .A1(wr_dat[52]), .Z(n264));
Q_MX02 U339 ( .S(n509), .A0(n264), .A1(sw_rdat[52]), .Z(n265));
Q_AN02 U340 ( .A0(n508), .A1(wr_dat[53]), .Z(n266));
Q_MX02 U341 ( .S(n509), .A0(n266), .A1(sw_rdat[53]), .Z(n267));
Q_AN02 U342 ( .A0(n508), .A1(wr_dat[54]), .Z(n268));
Q_MX02 U343 ( .S(n509), .A0(n268), .A1(sw_rdat[54]), .Z(n269));
Q_AN02 U344 ( .A0(n508), .A1(wr_dat[55]), .Z(n270));
Q_MX02 U345 ( .S(n509), .A0(n270), .A1(sw_rdat[55]), .Z(n271));
Q_AN02 U346 ( .A0(n508), .A1(wr_dat[56]), .Z(n272));
Q_MX02 U347 ( .S(n509), .A0(n272), .A1(sw_rdat[56]), .Z(n273));
Q_AN02 U348 ( .A0(n508), .A1(wr_dat[57]), .Z(n274));
Q_MX02 U349 ( .S(n509), .A0(n274), .A1(sw_rdat[57]), .Z(n275));
Q_AN02 U350 ( .A0(n508), .A1(wr_dat[58]), .Z(n276));
Q_MX02 U351 ( .S(n509), .A0(n276), .A1(sw_rdat[58]), .Z(n277));
Q_AN02 U352 ( .A0(n508), .A1(wr_dat[59]), .Z(n278));
Q_MX02 U353 ( .S(n509), .A0(n278), .A1(sw_rdat[59]), .Z(n279));
Q_AN02 U354 ( .A0(n508), .A1(wr_dat[60]), .Z(n280));
Q_MX02 U355 ( .S(n509), .A0(n280), .A1(sw_rdat[60]), .Z(n281));
Q_AN02 U356 ( .A0(n508), .A1(wr_dat[61]), .Z(n282));
Q_MX02 U357 ( .S(n509), .A0(n282), .A1(sw_rdat[61]), .Z(n283));
Q_AN02 U358 ( .A0(n508), .A1(wr_dat[62]), .Z(n284));
Q_MX02 U359 ( .S(n509), .A0(n284), .A1(sw_rdat[62]), .Z(n285));
Q_AN02 U360 ( .A0(n508), .A1(wr_dat[63]), .Z(n286));
Q_MX02 U361 ( .S(n509), .A0(n286), .A1(sw_rdat[63]), .Z(n287));
Q_AN02 U362 ( .A0(n508), .A1(wr_dat[64]), .Z(n288));
Q_MX02 U363 ( .S(n509), .A0(n288), .A1(sw_rdat[64]), .Z(n289));
Q_AN02 U364 ( .A0(n508), .A1(wr_dat[65]), .Z(n290));
Q_MX02 U365 ( .S(n509), .A0(n290), .A1(sw_rdat[65]), .Z(n291));
Q_AN02 U366 ( .A0(n508), .A1(wr_dat[66]), .Z(n292));
Q_MX02 U367 ( .S(n509), .A0(n292), .A1(sw_rdat[66]), .Z(n293));
Q_AN02 U368 ( .A0(n508), .A1(wr_dat[67]), .Z(n294));
Q_MX02 U369 ( .S(n509), .A0(n294), .A1(sw_rdat[67]), .Z(n295));
Q_AN02 U370 ( .A0(n508), .A1(wr_dat[68]), .Z(n296));
Q_MX02 U371 ( .S(n509), .A0(n296), .A1(sw_rdat[68]), .Z(n297));
Q_AN02 U372 ( .A0(n508), .A1(wr_dat[69]), .Z(n298));
Q_MX02 U373 ( .S(n509), .A0(n298), .A1(sw_rdat[69]), .Z(n299));
Q_AN02 U374 ( .A0(n508), .A1(wr_dat[70]), .Z(n300));
Q_MX02 U375 ( .S(n509), .A0(n300), .A1(sw_rdat[70]), .Z(n301));
Q_AN02 U376 ( .A0(n508), .A1(wr_dat[71]), .Z(n302));
Q_MX02 U377 ( .S(n509), .A0(n302), .A1(sw_rdat[71]), .Z(n303));
Q_AN02 U378 ( .A0(n508), .A1(wr_dat[72]), .Z(n304));
Q_MX02 U379 ( .S(n509), .A0(n304), .A1(sw_rdat[72]), .Z(n305));
Q_AN02 U380 ( .A0(n508), .A1(wr_dat[73]), .Z(n306));
Q_MX02 U381 ( .S(n509), .A0(n306), .A1(sw_rdat[73]), .Z(n307));
Q_AN02 U382 ( .A0(n508), .A1(wr_dat[74]), .Z(n308));
Q_MX02 U383 ( .S(n509), .A0(n308), .A1(sw_rdat[74]), .Z(n309));
Q_AN02 U384 ( .A0(n508), .A1(wr_dat[75]), .Z(n310));
Q_MX02 U385 ( .S(n509), .A0(n310), .A1(sw_rdat[75]), .Z(n311));
Q_AN02 U386 ( .A0(n508), .A1(wr_dat[76]), .Z(n312));
Q_MX02 U387 ( .S(n509), .A0(n312), .A1(sw_rdat[76]), .Z(n313));
Q_AN02 U388 ( .A0(n508), .A1(wr_dat[77]), .Z(n314));
Q_MX02 U389 ( .S(n509), .A0(n314), .A1(sw_rdat[77]), .Z(n315));
Q_AN02 U390 ( .A0(n508), .A1(wr_dat[78]), .Z(n316));
Q_MX02 U391 ( .S(n509), .A0(n316), .A1(sw_rdat[78]), .Z(n317));
Q_AN02 U392 ( .A0(n508), .A1(wr_dat[79]), .Z(n318));
Q_MX02 U393 ( .S(n509), .A0(n318), .A1(sw_rdat[79]), .Z(n319));
Q_AN02 U394 ( .A0(n508), .A1(wr_dat[80]), .Z(n320));
Q_MX02 U395 ( .S(n509), .A0(n320), .A1(sw_rdat[80]), .Z(n321));
Q_AN02 U396 ( .A0(n508), .A1(wr_dat[81]), .Z(n322));
Q_MX02 U397 ( .S(n509), .A0(n322), .A1(sw_rdat[81]), .Z(n323));
Q_AN02 U398 ( .A0(n508), .A1(wr_dat[82]), .Z(n324));
Q_MX02 U399 ( .S(n509), .A0(n324), .A1(sw_rdat[82]), .Z(n325));
Q_AN02 U400 ( .A0(n508), .A1(wr_dat[83]), .Z(n326));
Q_MX02 U401 ( .S(n509), .A0(n326), .A1(sw_rdat[83]), .Z(n327));
Q_AN02 U402 ( .A0(n508), .A1(wr_dat[84]), .Z(n328));
Q_MX02 U403 ( .S(n509), .A0(n328), .A1(sw_rdat[84]), .Z(n329));
Q_AN02 U404 ( .A0(n508), .A1(wr_dat[85]), .Z(n330));
Q_MX02 U405 ( .S(n509), .A0(n330), .A1(sw_rdat[85]), .Z(n331));
Q_AN02 U406 ( .A0(n508), .A1(wr_dat[86]), .Z(n332));
Q_MX02 U407 ( .S(n509), .A0(n332), .A1(sw_rdat[86]), .Z(n333));
Q_AN02 U408 ( .A0(n508), .A1(wr_dat[87]), .Z(n334));
Q_MX02 U409 ( .S(n509), .A0(n334), .A1(sw_rdat[87]), .Z(n335));
Q_AN02 U410 ( .A0(n508), .A1(wr_dat[88]), .Z(n336));
Q_MX02 U411 ( .S(n509), .A0(n336), .A1(sw_rdat[88]), .Z(n337));
Q_AN02 U412 ( .A0(n508), .A1(wr_dat[89]), .Z(n338));
Q_MX02 U413 ( .S(n509), .A0(n338), .A1(sw_rdat[89]), .Z(n339));
Q_AN02 U414 ( .A0(n508), .A1(wr_dat[90]), .Z(n340));
Q_MX02 U415 ( .S(n509), .A0(n340), .A1(sw_rdat[90]), .Z(n341));
Q_AN02 U416 ( .A0(n508), .A1(wr_dat[91]), .Z(n342));
Q_MX02 U417 ( .S(n509), .A0(n342), .A1(sw_rdat[91]), .Z(n343));
Q_AN02 U418 ( .A0(n508), .A1(wr_dat[92]), .Z(n344));
Q_MX02 U419 ( .S(n509), .A0(n344), .A1(sw_rdat[92]), .Z(n345));
Q_AN02 U420 ( .A0(n508), .A1(wr_dat[93]), .Z(n346));
Q_MX02 U421 ( .S(n509), .A0(n346), .A1(sw_rdat[93]), .Z(n347));
Q_AN02 U422 ( .A0(n508), .A1(wr_dat[94]), .Z(n348));
Q_MX02 U423 ( .S(n509), .A0(n348), .A1(sw_rdat[94]), .Z(n349));
Q_AN02 U424 ( .A0(n508), .A1(wr_dat[95]), .Z(n350));
Q_MX02 U425 ( .S(n509), .A0(n350), .A1(sw_rdat[95]), .Z(n351));
Q_FDP1 \state_r_REG[3] ( .CK(clk), .R(rst_n), .D(n523), .Q(state_r[3]), .QN(n409));
Q_FDP1 \state_r_REG[2] ( .CK(clk), .R(rst_n), .D(n522), .Q(state_r[2]), .QN(n410));
Q_FDP1 \state_r_REG[1] ( .CK(clk), .R(rst_n), .D(n521), .Q(state_r[1]), .QN(n412));
Q_FDP1 \state_r_REG[0] ( .CK(clk), .R(rst_n), .D(n520), .Q(state_r[0]), .QN(n381));
Q_FDP1 \timer_r_REG[5] ( .CK(clk), .R(rst_n), .D(n149), .Q(timer_r[5]), .QN( ));
Q_FDP1 \timer_r_REG[4] ( .CK(clk), .R(rst_n), .D(n148), .Q(timer_r[4]), .QN( ));
Q_FDP1 \timer_r_REG[3] ( .CK(clk), .R(rst_n), .D(n147), .Q(timer_r[3]), .QN( ));
Q_FDP1 \timer_r_REG[2] ( .CK(clk), .R(rst_n), .D(n146), .Q(timer_r[2]), .QN( ));
Q_FDP1 \timer_r_REG[1] ( .CK(clk), .R(rst_n), .D(n145), .Q(timer_r[1]), .QN( ));
Q_FDP1 \timer_r_REG[0] ( .CK(clk), .R(rst_n), .D(n144), .Q(timer_r[0]), .QN(n113));
Q_ND02 U436 ( .A0(n353), .A1(n354), .Z(n352));
Q_ND02 U437 ( .A0(n355), .A1(n467), .Z(n354));
Q_OR02 U438 ( .A0(n356), .A1(n511), .Z(n355));
Q_INV U439 ( .A(n510), .Z(n356));
Q_ND02 U440 ( .A0(n353), .A1(n358), .Z(n357));
Q_ND02 U441 ( .A0(n510), .A1(n467), .Z(n358));
Q_OR03 U442 ( .A0(n510), .A1(n511), .A2(n467), .Z(n353));
Q_MX02 U443 ( .S(n467), .A0(n510), .A1(n511), .Z(n359));
Q_FDP2 \stat_code_REG[2] ( .CK(clk), .S(rst_n), .D(n360), .Q(stat_code[2]), .QN( ));
Q_MX02 U445 ( .S(n482), .A0(stat_code[2]), .A1(n359), .Z(n360));
Q_FDP2 \stat_code_REG[1] ( .CK(clk), .S(rst_n), .D(n361), .Q(stat_code[1]), .QN( ));
Q_MX02 U447 ( .S(n482), .A0(stat_code[1]), .A1(n357), .Z(n361));
Q_FDP2 \stat_code_REG[0] ( .CK(clk), .S(rst_n), .D(n362), .Q(stat_code[0]), .QN( ));
Q_MX02 U449 ( .S(n482), .A0(stat_code[0]), .A1(n352), .Z(n362));
Q_FDP2 init_r_REG  ( .CK(clk), .S(rst_n), .D(n363), .Q(init_r), .QN(enable));
Q_MX02 U451 ( .S(n513), .A0(init_r), .A1(n507), .Z(n363));
Q_FDP1 sw_cs_r_REG  ( .CK(clk), .R(rst_n), .D(n505), .Q(sw_cs_r), .QN( ));
Q_FDP1 sw_ce_r_REG  ( .CK(clk), .R(rst_n), .D(n504), .Q(sw_ce_r), .QN( ));
Q_FDP1 rst_r_REG  ( .CK(clk), .R(rst_n), .D(n503), .Q(rst_r), .QN(n524));
Q_FDP1 rst_or_ini_r_REG  ( .CK(clk), .R(rst_n), .D(n502), .Q(rst_or_ini_r), .QN( ));
Q_FDP1 sw_we_r_REG  ( .CK(clk), .R(rst_n), .D(n499), .Q(sw_we_r), .QN( ));
Q_OA21 U457 ( .A0(n365), .A1(n366), .B0(n364), .Z(n494));
Q_OR03 U458 ( .A0(n368), .A1(n369), .A2(n367), .Z(n366));
Q_AN03 U459 ( .A0(state_r[0]), .A1(n372), .A2(n370), .Z(n371));
Q_AN02 U460 ( .A0(n67), .A1(cmnd_rd_stb), .Z(n372));
Q_AN02 U461 ( .A0(n375), .A1(n64), .Z(n376));
Q_AN03 U462 ( .A0(n377), .A1(n376), .A2(n373), .Z(n374));
Q_AN02 U463 ( .A0(n378), .A1(state_r[0]), .Z(n377));
Q_OR03 U464 ( .A0(n374), .A1(n379), .A2(n371), .Z(n369));
Q_AN02 U465 ( .A0(n370), .A1(n380), .Z(n379));
Q_NR02 U466 ( .A0(state_r[0]), .A1(cmnd_ena_stb), .Z(n380));
Q_OA21 U467 ( .A0(n383), .A1(n384), .B0(n382), .Z(n368));
Q_AN02 U468 ( .A0(n385), .A1(n386), .Z(n384));
Q_NR02 U469 ( .A0(state_r[0]), .A1(igrant), .Z(n386));
Q_OA21 U470 ( .A0(n389), .A1(n390), .B0(n388), .Z(n383));
Q_AN02 U471 ( .A0(n391), .A1(n387), .Z(n390));
Q_NR02 U472 ( .A0(n392), .A1(n519), .Z(n389));
Q_INV U473 ( .A(n393), .Z(n375));
Q_AN03 U474 ( .A0(cmnd_rst_stb), .A1(n370), .A2(n395), .Z(n396));
Q_OR03 U475 ( .A0(n397), .A1(n396), .A2(n394), .Z(n365));
Q_AN03 U476 ( .A0(n381), .A1(n399), .A2(n398), .Z(n397));
Q_INV U477 ( .A(n400), .Z(n495));
Q_OA21 U478 ( .A0(n401), .A1(n367), .B0(n364), .Z(n400));
Q_AO21 U479 ( .A0(n370), .A1(n404), .B0(n403), .Z(n401));
Q_AN02 U480 ( .A0(state_r[0]), .A1(cmnd_wr_stb), .Z(n404));
Q_AN03 U481 ( .A0(n408), .A1(n381), .A2(n406), .Z(n407));
Q_NR02 U482 ( .A0(state_r[3]), .A1(state_r[2]), .Z(n408));
Q_MX02 U483 ( .S(state_r[1]), .A0(cmnd_ena_stb), .A1(n411), .Z(n406));
Q_OR03 U484 ( .A0(n413), .A1(n407), .A2(n405), .Z(n367));
Q_AN02 U485 ( .A0(n414), .A1(n382), .Z(n405));
Q_AN02 U486 ( .A0(n378), .A1(n64), .Z(n382));
Q_AN02 U487 ( .A0(n415), .A1(n416), .Z(n413));
Q_NR02 U488 ( .A0(cmnd_dis_stb), .A1(unsupported_op), .Z(n416));
Q_MX02 U489 ( .S(state_r[3]), .A0(n418), .A1(n417), .Z(n414));
Q_AN02 U490 ( .A0(n453), .A1(n411), .Z(n419));
Q_AN02 U491 ( .A0(ack_error), .A1(enable), .Z(n411));
Q_AO21 U492 ( .A0(n420), .A1(n381), .B0(n419), .Z(n417));
Q_AN02 U493 ( .A0(state_r[2]), .A1(igrant), .Z(n422));
Q_AO21 U494 ( .A0(n423), .A1(n424), .B0(n421), .Z(n418));
Q_OA21 U495 ( .A0(state_r[0]), .A1(n425), .B0(n422), .Z(n421));
Q_AN02 U496 ( .A0(n412), .A1(n519), .Z(n425));
Q_OR02 U497 ( .A0(state_r[2]), .A1(n393), .Z(n423));
Q_AN02 U498 ( .A0(igrant), .A1(n518), .Z(n393));
Q_OA21 U499 ( .A0(n426), .A1(n427), .B0(n402), .Z(n403));
Q_AN03 U500 ( .A0(n428), .A1(n409), .A2(n395), .Z(n427));
Q_AN02 U501 ( .A0(n429), .A1(n430), .Z(n426));
Q_AN03 U502 ( .A0(n432), .A1(n433), .A2(n431), .Z(n496));
Q_AO21 U503 ( .A0(n428), .A1(n435), .B0(n434), .Z(n431));
Q_INV U504 ( .A(n434), .Z(n435));
Q_INV U505 ( .A(n436), .Z(n497));
Q_OA21 U506 ( .A0(n437), .A1(n394), .B0(n364), .Z(n436));
Q_AN03 U507 ( .A0(n434), .A1(n433), .A2(n370), .Z(n438));
Q_AN02 U508 ( .A0(state_r[0]), .A1(n67), .Z(n433));
Q_AO21 U509 ( .A0(n68), .A1(cmnd_cmp_stb), .B0(cmnd_rd_stb), .Z(n434));
Q_AN03 U510 ( .A0(n428), .A1(n370), .A2(n395), .Z(n439));
Q_AN02 U511 ( .A0(n440), .A1(n65), .Z(n395));
Q_AO21 U512 ( .A0(n66), .A1(n517), .B0(cmnd_rst_stb), .Z(n428));
Q_AN03 U513 ( .A0(n429), .A1(n64), .A2(n398), .Z(n442));
Q_AN02 U514 ( .A0(n378), .A1(n385), .Z(n398));
Q_AN02 U515 ( .A0(state_r[3]), .A1(n402), .Z(n385));
Q_OR03 U516 ( .A0(n442), .A1(n441), .A2(n438), .Z(n437));
Q_AO21 U517 ( .A0(n443), .A1(n444), .B0(n439), .Z(n441));
Q_AN02 U518 ( .A0(igrant), .A1(n64), .Z(n399));
Q_AN02 U519 ( .A0(n445), .A1(n399), .Z(n443));
Q_NR02 U520 ( .A0(timeout), .A1(state_r[0]), .Z(n445));
Q_AN02 U521 ( .A0(ack_error), .A1(init_r), .Z(n447));
Q_AO21 U522 ( .A0(n415), .A1(cmnd_dis_stb), .B0(n446), .Z(n394));
Q_AN02 U523 ( .A0(n440), .A1(n449), .Z(n448));
Q_NR02 U524 ( .A0(cmnd_cmp_stb), .A1(n517), .Z(n449));
Q_AN02 U525 ( .A0(state_r[0]), .A1(n450), .Z(n440));
Q_NR02 U526 ( .A0(cmnd_wr_stb), .A1(cmnd_rd_stb), .Z(n450));
Q_AN03 U527 ( .A0(n66), .A1(n370), .A2(n448), .Z(n415));
Q_OA21 U528 ( .A0(n451), .A1(n452), .B0(n447), .Z(n446));
Q_AN02 U529 ( .A0(n453), .A1(n430), .Z(n451));
Q_AN03 U530 ( .A0(n378), .A1(state_r[3]), .A2(n64), .Z(n430));
Q_INV U531 ( .A(n391), .Z(n424));
Q_AO21 U532 ( .A0(n381), .A1(igrant), .B0(state_r[0]), .Z(n429));
Q_AN02 U533 ( .A0(n387), .A1(n505), .Z(n498));
Q_INV U534 ( .A(igrant), .Z(n387));
Q_OA21 U535 ( .A0(n455), .A1(n456), .B0(n454), .Z(n499));
Q_AN02 U536 ( .A0(n522), .A1(n457), .Z(n456));
Q_AN02 U537 ( .A0(cmnd_sis_stb), .A1(n458), .Z(n500));
Q_INV U538 ( .A(n501), .Z(n458));
Q_ND02 U539 ( .A0(n391), .A1(n410), .Z(n453));
Q_OR02 U540 ( .A0(state_r[0]), .A1(state_r[1]), .Z(n392));
Q_ND02 U541 ( .A0(state_r[1]), .A1(state_r[0]), .Z(n391));
Q_OA21 U542 ( .A0(n455), .A1(n459), .B0(n454), .Z(n502));
Q_AN02 U543 ( .A0(n522), .A1(n460), .Z(n459));
Q_AN02 U544 ( .A0(n461), .A1(n462), .Z(n455));
Q_AN02 U545 ( .A0(n463), .A1(n462), .Z(n503));
Q_OR03 U546 ( .A0(n464), .A1(n504), .A2(n503), .Z(n505));
Q_AN03 U547 ( .A0(n523), .A1(n461), .A2(n460), .Z(n504));
Q_AN03 U548 ( .A0(n454), .A1(n522), .A2(n465), .Z(n464));
Q_INV U549 ( .A(n462), .Z(n465));
Q_INV U550 ( .A(n466), .Z(n506));
Q_AN02 U551 ( .A0(n444), .A1(state_r[0]), .Z(n509));
Q_AN03 U552 ( .A0(state_r[2]), .A1(state_r[1]), .A2(n409), .Z(n444));
Q_AN02 U553 ( .A0(n469), .A1(n470), .Z(n471));
Q_INV U554 ( .A(n472), .Z(n469));
Q_OR03 U555 ( .A0(n473), .A1(n471), .A2(n468), .Z(n467));
Q_AN03 U556 ( .A0(n475), .A1(n63), .A2(n474), .Z(n468));
Q_OR02 U557 ( .A0(n462), .A1(n476), .Z(n473));
Q_AN02 U558 ( .A0(n521), .A1(n520), .Z(n462));
Q_INV U559 ( .A(n463), .Z(n476));
Q_AN02 U560 ( .A0(n463), .A1(n477), .Z(n470));
Q_OA21 U561 ( .A0(n478), .A1(n457), .B0(n470), .Z(n510));
Q_AN02 U562 ( .A0(n63), .A1(n521), .Z(n472));
Q_OA21 U563 ( .A0(n475), .A1(badaddr), .B0(n472), .Z(n478));
Q_AN02 U564 ( .A0(timeout), .A1(n364), .Z(n475));
Q_OA21 U565 ( .A0(n479), .A1(n480), .B0(n463), .Z(n511));
Q_AO21 U566 ( .A0(n457), .A1(n520), .B0(n460), .Z(n480));
Q_AN02 U567 ( .A0(unsupported_op), .A1(n481), .Z(n479));
Q_ND02 U568 ( .A0(n452), .A1(n474), .Z(n482));
Q_AN02 U569 ( .A0(n463), .A1(n481), .Z(n474));
Q_AN02 U570 ( .A0(n521), .A1(n477), .Z(n481));
Q_AN02 U571 ( .A0(n373), .A1(n381), .Z(n452));
Q_AN02 U572 ( .A0(n409), .A1(n420), .Z(n373));
Q_OA21 U573 ( .A0(n508), .A1(n483), .B0(n364), .Z(n512));
Q_AN02 U574 ( .A0(n484), .A1(state_r[1]), .Z(n483));
Q_INV U575 ( .A(n507), .Z(n508));
Q_AN02 U576 ( .A0(n409), .A1(n402), .Z(n370));
Q_MX02 U577 ( .S(state_r[0]), .A0(n485), .A1(n388), .Z(n484));
Q_AN02 U578 ( .A0(state_r[3]), .A1(n410), .Z(n485));
Q_AN02 U579 ( .A0(n409), .A1(state_r[2]), .Z(n388));
Q_AN03 U580 ( .A0(n463), .A1(n460), .A2(n507), .Z(n486));
Q_NR02 U581 ( .A0(n521), .A1(n520), .Z(n460));
Q_INV U582 ( .A(n520), .Z(n477));
Q_INV U583 ( .A(n521), .Z(n457));
Q_NR02 U584 ( .A0(n523), .A1(n522), .Z(n463));
Q_INV U585 ( .A(n522), .Z(n461));
Q_INV U586 ( .A(n523), .Z(n454));
Q_AO21 U587 ( .A0(n432), .A1(n487), .B0(n486), .Z(n513));
Q_AN02 U588 ( .A0(n381), .A1(cmnd_ena_stb), .Z(n487));
Q_OR02 U589 ( .A0(state_r[3]), .A1(state_r[1]), .Z(n488));
Q_OR03 U590 ( .A0(state_r[2]), .A1(state_r[0]), .A2(n488), .Z(n507));
Q_AN03 U591 ( .A0(n490), .A1(n412), .A2(n489), .Z(n514));
Q_AO21 U592 ( .A0(state_r[2]), .A1(n381), .B0(n466), .Z(n489));
Q_AN02 U593 ( .A0(n410), .A1(state_r[0]), .Z(n466));
Q_ND02 U594 ( .A0(n432), .A1(state_r[0]), .Z(n515));
Q_AN02 U595 ( .A0(n490), .A1(n402), .Z(n432));
Q_NR02 U596 ( .A0(state_r[2]), .A1(state_r[1]), .Z(n402));
Q_AN02 U597 ( .A0(n491), .A1(n490), .Z(n501));
Q_NR02 U598 ( .A0(badaddr), .A1(state_r[3]), .Z(n490));
Q_INV U599 ( .A(badaddr), .Z(n364));
Q_OR03 U600 ( .A0(cmnd_rst_stb), .A1(cmnd_sis_stb), .A2(n501), .Z(n516));
Q_MX02 U601 ( .S(state_r[0]), .A0(n492), .A1(n420), .Z(n491));
Q_AN02 U602 ( .A0(state_r[2]), .A1(n412), .Z(n492));
Q_AN02 U603 ( .A0(n410), .A1(state_r[1]), .Z(n420));
Q_OR02 U604 ( .A0(cmnd_tmo_stb), .A1(timeout), .Z(n493));
Q_INV U605 ( .A(timeout), .Z(n378));
Q_AN02 U606 ( .A0(n524), .A1(wr_dat[0]), .Z(sw_wdat[0]));
Q_AN02 U607 ( .A0(n524), .A1(wr_dat[1]), .Z(sw_wdat[1]));
Q_AN02 U608 ( .A0(n524), .A1(wr_dat[2]), .Z(sw_wdat[2]));
Q_AN02 U609 ( .A0(n524), .A1(wr_dat[3]), .Z(sw_wdat[3]));
Q_AN02 U610 ( .A0(n524), .A1(wr_dat[4]), .Z(sw_wdat[4]));
Q_AN02 U611 ( .A0(n524), .A1(wr_dat[5]), .Z(sw_wdat[5]));
Q_AN02 U612 ( .A0(n524), .A1(wr_dat[6]), .Z(sw_wdat[6]));
Q_AN02 U613 ( .A0(n524), .A1(wr_dat[7]), .Z(sw_wdat[7]));
Q_AN02 U614 ( .A0(n524), .A1(wr_dat[8]), .Z(sw_wdat[8]));
Q_AN02 U615 ( .A0(n524), .A1(wr_dat[9]), .Z(sw_wdat[9]));
Q_AN02 U616 ( .A0(n524), .A1(wr_dat[10]), .Z(sw_wdat[10]));
Q_AN02 U617 ( .A0(n524), .A1(wr_dat[11]), .Z(sw_wdat[11]));
Q_AN02 U618 ( .A0(n524), .A1(wr_dat[12]), .Z(sw_wdat[12]));
Q_AN02 U619 ( .A0(n524), .A1(wr_dat[13]), .Z(sw_wdat[13]));
Q_AN02 U620 ( .A0(n524), .A1(wr_dat[14]), .Z(sw_wdat[14]));
Q_AN02 U621 ( .A0(n524), .A1(wr_dat[15]), .Z(sw_wdat[15]));
Q_AN02 U622 ( .A0(n524), .A1(wr_dat[16]), .Z(sw_wdat[16]));
Q_AN02 U623 ( .A0(n524), .A1(wr_dat[17]), .Z(sw_wdat[17]));
Q_AN02 U624 ( .A0(n524), .A1(wr_dat[18]), .Z(sw_wdat[18]));
Q_AN02 U625 ( .A0(n524), .A1(wr_dat[19]), .Z(sw_wdat[19]));
Q_AN02 U626 ( .A0(n524), .A1(wr_dat[20]), .Z(sw_wdat[20]));
Q_AN02 U627 ( .A0(n524), .A1(wr_dat[21]), .Z(sw_wdat[21]));
Q_AN02 U628 ( .A0(n524), .A1(wr_dat[22]), .Z(sw_wdat[22]));
Q_AN02 U629 ( .A0(n524), .A1(wr_dat[23]), .Z(sw_wdat[23]));
Q_AN02 U630 ( .A0(n524), .A1(wr_dat[24]), .Z(sw_wdat[24]));
Q_AN02 U631 ( .A0(n524), .A1(wr_dat[25]), .Z(sw_wdat[25]));
Q_AN02 U632 ( .A0(n524), .A1(wr_dat[26]), .Z(sw_wdat[26]));
Q_AN02 U633 ( .A0(n524), .A1(wr_dat[27]), .Z(sw_wdat[27]));
Q_AN02 U634 ( .A0(n524), .A1(wr_dat[28]), .Z(sw_wdat[28]));
Q_AN02 U635 ( .A0(n524), .A1(wr_dat[29]), .Z(sw_wdat[29]));
Q_AN02 U636 ( .A0(n524), .A1(wr_dat[30]), .Z(sw_wdat[30]));
Q_AN02 U637 ( .A0(n524), .A1(wr_dat[31]), .Z(sw_wdat[31]));
Q_AN02 U638 ( .A0(n524), .A1(wr_dat[32]), .Z(sw_wdat[32]));
Q_AN02 U639 ( .A0(n524), .A1(wr_dat[33]), .Z(sw_wdat[33]));
Q_AN02 U640 ( .A0(n524), .A1(wr_dat[34]), .Z(sw_wdat[34]));
Q_AN02 U641 ( .A0(n524), .A1(wr_dat[35]), .Z(sw_wdat[35]));
Q_AN02 U642 ( .A0(n524), .A1(wr_dat[36]), .Z(sw_wdat[36]));
Q_AN02 U643 ( .A0(n524), .A1(wr_dat[37]), .Z(sw_wdat[37]));
Q_AN02 U644 ( .A0(n524), .A1(wr_dat[38]), .Z(sw_wdat[38]));
Q_AN02 U645 ( .A0(n524), .A1(wr_dat[39]), .Z(sw_wdat[39]));
Q_AN02 U646 ( .A0(n524), .A1(wr_dat[40]), .Z(sw_wdat[40]));
Q_AN02 U647 ( .A0(n524), .A1(wr_dat[41]), .Z(sw_wdat[41]));
Q_AN02 U648 ( .A0(n524), .A1(wr_dat[42]), .Z(sw_wdat[42]));
Q_AN02 U649 ( .A0(n524), .A1(wr_dat[43]), .Z(sw_wdat[43]));
Q_AN02 U650 ( .A0(n524), .A1(wr_dat[44]), .Z(sw_wdat[44]));
Q_AN02 U651 ( .A0(n524), .A1(wr_dat[45]), .Z(sw_wdat[45]));
Q_AN02 U652 ( .A0(n524), .A1(wr_dat[46]), .Z(sw_wdat[46]));
Q_AN02 U653 ( .A0(n524), .A1(wr_dat[47]), .Z(sw_wdat[47]));
Q_AN02 U654 ( .A0(n524), .A1(wr_dat[48]), .Z(sw_wdat[48]));
Q_AN02 U655 ( .A0(n524), .A1(wr_dat[49]), .Z(sw_wdat[49]));
Q_AN02 U656 ( .A0(n524), .A1(wr_dat[50]), .Z(sw_wdat[50]));
Q_AN02 U657 ( .A0(n524), .A1(wr_dat[51]), .Z(sw_wdat[51]));
Q_AN02 U658 ( .A0(n524), .A1(wr_dat[52]), .Z(sw_wdat[52]));
Q_AN02 U659 ( .A0(n524), .A1(wr_dat[53]), .Z(sw_wdat[53]));
Q_AN02 U660 ( .A0(n524), .A1(wr_dat[54]), .Z(sw_wdat[54]));
Q_AN02 U661 ( .A0(n524), .A1(wr_dat[55]), .Z(sw_wdat[55]));
Q_AN02 U662 ( .A0(n524), .A1(wr_dat[56]), .Z(sw_wdat[56]));
Q_AN02 U663 ( .A0(n524), .A1(wr_dat[57]), .Z(sw_wdat[57]));
Q_AN02 U664 ( .A0(n524), .A1(wr_dat[58]), .Z(sw_wdat[58]));
Q_AN02 U665 ( .A0(n524), .A1(wr_dat[59]), .Z(sw_wdat[59]));
Q_AN02 U666 ( .A0(n524), .A1(wr_dat[60]), .Z(sw_wdat[60]));
Q_AN02 U667 ( .A0(n524), .A1(wr_dat[61]), .Z(sw_wdat[61]));
Q_AN02 U668 ( .A0(n524), .A1(wr_dat[62]), .Z(sw_wdat[62]));
Q_AN02 U669 ( .A0(n524), .A1(wr_dat[63]), .Z(sw_wdat[63]));
Q_AN02 U670 ( .A0(n524), .A1(wr_dat[64]), .Z(sw_wdat[64]));
Q_AN02 U671 ( .A0(n524), .A1(wr_dat[65]), .Z(sw_wdat[65]));
Q_AN02 U672 ( .A0(n524), .A1(wr_dat[66]), .Z(sw_wdat[66]));
Q_AN02 U673 ( .A0(n524), .A1(wr_dat[67]), .Z(sw_wdat[67]));
Q_AN02 U674 ( .A0(n524), .A1(wr_dat[68]), .Z(sw_wdat[68]));
Q_AN02 U675 ( .A0(n524), .A1(wr_dat[69]), .Z(sw_wdat[69]));
Q_AN02 U676 ( .A0(n524), .A1(wr_dat[70]), .Z(sw_wdat[70]));
Q_AN02 U677 ( .A0(n524), .A1(wr_dat[71]), .Z(sw_wdat[71]));
Q_AN02 U678 ( .A0(n524), .A1(wr_dat[72]), .Z(sw_wdat[72]));
Q_AN02 U679 ( .A0(n524), .A1(wr_dat[73]), .Z(sw_wdat[73]));
Q_AN02 U680 ( .A0(n524), .A1(wr_dat[74]), .Z(sw_wdat[74]));
Q_AN02 U681 ( .A0(n524), .A1(wr_dat[75]), .Z(sw_wdat[75]));
Q_AN02 U682 ( .A0(n524), .A1(wr_dat[76]), .Z(sw_wdat[76]));
Q_AN02 U683 ( .A0(n524), .A1(wr_dat[77]), .Z(sw_wdat[77]));
Q_AN02 U684 ( .A0(n524), .A1(wr_dat[78]), .Z(sw_wdat[78]));
Q_AN02 U685 ( .A0(n524), .A1(wr_dat[79]), .Z(sw_wdat[79]));
Q_AN02 U686 ( .A0(n524), .A1(wr_dat[80]), .Z(sw_wdat[80]));
Q_AN02 U687 ( .A0(n524), .A1(wr_dat[81]), .Z(sw_wdat[81]));
Q_AN02 U688 ( .A0(n524), .A1(wr_dat[82]), .Z(sw_wdat[82]));
Q_AN02 U689 ( .A0(n524), .A1(wr_dat[83]), .Z(sw_wdat[83]));
Q_AN02 U690 ( .A0(n524), .A1(wr_dat[84]), .Z(sw_wdat[84]));
Q_AN02 U691 ( .A0(n524), .A1(wr_dat[85]), .Z(sw_wdat[85]));
Q_AN02 U692 ( .A0(n524), .A1(wr_dat[86]), .Z(sw_wdat[86]));
Q_AN02 U693 ( .A0(n524), .A1(wr_dat[87]), .Z(sw_wdat[87]));
Q_AN02 U694 ( .A0(n524), .A1(wr_dat[88]), .Z(sw_wdat[88]));
Q_AN02 U695 ( .A0(n524), .A1(wr_dat[89]), .Z(sw_wdat[89]));
Q_AN02 U696 ( .A0(n524), .A1(wr_dat[90]), .Z(sw_wdat[90]));
Q_AN02 U697 ( .A0(n524), .A1(wr_dat[91]), .Z(sw_wdat[91]));
Q_AN02 U698 ( .A0(n524), .A1(wr_dat[92]), .Z(sw_wdat[92]));
Q_AN02 U699 ( .A0(n524), .A1(wr_dat[93]), .Z(sw_wdat[93]));
Q_AN02 U700 ( .A0(n524), .A1(wr_dat[94]), .Z(sw_wdat[94]));
Q_AN02 U701 ( .A0(n524), .A1(wr_dat[95]), .Z(sw_wdat[95]));
Q_FDP4EP sim_tmo_r_REG  ( .CK(clk), .CE(n493), .R(n525), .D(cmnd_tmo_stb), .Q(sim_tmo_r));
Q_INV U703 ( .A(rst_n), .Z(n525));
Q_INV U704 ( .A(sim_tmo_r), .Z(n36));
Q_FDP4EP \rst_addr_r_REG[0] ( .CK(clk), .CE(n516), .R(n525), .D(n151), .Q(rst_addr_r[0]));
Q_FDP4EP \rst_addr_r_REG[1] ( .CK(clk), .CE(n516), .R(n525), .D(n153), .Q(rst_addr_r[1]));
Q_FDP4EP \rst_addr_r_REG[2] ( .CK(clk), .CE(n516), .R(n525), .D(n155), .Q(rst_addr_r[2]));
Q_FDP4EP \rst_addr_r_REG[3] ( .CK(clk), .CE(n516), .R(n525), .D(n157), .Q(rst_addr_r[3]));
Q_FDP4EP \rst_addr_r_REG[4] ( .CK(clk), .CE(n516), .R(n525), .D(n159), .Q(rst_addr_r[4]));
Q_FDP4EP \rst_addr_r_REG[5] ( .CK(clk), .CE(n516), .R(n525), .D(n161), .Q(rst_addr_r[5]));
Q_FDP4EP \rst_addr_r_REG[6] ( .CK(clk), .CE(n516), .R(n525), .D(n163), .Q(rst_addr_r[6]));
Q_FDP4EP \rst_addr_r_REG[7] ( .CK(clk), .CE(n516), .R(n525), .D(n165), .Q(rst_addr_r[7]));
Q_FDP4EP \rst_addr_r_REG[8] ( .CK(clk), .CE(n516), .R(n525), .D(n167), .Q(rst_addr_r[8]));
Q_FDP4EP \inc_r_REG[0] ( .CK(clk), .CE(n514), .R(n525), .D(n168), .Q(inc_r[0]));
Q_FDP4EP \rd_dat_REG[0] ( .CK(clk), .CE(n512), .R(n525), .D(n169), .Q(rd_dat[0]));
Q_FDP4EP \rd_dat_REG[1] ( .CK(clk), .CE(n512), .R(n525), .D(n170), .Q(rd_dat[1]));
Q_FDP4EP \rd_dat_REG[2] ( .CK(clk), .CE(n512), .R(n525), .D(n171), .Q(rd_dat[2]));
Q_FDP4EP \rd_dat_REG[3] ( .CK(clk), .CE(n512), .R(n525), .D(n172), .Q(rd_dat[3]));
Q_FDP4EP \rd_dat_REG[4] ( .CK(clk), .CE(n512), .R(n525), .D(n173), .Q(rd_dat[4]));
Q_FDP4EP \rd_dat_REG[5] ( .CK(clk), .CE(n512), .R(n525), .D(n174), .Q(rd_dat[5]));
Q_FDP4EP \rd_dat_REG[6] ( .CK(clk), .CE(n512), .R(n525), .D(n175), .Q(rd_dat[6]));
Q_FDP4EP \rd_dat_REG[7] ( .CK(clk), .CE(n512), .R(n525), .D(n176), .Q(rd_dat[7]));
Q_FDP4EP \rd_dat_REG[8] ( .CK(clk), .CE(n512), .R(n525), .D(n177), .Q(rd_dat[8]));
Q_FDP4EP \rd_dat_REG[9] ( .CK(clk), .CE(n512), .R(n525), .D(n179), .Q(rd_dat[9]));
Q_FDP4EP \rd_dat_REG[10] ( .CK(clk), .CE(n512), .R(n525), .D(n181), .Q(rd_dat[10]));
Q_FDP4EP \rd_dat_REG[11] ( .CK(clk), .CE(n512), .R(n525), .D(n183), .Q(rd_dat[11]));
Q_FDP4EP \rd_dat_REG[12] ( .CK(clk), .CE(n512), .R(n525), .D(n185), .Q(rd_dat[12]));
Q_FDP4EP \rd_dat_REG[13] ( .CK(clk), .CE(n512), .R(n525), .D(n187), .Q(rd_dat[13]));
Q_FDP4EP \rd_dat_REG[14] ( .CK(clk), .CE(n512), .R(n525), .D(n189), .Q(rd_dat[14]));
Q_FDP4EP \rd_dat_REG[15] ( .CK(clk), .CE(n512), .R(n525), .D(n191), .Q(rd_dat[15]));
Q_FDP4EP \rd_dat_REG[16] ( .CK(clk), .CE(n512), .R(n525), .D(n193), .Q(rd_dat[16]));
Q_FDP4EP \rd_dat_REG[17] ( .CK(clk), .CE(n512), .R(n525), .D(n195), .Q(rd_dat[17]));
Q_FDP4EP \rd_dat_REG[18] ( .CK(clk), .CE(n512), .R(n525), .D(n197), .Q(rd_dat[18]));
Q_FDP4EP \rd_dat_REG[19] ( .CK(clk), .CE(n512), .R(n525), .D(n199), .Q(rd_dat[19]));
Q_FDP4EP \rd_dat_REG[20] ( .CK(clk), .CE(n512), .R(n525), .D(n201), .Q(rd_dat[20]));
Q_FDP4EP \rd_dat_REG[21] ( .CK(clk), .CE(n512), .R(n525), .D(n203), .Q(rd_dat[21]));
Q_FDP4EP \rd_dat_REG[22] ( .CK(clk), .CE(n512), .R(n525), .D(n205), .Q(rd_dat[22]));
Q_FDP4EP \rd_dat_REG[23] ( .CK(clk), .CE(n512), .R(n525), .D(n207), .Q(rd_dat[23]));
Q_FDP4EP \rd_dat_REG[24] ( .CK(clk), .CE(n512), .R(n525), .D(n209), .Q(rd_dat[24]));
Q_FDP4EP \rd_dat_REG[25] ( .CK(clk), .CE(n512), .R(n525), .D(n211), .Q(rd_dat[25]));
Q_FDP4EP \rd_dat_REG[26] ( .CK(clk), .CE(n512), .R(n525), .D(n213), .Q(rd_dat[26]));
Q_FDP4EP \rd_dat_REG[27] ( .CK(clk), .CE(n512), .R(n525), .D(n215), .Q(rd_dat[27]));
Q_FDP4EP \rd_dat_REG[28] ( .CK(clk), .CE(n512), .R(n525), .D(n217), .Q(rd_dat[28]));
Q_FDP4EP \rd_dat_REG[29] ( .CK(clk), .CE(n512), .R(n525), .D(n219), .Q(rd_dat[29]));
Q_FDP4EP \rd_dat_REG[30] ( .CK(clk), .CE(n512), .R(n525), .D(n221), .Q(rd_dat[30]));
Q_FDP4EP \rd_dat_REG[31] ( .CK(clk), .CE(n512), .R(n525), .D(n223), .Q(rd_dat[31]));
Q_FDP4EP \rd_dat_REG[32] ( .CK(clk), .CE(n512), .R(n525), .D(n225), .Q(rd_dat[32]));
Q_FDP4EP \rd_dat_REG[33] ( .CK(clk), .CE(n512), .R(n525), .D(n227), .Q(rd_dat[33]));
Q_FDP4EP \rd_dat_REG[34] ( .CK(clk), .CE(n512), .R(n525), .D(n229), .Q(rd_dat[34]));
Q_FDP4EP \rd_dat_REG[35] ( .CK(clk), .CE(n512), .R(n525), .D(n231), .Q(rd_dat[35]));
Q_FDP4EP \rd_dat_REG[36] ( .CK(clk), .CE(n512), .R(n525), .D(n233), .Q(rd_dat[36]));
Q_FDP4EP \rd_dat_REG[37] ( .CK(clk), .CE(n512), .R(n525), .D(n235), .Q(rd_dat[37]));
Q_FDP4EP \rd_dat_REG[38] ( .CK(clk), .CE(n512), .R(n525), .D(n237), .Q(rd_dat[38]));
Q_FDP4EP \rd_dat_REG[39] ( .CK(clk), .CE(n512), .R(n525), .D(n239), .Q(rd_dat[39]));
Q_FDP4EP \rd_dat_REG[40] ( .CK(clk), .CE(n512), .R(n525), .D(n241), .Q(rd_dat[40]));
Q_FDP4EP \rd_dat_REG[41] ( .CK(clk), .CE(n512), .R(n525), .D(n243), .Q(rd_dat[41]));
Q_FDP4EP \rd_dat_REG[42] ( .CK(clk), .CE(n512), .R(n525), .D(n245), .Q(rd_dat[42]));
Q_FDP4EP \rd_dat_REG[43] ( .CK(clk), .CE(n512), .R(n525), .D(n247), .Q(rd_dat[43]));
Q_FDP4EP \rd_dat_REG[44] ( .CK(clk), .CE(n512), .R(n525), .D(n249), .Q(rd_dat[44]));
Q_FDP4EP \rd_dat_REG[45] ( .CK(clk), .CE(n512), .R(n525), .D(n251), .Q(rd_dat[45]));
Q_FDP4EP \rd_dat_REG[46] ( .CK(clk), .CE(n512), .R(n525), .D(n253), .Q(rd_dat[46]));
Q_FDP4EP \rd_dat_REG[47] ( .CK(clk), .CE(n512), .R(n525), .D(n255), .Q(rd_dat[47]));
Q_FDP4EP \rd_dat_REG[48] ( .CK(clk), .CE(n512), .R(n525), .D(n257), .Q(rd_dat[48]));
Q_FDP4EP \rd_dat_REG[49] ( .CK(clk), .CE(n512), .R(n525), .D(n259), .Q(rd_dat[49]));
Q_FDP4EP \rd_dat_REG[50] ( .CK(clk), .CE(n512), .R(n525), .D(n261), .Q(rd_dat[50]));
Q_FDP4EP \rd_dat_REG[51] ( .CK(clk), .CE(n512), .R(n525), .D(n263), .Q(rd_dat[51]));
Q_FDP4EP \rd_dat_REG[52] ( .CK(clk), .CE(n512), .R(n525), .D(n265), .Q(rd_dat[52]));
Q_FDP4EP \rd_dat_REG[53] ( .CK(clk), .CE(n512), .R(n525), .D(n267), .Q(rd_dat[53]));
Q_FDP4EP \rd_dat_REG[54] ( .CK(clk), .CE(n512), .R(n525), .D(n269), .Q(rd_dat[54]));
Q_FDP4EP \rd_dat_REG[55] ( .CK(clk), .CE(n512), .R(n525), .D(n271), .Q(rd_dat[55]));
Q_FDP4EP \rd_dat_REG[56] ( .CK(clk), .CE(n512), .R(n525), .D(n273), .Q(rd_dat[56]));
Q_FDP4EP \rd_dat_REG[57] ( .CK(clk), .CE(n512), .R(n525), .D(n275), .Q(rd_dat[57]));
Q_FDP4EP \rd_dat_REG[58] ( .CK(clk), .CE(n512), .R(n525), .D(n277), .Q(rd_dat[58]));
Q_FDP4EP \rd_dat_REG[59] ( .CK(clk), .CE(n512), .R(n525), .D(n279), .Q(rd_dat[59]));
Q_FDP4EP \rd_dat_REG[60] ( .CK(clk), .CE(n512), .R(n525), .D(n281), .Q(rd_dat[60]));
Q_FDP4EP \rd_dat_REG[61] ( .CK(clk), .CE(n512), .R(n525), .D(n283), .Q(rd_dat[61]));
Q_FDP4EP \rd_dat_REG[62] ( .CK(clk), .CE(n512), .R(n525), .D(n285), .Q(rd_dat[62]));
Q_FDP4EP \rd_dat_REG[63] ( .CK(clk), .CE(n512), .R(n525), .D(n287), .Q(rd_dat[63]));
Q_FDP4EP \rd_dat_REG[64] ( .CK(clk), .CE(n512), .R(n525), .D(n289), .Q(rd_dat[64]));
Q_FDP4EP \rd_dat_REG[65] ( .CK(clk), .CE(n512), .R(n525), .D(n291), .Q(rd_dat[65]));
Q_FDP4EP \rd_dat_REG[66] ( .CK(clk), .CE(n512), .R(n525), .D(n293), .Q(rd_dat[66]));
Q_FDP4EP \rd_dat_REG[67] ( .CK(clk), .CE(n512), .R(n525), .D(n295), .Q(rd_dat[67]));
Q_FDP4EP \rd_dat_REG[68] ( .CK(clk), .CE(n512), .R(n525), .D(n297), .Q(rd_dat[68]));
Q_FDP4EP \rd_dat_REG[69] ( .CK(clk), .CE(n512), .R(n525), .D(n299), .Q(rd_dat[69]));
Q_FDP4EP \rd_dat_REG[70] ( .CK(clk), .CE(n512), .R(n525), .D(n301), .Q(rd_dat[70]));
Q_FDP4EP \rd_dat_REG[71] ( .CK(clk), .CE(n512), .R(n525), .D(n303), .Q(rd_dat[71]));
Q_FDP4EP \rd_dat_REG[72] ( .CK(clk), .CE(n512), .R(n525), .D(n305), .Q(rd_dat[72]));
Q_FDP4EP \rd_dat_REG[73] ( .CK(clk), .CE(n512), .R(n525), .D(n307), .Q(rd_dat[73]));
Q_FDP4EP \rd_dat_REG[74] ( .CK(clk), .CE(n512), .R(n525), .D(n309), .Q(rd_dat[74]));
Q_FDP4EP \rd_dat_REG[75] ( .CK(clk), .CE(n512), .R(n525), .D(n311), .Q(rd_dat[75]));
Q_FDP4EP \rd_dat_REG[76] ( .CK(clk), .CE(n512), .R(n525), .D(n313), .Q(rd_dat[76]));
Q_FDP4EP \rd_dat_REG[77] ( .CK(clk), .CE(n512), .R(n525), .D(n315), .Q(rd_dat[77]));
Q_FDP4EP \rd_dat_REG[78] ( .CK(clk), .CE(n512), .R(n525), .D(n317), .Q(rd_dat[78]));
Q_FDP4EP \rd_dat_REG[79] ( .CK(clk), .CE(n512), .R(n525), .D(n319), .Q(rd_dat[79]));
Q_FDP4EP \rd_dat_REG[80] ( .CK(clk), .CE(n512), .R(n525), .D(n321), .Q(rd_dat[80]));
Q_FDP4EP \rd_dat_REG[81] ( .CK(clk), .CE(n512), .R(n525), .D(n323), .Q(rd_dat[81]));
Q_FDP4EP \rd_dat_REG[82] ( .CK(clk), .CE(n512), .R(n525), .D(n325), .Q(rd_dat[82]));
Q_FDP4EP \rd_dat_REG[83] ( .CK(clk), .CE(n512), .R(n525), .D(n327), .Q(rd_dat[83]));
Q_FDP4EP \rd_dat_REG[84] ( .CK(clk), .CE(n512), .R(n525), .D(n329), .Q(rd_dat[84]));
Q_FDP4EP \rd_dat_REG[85] ( .CK(clk), .CE(n512), .R(n525), .D(n331), .Q(rd_dat[85]));
Q_FDP4EP \rd_dat_REG[86] ( .CK(clk), .CE(n512), .R(n525), .D(n333), .Q(rd_dat[86]));
Q_FDP4EP \rd_dat_REG[87] ( .CK(clk), .CE(n512), .R(n525), .D(n335), .Q(rd_dat[87]));
Q_FDP4EP \rd_dat_REG[88] ( .CK(clk), .CE(n512), .R(n525), .D(n337), .Q(rd_dat[88]));
Q_FDP4EP \rd_dat_REG[89] ( .CK(clk), .CE(n512), .R(n525), .D(n339), .Q(rd_dat[89]));
Q_FDP4EP \rd_dat_REG[90] ( .CK(clk), .CE(n512), .R(n525), .D(n341), .Q(rd_dat[90]));
Q_FDP4EP \rd_dat_REG[91] ( .CK(clk), .CE(n512), .R(n525), .D(n343), .Q(rd_dat[91]));
Q_FDP4EP \rd_dat_REG[92] ( .CK(clk), .CE(n512), .R(n525), .D(n345), .Q(rd_dat[92]));
Q_FDP4EP \rd_dat_REG[93] ( .CK(clk), .CE(n512), .R(n525), .D(n347), .Q(rd_dat[93]));
Q_FDP4EP \rd_dat_REG[94] ( .CK(clk), .CE(n512), .R(n525), .D(n349), .Q(rd_dat[94]));
Q_FDP4EP \rd_dat_REG[95] ( .CK(clk), .CE(n512), .R(n525), .D(n351), .Q(rd_dat[95]));
Q_INV U811 ( .A(n515), .Z(n526));
Q_FDP4EP init_inc_r_REG  ( .CK(clk), .CE(n526), .R(n525), .D(n1), .Q(init_inc_r));
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "addr_limit (2,0) 1 8 0 0 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "1"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_1 "-1 genblk2  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_0 "-1 genblk1  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "genblk2"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "genblk1"
endmodule
