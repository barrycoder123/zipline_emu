
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
(* celldefine = 1 *) 
module nx_ram_1rw_xcm109 ( clk, rst_n, ovstb, lvm, mlvm, mrdten, bimc_rst_n, 
	bimc_isync, bimc_idat, bimc_odat, bimc_osync, 
	ro_uncorrectable_ecc_error, bwe, din, add, cs, we, dout);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
input clk;
input rst_n;
input ovstb;
input lvm;
input mlvm;
input mrdten;
input bimc_rst_n;
input bimc_isync;
input bimc_idat;
output bimc_odat;
output bimc_osync;
output ro_uncorrectable_ecc_error;
input [63:0] bwe;
input [63:0] din;
input [14:0] add;
input cs;
input we;
output [63:0] dout;
wire _zy_simnet_bimc_odat_0_w$;
wire _zy_simnet_bimc_osync_1_w$;
wire _zy_simnet_ro_uncorrectable_ecc_error_2_w$;
wire bimc_iclk;
wire bimc_irstn;
wire rst_clk_n;
wire p_mode_disable_ecc_mem;
wire byp;
wire se;
wire rds;
wire [1:0] ecc_corrupt;
wire rst_rclk_n;
wire sew;
wire web;
wire ro_mem_ecc_error_ev;
wire ro_mem_ecc_corrected;
wire [14:0] ro_mem_ecc_error_addr;
wire [63:0] \g.dout_i ;
wire [63:0] \g.dat_r ;
wire [63:0] \g.din_i ;
wire [32767:0] \g.we_clk ;
wire [31:0] \g.u_ram._zyictd_sysfunc_11_L263_9 ;
wire [32767:0] \g.we_gate ;
wire [14:0] \g.add_r ;
supply0 n217;
Q_BUF U0 ( .A(n217), .Z(p_mode_disable_ecc_mem));
Q_BUF U1 ( .A(n217), .Z(byp));
Q_BUF U2 ( .A(n217), .Z(se));
Q_BUF U3 ( .A(n217), .Z(rds));
Q_BUF U4 ( .A(n217), .Z(ecc_corrupt[1]));
Q_BUF U5 ( .A(n217), .Z(ecc_corrupt[0]));
Q_BUF U6 ( .A(n217), .Z(sew));
Q_ASSIGN U7 ( .B(clk), .A(\g.we_clk [32767]));
Q_ASSIGN U8 ( .B(clk), .A(\g.we_clk [32766]));
Q_ASSIGN U9 ( .B(clk), .A(\g.we_clk [32765]));
Q_ASSIGN U10 ( .B(clk), .A(\g.we_clk [32764]));
Q_ASSIGN U11 ( .B(clk), .A(\g.we_clk [32763]));
Q_ASSIGN U12 ( .B(clk), .A(\g.we_clk [32762]));
Q_ASSIGN U13 ( .B(clk), .A(\g.we_clk [32761]));
Q_ASSIGN U14 ( .B(clk), .A(\g.we_clk [32760]));
Q_ASSIGN U15 ( .B(clk), .A(\g.we_clk [32759]));
Q_ASSIGN U16 ( .B(clk), .A(\g.we_clk [32758]));
Q_ASSIGN U17 ( .B(clk), .A(\g.we_clk [32757]));
Q_ASSIGN U18 ( .B(clk), .A(\g.we_clk [32756]));
Q_ASSIGN U19 ( .B(clk), .A(\g.we_clk [32755]));
Q_ASSIGN U20 ( .B(clk), .A(\g.we_clk [32754]));
Q_ASSIGN U21 ( .B(clk), .A(\g.we_clk [32753]));
Q_ASSIGN U22 ( .B(clk), .A(\g.we_clk [32752]));
Q_ASSIGN U23 ( .B(clk), .A(\g.we_clk [32751]));
Q_ASSIGN U24 ( .B(clk), .A(\g.we_clk [32750]));
Q_ASSIGN U25 ( .B(clk), .A(\g.we_clk [32749]));
Q_ASSIGN U26 ( .B(clk), .A(\g.we_clk [32748]));
Q_ASSIGN U27 ( .B(clk), .A(\g.we_clk [32747]));
Q_ASSIGN U28 ( .B(clk), .A(\g.we_clk [32746]));
Q_ASSIGN U29 ( .B(clk), .A(\g.we_clk [32745]));
Q_ASSIGN U30 ( .B(clk), .A(\g.we_clk [32744]));
Q_ASSIGN U31 ( .B(clk), .A(\g.we_clk [32743]));
Q_ASSIGN U32 ( .B(clk), .A(\g.we_clk [32742]));
Q_ASSIGN U33 ( .B(clk), .A(\g.we_clk [32741]));
Q_ASSIGN U34 ( .B(clk), .A(\g.we_clk [32740]));
Q_ASSIGN U35 ( .B(clk), .A(\g.we_clk [32739]));
Q_ASSIGN U36 ( .B(clk), .A(\g.we_clk [32738]));
Q_ASSIGN U37 ( .B(clk), .A(\g.we_clk [32737]));
Q_ASSIGN U38 ( .B(clk), .A(\g.we_clk [32736]));
Q_ASSIGN U39 ( .B(clk), .A(\g.we_clk [32735]));
Q_ASSIGN U40 ( .B(clk), .A(\g.we_clk [32734]));
Q_ASSIGN U41 ( .B(clk), .A(\g.we_clk [32733]));
Q_ASSIGN U42 ( .B(clk), .A(\g.we_clk [32732]));
Q_ASSIGN U43 ( .B(clk), .A(\g.we_clk [32731]));
Q_ASSIGN U44 ( .B(clk), .A(\g.we_clk [32730]));
Q_ASSIGN U45 ( .B(clk), .A(\g.we_clk [32729]));
Q_ASSIGN U46 ( .B(clk), .A(\g.we_clk [32728]));
Q_ASSIGN U47 ( .B(clk), .A(\g.we_clk [32727]));
Q_ASSIGN U48 ( .B(clk), .A(\g.we_clk [32726]));
Q_ASSIGN U49 ( .B(clk), .A(\g.we_clk [32725]));
Q_ASSIGN U50 ( .B(clk), .A(\g.we_clk [32724]));
Q_ASSIGN U51 ( .B(clk), .A(\g.we_clk [32723]));
Q_ASSIGN U52 ( .B(clk), .A(\g.we_clk [32722]));
Q_ASSIGN U53 ( .B(clk), .A(\g.we_clk [32721]));
Q_ASSIGN U54 ( .B(clk), .A(\g.we_clk [32720]));
Q_ASSIGN U55 ( .B(clk), .A(\g.we_clk [32719]));
Q_ASSIGN U56 ( .B(clk), .A(\g.we_clk [32718]));
Q_ASSIGN U57 ( .B(clk), .A(\g.we_clk [32717]));
Q_ASSIGN U58 ( .B(clk), .A(\g.we_clk [32716]));
Q_ASSIGN U59 ( .B(clk), .A(\g.we_clk [32715]));
Q_ASSIGN U60 ( .B(clk), .A(\g.we_clk [32714]));
Q_ASSIGN U61 ( .B(clk), .A(\g.we_clk [32713]));
Q_ASSIGN U62 ( .B(clk), .A(\g.we_clk [32712]));
Q_ASSIGN U63 ( .B(clk), .A(\g.we_clk [32711]));
Q_ASSIGN U64 ( .B(clk), .A(\g.we_clk [32710]));
Q_ASSIGN U65 ( .B(clk), .A(\g.we_clk [32709]));
Q_ASSIGN U66 ( .B(clk), .A(\g.we_clk [32708]));
Q_ASSIGN U67 ( .B(clk), .A(\g.we_clk [32707]));
Q_ASSIGN U68 ( .B(clk), .A(\g.we_clk [32706]));
Q_ASSIGN U69 ( .B(clk), .A(\g.we_clk [32705]));
Q_ASSIGN U70 ( .B(clk), .A(\g.we_clk [32704]));
Q_ASSIGN U71 ( .B(clk), .A(\g.we_clk [32703]));
Q_ASSIGN U72 ( .B(clk), .A(\g.we_clk [32702]));
Q_ASSIGN U73 ( .B(clk), .A(\g.we_clk [32701]));
Q_ASSIGN U74 ( .B(clk), .A(\g.we_clk [32700]));
Q_ASSIGN U75 ( .B(clk), .A(\g.we_clk [32699]));
Q_ASSIGN U76 ( .B(clk), .A(\g.we_clk [32698]));
Q_ASSIGN U77 ( .B(clk), .A(\g.we_clk [32697]));
Q_ASSIGN U78 ( .B(clk), .A(\g.we_clk [32696]));
Q_ASSIGN U79 ( .B(clk), .A(\g.we_clk [32695]));
Q_ASSIGN U80 ( .B(clk), .A(\g.we_clk [32694]));
Q_ASSIGN U81 ( .B(clk), .A(\g.we_clk [32693]));
Q_ASSIGN U82 ( .B(clk), .A(\g.we_clk [32692]));
Q_ASSIGN U83 ( .B(clk), .A(\g.we_clk [32691]));
Q_ASSIGN U84 ( .B(clk), .A(\g.we_clk [32690]));
Q_ASSIGN U85 ( .B(clk), .A(\g.we_clk [32689]));
Q_ASSIGN U86 ( .B(clk), .A(\g.we_clk [32688]));
Q_ASSIGN U87 ( .B(clk), .A(\g.we_clk [32687]));
Q_ASSIGN U88 ( .B(clk), .A(\g.we_clk [32686]));
Q_ASSIGN U89 ( .B(clk), .A(\g.we_clk [32685]));
Q_ASSIGN U90 ( .B(clk), .A(\g.we_clk [32684]));
Q_ASSIGN U91 ( .B(clk), .A(\g.we_clk [32683]));
Q_ASSIGN U92 ( .B(clk), .A(\g.we_clk [32682]));
Q_ASSIGN U93 ( .B(clk), .A(\g.we_clk [32681]));
Q_ASSIGN U94 ( .B(clk), .A(\g.we_clk [32680]));
Q_ASSIGN U95 ( .B(clk), .A(\g.we_clk [32679]));
Q_ASSIGN U96 ( .B(clk), .A(\g.we_clk [32678]));
Q_ASSIGN U97 ( .B(clk), .A(\g.we_clk [32677]));
Q_ASSIGN U98 ( .B(clk), .A(\g.we_clk [32676]));
Q_ASSIGN U99 ( .B(clk), .A(\g.we_clk [32675]));
Q_ASSIGN U100 ( .B(clk), .A(\g.we_clk [32674]));
Q_ASSIGN U101 ( .B(clk), .A(\g.we_clk [32673]));
Q_ASSIGN U102 ( .B(clk), .A(\g.we_clk [32672]));
Q_ASSIGN U103 ( .B(clk), .A(\g.we_clk [32671]));
Q_ASSIGN U104 ( .B(clk), .A(\g.we_clk [32670]));
Q_ASSIGN U105 ( .B(clk), .A(\g.we_clk [32669]));
Q_ASSIGN U106 ( .B(clk), .A(\g.we_clk [32668]));
Q_ASSIGN U107 ( .B(clk), .A(\g.we_clk [32667]));
Q_ASSIGN U108 ( .B(clk), .A(\g.we_clk [32666]));
Q_ASSIGN U109 ( .B(clk), .A(\g.we_clk [32665]));
Q_ASSIGN U110 ( .B(clk), .A(\g.we_clk [32664]));
Q_ASSIGN U111 ( .B(clk), .A(\g.we_clk [32663]));
Q_ASSIGN U112 ( .B(clk), .A(\g.we_clk [32662]));
Q_ASSIGN U113 ( .B(clk), .A(\g.we_clk [32661]));
Q_ASSIGN U114 ( .B(clk), .A(\g.we_clk [32660]));
Q_ASSIGN U115 ( .B(clk), .A(\g.we_clk [32659]));
Q_ASSIGN U116 ( .B(clk), .A(\g.we_clk [32658]));
Q_ASSIGN U117 ( .B(clk), .A(\g.we_clk [32657]));
Q_ASSIGN U118 ( .B(clk), .A(\g.we_clk [32656]));
Q_ASSIGN U119 ( .B(clk), .A(\g.we_clk [32655]));
Q_ASSIGN U120 ( .B(clk), .A(\g.we_clk [32654]));
Q_ASSIGN U121 ( .B(clk), .A(\g.we_clk [32653]));
Q_ASSIGN U122 ( .B(clk), .A(\g.we_clk [32652]));
Q_ASSIGN U123 ( .B(clk), .A(\g.we_clk [32651]));
Q_ASSIGN U124 ( .B(clk), .A(\g.we_clk [32650]));
Q_ASSIGN U125 ( .B(clk), .A(\g.we_clk [32649]));
Q_ASSIGN U126 ( .B(clk), .A(\g.we_clk [32648]));
Q_ASSIGN U127 ( .B(clk), .A(\g.we_clk [32647]));
Q_ASSIGN U128 ( .B(clk), .A(\g.we_clk [32646]));
Q_ASSIGN U129 ( .B(clk), .A(\g.we_clk [32645]));
Q_ASSIGN U130 ( .B(clk), .A(\g.we_clk [32644]));
Q_ASSIGN U131 ( .B(clk), .A(\g.we_clk [32643]));
Q_ASSIGN U132 ( .B(clk), .A(\g.we_clk [32642]));
Q_ASSIGN U133 ( .B(clk), .A(\g.we_clk [32641]));
Q_ASSIGN U134 ( .B(clk), .A(\g.we_clk [32640]));
Q_ASSIGN U135 ( .B(clk), .A(\g.we_clk [32639]));
Q_ASSIGN U136 ( .B(clk), .A(\g.we_clk [32638]));
Q_ASSIGN U137 ( .B(clk), .A(\g.we_clk [32637]));
Q_ASSIGN U138 ( .B(clk), .A(\g.we_clk [32636]));
Q_ASSIGN U139 ( .B(clk), .A(\g.we_clk [32635]));
Q_ASSIGN U140 ( .B(clk), .A(\g.we_clk [32634]));
Q_ASSIGN U141 ( .B(clk), .A(\g.we_clk [32633]));
Q_ASSIGN U142 ( .B(clk), .A(\g.we_clk [32632]));
Q_ASSIGN U143 ( .B(clk), .A(\g.we_clk [32631]));
Q_ASSIGN U144 ( .B(clk), .A(\g.we_clk [32630]));
Q_ASSIGN U145 ( .B(clk), .A(\g.we_clk [32629]));
Q_ASSIGN U146 ( .B(clk), .A(\g.we_clk [32628]));
Q_ASSIGN U147 ( .B(clk), .A(\g.we_clk [32627]));
Q_ASSIGN U148 ( .B(clk), .A(\g.we_clk [32626]));
Q_ASSIGN U149 ( .B(clk), .A(\g.we_clk [32625]));
Q_ASSIGN U150 ( .B(clk), .A(\g.we_clk [32624]));
Q_ASSIGN U151 ( .B(clk), .A(\g.we_clk [32623]));
Q_ASSIGN U152 ( .B(clk), .A(\g.we_clk [32622]));
Q_ASSIGN U153 ( .B(clk), .A(\g.we_clk [32621]));
Q_ASSIGN U154 ( .B(clk), .A(\g.we_clk [32620]));
Q_ASSIGN U155 ( .B(clk), .A(\g.we_clk [32619]));
Q_ASSIGN U156 ( .B(clk), .A(\g.we_clk [32618]));
Q_ASSIGN U157 ( .B(clk), .A(\g.we_clk [32617]));
Q_ASSIGN U158 ( .B(clk), .A(\g.we_clk [32616]));
Q_ASSIGN U159 ( .B(clk), .A(\g.we_clk [32615]));
Q_ASSIGN U160 ( .B(clk), .A(\g.we_clk [32614]));
Q_ASSIGN U161 ( .B(clk), .A(\g.we_clk [32613]));
Q_ASSIGN U162 ( .B(clk), .A(\g.we_clk [32612]));
Q_ASSIGN U163 ( .B(clk), .A(\g.we_clk [32611]));
Q_ASSIGN U164 ( .B(clk), .A(\g.we_clk [32610]));
Q_ASSIGN U165 ( .B(clk), .A(\g.we_clk [32609]));
Q_ASSIGN U166 ( .B(clk), .A(\g.we_clk [32608]));
Q_ASSIGN U167 ( .B(clk), .A(\g.we_clk [32607]));
Q_ASSIGN U168 ( .B(clk), .A(\g.we_clk [32606]));
Q_ASSIGN U169 ( .B(clk), .A(\g.we_clk [32605]));
Q_ASSIGN U170 ( .B(clk), .A(\g.we_clk [32604]));
Q_ASSIGN U171 ( .B(clk), .A(\g.we_clk [32603]));
Q_ASSIGN U172 ( .B(clk), .A(\g.we_clk [32602]));
Q_ASSIGN U173 ( .B(clk), .A(\g.we_clk [32601]));
Q_ASSIGN U174 ( .B(clk), .A(\g.we_clk [32600]));
Q_ASSIGN U175 ( .B(clk), .A(\g.we_clk [32599]));
Q_ASSIGN U176 ( .B(clk), .A(\g.we_clk [32598]));
Q_ASSIGN U177 ( .B(clk), .A(\g.we_clk [32597]));
Q_ASSIGN U178 ( .B(clk), .A(\g.we_clk [32596]));
Q_ASSIGN U179 ( .B(clk), .A(\g.we_clk [32595]));
Q_ASSIGN U180 ( .B(clk), .A(\g.we_clk [32594]));
Q_ASSIGN U181 ( .B(clk), .A(\g.we_clk [32593]));
Q_ASSIGN U182 ( .B(clk), .A(\g.we_clk [32592]));
Q_ASSIGN U183 ( .B(clk), .A(\g.we_clk [32591]));
Q_ASSIGN U184 ( .B(clk), .A(\g.we_clk [32590]));
Q_ASSIGN U185 ( .B(clk), .A(\g.we_clk [32589]));
Q_ASSIGN U186 ( .B(clk), .A(\g.we_clk [32588]));
Q_ASSIGN U187 ( .B(clk), .A(\g.we_clk [32587]));
Q_ASSIGN U188 ( .B(clk), .A(\g.we_clk [32586]));
Q_ASSIGN U189 ( .B(clk), .A(\g.we_clk [32585]));
Q_ASSIGN U190 ( .B(clk), .A(\g.we_clk [32584]));
Q_ASSIGN U191 ( .B(clk), .A(\g.we_clk [32583]));
Q_ASSIGN U192 ( .B(clk), .A(\g.we_clk [32582]));
Q_ASSIGN U193 ( .B(clk), .A(\g.we_clk [32581]));
Q_ASSIGN U194 ( .B(clk), .A(\g.we_clk [32580]));
Q_ASSIGN U195 ( .B(clk), .A(\g.we_clk [32579]));
Q_ASSIGN U196 ( .B(clk), .A(\g.we_clk [32578]));
Q_ASSIGN U197 ( .B(clk), .A(\g.we_clk [32577]));
Q_ASSIGN U198 ( .B(clk), .A(\g.we_clk [32576]));
Q_ASSIGN U199 ( .B(clk), .A(\g.we_clk [32575]));
Q_ASSIGN U200 ( .B(clk), .A(\g.we_clk [32574]));
Q_ASSIGN U201 ( .B(clk), .A(\g.we_clk [32573]));
Q_ASSIGN U202 ( .B(clk), .A(\g.we_clk [32572]));
Q_ASSIGN U203 ( .B(clk), .A(\g.we_clk [32571]));
Q_ASSIGN U204 ( .B(clk), .A(\g.we_clk [32570]));
Q_ASSIGN U205 ( .B(clk), .A(\g.we_clk [32569]));
Q_ASSIGN U206 ( .B(clk), .A(\g.we_clk [32568]));
Q_ASSIGN U207 ( .B(clk), .A(\g.we_clk [32567]));
Q_ASSIGN U208 ( .B(clk), .A(\g.we_clk [32566]));
Q_ASSIGN U209 ( .B(clk), .A(\g.we_clk [32565]));
Q_ASSIGN U210 ( .B(clk), .A(\g.we_clk [32564]));
Q_ASSIGN U211 ( .B(clk), .A(\g.we_clk [32563]));
Q_ASSIGN U212 ( .B(clk), .A(\g.we_clk [32562]));
Q_ASSIGN U213 ( .B(clk), .A(\g.we_clk [32561]));
Q_ASSIGN U214 ( .B(clk), .A(\g.we_clk [32560]));
Q_ASSIGN U215 ( .B(clk), .A(\g.we_clk [32559]));
Q_ASSIGN U216 ( .B(clk), .A(\g.we_clk [32558]));
Q_ASSIGN U217 ( .B(clk), .A(\g.we_clk [32557]));
Q_ASSIGN U218 ( .B(clk), .A(\g.we_clk [32556]));
Q_ASSIGN U219 ( .B(clk), .A(\g.we_clk [32555]));
Q_ASSIGN U220 ( .B(clk), .A(\g.we_clk [32554]));
Q_ASSIGN U221 ( .B(clk), .A(\g.we_clk [32553]));
Q_ASSIGN U222 ( .B(clk), .A(\g.we_clk [32552]));
Q_ASSIGN U223 ( .B(clk), .A(\g.we_clk [32551]));
Q_ASSIGN U224 ( .B(clk), .A(\g.we_clk [32550]));
Q_ASSIGN U225 ( .B(clk), .A(\g.we_clk [32549]));
Q_ASSIGN U226 ( .B(clk), .A(\g.we_clk [32548]));
Q_ASSIGN U227 ( .B(clk), .A(\g.we_clk [32547]));
Q_ASSIGN U228 ( .B(clk), .A(\g.we_clk [32546]));
Q_ASSIGN U229 ( .B(clk), .A(\g.we_clk [32545]));
Q_ASSIGN U230 ( .B(clk), .A(\g.we_clk [32544]));
Q_ASSIGN U231 ( .B(clk), .A(\g.we_clk [32543]));
Q_ASSIGN U232 ( .B(clk), .A(\g.we_clk [32542]));
Q_ASSIGN U233 ( .B(clk), .A(\g.we_clk [32541]));
Q_ASSIGN U234 ( .B(clk), .A(\g.we_clk [32540]));
Q_ASSIGN U235 ( .B(clk), .A(\g.we_clk [32539]));
Q_ASSIGN U236 ( .B(clk), .A(\g.we_clk [32538]));
Q_ASSIGN U237 ( .B(clk), .A(\g.we_clk [32537]));
Q_ASSIGN U238 ( .B(clk), .A(\g.we_clk [32536]));
Q_ASSIGN U239 ( .B(clk), .A(\g.we_clk [32535]));
Q_ASSIGN U240 ( .B(clk), .A(\g.we_clk [32534]));
Q_ASSIGN U241 ( .B(clk), .A(\g.we_clk [32533]));
Q_ASSIGN U242 ( .B(clk), .A(\g.we_clk [32532]));
Q_ASSIGN U243 ( .B(clk), .A(\g.we_clk [32531]));
Q_ASSIGN U244 ( .B(clk), .A(\g.we_clk [32530]));
Q_ASSIGN U245 ( .B(clk), .A(\g.we_clk [32529]));
Q_ASSIGN U246 ( .B(clk), .A(\g.we_clk [32528]));
Q_ASSIGN U247 ( .B(clk), .A(\g.we_clk [32527]));
Q_ASSIGN U248 ( .B(clk), .A(\g.we_clk [32526]));
Q_ASSIGN U249 ( .B(clk), .A(\g.we_clk [32525]));
Q_ASSIGN U250 ( .B(clk), .A(\g.we_clk [32524]));
Q_ASSIGN U251 ( .B(clk), .A(\g.we_clk [32523]));
Q_ASSIGN U252 ( .B(clk), .A(\g.we_clk [32522]));
Q_ASSIGN U253 ( .B(clk), .A(\g.we_clk [32521]));
Q_ASSIGN U254 ( .B(clk), .A(\g.we_clk [32520]));
Q_ASSIGN U255 ( .B(clk), .A(\g.we_clk [32519]));
Q_ASSIGN U256 ( .B(clk), .A(\g.we_clk [32518]));
Q_ASSIGN U257 ( .B(clk), .A(\g.we_clk [32517]));
Q_ASSIGN U258 ( .B(clk), .A(\g.we_clk [32516]));
Q_ASSIGN U259 ( .B(clk), .A(\g.we_clk [32515]));
Q_ASSIGN U260 ( .B(clk), .A(\g.we_clk [32514]));
Q_ASSIGN U261 ( .B(clk), .A(\g.we_clk [32513]));
Q_ASSIGN U262 ( .B(clk), .A(\g.we_clk [32512]));
Q_ASSIGN U263 ( .B(clk), .A(\g.we_clk [32511]));
Q_ASSIGN U264 ( .B(clk), .A(\g.we_clk [32510]));
Q_ASSIGN U265 ( .B(clk), .A(\g.we_clk [32509]));
Q_ASSIGN U266 ( .B(clk), .A(\g.we_clk [32508]));
Q_ASSIGN U267 ( .B(clk), .A(\g.we_clk [32507]));
Q_ASSIGN U268 ( .B(clk), .A(\g.we_clk [32506]));
Q_ASSIGN U269 ( .B(clk), .A(\g.we_clk [32505]));
Q_ASSIGN U270 ( .B(clk), .A(\g.we_clk [32504]));
Q_ASSIGN U271 ( .B(clk), .A(\g.we_clk [32503]));
Q_ASSIGN U272 ( .B(clk), .A(\g.we_clk [32502]));
Q_ASSIGN U273 ( .B(clk), .A(\g.we_clk [32501]));
Q_ASSIGN U274 ( .B(clk), .A(\g.we_clk [32500]));
Q_ASSIGN U275 ( .B(clk), .A(\g.we_clk [32499]));
Q_ASSIGN U276 ( .B(clk), .A(\g.we_clk [32498]));
Q_ASSIGN U277 ( .B(clk), .A(\g.we_clk [32497]));
Q_ASSIGN U278 ( .B(clk), .A(\g.we_clk [32496]));
Q_ASSIGN U279 ( .B(clk), .A(\g.we_clk [32495]));
Q_ASSIGN U280 ( .B(clk), .A(\g.we_clk [32494]));
Q_ASSIGN U281 ( .B(clk), .A(\g.we_clk [32493]));
Q_ASSIGN U282 ( .B(clk), .A(\g.we_clk [32492]));
Q_ASSIGN U283 ( .B(clk), .A(\g.we_clk [32491]));
Q_ASSIGN U284 ( .B(clk), .A(\g.we_clk [32490]));
Q_ASSIGN U285 ( .B(clk), .A(\g.we_clk [32489]));
Q_ASSIGN U286 ( .B(clk), .A(\g.we_clk [32488]));
Q_ASSIGN U287 ( .B(clk), .A(\g.we_clk [32487]));
Q_ASSIGN U288 ( .B(clk), .A(\g.we_clk [32486]));
Q_ASSIGN U289 ( .B(clk), .A(\g.we_clk [32485]));
Q_ASSIGN U290 ( .B(clk), .A(\g.we_clk [32484]));
Q_ASSIGN U291 ( .B(clk), .A(\g.we_clk [32483]));
Q_ASSIGN U292 ( .B(clk), .A(\g.we_clk [32482]));
Q_ASSIGN U293 ( .B(clk), .A(\g.we_clk [32481]));
Q_ASSIGN U294 ( .B(clk), .A(\g.we_clk [32480]));
Q_ASSIGN U295 ( .B(clk), .A(\g.we_clk [32479]));
Q_ASSIGN U296 ( .B(clk), .A(\g.we_clk [32478]));
Q_ASSIGN U297 ( .B(clk), .A(\g.we_clk [32477]));
Q_ASSIGN U298 ( .B(clk), .A(\g.we_clk [32476]));
Q_ASSIGN U299 ( .B(clk), .A(\g.we_clk [32475]));
Q_ASSIGN U300 ( .B(clk), .A(\g.we_clk [32474]));
Q_ASSIGN U301 ( .B(clk), .A(\g.we_clk [32473]));
Q_ASSIGN U302 ( .B(clk), .A(\g.we_clk [32472]));
Q_ASSIGN U303 ( .B(clk), .A(\g.we_clk [32471]));
Q_ASSIGN U304 ( .B(clk), .A(\g.we_clk [32470]));
Q_ASSIGN U305 ( .B(clk), .A(\g.we_clk [32469]));
Q_ASSIGN U306 ( .B(clk), .A(\g.we_clk [32468]));
Q_ASSIGN U307 ( .B(clk), .A(\g.we_clk [32467]));
Q_ASSIGN U308 ( .B(clk), .A(\g.we_clk [32466]));
Q_ASSIGN U309 ( .B(clk), .A(\g.we_clk [32465]));
Q_ASSIGN U310 ( .B(clk), .A(\g.we_clk [32464]));
Q_ASSIGN U311 ( .B(clk), .A(\g.we_clk [32463]));
Q_ASSIGN U312 ( .B(clk), .A(\g.we_clk [32462]));
Q_ASSIGN U313 ( .B(clk), .A(\g.we_clk [32461]));
Q_ASSIGN U314 ( .B(clk), .A(\g.we_clk [32460]));
Q_ASSIGN U315 ( .B(clk), .A(\g.we_clk [32459]));
Q_ASSIGN U316 ( .B(clk), .A(\g.we_clk [32458]));
Q_ASSIGN U317 ( .B(clk), .A(\g.we_clk [32457]));
Q_ASSIGN U318 ( .B(clk), .A(\g.we_clk [32456]));
Q_ASSIGN U319 ( .B(clk), .A(\g.we_clk [32455]));
Q_ASSIGN U320 ( .B(clk), .A(\g.we_clk [32454]));
Q_ASSIGN U321 ( .B(clk), .A(\g.we_clk [32453]));
Q_ASSIGN U322 ( .B(clk), .A(\g.we_clk [32452]));
Q_ASSIGN U323 ( .B(clk), .A(\g.we_clk [32451]));
Q_ASSIGN U324 ( .B(clk), .A(\g.we_clk [32450]));
Q_ASSIGN U325 ( .B(clk), .A(\g.we_clk [32449]));
Q_ASSIGN U326 ( .B(clk), .A(\g.we_clk [32448]));
Q_ASSIGN U327 ( .B(clk), .A(\g.we_clk [32447]));
Q_ASSIGN U328 ( .B(clk), .A(\g.we_clk [32446]));
Q_ASSIGN U329 ( .B(clk), .A(\g.we_clk [32445]));
Q_ASSIGN U330 ( .B(clk), .A(\g.we_clk [32444]));
Q_ASSIGN U331 ( .B(clk), .A(\g.we_clk [32443]));
Q_ASSIGN U332 ( .B(clk), .A(\g.we_clk [32442]));
Q_ASSIGN U333 ( .B(clk), .A(\g.we_clk [32441]));
Q_ASSIGN U334 ( .B(clk), .A(\g.we_clk [32440]));
Q_ASSIGN U335 ( .B(clk), .A(\g.we_clk [32439]));
Q_ASSIGN U336 ( .B(clk), .A(\g.we_clk [32438]));
Q_ASSIGN U337 ( .B(clk), .A(\g.we_clk [32437]));
Q_ASSIGN U338 ( .B(clk), .A(\g.we_clk [32436]));
Q_ASSIGN U339 ( .B(clk), .A(\g.we_clk [32435]));
Q_ASSIGN U340 ( .B(clk), .A(\g.we_clk [32434]));
Q_ASSIGN U341 ( .B(clk), .A(\g.we_clk [32433]));
Q_ASSIGN U342 ( .B(clk), .A(\g.we_clk [32432]));
Q_ASSIGN U343 ( .B(clk), .A(\g.we_clk [32431]));
Q_ASSIGN U344 ( .B(clk), .A(\g.we_clk [32430]));
Q_ASSIGN U345 ( .B(clk), .A(\g.we_clk [32429]));
Q_ASSIGN U346 ( .B(clk), .A(\g.we_clk [32428]));
Q_ASSIGN U347 ( .B(clk), .A(\g.we_clk [32427]));
Q_ASSIGN U348 ( .B(clk), .A(\g.we_clk [32426]));
Q_ASSIGN U349 ( .B(clk), .A(\g.we_clk [32425]));
Q_ASSIGN U350 ( .B(clk), .A(\g.we_clk [32424]));
Q_ASSIGN U351 ( .B(clk), .A(\g.we_clk [32423]));
Q_ASSIGN U352 ( .B(clk), .A(\g.we_clk [32422]));
Q_ASSIGN U353 ( .B(clk), .A(\g.we_clk [32421]));
Q_ASSIGN U354 ( .B(clk), .A(\g.we_clk [32420]));
Q_ASSIGN U355 ( .B(clk), .A(\g.we_clk [32419]));
Q_ASSIGN U356 ( .B(clk), .A(\g.we_clk [32418]));
Q_ASSIGN U357 ( .B(clk), .A(\g.we_clk [32417]));
Q_ASSIGN U358 ( .B(clk), .A(\g.we_clk [32416]));
Q_ASSIGN U359 ( .B(clk), .A(\g.we_clk [32415]));
Q_ASSIGN U360 ( .B(clk), .A(\g.we_clk [32414]));
Q_ASSIGN U361 ( .B(clk), .A(\g.we_clk [32413]));
Q_ASSIGN U362 ( .B(clk), .A(\g.we_clk [32412]));
Q_ASSIGN U363 ( .B(clk), .A(\g.we_clk [32411]));
Q_ASSIGN U364 ( .B(clk), .A(\g.we_clk [32410]));
Q_ASSIGN U365 ( .B(clk), .A(\g.we_clk [32409]));
Q_ASSIGN U366 ( .B(clk), .A(\g.we_clk [32408]));
Q_ASSIGN U367 ( .B(clk), .A(\g.we_clk [32407]));
Q_ASSIGN U368 ( .B(clk), .A(\g.we_clk [32406]));
Q_ASSIGN U369 ( .B(clk), .A(\g.we_clk [32405]));
Q_ASSIGN U370 ( .B(clk), .A(\g.we_clk [32404]));
Q_ASSIGN U371 ( .B(clk), .A(\g.we_clk [32403]));
Q_ASSIGN U372 ( .B(clk), .A(\g.we_clk [32402]));
Q_ASSIGN U373 ( .B(clk), .A(\g.we_clk [32401]));
Q_ASSIGN U374 ( .B(clk), .A(\g.we_clk [32400]));
Q_ASSIGN U375 ( .B(clk), .A(\g.we_clk [32399]));
Q_ASSIGN U376 ( .B(clk), .A(\g.we_clk [32398]));
Q_ASSIGN U377 ( .B(clk), .A(\g.we_clk [32397]));
Q_ASSIGN U378 ( .B(clk), .A(\g.we_clk [32396]));
Q_ASSIGN U379 ( .B(clk), .A(\g.we_clk [32395]));
Q_ASSIGN U380 ( .B(clk), .A(\g.we_clk [32394]));
Q_ASSIGN U381 ( .B(clk), .A(\g.we_clk [32393]));
Q_ASSIGN U382 ( .B(clk), .A(\g.we_clk [32392]));
Q_ASSIGN U383 ( .B(clk), .A(\g.we_clk [32391]));
Q_ASSIGN U384 ( .B(clk), .A(\g.we_clk [32390]));
Q_ASSIGN U385 ( .B(clk), .A(\g.we_clk [32389]));
Q_ASSIGN U386 ( .B(clk), .A(\g.we_clk [32388]));
Q_ASSIGN U387 ( .B(clk), .A(\g.we_clk [32387]));
Q_ASSIGN U388 ( .B(clk), .A(\g.we_clk [32386]));
Q_ASSIGN U389 ( .B(clk), .A(\g.we_clk [32385]));
Q_ASSIGN U390 ( .B(clk), .A(\g.we_clk [32384]));
Q_ASSIGN U391 ( .B(clk), .A(\g.we_clk [32383]));
Q_ASSIGN U392 ( .B(clk), .A(\g.we_clk [32382]));
Q_ASSIGN U393 ( .B(clk), .A(\g.we_clk [32381]));
Q_ASSIGN U394 ( .B(clk), .A(\g.we_clk [32380]));
Q_ASSIGN U395 ( .B(clk), .A(\g.we_clk [32379]));
Q_ASSIGN U396 ( .B(clk), .A(\g.we_clk [32378]));
Q_ASSIGN U397 ( .B(clk), .A(\g.we_clk [32377]));
Q_ASSIGN U398 ( .B(clk), .A(\g.we_clk [32376]));
Q_ASSIGN U399 ( .B(clk), .A(\g.we_clk [32375]));
Q_ASSIGN U400 ( .B(clk), .A(\g.we_clk [32374]));
Q_ASSIGN U401 ( .B(clk), .A(\g.we_clk [32373]));
Q_ASSIGN U402 ( .B(clk), .A(\g.we_clk [32372]));
Q_ASSIGN U403 ( .B(clk), .A(\g.we_clk [32371]));
Q_ASSIGN U404 ( .B(clk), .A(\g.we_clk [32370]));
Q_ASSIGN U405 ( .B(clk), .A(\g.we_clk [32369]));
Q_ASSIGN U406 ( .B(clk), .A(\g.we_clk [32368]));
Q_ASSIGN U407 ( .B(clk), .A(\g.we_clk [32367]));
Q_ASSIGN U408 ( .B(clk), .A(\g.we_clk [32366]));
Q_ASSIGN U409 ( .B(clk), .A(\g.we_clk [32365]));
Q_ASSIGN U410 ( .B(clk), .A(\g.we_clk [32364]));
Q_ASSIGN U411 ( .B(clk), .A(\g.we_clk [32363]));
Q_ASSIGN U412 ( .B(clk), .A(\g.we_clk [32362]));
Q_ASSIGN U413 ( .B(clk), .A(\g.we_clk [32361]));
Q_ASSIGN U414 ( .B(clk), .A(\g.we_clk [32360]));
Q_ASSIGN U415 ( .B(clk), .A(\g.we_clk [32359]));
Q_ASSIGN U416 ( .B(clk), .A(\g.we_clk [32358]));
Q_ASSIGN U417 ( .B(clk), .A(\g.we_clk [32357]));
Q_ASSIGN U418 ( .B(clk), .A(\g.we_clk [32356]));
Q_ASSIGN U419 ( .B(clk), .A(\g.we_clk [32355]));
Q_ASSIGN U420 ( .B(clk), .A(\g.we_clk [32354]));
Q_ASSIGN U421 ( .B(clk), .A(\g.we_clk [32353]));
Q_ASSIGN U422 ( .B(clk), .A(\g.we_clk [32352]));
Q_ASSIGN U423 ( .B(clk), .A(\g.we_clk [32351]));
Q_ASSIGN U424 ( .B(clk), .A(\g.we_clk [32350]));
Q_ASSIGN U425 ( .B(clk), .A(\g.we_clk [32349]));
Q_ASSIGN U426 ( .B(clk), .A(\g.we_clk [32348]));
Q_ASSIGN U427 ( .B(clk), .A(\g.we_clk [32347]));
Q_ASSIGN U428 ( .B(clk), .A(\g.we_clk [32346]));
Q_ASSIGN U429 ( .B(clk), .A(\g.we_clk [32345]));
Q_ASSIGN U430 ( .B(clk), .A(\g.we_clk [32344]));
Q_ASSIGN U431 ( .B(clk), .A(\g.we_clk [32343]));
Q_ASSIGN U432 ( .B(clk), .A(\g.we_clk [32342]));
Q_ASSIGN U433 ( .B(clk), .A(\g.we_clk [32341]));
Q_ASSIGN U434 ( .B(clk), .A(\g.we_clk [32340]));
Q_ASSIGN U435 ( .B(clk), .A(\g.we_clk [32339]));
Q_ASSIGN U436 ( .B(clk), .A(\g.we_clk [32338]));
Q_ASSIGN U437 ( .B(clk), .A(\g.we_clk [32337]));
Q_ASSIGN U438 ( .B(clk), .A(\g.we_clk [32336]));
Q_ASSIGN U439 ( .B(clk), .A(\g.we_clk [32335]));
Q_ASSIGN U440 ( .B(clk), .A(\g.we_clk [32334]));
Q_ASSIGN U441 ( .B(clk), .A(\g.we_clk [32333]));
Q_ASSIGN U442 ( .B(clk), .A(\g.we_clk [32332]));
Q_ASSIGN U443 ( .B(clk), .A(\g.we_clk [32331]));
Q_ASSIGN U444 ( .B(clk), .A(\g.we_clk [32330]));
Q_ASSIGN U445 ( .B(clk), .A(\g.we_clk [32329]));
Q_ASSIGN U446 ( .B(clk), .A(\g.we_clk [32328]));
Q_ASSIGN U447 ( .B(clk), .A(\g.we_clk [32327]));
Q_ASSIGN U448 ( .B(clk), .A(\g.we_clk [32326]));
Q_ASSIGN U449 ( .B(clk), .A(\g.we_clk [32325]));
Q_ASSIGN U450 ( .B(clk), .A(\g.we_clk [32324]));
Q_ASSIGN U451 ( .B(clk), .A(\g.we_clk [32323]));
Q_ASSIGN U452 ( .B(clk), .A(\g.we_clk [32322]));
Q_ASSIGN U453 ( .B(clk), .A(\g.we_clk [32321]));
Q_ASSIGN U454 ( .B(clk), .A(\g.we_clk [32320]));
Q_ASSIGN U455 ( .B(clk), .A(\g.we_clk [32319]));
Q_ASSIGN U456 ( .B(clk), .A(\g.we_clk [32318]));
Q_ASSIGN U457 ( .B(clk), .A(\g.we_clk [32317]));
Q_ASSIGN U458 ( .B(clk), .A(\g.we_clk [32316]));
Q_ASSIGN U459 ( .B(clk), .A(\g.we_clk [32315]));
Q_ASSIGN U460 ( .B(clk), .A(\g.we_clk [32314]));
Q_ASSIGN U461 ( .B(clk), .A(\g.we_clk [32313]));
Q_ASSIGN U462 ( .B(clk), .A(\g.we_clk [32312]));
Q_ASSIGN U463 ( .B(clk), .A(\g.we_clk [32311]));
Q_ASSIGN U464 ( .B(clk), .A(\g.we_clk [32310]));
Q_ASSIGN U465 ( .B(clk), .A(\g.we_clk [32309]));
Q_ASSIGN U466 ( .B(clk), .A(\g.we_clk [32308]));
Q_ASSIGN U467 ( .B(clk), .A(\g.we_clk [32307]));
Q_ASSIGN U468 ( .B(clk), .A(\g.we_clk [32306]));
Q_ASSIGN U469 ( .B(clk), .A(\g.we_clk [32305]));
Q_ASSIGN U470 ( .B(clk), .A(\g.we_clk [32304]));
Q_ASSIGN U471 ( .B(clk), .A(\g.we_clk [32303]));
Q_ASSIGN U472 ( .B(clk), .A(\g.we_clk [32302]));
Q_ASSIGN U473 ( .B(clk), .A(\g.we_clk [32301]));
Q_ASSIGN U474 ( .B(clk), .A(\g.we_clk [32300]));
Q_ASSIGN U475 ( .B(clk), .A(\g.we_clk [32299]));
Q_ASSIGN U476 ( .B(clk), .A(\g.we_clk [32298]));
Q_ASSIGN U477 ( .B(clk), .A(\g.we_clk [32297]));
Q_ASSIGN U478 ( .B(clk), .A(\g.we_clk [32296]));
Q_ASSIGN U479 ( .B(clk), .A(\g.we_clk [32295]));
Q_ASSIGN U480 ( .B(clk), .A(\g.we_clk [32294]));
Q_ASSIGN U481 ( .B(clk), .A(\g.we_clk [32293]));
Q_ASSIGN U482 ( .B(clk), .A(\g.we_clk [32292]));
Q_ASSIGN U483 ( .B(clk), .A(\g.we_clk [32291]));
Q_ASSIGN U484 ( .B(clk), .A(\g.we_clk [32290]));
Q_ASSIGN U485 ( .B(clk), .A(\g.we_clk [32289]));
Q_ASSIGN U486 ( .B(clk), .A(\g.we_clk [32288]));
Q_ASSIGN U487 ( .B(clk), .A(\g.we_clk [32287]));
Q_ASSIGN U488 ( .B(clk), .A(\g.we_clk [32286]));
Q_ASSIGN U489 ( .B(clk), .A(\g.we_clk [32285]));
Q_ASSIGN U490 ( .B(clk), .A(\g.we_clk [32284]));
Q_ASSIGN U491 ( .B(clk), .A(\g.we_clk [32283]));
Q_ASSIGN U492 ( .B(clk), .A(\g.we_clk [32282]));
Q_ASSIGN U493 ( .B(clk), .A(\g.we_clk [32281]));
Q_ASSIGN U494 ( .B(clk), .A(\g.we_clk [32280]));
Q_ASSIGN U495 ( .B(clk), .A(\g.we_clk [32279]));
Q_ASSIGN U496 ( .B(clk), .A(\g.we_clk [32278]));
Q_ASSIGN U497 ( .B(clk), .A(\g.we_clk [32277]));
Q_ASSIGN U498 ( .B(clk), .A(\g.we_clk [32276]));
Q_ASSIGN U499 ( .B(clk), .A(\g.we_clk [32275]));
Q_ASSIGN U500 ( .B(clk), .A(\g.we_clk [32274]));
Q_ASSIGN U501 ( .B(clk), .A(\g.we_clk [32273]));
Q_ASSIGN U502 ( .B(clk), .A(\g.we_clk [32272]));
Q_ASSIGN U503 ( .B(clk), .A(\g.we_clk [32271]));
Q_ASSIGN U504 ( .B(clk), .A(\g.we_clk [32270]));
Q_ASSIGN U505 ( .B(clk), .A(\g.we_clk [32269]));
Q_ASSIGN U506 ( .B(clk), .A(\g.we_clk [32268]));
Q_ASSIGN U507 ( .B(clk), .A(\g.we_clk [32267]));
Q_ASSIGN U508 ( .B(clk), .A(\g.we_clk [32266]));
Q_ASSIGN U509 ( .B(clk), .A(\g.we_clk [32265]));
Q_ASSIGN U510 ( .B(clk), .A(\g.we_clk [32264]));
Q_ASSIGN U511 ( .B(clk), .A(\g.we_clk [32263]));
Q_ASSIGN U512 ( .B(clk), .A(\g.we_clk [32262]));
Q_ASSIGN U513 ( .B(clk), .A(\g.we_clk [32261]));
Q_ASSIGN U514 ( .B(clk), .A(\g.we_clk [32260]));
Q_ASSIGN U515 ( .B(clk), .A(\g.we_clk [32259]));
Q_ASSIGN U516 ( .B(clk), .A(\g.we_clk [32258]));
Q_ASSIGN U517 ( .B(clk), .A(\g.we_clk [32257]));
Q_ASSIGN U518 ( .B(clk), .A(\g.we_clk [32256]));
Q_ASSIGN U519 ( .B(clk), .A(\g.we_clk [32255]));
Q_ASSIGN U520 ( .B(clk), .A(\g.we_clk [32254]));
Q_ASSIGN U521 ( .B(clk), .A(\g.we_clk [32253]));
Q_ASSIGN U522 ( .B(clk), .A(\g.we_clk [32252]));
Q_ASSIGN U523 ( .B(clk), .A(\g.we_clk [32251]));
Q_ASSIGN U524 ( .B(clk), .A(\g.we_clk [32250]));
Q_ASSIGN U525 ( .B(clk), .A(\g.we_clk [32249]));
Q_ASSIGN U526 ( .B(clk), .A(\g.we_clk [32248]));
Q_ASSIGN U527 ( .B(clk), .A(\g.we_clk [32247]));
Q_ASSIGN U528 ( .B(clk), .A(\g.we_clk [32246]));
Q_ASSIGN U529 ( .B(clk), .A(\g.we_clk [32245]));
Q_ASSIGN U530 ( .B(clk), .A(\g.we_clk [32244]));
Q_ASSIGN U531 ( .B(clk), .A(\g.we_clk [32243]));
Q_ASSIGN U532 ( .B(clk), .A(\g.we_clk [32242]));
Q_ASSIGN U533 ( .B(clk), .A(\g.we_clk [32241]));
Q_ASSIGN U534 ( .B(clk), .A(\g.we_clk [32240]));
Q_ASSIGN U535 ( .B(clk), .A(\g.we_clk [32239]));
Q_ASSIGN U536 ( .B(clk), .A(\g.we_clk [32238]));
Q_ASSIGN U537 ( .B(clk), .A(\g.we_clk [32237]));
Q_ASSIGN U538 ( .B(clk), .A(\g.we_clk [32236]));
Q_ASSIGN U539 ( .B(clk), .A(\g.we_clk [32235]));
Q_ASSIGN U540 ( .B(clk), .A(\g.we_clk [32234]));
Q_ASSIGN U541 ( .B(clk), .A(\g.we_clk [32233]));
Q_ASSIGN U542 ( .B(clk), .A(\g.we_clk [32232]));
Q_ASSIGN U543 ( .B(clk), .A(\g.we_clk [32231]));
Q_ASSIGN U544 ( .B(clk), .A(\g.we_clk [32230]));
Q_ASSIGN U545 ( .B(clk), .A(\g.we_clk [32229]));
Q_ASSIGN U546 ( .B(clk), .A(\g.we_clk [32228]));
Q_ASSIGN U547 ( .B(clk), .A(\g.we_clk [32227]));
Q_ASSIGN U548 ( .B(clk), .A(\g.we_clk [32226]));
Q_ASSIGN U549 ( .B(clk), .A(\g.we_clk [32225]));
Q_ASSIGN U550 ( .B(clk), .A(\g.we_clk [32224]));
Q_ASSIGN U551 ( .B(clk), .A(\g.we_clk [32223]));
Q_ASSIGN U552 ( .B(clk), .A(\g.we_clk [32222]));
Q_ASSIGN U553 ( .B(clk), .A(\g.we_clk [32221]));
Q_ASSIGN U554 ( .B(clk), .A(\g.we_clk [32220]));
Q_ASSIGN U555 ( .B(clk), .A(\g.we_clk [32219]));
Q_ASSIGN U556 ( .B(clk), .A(\g.we_clk [32218]));
Q_ASSIGN U557 ( .B(clk), .A(\g.we_clk [32217]));
Q_ASSIGN U558 ( .B(clk), .A(\g.we_clk [32216]));
Q_ASSIGN U559 ( .B(clk), .A(\g.we_clk [32215]));
Q_ASSIGN U560 ( .B(clk), .A(\g.we_clk [32214]));
Q_ASSIGN U561 ( .B(clk), .A(\g.we_clk [32213]));
Q_ASSIGN U562 ( .B(clk), .A(\g.we_clk [32212]));
Q_ASSIGN U563 ( .B(clk), .A(\g.we_clk [32211]));
Q_ASSIGN U564 ( .B(clk), .A(\g.we_clk [32210]));
Q_ASSIGN U565 ( .B(clk), .A(\g.we_clk [32209]));
Q_ASSIGN U566 ( .B(clk), .A(\g.we_clk [32208]));
Q_ASSIGN U567 ( .B(clk), .A(\g.we_clk [32207]));
Q_ASSIGN U568 ( .B(clk), .A(\g.we_clk [32206]));
Q_ASSIGN U569 ( .B(clk), .A(\g.we_clk [32205]));
Q_ASSIGN U570 ( .B(clk), .A(\g.we_clk [32204]));
Q_ASSIGN U571 ( .B(clk), .A(\g.we_clk [32203]));
Q_ASSIGN U572 ( .B(clk), .A(\g.we_clk [32202]));
Q_ASSIGN U573 ( .B(clk), .A(\g.we_clk [32201]));
Q_ASSIGN U574 ( .B(clk), .A(\g.we_clk [32200]));
Q_ASSIGN U575 ( .B(clk), .A(\g.we_clk [32199]));
Q_ASSIGN U576 ( .B(clk), .A(\g.we_clk [32198]));
Q_ASSIGN U577 ( .B(clk), .A(\g.we_clk [32197]));
Q_ASSIGN U578 ( .B(clk), .A(\g.we_clk [32196]));
Q_ASSIGN U579 ( .B(clk), .A(\g.we_clk [32195]));
Q_ASSIGN U580 ( .B(clk), .A(\g.we_clk [32194]));
Q_ASSIGN U581 ( .B(clk), .A(\g.we_clk [32193]));
Q_ASSIGN U582 ( .B(clk), .A(\g.we_clk [32192]));
Q_ASSIGN U583 ( .B(clk), .A(\g.we_clk [32191]));
Q_ASSIGN U584 ( .B(clk), .A(\g.we_clk [32190]));
Q_ASSIGN U585 ( .B(clk), .A(\g.we_clk [32189]));
Q_ASSIGN U586 ( .B(clk), .A(\g.we_clk [32188]));
Q_ASSIGN U587 ( .B(clk), .A(\g.we_clk [32187]));
Q_ASSIGN U588 ( .B(clk), .A(\g.we_clk [32186]));
Q_ASSIGN U589 ( .B(clk), .A(\g.we_clk [32185]));
Q_ASSIGN U590 ( .B(clk), .A(\g.we_clk [32184]));
Q_ASSIGN U591 ( .B(clk), .A(\g.we_clk [32183]));
Q_ASSIGN U592 ( .B(clk), .A(\g.we_clk [32182]));
Q_ASSIGN U593 ( .B(clk), .A(\g.we_clk [32181]));
Q_ASSIGN U594 ( .B(clk), .A(\g.we_clk [32180]));
Q_ASSIGN U595 ( .B(clk), .A(\g.we_clk [32179]));
Q_ASSIGN U596 ( .B(clk), .A(\g.we_clk [32178]));
Q_ASSIGN U597 ( .B(clk), .A(\g.we_clk [32177]));
Q_ASSIGN U598 ( .B(clk), .A(\g.we_clk [32176]));
Q_ASSIGN U599 ( .B(clk), .A(\g.we_clk [32175]));
Q_ASSIGN U600 ( .B(clk), .A(\g.we_clk [32174]));
Q_ASSIGN U601 ( .B(clk), .A(\g.we_clk [32173]));
Q_ASSIGN U602 ( .B(clk), .A(\g.we_clk [32172]));
Q_ASSIGN U603 ( .B(clk), .A(\g.we_clk [32171]));
Q_ASSIGN U604 ( .B(clk), .A(\g.we_clk [32170]));
Q_ASSIGN U605 ( .B(clk), .A(\g.we_clk [32169]));
Q_ASSIGN U606 ( .B(clk), .A(\g.we_clk [32168]));
Q_ASSIGN U607 ( .B(clk), .A(\g.we_clk [32167]));
Q_ASSIGN U608 ( .B(clk), .A(\g.we_clk [32166]));
Q_ASSIGN U609 ( .B(clk), .A(\g.we_clk [32165]));
Q_ASSIGN U610 ( .B(clk), .A(\g.we_clk [32164]));
Q_ASSIGN U611 ( .B(clk), .A(\g.we_clk [32163]));
Q_ASSIGN U612 ( .B(clk), .A(\g.we_clk [32162]));
Q_ASSIGN U613 ( .B(clk), .A(\g.we_clk [32161]));
Q_ASSIGN U614 ( .B(clk), .A(\g.we_clk [32160]));
Q_ASSIGN U615 ( .B(clk), .A(\g.we_clk [32159]));
Q_ASSIGN U616 ( .B(clk), .A(\g.we_clk [32158]));
Q_ASSIGN U617 ( .B(clk), .A(\g.we_clk [32157]));
Q_ASSIGN U618 ( .B(clk), .A(\g.we_clk [32156]));
Q_ASSIGN U619 ( .B(clk), .A(\g.we_clk [32155]));
Q_ASSIGN U620 ( .B(clk), .A(\g.we_clk [32154]));
Q_ASSIGN U621 ( .B(clk), .A(\g.we_clk [32153]));
Q_ASSIGN U622 ( .B(clk), .A(\g.we_clk [32152]));
Q_ASSIGN U623 ( .B(clk), .A(\g.we_clk [32151]));
Q_ASSIGN U624 ( .B(clk), .A(\g.we_clk [32150]));
Q_ASSIGN U625 ( .B(clk), .A(\g.we_clk [32149]));
Q_ASSIGN U626 ( .B(clk), .A(\g.we_clk [32148]));
Q_ASSIGN U627 ( .B(clk), .A(\g.we_clk [32147]));
Q_ASSIGN U628 ( .B(clk), .A(\g.we_clk [32146]));
Q_ASSIGN U629 ( .B(clk), .A(\g.we_clk [32145]));
Q_ASSIGN U630 ( .B(clk), .A(\g.we_clk [32144]));
Q_ASSIGN U631 ( .B(clk), .A(\g.we_clk [32143]));
Q_ASSIGN U632 ( .B(clk), .A(\g.we_clk [32142]));
Q_ASSIGN U633 ( .B(clk), .A(\g.we_clk [32141]));
Q_ASSIGN U634 ( .B(clk), .A(\g.we_clk [32140]));
Q_ASSIGN U635 ( .B(clk), .A(\g.we_clk [32139]));
Q_ASSIGN U636 ( .B(clk), .A(\g.we_clk [32138]));
Q_ASSIGN U637 ( .B(clk), .A(\g.we_clk [32137]));
Q_ASSIGN U638 ( .B(clk), .A(\g.we_clk [32136]));
Q_ASSIGN U639 ( .B(clk), .A(\g.we_clk [32135]));
Q_ASSIGN U640 ( .B(clk), .A(\g.we_clk [32134]));
Q_ASSIGN U641 ( .B(clk), .A(\g.we_clk [32133]));
Q_ASSIGN U642 ( .B(clk), .A(\g.we_clk [32132]));
Q_ASSIGN U643 ( .B(clk), .A(\g.we_clk [32131]));
Q_ASSIGN U644 ( .B(clk), .A(\g.we_clk [32130]));
Q_ASSIGN U645 ( .B(clk), .A(\g.we_clk [32129]));
Q_ASSIGN U646 ( .B(clk), .A(\g.we_clk [32128]));
Q_ASSIGN U647 ( .B(clk), .A(\g.we_clk [32127]));
Q_ASSIGN U648 ( .B(clk), .A(\g.we_clk [32126]));
Q_ASSIGN U649 ( .B(clk), .A(\g.we_clk [32125]));
Q_ASSIGN U650 ( .B(clk), .A(\g.we_clk [32124]));
Q_ASSIGN U651 ( .B(clk), .A(\g.we_clk [32123]));
Q_ASSIGN U652 ( .B(clk), .A(\g.we_clk [32122]));
Q_ASSIGN U653 ( .B(clk), .A(\g.we_clk [32121]));
Q_ASSIGN U654 ( .B(clk), .A(\g.we_clk [32120]));
Q_ASSIGN U655 ( .B(clk), .A(\g.we_clk [32119]));
Q_ASSIGN U656 ( .B(clk), .A(\g.we_clk [32118]));
Q_ASSIGN U657 ( .B(clk), .A(\g.we_clk [32117]));
Q_ASSIGN U658 ( .B(clk), .A(\g.we_clk [32116]));
Q_ASSIGN U659 ( .B(clk), .A(\g.we_clk [32115]));
Q_ASSIGN U660 ( .B(clk), .A(\g.we_clk [32114]));
Q_ASSIGN U661 ( .B(clk), .A(\g.we_clk [32113]));
Q_ASSIGN U662 ( .B(clk), .A(\g.we_clk [32112]));
Q_ASSIGN U663 ( .B(clk), .A(\g.we_clk [32111]));
Q_ASSIGN U664 ( .B(clk), .A(\g.we_clk [32110]));
Q_ASSIGN U665 ( .B(clk), .A(\g.we_clk [32109]));
Q_ASSIGN U666 ( .B(clk), .A(\g.we_clk [32108]));
Q_ASSIGN U667 ( .B(clk), .A(\g.we_clk [32107]));
Q_ASSIGN U668 ( .B(clk), .A(\g.we_clk [32106]));
Q_ASSIGN U669 ( .B(clk), .A(\g.we_clk [32105]));
Q_ASSIGN U670 ( .B(clk), .A(\g.we_clk [32104]));
Q_ASSIGN U671 ( .B(clk), .A(\g.we_clk [32103]));
Q_ASSIGN U672 ( .B(clk), .A(\g.we_clk [32102]));
Q_ASSIGN U673 ( .B(clk), .A(\g.we_clk [32101]));
Q_ASSIGN U674 ( .B(clk), .A(\g.we_clk [32100]));
Q_ASSIGN U675 ( .B(clk), .A(\g.we_clk [32099]));
Q_ASSIGN U676 ( .B(clk), .A(\g.we_clk [32098]));
Q_ASSIGN U677 ( .B(clk), .A(\g.we_clk [32097]));
Q_ASSIGN U678 ( .B(clk), .A(\g.we_clk [32096]));
Q_ASSIGN U679 ( .B(clk), .A(\g.we_clk [32095]));
Q_ASSIGN U680 ( .B(clk), .A(\g.we_clk [32094]));
Q_ASSIGN U681 ( .B(clk), .A(\g.we_clk [32093]));
Q_ASSIGN U682 ( .B(clk), .A(\g.we_clk [32092]));
Q_ASSIGN U683 ( .B(clk), .A(\g.we_clk [32091]));
Q_ASSIGN U684 ( .B(clk), .A(\g.we_clk [32090]));
Q_ASSIGN U685 ( .B(clk), .A(\g.we_clk [32089]));
Q_ASSIGN U686 ( .B(clk), .A(\g.we_clk [32088]));
Q_ASSIGN U687 ( .B(clk), .A(\g.we_clk [32087]));
Q_ASSIGN U688 ( .B(clk), .A(\g.we_clk [32086]));
Q_ASSIGN U689 ( .B(clk), .A(\g.we_clk [32085]));
Q_ASSIGN U690 ( .B(clk), .A(\g.we_clk [32084]));
Q_ASSIGN U691 ( .B(clk), .A(\g.we_clk [32083]));
Q_ASSIGN U692 ( .B(clk), .A(\g.we_clk [32082]));
Q_ASSIGN U693 ( .B(clk), .A(\g.we_clk [32081]));
Q_ASSIGN U694 ( .B(clk), .A(\g.we_clk [32080]));
Q_ASSIGN U695 ( .B(clk), .A(\g.we_clk [32079]));
Q_ASSIGN U696 ( .B(clk), .A(\g.we_clk [32078]));
Q_ASSIGN U697 ( .B(clk), .A(\g.we_clk [32077]));
Q_ASSIGN U698 ( .B(clk), .A(\g.we_clk [32076]));
Q_ASSIGN U699 ( .B(clk), .A(\g.we_clk [32075]));
Q_ASSIGN U700 ( .B(clk), .A(\g.we_clk [32074]));
Q_ASSIGN U701 ( .B(clk), .A(\g.we_clk [32073]));
Q_ASSIGN U702 ( .B(clk), .A(\g.we_clk [32072]));
Q_ASSIGN U703 ( .B(clk), .A(\g.we_clk [32071]));
Q_ASSIGN U704 ( .B(clk), .A(\g.we_clk [32070]));
Q_ASSIGN U705 ( .B(clk), .A(\g.we_clk [32069]));
Q_ASSIGN U706 ( .B(clk), .A(\g.we_clk [32068]));
Q_ASSIGN U707 ( .B(clk), .A(\g.we_clk [32067]));
Q_ASSIGN U708 ( .B(clk), .A(\g.we_clk [32066]));
Q_ASSIGN U709 ( .B(clk), .A(\g.we_clk [32065]));
Q_ASSIGN U710 ( .B(clk), .A(\g.we_clk [32064]));
Q_ASSIGN U711 ( .B(clk), .A(\g.we_clk [32063]));
Q_ASSIGN U712 ( .B(clk), .A(\g.we_clk [32062]));
Q_ASSIGN U713 ( .B(clk), .A(\g.we_clk [32061]));
Q_ASSIGN U714 ( .B(clk), .A(\g.we_clk [32060]));
Q_ASSIGN U715 ( .B(clk), .A(\g.we_clk [32059]));
Q_ASSIGN U716 ( .B(clk), .A(\g.we_clk [32058]));
Q_ASSIGN U717 ( .B(clk), .A(\g.we_clk [32057]));
Q_ASSIGN U718 ( .B(clk), .A(\g.we_clk [32056]));
Q_ASSIGN U719 ( .B(clk), .A(\g.we_clk [32055]));
Q_ASSIGN U720 ( .B(clk), .A(\g.we_clk [32054]));
Q_ASSIGN U721 ( .B(clk), .A(\g.we_clk [32053]));
Q_ASSIGN U722 ( .B(clk), .A(\g.we_clk [32052]));
Q_ASSIGN U723 ( .B(clk), .A(\g.we_clk [32051]));
Q_ASSIGN U724 ( .B(clk), .A(\g.we_clk [32050]));
Q_ASSIGN U725 ( .B(clk), .A(\g.we_clk [32049]));
Q_ASSIGN U726 ( .B(clk), .A(\g.we_clk [32048]));
Q_ASSIGN U727 ( .B(clk), .A(\g.we_clk [32047]));
Q_ASSIGN U728 ( .B(clk), .A(\g.we_clk [32046]));
Q_ASSIGN U729 ( .B(clk), .A(\g.we_clk [32045]));
Q_ASSIGN U730 ( .B(clk), .A(\g.we_clk [32044]));
Q_ASSIGN U731 ( .B(clk), .A(\g.we_clk [32043]));
Q_ASSIGN U732 ( .B(clk), .A(\g.we_clk [32042]));
Q_ASSIGN U733 ( .B(clk), .A(\g.we_clk [32041]));
Q_ASSIGN U734 ( .B(clk), .A(\g.we_clk [32040]));
Q_ASSIGN U735 ( .B(clk), .A(\g.we_clk [32039]));
Q_ASSIGN U736 ( .B(clk), .A(\g.we_clk [32038]));
Q_ASSIGN U737 ( .B(clk), .A(\g.we_clk [32037]));
Q_ASSIGN U738 ( .B(clk), .A(\g.we_clk [32036]));
Q_ASSIGN U739 ( .B(clk), .A(\g.we_clk [32035]));
Q_ASSIGN U740 ( .B(clk), .A(\g.we_clk [32034]));
Q_ASSIGN U741 ( .B(clk), .A(\g.we_clk [32033]));
Q_ASSIGN U742 ( .B(clk), .A(\g.we_clk [32032]));
Q_ASSIGN U743 ( .B(clk), .A(\g.we_clk [32031]));
Q_ASSIGN U744 ( .B(clk), .A(\g.we_clk [32030]));
Q_ASSIGN U745 ( .B(clk), .A(\g.we_clk [32029]));
Q_ASSIGN U746 ( .B(clk), .A(\g.we_clk [32028]));
Q_ASSIGN U747 ( .B(clk), .A(\g.we_clk [32027]));
Q_ASSIGN U748 ( .B(clk), .A(\g.we_clk [32026]));
Q_ASSIGN U749 ( .B(clk), .A(\g.we_clk [32025]));
Q_ASSIGN U750 ( .B(clk), .A(\g.we_clk [32024]));
Q_ASSIGN U751 ( .B(clk), .A(\g.we_clk [32023]));
Q_ASSIGN U752 ( .B(clk), .A(\g.we_clk [32022]));
Q_ASSIGN U753 ( .B(clk), .A(\g.we_clk [32021]));
Q_ASSIGN U754 ( .B(clk), .A(\g.we_clk [32020]));
Q_ASSIGN U755 ( .B(clk), .A(\g.we_clk [32019]));
Q_ASSIGN U756 ( .B(clk), .A(\g.we_clk [32018]));
Q_ASSIGN U757 ( .B(clk), .A(\g.we_clk [32017]));
Q_ASSIGN U758 ( .B(clk), .A(\g.we_clk [32016]));
Q_ASSIGN U759 ( .B(clk), .A(\g.we_clk [32015]));
Q_ASSIGN U760 ( .B(clk), .A(\g.we_clk [32014]));
Q_ASSIGN U761 ( .B(clk), .A(\g.we_clk [32013]));
Q_ASSIGN U762 ( .B(clk), .A(\g.we_clk [32012]));
Q_ASSIGN U763 ( .B(clk), .A(\g.we_clk [32011]));
Q_ASSIGN U764 ( .B(clk), .A(\g.we_clk [32010]));
Q_ASSIGN U765 ( .B(clk), .A(\g.we_clk [32009]));
Q_ASSIGN U766 ( .B(clk), .A(\g.we_clk [32008]));
Q_ASSIGN U767 ( .B(clk), .A(\g.we_clk [32007]));
Q_ASSIGN U768 ( .B(clk), .A(\g.we_clk [32006]));
Q_ASSIGN U769 ( .B(clk), .A(\g.we_clk [32005]));
Q_ASSIGN U770 ( .B(clk), .A(\g.we_clk [32004]));
Q_ASSIGN U771 ( .B(clk), .A(\g.we_clk [32003]));
Q_ASSIGN U772 ( .B(clk), .A(\g.we_clk [32002]));
Q_ASSIGN U773 ( .B(clk), .A(\g.we_clk [32001]));
Q_ASSIGN U774 ( .B(clk), .A(\g.we_clk [32000]));
Q_ASSIGN U775 ( .B(clk), .A(\g.we_clk [31999]));
Q_ASSIGN U776 ( .B(clk), .A(\g.we_clk [31998]));
Q_ASSIGN U777 ( .B(clk), .A(\g.we_clk [31997]));
Q_ASSIGN U778 ( .B(clk), .A(\g.we_clk [31996]));
Q_ASSIGN U779 ( .B(clk), .A(\g.we_clk [31995]));
Q_ASSIGN U780 ( .B(clk), .A(\g.we_clk [31994]));
Q_ASSIGN U781 ( .B(clk), .A(\g.we_clk [31993]));
Q_ASSIGN U782 ( .B(clk), .A(\g.we_clk [31992]));
Q_ASSIGN U783 ( .B(clk), .A(\g.we_clk [31991]));
Q_ASSIGN U784 ( .B(clk), .A(\g.we_clk [31990]));
Q_ASSIGN U785 ( .B(clk), .A(\g.we_clk [31989]));
Q_ASSIGN U786 ( .B(clk), .A(\g.we_clk [31988]));
Q_ASSIGN U787 ( .B(clk), .A(\g.we_clk [31987]));
Q_ASSIGN U788 ( .B(clk), .A(\g.we_clk [31986]));
Q_ASSIGN U789 ( .B(clk), .A(\g.we_clk [31985]));
Q_ASSIGN U790 ( .B(clk), .A(\g.we_clk [31984]));
Q_ASSIGN U791 ( .B(clk), .A(\g.we_clk [31983]));
Q_ASSIGN U792 ( .B(clk), .A(\g.we_clk [31982]));
Q_ASSIGN U793 ( .B(clk), .A(\g.we_clk [31981]));
Q_ASSIGN U794 ( .B(clk), .A(\g.we_clk [31980]));
Q_ASSIGN U795 ( .B(clk), .A(\g.we_clk [31979]));
Q_ASSIGN U796 ( .B(clk), .A(\g.we_clk [31978]));
Q_ASSIGN U797 ( .B(clk), .A(\g.we_clk [31977]));
Q_ASSIGN U798 ( .B(clk), .A(\g.we_clk [31976]));
Q_ASSIGN U799 ( .B(clk), .A(\g.we_clk [31975]));
Q_ASSIGN U800 ( .B(clk), .A(\g.we_clk [31974]));
Q_ASSIGN U801 ( .B(clk), .A(\g.we_clk [31973]));
Q_ASSIGN U802 ( .B(clk), .A(\g.we_clk [31972]));
Q_ASSIGN U803 ( .B(clk), .A(\g.we_clk [31971]));
Q_ASSIGN U804 ( .B(clk), .A(\g.we_clk [31970]));
Q_ASSIGN U805 ( .B(clk), .A(\g.we_clk [31969]));
Q_ASSIGN U806 ( .B(clk), .A(\g.we_clk [31968]));
Q_ASSIGN U807 ( .B(clk), .A(\g.we_clk [31967]));
Q_ASSIGN U808 ( .B(clk), .A(\g.we_clk [31966]));
Q_ASSIGN U809 ( .B(clk), .A(\g.we_clk [31965]));
Q_ASSIGN U810 ( .B(clk), .A(\g.we_clk [31964]));
Q_ASSIGN U811 ( .B(clk), .A(\g.we_clk [31963]));
Q_ASSIGN U812 ( .B(clk), .A(\g.we_clk [31962]));
Q_ASSIGN U813 ( .B(clk), .A(\g.we_clk [31961]));
Q_ASSIGN U814 ( .B(clk), .A(\g.we_clk [31960]));
Q_ASSIGN U815 ( .B(clk), .A(\g.we_clk [31959]));
Q_ASSIGN U816 ( .B(clk), .A(\g.we_clk [31958]));
Q_ASSIGN U817 ( .B(clk), .A(\g.we_clk [31957]));
Q_ASSIGN U818 ( .B(clk), .A(\g.we_clk [31956]));
Q_ASSIGN U819 ( .B(clk), .A(\g.we_clk [31955]));
Q_ASSIGN U820 ( .B(clk), .A(\g.we_clk [31954]));
Q_ASSIGN U821 ( .B(clk), .A(\g.we_clk [31953]));
Q_ASSIGN U822 ( .B(clk), .A(\g.we_clk [31952]));
Q_ASSIGN U823 ( .B(clk), .A(\g.we_clk [31951]));
Q_ASSIGN U824 ( .B(clk), .A(\g.we_clk [31950]));
Q_ASSIGN U825 ( .B(clk), .A(\g.we_clk [31949]));
Q_ASSIGN U826 ( .B(clk), .A(\g.we_clk [31948]));
Q_ASSIGN U827 ( .B(clk), .A(\g.we_clk [31947]));
Q_ASSIGN U828 ( .B(clk), .A(\g.we_clk [31946]));
Q_ASSIGN U829 ( .B(clk), .A(\g.we_clk [31945]));
Q_ASSIGN U830 ( .B(clk), .A(\g.we_clk [31944]));
Q_ASSIGN U831 ( .B(clk), .A(\g.we_clk [31943]));
Q_ASSIGN U832 ( .B(clk), .A(\g.we_clk [31942]));
Q_ASSIGN U833 ( .B(clk), .A(\g.we_clk [31941]));
Q_ASSIGN U834 ( .B(clk), .A(\g.we_clk [31940]));
Q_ASSIGN U835 ( .B(clk), .A(\g.we_clk [31939]));
Q_ASSIGN U836 ( .B(clk), .A(\g.we_clk [31938]));
Q_ASSIGN U837 ( .B(clk), .A(\g.we_clk [31937]));
Q_ASSIGN U838 ( .B(clk), .A(\g.we_clk [31936]));
Q_ASSIGN U839 ( .B(clk), .A(\g.we_clk [31935]));
Q_ASSIGN U840 ( .B(clk), .A(\g.we_clk [31934]));
Q_ASSIGN U841 ( .B(clk), .A(\g.we_clk [31933]));
Q_ASSIGN U842 ( .B(clk), .A(\g.we_clk [31932]));
Q_ASSIGN U843 ( .B(clk), .A(\g.we_clk [31931]));
Q_ASSIGN U844 ( .B(clk), .A(\g.we_clk [31930]));
Q_ASSIGN U845 ( .B(clk), .A(\g.we_clk [31929]));
Q_ASSIGN U846 ( .B(clk), .A(\g.we_clk [31928]));
Q_ASSIGN U847 ( .B(clk), .A(\g.we_clk [31927]));
Q_ASSIGN U848 ( .B(clk), .A(\g.we_clk [31926]));
Q_ASSIGN U849 ( .B(clk), .A(\g.we_clk [31925]));
Q_ASSIGN U850 ( .B(clk), .A(\g.we_clk [31924]));
Q_ASSIGN U851 ( .B(clk), .A(\g.we_clk [31923]));
Q_ASSIGN U852 ( .B(clk), .A(\g.we_clk [31922]));
Q_ASSIGN U853 ( .B(clk), .A(\g.we_clk [31921]));
Q_ASSIGN U854 ( .B(clk), .A(\g.we_clk [31920]));
Q_ASSIGN U855 ( .B(clk), .A(\g.we_clk [31919]));
Q_ASSIGN U856 ( .B(clk), .A(\g.we_clk [31918]));
Q_ASSIGN U857 ( .B(clk), .A(\g.we_clk [31917]));
Q_ASSIGN U858 ( .B(clk), .A(\g.we_clk [31916]));
Q_ASSIGN U859 ( .B(clk), .A(\g.we_clk [31915]));
Q_ASSIGN U860 ( .B(clk), .A(\g.we_clk [31914]));
Q_ASSIGN U861 ( .B(clk), .A(\g.we_clk [31913]));
Q_ASSIGN U862 ( .B(clk), .A(\g.we_clk [31912]));
Q_ASSIGN U863 ( .B(clk), .A(\g.we_clk [31911]));
Q_ASSIGN U864 ( .B(clk), .A(\g.we_clk [31910]));
Q_ASSIGN U865 ( .B(clk), .A(\g.we_clk [31909]));
Q_ASSIGN U866 ( .B(clk), .A(\g.we_clk [31908]));
Q_ASSIGN U867 ( .B(clk), .A(\g.we_clk [31907]));
Q_ASSIGN U868 ( .B(clk), .A(\g.we_clk [31906]));
Q_ASSIGN U869 ( .B(clk), .A(\g.we_clk [31905]));
Q_ASSIGN U870 ( .B(clk), .A(\g.we_clk [31904]));
Q_ASSIGN U871 ( .B(clk), .A(\g.we_clk [31903]));
Q_ASSIGN U872 ( .B(clk), .A(\g.we_clk [31902]));
Q_ASSIGN U873 ( .B(clk), .A(\g.we_clk [31901]));
Q_ASSIGN U874 ( .B(clk), .A(\g.we_clk [31900]));
Q_ASSIGN U875 ( .B(clk), .A(\g.we_clk [31899]));
Q_ASSIGN U876 ( .B(clk), .A(\g.we_clk [31898]));
Q_ASSIGN U877 ( .B(clk), .A(\g.we_clk [31897]));
Q_ASSIGN U878 ( .B(clk), .A(\g.we_clk [31896]));
Q_ASSIGN U879 ( .B(clk), .A(\g.we_clk [31895]));
Q_ASSIGN U880 ( .B(clk), .A(\g.we_clk [31894]));
Q_ASSIGN U881 ( .B(clk), .A(\g.we_clk [31893]));
Q_ASSIGN U882 ( .B(clk), .A(\g.we_clk [31892]));
Q_ASSIGN U883 ( .B(clk), .A(\g.we_clk [31891]));
Q_ASSIGN U884 ( .B(clk), .A(\g.we_clk [31890]));
Q_ASSIGN U885 ( .B(clk), .A(\g.we_clk [31889]));
Q_ASSIGN U886 ( .B(clk), .A(\g.we_clk [31888]));
Q_ASSIGN U887 ( .B(clk), .A(\g.we_clk [31887]));
Q_ASSIGN U888 ( .B(clk), .A(\g.we_clk [31886]));
Q_ASSIGN U889 ( .B(clk), .A(\g.we_clk [31885]));
Q_ASSIGN U890 ( .B(clk), .A(\g.we_clk [31884]));
Q_ASSIGN U891 ( .B(clk), .A(\g.we_clk [31883]));
Q_ASSIGN U892 ( .B(clk), .A(\g.we_clk [31882]));
Q_ASSIGN U893 ( .B(clk), .A(\g.we_clk [31881]));
Q_ASSIGN U894 ( .B(clk), .A(\g.we_clk [31880]));
Q_ASSIGN U895 ( .B(clk), .A(\g.we_clk [31879]));
Q_ASSIGN U896 ( .B(clk), .A(\g.we_clk [31878]));
Q_ASSIGN U897 ( .B(clk), .A(\g.we_clk [31877]));
Q_ASSIGN U898 ( .B(clk), .A(\g.we_clk [31876]));
Q_ASSIGN U899 ( .B(clk), .A(\g.we_clk [31875]));
Q_ASSIGN U900 ( .B(clk), .A(\g.we_clk [31874]));
Q_ASSIGN U901 ( .B(clk), .A(\g.we_clk [31873]));
Q_ASSIGN U902 ( .B(clk), .A(\g.we_clk [31872]));
Q_ASSIGN U903 ( .B(clk), .A(\g.we_clk [31871]));
Q_ASSIGN U904 ( .B(clk), .A(\g.we_clk [31870]));
Q_ASSIGN U905 ( .B(clk), .A(\g.we_clk [31869]));
Q_ASSIGN U906 ( .B(clk), .A(\g.we_clk [31868]));
Q_ASSIGN U907 ( .B(clk), .A(\g.we_clk [31867]));
Q_ASSIGN U908 ( .B(clk), .A(\g.we_clk [31866]));
Q_ASSIGN U909 ( .B(clk), .A(\g.we_clk [31865]));
Q_ASSIGN U910 ( .B(clk), .A(\g.we_clk [31864]));
Q_ASSIGN U911 ( .B(clk), .A(\g.we_clk [31863]));
Q_ASSIGN U912 ( .B(clk), .A(\g.we_clk [31862]));
Q_ASSIGN U913 ( .B(clk), .A(\g.we_clk [31861]));
Q_ASSIGN U914 ( .B(clk), .A(\g.we_clk [31860]));
Q_ASSIGN U915 ( .B(clk), .A(\g.we_clk [31859]));
Q_ASSIGN U916 ( .B(clk), .A(\g.we_clk [31858]));
Q_ASSIGN U917 ( .B(clk), .A(\g.we_clk [31857]));
Q_ASSIGN U918 ( .B(clk), .A(\g.we_clk [31856]));
Q_ASSIGN U919 ( .B(clk), .A(\g.we_clk [31855]));
Q_ASSIGN U920 ( .B(clk), .A(\g.we_clk [31854]));
Q_ASSIGN U921 ( .B(clk), .A(\g.we_clk [31853]));
Q_ASSIGN U922 ( .B(clk), .A(\g.we_clk [31852]));
Q_ASSIGN U923 ( .B(clk), .A(\g.we_clk [31851]));
Q_ASSIGN U924 ( .B(clk), .A(\g.we_clk [31850]));
Q_ASSIGN U925 ( .B(clk), .A(\g.we_clk [31849]));
Q_ASSIGN U926 ( .B(clk), .A(\g.we_clk [31848]));
Q_ASSIGN U927 ( .B(clk), .A(\g.we_clk [31847]));
Q_ASSIGN U928 ( .B(clk), .A(\g.we_clk [31846]));
Q_ASSIGN U929 ( .B(clk), .A(\g.we_clk [31845]));
Q_ASSIGN U930 ( .B(clk), .A(\g.we_clk [31844]));
Q_ASSIGN U931 ( .B(clk), .A(\g.we_clk [31843]));
Q_ASSIGN U932 ( .B(clk), .A(\g.we_clk [31842]));
Q_ASSIGN U933 ( .B(clk), .A(\g.we_clk [31841]));
Q_ASSIGN U934 ( .B(clk), .A(\g.we_clk [31840]));
Q_ASSIGN U935 ( .B(clk), .A(\g.we_clk [31839]));
Q_ASSIGN U936 ( .B(clk), .A(\g.we_clk [31838]));
Q_ASSIGN U937 ( .B(clk), .A(\g.we_clk [31837]));
Q_ASSIGN U938 ( .B(clk), .A(\g.we_clk [31836]));
Q_ASSIGN U939 ( .B(clk), .A(\g.we_clk [31835]));
Q_ASSIGN U940 ( .B(clk), .A(\g.we_clk [31834]));
Q_ASSIGN U941 ( .B(clk), .A(\g.we_clk [31833]));
Q_ASSIGN U942 ( .B(clk), .A(\g.we_clk [31832]));
Q_ASSIGN U943 ( .B(clk), .A(\g.we_clk [31831]));
Q_ASSIGN U944 ( .B(clk), .A(\g.we_clk [31830]));
Q_ASSIGN U945 ( .B(clk), .A(\g.we_clk [31829]));
Q_ASSIGN U946 ( .B(clk), .A(\g.we_clk [31828]));
Q_ASSIGN U947 ( .B(clk), .A(\g.we_clk [31827]));
Q_ASSIGN U948 ( .B(clk), .A(\g.we_clk [31826]));
Q_ASSIGN U949 ( .B(clk), .A(\g.we_clk [31825]));
Q_ASSIGN U950 ( .B(clk), .A(\g.we_clk [31824]));
Q_ASSIGN U951 ( .B(clk), .A(\g.we_clk [31823]));
Q_ASSIGN U952 ( .B(clk), .A(\g.we_clk [31822]));
Q_ASSIGN U953 ( .B(clk), .A(\g.we_clk [31821]));
Q_ASSIGN U954 ( .B(clk), .A(\g.we_clk [31820]));
Q_ASSIGN U955 ( .B(clk), .A(\g.we_clk [31819]));
Q_ASSIGN U956 ( .B(clk), .A(\g.we_clk [31818]));
Q_ASSIGN U957 ( .B(clk), .A(\g.we_clk [31817]));
Q_ASSIGN U958 ( .B(clk), .A(\g.we_clk [31816]));
Q_ASSIGN U959 ( .B(clk), .A(\g.we_clk [31815]));
Q_ASSIGN U960 ( .B(clk), .A(\g.we_clk [31814]));
Q_ASSIGN U961 ( .B(clk), .A(\g.we_clk [31813]));
Q_ASSIGN U962 ( .B(clk), .A(\g.we_clk [31812]));
Q_ASSIGN U963 ( .B(clk), .A(\g.we_clk [31811]));
Q_ASSIGN U964 ( .B(clk), .A(\g.we_clk [31810]));
Q_ASSIGN U965 ( .B(clk), .A(\g.we_clk [31809]));
Q_ASSIGN U966 ( .B(clk), .A(\g.we_clk [31808]));
Q_ASSIGN U967 ( .B(clk), .A(\g.we_clk [31807]));
Q_ASSIGN U968 ( .B(clk), .A(\g.we_clk [31806]));
Q_ASSIGN U969 ( .B(clk), .A(\g.we_clk [31805]));
Q_ASSIGN U970 ( .B(clk), .A(\g.we_clk [31804]));
Q_ASSIGN U971 ( .B(clk), .A(\g.we_clk [31803]));
Q_ASSIGN U972 ( .B(clk), .A(\g.we_clk [31802]));
Q_ASSIGN U973 ( .B(clk), .A(\g.we_clk [31801]));
Q_ASSIGN U974 ( .B(clk), .A(\g.we_clk [31800]));
Q_ASSIGN U975 ( .B(clk), .A(\g.we_clk [31799]));
Q_ASSIGN U976 ( .B(clk), .A(\g.we_clk [31798]));
Q_ASSIGN U977 ( .B(clk), .A(\g.we_clk [31797]));
Q_ASSIGN U978 ( .B(clk), .A(\g.we_clk [31796]));
Q_ASSIGN U979 ( .B(clk), .A(\g.we_clk [31795]));
Q_ASSIGN U980 ( .B(clk), .A(\g.we_clk [31794]));
Q_ASSIGN U981 ( .B(clk), .A(\g.we_clk [31793]));
Q_ASSIGN U982 ( .B(clk), .A(\g.we_clk [31792]));
Q_ASSIGN U983 ( .B(clk), .A(\g.we_clk [31791]));
Q_ASSIGN U984 ( .B(clk), .A(\g.we_clk [31790]));
Q_ASSIGN U985 ( .B(clk), .A(\g.we_clk [31789]));
Q_ASSIGN U986 ( .B(clk), .A(\g.we_clk [31788]));
Q_ASSIGN U987 ( .B(clk), .A(\g.we_clk [31787]));
Q_ASSIGN U988 ( .B(clk), .A(\g.we_clk [31786]));
Q_ASSIGN U989 ( .B(clk), .A(\g.we_clk [31785]));
Q_ASSIGN U990 ( .B(clk), .A(\g.we_clk [31784]));
Q_ASSIGN U991 ( .B(clk), .A(\g.we_clk [31783]));
Q_ASSIGN U992 ( .B(clk), .A(\g.we_clk [31782]));
Q_ASSIGN U993 ( .B(clk), .A(\g.we_clk [31781]));
Q_ASSIGN U994 ( .B(clk), .A(\g.we_clk [31780]));
Q_ASSIGN U995 ( .B(clk), .A(\g.we_clk [31779]));
Q_ASSIGN U996 ( .B(clk), .A(\g.we_clk [31778]));
Q_ASSIGN U997 ( .B(clk), .A(\g.we_clk [31777]));
Q_ASSIGN U998 ( .B(clk), .A(\g.we_clk [31776]));
Q_ASSIGN U999 ( .B(clk), .A(\g.we_clk [31775]));
Q_ASSIGN U1000 ( .B(clk), .A(\g.we_clk [31774]));
Q_ASSIGN U1001 ( .B(clk), .A(\g.we_clk [31773]));
Q_ASSIGN U1002 ( .B(clk), .A(\g.we_clk [31772]));
Q_ASSIGN U1003 ( .B(clk), .A(\g.we_clk [31771]));
Q_ASSIGN U1004 ( .B(clk), .A(\g.we_clk [31770]));
Q_ASSIGN U1005 ( .B(clk), .A(\g.we_clk [31769]));
Q_ASSIGN U1006 ( .B(clk), .A(\g.we_clk [31768]));
Q_ASSIGN U1007 ( .B(clk), .A(\g.we_clk [31767]));
Q_ASSIGN U1008 ( .B(clk), .A(\g.we_clk [31766]));
Q_ASSIGN U1009 ( .B(clk), .A(\g.we_clk [31765]));
Q_ASSIGN U1010 ( .B(clk), .A(\g.we_clk [31764]));
Q_ASSIGN U1011 ( .B(clk), .A(\g.we_clk [31763]));
Q_ASSIGN U1012 ( .B(clk), .A(\g.we_clk [31762]));
Q_ASSIGN U1013 ( .B(clk), .A(\g.we_clk [31761]));
Q_ASSIGN U1014 ( .B(clk), .A(\g.we_clk [31760]));
Q_ASSIGN U1015 ( .B(clk), .A(\g.we_clk [31759]));
Q_ASSIGN U1016 ( .B(clk), .A(\g.we_clk [31758]));
Q_ASSIGN U1017 ( .B(clk), .A(\g.we_clk [31757]));
Q_ASSIGN U1018 ( .B(clk), .A(\g.we_clk [31756]));
Q_ASSIGN U1019 ( .B(clk), .A(\g.we_clk [31755]));
Q_ASSIGN U1020 ( .B(clk), .A(\g.we_clk [31754]));
Q_ASSIGN U1021 ( .B(clk), .A(\g.we_clk [31753]));
Q_ASSIGN U1022 ( .B(clk), .A(\g.we_clk [31752]));
Q_ASSIGN U1023 ( .B(clk), .A(\g.we_clk [31751]));
Q_ASSIGN U1024 ( .B(clk), .A(\g.we_clk [31750]));
Q_ASSIGN U1025 ( .B(clk), .A(\g.we_clk [31749]));
Q_ASSIGN U1026 ( .B(clk), .A(\g.we_clk [31748]));
Q_ASSIGN U1027 ( .B(clk), .A(\g.we_clk [31747]));
Q_ASSIGN U1028 ( .B(clk), .A(\g.we_clk [31746]));
Q_ASSIGN U1029 ( .B(clk), .A(\g.we_clk [31745]));
Q_ASSIGN U1030 ( .B(clk), .A(\g.we_clk [31744]));
Q_ASSIGN U1031 ( .B(clk), .A(\g.we_clk [31743]));
Q_ASSIGN U1032 ( .B(clk), .A(\g.we_clk [31742]));
Q_ASSIGN U1033 ( .B(clk), .A(\g.we_clk [31741]));
Q_ASSIGN U1034 ( .B(clk), .A(\g.we_clk [31740]));
Q_ASSIGN U1035 ( .B(clk), .A(\g.we_clk [31739]));
Q_ASSIGN U1036 ( .B(clk), .A(\g.we_clk [31738]));
Q_ASSIGN U1037 ( .B(clk), .A(\g.we_clk [31737]));
Q_ASSIGN U1038 ( .B(clk), .A(\g.we_clk [31736]));
Q_ASSIGN U1039 ( .B(clk), .A(\g.we_clk [31735]));
Q_ASSIGN U1040 ( .B(clk), .A(\g.we_clk [31734]));
Q_ASSIGN U1041 ( .B(clk), .A(\g.we_clk [31733]));
Q_ASSIGN U1042 ( .B(clk), .A(\g.we_clk [31732]));
Q_ASSIGN U1043 ( .B(clk), .A(\g.we_clk [31731]));
Q_ASSIGN U1044 ( .B(clk), .A(\g.we_clk [31730]));
Q_ASSIGN U1045 ( .B(clk), .A(\g.we_clk [31729]));
Q_ASSIGN U1046 ( .B(clk), .A(\g.we_clk [31728]));
Q_ASSIGN U1047 ( .B(clk), .A(\g.we_clk [31727]));
Q_ASSIGN U1048 ( .B(clk), .A(\g.we_clk [31726]));
Q_ASSIGN U1049 ( .B(clk), .A(\g.we_clk [31725]));
Q_ASSIGN U1050 ( .B(clk), .A(\g.we_clk [31724]));
Q_ASSIGN U1051 ( .B(clk), .A(\g.we_clk [31723]));
Q_ASSIGN U1052 ( .B(clk), .A(\g.we_clk [31722]));
Q_ASSIGN U1053 ( .B(clk), .A(\g.we_clk [31721]));
Q_ASSIGN U1054 ( .B(clk), .A(\g.we_clk [31720]));
Q_ASSIGN U1055 ( .B(clk), .A(\g.we_clk [31719]));
Q_ASSIGN U1056 ( .B(clk), .A(\g.we_clk [31718]));
Q_ASSIGN U1057 ( .B(clk), .A(\g.we_clk [31717]));
Q_ASSIGN U1058 ( .B(clk), .A(\g.we_clk [31716]));
Q_ASSIGN U1059 ( .B(clk), .A(\g.we_clk [31715]));
Q_ASSIGN U1060 ( .B(clk), .A(\g.we_clk [31714]));
Q_ASSIGN U1061 ( .B(clk), .A(\g.we_clk [31713]));
Q_ASSIGN U1062 ( .B(clk), .A(\g.we_clk [31712]));
Q_ASSIGN U1063 ( .B(clk), .A(\g.we_clk [31711]));
Q_ASSIGN U1064 ( .B(clk), .A(\g.we_clk [31710]));
Q_ASSIGN U1065 ( .B(clk), .A(\g.we_clk [31709]));
Q_ASSIGN U1066 ( .B(clk), .A(\g.we_clk [31708]));
Q_ASSIGN U1067 ( .B(clk), .A(\g.we_clk [31707]));
Q_ASSIGN U1068 ( .B(clk), .A(\g.we_clk [31706]));
Q_ASSIGN U1069 ( .B(clk), .A(\g.we_clk [31705]));
Q_ASSIGN U1070 ( .B(clk), .A(\g.we_clk [31704]));
Q_ASSIGN U1071 ( .B(clk), .A(\g.we_clk [31703]));
Q_ASSIGN U1072 ( .B(clk), .A(\g.we_clk [31702]));
Q_ASSIGN U1073 ( .B(clk), .A(\g.we_clk [31701]));
Q_ASSIGN U1074 ( .B(clk), .A(\g.we_clk [31700]));
Q_ASSIGN U1075 ( .B(clk), .A(\g.we_clk [31699]));
Q_ASSIGN U1076 ( .B(clk), .A(\g.we_clk [31698]));
Q_ASSIGN U1077 ( .B(clk), .A(\g.we_clk [31697]));
Q_ASSIGN U1078 ( .B(clk), .A(\g.we_clk [31696]));
Q_ASSIGN U1079 ( .B(clk), .A(\g.we_clk [31695]));
Q_ASSIGN U1080 ( .B(clk), .A(\g.we_clk [31694]));
Q_ASSIGN U1081 ( .B(clk), .A(\g.we_clk [31693]));
Q_ASSIGN U1082 ( .B(clk), .A(\g.we_clk [31692]));
Q_ASSIGN U1083 ( .B(clk), .A(\g.we_clk [31691]));
Q_ASSIGN U1084 ( .B(clk), .A(\g.we_clk [31690]));
Q_ASSIGN U1085 ( .B(clk), .A(\g.we_clk [31689]));
Q_ASSIGN U1086 ( .B(clk), .A(\g.we_clk [31688]));
Q_ASSIGN U1087 ( .B(clk), .A(\g.we_clk [31687]));
Q_ASSIGN U1088 ( .B(clk), .A(\g.we_clk [31686]));
Q_ASSIGN U1089 ( .B(clk), .A(\g.we_clk [31685]));
Q_ASSIGN U1090 ( .B(clk), .A(\g.we_clk [31684]));
Q_ASSIGN U1091 ( .B(clk), .A(\g.we_clk [31683]));
Q_ASSIGN U1092 ( .B(clk), .A(\g.we_clk [31682]));
Q_ASSIGN U1093 ( .B(clk), .A(\g.we_clk [31681]));
Q_ASSIGN U1094 ( .B(clk), .A(\g.we_clk [31680]));
Q_ASSIGN U1095 ( .B(clk), .A(\g.we_clk [31679]));
Q_ASSIGN U1096 ( .B(clk), .A(\g.we_clk [31678]));
Q_ASSIGN U1097 ( .B(clk), .A(\g.we_clk [31677]));
Q_ASSIGN U1098 ( .B(clk), .A(\g.we_clk [31676]));
Q_ASSIGN U1099 ( .B(clk), .A(\g.we_clk [31675]));
Q_ASSIGN U1100 ( .B(clk), .A(\g.we_clk [31674]));
Q_ASSIGN U1101 ( .B(clk), .A(\g.we_clk [31673]));
Q_ASSIGN U1102 ( .B(clk), .A(\g.we_clk [31672]));
Q_ASSIGN U1103 ( .B(clk), .A(\g.we_clk [31671]));
Q_ASSIGN U1104 ( .B(clk), .A(\g.we_clk [31670]));
Q_ASSIGN U1105 ( .B(clk), .A(\g.we_clk [31669]));
Q_ASSIGN U1106 ( .B(clk), .A(\g.we_clk [31668]));
Q_ASSIGN U1107 ( .B(clk), .A(\g.we_clk [31667]));
Q_ASSIGN U1108 ( .B(clk), .A(\g.we_clk [31666]));
Q_ASSIGN U1109 ( .B(clk), .A(\g.we_clk [31665]));
Q_ASSIGN U1110 ( .B(clk), .A(\g.we_clk [31664]));
Q_ASSIGN U1111 ( .B(clk), .A(\g.we_clk [31663]));
Q_ASSIGN U1112 ( .B(clk), .A(\g.we_clk [31662]));
Q_ASSIGN U1113 ( .B(clk), .A(\g.we_clk [31661]));
Q_ASSIGN U1114 ( .B(clk), .A(\g.we_clk [31660]));
Q_ASSIGN U1115 ( .B(clk), .A(\g.we_clk [31659]));
Q_ASSIGN U1116 ( .B(clk), .A(\g.we_clk [31658]));
Q_ASSIGN U1117 ( .B(clk), .A(\g.we_clk [31657]));
Q_ASSIGN U1118 ( .B(clk), .A(\g.we_clk [31656]));
Q_ASSIGN U1119 ( .B(clk), .A(\g.we_clk [31655]));
Q_ASSIGN U1120 ( .B(clk), .A(\g.we_clk [31654]));
Q_ASSIGN U1121 ( .B(clk), .A(\g.we_clk [31653]));
Q_ASSIGN U1122 ( .B(clk), .A(\g.we_clk [31652]));
Q_ASSIGN U1123 ( .B(clk), .A(\g.we_clk [31651]));
Q_ASSIGN U1124 ( .B(clk), .A(\g.we_clk [31650]));
Q_ASSIGN U1125 ( .B(clk), .A(\g.we_clk [31649]));
Q_ASSIGN U1126 ( .B(clk), .A(\g.we_clk [31648]));
Q_ASSIGN U1127 ( .B(clk), .A(\g.we_clk [31647]));
Q_ASSIGN U1128 ( .B(clk), .A(\g.we_clk [31646]));
Q_ASSIGN U1129 ( .B(clk), .A(\g.we_clk [31645]));
Q_ASSIGN U1130 ( .B(clk), .A(\g.we_clk [31644]));
Q_ASSIGN U1131 ( .B(clk), .A(\g.we_clk [31643]));
Q_ASSIGN U1132 ( .B(clk), .A(\g.we_clk [31642]));
Q_ASSIGN U1133 ( .B(clk), .A(\g.we_clk [31641]));
Q_ASSIGN U1134 ( .B(clk), .A(\g.we_clk [31640]));
Q_ASSIGN U1135 ( .B(clk), .A(\g.we_clk [31639]));
Q_ASSIGN U1136 ( .B(clk), .A(\g.we_clk [31638]));
Q_ASSIGN U1137 ( .B(clk), .A(\g.we_clk [31637]));
Q_ASSIGN U1138 ( .B(clk), .A(\g.we_clk [31636]));
Q_ASSIGN U1139 ( .B(clk), .A(\g.we_clk [31635]));
Q_ASSIGN U1140 ( .B(clk), .A(\g.we_clk [31634]));
Q_ASSIGN U1141 ( .B(clk), .A(\g.we_clk [31633]));
Q_ASSIGN U1142 ( .B(clk), .A(\g.we_clk [31632]));
Q_ASSIGN U1143 ( .B(clk), .A(\g.we_clk [31631]));
Q_ASSIGN U1144 ( .B(clk), .A(\g.we_clk [31630]));
Q_ASSIGN U1145 ( .B(clk), .A(\g.we_clk [31629]));
Q_ASSIGN U1146 ( .B(clk), .A(\g.we_clk [31628]));
Q_ASSIGN U1147 ( .B(clk), .A(\g.we_clk [31627]));
Q_ASSIGN U1148 ( .B(clk), .A(\g.we_clk [31626]));
Q_ASSIGN U1149 ( .B(clk), .A(\g.we_clk [31625]));
Q_ASSIGN U1150 ( .B(clk), .A(\g.we_clk [31624]));
Q_ASSIGN U1151 ( .B(clk), .A(\g.we_clk [31623]));
Q_ASSIGN U1152 ( .B(clk), .A(\g.we_clk [31622]));
Q_ASSIGN U1153 ( .B(clk), .A(\g.we_clk [31621]));
Q_ASSIGN U1154 ( .B(clk), .A(\g.we_clk [31620]));
Q_ASSIGN U1155 ( .B(clk), .A(\g.we_clk [31619]));
Q_ASSIGN U1156 ( .B(clk), .A(\g.we_clk [31618]));
Q_ASSIGN U1157 ( .B(clk), .A(\g.we_clk [31617]));
Q_ASSIGN U1158 ( .B(clk), .A(\g.we_clk [31616]));
Q_ASSIGN U1159 ( .B(clk), .A(\g.we_clk [31615]));
Q_ASSIGN U1160 ( .B(clk), .A(\g.we_clk [31614]));
Q_ASSIGN U1161 ( .B(clk), .A(\g.we_clk [31613]));
Q_ASSIGN U1162 ( .B(clk), .A(\g.we_clk [31612]));
Q_ASSIGN U1163 ( .B(clk), .A(\g.we_clk [31611]));
Q_ASSIGN U1164 ( .B(clk), .A(\g.we_clk [31610]));
Q_ASSIGN U1165 ( .B(clk), .A(\g.we_clk [31609]));
Q_ASSIGN U1166 ( .B(clk), .A(\g.we_clk [31608]));
Q_ASSIGN U1167 ( .B(clk), .A(\g.we_clk [31607]));
Q_ASSIGN U1168 ( .B(clk), .A(\g.we_clk [31606]));
Q_ASSIGN U1169 ( .B(clk), .A(\g.we_clk [31605]));
Q_ASSIGN U1170 ( .B(clk), .A(\g.we_clk [31604]));
Q_ASSIGN U1171 ( .B(clk), .A(\g.we_clk [31603]));
Q_ASSIGN U1172 ( .B(clk), .A(\g.we_clk [31602]));
Q_ASSIGN U1173 ( .B(clk), .A(\g.we_clk [31601]));
Q_ASSIGN U1174 ( .B(clk), .A(\g.we_clk [31600]));
Q_ASSIGN U1175 ( .B(clk), .A(\g.we_clk [31599]));
Q_ASSIGN U1176 ( .B(clk), .A(\g.we_clk [31598]));
Q_ASSIGN U1177 ( .B(clk), .A(\g.we_clk [31597]));
Q_ASSIGN U1178 ( .B(clk), .A(\g.we_clk [31596]));
Q_ASSIGN U1179 ( .B(clk), .A(\g.we_clk [31595]));
Q_ASSIGN U1180 ( .B(clk), .A(\g.we_clk [31594]));
Q_ASSIGN U1181 ( .B(clk), .A(\g.we_clk [31593]));
Q_ASSIGN U1182 ( .B(clk), .A(\g.we_clk [31592]));
Q_ASSIGN U1183 ( .B(clk), .A(\g.we_clk [31591]));
Q_ASSIGN U1184 ( .B(clk), .A(\g.we_clk [31590]));
Q_ASSIGN U1185 ( .B(clk), .A(\g.we_clk [31589]));
Q_ASSIGN U1186 ( .B(clk), .A(\g.we_clk [31588]));
Q_ASSIGN U1187 ( .B(clk), .A(\g.we_clk [31587]));
Q_ASSIGN U1188 ( .B(clk), .A(\g.we_clk [31586]));
Q_ASSIGN U1189 ( .B(clk), .A(\g.we_clk [31585]));
Q_ASSIGN U1190 ( .B(clk), .A(\g.we_clk [31584]));
Q_ASSIGN U1191 ( .B(clk), .A(\g.we_clk [31583]));
Q_ASSIGN U1192 ( .B(clk), .A(\g.we_clk [31582]));
Q_ASSIGN U1193 ( .B(clk), .A(\g.we_clk [31581]));
Q_ASSIGN U1194 ( .B(clk), .A(\g.we_clk [31580]));
Q_ASSIGN U1195 ( .B(clk), .A(\g.we_clk [31579]));
Q_ASSIGN U1196 ( .B(clk), .A(\g.we_clk [31578]));
Q_ASSIGN U1197 ( .B(clk), .A(\g.we_clk [31577]));
Q_ASSIGN U1198 ( .B(clk), .A(\g.we_clk [31576]));
Q_ASSIGN U1199 ( .B(clk), .A(\g.we_clk [31575]));
Q_ASSIGN U1200 ( .B(clk), .A(\g.we_clk [31574]));
Q_ASSIGN U1201 ( .B(clk), .A(\g.we_clk [31573]));
Q_ASSIGN U1202 ( .B(clk), .A(\g.we_clk [31572]));
Q_ASSIGN U1203 ( .B(clk), .A(\g.we_clk [31571]));
Q_ASSIGN U1204 ( .B(clk), .A(\g.we_clk [31570]));
Q_ASSIGN U1205 ( .B(clk), .A(\g.we_clk [31569]));
Q_ASSIGN U1206 ( .B(clk), .A(\g.we_clk [31568]));
Q_ASSIGN U1207 ( .B(clk), .A(\g.we_clk [31567]));
Q_ASSIGN U1208 ( .B(clk), .A(\g.we_clk [31566]));
Q_ASSIGN U1209 ( .B(clk), .A(\g.we_clk [31565]));
Q_ASSIGN U1210 ( .B(clk), .A(\g.we_clk [31564]));
Q_ASSIGN U1211 ( .B(clk), .A(\g.we_clk [31563]));
Q_ASSIGN U1212 ( .B(clk), .A(\g.we_clk [31562]));
Q_ASSIGN U1213 ( .B(clk), .A(\g.we_clk [31561]));
Q_ASSIGN U1214 ( .B(clk), .A(\g.we_clk [31560]));
Q_ASSIGN U1215 ( .B(clk), .A(\g.we_clk [31559]));
Q_ASSIGN U1216 ( .B(clk), .A(\g.we_clk [31558]));
Q_ASSIGN U1217 ( .B(clk), .A(\g.we_clk [31557]));
Q_ASSIGN U1218 ( .B(clk), .A(\g.we_clk [31556]));
Q_ASSIGN U1219 ( .B(clk), .A(\g.we_clk [31555]));
Q_ASSIGN U1220 ( .B(clk), .A(\g.we_clk [31554]));
Q_ASSIGN U1221 ( .B(clk), .A(\g.we_clk [31553]));
Q_ASSIGN U1222 ( .B(clk), .A(\g.we_clk [31552]));
Q_ASSIGN U1223 ( .B(clk), .A(\g.we_clk [31551]));
Q_ASSIGN U1224 ( .B(clk), .A(\g.we_clk [31550]));
Q_ASSIGN U1225 ( .B(clk), .A(\g.we_clk [31549]));
Q_ASSIGN U1226 ( .B(clk), .A(\g.we_clk [31548]));
Q_ASSIGN U1227 ( .B(clk), .A(\g.we_clk [31547]));
Q_ASSIGN U1228 ( .B(clk), .A(\g.we_clk [31546]));
Q_ASSIGN U1229 ( .B(clk), .A(\g.we_clk [31545]));
Q_ASSIGN U1230 ( .B(clk), .A(\g.we_clk [31544]));
Q_ASSIGN U1231 ( .B(clk), .A(\g.we_clk [31543]));
Q_ASSIGN U1232 ( .B(clk), .A(\g.we_clk [31542]));
Q_ASSIGN U1233 ( .B(clk), .A(\g.we_clk [31541]));
Q_ASSIGN U1234 ( .B(clk), .A(\g.we_clk [31540]));
Q_ASSIGN U1235 ( .B(clk), .A(\g.we_clk [31539]));
Q_ASSIGN U1236 ( .B(clk), .A(\g.we_clk [31538]));
Q_ASSIGN U1237 ( .B(clk), .A(\g.we_clk [31537]));
Q_ASSIGN U1238 ( .B(clk), .A(\g.we_clk [31536]));
Q_ASSIGN U1239 ( .B(clk), .A(\g.we_clk [31535]));
Q_ASSIGN U1240 ( .B(clk), .A(\g.we_clk [31534]));
Q_ASSIGN U1241 ( .B(clk), .A(\g.we_clk [31533]));
Q_ASSIGN U1242 ( .B(clk), .A(\g.we_clk [31532]));
Q_ASSIGN U1243 ( .B(clk), .A(\g.we_clk [31531]));
Q_ASSIGN U1244 ( .B(clk), .A(\g.we_clk [31530]));
Q_ASSIGN U1245 ( .B(clk), .A(\g.we_clk [31529]));
Q_ASSIGN U1246 ( .B(clk), .A(\g.we_clk [31528]));
Q_ASSIGN U1247 ( .B(clk), .A(\g.we_clk [31527]));
Q_ASSIGN U1248 ( .B(clk), .A(\g.we_clk [31526]));
Q_ASSIGN U1249 ( .B(clk), .A(\g.we_clk [31525]));
Q_ASSIGN U1250 ( .B(clk), .A(\g.we_clk [31524]));
Q_ASSIGN U1251 ( .B(clk), .A(\g.we_clk [31523]));
Q_ASSIGN U1252 ( .B(clk), .A(\g.we_clk [31522]));
Q_ASSIGN U1253 ( .B(clk), .A(\g.we_clk [31521]));
Q_ASSIGN U1254 ( .B(clk), .A(\g.we_clk [31520]));
Q_ASSIGN U1255 ( .B(clk), .A(\g.we_clk [31519]));
Q_ASSIGN U1256 ( .B(clk), .A(\g.we_clk [31518]));
Q_ASSIGN U1257 ( .B(clk), .A(\g.we_clk [31517]));
Q_ASSIGN U1258 ( .B(clk), .A(\g.we_clk [31516]));
Q_ASSIGN U1259 ( .B(clk), .A(\g.we_clk [31515]));
Q_ASSIGN U1260 ( .B(clk), .A(\g.we_clk [31514]));
Q_ASSIGN U1261 ( .B(clk), .A(\g.we_clk [31513]));
Q_ASSIGN U1262 ( .B(clk), .A(\g.we_clk [31512]));
Q_ASSIGN U1263 ( .B(clk), .A(\g.we_clk [31511]));
Q_ASSIGN U1264 ( .B(clk), .A(\g.we_clk [31510]));
Q_ASSIGN U1265 ( .B(clk), .A(\g.we_clk [31509]));
Q_ASSIGN U1266 ( .B(clk), .A(\g.we_clk [31508]));
Q_ASSIGN U1267 ( .B(clk), .A(\g.we_clk [31507]));
Q_ASSIGN U1268 ( .B(clk), .A(\g.we_clk [31506]));
Q_ASSIGN U1269 ( .B(clk), .A(\g.we_clk [31505]));
Q_ASSIGN U1270 ( .B(clk), .A(\g.we_clk [31504]));
Q_ASSIGN U1271 ( .B(clk), .A(\g.we_clk [31503]));
Q_ASSIGN U1272 ( .B(clk), .A(\g.we_clk [31502]));
Q_ASSIGN U1273 ( .B(clk), .A(\g.we_clk [31501]));
Q_ASSIGN U1274 ( .B(clk), .A(\g.we_clk [31500]));
Q_ASSIGN U1275 ( .B(clk), .A(\g.we_clk [31499]));
Q_ASSIGN U1276 ( .B(clk), .A(\g.we_clk [31498]));
Q_ASSIGN U1277 ( .B(clk), .A(\g.we_clk [31497]));
Q_ASSIGN U1278 ( .B(clk), .A(\g.we_clk [31496]));
Q_ASSIGN U1279 ( .B(clk), .A(\g.we_clk [31495]));
Q_ASSIGN U1280 ( .B(clk), .A(\g.we_clk [31494]));
Q_ASSIGN U1281 ( .B(clk), .A(\g.we_clk [31493]));
Q_ASSIGN U1282 ( .B(clk), .A(\g.we_clk [31492]));
Q_ASSIGN U1283 ( .B(clk), .A(\g.we_clk [31491]));
Q_ASSIGN U1284 ( .B(clk), .A(\g.we_clk [31490]));
Q_ASSIGN U1285 ( .B(clk), .A(\g.we_clk [31489]));
Q_ASSIGN U1286 ( .B(clk), .A(\g.we_clk [31488]));
Q_ASSIGN U1287 ( .B(clk), .A(\g.we_clk [31487]));
Q_ASSIGN U1288 ( .B(clk), .A(\g.we_clk [31486]));
Q_ASSIGN U1289 ( .B(clk), .A(\g.we_clk [31485]));
Q_ASSIGN U1290 ( .B(clk), .A(\g.we_clk [31484]));
Q_ASSIGN U1291 ( .B(clk), .A(\g.we_clk [31483]));
Q_ASSIGN U1292 ( .B(clk), .A(\g.we_clk [31482]));
Q_ASSIGN U1293 ( .B(clk), .A(\g.we_clk [31481]));
Q_ASSIGN U1294 ( .B(clk), .A(\g.we_clk [31480]));
Q_ASSIGN U1295 ( .B(clk), .A(\g.we_clk [31479]));
Q_ASSIGN U1296 ( .B(clk), .A(\g.we_clk [31478]));
Q_ASSIGN U1297 ( .B(clk), .A(\g.we_clk [31477]));
Q_ASSIGN U1298 ( .B(clk), .A(\g.we_clk [31476]));
Q_ASSIGN U1299 ( .B(clk), .A(\g.we_clk [31475]));
Q_ASSIGN U1300 ( .B(clk), .A(\g.we_clk [31474]));
Q_ASSIGN U1301 ( .B(clk), .A(\g.we_clk [31473]));
Q_ASSIGN U1302 ( .B(clk), .A(\g.we_clk [31472]));
Q_ASSIGN U1303 ( .B(clk), .A(\g.we_clk [31471]));
Q_ASSIGN U1304 ( .B(clk), .A(\g.we_clk [31470]));
Q_ASSIGN U1305 ( .B(clk), .A(\g.we_clk [31469]));
Q_ASSIGN U1306 ( .B(clk), .A(\g.we_clk [31468]));
Q_ASSIGN U1307 ( .B(clk), .A(\g.we_clk [31467]));
Q_ASSIGN U1308 ( .B(clk), .A(\g.we_clk [31466]));
Q_ASSIGN U1309 ( .B(clk), .A(\g.we_clk [31465]));
Q_ASSIGN U1310 ( .B(clk), .A(\g.we_clk [31464]));
Q_ASSIGN U1311 ( .B(clk), .A(\g.we_clk [31463]));
Q_ASSIGN U1312 ( .B(clk), .A(\g.we_clk [31462]));
Q_ASSIGN U1313 ( .B(clk), .A(\g.we_clk [31461]));
Q_ASSIGN U1314 ( .B(clk), .A(\g.we_clk [31460]));
Q_ASSIGN U1315 ( .B(clk), .A(\g.we_clk [31459]));
Q_ASSIGN U1316 ( .B(clk), .A(\g.we_clk [31458]));
Q_ASSIGN U1317 ( .B(clk), .A(\g.we_clk [31457]));
Q_ASSIGN U1318 ( .B(clk), .A(\g.we_clk [31456]));
Q_ASSIGN U1319 ( .B(clk), .A(\g.we_clk [31455]));
Q_ASSIGN U1320 ( .B(clk), .A(\g.we_clk [31454]));
Q_ASSIGN U1321 ( .B(clk), .A(\g.we_clk [31453]));
Q_ASSIGN U1322 ( .B(clk), .A(\g.we_clk [31452]));
Q_ASSIGN U1323 ( .B(clk), .A(\g.we_clk [31451]));
Q_ASSIGN U1324 ( .B(clk), .A(\g.we_clk [31450]));
Q_ASSIGN U1325 ( .B(clk), .A(\g.we_clk [31449]));
Q_ASSIGN U1326 ( .B(clk), .A(\g.we_clk [31448]));
Q_ASSIGN U1327 ( .B(clk), .A(\g.we_clk [31447]));
Q_ASSIGN U1328 ( .B(clk), .A(\g.we_clk [31446]));
Q_ASSIGN U1329 ( .B(clk), .A(\g.we_clk [31445]));
Q_ASSIGN U1330 ( .B(clk), .A(\g.we_clk [31444]));
Q_ASSIGN U1331 ( .B(clk), .A(\g.we_clk [31443]));
Q_ASSIGN U1332 ( .B(clk), .A(\g.we_clk [31442]));
Q_ASSIGN U1333 ( .B(clk), .A(\g.we_clk [31441]));
Q_ASSIGN U1334 ( .B(clk), .A(\g.we_clk [31440]));
Q_ASSIGN U1335 ( .B(clk), .A(\g.we_clk [31439]));
Q_ASSIGN U1336 ( .B(clk), .A(\g.we_clk [31438]));
Q_ASSIGN U1337 ( .B(clk), .A(\g.we_clk [31437]));
Q_ASSIGN U1338 ( .B(clk), .A(\g.we_clk [31436]));
Q_ASSIGN U1339 ( .B(clk), .A(\g.we_clk [31435]));
Q_ASSIGN U1340 ( .B(clk), .A(\g.we_clk [31434]));
Q_ASSIGN U1341 ( .B(clk), .A(\g.we_clk [31433]));
Q_ASSIGN U1342 ( .B(clk), .A(\g.we_clk [31432]));
Q_ASSIGN U1343 ( .B(clk), .A(\g.we_clk [31431]));
Q_ASSIGN U1344 ( .B(clk), .A(\g.we_clk [31430]));
Q_ASSIGN U1345 ( .B(clk), .A(\g.we_clk [31429]));
Q_ASSIGN U1346 ( .B(clk), .A(\g.we_clk [31428]));
Q_ASSIGN U1347 ( .B(clk), .A(\g.we_clk [31427]));
Q_ASSIGN U1348 ( .B(clk), .A(\g.we_clk [31426]));
Q_ASSIGN U1349 ( .B(clk), .A(\g.we_clk [31425]));
Q_ASSIGN U1350 ( .B(clk), .A(\g.we_clk [31424]));
Q_ASSIGN U1351 ( .B(clk), .A(\g.we_clk [31423]));
Q_ASSIGN U1352 ( .B(clk), .A(\g.we_clk [31422]));
Q_ASSIGN U1353 ( .B(clk), .A(\g.we_clk [31421]));
Q_ASSIGN U1354 ( .B(clk), .A(\g.we_clk [31420]));
Q_ASSIGN U1355 ( .B(clk), .A(\g.we_clk [31419]));
Q_ASSIGN U1356 ( .B(clk), .A(\g.we_clk [31418]));
Q_ASSIGN U1357 ( .B(clk), .A(\g.we_clk [31417]));
Q_ASSIGN U1358 ( .B(clk), .A(\g.we_clk [31416]));
Q_ASSIGN U1359 ( .B(clk), .A(\g.we_clk [31415]));
Q_ASSIGN U1360 ( .B(clk), .A(\g.we_clk [31414]));
Q_ASSIGN U1361 ( .B(clk), .A(\g.we_clk [31413]));
Q_ASSIGN U1362 ( .B(clk), .A(\g.we_clk [31412]));
Q_ASSIGN U1363 ( .B(clk), .A(\g.we_clk [31411]));
Q_ASSIGN U1364 ( .B(clk), .A(\g.we_clk [31410]));
Q_ASSIGN U1365 ( .B(clk), .A(\g.we_clk [31409]));
Q_ASSIGN U1366 ( .B(clk), .A(\g.we_clk [31408]));
Q_ASSIGN U1367 ( .B(clk), .A(\g.we_clk [31407]));
Q_ASSIGN U1368 ( .B(clk), .A(\g.we_clk [31406]));
Q_ASSIGN U1369 ( .B(clk), .A(\g.we_clk [31405]));
Q_ASSIGN U1370 ( .B(clk), .A(\g.we_clk [31404]));
Q_ASSIGN U1371 ( .B(clk), .A(\g.we_clk [31403]));
Q_ASSIGN U1372 ( .B(clk), .A(\g.we_clk [31402]));
Q_ASSIGN U1373 ( .B(clk), .A(\g.we_clk [31401]));
Q_ASSIGN U1374 ( .B(clk), .A(\g.we_clk [31400]));
Q_ASSIGN U1375 ( .B(clk), .A(\g.we_clk [31399]));
Q_ASSIGN U1376 ( .B(clk), .A(\g.we_clk [31398]));
Q_ASSIGN U1377 ( .B(clk), .A(\g.we_clk [31397]));
Q_ASSIGN U1378 ( .B(clk), .A(\g.we_clk [31396]));
Q_ASSIGN U1379 ( .B(clk), .A(\g.we_clk [31395]));
Q_ASSIGN U1380 ( .B(clk), .A(\g.we_clk [31394]));
Q_ASSIGN U1381 ( .B(clk), .A(\g.we_clk [31393]));
Q_ASSIGN U1382 ( .B(clk), .A(\g.we_clk [31392]));
Q_ASSIGN U1383 ( .B(clk), .A(\g.we_clk [31391]));
Q_ASSIGN U1384 ( .B(clk), .A(\g.we_clk [31390]));
Q_ASSIGN U1385 ( .B(clk), .A(\g.we_clk [31389]));
Q_ASSIGN U1386 ( .B(clk), .A(\g.we_clk [31388]));
Q_ASSIGN U1387 ( .B(clk), .A(\g.we_clk [31387]));
Q_ASSIGN U1388 ( .B(clk), .A(\g.we_clk [31386]));
Q_ASSIGN U1389 ( .B(clk), .A(\g.we_clk [31385]));
Q_ASSIGN U1390 ( .B(clk), .A(\g.we_clk [31384]));
Q_ASSIGN U1391 ( .B(clk), .A(\g.we_clk [31383]));
Q_ASSIGN U1392 ( .B(clk), .A(\g.we_clk [31382]));
Q_ASSIGN U1393 ( .B(clk), .A(\g.we_clk [31381]));
Q_ASSIGN U1394 ( .B(clk), .A(\g.we_clk [31380]));
Q_ASSIGN U1395 ( .B(clk), .A(\g.we_clk [31379]));
Q_ASSIGN U1396 ( .B(clk), .A(\g.we_clk [31378]));
Q_ASSIGN U1397 ( .B(clk), .A(\g.we_clk [31377]));
Q_ASSIGN U1398 ( .B(clk), .A(\g.we_clk [31376]));
Q_ASSIGN U1399 ( .B(clk), .A(\g.we_clk [31375]));
Q_ASSIGN U1400 ( .B(clk), .A(\g.we_clk [31374]));
Q_ASSIGN U1401 ( .B(clk), .A(\g.we_clk [31373]));
Q_ASSIGN U1402 ( .B(clk), .A(\g.we_clk [31372]));
Q_ASSIGN U1403 ( .B(clk), .A(\g.we_clk [31371]));
Q_ASSIGN U1404 ( .B(clk), .A(\g.we_clk [31370]));
Q_ASSIGN U1405 ( .B(clk), .A(\g.we_clk [31369]));
Q_ASSIGN U1406 ( .B(clk), .A(\g.we_clk [31368]));
Q_ASSIGN U1407 ( .B(clk), .A(\g.we_clk [31367]));
Q_ASSIGN U1408 ( .B(clk), .A(\g.we_clk [31366]));
Q_ASSIGN U1409 ( .B(clk), .A(\g.we_clk [31365]));
Q_ASSIGN U1410 ( .B(clk), .A(\g.we_clk [31364]));
Q_ASSIGN U1411 ( .B(clk), .A(\g.we_clk [31363]));
Q_ASSIGN U1412 ( .B(clk), .A(\g.we_clk [31362]));
Q_ASSIGN U1413 ( .B(clk), .A(\g.we_clk [31361]));
Q_ASSIGN U1414 ( .B(clk), .A(\g.we_clk [31360]));
Q_ASSIGN U1415 ( .B(clk), .A(\g.we_clk [31359]));
Q_ASSIGN U1416 ( .B(clk), .A(\g.we_clk [31358]));
Q_ASSIGN U1417 ( .B(clk), .A(\g.we_clk [31357]));
Q_ASSIGN U1418 ( .B(clk), .A(\g.we_clk [31356]));
Q_ASSIGN U1419 ( .B(clk), .A(\g.we_clk [31355]));
Q_ASSIGN U1420 ( .B(clk), .A(\g.we_clk [31354]));
Q_ASSIGN U1421 ( .B(clk), .A(\g.we_clk [31353]));
Q_ASSIGN U1422 ( .B(clk), .A(\g.we_clk [31352]));
Q_ASSIGN U1423 ( .B(clk), .A(\g.we_clk [31351]));
Q_ASSIGN U1424 ( .B(clk), .A(\g.we_clk [31350]));
Q_ASSIGN U1425 ( .B(clk), .A(\g.we_clk [31349]));
Q_ASSIGN U1426 ( .B(clk), .A(\g.we_clk [31348]));
Q_ASSIGN U1427 ( .B(clk), .A(\g.we_clk [31347]));
Q_ASSIGN U1428 ( .B(clk), .A(\g.we_clk [31346]));
Q_ASSIGN U1429 ( .B(clk), .A(\g.we_clk [31345]));
Q_ASSIGN U1430 ( .B(clk), .A(\g.we_clk [31344]));
Q_ASSIGN U1431 ( .B(clk), .A(\g.we_clk [31343]));
Q_ASSIGN U1432 ( .B(clk), .A(\g.we_clk [31342]));
Q_ASSIGN U1433 ( .B(clk), .A(\g.we_clk [31341]));
Q_ASSIGN U1434 ( .B(clk), .A(\g.we_clk [31340]));
Q_ASSIGN U1435 ( .B(clk), .A(\g.we_clk [31339]));
Q_ASSIGN U1436 ( .B(clk), .A(\g.we_clk [31338]));
Q_ASSIGN U1437 ( .B(clk), .A(\g.we_clk [31337]));
Q_ASSIGN U1438 ( .B(clk), .A(\g.we_clk [31336]));
Q_ASSIGN U1439 ( .B(clk), .A(\g.we_clk [31335]));
Q_ASSIGN U1440 ( .B(clk), .A(\g.we_clk [31334]));
Q_ASSIGN U1441 ( .B(clk), .A(\g.we_clk [31333]));
Q_ASSIGN U1442 ( .B(clk), .A(\g.we_clk [31332]));
Q_ASSIGN U1443 ( .B(clk), .A(\g.we_clk [31331]));
Q_ASSIGN U1444 ( .B(clk), .A(\g.we_clk [31330]));
Q_ASSIGN U1445 ( .B(clk), .A(\g.we_clk [31329]));
Q_ASSIGN U1446 ( .B(clk), .A(\g.we_clk [31328]));
Q_ASSIGN U1447 ( .B(clk), .A(\g.we_clk [31327]));
Q_ASSIGN U1448 ( .B(clk), .A(\g.we_clk [31326]));
Q_ASSIGN U1449 ( .B(clk), .A(\g.we_clk [31325]));
Q_ASSIGN U1450 ( .B(clk), .A(\g.we_clk [31324]));
Q_ASSIGN U1451 ( .B(clk), .A(\g.we_clk [31323]));
Q_ASSIGN U1452 ( .B(clk), .A(\g.we_clk [31322]));
Q_ASSIGN U1453 ( .B(clk), .A(\g.we_clk [31321]));
Q_ASSIGN U1454 ( .B(clk), .A(\g.we_clk [31320]));
Q_ASSIGN U1455 ( .B(clk), .A(\g.we_clk [31319]));
Q_ASSIGN U1456 ( .B(clk), .A(\g.we_clk [31318]));
Q_ASSIGN U1457 ( .B(clk), .A(\g.we_clk [31317]));
Q_ASSIGN U1458 ( .B(clk), .A(\g.we_clk [31316]));
Q_ASSIGN U1459 ( .B(clk), .A(\g.we_clk [31315]));
Q_ASSIGN U1460 ( .B(clk), .A(\g.we_clk [31314]));
Q_ASSIGN U1461 ( .B(clk), .A(\g.we_clk [31313]));
Q_ASSIGN U1462 ( .B(clk), .A(\g.we_clk [31312]));
Q_ASSIGN U1463 ( .B(clk), .A(\g.we_clk [31311]));
Q_ASSIGN U1464 ( .B(clk), .A(\g.we_clk [31310]));
Q_ASSIGN U1465 ( .B(clk), .A(\g.we_clk [31309]));
Q_ASSIGN U1466 ( .B(clk), .A(\g.we_clk [31308]));
Q_ASSIGN U1467 ( .B(clk), .A(\g.we_clk [31307]));
Q_ASSIGN U1468 ( .B(clk), .A(\g.we_clk [31306]));
Q_ASSIGN U1469 ( .B(clk), .A(\g.we_clk [31305]));
Q_ASSIGN U1470 ( .B(clk), .A(\g.we_clk [31304]));
Q_ASSIGN U1471 ( .B(clk), .A(\g.we_clk [31303]));
Q_ASSIGN U1472 ( .B(clk), .A(\g.we_clk [31302]));
Q_ASSIGN U1473 ( .B(clk), .A(\g.we_clk [31301]));
Q_ASSIGN U1474 ( .B(clk), .A(\g.we_clk [31300]));
Q_ASSIGN U1475 ( .B(clk), .A(\g.we_clk [31299]));
Q_ASSIGN U1476 ( .B(clk), .A(\g.we_clk [31298]));
Q_ASSIGN U1477 ( .B(clk), .A(\g.we_clk [31297]));
Q_ASSIGN U1478 ( .B(clk), .A(\g.we_clk [31296]));
Q_ASSIGN U1479 ( .B(clk), .A(\g.we_clk [31295]));
Q_ASSIGN U1480 ( .B(clk), .A(\g.we_clk [31294]));
Q_ASSIGN U1481 ( .B(clk), .A(\g.we_clk [31293]));
Q_ASSIGN U1482 ( .B(clk), .A(\g.we_clk [31292]));
Q_ASSIGN U1483 ( .B(clk), .A(\g.we_clk [31291]));
Q_ASSIGN U1484 ( .B(clk), .A(\g.we_clk [31290]));
Q_ASSIGN U1485 ( .B(clk), .A(\g.we_clk [31289]));
Q_ASSIGN U1486 ( .B(clk), .A(\g.we_clk [31288]));
Q_ASSIGN U1487 ( .B(clk), .A(\g.we_clk [31287]));
Q_ASSIGN U1488 ( .B(clk), .A(\g.we_clk [31286]));
Q_ASSIGN U1489 ( .B(clk), .A(\g.we_clk [31285]));
Q_ASSIGN U1490 ( .B(clk), .A(\g.we_clk [31284]));
Q_ASSIGN U1491 ( .B(clk), .A(\g.we_clk [31283]));
Q_ASSIGN U1492 ( .B(clk), .A(\g.we_clk [31282]));
Q_ASSIGN U1493 ( .B(clk), .A(\g.we_clk [31281]));
Q_ASSIGN U1494 ( .B(clk), .A(\g.we_clk [31280]));
Q_ASSIGN U1495 ( .B(clk), .A(\g.we_clk [31279]));
Q_ASSIGN U1496 ( .B(clk), .A(\g.we_clk [31278]));
Q_ASSIGN U1497 ( .B(clk), .A(\g.we_clk [31277]));
Q_ASSIGN U1498 ( .B(clk), .A(\g.we_clk [31276]));
Q_ASSIGN U1499 ( .B(clk), .A(\g.we_clk [31275]));
Q_ASSIGN U1500 ( .B(clk), .A(\g.we_clk [31274]));
Q_ASSIGN U1501 ( .B(clk), .A(\g.we_clk [31273]));
Q_ASSIGN U1502 ( .B(clk), .A(\g.we_clk [31272]));
Q_ASSIGN U1503 ( .B(clk), .A(\g.we_clk [31271]));
Q_ASSIGN U1504 ( .B(clk), .A(\g.we_clk [31270]));
Q_ASSIGN U1505 ( .B(clk), .A(\g.we_clk [31269]));
Q_ASSIGN U1506 ( .B(clk), .A(\g.we_clk [31268]));
Q_ASSIGN U1507 ( .B(clk), .A(\g.we_clk [31267]));
Q_ASSIGN U1508 ( .B(clk), .A(\g.we_clk [31266]));
Q_ASSIGN U1509 ( .B(clk), .A(\g.we_clk [31265]));
Q_ASSIGN U1510 ( .B(clk), .A(\g.we_clk [31264]));
Q_ASSIGN U1511 ( .B(clk), .A(\g.we_clk [31263]));
Q_ASSIGN U1512 ( .B(clk), .A(\g.we_clk [31262]));
Q_ASSIGN U1513 ( .B(clk), .A(\g.we_clk [31261]));
Q_ASSIGN U1514 ( .B(clk), .A(\g.we_clk [31260]));
Q_ASSIGN U1515 ( .B(clk), .A(\g.we_clk [31259]));
Q_ASSIGN U1516 ( .B(clk), .A(\g.we_clk [31258]));
Q_ASSIGN U1517 ( .B(clk), .A(\g.we_clk [31257]));
Q_ASSIGN U1518 ( .B(clk), .A(\g.we_clk [31256]));
Q_ASSIGN U1519 ( .B(clk), .A(\g.we_clk [31255]));
Q_ASSIGN U1520 ( .B(clk), .A(\g.we_clk [31254]));
Q_ASSIGN U1521 ( .B(clk), .A(\g.we_clk [31253]));
Q_ASSIGN U1522 ( .B(clk), .A(\g.we_clk [31252]));
Q_ASSIGN U1523 ( .B(clk), .A(\g.we_clk [31251]));
Q_ASSIGN U1524 ( .B(clk), .A(\g.we_clk [31250]));
Q_ASSIGN U1525 ( .B(clk), .A(\g.we_clk [31249]));
Q_ASSIGN U1526 ( .B(clk), .A(\g.we_clk [31248]));
Q_ASSIGN U1527 ( .B(clk), .A(\g.we_clk [31247]));
Q_ASSIGN U1528 ( .B(clk), .A(\g.we_clk [31246]));
Q_ASSIGN U1529 ( .B(clk), .A(\g.we_clk [31245]));
Q_ASSIGN U1530 ( .B(clk), .A(\g.we_clk [31244]));
Q_ASSIGN U1531 ( .B(clk), .A(\g.we_clk [31243]));
Q_ASSIGN U1532 ( .B(clk), .A(\g.we_clk [31242]));
Q_ASSIGN U1533 ( .B(clk), .A(\g.we_clk [31241]));
Q_ASSIGN U1534 ( .B(clk), .A(\g.we_clk [31240]));
Q_ASSIGN U1535 ( .B(clk), .A(\g.we_clk [31239]));
Q_ASSIGN U1536 ( .B(clk), .A(\g.we_clk [31238]));
Q_ASSIGN U1537 ( .B(clk), .A(\g.we_clk [31237]));
Q_ASSIGN U1538 ( .B(clk), .A(\g.we_clk [31236]));
Q_ASSIGN U1539 ( .B(clk), .A(\g.we_clk [31235]));
Q_ASSIGN U1540 ( .B(clk), .A(\g.we_clk [31234]));
Q_ASSIGN U1541 ( .B(clk), .A(\g.we_clk [31233]));
Q_ASSIGN U1542 ( .B(clk), .A(\g.we_clk [31232]));
Q_ASSIGN U1543 ( .B(clk), .A(\g.we_clk [31231]));
Q_ASSIGN U1544 ( .B(clk), .A(\g.we_clk [31230]));
Q_ASSIGN U1545 ( .B(clk), .A(\g.we_clk [31229]));
Q_ASSIGN U1546 ( .B(clk), .A(\g.we_clk [31228]));
Q_ASSIGN U1547 ( .B(clk), .A(\g.we_clk [31227]));
Q_ASSIGN U1548 ( .B(clk), .A(\g.we_clk [31226]));
Q_ASSIGN U1549 ( .B(clk), .A(\g.we_clk [31225]));
Q_ASSIGN U1550 ( .B(clk), .A(\g.we_clk [31224]));
Q_ASSIGN U1551 ( .B(clk), .A(\g.we_clk [31223]));
Q_ASSIGN U1552 ( .B(clk), .A(\g.we_clk [31222]));
Q_ASSIGN U1553 ( .B(clk), .A(\g.we_clk [31221]));
Q_ASSIGN U1554 ( .B(clk), .A(\g.we_clk [31220]));
Q_ASSIGN U1555 ( .B(clk), .A(\g.we_clk [31219]));
Q_ASSIGN U1556 ( .B(clk), .A(\g.we_clk [31218]));
Q_ASSIGN U1557 ( .B(clk), .A(\g.we_clk [31217]));
Q_ASSIGN U1558 ( .B(clk), .A(\g.we_clk [31216]));
Q_ASSIGN U1559 ( .B(clk), .A(\g.we_clk [31215]));
Q_ASSIGN U1560 ( .B(clk), .A(\g.we_clk [31214]));
Q_ASSIGN U1561 ( .B(clk), .A(\g.we_clk [31213]));
Q_ASSIGN U1562 ( .B(clk), .A(\g.we_clk [31212]));
Q_ASSIGN U1563 ( .B(clk), .A(\g.we_clk [31211]));
Q_ASSIGN U1564 ( .B(clk), .A(\g.we_clk [31210]));
Q_ASSIGN U1565 ( .B(clk), .A(\g.we_clk [31209]));
Q_ASSIGN U1566 ( .B(clk), .A(\g.we_clk [31208]));
Q_ASSIGN U1567 ( .B(clk), .A(\g.we_clk [31207]));
Q_ASSIGN U1568 ( .B(clk), .A(\g.we_clk [31206]));
Q_ASSIGN U1569 ( .B(clk), .A(\g.we_clk [31205]));
Q_ASSIGN U1570 ( .B(clk), .A(\g.we_clk [31204]));
Q_ASSIGN U1571 ( .B(clk), .A(\g.we_clk [31203]));
Q_ASSIGN U1572 ( .B(clk), .A(\g.we_clk [31202]));
Q_ASSIGN U1573 ( .B(clk), .A(\g.we_clk [31201]));
Q_ASSIGN U1574 ( .B(clk), .A(\g.we_clk [31200]));
Q_ASSIGN U1575 ( .B(clk), .A(\g.we_clk [31199]));
Q_ASSIGN U1576 ( .B(clk), .A(\g.we_clk [31198]));
Q_ASSIGN U1577 ( .B(clk), .A(\g.we_clk [31197]));
Q_ASSIGN U1578 ( .B(clk), .A(\g.we_clk [31196]));
Q_ASSIGN U1579 ( .B(clk), .A(\g.we_clk [31195]));
Q_ASSIGN U1580 ( .B(clk), .A(\g.we_clk [31194]));
Q_ASSIGN U1581 ( .B(clk), .A(\g.we_clk [31193]));
Q_ASSIGN U1582 ( .B(clk), .A(\g.we_clk [31192]));
Q_ASSIGN U1583 ( .B(clk), .A(\g.we_clk [31191]));
Q_ASSIGN U1584 ( .B(clk), .A(\g.we_clk [31190]));
Q_ASSIGN U1585 ( .B(clk), .A(\g.we_clk [31189]));
Q_ASSIGN U1586 ( .B(clk), .A(\g.we_clk [31188]));
Q_ASSIGN U1587 ( .B(clk), .A(\g.we_clk [31187]));
Q_ASSIGN U1588 ( .B(clk), .A(\g.we_clk [31186]));
Q_ASSIGN U1589 ( .B(clk), .A(\g.we_clk [31185]));
Q_ASSIGN U1590 ( .B(clk), .A(\g.we_clk [31184]));
Q_ASSIGN U1591 ( .B(clk), .A(\g.we_clk [31183]));
Q_ASSIGN U1592 ( .B(clk), .A(\g.we_clk [31182]));
Q_ASSIGN U1593 ( .B(clk), .A(\g.we_clk [31181]));
Q_ASSIGN U1594 ( .B(clk), .A(\g.we_clk [31180]));
Q_ASSIGN U1595 ( .B(clk), .A(\g.we_clk [31179]));
Q_ASSIGN U1596 ( .B(clk), .A(\g.we_clk [31178]));
Q_ASSIGN U1597 ( .B(clk), .A(\g.we_clk [31177]));
Q_ASSIGN U1598 ( .B(clk), .A(\g.we_clk [31176]));
Q_ASSIGN U1599 ( .B(clk), .A(\g.we_clk [31175]));
Q_ASSIGN U1600 ( .B(clk), .A(\g.we_clk [31174]));
Q_ASSIGN U1601 ( .B(clk), .A(\g.we_clk [31173]));
Q_ASSIGN U1602 ( .B(clk), .A(\g.we_clk [31172]));
Q_ASSIGN U1603 ( .B(clk), .A(\g.we_clk [31171]));
Q_ASSIGN U1604 ( .B(clk), .A(\g.we_clk [31170]));
Q_ASSIGN U1605 ( .B(clk), .A(\g.we_clk [31169]));
Q_ASSIGN U1606 ( .B(clk), .A(\g.we_clk [31168]));
Q_ASSIGN U1607 ( .B(clk), .A(\g.we_clk [31167]));
Q_ASSIGN U1608 ( .B(clk), .A(\g.we_clk [31166]));
Q_ASSIGN U1609 ( .B(clk), .A(\g.we_clk [31165]));
Q_ASSIGN U1610 ( .B(clk), .A(\g.we_clk [31164]));
Q_ASSIGN U1611 ( .B(clk), .A(\g.we_clk [31163]));
Q_ASSIGN U1612 ( .B(clk), .A(\g.we_clk [31162]));
Q_ASSIGN U1613 ( .B(clk), .A(\g.we_clk [31161]));
Q_ASSIGN U1614 ( .B(clk), .A(\g.we_clk [31160]));
Q_ASSIGN U1615 ( .B(clk), .A(\g.we_clk [31159]));
Q_ASSIGN U1616 ( .B(clk), .A(\g.we_clk [31158]));
Q_ASSIGN U1617 ( .B(clk), .A(\g.we_clk [31157]));
Q_ASSIGN U1618 ( .B(clk), .A(\g.we_clk [31156]));
Q_ASSIGN U1619 ( .B(clk), .A(\g.we_clk [31155]));
Q_ASSIGN U1620 ( .B(clk), .A(\g.we_clk [31154]));
Q_ASSIGN U1621 ( .B(clk), .A(\g.we_clk [31153]));
Q_ASSIGN U1622 ( .B(clk), .A(\g.we_clk [31152]));
Q_ASSIGN U1623 ( .B(clk), .A(\g.we_clk [31151]));
Q_ASSIGN U1624 ( .B(clk), .A(\g.we_clk [31150]));
Q_ASSIGN U1625 ( .B(clk), .A(\g.we_clk [31149]));
Q_ASSIGN U1626 ( .B(clk), .A(\g.we_clk [31148]));
Q_ASSIGN U1627 ( .B(clk), .A(\g.we_clk [31147]));
Q_ASSIGN U1628 ( .B(clk), .A(\g.we_clk [31146]));
Q_ASSIGN U1629 ( .B(clk), .A(\g.we_clk [31145]));
Q_ASSIGN U1630 ( .B(clk), .A(\g.we_clk [31144]));
Q_ASSIGN U1631 ( .B(clk), .A(\g.we_clk [31143]));
Q_ASSIGN U1632 ( .B(clk), .A(\g.we_clk [31142]));
Q_ASSIGN U1633 ( .B(clk), .A(\g.we_clk [31141]));
Q_ASSIGN U1634 ( .B(clk), .A(\g.we_clk [31140]));
Q_ASSIGN U1635 ( .B(clk), .A(\g.we_clk [31139]));
Q_ASSIGN U1636 ( .B(clk), .A(\g.we_clk [31138]));
Q_ASSIGN U1637 ( .B(clk), .A(\g.we_clk [31137]));
Q_ASSIGN U1638 ( .B(clk), .A(\g.we_clk [31136]));
Q_ASSIGN U1639 ( .B(clk), .A(\g.we_clk [31135]));
Q_ASSIGN U1640 ( .B(clk), .A(\g.we_clk [31134]));
Q_ASSIGN U1641 ( .B(clk), .A(\g.we_clk [31133]));
Q_ASSIGN U1642 ( .B(clk), .A(\g.we_clk [31132]));
Q_ASSIGN U1643 ( .B(clk), .A(\g.we_clk [31131]));
Q_ASSIGN U1644 ( .B(clk), .A(\g.we_clk [31130]));
Q_ASSIGN U1645 ( .B(clk), .A(\g.we_clk [31129]));
Q_ASSIGN U1646 ( .B(clk), .A(\g.we_clk [31128]));
Q_ASSIGN U1647 ( .B(clk), .A(\g.we_clk [31127]));
Q_ASSIGN U1648 ( .B(clk), .A(\g.we_clk [31126]));
Q_ASSIGN U1649 ( .B(clk), .A(\g.we_clk [31125]));
Q_ASSIGN U1650 ( .B(clk), .A(\g.we_clk [31124]));
Q_ASSIGN U1651 ( .B(clk), .A(\g.we_clk [31123]));
Q_ASSIGN U1652 ( .B(clk), .A(\g.we_clk [31122]));
Q_ASSIGN U1653 ( .B(clk), .A(\g.we_clk [31121]));
Q_ASSIGN U1654 ( .B(clk), .A(\g.we_clk [31120]));
Q_ASSIGN U1655 ( .B(clk), .A(\g.we_clk [31119]));
Q_ASSIGN U1656 ( .B(clk), .A(\g.we_clk [31118]));
Q_ASSIGN U1657 ( .B(clk), .A(\g.we_clk [31117]));
Q_ASSIGN U1658 ( .B(clk), .A(\g.we_clk [31116]));
Q_ASSIGN U1659 ( .B(clk), .A(\g.we_clk [31115]));
Q_ASSIGN U1660 ( .B(clk), .A(\g.we_clk [31114]));
Q_ASSIGN U1661 ( .B(clk), .A(\g.we_clk [31113]));
Q_ASSIGN U1662 ( .B(clk), .A(\g.we_clk [31112]));
Q_ASSIGN U1663 ( .B(clk), .A(\g.we_clk [31111]));
Q_ASSIGN U1664 ( .B(clk), .A(\g.we_clk [31110]));
Q_ASSIGN U1665 ( .B(clk), .A(\g.we_clk [31109]));
Q_ASSIGN U1666 ( .B(clk), .A(\g.we_clk [31108]));
Q_ASSIGN U1667 ( .B(clk), .A(\g.we_clk [31107]));
Q_ASSIGN U1668 ( .B(clk), .A(\g.we_clk [31106]));
Q_ASSIGN U1669 ( .B(clk), .A(\g.we_clk [31105]));
Q_ASSIGN U1670 ( .B(clk), .A(\g.we_clk [31104]));
Q_ASSIGN U1671 ( .B(clk), .A(\g.we_clk [31103]));
Q_ASSIGN U1672 ( .B(clk), .A(\g.we_clk [31102]));
Q_ASSIGN U1673 ( .B(clk), .A(\g.we_clk [31101]));
Q_ASSIGN U1674 ( .B(clk), .A(\g.we_clk [31100]));
Q_ASSIGN U1675 ( .B(clk), .A(\g.we_clk [31099]));
Q_ASSIGN U1676 ( .B(clk), .A(\g.we_clk [31098]));
Q_ASSIGN U1677 ( .B(clk), .A(\g.we_clk [31097]));
Q_ASSIGN U1678 ( .B(clk), .A(\g.we_clk [31096]));
Q_ASSIGN U1679 ( .B(clk), .A(\g.we_clk [31095]));
Q_ASSIGN U1680 ( .B(clk), .A(\g.we_clk [31094]));
Q_ASSIGN U1681 ( .B(clk), .A(\g.we_clk [31093]));
Q_ASSIGN U1682 ( .B(clk), .A(\g.we_clk [31092]));
Q_ASSIGN U1683 ( .B(clk), .A(\g.we_clk [31091]));
Q_ASSIGN U1684 ( .B(clk), .A(\g.we_clk [31090]));
Q_ASSIGN U1685 ( .B(clk), .A(\g.we_clk [31089]));
Q_ASSIGN U1686 ( .B(clk), .A(\g.we_clk [31088]));
Q_ASSIGN U1687 ( .B(clk), .A(\g.we_clk [31087]));
Q_ASSIGN U1688 ( .B(clk), .A(\g.we_clk [31086]));
Q_ASSIGN U1689 ( .B(clk), .A(\g.we_clk [31085]));
Q_ASSIGN U1690 ( .B(clk), .A(\g.we_clk [31084]));
Q_ASSIGN U1691 ( .B(clk), .A(\g.we_clk [31083]));
Q_ASSIGN U1692 ( .B(clk), .A(\g.we_clk [31082]));
Q_ASSIGN U1693 ( .B(clk), .A(\g.we_clk [31081]));
Q_ASSIGN U1694 ( .B(clk), .A(\g.we_clk [31080]));
Q_ASSIGN U1695 ( .B(clk), .A(\g.we_clk [31079]));
Q_ASSIGN U1696 ( .B(clk), .A(\g.we_clk [31078]));
Q_ASSIGN U1697 ( .B(clk), .A(\g.we_clk [31077]));
Q_ASSIGN U1698 ( .B(clk), .A(\g.we_clk [31076]));
Q_ASSIGN U1699 ( .B(clk), .A(\g.we_clk [31075]));
Q_ASSIGN U1700 ( .B(clk), .A(\g.we_clk [31074]));
Q_ASSIGN U1701 ( .B(clk), .A(\g.we_clk [31073]));
Q_ASSIGN U1702 ( .B(clk), .A(\g.we_clk [31072]));
Q_ASSIGN U1703 ( .B(clk), .A(\g.we_clk [31071]));
Q_ASSIGN U1704 ( .B(clk), .A(\g.we_clk [31070]));
Q_ASSIGN U1705 ( .B(clk), .A(\g.we_clk [31069]));
Q_ASSIGN U1706 ( .B(clk), .A(\g.we_clk [31068]));
Q_ASSIGN U1707 ( .B(clk), .A(\g.we_clk [31067]));
Q_ASSIGN U1708 ( .B(clk), .A(\g.we_clk [31066]));
Q_ASSIGN U1709 ( .B(clk), .A(\g.we_clk [31065]));
Q_ASSIGN U1710 ( .B(clk), .A(\g.we_clk [31064]));
Q_ASSIGN U1711 ( .B(clk), .A(\g.we_clk [31063]));
Q_ASSIGN U1712 ( .B(clk), .A(\g.we_clk [31062]));
Q_ASSIGN U1713 ( .B(clk), .A(\g.we_clk [31061]));
Q_ASSIGN U1714 ( .B(clk), .A(\g.we_clk [31060]));
Q_ASSIGN U1715 ( .B(clk), .A(\g.we_clk [31059]));
Q_ASSIGN U1716 ( .B(clk), .A(\g.we_clk [31058]));
Q_ASSIGN U1717 ( .B(clk), .A(\g.we_clk [31057]));
Q_ASSIGN U1718 ( .B(clk), .A(\g.we_clk [31056]));
Q_ASSIGN U1719 ( .B(clk), .A(\g.we_clk [31055]));
Q_ASSIGN U1720 ( .B(clk), .A(\g.we_clk [31054]));
Q_ASSIGN U1721 ( .B(clk), .A(\g.we_clk [31053]));
Q_ASSIGN U1722 ( .B(clk), .A(\g.we_clk [31052]));
Q_ASSIGN U1723 ( .B(clk), .A(\g.we_clk [31051]));
Q_ASSIGN U1724 ( .B(clk), .A(\g.we_clk [31050]));
Q_ASSIGN U1725 ( .B(clk), .A(\g.we_clk [31049]));
Q_ASSIGN U1726 ( .B(clk), .A(\g.we_clk [31048]));
Q_ASSIGN U1727 ( .B(clk), .A(\g.we_clk [31047]));
Q_ASSIGN U1728 ( .B(clk), .A(\g.we_clk [31046]));
Q_ASSIGN U1729 ( .B(clk), .A(\g.we_clk [31045]));
Q_ASSIGN U1730 ( .B(clk), .A(\g.we_clk [31044]));
Q_ASSIGN U1731 ( .B(clk), .A(\g.we_clk [31043]));
Q_ASSIGN U1732 ( .B(clk), .A(\g.we_clk [31042]));
Q_ASSIGN U1733 ( .B(clk), .A(\g.we_clk [31041]));
Q_ASSIGN U1734 ( .B(clk), .A(\g.we_clk [31040]));
Q_ASSIGN U1735 ( .B(clk), .A(\g.we_clk [31039]));
Q_ASSIGN U1736 ( .B(clk), .A(\g.we_clk [31038]));
Q_ASSIGN U1737 ( .B(clk), .A(\g.we_clk [31037]));
Q_ASSIGN U1738 ( .B(clk), .A(\g.we_clk [31036]));
Q_ASSIGN U1739 ( .B(clk), .A(\g.we_clk [31035]));
Q_ASSIGN U1740 ( .B(clk), .A(\g.we_clk [31034]));
Q_ASSIGN U1741 ( .B(clk), .A(\g.we_clk [31033]));
Q_ASSIGN U1742 ( .B(clk), .A(\g.we_clk [31032]));
Q_ASSIGN U1743 ( .B(clk), .A(\g.we_clk [31031]));
Q_ASSIGN U1744 ( .B(clk), .A(\g.we_clk [31030]));
Q_ASSIGN U1745 ( .B(clk), .A(\g.we_clk [31029]));
Q_ASSIGN U1746 ( .B(clk), .A(\g.we_clk [31028]));
Q_ASSIGN U1747 ( .B(clk), .A(\g.we_clk [31027]));
Q_ASSIGN U1748 ( .B(clk), .A(\g.we_clk [31026]));
Q_ASSIGN U1749 ( .B(clk), .A(\g.we_clk [31025]));
Q_ASSIGN U1750 ( .B(clk), .A(\g.we_clk [31024]));
Q_ASSIGN U1751 ( .B(clk), .A(\g.we_clk [31023]));
Q_ASSIGN U1752 ( .B(clk), .A(\g.we_clk [31022]));
Q_ASSIGN U1753 ( .B(clk), .A(\g.we_clk [31021]));
Q_ASSIGN U1754 ( .B(clk), .A(\g.we_clk [31020]));
Q_ASSIGN U1755 ( .B(clk), .A(\g.we_clk [31019]));
Q_ASSIGN U1756 ( .B(clk), .A(\g.we_clk [31018]));
Q_ASSIGN U1757 ( .B(clk), .A(\g.we_clk [31017]));
Q_ASSIGN U1758 ( .B(clk), .A(\g.we_clk [31016]));
Q_ASSIGN U1759 ( .B(clk), .A(\g.we_clk [31015]));
Q_ASSIGN U1760 ( .B(clk), .A(\g.we_clk [31014]));
Q_ASSIGN U1761 ( .B(clk), .A(\g.we_clk [31013]));
Q_ASSIGN U1762 ( .B(clk), .A(\g.we_clk [31012]));
Q_ASSIGN U1763 ( .B(clk), .A(\g.we_clk [31011]));
Q_ASSIGN U1764 ( .B(clk), .A(\g.we_clk [31010]));
Q_ASSIGN U1765 ( .B(clk), .A(\g.we_clk [31009]));
Q_ASSIGN U1766 ( .B(clk), .A(\g.we_clk [31008]));
Q_ASSIGN U1767 ( .B(clk), .A(\g.we_clk [31007]));
Q_ASSIGN U1768 ( .B(clk), .A(\g.we_clk [31006]));
Q_ASSIGN U1769 ( .B(clk), .A(\g.we_clk [31005]));
Q_ASSIGN U1770 ( .B(clk), .A(\g.we_clk [31004]));
Q_ASSIGN U1771 ( .B(clk), .A(\g.we_clk [31003]));
Q_ASSIGN U1772 ( .B(clk), .A(\g.we_clk [31002]));
Q_ASSIGN U1773 ( .B(clk), .A(\g.we_clk [31001]));
Q_ASSIGN U1774 ( .B(clk), .A(\g.we_clk [31000]));
Q_ASSIGN U1775 ( .B(clk), .A(\g.we_clk [30999]));
Q_ASSIGN U1776 ( .B(clk), .A(\g.we_clk [30998]));
Q_ASSIGN U1777 ( .B(clk), .A(\g.we_clk [30997]));
Q_ASSIGN U1778 ( .B(clk), .A(\g.we_clk [30996]));
Q_ASSIGN U1779 ( .B(clk), .A(\g.we_clk [30995]));
Q_ASSIGN U1780 ( .B(clk), .A(\g.we_clk [30994]));
Q_ASSIGN U1781 ( .B(clk), .A(\g.we_clk [30993]));
Q_ASSIGN U1782 ( .B(clk), .A(\g.we_clk [30992]));
Q_ASSIGN U1783 ( .B(clk), .A(\g.we_clk [30991]));
Q_ASSIGN U1784 ( .B(clk), .A(\g.we_clk [30990]));
Q_ASSIGN U1785 ( .B(clk), .A(\g.we_clk [30989]));
Q_ASSIGN U1786 ( .B(clk), .A(\g.we_clk [30988]));
Q_ASSIGN U1787 ( .B(clk), .A(\g.we_clk [30987]));
Q_ASSIGN U1788 ( .B(clk), .A(\g.we_clk [30986]));
Q_ASSIGN U1789 ( .B(clk), .A(\g.we_clk [30985]));
Q_ASSIGN U1790 ( .B(clk), .A(\g.we_clk [30984]));
Q_ASSIGN U1791 ( .B(clk), .A(\g.we_clk [30983]));
Q_ASSIGN U1792 ( .B(clk), .A(\g.we_clk [30982]));
Q_ASSIGN U1793 ( .B(clk), .A(\g.we_clk [30981]));
Q_ASSIGN U1794 ( .B(clk), .A(\g.we_clk [30980]));
Q_ASSIGN U1795 ( .B(clk), .A(\g.we_clk [30979]));
Q_ASSIGN U1796 ( .B(clk), .A(\g.we_clk [30978]));
Q_ASSIGN U1797 ( .B(clk), .A(\g.we_clk [30977]));
Q_ASSIGN U1798 ( .B(clk), .A(\g.we_clk [30976]));
Q_ASSIGN U1799 ( .B(clk), .A(\g.we_clk [30975]));
Q_ASSIGN U1800 ( .B(clk), .A(\g.we_clk [30974]));
Q_ASSIGN U1801 ( .B(clk), .A(\g.we_clk [30973]));
Q_ASSIGN U1802 ( .B(clk), .A(\g.we_clk [30972]));
Q_ASSIGN U1803 ( .B(clk), .A(\g.we_clk [30971]));
Q_ASSIGN U1804 ( .B(clk), .A(\g.we_clk [30970]));
Q_ASSIGN U1805 ( .B(clk), .A(\g.we_clk [30969]));
Q_ASSIGN U1806 ( .B(clk), .A(\g.we_clk [30968]));
Q_ASSIGN U1807 ( .B(clk), .A(\g.we_clk [30967]));
Q_ASSIGN U1808 ( .B(clk), .A(\g.we_clk [30966]));
Q_ASSIGN U1809 ( .B(clk), .A(\g.we_clk [30965]));
Q_ASSIGN U1810 ( .B(clk), .A(\g.we_clk [30964]));
Q_ASSIGN U1811 ( .B(clk), .A(\g.we_clk [30963]));
Q_ASSIGN U1812 ( .B(clk), .A(\g.we_clk [30962]));
Q_ASSIGN U1813 ( .B(clk), .A(\g.we_clk [30961]));
Q_ASSIGN U1814 ( .B(clk), .A(\g.we_clk [30960]));
Q_ASSIGN U1815 ( .B(clk), .A(\g.we_clk [30959]));
Q_ASSIGN U1816 ( .B(clk), .A(\g.we_clk [30958]));
Q_ASSIGN U1817 ( .B(clk), .A(\g.we_clk [30957]));
Q_ASSIGN U1818 ( .B(clk), .A(\g.we_clk [30956]));
Q_ASSIGN U1819 ( .B(clk), .A(\g.we_clk [30955]));
Q_ASSIGN U1820 ( .B(clk), .A(\g.we_clk [30954]));
Q_ASSIGN U1821 ( .B(clk), .A(\g.we_clk [30953]));
Q_ASSIGN U1822 ( .B(clk), .A(\g.we_clk [30952]));
Q_ASSIGN U1823 ( .B(clk), .A(\g.we_clk [30951]));
Q_ASSIGN U1824 ( .B(clk), .A(\g.we_clk [30950]));
Q_ASSIGN U1825 ( .B(clk), .A(\g.we_clk [30949]));
Q_ASSIGN U1826 ( .B(clk), .A(\g.we_clk [30948]));
Q_ASSIGN U1827 ( .B(clk), .A(\g.we_clk [30947]));
Q_ASSIGN U1828 ( .B(clk), .A(\g.we_clk [30946]));
Q_ASSIGN U1829 ( .B(clk), .A(\g.we_clk [30945]));
Q_ASSIGN U1830 ( .B(clk), .A(\g.we_clk [30944]));
Q_ASSIGN U1831 ( .B(clk), .A(\g.we_clk [30943]));
Q_ASSIGN U1832 ( .B(clk), .A(\g.we_clk [30942]));
Q_ASSIGN U1833 ( .B(clk), .A(\g.we_clk [30941]));
Q_ASSIGN U1834 ( .B(clk), .A(\g.we_clk [30940]));
Q_ASSIGN U1835 ( .B(clk), .A(\g.we_clk [30939]));
Q_ASSIGN U1836 ( .B(clk), .A(\g.we_clk [30938]));
Q_ASSIGN U1837 ( .B(clk), .A(\g.we_clk [30937]));
Q_ASSIGN U1838 ( .B(clk), .A(\g.we_clk [30936]));
Q_ASSIGN U1839 ( .B(clk), .A(\g.we_clk [30935]));
Q_ASSIGN U1840 ( .B(clk), .A(\g.we_clk [30934]));
Q_ASSIGN U1841 ( .B(clk), .A(\g.we_clk [30933]));
Q_ASSIGN U1842 ( .B(clk), .A(\g.we_clk [30932]));
Q_ASSIGN U1843 ( .B(clk), .A(\g.we_clk [30931]));
Q_ASSIGN U1844 ( .B(clk), .A(\g.we_clk [30930]));
Q_ASSIGN U1845 ( .B(clk), .A(\g.we_clk [30929]));
Q_ASSIGN U1846 ( .B(clk), .A(\g.we_clk [30928]));
Q_ASSIGN U1847 ( .B(clk), .A(\g.we_clk [30927]));
Q_ASSIGN U1848 ( .B(clk), .A(\g.we_clk [30926]));
Q_ASSIGN U1849 ( .B(clk), .A(\g.we_clk [30925]));
Q_ASSIGN U1850 ( .B(clk), .A(\g.we_clk [30924]));
Q_ASSIGN U1851 ( .B(clk), .A(\g.we_clk [30923]));
Q_ASSIGN U1852 ( .B(clk), .A(\g.we_clk [30922]));
Q_ASSIGN U1853 ( .B(clk), .A(\g.we_clk [30921]));
Q_ASSIGN U1854 ( .B(clk), .A(\g.we_clk [30920]));
Q_ASSIGN U1855 ( .B(clk), .A(\g.we_clk [30919]));
Q_ASSIGN U1856 ( .B(clk), .A(\g.we_clk [30918]));
Q_ASSIGN U1857 ( .B(clk), .A(\g.we_clk [30917]));
Q_ASSIGN U1858 ( .B(clk), .A(\g.we_clk [30916]));
Q_ASSIGN U1859 ( .B(clk), .A(\g.we_clk [30915]));
Q_ASSIGN U1860 ( .B(clk), .A(\g.we_clk [30914]));
Q_ASSIGN U1861 ( .B(clk), .A(\g.we_clk [30913]));
Q_ASSIGN U1862 ( .B(clk), .A(\g.we_clk [30912]));
Q_ASSIGN U1863 ( .B(clk), .A(\g.we_clk [30911]));
Q_ASSIGN U1864 ( .B(clk), .A(\g.we_clk [30910]));
Q_ASSIGN U1865 ( .B(clk), .A(\g.we_clk [30909]));
Q_ASSIGN U1866 ( .B(clk), .A(\g.we_clk [30908]));
Q_ASSIGN U1867 ( .B(clk), .A(\g.we_clk [30907]));
Q_ASSIGN U1868 ( .B(clk), .A(\g.we_clk [30906]));
Q_ASSIGN U1869 ( .B(clk), .A(\g.we_clk [30905]));
Q_ASSIGN U1870 ( .B(clk), .A(\g.we_clk [30904]));
Q_ASSIGN U1871 ( .B(clk), .A(\g.we_clk [30903]));
Q_ASSIGN U1872 ( .B(clk), .A(\g.we_clk [30902]));
Q_ASSIGN U1873 ( .B(clk), .A(\g.we_clk [30901]));
Q_ASSIGN U1874 ( .B(clk), .A(\g.we_clk [30900]));
Q_ASSIGN U1875 ( .B(clk), .A(\g.we_clk [30899]));
Q_ASSIGN U1876 ( .B(clk), .A(\g.we_clk [30898]));
Q_ASSIGN U1877 ( .B(clk), .A(\g.we_clk [30897]));
Q_ASSIGN U1878 ( .B(clk), .A(\g.we_clk [30896]));
Q_ASSIGN U1879 ( .B(clk), .A(\g.we_clk [30895]));
Q_ASSIGN U1880 ( .B(clk), .A(\g.we_clk [30894]));
Q_ASSIGN U1881 ( .B(clk), .A(\g.we_clk [30893]));
Q_ASSIGN U1882 ( .B(clk), .A(\g.we_clk [30892]));
Q_ASSIGN U1883 ( .B(clk), .A(\g.we_clk [30891]));
Q_ASSIGN U1884 ( .B(clk), .A(\g.we_clk [30890]));
Q_ASSIGN U1885 ( .B(clk), .A(\g.we_clk [30889]));
Q_ASSIGN U1886 ( .B(clk), .A(\g.we_clk [30888]));
Q_ASSIGN U1887 ( .B(clk), .A(\g.we_clk [30887]));
Q_ASSIGN U1888 ( .B(clk), .A(\g.we_clk [30886]));
Q_ASSIGN U1889 ( .B(clk), .A(\g.we_clk [30885]));
Q_ASSIGN U1890 ( .B(clk), .A(\g.we_clk [30884]));
Q_ASSIGN U1891 ( .B(clk), .A(\g.we_clk [30883]));
Q_ASSIGN U1892 ( .B(clk), .A(\g.we_clk [30882]));
Q_ASSIGN U1893 ( .B(clk), .A(\g.we_clk [30881]));
Q_ASSIGN U1894 ( .B(clk), .A(\g.we_clk [30880]));
Q_ASSIGN U1895 ( .B(clk), .A(\g.we_clk [30879]));
Q_ASSIGN U1896 ( .B(clk), .A(\g.we_clk [30878]));
Q_ASSIGN U1897 ( .B(clk), .A(\g.we_clk [30877]));
Q_ASSIGN U1898 ( .B(clk), .A(\g.we_clk [30876]));
Q_ASSIGN U1899 ( .B(clk), .A(\g.we_clk [30875]));
Q_ASSIGN U1900 ( .B(clk), .A(\g.we_clk [30874]));
Q_ASSIGN U1901 ( .B(clk), .A(\g.we_clk [30873]));
Q_ASSIGN U1902 ( .B(clk), .A(\g.we_clk [30872]));
Q_ASSIGN U1903 ( .B(clk), .A(\g.we_clk [30871]));
Q_ASSIGN U1904 ( .B(clk), .A(\g.we_clk [30870]));
Q_ASSIGN U1905 ( .B(clk), .A(\g.we_clk [30869]));
Q_ASSIGN U1906 ( .B(clk), .A(\g.we_clk [30868]));
Q_ASSIGN U1907 ( .B(clk), .A(\g.we_clk [30867]));
Q_ASSIGN U1908 ( .B(clk), .A(\g.we_clk [30866]));
Q_ASSIGN U1909 ( .B(clk), .A(\g.we_clk [30865]));
Q_ASSIGN U1910 ( .B(clk), .A(\g.we_clk [30864]));
Q_ASSIGN U1911 ( .B(clk), .A(\g.we_clk [30863]));
Q_ASSIGN U1912 ( .B(clk), .A(\g.we_clk [30862]));
Q_ASSIGN U1913 ( .B(clk), .A(\g.we_clk [30861]));
Q_ASSIGN U1914 ( .B(clk), .A(\g.we_clk [30860]));
Q_ASSIGN U1915 ( .B(clk), .A(\g.we_clk [30859]));
Q_ASSIGN U1916 ( .B(clk), .A(\g.we_clk [30858]));
Q_ASSIGN U1917 ( .B(clk), .A(\g.we_clk [30857]));
Q_ASSIGN U1918 ( .B(clk), .A(\g.we_clk [30856]));
Q_ASSIGN U1919 ( .B(clk), .A(\g.we_clk [30855]));
Q_ASSIGN U1920 ( .B(clk), .A(\g.we_clk [30854]));
Q_ASSIGN U1921 ( .B(clk), .A(\g.we_clk [30853]));
Q_ASSIGN U1922 ( .B(clk), .A(\g.we_clk [30852]));
Q_ASSIGN U1923 ( .B(clk), .A(\g.we_clk [30851]));
Q_ASSIGN U1924 ( .B(clk), .A(\g.we_clk [30850]));
Q_ASSIGN U1925 ( .B(clk), .A(\g.we_clk [30849]));
Q_ASSIGN U1926 ( .B(clk), .A(\g.we_clk [30848]));
Q_ASSIGN U1927 ( .B(clk), .A(\g.we_clk [30847]));
Q_ASSIGN U1928 ( .B(clk), .A(\g.we_clk [30846]));
Q_ASSIGN U1929 ( .B(clk), .A(\g.we_clk [30845]));
Q_ASSIGN U1930 ( .B(clk), .A(\g.we_clk [30844]));
Q_ASSIGN U1931 ( .B(clk), .A(\g.we_clk [30843]));
Q_ASSIGN U1932 ( .B(clk), .A(\g.we_clk [30842]));
Q_ASSIGN U1933 ( .B(clk), .A(\g.we_clk [30841]));
Q_ASSIGN U1934 ( .B(clk), .A(\g.we_clk [30840]));
Q_ASSIGN U1935 ( .B(clk), .A(\g.we_clk [30839]));
Q_ASSIGN U1936 ( .B(clk), .A(\g.we_clk [30838]));
Q_ASSIGN U1937 ( .B(clk), .A(\g.we_clk [30837]));
Q_ASSIGN U1938 ( .B(clk), .A(\g.we_clk [30836]));
Q_ASSIGN U1939 ( .B(clk), .A(\g.we_clk [30835]));
Q_ASSIGN U1940 ( .B(clk), .A(\g.we_clk [30834]));
Q_ASSIGN U1941 ( .B(clk), .A(\g.we_clk [30833]));
Q_ASSIGN U1942 ( .B(clk), .A(\g.we_clk [30832]));
Q_ASSIGN U1943 ( .B(clk), .A(\g.we_clk [30831]));
Q_ASSIGN U1944 ( .B(clk), .A(\g.we_clk [30830]));
Q_ASSIGN U1945 ( .B(clk), .A(\g.we_clk [30829]));
Q_ASSIGN U1946 ( .B(clk), .A(\g.we_clk [30828]));
Q_ASSIGN U1947 ( .B(clk), .A(\g.we_clk [30827]));
Q_ASSIGN U1948 ( .B(clk), .A(\g.we_clk [30826]));
Q_ASSIGN U1949 ( .B(clk), .A(\g.we_clk [30825]));
Q_ASSIGN U1950 ( .B(clk), .A(\g.we_clk [30824]));
Q_ASSIGN U1951 ( .B(clk), .A(\g.we_clk [30823]));
Q_ASSIGN U1952 ( .B(clk), .A(\g.we_clk [30822]));
Q_ASSIGN U1953 ( .B(clk), .A(\g.we_clk [30821]));
Q_ASSIGN U1954 ( .B(clk), .A(\g.we_clk [30820]));
Q_ASSIGN U1955 ( .B(clk), .A(\g.we_clk [30819]));
Q_ASSIGN U1956 ( .B(clk), .A(\g.we_clk [30818]));
Q_ASSIGN U1957 ( .B(clk), .A(\g.we_clk [30817]));
Q_ASSIGN U1958 ( .B(clk), .A(\g.we_clk [30816]));
Q_ASSIGN U1959 ( .B(clk), .A(\g.we_clk [30815]));
Q_ASSIGN U1960 ( .B(clk), .A(\g.we_clk [30814]));
Q_ASSIGN U1961 ( .B(clk), .A(\g.we_clk [30813]));
Q_ASSIGN U1962 ( .B(clk), .A(\g.we_clk [30812]));
Q_ASSIGN U1963 ( .B(clk), .A(\g.we_clk [30811]));
Q_ASSIGN U1964 ( .B(clk), .A(\g.we_clk [30810]));
Q_ASSIGN U1965 ( .B(clk), .A(\g.we_clk [30809]));
Q_ASSIGN U1966 ( .B(clk), .A(\g.we_clk [30808]));
Q_ASSIGN U1967 ( .B(clk), .A(\g.we_clk [30807]));
Q_ASSIGN U1968 ( .B(clk), .A(\g.we_clk [30806]));
Q_ASSIGN U1969 ( .B(clk), .A(\g.we_clk [30805]));
Q_ASSIGN U1970 ( .B(clk), .A(\g.we_clk [30804]));
Q_ASSIGN U1971 ( .B(clk), .A(\g.we_clk [30803]));
Q_ASSIGN U1972 ( .B(clk), .A(\g.we_clk [30802]));
Q_ASSIGN U1973 ( .B(clk), .A(\g.we_clk [30801]));
Q_ASSIGN U1974 ( .B(clk), .A(\g.we_clk [30800]));
Q_ASSIGN U1975 ( .B(clk), .A(\g.we_clk [30799]));
Q_ASSIGN U1976 ( .B(clk), .A(\g.we_clk [30798]));
Q_ASSIGN U1977 ( .B(clk), .A(\g.we_clk [30797]));
Q_ASSIGN U1978 ( .B(clk), .A(\g.we_clk [30796]));
Q_ASSIGN U1979 ( .B(clk), .A(\g.we_clk [30795]));
Q_ASSIGN U1980 ( .B(clk), .A(\g.we_clk [30794]));
Q_ASSIGN U1981 ( .B(clk), .A(\g.we_clk [30793]));
Q_ASSIGN U1982 ( .B(clk), .A(\g.we_clk [30792]));
Q_ASSIGN U1983 ( .B(clk), .A(\g.we_clk [30791]));
Q_ASSIGN U1984 ( .B(clk), .A(\g.we_clk [30790]));
Q_ASSIGN U1985 ( .B(clk), .A(\g.we_clk [30789]));
Q_ASSIGN U1986 ( .B(clk), .A(\g.we_clk [30788]));
Q_ASSIGN U1987 ( .B(clk), .A(\g.we_clk [30787]));
Q_ASSIGN U1988 ( .B(clk), .A(\g.we_clk [30786]));
Q_ASSIGN U1989 ( .B(clk), .A(\g.we_clk [30785]));
Q_ASSIGN U1990 ( .B(clk), .A(\g.we_clk [30784]));
Q_ASSIGN U1991 ( .B(clk), .A(\g.we_clk [30783]));
Q_ASSIGN U1992 ( .B(clk), .A(\g.we_clk [30782]));
Q_ASSIGN U1993 ( .B(clk), .A(\g.we_clk [30781]));
Q_ASSIGN U1994 ( .B(clk), .A(\g.we_clk [30780]));
Q_ASSIGN U1995 ( .B(clk), .A(\g.we_clk [30779]));
Q_ASSIGN U1996 ( .B(clk), .A(\g.we_clk [30778]));
Q_ASSIGN U1997 ( .B(clk), .A(\g.we_clk [30777]));
Q_ASSIGN U1998 ( .B(clk), .A(\g.we_clk [30776]));
Q_ASSIGN U1999 ( .B(clk), .A(\g.we_clk [30775]));
Q_ASSIGN U2000 ( .B(clk), .A(\g.we_clk [30774]));
Q_ASSIGN U2001 ( .B(clk), .A(\g.we_clk [30773]));
Q_ASSIGN U2002 ( .B(clk), .A(\g.we_clk [30772]));
Q_ASSIGN U2003 ( .B(clk), .A(\g.we_clk [30771]));
Q_ASSIGN U2004 ( .B(clk), .A(\g.we_clk [30770]));
Q_ASSIGN U2005 ( .B(clk), .A(\g.we_clk [30769]));
Q_ASSIGN U2006 ( .B(clk), .A(\g.we_clk [30768]));
Q_ASSIGN U2007 ( .B(clk), .A(\g.we_clk [30767]));
Q_ASSIGN U2008 ( .B(clk), .A(\g.we_clk [30766]));
Q_ASSIGN U2009 ( .B(clk), .A(\g.we_clk [30765]));
Q_ASSIGN U2010 ( .B(clk), .A(\g.we_clk [30764]));
Q_ASSIGN U2011 ( .B(clk), .A(\g.we_clk [30763]));
Q_ASSIGN U2012 ( .B(clk), .A(\g.we_clk [30762]));
Q_ASSIGN U2013 ( .B(clk), .A(\g.we_clk [30761]));
Q_ASSIGN U2014 ( .B(clk), .A(\g.we_clk [30760]));
Q_ASSIGN U2015 ( .B(clk), .A(\g.we_clk [30759]));
Q_ASSIGN U2016 ( .B(clk), .A(\g.we_clk [30758]));
Q_ASSIGN U2017 ( .B(clk), .A(\g.we_clk [30757]));
Q_ASSIGN U2018 ( .B(clk), .A(\g.we_clk [30756]));
Q_ASSIGN U2019 ( .B(clk), .A(\g.we_clk [30755]));
Q_ASSIGN U2020 ( .B(clk), .A(\g.we_clk [30754]));
Q_ASSIGN U2021 ( .B(clk), .A(\g.we_clk [30753]));
Q_ASSIGN U2022 ( .B(clk), .A(\g.we_clk [30752]));
Q_ASSIGN U2023 ( .B(clk), .A(\g.we_clk [30751]));
Q_ASSIGN U2024 ( .B(clk), .A(\g.we_clk [30750]));
Q_ASSIGN U2025 ( .B(clk), .A(\g.we_clk [30749]));
Q_ASSIGN U2026 ( .B(clk), .A(\g.we_clk [30748]));
Q_ASSIGN U2027 ( .B(clk), .A(\g.we_clk [30747]));
Q_ASSIGN U2028 ( .B(clk), .A(\g.we_clk [30746]));
Q_ASSIGN U2029 ( .B(clk), .A(\g.we_clk [30745]));
Q_ASSIGN U2030 ( .B(clk), .A(\g.we_clk [30744]));
Q_ASSIGN U2031 ( .B(clk), .A(\g.we_clk [30743]));
Q_ASSIGN U2032 ( .B(clk), .A(\g.we_clk [30742]));
Q_ASSIGN U2033 ( .B(clk), .A(\g.we_clk [30741]));
Q_ASSIGN U2034 ( .B(clk), .A(\g.we_clk [30740]));
Q_ASSIGN U2035 ( .B(clk), .A(\g.we_clk [30739]));
Q_ASSIGN U2036 ( .B(clk), .A(\g.we_clk [30738]));
Q_ASSIGN U2037 ( .B(clk), .A(\g.we_clk [30737]));
Q_ASSIGN U2038 ( .B(clk), .A(\g.we_clk [30736]));
Q_ASSIGN U2039 ( .B(clk), .A(\g.we_clk [30735]));
Q_ASSIGN U2040 ( .B(clk), .A(\g.we_clk [30734]));
Q_ASSIGN U2041 ( .B(clk), .A(\g.we_clk [30733]));
Q_ASSIGN U2042 ( .B(clk), .A(\g.we_clk [30732]));
Q_ASSIGN U2043 ( .B(clk), .A(\g.we_clk [30731]));
Q_ASSIGN U2044 ( .B(clk), .A(\g.we_clk [30730]));
Q_ASSIGN U2045 ( .B(clk), .A(\g.we_clk [30729]));
Q_ASSIGN U2046 ( .B(clk), .A(\g.we_clk [30728]));
Q_ASSIGN U2047 ( .B(clk), .A(\g.we_clk [30727]));
Q_ASSIGN U2048 ( .B(clk), .A(\g.we_clk [30726]));
Q_ASSIGN U2049 ( .B(clk), .A(\g.we_clk [30725]));
Q_ASSIGN U2050 ( .B(clk), .A(\g.we_clk [30724]));
Q_ASSIGN U2051 ( .B(clk), .A(\g.we_clk [30723]));
Q_ASSIGN U2052 ( .B(clk), .A(\g.we_clk [30722]));
Q_ASSIGN U2053 ( .B(clk), .A(\g.we_clk [30721]));
Q_ASSIGN U2054 ( .B(clk), .A(\g.we_clk [30720]));
Q_ASSIGN U2055 ( .B(clk), .A(\g.we_clk [30719]));
Q_ASSIGN U2056 ( .B(clk), .A(\g.we_clk [30718]));
Q_ASSIGN U2057 ( .B(clk), .A(\g.we_clk [30717]));
Q_ASSIGN U2058 ( .B(clk), .A(\g.we_clk [30716]));
Q_ASSIGN U2059 ( .B(clk), .A(\g.we_clk [30715]));
Q_ASSIGN U2060 ( .B(clk), .A(\g.we_clk [30714]));
Q_ASSIGN U2061 ( .B(clk), .A(\g.we_clk [30713]));
Q_ASSIGN U2062 ( .B(clk), .A(\g.we_clk [30712]));
Q_ASSIGN U2063 ( .B(clk), .A(\g.we_clk [30711]));
Q_ASSIGN U2064 ( .B(clk), .A(\g.we_clk [30710]));
Q_ASSIGN U2065 ( .B(clk), .A(\g.we_clk [30709]));
Q_ASSIGN U2066 ( .B(clk), .A(\g.we_clk [30708]));
Q_ASSIGN U2067 ( .B(clk), .A(\g.we_clk [30707]));
Q_ASSIGN U2068 ( .B(clk), .A(\g.we_clk [30706]));
Q_ASSIGN U2069 ( .B(clk), .A(\g.we_clk [30705]));
Q_ASSIGN U2070 ( .B(clk), .A(\g.we_clk [30704]));
Q_ASSIGN U2071 ( .B(clk), .A(\g.we_clk [30703]));
Q_ASSIGN U2072 ( .B(clk), .A(\g.we_clk [30702]));
Q_ASSIGN U2073 ( .B(clk), .A(\g.we_clk [30701]));
Q_ASSIGN U2074 ( .B(clk), .A(\g.we_clk [30700]));
Q_ASSIGN U2075 ( .B(clk), .A(\g.we_clk [30699]));
Q_ASSIGN U2076 ( .B(clk), .A(\g.we_clk [30698]));
Q_ASSIGN U2077 ( .B(clk), .A(\g.we_clk [30697]));
Q_ASSIGN U2078 ( .B(clk), .A(\g.we_clk [30696]));
Q_ASSIGN U2079 ( .B(clk), .A(\g.we_clk [30695]));
Q_ASSIGN U2080 ( .B(clk), .A(\g.we_clk [30694]));
Q_ASSIGN U2081 ( .B(clk), .A(\g.we_clk [30693]));
Q_ASSIGN U2082 ( .B(clk), .A(\g.we_clk [30692]));
Q_ASSIGN U2083 ( .B(clk), .A(\g.we_clk [30691]));
Q_ASSIGN U2084 ( .B(clk), .A(\g.we_clk [30690]));
Q_ASSIGN U2085 ( .B(clk), .A(\g.we_clk [30689]));
Q_ASSIGN U2086 ( .B(clk), .A(\g.we_clk [30688]));
Q_ASSIGN U2087 ( .B(clk), .A(\g.we_clk [30687]));
Q_ASSIGN U2088 ( .B(clk), .A(\g.we_clk [30686]));
Q_ASSIGN U2089 ( .B(clk), .A(\g.we_clk [30685]));
Q_ASSIGN U2090 ( .B(clk), .A(\g.we_clk [30684]));
Q_ASSIGN U2091 ( .B(clk), .A(\g.we_clk [30683]));
Q_ASSIGN U2092 ( .B(clk), .A(\g.we_clk [30682]));
Q_ASSIGN U2093 ( .B(clk), .A(\g.we_clk [30681]));
Q_ASSIGN U2094 ( .B(clk), .A(\g.we_clk [30680]));
Q_ASSIGN U2095 ( .B(clk), .A(\g.we_clk [30679]));
Q_ASSIGN U2096 ( .B(clk), .A(\g.we_clk [30678]));
Q_ASSIGN U2097 ( .B(clk), .A(\g.we_clk [30677]));
Q_ASSIGN U2098 ( .B(clk), .A(\g.we_clk [30676]));
Q_ASSIGN U2099 ( .B(clk), .A(\g.we_clk [30675]));
Q_ASSIGN U2100 ( .B(clk), .A(\g.we_clk [30674]));
Q_ASSIGN U2101 ( .B(clk), .A(\g.we_clk [30673]));
Q_ASSIGN U2102 ( .B(clk), .A(\g.we_clk [30672]));
Q_ASSIGN U2103 ( .B(clk), .A(\g.we_clk [30671]));
Q_ASSIGN U2104 ( .B(clk), .A(\g.we_clk [30670]));
Q_ASSIGN U2105 ( .B(clk), .A(\g.we_clk [30669]));
Q_ASSIGN U2106 ( .B(clk), .A(\g.we_clk [30668]));
Q_ASSIGN U2107 ( .B(clk), .A(\g.we_clk [30667]));
Q_ASSIGN U2108 ( .B(clk), .A(\g.we_clk [30666]));
Q_ASSIGN U2109 ( .B(clk), .A(\g.we_clk [30665]));
Q_ASSIGN U2110 ( .B(clk), .A(\g.we_clk [30664]));
Q_ASSIGN U2111 ( .B(clk), .A(\g.we_clk [30663]));
Q_ASSIGN U2112 ( .B(clk), .A(\g.we_clk [30662]));
Q_ASSIGN U2113 ( .B(clk), .A(\g.we_clk [30661]));
Q_ASSIGN U2114 ( .B(clk), .A(\g.we_clk [30660]));
Q_ASSIGN U2115 ( .B(clk), .A(\g.we_clk [30659]));
Q_ASSIGN U2116 ( .B(clk), .A(\g.we_clk [30658]));
Q_ASSIGN U2117 ( .B(clk), .A(\g.we_clk [30657]));
Q_ASSIGN U2118 ( .B(clk), .A(\g.we_clk [30656]));
Q_ASSIGN U2119 ( .B(clk), .A(\g.we_clk [30655]));
Q_ASSIGN U2120 ( .B(clk), .A(\g.we_clk [30654]));
Q_ASSIGN U2121 ( .B(clk), .A(\g.we_clk [30653]));
Q_ASSIGN U2122 ( .B(clk), .A(\g.we_clk [30652]));
Q_ASSIGN U2123 ( .B(clk), .A(\g.we_clk [30651]));
Q_ASSIGN U2124 ( .B(clk), .A(\g.we_clk [30650]));
Q_ASSIGN U2125 ( .B(clk), .A(\g.we_clk [30649]));
Q_ASSIGN U2126 ( .B(clk), .A(\g.we_clk [30648]));
Q_ASSIGN U2127 ( .B(clk), .A(\g.we_clk [30647]));
Q_ASSIGN U2128 ( .B(clk), .A(\g.we_clk [30646]));
Q_ASSIGN U2129 ( .B(clk), .A(\g.we_clk [30645]));
Q_ASSIGN U2130 ( .B(clk), .A(\g.we_clk [30644]));
Q_ASSIGN U2131 ( .B(clk), .A(\g.we_clk [30643]));
Q_ASSIGN U2132 ( .B(clk), .A(\g.we_clk [30642]));
Q_ASSIGN U2133 ( .B(clk), .A(\g.we_clk [30641]));
Q_ASSIGN U2134 ( .B(clk), .A(\g.we_clk [30640]));
Q_ASSIGN U2135 ( .B(clk), .A(\g.we_clk [30639]));
Q_ASSIGN U2136 ( .B(clk), .A(\g.we_clk [30638]));
Q_ASSIGN U2137 ( .B(clk), .A(\g.we_clk [30637]));
Q_ASSIGN U2138 ( .B(clk), .A(\g.we_clk [30636]));
Q_ASSIGN U2139 ( .B(clk), .A(\g.we_clk [30635]));
Q_ASSIGN U2140 ( .B(clk), .A(\g.we_clk [30634]));
Q_ASSIGN U2141 ( .B(clk), .A(\g.we_clk [30633]));
Q_ASSIGN U2142 ( .B(clk), .A(\g.we_clk [30632]));
Q_ASSIGN U2143 ( .B(clk), .A(\g.we_clk [30631]));
Q_ASSIGN U2144 ( .B(clk), .A(\g.we_clk [30630]));
Q_ASSIGN U2145 ( .B(clk), .A(\g.we_clk [30629]));
Q_ASSIGN U2146 ( .B(clk), .A(\g.we_clk [30628]));
Q_ASSIGN U2147 ( .B(clk), .A(\g.we_clk [30627]));
Q_ASSIGN U2148 ( .B(clk), .A(\g.we_clk [30626]));
Q_ASSIGN U2149 ( .B(clk), .A(\g.we_clk [30625]));
Q_ASSIGN U2150 ( .B(clk), .A(\g.we_clk [30624]));
Q_ASSIGN U2151 ( .B(clk), .A(\g.we_clk [30623]));
Q_ASSIGN U2152 ( .B(clk), .A(\g.we_clk [30622]));
Q_ASSIGN U2153 ( .B(clk), .A(\g.we_clk [30621]));
Q_ASSIGN U2154 ( .B(clk), .A(\g.we_clk [30620]));
Q_ASSIGN U2155 ( .B(clk), .A(\g.we_clk [30619]));
Q_ASSIGN U2156 ( .B(clk), .A(\g.we_clk [30618]));
Q_ASSIGN U2157 ( .B(clk), .A(\g.we_clk [30617]));
Q_ASSIGN U2158 ( .B(clk), .A(\g.we_clk [30616]));
Q_ASSIGN U2159 ( .B(clk), .A(\g.we_clk [30615]));
Q_ASSIGN U2160 ( .B(clk), .A(\g.we_clk [30614]));
Q_ASSIGN U2161 ( .B(clk), .A(\g.we_clk [30613]));
Q_ASSIGN U2162 ( .B(clk), .A(\g.we_clk [30612]));
Q_ASSIGN U2163 ( .B(clk), .A(\g.we_clk [30611]));
Q_ASSIGN U2164 ( .B(clk), .A(\g.we_clk [30610]));
Q_ASSIGN U2165 ( .B(clk), .A(\g.we_clk [30609]));
Q_ASSIGN U2166 ( .B(clk), .A(\g.we_clk [30608]));
Q_ASSIGN U2167 ( .B(clk), .A(\g.we_clk [30607]));
Q_ASSIGN U2168 ( .B(clk), .A(\g.we_clk [30606]));
Q_ASSIGN U2169 ( .B(clk), .A(\g.we_clk [30605]));
Q_ASSIGN U2170 ( .B(clk), .A(\g.we_clk [30604]));
Q_ASSIGN U2171 ( .B(clk), .A(\g.we_clk [30603]));
Q_ASSIGN U2172 ( .B(clk), .A(\g.we_clk [30602]));
Q_ASSIGN U2173 ( .B(clk), .A(\g.we_clk [30601]));
Q_ASSIGN U2174 ( .B(clk), .A(\g.we_clk [30600]));
Q_ASSIGN U2175 ( .B(clk), .A(\g.we_clk [30599]));
Q_ASSIGN U2176 ( .B(clk), .A(\g.we_clk [30598]));
Q_ASSIGN U2177 ( .B(clk), .A(\g.we_clk [30597]));
Q_ASSIGN U2178 ( .B(clk), .A(\g.we_clk [30596]));
Q_ASSIGN U2179 ( .B(clk), .A(\g.we_clk [30595]));
Q_ASSIGN U2180 ( .B(clk), .A(\g.we_clk [30594]));
Q_ASSIGN U2181 ( .B(clk), .A(\g.we_clk [30593]));
Q_ASSIGN U2182 ( .B(clk), .A(\g.we_clk [30592]));
Q_ASSIGN U2183 ( .B(clk), .A(\g.we_clk [30591]));
Q_ASSIGN U2184 ( .B(clk), .A(\g.we_clk [30590]));
Q_ASSIGN U2185 ( .B(clk), .A(\g.we_clk [30589]));
Q_ASSIGN U2186 ( .B(clk), .A(\g.we_clk [30588]));
Q_ASSIGN U2187 ( .B(clk), .A(\g.we_clk [30587]));
Q_ASSIGN U2188 ( .B(clk), .A(\g.we_clk [30586]));
Q_ASSIGN U2189 ( .B(clk), .A(\g.we_clk [30585]));
Q_ASSIGN U2190 ( .B(clk), .A(\g.we_clk [30584]));
Q_ASSIGN U2191 ( .B(clk), .A(\g.we_clk [30583]));
Q_ASSIGN U2192 ( .B(clk), .A(\g.we_clk [30582]));
Q_ASSIGN U2193 ( .B(clk), .A(\g.we_clk [30581]));
Q_ASSIGN U2194 ( .B(clk), .A(\g.we_clk [30580]));
Q_ASSIGN U2195 ( .B(clk), .A(\g.we_clk [30579]));
Q_ASSIGN U2196 ( .B(clk), .A(\g.we_clk [30578]));
Q_ASSIGN U2197 ( .B(clk), .A(\g.we_clk [30577]));
Q_ASSIGN U2198 ( .B(clk), .A(\g.we_clk [30576]));
Q_ASSIGN U2199 ( .B(clk), .A(\g.we_clk [30575]));
Q_ASSIGN U2200 ( .B(clk), .A(\g.we_clk [30574]));
Q_ASSIGN U2201 ( .B(clk), .A(\g.we_clk [30573]));
Q_ASSIGN U2202 ( .B(clk), .A(\g.we_clk [30572]));
Q_ASSIGN U2203 ( .B(clk), .A(\g.we_clk [30571]));
Q_ASSIGN U2204 ( .B(clk), .A(\g.we_clk [30570]));
Q_ASSIGN U2205 ( .B(clk), .A(\g.we_clk [30569]));
Q_ASSIGN U2206 ( .B(clk), .A(\g.we_clk [30568]));
Q_ASSIGN U2207 ( .B(clk), .A(\g.we_clk [30567]));
Q_ASSIGN U2208 ( .B(clk), .A(\g.we_clk [30566]));
Q_ASSIGN U2209 ( .B(clk), .A(\g.we_clk [30565]));
Q_ASSIGN U2210 ( .B(clk), .A(\g.we_clk [30564]));
Q_ASSIGN U2211 ( .B(clk), .A(\g.we_clk [30563]));
Q_ASSIGN U2212 ( .B(clk), .A(\g.we_clk [30562]));
Q_ASSIGN U2213 ( .B(clk), .A(\g.we_clk [30561]));
Q_ASSIGN U2214 ( .B(clk), .A(\g.we_clk [30560]));
Q_ASSIGN U2215 ( .B(clk), .A(\g.we_clk [30559]));
Q_ASSIGN U2216 ( .B(clk), .A(\g.we_clk [30558]));
Q_ASSIGN U2217 ( .B(clk), .A(\g.we_clk [30557]));
Q_ASSIGN U2218 ( .B(clk), .A(\g.we_clk [30556]));
Q_ASSIGN U2219 ( .B(clk), .A(\g.we_clk [30555]));
Q_ASSIGN U2220 ( .B(clk), .A(\g.we_clk [30554]));
Q_ASSIGN U2221 ( .B(clk), .A(\g.we_clk [30553]));
Q_ASSIGN U2222 ( .B(clk), .A(\g.we_clk [30552]));
Q_ASSIGN U2223 ( .B(clk), .A(\g.we_clk [30551]));
Q_ASSIGN U2224 ( .B(clk), .A(\g.we_clk [30550]));
Q_ASSIGN U2225 ( .B(clk), .A(\g.we_clk [30549]));
Q_ASSIGN U2226 ( .B(clk), .A(\g.we_clk [30548]));
Q_ASSIGN U2227 ( .B(clk), .A(\g.we_clk [30547]));
Q_ASSIGN U2228 ( .B(clk), .A(\g.we_clk [30546]));
Q_ASSIGN U2229 ( .B(clk), .A(\g.we_clk [30545]));
Q_ASSIGN U2230 ( .B(clk), .A(\g.we_clk [30544]));
Q_ASSIGN U2231 ( .B(clk), .A(\g.we_clk [30543]));
Q_ASSIGN U2232 ( .B(clk), .A(\g.we_clk [30542]));
Q_ASSIGN U2233 ( .B(clk), .A(\g.we_clk [30541]));
Q_ASSIGN U2234 ( .B(clk), .A(\g.we_clk [30540]));
Q_ASSIGN U2235 ( .B(clk), .A(\g.we_clk [30539]));
Q_ASSIGN U2236 ( .B(clk), .A(\g.we_clk [30538]));
Q_ASSIGN U2237 ( .B(clk), .A(\g.we_clk [30537]));
Q_ASSIGN U2238 ( .B(clk), .A(\g.we_clk [30536]));
Q_ASSIGN U2239 ( .B(clk), .A(\g.we_clk [30535]));
Q_ASSIGN U2240 ( .B(clk), .A(\g.we_clk [30534]));
Q_ASSIGN U2241 ( .B(clk), .A(\g.we_clk [30533]));
Q_ASSIGN U2242 ( .B(clk), .A(\g.we_clk [30532]));
Q_ASSIGN U2243 ( .B(clk), .A(\g.we_clk [30531]));
Q_ASSIGN U2244 ( .B(clk), .A(\g.we_clk [30530]));
Q_ASSIGN U2245 ( .B(clk), .A(\g.we_clk [30529]));
Q_ASSIGN U2246 ( .B(clk), .A(\g.we_clk [30528]));
Q_ASSIGN U2247 ( .B(clk), .A(\g.we_clk [30527]));
Q_ASSIGN U2248 ( .B(clk), .A(\g.we_clk [30526]));
Q_ASSIGN U2249 ( .B(clk), .A(\g.we_clk [30525]));
Q_ASSIGN U2250 ( .B(clk), .A(\g.we_clk [30524]));
Q_ASSIGN U2251 ( .B(clk), .A(\g.we_clk [30523]));
Q_ASSIGN U2252 ( .B(clk), .A(\g.we_clk [30522]));
Q_ASSIGN U2253 ( .B(clk), .A(\g.we_clk [30521]));
Q_ASSIGN U2254 ( .B(clk), .A(\g.we_clk [30520]));
Q_ASSIGN U2255 ( .B(clk), .A(\g.we_clk [30519]));
Q_ASSIGN U2256 ( .B(clk), .A(\g.we_clk [30518]));
Q_ASSIGN U2257 ( .B(clk), .A(\g.we_clk [30517]));
Q_ASSIGN U2258 ( .B(clk), .A(\g.we_clk [30516]));
Q_ASSIGN U2259 ( .B(clk), .A(\g.we_clk [30515]));
Q_ASSIGN U2260 ( .B(clk), .A(\g.we_clk [30514]));
Q_ASSIGN U2261 ( .B(clk), .A(\g.we_clk [30513]));
Q_ASSIGN U2262 ( .B(clk), .A(\g.we_clk [30512]));
Q_ASSIGN U2263 ( .B(clk), .A(\g.we_clk [30511]));
Q_ASSIGN U2264 ( .B(clk), .A(\g.we_clk [30510]));
Q_ASSIGN U2265 ( .B(clk), .A(\g.we_clk [30509]));
Q_ASSIGN U2266 ( .B(clk), .A(\g.we_clk [30508]));
Q_ASSIGN U2267 ( .B(clk), .A(\g.we_clk [30507]));
Q_ASSIGN U2268 ( .B(clk), .A(\g.we_clk [30506]));
Q_ASSIGN U2269 ( .B(clk), .A(\g.we_clk [30505]));
Q_ASSIGN U2270 ( .B(clk), .A(\g.we_clk [30504]));
Q_ASSIGN U2271 ( .B(clk), .A(\g.we_clk [30503]));
Q_ASSIGN U2272 ( .B(clk), .A(\g.we_clk [30502]));
Q_ASSIGN U2273 ( .B(clk), .A(\g.we_clk [30501]));
Q_ASSIGN U2274 ( .B(clk), .A(\g.we_clk [30500]));
Q_ASSIGN U2275 ( .B(clk), .A(\g.we_clk [30499]));
Q_ASSIGN U2276 ( .B(clk), .A(\g.we_clk [30498]));
Q_ASSIGN U2277 ( .B(clk), .A(\g.we_clk [30497]));
Q_ASSIGN U2278 ( .B(clk), .A(\g.we_clk [30496]));
Q_ASSIGN U2279 ( .B(clk), .A(\g.we_clk [30495]));
Q_ASSIGN U2280 ( .B(clk), .A(\g.we_clk [30494]));
Q_ASSIGN U2281 ( .B(clk), .A(\g.we_clk [30493]));
Q_ASSIGN U2282 ( .B(clk), .A(\g.we_clk [30492]));
Q_ASSIGN U2283 ( .B(clk), .A(\g.we_clk [30491]));
Q_ASSIGN U2284 ( .B(clk), .A(\g.we_clk [30490]));
Q_ASSIGN U2285 ( .B(clk), .A(\g.we_clk [30489]));
Q_ASSIGN U2286 ( .B(clk), .A(\g.we_clk [30488]));
Q_ASSIGN U2287 ( .B(clk), .A(\g.we_clk [30487]));
Q_ASSIGN U2288 ( .B(clk), .A(\g.we_clk [30486]));
Q_ASSIGN U2289 ( .B(clk), .A(\g.we_clk [30485]));
Q_ASSIGN U2290 ( .B(clk), .A(\g.we_clk [30484]));
Q_ASSIGN U2291 ( .B(clk), .A(\g.we_clk [30483]));
Q_ASSIGN U2292 ( .B(clk), .A(\g.we_clk [30482]));
Q_ASSIGN U2293 ( .B(clk), .A(\g.we_clk [30481]));
Q_ASSIGN U2294 ( .B(clk), .A(\g.we_clk [30480]));
Q_ASSIGN U2295 ( .B(clk), .A(\g.we_clk [30479]));
Q_ASSIGN U2296 ( .B(clk), .A(\g.we_clk [30478]));
Q_ASSIGN U2297 ( .B(clk), .A(\g.we_clk [30477]));
Q_ASSIGN U2298 ( .B(clk), .A(\g.we_clk [30476]));
Q_ASSIGN U2299 ( .B(clk), .A(\g.we_clk [30475]));
Q_ASSIGN U2300 ( .B(clk), .A(\g.we_clk [30474]));
Q_ASSIGN U2301 ( .B(clk), .A(\g.we_clk [30473]));
Q_ASSIGN U2302 ( .B(clk), .A(\g.we_clk [30472]));
Q_ASSIGN U2303 ( .B(clk), .A(\g.we_clk [30471]));
Q_ASSIGN U2304 ( .B(clk), .A(\g.we_clk [30470]));
Q_ASSIGN U2305 ( .B(clk), .A(\g.we_clk [30469]));
Q_ASSIGN U2306 ( .B(clk), .A(\g.we_clk [30468]));
Q_ASSIGN U2307 ( .B(clk), .A(\g.we_clk [30467]));
Q_ASSIGN U2308 ( .B(clk), .A(\g.we_clk [30466]));
Q_ASSIGN U2309 ( .B(clk), .A(\g.we_clk [30465]));
Q_ASSIGN U2310 ( .B(clk), .A(\g.we_clk [30464]));
Q_ASSIGN U2311 ( .B(clk), .A(\g.we_clk [30463]));
Q_ASSIGN U2312 ( .B(clk), .A(\g.we_clk [30462]));
Q_ASSIGN U2313 ( .B(clk), .A(\g.we_clk [30461]));
Q_ASSIGN U2314 ( .B(clk), .A(\g.we_clk [30460]));
Q_ASSIGN U2315 ( .B(clk), .A(\g.we_clk [30459]));
Q_ASSIGN U2316 ( .B(clk), .A(\g.we_clk [30458]));
Q_ASSIGN U2317 ( .B(clk), .A(\g.we_clk [30457]));
Q_ASSIGN U2318 ( .B(clk), .A(\g.we_clk [30456]));
Q_ASSIGN U2319 ( .B(clk), .A(\g.we_clk [30455]));
Q_ASSIGN U2320 ( .B(clk), .A(\g.we_clk [30454]));
Q_ASSIGN U2321 ( .B(clk), .A(\g.we_clk [30453]));
Q_ASSIGN U2322 ( .B(clk), .A(\g.we_clk [30452]));
Q_ASSIGN U2323 ( .B(clk), .A(\g.we_clk [30451]));
Q_ASSIGN U2324 ( .B(clk), .A(\g.we_clk [30450]));
Q_ASSIGN U2325 ( .B(clk), .A(\g.we_clk [30449]));
Q_ASSIGN U2326 ( .B(clk), .A(\g.we_clk [30448]));
Q_ASSIGN U2327 ( .B(clk), .A(\g.we_clk [30447]));
Q_ASSIGN U2328 ( .B(clk), .A(\g.we_clk [30446]));
Q_ASSIGN U2329 ( .B(clk), .A(\g.we_clk [30445]));
Q_ASSIGN U2330 ( .B(clk), .A(\g.we_clk [30444]));
Q_ASSIGN U2331 ( .B(clk), .A(\g.we_clk [30443]));
Q_ASSIGN U2332 ( .B(clk), .A(\g.we_clk [30442]));
Q_ASSIGN U2333 ( .B(clk), .A(\g.we_clk [30441]));
Q_ASSIGN U2334 ( .B(clk), .A(\g.we_clk [30440]));
Q_ASSIGN U2335 ( .B(clk), .A(\g.we_clk [30439]));
Q_ASSIGN U2336 ( .B(clk), .A(\g.we_clk [30438]));
Q_ASSIGN U2337 ( .B(clk), .A(\g.we_clk [30437]));
Q_ASSIGN U2338 ( .B(clk), .A(\g.we_clk [30436]));
Q_ASSIGN U2339 ( .B(clk), .A(\g.we_clk [30435]));
Q_ASSIGN U2340 ( .B(clk), .A(\g.we_clk [30434]));
Q_ASSIGN U2341 ( .B(clk), .A(\g.we_clk [30433]));
Q_ASSIGN U2342 ( .B(clk), .A(\g.we_clk [30432]));
Q_ASSIGN U2343 ( .B(clk), .A(\g.we_clk [30431]));
Q_ASSIGN U2344 ( .B(clk), .A(\g.we_clk [30430]));
Q_ASSIGN U2345 ( .B(clk), .A(\g.we_clk [30429]));
Q_ASSIGN U2346 ( .B(clk), .A(\g.we_clk [30428]));
Q_ASSIGN U2347 ( .B(clk), .A(\g.we_clk [30427]));
Q_ASSIGN U2348 ( .B(clk), .A(\g.we_clk [30426]));
Q_ASSIGN U2349 ( .B(clk), .A(\g.we_clk [30425]));
Q_ASSIGN U2350 ( .B(clk), .A(\g.we_clk [30424]));
Q_ASSIGN U2351 ( .B(clk), .A(\g.we_clk [30423]));
Q_ASSIGN U2352 ( .B(clk), .A(\g.we_clk [30422]));
Q_ASSIGN U2353 ( .B(clk), .A(\g.we_clk [30421]));
Q_ASSIGN U2354 ( .B(clk), .A(\g.we_clk [30420]));
Q_ASSIGN U2355 ( .B(clk), .A(\g.we_clk [30419]));
Q_ASSIGN U2356 ( .B(clk), .A(\g.we_clk [30418]));
Q_ASSIGN U2357 ( .B(clk), .A(\g.we_clk [30417]));
Q_ASSIGN U2358 ( .B(clk), .A(\g.we_clk [30416]));
Q_ASSIGN U2359 ( .B(clk), .A(\g.we_clk [30415]));
Q_ASSIGN U2360 ( .B(clk), .A(\g.we_clk [30414]));
Q_ASSIGN U2361 ( .B(clk), .A(\g.we_clk [30413]));
Q_ASSIGN U2362 ( .B(clk), .A(\g.we_clk [30412]));
Q_ASSIGN U2363 ( .B(clk), .A(\g.we_clk [30411]));
Q_ASSIGN U2364 ( .B(clk), .A(\g.we_clk [30410]));
Q_ASSIGN U2365 ( .B(clk), .A(\g.we_clk [30409]));
Q_ASSIGN U2366 ( .B(clk), .A(\g.we_clk [30408]));
Q_ASSIGN U2367 ( .B(clk), .A(\g.we_clk [30407]));
Q_ASSIGN U2368 ( .B(clk), .A(\g.we_clk [30406]));
Q_ASSIGN U2369 ( .B(clk), .A(\g.we_clk [30405]));
Q_ASSIGN U2370 ( .B(clk), .A(\g.we_clk [30404]));
Q_ASSIGN U2371 ( .B(clk), .A(\g.we_clk [30403]));
Q_ASSIGN U2372 ( .B(clk), .A(\g.we_clk [30402]));
Q_ASSIGN U2373 ( .B(clk), .A(\g.we_clk [30401]));
Q_ASSIGN U2374 ( .B(clk), .A(\g.we_clk [30400]));
Q_ASSIGN U2375 ( .B(clk), .A(\g.we_clk [30399]));
Q_ASSIGN U2376 ( .B(clk), .A(\g.we_clk [30398]));
Q_ASSIGN U2377 ( .B(clk), .A(\g.we_clk [30397]));
Q_ASSIGN U2378 ( .B(clk), .A(\g.we_clk [30396]));
Q_ASSIGN U2379 ( .B(clk), .A(\g.we_clk [30395]));
Q_ASSIGN U2380 ( .B(clk), .A(\g.we_clk [30394]));
Q_ASSIGN U2381 ( .B(clk), .A(\g.we_clk [30393]));
Q_ASSIGN U2382 ( .B(clk), .A(\g.we_clk [30392]));
Q_ASSIGN U2383 ( .B(clk), .A(\g.we_clk [30391]));
Q_ASSIGN U2384 ( .B(clk), .A(\g.we_clk [30390]));
Q_ASSIGN U2385 ( .B(clk), .A(\g.we_clk [30389]));
Q_ASSIGN U2386 ( .B(clk), .A(\g.we_clk [30388]));
Q_ASSIGN U2387 ( .B(clk), .A(\g.we_clk [30387]));
Q_ASSIGN U2388 ( .B(clk), .A(\g.we_clk [30386]));
Q_ASSIGN U2389 ( .B(clk), .A(\g.we_clk [30385]));
Q_ASSIGN U2390 ( .B(clk), .A(\g.we_clk [30384]));
Q_ASSIGN U2391 ( .B(clk), .A(\g.we_clk [30383]));
Q_ASSIGN U2392 ( .B(clk), .A(\g.we_clk [30382]));
Q_ASSIGN U2393 ( .B(clk), .A(\g.we_clk [30381]));
Q_ASSIGN U2394 ( .B(clk), .A(\g.we_clk [30380]));
Q_ASSIGN U2395 ( .B(clk), .A(\g.we_clk [30379]));
Q_ASSIGN U2396 ( .B(clk), .A(\g.we_clk [30378]));
Q_ASSIGN U2397 ( .B(clk), .A(\g.we_clk [30377]));
Q_ASSIGN U2398 ( .B(clk), .A(\g.we_clk [30376]));
Q_ASSIGN U2399 ( .B(clk), .A(\g.we_clk [30375]));
Q_ASSIGN U2400 ( .B(clk), .A(\g.we_clk [30374]));
Q_ASSIGN U2401 ( .B(clk), .A(\g.we_clk [30373]));
Q_ASSIGN U2402 ( .B(clk), .A(\g.we_clk [30372]));
Q_ASSIGN U2403 ( .B(clk), .A(\g.we_clk [30371]));
Q_ASSIGN U2404 ( .B(clk), .A(\g.we_clk [30370]));
Q_ASSIGN U2405 ( .B(clk), .A(\g.we_clk [30369]));
Q_ASSIGN U2406 ( .B(clk), .A(\g.we_clk [30368]));
Q_ASSIGN U2407 ( .B(clk), .A(\g.we_clk [30367]));
Q_ASSIGN U2408 ( .B(clk), .A(\g.we_clk [30366]));
Q_ASSIGN U2409 ( .B(clk), .A(\g.we_clk [30365]));
Q_ASSIGN U2410 ( .B(clk), .A(\g.we_clk [30364]));
Q_ASSIGN U2411 ( .B(clk), .A(\g.we_clk [30363]));
Q_ASSIGN U2412 ( .B(clk), .A(\g.we_clk [30362]));
Q_ASSIGN U2413 ( .B(clk), .A(\g.we_clk [30361]));
Q_ASSIGN U2414 ( .B(clk), .A(\g.we_clk [30360]));
Q_ASSIGN U2415 ( .B(clk), .A(\g.we_clk [30359]));
Q_ASSIGN U2416 ( .B(clk), .A(\g.we_clk [30358]));
Q_ASSIGN U2417 ( .B(clk), .A(\g.we_clk [30357]));
Q_ASSIGN U2418 ( .B(clk), .A(\g.we_clk [30356]));
Q_ASSIGN U2419 ( .B(clk), .A(\g.we_clk [30355]));
Q_ASSIGN U2420 ( .B(clk), .A(\g.we_clk [30354]));
Q_ASSIGN U2421 ( .B(clk), .A(\g.we_clk [30353]));
Q_ASSIGN U2422 ( .B(clk), .A(\g.we_clk [30352]));
Q_ASSIGN U2423 ( .B(clk), .A(\g.we_clk [30351]));
Q_ASSIGN U2424 ( .B(clk), .A(\g.we_clk [30350]));
Q_ASSIGN U2425 ( .B(clk), .A(\g.we_clk [30349]));
Q_ASSIGN U2426 ( .B(clk), .A(\g.we_clk [30348]));
Q_ASSIGN U2427 ( .B(clk), .A(\g.we_clk [30347]));
Q_ASSIGN U2428 ( .B(clk), .A(\g.we_clk [30346]));
Q_ASSIGN U2429 ( .B(clk), .A(\g.we_clk [30345]));
Q_ASSIGN U2430 ( .B(clk), .A(\g.we_clk [30344]));
Q_ASSIGN U2431 ( .B(clk), .A(\g.we_clk [30343]));
Q_ASSIGN U2432 ( .B(clk), .A(\g.we_clk [30342]));
Q_ASSIGN U2433 ( .B(clk), .A(\g.we_clk [30341]));
Q_ASSIGN U2434 ( .B(clk), .A(\g.we_clk [30340]));
Q_ASSIGN U2435 ( .B(clk), .A(\g.we_clk [30339]));
Q_ASSIGN U2436 ( .B(clk), .A(\g.we_clk [30338]));
Q_ASSIGN U2437 ( .B(clk), .A(\g.we_clk [30337]));
Q_ASSIGN U2438 ( .B(clk), .A(\g.we_clk [30336]));
Q_ASSIGN U2439 ( .B(clk), .A(\g.we_clk [30335]));
Q_ASSIGN U2440 ( .B(clk), .A(\g.we_clk [30334]));
Q_ASSIGN U2441 ( .B(clk), .A(\g.we_clk [30333]));
Q_ASSIGN U2442 ( .B(clk), .A(\g.we_clk [30332]));
Q_ASSIGN U2443 ( .B(clk), .A(\g.we_clk [30331]));
Q_ASSIGN U2444 ( .B(clk), .A(\g.we_clk [30330]));
Q_ASSIGN U2445 ( .B(clk), .A(\g.we_clk [30329]));
Q_ASSIGN U2446 ( .B(clk), .A(\g.we_clk [30328]));
Q_ASSIGN U2447 ( .B(clk), .A(\g.we_clk [30327]));
Q_ASSIGN U2448 ( .B(clk), .A(\g.we_clk [30326]));
Q_ASSIGN U2449 ( .B(clk), .A(\g.we_clk [30325]));
Q_ASSIGN U2450 ( .B(clk), .A(\g.we_clk [30324]));
Q_ASSIGN U2451 ( .B(clk), .A(\g.we_clk [30323]));
Q_ASSIGN U2452 ( .B(clk), .A(\g.we_clk [30322]));
Q_ASSIGN U2453 ( .B(clk), .A(\g.we_clk [30321]));
Q_ASSIGN U2454 ( .B(clk), .A(\g.we_clk [30320]));
Q_ASSIGN U2455 ( .B(clk), .A(\g.we_clk [30319]));
Q_ASSIGN U2456 ( .B(clk), .A(\g.we_clk [30318]));
Q_ASSIGN U2457 ( .B(clk), .A(\g.we_clk [30317]));
Q_ASSIGN U2458 ( .B(clk), .A(\g.we_clk [30316]));
Q_ASSIGN U2459 ( .B(clk), .A(\g.we_clk [30315]));
Q_ASSIGN U2460 ( .B(clk), .A(\g.we_clk [30314]));
Q_ASSIGN U2461 ( .B(clk), .A(\g.we_clk [30313]));
Q_ASSIGN U2462 ( .B(clk), .A(\g.we_clk [30312]));
Q_ASSIGN U2463 ( .B(clk), .A(\g.we_clk [30311]));
Q_ASSIGN U2464 ( .B(clk), .A(\g.we_clk [30310]));
Q_ASSIGN U2465 ( .B(clk), .A(\g.we_clk [30309]));
Q_ASSIGN U2466 ( .B(clk), .A(\g.we_clk [30308]));
Q_ASSIGN U2467 ( .B(clk), .A(\g.we_clk [30307]));
Q_ASSIGN U2468 ( .B(clk), .A(\g.we_clk [30306]));
Q_ASSIGN U2469 ( .B(clk), .A(\g.we_clk [30305]));
Q_ASSIGN U2470 ( .B(clk), .A(\g.we_clk [30304]));
Q_ASSIGN U2471 ( .B(clk), .A(\g.we_clk [30303]));
Q_ASSIGN U2472 ( .B(clk), .A(\g.we_clk [30302]));
Q_ASSIGN U2473 ( .B(clk), .A(\g.we_clk [30301]));
Q_ASSIGN U2474 ( .B(clk), .A(\g.we_clk [30300]));
Q_ASSIGN U2475 ( .B(clk), .A(\g.we_clk [30299]));
Q_ASSIGN U2476 ( .B(clk), .A(\g.we_clk [30298]));
Q_ASSIGN U2477 ( .B(clk), .A(\g.we_clk [30297]));
Q_ASSIGN U2478 ( .B(clk), .A(\g.we_clk [30296]));
Q_ASSIGN U2479 ( .B(clk), .A(\g.we_clk [30295]));
Q_ASSIGN U2480 ( .B(clk), .A(\g.we_clk [30294]));
Q_ASSIGN U2481 ( .B(clk), .A(\g.we_clk [30293]));
Q_ASSIGN U2482 ( .B(clk), .A(\g.we_clk [30292]));
Q_ASSIGN U2483 ( .B(clk), .A(\g.we_clk [30291]));
Q_ASSIGN U2484 ( .B(clk), .A(\g.we_clk [30290]));
Q_ASSIGN U2485 ( .B(clk), .A(\g.we_clk [30289]));
Q_ASSIGN U2486 ( .B(clk), .A(\g.we_clk [30288]));
Q_ASSIGN U2487 ( .B(clk), .A(\g.we_clk [30287]));
Q_ASSIGN U2488 ( .B(clk), .A(\g.we_clk [30286]));
Q_ASSIGN U2489 ( .B(clk), .A(\g.we_clk [30285]));
Q_ASSIGN U2490 ( .B(clk), .A(\g.we_clk [30284]));
Q_ASSIGN U2491 ( .B(clk), .A(\g.we_clk [30283]));
Q_ASSIGN U2492 ( .B(clk), .A(\g.we_clk [30282]));
Q_ASSIGN U2493 ( .B(clk), .A(\g.we_clk [30281]));
Q_ASSIGN U2494 ( .B(clk), .A(\g.we_clk [30280]));
Q_ASSIGN U2495 ( .B(clk), .A(\g.we_clk [30279]));
Q_ASSIGN U2496 ( .B(clk), .A(\g.we_clk [30278]));
Q_ASSIGN U2497 ( .B(clk), .A(\g.we_clk [30277]));
Q_ASSIGN U2498 ( .B(clk), .A(\g.we_clk [30276]));
Q_ASSIGN U2499 ( .B(clk), .A(\g.we_clk [30275]));
Q_ASSIGN U2500 ( .B(clk), .A(\g.we_clk [30274]));
Q_ASSIGN U2501 ( .B(clk), .A(\g.we_clk [30273]));
Q_ASSIGN U2502 ( .B(clk), .A(\g.we_clk [30272]));
Q_ASSIGN U2503 ( .B(clk), .A(\g.we_clk [30271]));
Q_ASSIGN U2504 ( .B(clk), .A(\g.we_clk [30270]));
Q_ASSIGN U2505 ( .B(clk), .A(\g.we_clk [30269]));
Q_ASSIGN U2506 ( .B(clk), .A(\g.we_clk [30268]));
Q_ASSIGN U2507 ( .B(clk), .A(\g.we_clk [30267]));
Q_ASSIGN U2508 ( .B(clk), .A(\g.we_clk [30266]));
Q_ASSIGN U2509 ( .B(clk), .A(\g.we_clk [30265]));
Q_ASSIGN U2510 ( .B(clk), .A(\g.we_clk [30264]));
Q_ASSIGN U2511 ( .B(clk), .A(\g.we_clk [30263]));
Q_ASSIGN U2512 ( .B(clk), .A(\g.we_clk [30262]));
Q_ASSIGN U2513 ( .B(clk), .A(\g.we_clk [30261]));
Q_ASSIGN U2514 ( .B(clk), .A(\g.we_clk [30260]));
Q_ASSIGN U2515 ( .B(clk), .A(\g.we_clk [30259]));
Q_ASSIGN U2516 ( .B(clk), .A(\g.we_clk [30258]));
Q_ASSIGN U2517 ( .B(clk), .A(\g.we_clk [30257]));
Q_ASSIGN U2518 ( .B(clk), .A(\g.we_clk [30256]));
Q_ASSIGN U2519 ( .B(clk), .A(\g.we_clk [30255]));
Q_ASSIGN U2520 ( .B(clk), .A(\g.we_clk [30254]));
Q_ASSIGN U2521 ( .B(clk), .A(\g.we_clk [30253]));
Q_ASSIGN U2522 ( .B(clk), .A(\g.we_clk [30252]));
Q_ASSIGN U2523 ( .B(clk), .A(\g.we_clk [30251]));
Q_ASSIGN U2524 ( .B(clk), .A(\g.we_clk [30250]));
Q_ASSIGN U2525 ( .B(clk), .A(\g.we_clk [30249]));
Q_ASSIGN U2526 ( .B(clk), .A(\g.we_clk [30248]));
Q_ASSIGN U2527 ( .B(clk), .A(\g.we_clk [30247]));
Q_ASSIGN U2528 ( .B(clk), .A(\g.we_clk [30246]));
Q_ASSIGN U2529 ( .B(clk), .A(\g.we_clk [30245]));
Q_ASSIGN U2530 ( .B(clk), .A(\g.we_clk [30244]));
Q_ASSIGN U2531 ( .B(clk), .A(\g.we_clk [30243]));
Q_ASSIGN U2532 ( .B(clk), .A(\g.we_clk [30242]));
Q_ASSIGN U2533 ( .B(clk), .A(\g.we_clk [30241]));
Q_ASSIGN U2534 ( .B(clk), .A(\g.we_clk [30240]));
Q_ASSIGN U2535 ( .B(clk), .A(\g.we_clk [30239]));
Q_ASSIGN U2536 ( .B(clk), .A(\g.we_clk [30238]));
Q_ASSIGN U2537 ( .B(clk), .A(\g.we_clk [30237]));
Q_ASSIGN U2538 ( .B(clk), .A(\g.we_clk [30236]));
Q_ASSIGN U2539 ( .B(clk), .A(\g.we_clk [30235]));
Q_ASSIGN U2540 ( .B(clk), .A(\g.we_clk [30234]));
Q_ASSIGN U2541 ( .B(clk), .A(\g.we_clk [30233]));
Q_ASSIGN U2542 ( .B(clk), .A(\g.we_clk [30232]));
Q_ASSIGN U2543 ( .B(clk), .A(\g.we_clk [30231]));
Q_ASSIGN U2544 ( .B(clk), .A(\g.we_clk [30230]));
Q_ASSIGN U2545 ( .B(clk), .A(\g.we_clk [30229]));
Q_ASSIGN U2546 ( .B(clk), .A(\g.we_clk [30228]));
Q_ASSIGN U2547 ( .B(clk), .A(\g.we_clk [30227]));
Q_ASSIGN U2548 ( .B(clk), .A(\g.we_clk [30226]));
Q_ASSIGN U2549 ( .B(clk), .A(\g.we_clk [30225]));
Q_ASSIGN U2550 ( .B(clk), .A(\g.we_clk [30224]));
Q_ASSIGN U2551 ( .B(clk), .A(\g.we_clk [30223]));
Q_ASSIGN U2552 ( .B(clk), .A(\g.we_clk [30222]));
Q_ASSIGN U2553 ( .B(clk), .A(\g.we_clk [30221]));
Q_ASSIGN U2554 ( .B(clk), .A(\g.we_clk [30220]));
Q_ASSIGN U2555 ( .B(clk), .A(\g.we_clk [30219]));
Q_ASSIGN U2556 ( .B(clk), .A(\g.we_clk [30218]));
Q_ASSIGN U2557 ( .B(clk), .A(\g.we_clk [30217]));
Q_ASSIGN U2558 ( .B(clk), .A(\g.we_clk [30216]));
Q_ASSIGN U2559 ( .B(clk), .A(\g.we_clk [30215]));
Q_ASSIGN U2560 ( .B(clk), .A(\g.we_clk [30214]));
Q_ASSIGN U2561 ( .B(clk), .A(\g.we_clk [30213]));
Q_ASSIGN U2562 ( .B(clk), .A(\g.we_clk [30212]));
Q_ASSIGN U2563 ( .B(clk), .A(\g.we_clk [30211]));
Q_ASSIGN U2564 ( .B(clk), .A(\g.we_clk [30210]));
Q_ASSIGN U2565 ( .B(clk), .A(\g.we_clk [30209]));
Q_ASSIGN U2566 ( .B(clk), .A(\g.we_clk [30208]));
Q_ASSIGN U2567 ( .B(clk), .A(\g.we_clk [30207]));
Q_ASSIGN U2568 ( .B(clk), .A(\g.we_clk [30206]));
Q_ASSIGN U2569 ( .B(clk), .A(\g.we_clk [30205]));
Q_ASSIGN U2570 ( .B(clk), .A(\g.we_clk [30204]));
Q_ASSIGN U2571 ( .B(clk), .A(\g.we_clk [30203]));
Q_ASSIGN U2572 ( .B(clk), .A(\g.we_clk [30202]));
Q_ASSIGN U2573 ( .B(clk), .A(\g.we_clk [30201]));
Q_ASSIGN U2574 ( .B(clk), .A(\g.we_clk [30200]));
Q_ASSIGN U2575 ( .B(clk), .A(\g.we_clk [30199]));
Q_ASSIGN U2576 ( .B(clk), .A(\g.we_clk [30198]));
Q_ASSIGN U2577 ( .B(clk), .A(\g.we_clk [30197]));
Q_ASSIGN U2578 ( .B(clk), .A(\g.we_clk [30196]));
Q_ASSIGN U2579 ( .B(clk), .A(\g.we_clk [30195]));
Q_ASSIGN U2580 ( .B(clk), .A(\g.we_clk [30194]));
Q_ASSIGN U2581 ( .B(clk), .A(\g.we_clk [30193]));
Q_ASSIGN U2582 ( .B(clk), .A(\g.we_clk [30192]));
Q_ASSIGN U2583 ( .B(clk), .A(\g.we_clk [30191]));
Q_ASSIGN U2584 ( .B(clk), .A(\g.we_clk [30190]));
Q_ASSIGN U2585 ( .B(clk), .A(\g.we_clk [30189]));
Q_ASSIGN U2586 ( .B(clk), .A(\g.we_clk [30188]));
Q_ASSIGN U2587 ( .B(clk), .A(\g.we_clk [30187]));
Q_ASSIGN U2588 ( .B(clk), .A(\g.we_clk [30186]));
Q_ASSIGN U2589 ( .B(clk), .A(\g.we_clk [30185]));
Q_ASSIGN U2590 ( .B(clk), .A(\g.we_clk [30184]));
Q_ASSIGN U2591 ( .B(clk), .A(\g.we_clk [30183]));
Q_ASSIGN U2592 ( .B(clk), .A(\g.we_clk [30182]));
Q_ASSIGN U2593 ( .B(clk), .A(\g.we_clk [30181]));
Q_ASSIGN U2594 ( .B(clk), .A(\g.we_clk [30180]));
Q_ASSIGN U2595 ( .B(clk), .A(\g.we_clk [30179]));
Q_ASSIGN U2596 ( .B(clk), .A(\g.we_clk [30178]));
Q_ASSIGN U2597 ( .B(clk), .A(\g.we_clk [30177]));
Q_ASSIGN U2598 ( .B(clk), .A(\g.we_clk [30176]));
Q_ASSIGN U2599 ( .B(clk), .A(\g.we_clk [30175]));
Q_ASSIGN U2600 ( .B(clk), .A(\g.we_clk [30174]));
Q_ASSIGN U2601 ( .B(clk), .A(\g.we_clk [30173]));
Q_ASSIGN U2602 ( .B(clk), .A(\g.we_clk [30172]));
Q_ASSIGN U2603 ( .B(clk), .A(\g.we_clk [30171]));
Q_ASSIGN U2604 ( .B(clk), .A(\g.we_clk [30170]));
Q_ASSIGN U2605 ( .B(clk), .A(\g.we_clk [30169]));
Q_ASSIGN U2606 ( .B(clk), .A(\g.we_clk [30168]));
Q_ASSIGN U2607 ( .B(clk), .A(\g.we_clk [30167]));
Q_ASSIGN U2608 ( .B(clk), .A(\g.we_clk [30166]));
Q_ASSIGN U2609 ( .B(clk), .A(\g.we_clk [30165]));
Q_ASSIGN U2610 ( .B(clk), .A(\g.we_clk [30164]));
Q_ASSIGN U2611 ( .B(clk), .A(\g.we_clk [30163]));
Q_ASSIGN U2612 ( .B(clk), .A(\g.we_clk [30162]));
Q_ASSIGN U2613 ( .B(clk), .A(\g.we_clk [30161]));
Q_ASSIGN U2614 ( .B(clk), .A(\g.we_clk [30160]));
Q_ASSIGN U2615 ( .B(clk), .A(\g.we_clk [30159]));
Q_ASSIGN U2616 ( .B(clk), .A(\g.we_clk [30158]));
Q_ASSIGN U2617 ( .B(clk), .A(\g.we_clk [30157]));
Q_ASSIGN U2618 ( .B(clk), .A(\g.we_clk [30156]));
Q_ASSIGN U2619 ( .B(clk), .A(\g.we_clk [30155]));
Q_ASSIGN U2620 ( .B(clk), .A(\g.we_clk [30154]));
Q_ASSIGN U2621 ( .B(clk), .A(\g.we_clk [30153]));
Q_ASSIGN U2622 ( .B(clk), .A(\g.we_clk [30152]));
Q_ASSIGN U2623 ( .B(clk), .A(\g.we_clk [30151]));
Q_ASSIGN U2624 ( .B(clk), .A(\g.we_clk [30150]));
Q_ASSIGN U2625 ( .B(clk), .A(\g.we_clk [30149]));
Q_ASSIGN U2626 ( .B(clk), .A(\g.we_clk [30148]));
Q_ASSIGN U2627 ( .B(clk), .A(\g.we_clk [30147]));
Q_ASSIGN U2628 ( .B(clk), .A(\g.we_clk [30146]));
Q_ASSIGN U2629 ( .B(clk), .A(\g.we_clk [30145]));
Q_ASSIGN U2630 ( .B(clk), .A(\g.we_clk [30144]));
Q_ASSIGN U2631 ( .B(clk), .A(\g.we_clk [30143]));
Q_ASSIGN U2632 ( .B(clk), .A(\g.we_clk [30142]));
Q_ASSIGN U2633 ( .B(clk), .A(\g.we_clk [30141]));
Q_ASSIGN U2634 ( .B(clk), .A(\g.we_clk [30140]));
Q_ASSIGN U2635 ( .B(clk), .A(\g.we_clk [30139]));
Q_ASSIGN U2636 ( .B(clk), .A(\g.we_clk [30138]));
Q_ASSIGN U2637 ( .B(clk), .A(\g.we_clk [30137]));
Q_ASSIGN U2638 ( .B(clk), .A(\g.we_clk [30136]));
Q_ASSIGN U2639 ( .B(clk), .A(\g.we_clk [30135]));
Q_ASSIGN U2640 ( .B(clk), .A(\g.we_clk [30134]));
Q_ASSIGN U2641 ( .B(clk), .A(\g.we_clk [30133]));
Q_ASSIGN U2642 ( .B(clk), .A(\g.we_clk [30132]));
Q_ASSIGN U2643 ( .B(clk), .A(\g.we_clk [30131]));
Q_ASSIGN U2644 ( .B(clk), .A(\g.we_clk [30130]));
Q_ASSIGN U2645 ( .B(clk), .A(\g.we_clk [30129]));
Q_ASSIGN U2646 ( .B(clk), .A(\g.we_clk [30128]));
Q_ASSIGN U2647 ( .B(clk), .A(\g.we_clk [30127]));
Q_ASSIGN U2648 ( .B(clk), .A(\g.we_clk [30126]));
Q_ASSIGN U2649 ( .B(clk), .A(\g.we_clk [30125]));
Q_ASSIGN U2650 ( .B(clk), .A(\g.we_clk [30124]));
Q_ASSIGN U2651 ( .B(clk), .A(\g.we_clk [30123]));
Q_ASSIGN U2652 ( .B(clk), .A(\g.we_clk [30122]));
Q_ASSIGN U2653 ( .B(clk), .A(\g.we_clk [30121]));
Q_ASSIGN U2654 ( .B(clk), .A(\g.we_clk [30120]));
Q_ASSIGN U2655 ( .B(clk), .A(\g.we_clk [30119]));
Q_ASSIGN U2656 ( .B(clk), .A(\g.we_clk [30118]));
Q_ASSIGN U2657 ( .B(clk), .A(\g.we_clk [30117]));
Q_ASSIGN U2658 ( .B(clk), .A(\g.we_clk [30116]));
Q_ASSIGN U2659 ( .B(clk), .A(\g.we_clk [30115]));
Q_ASSIGN U2660 ( .B(clk), .A(\g.we_clk [30114]));
Q_ASSIGN U2661 ( .B(clk), .A(\g.we_clk [30113]));
Q_ASSIGN U2662 ( .B(clk), .A(\g.we_clk [30112]));
Q_ASSIGN U2663 ( .B(clk), .A(\g.we_clk [30111]));
Q_ASSIGN U2664 ( .B(clk), .A(\g.we_clk [30110]));
Q_ASSIGN U2665 ( .B(clk), .A(\g.we_clk [30109]));
Q_ASSIGN U2666 ( .B(clk), .A(\g.we_clk [30108]));
Q_ASSIGN U2667 ( .B(clk), .A(\g.we_clk [30107]));
Q_ASSIGN U2668 ( .B(clk), .A(\g.we_clk [30106]));
Q_ASSIGN U2669 ( .B(clk), .A(\g.we_clk [30105]));
Q_ASSIGN U2670 ( .B(clk), .A(\g.we_clk [30104]));
Q_ASSIGN U2671 ( .B(clk), .A(\g.we_clk [30103]));
Q_ASSIGN U2672 ( .B(clk), .A(\g.we_clk [30102]));
Q_ASSIGN U2673 ( .B(clk), .A(\g.we_clk [30101]));
Q_ASSIGN U2674 ( .B(clk), .A(\g.we_clk [30100]));
Q_ASSIGN U2675 ( .B(clk), .A(\g.we_clk [30099]));
Q_ASSIGN U2676 ( .B(clk), .A(\g.we_clk [30098]));
Q_ASSIGN U2677 ( .B(clk), .A(\g.we_clk [30097]));
Q_ASSIGN U2678 ( .B(clk), .A(\g.we_clk [30096]));
Q_ASSIGN U2679 ( .B(clk), .A(\g.we_clk [30095]));
Q_ASSIGN U2680 ( .B(clk), .A(\g.we_clk [30094]));
Q_ASSIGN U2681 ( .B(clk), .A(\g.we_clk [30093]));
Q_ASSIGN U2682 ( .B(clk), .A(\g.we_clk [30092]));
Q_ASSIGN U2683 ( .B(clk), .A(\g.we_clk [30091]));
Q_ASSIGN U2684 ( .B(clk), .A(\g.we_clk [30090]));
Q_ASSIGN U2685 ( .B(clk), .A(\g.we_clk [30089]));
Q_ASSIGN U2686 ( .B(clk), .A(\g.we_clk [30088]));
Q_ASSIGN U2687 ( .B(clk), .A(\g.we_clk [30087]));
Q_ASSIGN U2688 ( .B(clk), .A(\g.we_clk [30086]));
Q_ASSIGN U2689 ( .B(clk), .A(\g.we_clk [30085]));
Q_ASSIGN U2690 ( .B(clk), .A(\g.we_clk [30084]));
Q_ASSIGN U2691 ( .B(clk), .A(\g.we_clk [30083]));
Q_ASSIGN U2692 ( .B(clk), .A(\g.we_clk [30082]));
Q_ASSIGN U2693 ( .B(clk), .A(\g.we_clk [30081]));
Q_ASSIGN U2694 ( .B(clk), .A(\g.we_clk [30080]));
Q_ASSIGN U2695 ( .B(clk), .A(\g.we_clk [30079]));
Q_ASSIGN U2696 ( .B(clk), .A(\g.we_clk [30078]));
Q_ASSIGN U2697 ( .B(clk), .A(\g.we_clk [30077]));
Q_ASSIGN U2698 ( .B(clk), .A(\g.we_clk [30076]));
Q_ASSIGN U2699 ( .B(clk), .A(\g.we_clk [30075]));
Q_ASSIGN U2700 ( .B(clk), .A(\g.we_clk [30074]));
Q_ASSIGN U2701 ( .B(clk), .A(\g.we_clk [30073]));
Q_ASSIGN U2702 ( .B(clk), .A(\g.we_clk [30072]));
Q_ASSIGN U2703 ( .B(clk), .A(\g.we_clk [30071]));
Q_ASSIGN U2704 ( .B(clk), .A(\g.we_clk [30070]));
Q_ASSIGN U2705 ( .B(clk), .A(\g.we_clk [30069]));
Q_ASSIGN U2706 ( .B(clk), .A(\g.we_clk [30068]));
Q_ASSIGN U2707 ( .B(clk), .A(\g.we_clk [30067]));
Q_ASSIGN U2708 ( .B(clk), .A(\g.we_clk [30066]));
Q_ASSIGN U2709 ( .B(clk), .A(\g.we_clk [30065]));
Q_ASSIGN U2710 ( .B(clk), .A(\g.we_clk [30064]));
Q_ASSIGN U2711 ( .B(clk), .A(\g.we_clk [30063]));
Q_ASSIGN U2712 ( .B(clk), .A(\g.we_clk [30062]));
Q_ASSIGN U2713 ( .B(clk), .A(\g.we_clk [30061]));
Q_ASSIGN U2714 ( .B(clk), .A(\g.we_clk [30060]));
Q_ASSIGN U2715 ( .B(clk), .A(\g.we_clk [30059]));
Q_ASSIGN U2716 ( .B(clk), .A(\g.we_clk [30058]));
Q_ASSIGN U2717 ( .B(clk), .A(\g.we_clk [30057]));
Q_ASSIGN U2718 ( .B(clk), .A(\g.we_clk [30056]));
Q_ASSIGN U2719 ( .B(clk), .A(\g.we_clk [30055]));
Q_ASSIGN U2720 ( .B(clk), .A(\g.we_clk [30054]));
Q_ASSIGN U2721 ( .B(clk), .A(\g.we_clk [30053]));
Q_ASSIGN U2722 ( .B(clk), .A(\g.we_clk [30052]));
Q_ASSIGN U2723 ( .B(clk), .A(\g.we_clk [30051]));
Q_ASSIGN U2724 ( .B(clk), .A(\g.we_clk [30050]));
Q_ASSIGN U2725 ( .B(clk), .A(\g.we_clk [30049]));
Q_ASSIGN U2726 ( .B(clk), .A(\g.we_clk [30048]));
Q_ASSIGN U2727 ( .B(clk), .A(\g.we_clk [30047]));
Q_ASSIGN U2728 ( .B(clk), .A(\g.we_clk [30046]));
Q_ASSIGN U2729 ( .B(clk), .A(\g.we_clk [30045]));
Q_ASSIGN U2730 ( .B(clk), .A(\g.we_clk [30044]));
Q_ASSIGN U2731 ( .B(clk), .A(\g.we_clk [30043]));
Q_ASSIGN U2732 ( .B(clk), .A(\g.we_clk [30042]));
Q_ASSIGN U2733 ( .B(clk), .A(\g.we_clk [30041]));
Q_ASSIGN U2734 ( .B(clk), .A(\g.we_clk [30040]));
Q_ASSIGN U2735 ( .B(clk), .A(\g.we_clk [30039]));
Q_ASSIGN U2736 ( .B(clk), .A(\g.we_clk [30038]));
Q_ASSIGN U2737 ( .B(clk), .A(\g.we_clk [30037]));
Q_ASSIGN U2738 ( .B(clk), .A(\g.we_clk [30036]));
Q_ASSIGN U2739 ( .B(clk), .A(\g.we_clk [30035]));
Q_ASSIGN U2740 ( .B(clk), .A(\g.we_clk [30034]));
Q_ASSIGN U2741 ( .B(clk), .A(\g.we_clk [30033]));
Q_ASSIGN U2742 ( .B(clk), .A(\g.we_clk [30032]));
Q_ASSIGN U2743 ( .B(clk), .A(\g.we_clk [30031]));
Q_ASSIGN U2744 ( .B(clk), .A(\g.we_clk [30030]));
Q_ASSIGN U2745 ( .B(clk), .A(\g.we_clk [30029]));
Q_ASSIGN U2746 ( .B(clk), .A(\g.we_clk [30028]));
Q_ASSIGN U2747 ( .B(clk), .A(\g.we_clk [30027]));
Q_ASSIGN U2748 ( .B(clk), .A(\g.we_clk [30026]));
Q_ASSIGN U2749 ( .B(clk), .A(\g.we_clk [30025]));
Q_ASSIGN U2750 ( .B(clk), .A(\g.we_clk [30024]));
Q_ASSIGN U2751 ( .B(clk), .A(\g.we_clk [30023]));
Q_ASSIGN U2752 ( .B(clk), .A(\g.we_clk [30022]));
Q_ASSIGN U2753 ( .B(clk), .A(\g.we_clk [30021]));
Q_ASSIGN U2754 ( .B(clk), .A(\g.we_clk [30020]));
Q_ASSIGN U2755 ( .B(clk), .A(\g.we_clk [30019]));
Q_ASSIGN U2756 ( .B(clk), .A(\g.we_clk [30018]));
Q_ASSIGN U2757 ( .B(clk), .A(\g.we_clk [30017]));
Q_ASSIGN U2758 ( .B(clk), .A(\g.we_clk [30016]));
Q_ASSIGN U2759 ( .B(clk), .A(\g.we_clk [30015]));
Q_ASSIGN U2760 ( .B(clk), .A(\g.we_clk [30014]));
Q_ASSIGN U2761 ( .B(clk), .A(\g.we_clk [30013]));
Q_ASSIGN U2762 ( .B(clk), .A(\g.we_clk [30012]));
Q_ASSIGN U2763 ( .B(clk), .A(\g.we_clk [30011]));
Q_ASSIGN U2764 ( .B(clk), .A(\g.we_clk [30010]));
Q_ASSIGN U2765 ( .B(clk), .A(\g.we_clk [30009]));
Q_ASSIGN U2766 ( .B(clk), .A(\g.we_clk [30008]));
Q_ASSIGN U2767 ( .B(clk), .A(\g.we_clk [30007]));
Q_ASSIGN U2768 ( .B(clk), .A(\g.we_clk [30006]));
Q_ASSIGN U2769 ( .B(clk), .A(\g.we_clk [30005]));
Q_ASSIGN U2770 ( .B(clk), .A(\g.we_clk [30004]));
Q_ASSIGN U2771 ( .B(clk), .A(\g.we_clk [30003]));
Q_ASSIGN U2772 ( .B(clk), .A(\g.we_clk [30002]));
Q_ASSIGN U2773 ( .B(clk), .A(\g.we_clk [30001]));
Q_ASSIGN U2774 ( .B(clk), .A(\g.we_clk [30000]));
Q_ASSIGN U2775 ( .B(clk), .A(\g.we_clk [29999]));
Q_ASSIGN U2776 ( .B(clk), .A(\g.we_clk [29998]));
Q_ASSIGN U2777 ( .B(clk), .A(\g.we_clk [29997]));
Q_ASSIGN U2778 ( .B(clk), .A(\g.we_clk [29996]));
Q_ASSIGN U2779 ( .B(clk), .A(\g.we_clk [29995]));
Q_ASSIGN U2780 ( .B(clk), .A(\g.we_clk [29994]));
Q_ASSIGN U2781 ( .B(clk), .A(\g.we_clk [29993]));
Q_ASSIGN U2782 ( .B(clk), .A(\g.we_clk [29992]));
Q_ASSIGN U2783 ( .B(clk), .A(\g.we_clk [29991]));
Q_ASSIGN U2784 ( .B(clk), .A(\g.we_clk [29990]));
Q_ASSIGN U2785 ( .B(clk), .A(\g.we_clk [29989]));
Q_ASSIGN U2786 ( .B(clk), .A(\g.we_clk [29988]));
Q_ASSIGN U2787 ( .B(clk), .A(\g.we_clk [29987]));
Q_ASSIGN U2788 ( .B(clk), .A(\g.we_clk [29986]));
Q_ASSIGN U2789 ( .B(clk), .A(\g.we_clk [29985]));
Q_ASSIGN U2790 ( .B(clk), .A(\g.we_clk [29984]));
Q_ASSIGN U2791 ( .B(clk), .A(\g.we_clk [29983]));
Q_ASSIGN U2792 ( .B(clk), .A(\g.we_clk [29982]));
Q_ASSIGN U2793 ( .B(clk), .A(\g.we_clk [29981]));
Q_ASSIGN U2794 ( .B(clk), .A(\g.we_clk [29980]));
Q_ASSIGN U2795 ( .B(clk), .A(\g.we_clk [29979]));
Q_ASSIGN U2796 ( .B(clk), .A(\g.we_clk [29978]));
Q_ASSIGN U2797 ( .B(clk), .A(\g.we_clk [29977]));
Q_ASSIGN U2798 ( .B(clk), .A(\g.we_clk [29976]));
Q_ASSIGN U2799 ( .B(clk), .A(\g.we_clk [29975]));
Q_ASSIGN U2800 ( .B(clk), .A(\g.we_clk [29974]));
Q_ASSIGN U2801 ( .B(clk), .A(\g.we_clk [29973]));
Q_ASSIGN U2802 ( .B(clk), .A(\g.we_clk [29972]));
Q_ASSIGN U2803 ( .B(clk), .A(\g.we_clk [29971]));
Q_ASSIGN U2804 ( .B(clk), .A(\g.we_clk [29970]));
Q_ASSIGN U2805 ( .B(clk), .A(\g.we_clk [29969]));
Q_ASSIGN U2806 ( .B(clk), .A(\g.we_clk [29968]));
Q_ASSIGN U2807 ( .B(clk), .A(\g.we_clk [29967]));
Q_ASSIGN U2808 ( .B(clk), .A(\g.we_clk [29966]));
Q_ASSIGN U2809 ( .B(clk), .A(\g.we_clk [29965]));
Q_ASSIGN U2810 ( .B(clk), .A(\g.we_clk [29964]));
Q_ASSIGN U2811 ( .B(clk), .A(\g.we_clk [29963]));
Q_ASSIGN U2812 ( .B(clk), .A(\g.we_clk [29962]));
Q_ASSIGN U2813 ( .B(clk), .A(\g.we_clk [29961]));
Q_ASSIGN U2814 ( .B(clk), .A(\g.we_clk [29960]));
Q_ASSIGN U2815 ( .B(clk), .A(\g.we_clk [29959]));
Q_ASSIGN U2816 ( .B(clk), .A(\g.we_clk [29958]));
Q_ASSIGN U2817 ( .B(clk), .A(\g.we_clk [29957]));
Q_ASSIGN U2818 ( .B(clk), .A(\g.we_clk [29956]));
Q_ASSIGN U2819 ( .B(clk), .A(\g.we_clk [29955]));
Q_ASSIGN U2820 ( .B(clk), .A(\g.we_clk [29954]));
Q_ASSIGN U2821 ( .B(clk), .A(\g.we_clk [29953]));
Q_ASSIGN U2822 ( .B(clk), .A(\g.we_clk [29952]));
Q_ASSIGN U2823 ( .B(clk), .A(\g.we_clk [29951]));
Q_ASSIGN U2824 ( .B(clk), .A(\g.we_clk [29950]));
Q_ASSIGN U2825 ( .B(clk), .A(\g.we_clk [29949]));
Q_ASSIGN U2826 ( .B(clk), .A(\g.we_clk [29948]));
Q_ASSIGN U2827 ( .B(clk), .A(\g.we_clk [29947]));
Q_ASSIGN U2828 ( .B(clk), .A(\g.we_clk [29946]));
Q_ASSIGN U2829 ( .B(clk), .A(\g.we_clk [29945]));
Q_ASSIGN U2830 ( .B(clk), .A(\g.we_clk [29944]));
Q_ASSIGN U2831 ( .B(clk), .A(\g.we_clk [29943]));
Q_ASSIGN U2832 ( .B(clk), .A(\g.we_clk [29942]));
Q_ASSIGN U2833 ( .B(clk), .A(\g.we_clk [29941]));
Q_ASSIGN U2834 ( .B(clk), .A(\g.we_clk [29940]));
Q_ASSIGN U2835 ( .B(clk), .A(\g.we_clk [29939]));
Q_ASSIGN U2836 ( .B(clk), .A(\g.we_clk [29938]));
Q_ASSIGN U2837 ( .B(clk), .A(\g.we_clk [29937]));
Q_ASSIGN U2838 ( .B(clk), .A(\g.we_clk [29936]));
Q_ASSIGN U2839 ( .B(clk), .A(\g.we_clk [29935]));
Q_ASSIGN U2840 ( .B(clk), .A(\g.we_clk [29934]));
Q_ASSIGN U2841 ( .B(clk), .A(\g.we_clk [29933]));
Q_ASSIGN U2842 ( .B(clk), .A(\g.we_clk [29932]));
Q_ASSIGN U2843 ( .B(clk), .A(\g.we_clk [29931]));
Q_ASSIGN U2844 ( .B(clk), .A(\g.we_clk [29930]));
Q_ASSIGN U2845 ( .B(clk), .A(\g.we_clk [29929]));
Q_ASSIGN U2846 ( .B(clk), .A(\g.we_clk [29928]));
Q_ASSIGN U2847 ( .B(clk), .A(\g.we_clk [29927]));
Q_ASSIGN U2848 ( .B(clk), .A(\g.we_clk [29926]));
Q_ASSIGN U2849 ( .B(clk), .A(\g.we_clk [29925]));
Q_ASSIGN U2850 ( .B(clk), .A(\g.we_clk [29924]));
Q_ASSIGN U2851 ( .B(clk), .A(\g.we_clk [29923]));
Q_ASSIGN U2852 ( .B(clk), .A(\g.we_clk [29922]));
Q_ASSIGN U2853 ( .B(clk), .A(\g.we_clk [29921]));
Q_ASSIGN U2854 ( .B(clk), .A(\g.we_clk [29920]));
Q_ASSIGN U2855 ( .B(clk), .A(\g.we_clk [29919]));
Q_ASSIGN U2856 ( .B(clk), .A(\g.we_clk [29918]));
Q_ASSIGN U2857 ( .B(clk), .A(\g.we_clk [29917]));
Q_ASSIGN U2858 ( .B(clk), .A(\g.we_clk [29916]));
Q_ASSIGN U2859 ( .B(clk), .A(\g.we_clk [29915]));
Q_ASSIGN U2860 ( .B(clk), .A(\g.we_clk [29914]));
Q_ASSIGN U2861 ( .B(clk), .A(\g.we_clk [29913]));
Q_ASSIGN U2862 ( .B(clk), .A(\g.we_clk [29912]));
Q_ASSIGN U2863 ( .B(clk), .A(\g.we_clk [29911]));
Q_ASSIGN U2864 ( .B(clk), .A(\g.we_clk [29910]));
Q_ASSIGN U2865 ( .B(clk), .A(\g.we_clk [29909]));
Q_ASSIGN U2866 ( .B(clk), .A(\g.we_clk [29908]));
Q_ASSIGN U2867 ( .B(clk), .A(\g.we_clk [29907]));
Q_ASSIGN U2868 ( .B(clk), .A(\g.we_clk [29906]));
Q_ASSIGN U2869 ( .B(clk), .A(\g.we_clk [29905]));
Q_ASSIGN U2870 ( .B(clk), .A(\g.we_clk [29904]));
Q_ASSIGN U2871 ( .B(clk), .A(\g.we_clk [29903]));
Q_ASSIGN U2872 ( .B(clk), .A(\g.we_clk [29902]));
Q_ASSIGN U2873 ( .B(clk), .A(\g.we_clk [29901]));
Q_ASSIGN U2874 ( .B(clk), .A(\g.we_clk [29900]));
Q_ASSIGN U2875 ( .B(clk), .A(\g.we_clk [29899]));
Q_ASSIGN U2876 ( .B(clk), .A(\g.we_clk [29898]));
Q_ASSIGN U2877 ( .B(clk), .A(\g.we_clk [29897]));
Q_ASSIGN U2878 ( .B(clk), .A(\g.we_clk [29896]));
Q_ASSIGN U2879 ( .B(clk), .A(\g.we_clk [29895]));
Q_ASSIGN U2880 ( .B(clk), .A(\g.we_clk [29894]));
Q_ASSIGN U2881 ( .B(clk), .A(\g.we_clk [29893]));
Q_ASSIGN U2882 ( .B(clk), .A(\g.we_clk [29892]));
Q_ASSIGN U2883 ( .B(clk), .A(\g.we_clk [29891]));
Q_ASSIGN U2884 ( .B(clk), .A(\g.we_clk [29890]));
Q_ASSIGN U2885 ( .B(clk), .A(\g.we_clk [29889]));
Q_ASSIGN U2886 ( .B(clk), .A(\g.we_clk [29888]));
Q_ASSIGN U2887 ( .B(clk), .A(\g.we_clk [29887]));
Q_ASSIGN U2888 ( .B(clk), .A(\g.we_clk [29886]));
Q_ASSIGN U2889 ( .B(clk), .A(\g.we_clk [29885]));
Q_ASSIGN U2890 ( .B(clk), .A(\g.we_clk [29884]));
Q_ASSIGN U2891 ( .B(clk), .A(\g.we_clk [29883]));
Q_ASSIGN U2892 ( .B(clk), .A(\g.we_clk [29882]));
Q_ASSIGN U2893 ( .B(clk), .A(\g.we_clk [29881]));
Q_ASSIGN U2894 ( .B(clk), .A(\g.we_clk [29880]));
Q_ASSIGN U2895 ( .B(clk), .A(\g.we_clk [29879]));
Q_ASSIGN U2896 ( .B(clk), .A(\g.we_clk [29878]));
Q_ASSIGN U2897 ( .B(clk), .A(\g.we_clk [29877]));
Q_ASSIGN U2898 ( .B(clk), .A(\g.we_clk [29876]));
Q_ASSIGN U2899 ( .B(clk), .A(\g.we_clk [29875]));
Q_ASSIGN U2900 ( .B(clk), .A(\g.we_clk [29874]));
Q_ASSIGN U2901 ( .B(clk), .A(\g.we_clk [29873]));
Q_ASSIGN U2902 ( .B(clk), .A(\g.we_clk [29872]));
Q_ASSIGN U2903 ( .B(clk), .A(\g.we_clk [29871]));
Q_ASSIGN U2904 ( .B(clk), .A(\g.we_clk [29870]));
Q_ASSIGN U2905 ( .B(clk), .A(\g.we_clk [29869]));
Q_ASSIGN U2906 ( .B(clk), .A(\g.we_clk [29868]));
Q_ASSIGN U2907 ( .B(clk), .A(\g.we_clk [29867]));
Q_ASSIGN U2908 ( .B(clk), .A(\g.we_clk [29866]));
Q_ASSIGN U2909 ( .B(clk), .A(\g.we_clk [29865]));
Q_ASSIGN U2910 ( .B(clk), .A(\g.we_clk [29864]));
Q_ASSIGN U2911 ( .B(clk), .A(\g.we_clk [29863]));
Q_ASSIGN U2912 ( .B(clk), .A(\g.we_clk [29862]));
Q_ASSIGN U2913 ( .B(clk), .A(\g.we_clk [29861]));
Q_ASSIGN U2914 ( .B(clk), .A(\g.we_clk [29860]));
Q_ASSIGN U2915 ( .B(clk), .A(\g.we_clk [29859]));
Q_ASSIGN U2916 ( .B(clk), .A(\g.we_clk [29858]));
Q_ASSIGN U2917 ( .B(clk), .A(\g.we_clk [29857]));
Q_ASSIGN U2918 ( .B(clk), .A(\g.we_clk [29856]));
Q_ASSIGN U2919 ( .B(clk), .A(\g.we_clk [29855]));
Q_ASSIGN U2920 ( .B(clk), .A(\g.we_clk [29854]));
Q_ASSIGN U2921 ( .B(clk), .A(\g.we_clk [29853]));
Q_ASSIGN U2922 ( .B(clk), .A(\g.we_clk [29852]));
Q_ASSIGN U2923 ( .B(clk), .A(\g.we_clk [29851]));
Q_ASSIGN U2924 ( .B(clk), .A(\g.we_clk [29850]));
Q_ASSIGN U2925 ( .B(clk), .A(\g.we_clk [29849]));
Q_ASSIGN U2926 ( .B(clk), .A(\g.we_clk [29848]));
Q_ASSIGN U2927 ( .B(clk), .A(\g.we_clk [29847]));
Q_ASSIGN U2928 ( .B(clk), .A(\g.we_clk [29846]));
Q_ASSIGN U2929 ( .B(clk), .A(\g.we_clk [29845]));
Q_ASSIGN U2930 ( .B(clk), .A(\g.we_clk [29844]));
Q_ASSIGN U2931 ( .B(clk), .A(\g.we_clk [29843]));
Q_ASSIGN U2932 ( .B(clk), .A(\g.we_clk [29842]));
Q_ASSIGN U2933 ( .B(clk), .A(\g.we_clk [29841]));
Q_ASSIGN U2934 ( .B(clk), .A(\g.we_clk [29840]));
Q_ASSIGN U2935 ( .B(clk), .A(\g.we_clk [29839]));
Q_ASSIGN U2936 ( .B(clk), .A(\g.we_clk [29838]));
Q_ASSIGN U2937 ( .B(clk), .A(\g.we_clk [29837]));
Q_ASSIGN U2938 ( .B(clk), .A(\g.we_clk [29836]));
Q_ASSIGN U2939 ( .B(clk), .A(\g.we_clk [29835]));
Q_ASSIGN U2940 ( .B(clk), .A(\g.we_clk [29834]));
Q_ASSIGN U2941 ( .B(clk), .A(\g.we_clk [29833]));
Q_ASSIGN U2942 ( .B(clk), .A(\g.we_clk [29832]));
Q_ASSIGN U2943 ( .B(clk), .A(\g.we_clk [29831]));
Q_ASSIGN U2944 ( .B(clk), .A(\g.we_clk [29830]));
Q_ASSIGN U2945 ( .B(clk), .A(\g.we_clk [29829]));
Q_ASSIGN U2946 ( .B(clk), .A(\g.we_clk [29828]));
Q_ASSIGN U2947 ( .B(clk), .A(\g.we_clk [29827]));
Q_ASSIGN U2948 ( .B(clk), .A(\g.we_clk [29826]));
Q_ASSIGN U2949 ( .B(clk), .A(\g.we_clk [29825]));
Q_ASSIGN U2950 ( .B(clk), .A(\g.we_clk [29824]));
Q_ASSIGN U2951 ( .B(clk), .A(\g.we_clk [29823]));
Q_ASSIGN U2952 ( .B(clk), .A(\g.we_clk [29822]));
Q_ASSIGN U2953 ( .B(clk), .A(\g.we_clk [29821]));
Q_ASSIGN U2954 ( .B(clk), .A(\g.we_clk [29820]));
Q_ASSIGN U2955 ( .B(clk), .A(\g.we_clk [29819]));
Q_ASSIGN U2956 ( .B(clk), .A(\g.we_clk [29818]));
Q_ASSIGN U2957 ( .B(clk), .A(\g.we_clk [29817]));
Q_ASSIGN U2958 ( .B(clk), .A(\g.we_clk [29816]));
Q_ASSIGN U2959 ( .B(clk), .A(\g.we_clk [29815]));
Q_ASSIGN U2960 ( .B(clk), .A(\g.we_clk [29814]));
Q_ASSIGN U2961 ( .B(clk), .A(\g.we_clk [29813]));
Q_ASSIGN U2962 ( .B(clk), .A(\g.we_clk [29812]));
Q_ASSIGN U2963 ( .B(clk), .A(\g.we_clk [29811]));
Q_ASSIGN U2964 ( .B(clk), .A(\g.we_clk [29810]));
Q_ASSIGN U2965 ( .B(clk), .A(\g.we_clk [29809]));
Q_ASSIGN U2966 ( .B(clk), .A(\g.we_clk [29808]));
Q_ASSIGN U2967 ( .B(clk), .A(\g.we_clk [29807]));
Q_ASSIGN U2968 ( .B(clk), .A(\g.we_clk [29806]));
Q_ASSIGN U2969 ( .B(clk), .A(\g.we_clk [29805]));
Q_ASSIGN U2970 ( .B(clk), .A(\g.we_clk [29804]));
Q_ASSIGN U2971 ( .B(clk), .A(\g.we_clk [29803]));
Q_ASSIGN U2972 ( .B(clk), .A(\g.we_clk [29802]));
Q_ASSIGN U2973 ( .B(clk), .A(\g.we_clk [29801]));
Q_ASSIGN U2974 ( .B(clk), .A(\g.we_clk [29800]));
Q_ASSIGN U2975 ( .B(clk), .A(\g.we_clk [29799]));
Q_ASSIGN U2976 ( .B(clk), .A(\g.we_clk [29798]));
Q_ASSIGN U2977 ( .B(clk), .A(\g.we_clk [29797]));
Q_ASSIGN U2978 ( .B(clk), .A(\g.we_clk [29796]));
Q_ASSIGN U2979 ( .B(clk), .A(\g.we_clk [29795]));
Q_ASSIGN U2980 ( .B(clk), .A(\g.we_clk [29794]));
Q_ASSIGN U2981 ( .B(clk), .A(\g.we_clk [29793]));
Q_ASSIGN U2982 ( .B(clk), .A(\g.we_clk [29792]));
Q_ASSIGN U2983 ( .B(clk), .A(\g.we_clk [29791]));
Q_ASSIGN U2984 ( .B(clk), .A(\g.we_clk [29790]));
Q_ASSIGN U2985 ( .B(clk), .A(\g.we_clk [29789]));
Q_ASSIGN U2986 ( .B(clk), .A(\g.we_clk [29788]));
Q_ASSIGN U2987 ( .B(clk), .A(\g.we_clk [29787]));
Q_ASSIGN U2988 ( .B(clk), .A(\g.we_clk [29786]));
Q_ASSIGN U2989 ( .B(clk), .A(\g.we_clk [29785]));
Q_ASSIGN U2990 ( .B(clk), .A(\g.we_clk [29784]));
Q_ASSIGN U2991 ( .B(clk), .A(\g.we_clk [29783]));
Q_ASSIGN U2992 ( .B(clk), .A(\g.we_clk [29782]));
Q_ASSIGN U2993 ( .B(clk), .A(\g.we_clk [29781]));
Q_ASSIGN U2994 ( .B(clk), .A(\g.we_clk [29780]));
Q_ASSIGN U2995 ( .B(clk), .A(\g.we_clk [29779]));
Q_ASSIGN U2996 ( .B(clk), .A(\g.we_clk [29778]));
Q_ASSIGN U2997 ( .B(clk), .A(\g.we_clk [29777]));
Q_ASSIGN U2998 ( .B(clk), .A(\g.we_clk [29776]));
Q_ASSIGN U2999 ( .B(clk), .A(\g.we_clk [29775]));
Q_ASSIGN U3000 ( .B(clk), .A(\g.we_clk [29774]));
Q_ASSIGN U3001 ( .B(clk), .A(\g.we_clk [29773]));
Q_ASSIGN U3002 ( .B(clk), .A(\g.we_clk [29772]));
Q_ASSIGN U3003 ( .B(clk), .A(\g.we_clk [29771]));
Q_ASSIGN U3004 ( .B(clk), .A(\g.we_clk [29770]));
Q_ASSIGN U3005 ( .B(clk), .A(\g.we_clk [29769]));
Q_ASSIGN U3006 ( .B(clk), .A(\g.we_clk [29768]));
Q_ASSIGN U3007 ( .B(clk), .A(\g.we_clk [29767]));
Q_ASSIGN U3008 ( .B(clk), .A(\g.we_clk [29766]));
Q_ASSIGN U3009 ( .B(clk), .A(\g.we_clk [29765]));
Q_ASSIGN U3010 ( .B(clk), .A(\g.we_clk [29764]));
Q_ASSIGN U3011 ( .B(clk), .A(\g.we_clk [29763]));
Q_ASSIGN U3012 ( .B(clk), .A(\g.we_clk [29762]));
Q_ASSIGN U3013 ( .B(clk), .A(\g.we_clk [29761]));
Q_ASSIGN U3014 ( .B(clk), .A(\g.we_clk [29760]));
Q_ASSIGN U3015 ( .B(clk), .A(\g.we_clk [29759]));
Q_ASSIGN U3016 ( .B(clk), .A(\g.we_clk [29758]));
Q_ASSIGN U3017 ( .B(clk), .A(\g.we_clk [29757]));
Q_ASSIGN U3018 ( .B(clk), .A(\g.we_clk [29756]));
Q_ASSIGN U3019 ( .B(clk), .A(\g.we_clk [29755]));
Q_ASSIGN U3020 ( .B(clk), .A(\g.we_clk [29754]));
Q_ASSIGN U3021 ( .B(clk), .A(\g.we_clk [29753]));
Q_ASSIGN U3022 ( .B(clk), .A(\g.we_clk [29752]));
Q_ASSIGN U3023 ( .B(clk), .A(\g.we_clk [29751]));
Q_ASSIGN U3024 ( .B(clk), .A(\g.we_clk [29750]));
Q_ASSIGN U3025 ( .B(clk), .A(\g.we_clk [29749]));
Q_ASSIGN U3026 ( .B(clk), .A(\g.we_clk [29748]));
Q_ASSIGN U3027 ( .B(clk), .A(\g.we_clk [29747]));
Q_ASSIGN U3028 ( .B(clk), .A(\g.we_clk [29746]));
Q_ASSIGN U3029 ( .B(clk), .A(\g.we_clk [29745]));
Q_ASSIGN U3030 ( .B(clk), .A(\g.we_clk [29744]));
Q_ASSIGN U3031 ( .B(clk), .A(\g.we_clk [29743]));
Q_ASSIGN U3032 ( .B(clk), .A(\g.we_clk [29742]));
Q_ASSIGN U3033 ( .B(clk), .A(\g.we_clk [29741]));
Q_ASSIGN U3034 ( .B(clk), .A(\g.we_clk [29740]));
Q_ASSIGN U3035 ( .B(clk), .A(\g.we_clk [29739]));
Q_ASSIGN U3036 ( .B(clk), .A(\g.we_clk [29738]));
Q_ASSIGN U3037 ( .B(clk), .A(\g.we_clk [29737]));
Q_ASSIGN U3038 ( .B(clk), .A(\g.we_clk [29736]));
Q_ASSIGN U3039 ( .B(clk), .A(\g.we_clk [29735]));
Q_ASSIGN U3040 ( .B(clk), .A(\g.we_clk [29734]));
Q_ASSIGN U3041 ( .B(clk), .A(\g.we_clk [29733]));
Q_ASSIGN U3042 ( .B(clk), .A(\g.we_clk [29732]));
Q_ASSIGN U3043 ( .B(clk), .A(\g.we_clk [29731]));
Q_ASSIGN U3044 ( .B(clk), .A(\g.we_clk [29730]));
Q_ASSIGN U3045 ( .B(clk), .A(\g.we_clk [29729]));
Q_ASSIGN U3046 ( .B(clk), .A(\g.we_clk [29728]));
Q_ASSIGN U3047 ( .B(clk), .A(\g.we_clk [29727]));
Q_ASSIGN U3048 ( .B(clk), .A(\g.we_clk [29726]));
Q_ASSIGN U3049 ( .B(clk), .A(\g.we_clk [29725]));
Q_ASSIGN U3050 ( .B(clk), .A(\g.we_clk [29724]));
Q_ASSIGN U3051 ( .B(clk), .A(\g.we_clk [29723]));
Q_ASSIGN U3052 ( .B(clk), .A(\g.we_clk [29722]));
Q_ASSIGN U3053 ( .B(clk), .A(\g.we_clk [29721]));
Q_ASSIGN U3054 ( .B(clk), .A(\g.we_clk [29720]));
Q_ASSIGN U3055 ( .B(clk), .A(\g.we_clk [29719]));
Q_ASSIGN U3056 ( .B(clk), .A(\g.we_clk [29718]));
Q_ASSIGN U3057 ( .B(clk), .A(\g.we_clk [29717]));
Q_ASSIGN U3058 ( .B(clk), .A(\g.we_clk [29716]));
Q_ASSIGN U3059 ( .B(clk), .A(\g.we_clk [29715]));
Q_ASSIGN U3060 ( .B(clk), .A(\g.we_clk [29714]));
Q_ASSIGN U3061 ( .B(clk), .A(\g.we_clk [29713]));
Q_ASSIGN U3062 ( .B(clk), .A(\g.we_clk [29712]));
Q_ASSIGN U3063 ( .B(clk), .A(\g.we_clk [29711]));
Q_ASSIGN U3064 ( .B(clk), .A(\g.we_clk [29710]));
Q_ASSIGN U3065 ( .B(clk), .A(\g.we_clk [29709]));
Q_ASSIGN U3066 ( .B(clk), .A(\g.we_clk [29708]));
Q_ASSIGN U3067 ( .B(clk), .A(\g.we_clk [29707]));
Q_ASSIGN U3068 ( .B(clk), .A(\g.we_clk [29706]));
Q_ASSIGN U3069 ( .B(clk), .A(\g.we_clk [29705]));
Q_ASSIGN U3070 ( .B(clk), .A(\g.we_clk [29704]));
Q_ASSIGN U3071 ( .B(clk), .A(\g.we_clk [29703]));
Q_ASSIGN U3072 ( .B(clk), .A(\g.we_clk [29702]));
Q_ASSIGN U3073 ( .B(clk), .A(\g.we_clk [29701]));
Q_ASSIGN U3074 ( .B(clk), .A(\g.we_clk [29700]));
Q_ASSIGN U3075 ( .B(clk), .A(\g.we_clk [29699]));
Q_ASSIGN U3076 ( .B(clk), .A(\g.we_clk [29698]));
Q_ASSIGN U3077 ( .B(clk), .A(\g.we_clk [29697]));
Q_ASSIGN U3078 ( .B(clk), .A(\g.we_clk [29696]));
Q_ASSIGN U3079 ( .B(clk), .A(\g.we_clk [29695]));
Q_ASSIGN U3080 ( .B(clk), .A(\g.we_clk [29694]));
Q_ASSIGN U3081 ( .B(clk), .A(\g.we_clk [29693]));
Q_ASSIGN U3082 ( .B(clk), .A(\g.we_clk [29692]));
Q_ASSIGN U3083 ( .B(clk), .A(\g.we_clk [29691]));
Q_ASSIGN U3084 ( .B(clk), .A(\g.we_clk [29690]));
Q_ASSIGN U3085 ( .B(clk), .A(\g.we_clk [29689]));
Q_ASSIGN U3086 ( .B(clk), .A(\g.we_clk [29688]));
Q_ASSIGN U3087 ( .B(clk), .A(\g.we_clk [29687]));
Q_ASSIGN U3088 ( .B(clk), .A(\g.we_clk [29686]));
Q_ASSIGN U3089 ( .B(clk), .A(\g.we_clk [29685]));
Q_ASSIGN U3090 ( .B(clk), .A(\g.we_clk [29684]));
Q_ASSIGN U3091 ( .B(clk), .A(\g.we_clk [29683]));
Q_ASSIGN U3092 ( .B(clk), .A(\g.we_clk [29682]));
Q_ASSIGN U3093 ( .B(clk), .A(\g.we_clk [29681]));
Q_ASSIGN U3094 ( .B(clk), .A(\g.we_clk [29680]));
Q_ASSIGN U3095 ( .B(clk), .A(\g.we_clk [29679]));
Q_ASSIGN U3096 ( .B(clk), .A(\g.we_clk [29678]));
Q_ASSIGN U3097 ( .B(clk), .A(\g.we_clk [29677]));
Q_ASSIGN U3098 ( .B(clk), .A(\g.we_clk [29676]));
Q_ASSIGN U3099 ( .B(clk), .A(\g.we_clk [29675]));
Q_ASSIGN U3100 ( .B(clk), .A(\g.we_clk [29674]));
Q_ASSIGN U3101 ( .B(clk), .A(\g.we_clk [29673]));
Q_ASSIGN U3102 ( .B(clk), .A(\g.we_clk [29672]));
Q_ASSIGN U3103 ( .B(clk), .A(\g.we_clk [29671]));
Q_ASSIGN U3104 ( .B(clk), .A(\g.we_clk [29670]));
Q_ASSIGN U3105 ( .B(clk), .A(\g.we_clk [29669]));
Q_ASSIGN U3106 ( .B(clk), .A(\g.we_clk [29668]));
Q_ASSIGN U3107 ( .B(clk), .A(\g.we_clk [29667]));
Q_ASSIGN U3108 ( .B(clk), .A(\g.we_clk [29666]));
Q_ASSIGN U3109 ( .B(clk), .A(\g.we_clk [29665]));
Q_ASSIGN U3110 ( .B(clk), .A(\g.we_clk [29664]));
Q_ASSIGN U3111 ( .B(clk), .A(\g.we_clk [29663]));
Q_ASSIGN U3112 ( .B(clk), .A(\g.we_clk [29662]));
Q_ASSIGN U3113 ( .B(clk), .A(\g.we_clk [29661]));
Q_ASSIGN U3114 ( .B(clk), .A(\g.we_clk [29660]));
Q_ASSIGN U3115 ( .B(clk), .A(\g.we_clk [29659]));
Q_ASSIGN U3116 ( .B(clk), .A(\g.we_clk [29658]));
Q_ASSIGN U3117 ( .B(clk), .A(\g.we_clk [29657]));
Q_ASSIGN U3118 ( .B(clk), .A(\g.we_clk [29656]));
Q_ASSIGN U3119 ( .B(clk), .A(\g.we_clk [29655]));
Q_ASSIGN U3120 ( .B(clk), .A(\g.we_clk [29654]));
Q_ASSIGN U3121 ( .B(clk), .A(\g.we_clk [29653]));
Q_ASSIGN U3122 ( .B(clk), .A(\g.we_clk [29652]));
Q_ASSIGN U3123 ( .B(clk), .A(\g.we_clk [29651]));
Q_ASSIGN U3124 ( .B(clk), .A(\g.we_clk [29650]));
Q_ASSIGN U3125 ( .B(clk), .A(\g.we_clk [29649]));
Q_ASSIGN U3126 ( .B(clk), .A(\g.we_clk [29648]));
Q_ASSIGN U3127 ( .B(clk), .A(\g.we_clk [29647]));
Q_ASSIGN U3128 ( .B(clk), .A(\g.we_clk [29646]));
Q_ASSIGN U3129 ( .B(clk), .A(\g.we_clk [29645]));
Q_ASSIGN U3130 ( .B(clk), .A(\g.we_clk [29644]));
Q_ASSIGN U3131 ( .B(clk), .A(\g.we_clk [29643]));
Q_ASSIGN U3132 ( .B(clk), .A(\g.we_clk [29642]));
Q_ASSIGN U3133 ( .B(clk), .A(\g.we_clk [29641]));
Q_ASSIGN U3134 ( .B(clk), .A(\g.we_clk [29640]));
Q_ASSIGN U3135 ( .B(clk), .A(\g.we_clk [29639]));
Q_ASSIGN U3136 ( .B(clk), .A(\g.we_clk [29638]));
Q_ASSIGN U3137 ( .B(clk), .A(\g.we_clk [29637]));
Q_ASSIGN U3138 ( .B(clk), .A(\g.we_clk [29636]));
Q_ASSIGN U3139 ( .B(clk), .A(\g.we_clk [29635]));
Q_ASSIGN U3140 ( .B(clk), .A(\g.we_clk [29634]));
Q_ASSIGN U3141 ( .B(clk), .A(\g.we_clk [29633]));
Q_ASSIGN U3142 ( .B(clk), .A(\g.we_clk [29632]));
Q_ASSIGN U3143 ( .B(clk), .A(\g.we_clk [29631]));
Q_ASSIGN U3144 ( .B(clk), .A(\g.we_clk [29630]));
Q_ASSIGN U3145 ( .B(clk), .A(\g.we_clk [29629]));
Q_ASSIGN U3146 ( .B(clk), .A(\g.we_clk [29628]));
Q_ASSIGN U3147 ( .B(clk), .A(\g.we_clk [29627]));
Q_ASSIGN U3148 ( .B(clk), .A(\g.we_clk [29626]));
Q_ASSIGN U3149 ( .B(clk), .A(\g.we_clk [29625]));
Q_ASSIGN U3150 ( .B(clk), .A(\g.we_clk [29624]));
Q_ASSIGN U3151 ( .B(clk), .A(\g.we_clk [29623]));
Q_ASSIGN U3152 ( .B(clk), .A(\g.we_clk [29622]));
Q_ASSIGN U3153 ( .B(clk), .A(\g.we_clk [29621]));
Q_ASSIGN U3154 ( .B(clk), .A(\g.we_clk [29620]));
Q_ASSIGN U3155 ( .B(clk), .A(\g.we_clk [29619]));
Q_ASSIGN U3156 ( .B(clk), .A(\g.we_clk [29618]));
Q_ASSIGN U3157 ( .B(clk), .A(\g.we_clk [29617]));
Q_ASSIGN U3158 ( .B(clk), .A(\g.we_clk [29616]));
Q_ASSIGN U3159 ( .B(clk), .A(\g.we_clk [29615]));
Q_ASSIGN U3160 ( .B(clk), .A(\g.we_clk [29614]));
Q_ASSIGN U3161 ( .B(clk), .A(\g.we_clk [29613]));
Q_ASSIGN U3162 ( .B(clk), .A(\g.we_clk [29612]));
Q_ASSIGN U3163 ( .B(clk), .A(\g.we_clk [29611]));
Q_ASSIGN U3164 ( .B(clk), .A(\g.we_clk [29610]));
Q_ASSIGN U3165 ( .B(clk), .A(\g.we_clk [29609]));
Q_ASSIGN U3166 ( .B(clk), .A(\g.we_clk [29608]));
Q_ASSIGN U3167 ( .B(clk), .A(\g.we_clk [29607]));
Q_ASSIGN U3168 ( .B(clk), .A(\g.we_clk [29606]));
Q_ASSIGN U3169 ( .B(clk), .A(\g.we_clk [29605]));
Q_ASSIGN U3170 ( .B(clk), .A(\g.we_clk [29604]));
Q_ASSIGN U3171 ( .B(clk), .A(\g.we_clk [29603]));
Q_ASSIGN U3172 ( .B(clk), .A(\g.we_clk [29602]));
Q_ASSIGN U3173 ( .B(clk), .A(\g.we_clk [29601]));
Q_ASSIGN U3174 ( .B(clk), .A(\g.we_clk [29600]));
Q_ASSIGN U3175 ( .B(clk), .A(\g.we_clk [29599]));
Q_ASSIGN U3176 ( .B(clk), .A(\g.we_clk [29598]));
Q_ASSIGN U3177 ( .B(clk), .A(\g.we_clk [29597]));
Q_ASSIGN U3178 ( .B(clk), .A(\g.we_clk [29596]));
Q_ASSIGN U3179 ( .B(clk), .A(\g.we_clk [29595]));
Q_ASSIGN U3180 ( .B(clk), .A(\g.we_clk [29594]));
Q_ASSIGN U3181 ( .B(clk), .A(\g.we_clk [29593]));
Q_ASSIGN U3182 ( .B(clk), .A(\g.we_clk [29592]));
Q_ASSIGN U3183 ( .B(clk), .A(\g.we_clk [29591]));
Q_ASSIGN U3184 ( .B(clk), .A(\g.we_clk [29590]));
Q_ASSIGN U3185 ( .B(clk), .A(\g.we_clk [29589]));
Q_ASSIGN U3186 ( .B(clk), .A(\g.we_clk [29588]));
Q_ASSIGN U3187 ( .B(clk), .A(\g.we_clk [29587]));
Q_ASSIGN U3188 ( .B(clk), .A(\g.we_clk [29586]));
Q_ASSIGN U3189 ( .B(clk), .A(\g.we_clk [29585]));
Q_ASSIGN U3190 ( .B(clk), .A(\g.we_clk [29584]));
Q_ASSIGN U3191 ( .B(clk), .A(\g.we_clk [29583]));
Q_ASSIGN U3192 ( .B(clk), .A(\g.we_clk [29582]));
Q_ASSIGN U3193 ( .B(clk), .A(\g.we_clk [29581]));
Q_ASSIGN U3194 ( .B(clk), .A(\g.we_clk [29580]));
Q_ASSIGN U3195 ( .B(clk), .A(\g.we_clk [29579]));
Q_ASSIGN U3196 ( .B(clk), .A(\g.we_clk [29578]));
Q_ASSIGN U3197 ( .B(clk), .A(\g.we_clk [29577]));
Q_ASSIGN U3198 ( .B(clk), .A(\g.we_clk [29576]));
Q_ASSIGN U3199 ( .B(clk), .A(\g.we_clk [29575]));
Q_ASSIGN U3200 ( .B(clk), .A(\g.we_clk [29574]));
Q_ASSIGN U3201 ( .B(clk), .A(\g.we_clk [29573]));
Q_ASSIGN U3202 ( .B(clk), .A(\g.we_clk [29572]));
Q_ASSIGN U3203 ( .B(clk), .A(\g.we_clk [29571]));
Q_ASSIGN U3204 ( .B(clk), .A(\g.we_clk [29570]));
Q_ASSIGN U3205 ( .B(clk), .A(\g.we_clk [29569]));
Q_ASSIGN U3206 ( .B(clk), .A(\g.we_clk [29568]));
Q_ASSIGN U3207 ( .B(clk), .A(\g.we_clk [29567]));
Q_ASSIGN U3208 ( .B(clk), .A(\g.we_clk [29566]));
Q_ASSIGN U3209 ( .B(clk), .A(\g.we_clk [29565]));
Q_ASSIGN U3210 ( .B(clk), .A(\g.we_clk [29564]));
Q_ASSIGN U3211 ( .B(clk), .A(\g.we_clk [29563]));
Q_ASSIGN U3212 ( .B(clk), .A(\g.we_clk [29562]));
Q_ASSIGN U3213 ( .B(clk), .A(\g.we_clk [29561]));
Q_ASSIGN U3214 ( .B(clk), .A(\g.we_clk [29560]));
Q_ASSIGN U3215 ( .B(clk), .A(\g.we_clk [29559]));
Q_ASSIGN U3216 ( .B(clk), .A(\g.we_clk [29558]));
Q_ASSIGN U3217 ( .B(clk), .A(\g.we_clk [29557]));
Q_ASSIGN U3218 ( .B(clk), .A(\g.we_clk [29556]));
Q_ASSIGN U3219 ( .B(clk), .A(\g.we_clk [29555]));
Q_ASSIGN U3220 ( .B(clk), .A(\g.we_clk [29554]));
Q_ASSIGN U3221 ( .B(clk), .A(\g.we_clk [29553]));
Q_ASSIGN U3222 ( .B(clk), .A(\g.we_clk [29552]));
Q_ASSIGN U3223 ( .B(clk), .A(\g.we_clk [29551]));
Q_ASSIGN U3224 ( .B(clk), .A(\g.we_clk [29550]));
Q_ASSIGN U3225 ( .B(clk), .A(\g.we_clk [29549]));
Q_ASSIGN U3226 ( .B(clk), .A(\g.we_clk [29548]));
Q_ASSIGN U3227 ( .B(clk), .A(\g.we_clk [29547]));
Q_ASSIGN U3228 ( .B(clk), .A(\g.we_clk [29546]));
Q_ASSIGN U3229 ( .B(clk), .A(\g.we_clk [29545]));
Q_ASSIGN U3230 ( .B(clk), .A(\g.we_clk [29544]));
Q_ASSIGN U3231 ( .B(clk), .A(\g.we_clk [29543]));
Q_ASSIGN U3232 ( .B(clk), .A(\g.we_clk [29542]));
Q_ASSIGN U3233 ( .B(clk), .A(\g.we_clk [29541]));
Q_ASSIGN U3234 ( .B(clk), .A(\g.we_clk [29540]));
Q_ASSIGN U3235 ( .B(clk), .A(\g.we_clk [29539]));
Q_ASSIGN U3236 ( .B(clk), .A(\g.we_clk [29538]));
Q_ASSIGN U3237 ( .B(clk), .A(\g.we_clk [29537]));
Q_ASSIGN U3238 ( .B(clk), .A(\g.we_clk [29536]));
Q_ASSIGN U3239 ( .B(clk), .A(\g.we_clk [29535]));
Q_ASSIGN U3240 ( .B(clk), .A(\g.we_clk [29534]));
Q_ASSIGN U3241 ( .B(clk), .A(\g.we_clk [29533]));
Q_ASSIGN U3242 ( .B(clk), .A(\g.we_clk [29532]));
Q_ASSIGN U3243 ( .B(clk), .A(\g.we_clk [29531]));
Q_ASSIGN U3244 ( .B(clk), .A(\g.we_clk [29530]));
Q_ASSIGN U3245 ( .B(clk), .A(\g.we_clk [29529]));
Q_ASSIGN U3246 ( .B(clk), .A(\g.we_clk [29528]));
Q_ASSIGN U3247 ( .B(clk), .A(\g.we_clk [29527]));
Q_ASSIGN U3248 ( .B(clk), .A(\g.we_clk [29526]));
Q_ASSIGN U3249 ( .B(clk), .A(\g.we_clk [29525]));
Q_ASSIGN U3250 ( .B(clk), .A(\g.we_clk [29524]));
Q_ASSIGN U3251 ( .B(clk), .A(\g.we_clk [29523]));
Q_ASSIGN U3252 ( .B(clk), .A(\g.we_clk [29522]));
Q_ASSIGN U3253 ( .B(clk), .A(\g.we_clk [29521]));
Q_ASSIGN U3254 ( .B(clk), .A(\g.we_clk [29520]));
Q_ASSIGN U3255 ( .B(clk), .A(\g.we_clk [29519]));
Q_ASSIGN U3256 ( .B(clk), .A(\g.we_clk [29518]));
Q_ASSIGN U3257 ( .B(clk), .A(\g.we_clk [29517]));
Q_ASSIGN U3258 ( .B(clk), .A(\g.we_clk [29516]));
Q_ASSIGN U3259 ( .B(clk), .A(\g.we_clk [29515]));
Q_ASSIGN U3260 ( .B(clk), .A(\g.we_clk [29514]));
Q_ASSIGN U3261 ( .B(clk), .A(\g.we_clk [29513]));
Q_ASSIGN U3262 ( .B(clk), .A(\g.we_clk [29512]));
Q_ASSIGN U3263 ( .B(clk), .A(\g.we_clk [29511]));
Q_ASSIGN U3264 ( .B(clk), .A(\g.we_clk [29510]));
Q_ASSIGN U3265 ( .B(clk), .A(\g.we_clk [29509]));
Q_ASSIGN U3266 ( .B(clk), .A(\g.we_clk [29508]));
Q_ASSIGN U3267 ( .B(clk), .A(\g.we_clk [29507]));
Q_ASSIGN U3268 ( .B(clk), .A(\g.we_clk [29506]));
Q_ASSIGN U3269 ( .B(clk), .A(\g.we_clk [29505]));
Q_ASSIGN U3270 ( .B(clk), .A(\g.we_clk [29504]));
Q_ASSIGN U3271 ( .B(clk), .A(\g.we_clk [29503]));
Q_ASSIGN U3272 ( .B(clk), .A(\g.we_clk [29502]));
Q_ASSIGN U3273 ( .B(clk), .A(\g.we_clk [29501]));
Q_ASSIGN U3274 ( .B(clk), .A(\g.we_clk [29500]));
Q_ASSIGN U3275 ( .B(clk), .A(\g.we_clk [29499]));
Q_ASSIGN U3276 ( .B(clk), .A(\g.we_clk [29498]));
Q_ASSIGN U3277 ( .B(clk), .A(\g.we_clk [29497]));
Q_ASSIGN U3278 ( .B(clk), .A(\g.we_clk [29496]));
Q_ASSIGN U3279 ( .B(clk), .A(\g.we_clk [29495]));
Q_ASSIGN U3280 ( .B(clk), .A(\g.we_clk [29494]));
Q_ASSIGN U3281 ( .B(clk), .A(\g.we_clk [29493]));
Q_ASSIGN U3282 ( .B(clk), .A(\g.we_clk [29492]));
Q_ASSIGN U3283 ( .B(clk), .A(\g.we_clk [29491]));
Q_ASSIGN U3284 ( .B(clk), .A(\g.we_clk [29490]));
Q_ASSIGN U3285 ( .B(clk), .A(\g.we_clk [29489]));
Q_ASSIGN U3286 ( .B(clk), .A(\g.we_clk [29488]));
Q_ASSIGN U3287 ( .B(clk), .A(\g.we_clk [29487]));
Q_ASSIGN U3288 ( .B(clk), .A(\g.we_clk [29486]));
Q_ASSIGN U3289 ( .B(clk), .A(\g.we_clk [29485]));
Q_ASSIGN U3290 ( .B(clk), .A(\g.we_clk [29484]));
Q_ASSIGN U3291 ( .B(clk), .A(\g.we_clk [29483]));
Q_ASSIGN U3292 ( .B(clk), .A(\g.we_clk [29482]));
Q_ASSIGN U3293 ( .B(clk), .A(\g.we_clk [29481]));
Q_ASSIGN U3294 ( .B(clk), .A(\g.we_clk [29480]));
Q_ASSIGN U3295 ( .B(clk), .A(\g.we_clk [29479]));
Q_ASSIGN U3296 ( .B(clk), .A(\g.we_clk [29478]));
Q_ASSIGN U3297 ( .B(clk), .A(\g.we_clk [29477]));
Q_ASSIGN U3298 ( .B(clk), .A(\g.we_clk [29476]));
Q_ASSIGN U3299 ( .B(clk), .A(\g.we_clk [29475]));
Q_ASSIGN U3300 ( .B(clk), .A(\g.we_clk [29474]));
Q_ASSIGN U3301 ( .B(clk), .A(\g.we_clk [29473]));
Q_ASSIGN U3302 ( .B(clk), .A(\g.we_clk [29472]));
Q_ASSIGN U3303 ( .B(clk), .A(\g.we_clk [29471]));
Q_ASSIGN U3304 ( .B(clk), .A(\g.we_clk [29470]));
Q_ASSIGN U3305 ( .B(clk), .A(\g.we_clk [29469]));
Q_ASSIGN U3306 ( .B(clk), .A(\g.we_clk [29468]));
Q_ASSIGN U3307 ( .B(clk), .A(\g.we_clk [29467]));
Q_ASSIGN U3308 ( .B(clk), .A(\g.we_clk [29466]));
Q_ASSIGN U3309 ( .B(clk), .A(\g.we_clk [29465]));
Q_ASSIGN U3310 ( .B(clk), .A(\g.we_clk [29464]));
Q_ASSIGN U3311 ( .B(clk), .A(\g.we_clk [29463]));
Q_ASSIGN U3312 ( .B(clk), .A(\g.we_clk [29462]));
Q_ASSIGN U3313 ( .B(clk), .A(\g.we_clk [29461]));
Q_ASSIGN U3314 ( .B(clk), .A(\g.we_clk [29460]));
Q_ASSIGN U3315 ( .B(clk), .A(\g.we_clk [29459]));
Q_ASSIGN U3316 ( .B(clk), .A(\g.we_clk [29458]));
Q_ASSIGN U3317 ( .B(clk), .A(\g.we_clk [29457]));
Q_ASSIGN U3318 ( .B(clk), .A(\g.we_clk [29456]));
Q_ASSIGN U3319 ( .B(clk), .A(\g.we_clk [29455]));
Q_ASSIGN U3320 ( .B(clk), .A(\g.we_clk [29454]));
Q_ASSIGN U3321 ( .B(clk), .A(\g.we_clk [29453]));
Q_ASSIGN U3322 ( .B(clk), .A(\g.we_clk [29452]));
Q_ASSIGN U3323 ( .B(clk), .A(\g.we_clk [29451]));
Q_ASSIGN U3324 ( .B(clk), .A(\g.we_clk [29450]));
Q_ASSIGN U3325 ( .B(clk), .A(\g.we_clk [29449]));
Q_ASSIGN U3326 ( .B(clk), .A(\g.we_clk [29448]));
Q_ASSIGN U3327 ( .B(clk), .A(\g.we_clk [29447]));
Q_ASSIGN U3328 ( .B(clk), .A(\g.we_clk [29446]));
Q_ASSIGN U3329 ( .B(clk), .A(\g.we_clk [29445]));
Q_ASSIGN U3330 ( .B(clk), .A(\g.we_clk [29444]));
Q_ASSIGN U3331 ( .B(clk), .A(\g.we_clk [29443]));
Q_ASSIGN U3332 ( .B(clk), .A(\g.we_clk [29442]));
Q_ASSIGN U3333 ( .B(clk), .A(\g.we_clk [29441]));
Q_ASSIGN U3334 ( .B(clk), .A(\g.we_clk [29440]));
Q_ASSIGN U3335 ( .B(clk), .A(\g.we_clk [29439]));
Q_ASSIGN U3336 ( .B(clk), .A(\g.we_clk [29438]));
Q_ASSIGN U3337 ( .B(clk), .A(\g.we_clk [29437]));
Q_ASSIGN U3338 ( .B(clk), .A(\g.we_clk [29436]));
Q_ASSIGN U3339 ( .B(clk), .A(\g.we_clk [29435]));
Q_ASSIGN U3340 ( .B(clk), .A(\g.we_clk [29434]));
Q_ASSIGN U3341 ( .B(clk), .A(\g.we_clk [29433]));
Q_ASSIGN U3342 ( .B(clk), .A(\g.we_clk [29432]));
Q_ASSIGN U3343 ( .B(clk), .A(\g.we_clk [29431]));
Q_ASSIGN U3344 ( .B(clk), .A(\g.we_clk [29430]));
Q_ASSIGN U3345 ( .B(clk), .A(\g.we_clk [29429]));
Q_ASSIGN U3346 ( .B(clk), .A(\g.we_clk [29428]));
Q_ASSIGN U3347 ( .B(clk), .A(\g.we_clk [29427]));
Q_ASSIGN U3348 ( .B(clk), .A(\g.we_clk [29426]));
Q_ASSIGN U3349 ( .B(clk), .A(\g.we_clk [29425]));
Q_ASSIGN U3350 ( .B(clk), .A(\g.we_clk [29424]));
Q_ASSIGN U3351 ( .B(clk), .A(\g.we_clk [29423]));
Q_ASSIGN U3352 ( .B(clk), .A(\g.we_clk [29422]));
Q_ASSIGN U3353 ( .B(clk), .A(\g.we_clk [29421]));
Q_ASSIGN U3354 ( .B(clk), .A(\g.we_clk [29420]));
Q_ASSIGN U3355 ( .B(clk), .A(\g.we_clk [29419]));
Q_ASSIGN U3356 ( .B(clk), .A(\g.we_clk [29418]));
Q_ASSIGN U3357 ( .B(clk), .A(\g.we_clk [29417]));
Q_ASSIGN U3358 ( .B(clk), .A(\g.we_clk [29416]));
Q_ASSIGN U3359 ( .B(clk), .A(\g.we_clk [29415]));
Q_ASSIGN U3360 ( .B(clk), .A(\g.we_clk [29414]));
Q_ASSIGN U3361 ( .B(clk), .A(\g.we_clk [29413]));
Q_ASSIGN U3362 ( .B(clk), .A(\g.we_clk [29412]));
Q_ASSIGN U3363 ( .B(clk), .A(\g.we_clk [29411]));
Q_ASSIGN U3364 ( .B(clk), .A(\g.we_clk [29410]));
Q_ASSIGN U3365 ( .B(clk), .A(\g.we_clk [29409]));
Q_ASSIGN U3366 ( .B(clk), .A(\g.we_clk [29408]));
Q_ASSIGN U3367 ( .B(clk), .A(\g.we_clk [29407]));
Q_ASSIGN U3368 ( .B(clk), .A(\g.we_clk [29406]));
Q_ASSIGN U3369 ( .B(clk), .A(\g.we_clk [29405]));
Q_ASSIGN U3370 ( .B(clk), .A(\g.we_clk [29404]));
Q_ASSIGN U3371 ( .B(clk), .A(\g.we_clk [29403]));
Q_ASSIGN U3372 ( .B(clk), .A(\g.we_clk [29402]));
Q_ASSIGN U3373 ( .B(clk), .A(\g.we_clk [29401]));
Q_ASSIGN U3374 ( .B(clk), .A(\g.we_clk [29400]));
Q_ASSIGN U3375 ( .B(clk), .A(\g.we_clk [29399]));
Q_ASSIGN U3376 ( .B(clk), .A(\g.we_clk [29398]));
Q_ASSIGN U3377 ( .B(clk), .A(\g.we_clk [29397]));
Q_ASSIGN U3378 ( .B(clk), .A(\g.we_clk [29396]));
Q_ASSIGN U3379 ( .B(clk), .A(\g.we_clk [29395]));
Q_ASSIGN U3380 ( .B(clk), .A(\g.we_clk [29394]));
Q_ASSIGN U3381 ( .B(clk), .A(\g.we_clk [29393]));
Q_ASSIGN U3382 ( .B(clk), .A(\g.we_clk [29392]));
Q_ASSIGN U3383 ( .B(clk), .A(\g.we_clk [29391]));
Q_ASSIGN U3384 ( .B(clk), .A(\g.we_clk [29390]));
Q_ASSIGN U3385 ( .B(clk), .A(\g.we_clk [29389]));
Q_ASSIGN U3386 ( .B(clk), .A(\g.we_clk [29388]));
Q_ASSIGN U3387 ( .B(clk), .A(\g.we_clk [29387]));
Q_ASSIGN U3388 ( .B(clk), .A(\g.we_clk [29386]));
Q_ASSIGN U3389 ( .B(clk), .A(\g.we_clk [29385]));
Q_ASSIGN U3390 ( .B(clk), .A(\g.we_clk [29384]));
Q_ASSIGN U3391 ( .B(clk), .A(\g.we_clk [29383]));
Q_ASSIGN U3392 ( .B(clk), .A(\g.we_clk [29382]));
Q_ASSIGN U3393 ( .B(clk), .A(\g.we_clk [29381]));
Q_ASSIGN U3394 ( .B(clk), .A(\g.we_clk [29380]));
Q_ASSIGN U3395 ( .B(clk), .A(\g.we_clk [29379]));
Q_ASSIGN U3396 ( .B(clk), .A(\g.we_clk [29378]));
Q_ASSIGN U3397 ( .B(clk), .A(\g.we_clk [29377]));
Q_ASSIGN U3398 ( .B(clk), .A(\g.we_clk [29376]));
Q_ASSIGN U3399 ( .B(clk), .A(\g.we_clk [29375]));
Q_ASSIGN U3400 ( .B(clk), .A(\g.we_clk [29374]));
Q_ASSIGN U3401 ( .B(clk), .A(\g.we_clk [29373]));
Q_ASSIGN U3402 ( .B(clk), .A(\g.we_clk [29372]));
Q_ASSIGN U3403 ( .B(clk), .A(\g.we_clk [29371]));
Q_ASSIGN U3404 ( .B(clk), .A(\g.we_clk [29370]));
Q_ASSIGN U3405 ( .B(clk), .A(\g.we_clk [29369]));
Q_ASSIGN U3406 ( .B(clk), .A(\g.we_clk [29368]));
Q_ASSIGN U3407 ( .B(clk), .A(\g.we_clk [29367]));
Q_ASSIGN U3408 ( .B(clk), .A(\g.we_clk [29366]));
Q_ASSIGN U3409 ( .B(clk), .A(\g.we_clk [29365]));
Q_ASSIGN U3410 ( .B(clk), .A(\g.we_clk [29364]));
Q_ASSIGN U3411 ( .B(clk), .A(\g.we_clk [29363]));
Q_ASSIGN U3412 ( .B(clk), .A(\g.we_clk [29362]));
Q_ASSIGN U3413 ( .B(clk), .A(\g.we_clk [29361]));
Q_ASSIGN U3414 ( .B(clk), .A(\g.we_clk [29360]));
Q_ASSIGN U3415 ( .B(clk), .A(\g.we_clk [29359]));
Q_ASSIGN U3416 ( .B(clk), .A(\g.we_clk [29358]));
Q_ASSIGN U3417 ( .B(clk), .A(\g.we_clk [29357]));
Q_ASSIGN U3418 ( .B(clk), .A(\g.we_clk [29356]));
Q_ASSIGN U3419 ( .B(clk), .A(\g.we_clk [29355]));
Q_ASSIGN U3420 ( .B(clk), .A(\g.we_clk [29354]));
Q_ASSIGN U3421 ( .B(clk), .A(\g.we_clk [29353]));
Q_ASSIGN U3422 ( .B(clk), .A(\g.we_clk [29352]));
Q_ASSIGN U3423 ( .B(clk), .A(\g.we_clk [29351]));
Q_ASSIGN U3424 ( .B(clk), .A(\g.we_clk [29350]));
Q_ASSIGN U3425 ( .B(clk), .A(\g.we_clk [29349]));
Q_ASSIGN U3426 ( .B(clk), .A(\g.we_clk [29348]));
Q_ASSIGN U3427 ( .B(clk), .A(\g.we_clk [29347]));
Q_ASSIGN U3428 ( .B(clk), .A(\g.we_clk [29346]));
Q_ASSIGN U3429 ( .B(clk), .A(\g.we_clk [29345]));
Q_ASSIGN U3430 ( .B(clk), .A(\g.we_clk [29344]));
Q_ASSIGN U3431 ( .B(clk), .A(\g.we_clk [29343]));
Q_ASSIGN U3432 ( .B(clk), .A(\g.we_clk [29342]));
Q_ASSIGN U3433 ( .B(clk), .A(\g.we_clk [29341]));
Q_ASSIGN U3434 ( .B(clk), .A(\g.we_clk [29340]));
Q_ASSIGN U3435 ( .B(clk), .A(\g.we_clk [29339]));
Q_ASSIGN U3436 ( .B(clk), .A(\g.we_clk [29338]));
Q_ASSIGN U3437 ( .B(clk), .A(\g.we_clk [29337]));
Q_ASSIGN U3438 ( .B(clk), .A(\g.we_clk [29336]));
Q_ASSIGN U3439 ( .B(clk), .A(\g.we_clk [29335]));
Q_ASSIGN U3440 ( .B(clk), .A(\g.we_clk [29334]));
Q_ASSIGN U3441 ( .B(clk), .A(\g.we_clk [29333]));
Q_ASSIGN U3442 ( .B(clk), .A(\g.we_clk [29332]));
Q_ASSIGN U3443 ( .B(clk), .A(\g.we_clk [29331]));
Q_ASSIGN U3444 ( .B(clk), .A(\g.we_clk [29330]));
Q_ASSIGN U3445 ( .B(clk), .A(\g.we_clk [29329]));
Q_ASSIGN U3446 ( .B(clk), .A(\g.we_clk [29328]));
Q_ASSIGN U3447 ( .B(clk), .A(\g.we_clk [29327]));
Q_ASSIGN U3448 ( .B(clk), .A(\g.we_clk [29326]));
Q_ASSIGN U3449 ( .B(clk), .A(\g.we_clk [29325]));
Q_ASSIGN U3450 ( .B(clk), .A(\g.we_clk [29324]));
Q_ASSIGN U3451 ( .B(clk), .A(\g.we_clk [29323]));
Q_ASSIGN U3452 ( .B(clk), .A(\g.we_clk [29322]));
Q_ASSIGN U3453 ( .B(clk), .A(\g.we_clk [29321]));
Q_ASSIGN U3454 ( .B(clk), .A(\g.we_clk [29320]));
Q_ASSIGN U3455 ( .B(clk), .A(\g.we_clk [29319]));
Q_ASSIGN U3456 ( .B(clk), .A(\g.we_clk [29318]));
Q_ASSIGN U3457 ( .B(clk), .A(\g.we_clk [29317]));
Q_ASSIGN U3458 ( .B(clk), .A(\g.we_clk [29316]));
Q_ASSIGN U3459 ( .B(clk), .A(\g.we_clk [29315]));
Q_ASSIGN U3460 ( .B(clk), .A(\g.we_clk [29314]));
Q_ASSIGN U3461 ( .B(clk), .A(\g.we_clk [29313]));
Q_ASSIGN U3462 ( .B(clk), .A(\g.we_clk [29312]));
Q_ASSIGN U3463 ( .B(clk), .A(\g.we_clk [29311]));
Q_ASSIGN U3464 ( .B(clk), .A(\g.we_clk [29310]));
Q_ASSIGN U3465 ( .B(clk), .A(\g.we_clk [29309]));
Q_ASSIGN U3466 ( .B(clk), .A(\g.we_clk [29308]));
Q_ASSIGN U3467 ( .B(clk), .A(\g.we_clk [29307]));
Q_ASSIGN U3468 ( .B(clk), .A(\g.we_clk [29306]));
Q_ASSIGN U3469 ( .B(clk), .A(\g.we_clk [29305]));
Q_ASSIGN U3470 ( .B(clk), .A(\g.we_clk [29304]));
Q_ASSIGN U3471 ( .B(clk), .A(\g.we_clk [29303]));
Q_ASSIGN U3472 ( .B(clk), .A(\g.we_clk [29302]));
Q_ASSIGN U3473 ( .B(clk), .A(\g.we_clk [29301]));
Q_ASSIGN U3474 ( .B(clk), .A(\g.we_clk [29300]));
Q_ASSIGN U3475 ( .B(clk), .A(\g.we_clk [29299]));
Q_ASSIGN U3476 ( .B(clk), .A(\g.we_clk [29298]));
Q_ASSIGN U3477 ( .B(clk), .A(\g.we_clk [29297]));
Q_ASSIGN U3478 ( .B(clk), .A(\g.we_clk [29296]));
Q_ASSIGN U3479 ( .B(clk), .A(\g.we_clk [29295]));
Q_ASSIGN U3480 ( .B(clk), .A(\g.we_clk [29294]));
Q_ASSIGN U3481 ( .B(clk), .A(\g.we_clk [29293]));
Q_ASSIGN U3482 ( .B(clk), .A(\g.we_clk [29292]));
Q_ASSIGN U3483 ( .B(clk), .A(\g.we_clk [29291]));
Q_ASSIGN U3484 ( .B(clk), .A(\g.we_clk [29290]));
Q_ASSIGN U3485 ( .B(clk), .A(\g.we_clk [29289]));
Q_ASSIGN U3486 ( .B(clk), .A(\g.we_clk [29288]));
Q_ASSIGN U3487 ( .B(clk), .A(\g.we_clk [29287]));
Q_ASSIGN U3488 ( .B(clk), .A(\g.we_clk [29286]));
Q_ASSIGN U3489 ( .B(clk), .A(\g.we_clk [29285]));
Q_ASSIGN U3490 ( .B(clk), .A(\g.we_clk [29284]));
Q_ASSIGN U3491 ( .B(clk), .A(\g.we_clk [29283]));
Q_ASSIGN U3492 ( .B(clk), .A(\g.we_clk [29282]));
Q_ASSIGN U3493 ( .B(clk), .A(\g.we_clk [29281]));
Q_ASSIGN U3494 ( .B(clk), .A(\g.we_clk [29280]));
Q_ASSIGN U3495 ( .B(clk), .A(\g.we_clk [29279]));
Q_ASSIGN U3496 ( .B(clk), .A(\g.we_clk [29278]));
Q_ASSIGN U3497 ( .B(clk), .A(\g.we_clk [29277]));
Q_ASSIGN U3498 ( .B(clk), .A(\g.we_clk [29276]));
Q_ASSIGN U3499 ( .B(clk), .A(\g.we_clk [29275]));
Q_ASSIGN U3500 ( .B(clk), .A(\g.we_clk [29274]));
Q_ASSIGN U3501 ( .B(clk), .A(\g.we_clk [29273]));
Q_ASSIGN U3502 ( .B(clk), .A(\g.we_clk [29272]));
Q_ASSIGN U3503 ( .B(clk), .A(\g.we_clk [29271]));
Q_ASSIGN U3504 ( .B(clk), .A(\g.we_clk [29270]));
Q_ASSIGN U3505 ( .B(clk), .A(\g.we_clk [29269]));
Q_ASSIGN U3506 ( .B(clk), .A(\g.we_clk [29268]));
Q_ASSIGN U3507 ( .B(clk), .A(\g.we_clk [29267]));
Q_ASSIGN U3508 ( .B(clk), .A(\g.we_clk [29266]));
Q_ASSIGN U3509 ( .B(clk), .A(\g.we_clk [29265]));
Q_ASSIGN U3510 ( .B(clk), .A(\g.we_clk [29264]));
Q_ASSIGN U3511 ( .B(clk), .A(\g.we_clk [29263]));
Q_ASSIGN U3512 ( .B(clk), .A(\g.we_clk [29262]));
Q_ASSIGN U3513 ( .B(clk), .A(\g.we_clk [29261]));
Q_ASSIGN U3514 ( .B(clk), .A(\g.we_clk [29260]));
Q_ASSIGN U3515 ( .B(clk), .A(\g.we_clk [29259]));
Q_ASSIGN U3516 ( .B(clk), .A(\g.we_clk [29258]));
Q_ASSIGN U3517 ( .B(clk), .A(\g.we_clk [29257]));
Q_ASSIGN U3518 ( .B(clk), .A(\g.we_clk [29256]));
Q_ASSIGN U3519 ( .B(clk), .A(\g.we_clk [29255]));
Q_ASSIGN U3520 ( .B(clk), .A(\g.we_clk [29254]));
Q_ASSIGN U3521 ( .B(clk), .A(\g.we_clk [29253]));
Q_ASSIGN U3522 ( .B(clk), .A(\g.we_clk [29252]));
Q_ASSIGN U3523 ( .B(clk), .A(\g.we_clk [29251]));
Q_ASSIGN U3524 ( .B(clk), .A(\g.we_clk [29250]));
Q_ASSIGN U3525 ( .B(clk), .A(\g.we_clk [29249]));
Q_ASSIGN U3526 ( .B(clk), .A(\g.we_clk [29248]));
Q_ASSIGN U3527 ( .B(clk), .A(\g.we_clk [29247]));
Q_ASSIGN U3528 ( .B(clk), .A(\g.we_clk [29246]));
Q_ASSIGN U3529 ( .B(clk), .A(\g.we_clk [29245]));
Q_ASSIGN U3530 ( .B(clk), .A(\g.we_clk [29244]));
Q_ASSIGN U3531 ( .B(clk), .A(\g.we_clk [29243]));
Q_ASSIGN U3532 ( .B(clk), .A(\g.we_clk [29242]));
Q_ASSIGN U3533 ( .B(clk), .A(\g.we_clk [29241]));
Q_ASSIGN U3534 ( .B(clk), .A(\g.we_clk [29240]));
Q_ASSIGN U3535 ( .B(clk), .A(\g.we_clk [29239]));
Q_ASSIGN U3536 ( .B(clk), .A(\g.we_clk [29238]));
Q_ASSIGN U3537 ( .B(clk), .A(\g.we_clk [29237]));
Q_ASSIGN U3538 ( .B(clk), .A(\g.we_clk [29236]));
Q_ASSIGN U3539 ( .B(clk), .A(\g.we_clk [29235]));
Q_ASSIGN U3540 ( .B(clk), .A(\g.we_clk [29234]));
Q_ASSIGN U3541 ( .B(clk), .A(\g.we_clk [29233]));
Q_ASSIGN U3542 ( .B(clk), .A(\g.we_clk [29232]));
Q_ASSIGN U3543 ( .B(clk), .A(\g.we_clk [29231]));
Q_ASSIGN U3544 ( .B(clk), .A(\g.we_clk [29230]));
Q_ASSIGN U3545 ( .B(clk), .A(\g.we_clk [29229]));
Q_ASSIGN U3546 ( .B(clk), .A(\g.we_clk [29228]));
Q_ASSIGN U3547 ( .B(clk), .A(\g.we_clk [29227]));
Q_ASSIGN U3548 ( .B(clk), .A(\g.we_clk [29226]));
Q_ASSIGN U3549 ( .B(clk), .A(\g.we_clk [29225]));
Q_ASSIGN U3550 ( .B(clk), .A(\g.we_clk [29224]));
Q_ASSIGN U3551 ( .B(clk), .A(\g.we_clk [29223]));
Q_ASSIGN U3552 ( .B(clk), .A(\g.we_clk [29222]));
Q_ASSIGN U3553 ( .B(clk), .A(\g.we_clk [29221]));
Q_ASSIGN U3554 ( .B(clk), .A(\g.we_clk [29220]));
Q_ASSIGN U3555 ( .B(clk), .A(\g.we_clk [29219]));
Q_ASSIGN U3556 ( .B(clk), .A(\g.we_clk [29218]));
Q_ASSIGN U3557 ( .B(clk), .A(\g.we_clk [29217]));
Q_ASSIGN U3558 ( .B(clk), .A(\g.we_clk [29216]));
Q_ASSIGN U3559 ( .B(clk), .A(\g.we_clk [29215]));
Q_ASSIGN U3560 ( .B(clk), .A(\g.we_clk [29214]));
Q_ASSIGN U3561 ( .B(clk), .A(\g.we_clk [29213]));
Q_ASSIGN U3562 ( .B(clk), .A(\g.we_clk [29212]));
Q_ASSIGN U3563 ( .B(clk), .A(\g.we_clk [29211]));
Q_ASSIGN U3564 ( .B(clk), .A(\g.we_clk [29210]));
Q_ASSIGN U3565 ( .B(clk), .A(\g.we_clk [29209]));
Q_ASSIGN U3566 ( .B(clk), .A(\g.we_clk [29208]));
Q_ASSIGN U3567 ( .B(clk), .A(\g.we_clk [29207]));
Q_ASSIGN U3568 ( .B(clk), .A(\g.we_clk [29206]));
Q_ASSIGN U3569 ( .B(clk), .A(\g.we_clk [29205]));
Q_ASSIGN U3570 ( .B(clk), .A(\g.we_clk [29204]));
Q_ASSIGN U3571 ( .B(clk), .A(\g.we_clk [29203]));
Q_ASSIGN U3572 ( .B(clk), .A(\g.we_clk [29202]));
Q_ASSIGN U3573 ( .B(clk), .A(\g.we_clk [29201]));
Q_ASSIGN U3574 ( .B(clk), .A(\g.we_clk [29200]));
Q_ASSIGN U3575 ( .B(clk), .A(\g.we_clk [29199]));
Q_ASSIGN U3576 ( .B(clk), .A(\g.we_clk [29198]));
Q_ASSIGN U3577 ( .B(clk), .A(\g.we_clk [29197]));
Q_ASSIGN U3578 ( .B(clk), .A(\g.we_clk [29196]));
Q_ASSIGN U3579 ( .B(clk), .A(\g.we_clk [29195]));
Q_ASSIGN U3580 ( .B(clk), .A(\g.we_clk [29194]));
Q_ASSIGN U3581 ( .B(clk), .A(\g.we_clk [29193]));
Q_ASSIGN U3582 ( .B(clk), .A(\g.we_clk [29192]));
Q_ASSIGN U3583 ( .B(clk), .A(\g.we_clk [29191]));
Q_ASSIGN U3584 ( .B(clk), .A(\g.we_clk [29190]));
Q_ASSIGN U3585 ( .B(clk), .A(\g.we_clk [29189]));
Q_ASSIGN U3586 ( .B(clk), .A(\g.we_clk [29188]));
Q_ASSIGN U3587 ( .B(clk), .A(\g.we_clk [29187]));
Q_ASSIGN U3588 ( .B(clk), .A(\g.we_clk [29186]));
Q_ASSIGN U3589 ( .B(clk), .A(\g.we_clk [29185]));
Q_ASSIGN U3590 ( .B(clk), .A(\g.we_clk [29184]));
Q_ASSIGN U3591 ( .B(clk), .A(\g.we_clk [29183]));
Q_ASSIGN U3592 ( .B(clk), .A(\g.we_clk [29182]));
Q_ASSIGN U3593 ( .B(clk), .A(\g.we_clk [29181]));
Q_ASSIGN U3594 ( .B(clk), .A(\g.we_clk [29180]));
Q_ASSIGN U3595 ( .B(clk), .A(\g.we_clk [29179]));
Q_ASSIGN U3596 ( .B(clk), .A(\g.we_clk [29178]));
Q_ASSIGN U3597 ( .B(clk), .A(\g.we_clk [29177]));
Q_ASSIGN U3598 ( .B(clk), .A(\g.we_clk [29176]));
Q_ASSIGN U3599 ( .B(clk), .A(\g.we_clk [29175]));
Q_ASSIGN U3600 ( .B(clk), .A(\g.we_clk [29174]));
Q_ASSIGN U3601 ( .B(clk), .A(\g.we_clk [29173]));
Q_ASSIGN U3602 ( .B(clk), .A(\g.we_clk [29172]));
Q_ASSIGN U3603 ( .B(clk), .A(\g.we_clk [29171]));
Q_ASSIGN U3604 ( .B(clk), .A(\g.we_clk [29170]));
Q_ASSIGN U3605 ( .B(clk), .A(\g.we_clk [29169]));
Q_ASSIGN U3606 ( .B(clk), .A(\g.we_clk [29168]));
Q_ASSIGN U3607 ( .B(clk), .A(\g.we_clk [29167]));
Q_ASSIGN U3608 ( .B(clk), .A(\g.we_clk [29166]));
Q_ASSIGN U3609 ( .B(clk), .A(\g.we_clk [29165]));
Q_ASSIGN U3610 ( .B(clk), .A(\g.we_clk [29164]));
Q_ASSIGN U3611 ( .B(clk), .A(\g.we_clk [29163]));
Q_ASSIGN U3612 ( .B(clk), .A(\g.we_clk [29162]));
Q_ASSIGN U3613 ( .B(clk), .A(\g.we_clk [29161]));
Q_ASSIGN U3614 ( .B(clk), .A(\g.we_clk [29160]));
Q_ASSIGN U3615 ( .B(clk), .A(\g.we_clk [29159]));
Q_ASSIGN U3616 ( .B(clk), .A(\g.we_clk [29158]));
Q_ASSIGN U3617 ( .B(clk), .A(\g.we_clk [29157]));
Q_ASSIGN U3618 ( .B(clk), .A(\g.we_clk [29156]));
Q_ASSIGN U3619 ( .B(clk), .A(\g.we_clk [29155]));
Q_ASSIGN U3620 ( .B(clk), .A(\g.we_clk [29154]));
Q_ASSIGN U3621 ( .B(clk), .A(\g.we_clk [29153]));
Q_ASSIGN U3622 ( .B(clk), .A(\g.we_clk [29152]));
Q_ASSIGN U3623 ( .B(clk), .A(\g.we_clk [29151]));
Q_ASSIGN U3624 ( .B(clk), .A(\g.we_clk [29150]));
Q_ASSIGN U3625 ( .B(clk), .A(\g.we_clk [29149]));
Q_ASSIGN U3626 ( .B(clk), .A(\g.we_clk [29148]));
Q_ASSIGN U3627 ( .B(clk), .A(\g.we_clk [29147]));
Q_ASSIGN U3628 ( .B(clk), .A(\g.we_clk [29146]));
Q_ASSIGN U3629 ( .B(clk), .A(\g.we_clk [29145]));
Q_ASSIGN U3630 ( .B(clk), .A(\g.we_clk [29144]));
Q_ASSIGN U3631 ( .B(clk), .A(\g.we_clk [29143]));
Q_ASSIGN U3632 ( .B(clk), .A(\g.we_clk [29142]));
Q_ASSIGN U3633 ( .B(clk), .A(\g.we_clk [29141]));
Q_ASSIGN U3634 ( .B(clk), .A(\g.we_clk [29140]));
Q_ASSIGN U3635 ( .B(clk), .A(\g.we_clk [29139]));
Q_ASSIGN U3636 ( .B(clk), .A(\g.we_clk [29138]));
Q_ASSIGN U3637 ( .B(clk), .A(\g.we_clk [29137]));
Q_ASSIGN U3638 ( .B(clk), .A(\g.we_clk [29136]));
Q_ASSIGN U3639 ( .B(clk), .A(\g.we_clk [29135]));
Q_ASSIGN U3640 ( .B(clk), .A(\g.we_clk [29134]));
Q_ASSIGN U3641 ( .B(clk), .A(\g.we_clk [29133]));
Q_ASSIGN U3642 ( .B(clk), .A(\g.we_clk [29132]));
Q_ASSIGN U3643 ( .B(clk), .A(\g.we_clk [29131]));
Q_ASSIGN U3644 ( .B(clk), .A(\g.we_clk [29130]));
Q_ASSIGN U3645 ( .B(clk), .A(\g.we_clk [29129]));
Q_ASSIGN U3646 ( .B(clk), .A(\g.we_clk [29128]));
Q_ASSIGN U3647 ( .B(clk), .A(\g.we_clk [29127]));
Q_ASSIGN U3648 ( .B(clk), .A(\g.we_clk [29126]));
Q_ASSIGN U3649 ( .B(clk), .A(\g.we_clk [29125]));
Q_ASSIGN U3650 ( .B(clk), .A(\g.we_clk [29124]));
Q_ASSIGN U3651 ( .B(clk), .A(\g.we_clk [29123]));
Q_ASSIGN U3652 ( .B(clk), .A(\g.we_clk [29122]));
Q_ASSIGN U3653 ( .B(clk), .A(\g.we_clk [29121]));
Q_ASSIGN U3654 ( .B(clk), .A(\g.we_clk [29120]));
Q_ASSIGN U3655 ( .B(clk), .A(\g.we_clk [29119]));
Q_ASSIGN U3656 ( .B(clk), .A(\g.we_clk [29118]));
Q_ASSIGN U3657 ( .B(clk), .A(\g.we_clk [29117]));
Q_ASSIGN U3658 ( .B(clk), .A(\g.we_clk [29116]));
Q_ASSIGN U3659 ( .B(clk), .A(\g.we_clk [29115]));
Q_ASSIGN U3660 ( .B(clk), .A(\g.we_clk [29114]));
Q_ASSIGN U3661 ( .B(clk), .A(\g.we_clk [29113]));
Q_ASSIGN U3662 ( .B(clk), .A(\g.we_clk [29112]));
Q_ASSIGN U3663 ( .B(clk), .A(\g.we_clk [29111]));
Q_ASSIGN U3664 ( .B(clk), .A(\g.we_clk [29110]));
Q_ASSIGN U3665 ( .B(clk), .A(\g.we_clk [29109]));
Q_ASSIGN U3666 ( .B(clk), .A(\g.we_clk [29108]));
Q_ASSIGN U3667 ( .B(clk), .A(\g.we_clk [29107]));
Q_ASSIGN U3668 ( .B(clk), .A(\g.we_clk [29106]));
Q_ASSIGN U3669 ( .B(clk), .A(\g.we_clk [29105]));
Q_ASSIGN U3670 ( .B(clk), .A(\g.we_clk [29104]));
Q_ASSIGN U3671 ( .B(clk), .A(\g.we_clk [29103]));
Q_ASSIGN U3672 ( .B(clk), .A(\g.we_clk [29102]));
Q_ASSIGN U3673 ( .B(clk), .A(\g.we_clk [29101]));
Q_ASSIGN U3674 ( .B(clk), .A(\g.we_clk [29100]));
Q_ASSIGN U3675 ( .B(clk), .A(\g.we_clk [29099]));
Q_ASSIGN U3676 ( .B(clk), .A(\g.we_clk [29098]));
Q_ASSIGN U3677 ( .B(clk), .A(\g.we_clk [29097]));
Q_ASSIGN U3678 ( .B(clk), .A(\g.we_clk [29096]));
Q_ASSIGN U3679 ( .B(clk), .A(\g.we_clk [29095]));
Q_ASSIGN U3680 ( .B(clk), .A(\g.we_clk [29094]));
Q_ASSIGN U3681 ( .B(clk), .A(\g.we_clk [29093]));
Q_ASSIGN U3682 ( .B(clk), .A(\g.we_clk [29092]));
Q_ASSIGN U3683 ( .B(clk), .A(\g.we_clk [29091]));
Q_ASSIGN U3684 ( .B(clk), .A(\g.we_clk [29090]));
Q_ASSIGN U3685 ( .B(clk), .A(\g.we_clk [29089]));
Q_ASSIGN U3686 ( .B(clk), .A(\g.we_clk [29088]));
Q_ASSIGN U3687 ( .B(clk), .A(\g.we_clk [29087]));
Q_ASSIGN U3688 ( .B(clk), .A(\g.we_clk [29086]));
Q_ASSIGN U3689 ( .B(clk), .A(\g.we_clk [29085]));
Q_ASSIGN U3690 ( .B(clk), .A(\g.we_clk [29084]));
Q_ASSIGN U3691 ( .B(clk), .A(\g.we_clk [29083]));
Q_ASSIGN U3692 ( .B(clk), .A(\g.we_clk [29082]));
Q_ASSIGN U3693 ( .B(clk), .A(\g.we_clk [29081]));
Q_ASSIGN U3694 ( .B(clk), .A(\g.we_clk [29080]));
Q_ASSIGN U3695 ( .B(clk), .A(\g.we_clk [29079]));
Q_ASSIGN U3696 ( .B(clk), .A(\g.we_clk [29078]));
Q_ASSIGN U3697 ( .B(clk), .A(\g.we_clk [29077]));
Q_ASSIGN U3698 ( .B(clk), .A(\g.we_clk [29076]));
Q_ASSIGN U3699 ( .B(clk), .A(\g.we_clk [29075]));
Q_ASSIGN U3700 ( .B(clk), .A(\g.we_clk [29074]));
Q_ASSIGN U3701 ( .B(clk), .A(\g.we_clk [29073]));
Q_ASSIGN U3702 ( .B(clk), .A(\g.we_clk [29072]));
Q_ASSIGN U3703 ( .B(clk), .A(\g.we_clk [29071]));
Q_ASSIGN U3704 ( .B(clk), .A(\g.we_clk [29070]));
Q_ASSIGN U3705 ( .B(clk), .A(\g.we_clk [29069]));
Q_ASSIGN U3706 ( .B(clk), .A(\g.we_clk [29068]));
Q_ASSIGN U3707 ( .B(clk), .A(\g.we_clk [29067]));
Q_ASSIGN U3708 ( .B(clk), .A(\g.we_clk [29066]));
Q_ASSIGN U3709 ( .B(clk), .A(\g.we_clk [29065]));
Q_ASSIGN U3710 ( .B(clk), .A(\g.we_clk [29064]));
Q_ASSIGN U3711 ( .B(clk), .A(\g.we_clk [29063]));
Q_ASSIGN U3712 ( .B(clk), .A(\g.we_clk [29062]));
Q_ASSIGN U3713 ( .B(clk), .A(\g.we_clk [29061]));
Q_ASSIGN U3714 ( .B(clk), .A(\g.we_clk [29060]));
Q_ASSIGN U3715 ( .B(clk), .A(\g.we_clk [29059]));
Q_ASSIGN U3716 ( .B(clk), .A(\g.we_clk [29058]));
Q_ASSIGN U3717 ( .B(clk), .A(\g.we_clk [29057]));
Q_ASSIGN U3718 ( .B(clk), .A(\g.we_clk [29056]));
Q_ASSIGN U3719 ( .B(clk), .A(\g.we_clk [29055]));
Q_ASSIGN U3720 ( .B(clk), .A(\g.we_clk [29054]));
Q_ASSIGN U3721 ( .B(clk), .A(\g.we_clk [29053]));
Q_ASSIGN U3722 ( .B(clk), .A(\g.we_clk [29052]));
Q_ASSIGN U3723 ( .B(clk), .A(\g.we_clk [29051]));
Q_ASSIGN U3724 ( .B(clk), .A(\g.we_clk [29050]));
Q_ASSIGN U3725 ( .B(clk), .A(\g.we_clk [29049]));
Q_ASSIGN U3726 ( .B(clk), .A(\g.we_clk [29048]));
Q_ASSIGN U3727 ( .B(clk), .A(\g.we_clk [29047]));
Q_ASSIGN U3728 ( .B(clk), .A(\g.we_clk [29046]));
Q_ASSIGN U3729 ( .B(clk), .A(\g.we_clk [29045]));
Q_ASSIGN U3730 ( .B(clk), .A(\g.we_clk [29044]));
Q_ASSIGN U3731 ( .B(clk), .A(\g.we_clk [29043]));
Q_ASSIGN U3732 ( .B(clk), .A(\g.we_clk [29042]));
Q_ASSIGN U3733 ( .B(clk), .A(\g.we_clk [29041]));
Q_ASSIGN U3734 ( .B(clk), .A(\g.we_clk [29040]));
Q_ASSIGN U3735 ( .B(clk), .A(\g.we_clk [29039]));
Q_ASSIGN U3736 ( .B(clk), .A(\g.we_clk [29038]));
Q_ASSIGN U3737 ( .B(clk), .A(\g.we_clk [29037]));
Q_ASSIGN U3738 ( .B(clk), .A(\g.we_clk [29036]));
Q_ASSIGN U3739 ( .B(clk), .A(\g.we_clk [29035]));
Q_ASSIGN U3740 ( .B(clk), .A(\g.we_clk [29034]));
Q_ASSIGN U3741 ( .B(clk), .A(\g.we_clk [29033]));
Q_ASSIGN U3742 ( .B(clk), .A(\g.we_clk [29032]));
Q_ASSIGN U3743 ( .B(clk), .A(\g.we_clk [29031]));
Q_ASSIGN U3744 ( .B(clk), .A(\g.we_clk [29030]));
Q_ASSIGN U3745 ( .B(clk), .A(\g.we_clk [29029]));
Q_ASSIGN U3746 ( .B(clk), .A(\g.we_clk [29028]));
Q_ASSIGN U3747 ( .B(clk), .A(\g.we_clk [29027]));
Q_ASSIGN U3748 ( .B(clk), .A(\g.we_clk [29026]));
Q_ASSIGN U3749 ( .B(clk), .A(\g.we_clk [29025]));
Q_ASSIGN U3750 ( .B(clk), .A(\g.we_clk [29024]));
Q_ASSIGN U3751 ( .B(clk), .A(\g.we_clk [29023]));
Q_ASSIGN U3752 ( .B(clk), .A(\g.we_clk [29022]));
Q_ASSIGN U3753 ( .B(clk), .A(\g.we_clk [29021]));
Q_ASSIGN U3754 ( .B(clk), .A(\g.we_clk [29020]));
Q_ASSIGN U3755 ( .B(clk), .A(\g.we_clk [29019]));
Q_ASSIGN U3756 ( .B(clk), .A(\g.we_clk [29018]));
Q_ASSIGN U3757 ( .B(clk), .A(\g.we_clk [29017]));
Q_ASSIGN U3758 ( .B(clk), .A(\g.we_clk [29016]));
Q_ASSIGN U3759 ( .B(clk), .A(\g.we_clk [29015]));
Q_ASSIGN U3760 ( .B(clk), .A(\g.we_clk [29014]));
Q_ASSIGN U3761 ( .B(clk), .A(\g.we_clk [29013]));
Q_ASSIGN U3762 ( .B(clk), .A(\g.we_clk [29012]));
Q_ASSIGN U3763 ( .B(clk), .A(\g.we_clk [29011]));
Q_ASSIGN U3764 ( .B(clk), .A(\g.we_clk [29010]));
Q_ASSIGN U3765 ( .B(clk), .A(\g.we_clk [29009]));
Q_ASSIGN U3766 ( .B(clk), .A(\g.we_clk [29008]));
Q_ASSIGN U3767 ( .B(clk), .A(\g.we_clk [29007]));
Q_ASSIGN U3768 ( .B(clk), .A(\g.we_clk [29006]));
Q_ASSIGN U3769 ( .B(clk), .A(\g.we_clk [29005]));
Q_ASSIGN U3770 ( .B(clk), .A(\g.we_clk [29004]));
Q_ASSIGN U3771 ( .B(clk), .A(\g.we_clk [29003]));
Q_ASSIGN U3772 ( .B(clk), .A(\g.we_clk [29002]));
Q_ASSIGN U3773 ( .B(clk), .A(\g.we_clk [29001]));
Q_ASSIGN U3774 ( .B(clk), .A(\g.we_clk [29000]));
Q_ASSIGN U3775 ( .B(clk), .A(\g.we_clk [28999]));
Q_ASSIGN U3776 ( .B(clk), .A(\g.we_clk [28998]));
Q_ASSIGN U3777 ( .B(clk), .A(\g.we_clk [28997]));
Q_ASSIGN U3778 ( .B(clk), .A(\g.we_clk [28996]));
Q_ASSIGN U3779 ( .B(clk), .A(\g.we_clk [28995]));
Q_ASSIGN U3780 ( .B(clk), .A(\g.we_clk [28994]));
Q_ASSIGN U3781 ( .B(clk), .A(\g.we_clk [28993]));
Q_ASSIGN U3782 ( .B(clk), .A(\g.we_clk [28992]));
Q_ASSIGN U3783 ( .B(clk), .A(\g.we_clk [28991]));
Q_ASSIGN U3784 ( .B(clk), .A(\g.we_clk [28990]));
Q_ASSIGN U3785 ( .B(clk), .A(\g.we_clk [28989]));
Q_ASSIGN U3786 ( .B(clk), .A(\g.we_clk [28988]));
Q_ASSIGN U3787 ( .B(clk), .A(\g.we_clk [28987]));
Q_ASSIGN U3788 ( .B(clk), .A(\g.we_clk [28986]));
Q_ASSIGN U3789 ( .B(clk), .A(\g.we_clk [28985]));
Q_ASSIGN U3790 ( .B(clk), .A(\g.we_clk [28984]));
Q_ASSIGN U3791 ( .B(clk), .A(\g.we_clk [28983]));
Q_ASSIGN U3792 ( .B(clk), .A(\g.we_clk [28982]));
Q_ASSIGN U3793 ( .B(clk), .A(\g.we_clk [28981]));
Q_ASSIGN U3794 ( .B(clk), .A(\g.we_clk [28980]));
Q_ASSIGN U3795 ( .B(clk), .A(\g.we_clk [28979]));
Q_ASSIGN U3796 ( .B(clk), .A(\g.we_clk [28978]));
Q_ASSIGN U3797 ( .B(clk), .A(\g.we_clk [28977]));
Q_ASSIGN U3798 ( .B(clk), .A(\g.we_clk [28976]));
Q_ASSIGN U3799 ( .B(clk), .A(\g.we_clk [28975]));
Q_ASSIGN U3800 ( .B(clk), .A(\g.we_clk [28974]));
Q_ASSIGN U3801 ( .B(clk), .A(\g.we_clk [28973]));
Q_ASSIGN U3802 ( .B(clk), .A(\g.we_clk [28972]));
Q_ASSIGN U3803 ( .B(clk), .A(\g.we_clk [28971]));
Q_ASSIGN U3804 ( .B(clk), .A(\g.we_clk [28970]));
Q_ASSIGN U3805 ( .B(clk), .A(\g.we_clk [28969]));
Q_ASSIGN U3806 ( .B(clk), .A(\g.we_clk [28968]));
Q_ASSIGN U3807 ( .B(clk), .A(\g.we_clk [28967]));
Q_ASSIGN U3808 ( .B(clk), .A(\g.we_clk [28966]));
Q_ASSIGN U3809 ( .B(clk), .A(\g.we_clk [28965]));
Q_ASSIGN U3810 ( .B(clk), .A(\g.we_clk [28964]));
Q_ASSIGN U3811 ( .B(clk), .A(\g.we_clk [28963]));
Q_ASSIGN U3812 ( .B(clk), .A(\g.we_clk [28962]));
Q_ASSIGN U3813 ( .B(clk), .A(\g.we_clk [28961]));
Q_ASSIGN U3814 ( .B(clk), .A(\g.we_clk [28960]));
Q_ASSIGN U3815 ( .B(clk), .A(\g.we_clk [28959]));
Q_ASSIGN U3816 ( .B(clk), .A(\g.we_clk [28958]));
Q_ASSIGN U3817 ( .B(clk), .A(\g.we_clk [28957]));
Q_ASSIGN U3818 ( .B(clk), .A(\g.we_clk [28956]));
Q_ASSIGN U3819 ( .B(clk), .A(\g.we_clk [28955]));
Q_ASSIGN U3820 ( .B(clk), .A(\g.we_clk [28954]));
Q_ASSIGN U3821 ( .B(clk), .A(\g.we_clk [28953]));
Q_ASSIGN U3822 ( .B(clk), .A(\g.we_clk [28952]));
Q_ASSIGN U3823 ( .B(clk), .A(\g.we_clk [28951]));
Q_ASSIGN U3824 ( .B(clk), .A(\g.we_clk [28950]));
Q_ASSIGN U3825 ( .B(clk), .A(\g.we_clk [28949]));
Q_ASSIGN U3826 ( .B(clk), .A(\g.we_clk [28948]));
Q_ASSIGN U3827 ( .B(clk), .A(\g.we_clk [28947]));
Q_ASSIGN U3828 ( .B(clk), .A(\g.we_clk [28946]));
Q_ASSIGN U3829 ( .B(clk), .A(\g.we_clk [28945]));
Q_ASSIGN U3830 ( .B(clk), .A(\g.we_clk [28944]));
Q_ASSIGN U3831 ( .B(clk), .A(\g.we_clk [28943]));
Q_ASSIGN U3832 ( .B(clk), .A(\g.we_clk [28942]));
Q_ASSIGN U3833 ( .B(clk), .A(\g.we_clk [28941]));
Q_ASSIGN U3834 ( .B(clk), .A(\g.we_clk [28940]));
Q_ASSIGN U3835 ( .B(clk), .A(\g.we_clk [28939]));
Q_ASSIGN U3836 ( .B(clk), .A(\g.we_clk [28938]));
Q_ASSIGN U3837 ( .B(clk), .A(\g.we_clk [28937]));
Q_ASSIGN U3838 ( .B(clk), .A(\g.we_clk [28936]));
Q_ASSIGN U3839 ( .B(clk), .A(\g.we_clk [28935]));
Q_ASSIGN U3840 ( .B(clk), .A(\g.we_clk [28934]));
Q_ASSIGN U3841 ( .B(clk), .A(\g.we_clk [28933]));
Q_ASSIGN U3842 ( .B(clk), .A(\g.we_clk [28932]));
Q_ASSIGN U3843 ( .B(clk), .A(\g.we_clk [28931]));
Q_ASSIGN U3844 ( .B(clk), .A(\g.we_clk [28930]));
Q_ASSIGN U3845 ( .B(clk), .A(\g.we_clk [28929]));
Q_ASSIGN U3846 ( .B(clk), .A(\g.we_clk [28928]));
Q_ASSIGN U3847 ( .B(clk), .A(\g.we_clk [28927]));
Q_ASSIGN U3848 ( .B(clk), .A(\g.we_clk [28926]));
Q_ASSIGN U3849 ( .B(clk), .A(\g.we_clk [28925]));
Q_ASSIGN U3850 ( .B(clk), .A(\g.we_clk [28924]));
Q_ASSIGN U3851 ( .B(clk), .A(\g.we_clk [28923]));
Q_ASSIGN U3852 ( .B(clk), .A(\g.we_clk [28922]));
Q_ASSIGN U3853 ( .B(clk), .A(\g.we_clk [28921]));
Q_ASSIGN U3854 ( .B(clk), .A(\g.we_clk [28920]));
Q_ASSIGN U3855 ( .B(clk), .A(\g.we_clk [28919]));
Q_ASSIGN U3856 ( .B(clk), .A(\g.we_clk [28918]));
Q_ASSIGN U3857 ( .B(clk), .A(\g.we_clk [28917]));
Q_ASSIGN U3858 ( .B(clk), .A(\g.we_clk [28916]));
Q_ASSIGN U3859 ( .B(clk), .A(\g.we_clk [28915]));
Q_ASSIGN U3860 ( .B(clk), .A(\g.we_clk [28914]));
Q_ASSIGN U3861 ( .B(clk), .A(\g.we_clk [28913]));
Q_ASSIGN U3862 ( .B(clk), .A(\g.we_clk [28912]));
Q_ASSIGN U3863 ( .B(clk), .A(\g.we_clk [28911]));
Q_ASSIGN U3864 ( .B(clk), .A(\g.we_clk [28910]));
Q_ASSIGN U3865 ( .B(clk), .A(\g.we_clk [28909]));
Q_ASSIGN U3866 ( .B(clk), .A(\g.we_clk [28908]));
Q_ASSIGN U3867 ( .B(clk), .A(\g.we_clk [28907]));
Q_ASSIGN U3868 ( .B(clk), .A(\g.we_clk [28906]));
Q_ASSIGN U3869 ( .B(clk), .A(\g.we_clk [28905]));
Q_ASSIGN U3870 ( .B(clk), .A(\g.we_clk [28904]));
Q_ASSIGN U3871 ( .B(clk), .A(\g.we_clk [28903]));
Q_ASSIGN U3872 ( .B(clk), .A(\g.we_clk [28902]));
Q_ASSIGN U3873 ( .B(clk), .A(\g.we_clk [28901]));
Q_ASSIGN U3874 ( .B(clk), .A(\g.we_clk [28900]));
Q_ASSIGN U3875 ( .B(clk), .A(\g.we_clk [28899]));
Q_ASSIGN U3876 ( .B(clk), .A(\g.we_clk [28898]));
Q_ASSIGN U3877 ( .B(clk), .A(\g.we_clk [28897]));
Q_ASSIGN U3878 ( .B(clk), .A(\g.we_clk [28896]));
Q_ASSIGN U3879 ( .B(clk), .A(\g.we_clk [28895]));
Q_ASSIGN U3880 ( .B(clk), .A(\g.we_clk [28894]));
Q_ASSIGN U3881 ( .B(clk), .A(\g.we_clk [28893]));
Q_ASSIGN U3882 ( .B(clk), .A(\g.we_clk [28892]));
Q_ASSIGN U3883 ( .B(clk), .A(\g.we_clk [28891]));
Q_ASSIGN U3884 ( .B(clk), .A(\g.we_clk [28890]));
Q_ASSIGN U3885 ( .B(clk), .A(\g.we_clk [28889]));
Q_ASSIGN U3886 ( .B(clk), .A(\g.we_clk [28888]));
Q_ASSIGN U3887 ( .B(clk), .A(\g.we_clk [28887]));
Q_ASSIGN U3888 ( .B(clk), .A(\g.we_clk [28886]));
Q_ASSIGN U3889 ( .B(clk), .A(\g.we_clk [28885]));
Q_ASSIGN U3890 ( .B(clk), .A(\g.we_clk [28884]));
Q_ASSIGN U3891 ( .B(clk), .A(\g.we_clk [28883]));
Q_ASSIGN U3892 ( .B(clk), .A(\g.we_clk [28882]));
Q_ASSIGN U3893 ( .B(clk), .A(\g.we_clk [28881]));
Q_ASSIGN U3894 ( .B(clk), .A(\g.we_clk [28880]));
Q_ASSIGN U3895 ( .B(clk), .A(\g.we_clk [28879]));
Q_ASSIGN U3896 ( .B(clk), .A(\g.we_clk [28878]));
Q_ASSIGN U3897 ( .B(clk), .A(\g.we_clk [28877]));
Q_ASSIGN U3898 ( .B(clk), .A(\g.we_clk [28876]));
Q_ASSIGN U3899 ( .B(clk), .A(\g.we_clk [28875]));
Q_ASSIGN U3900 ( .B(clk), .A(\g.we_clk [28874]));
Q_ASSIGN U3901 ( .B(clk), .A(\g.we_clk [28873]));
Q_ASSIGN U3902 ( .B(clk), .A(\g.we_clk [28872]));
Q_ASSIGN U3903 ( .B(clk), .A(\g.we_clk [28871]));
Q_ASSIGN U3904 ( .B(clk), .A(\g.we_clk [28870]));
Q_ASSIGN U3905 ( .B(clk), .A(\g.we_clk [28869]));
Q_ASSIGN U3906 ( .B(clk), .A(\g.we_clk [28868]));
Q_ASSIGN U3907 ( .B(clk), .A(\g.we_clk [28867]));
Q_ASSIGN U3908 ( .B(clk), .A(\g.we_clk [28866]));
Q_ASSIGN U3909 ( .B(clk), .A(\g.we_clk [28865]));
Q_ASSIGN U3910 ( .B(clk), .A(\g.we_clk [28864]));
Q_ASSIGN U3911 ( .B(clk), .A(\g.we_clk [28863]));
Q_ASSIGN U3912 ( .B(clk), .A(\g.we_clk [28862]));
Q_ASSIGN U3913 ( .B(clk), .A(\g.we_clk [28861]));
Q_ASSIGN U3914 ( .B(clk), .A(\g.we_clk [28860]));
Q_ASSIGN U3915 ( .B(clk), .A(\g.we_clk [28859]));
Q_ASSIGN U3916 ( .B(clk), .A(\g.we_clk [28858]));
Q_ASSIGN U3917 ( .B(clk), .A(\g.we_clk [28857]));
Q_ASSIGN U3918 ( .B(clk), .A(\g.we_clk [28856]));
Q_ASSIGN U3919 ( .B(clk), .A(\g.we_clk [28855]));
Q_ASSIGN U3920 ( .B(clk), .A(\g.we_clk [28854]));
Q_ASSIGN U3921 ( .B(clk), .A(\g.we_clk [28853]));
Q_ASSIGN U3922 ( .B(clk), .A(\g.we_clk [28852]));
Q_ASSIGN U3923 ( .B(clk), .A(\g.we_clk [28851]));
Q_ASSIGN U3924 ( .B(clk), .A(\g.we_clk [28850]));
Q_ASSIGN U3925 ( .B(clk), .A(\g.we_clk [28849]));
Q_ASSIGN U3926 ( .B(clk), .A(\g.we_clk [28848]));
Q_ASSIGN U3927 ( .B(clk), .A(\g.we_clk [28847]));
Q_ASSIGN U3928 ( .B(clk), .A(\g.we_clk [28846]));
Q_ASSIGN U3929 ( .B(clk), .A(\g.we_clk [28845]));
Q_ASSIGN U3930 ( .B(clk), .A(\g.we_clk [28844]));
Q_ASSIGN U3931 ( .B(clk), .A(\g.we_clk [28843]));
Q_ASSIGN U3932 ( .B(clk), .A(\g.we_clk [28842]));
Q_ASSIGN U3933 ( .B(clk), .A(\g.we_clk [28841]));
Q_ASSIGN U3934 ( .B(clk), .A(\g.we_clk [28840]));
Q_ASSIGN U3935 ( .B(clk), .A(\g.we_clk [28839]));
Q_ASSIGN U3936 ( .B(clk), .A(\g.we_clk [28838]));
Q_ASSIGN U3937 ( .B(clk), .A(\g.we_clk [28837]));
Q_ASSIGN U3938 ( .B(clk), .A(\g.we_clk [28836]));
Q_ASSIGN U3939 ( .B(clk), .A(\g.we_clk [28835]));
Q_ASSIGN U3940 ( .B(clk), .A(\g.we_clk [28834]));
Q_ASSIGN U3941 ( .B(clk), .A(\g.we_clk [28833]));
Q_ASSIGN U3942 ( .B(clk), .A(\g.we_clk [28832]));
Q_ASSIGN U3943 ( .B(clk), .A(\g.we_clk [28831]));
Q_ASSIGN U3944 ( .B(clk), .A(\g.we_clk [28830]));
Q_ASSIGN U3945 ( .B(clk), .A(\g.we_clk [28829]));
Q_ASSIGN U3946 ( .B(clk), .A(\g.we_clk [28828]));
Q_ASSIGN U3947 ( .B(clk), .A(\g.we_clk [28827]));
Q_ASSIGN U3948 ( .B(clk), .A(\g.we_clk [28826]));
Q_ASSIGN U3949 ( .B(clk), .A(\g.we_clk [28825]));
Q_ASSIGN U3950 ( .B(clk), .A(\g.we_clk [28824]));
Q_ASSIGN U3951 ( .B(clk), .A(\g.we_clk [28823]));
Q_ASSIGN U3952 ( .B(clk), .A(\g.we_clk [28822]));
Q_ASSIGN U3953 ( .B(clk), .A(\g.we_clk [28821]));
Q_ASSIGN U3954 ( .B(clk), .A(\g.we_clk [28820]));
Q_ASSIGN U3955 ( .B(clk), .A(\g.we_clk [28819]));
Q_ASSIGN U3956 ( .B(clk), .A(\g.we_clk [28818]));
Q_ASSIGN U3957 ( .B(clk), .A(\g.we_clk [28817]));
Q_ASSIGN U3958 ( .B(clk), .A(\g.we_clk [28816]));
Q_ASSIGN U3959 ( .B(clk), .A(\g.we_clk [28815]));
Q_ASSIGN U3960 ( .B(clk), .A(\g.we_clk [28814]));
Q_ASSIGN U3961 ( .B(clk), .A(\g.we_clk [28813]));
Q_ASSIGN U3962 ( .B(clk), .A(\g.we_clk [28812]));
Q_ASSIGN U3963 ( .B(clk), .A(\g.we_clk [28811]));
Q_ASSIGN U3964 ( .B(clk), .A(\g.we_clk [28810]));
Q_ASSIGN U3965 ( .B(clk), .A(\g.we_clk [28809]));
Q_ASSIGN U3966 ( .B(clk), .A(\g.we_clk [28808]));
Q_ASSIGN U3967 ( .B(clk), .A(\g.we_clk [28807]));
Q_ASSIGN U3968 ( .B(clk), .A(\g.we_clk [28806]));
Q_ASSIGN U3969 ( .B(clk), .A(\g.we_clk [28805]));
Q_ASSIGN U3970 ( .B(clk), .A(\g.we_clk [28804]));
Q_ASSIGN U3971 ( .B(clk), .A(\g.we_clk [28803]));
Q_ASSIGN U3972 ( .B(clk), .A(\g.we_clk [28802]));
Q_ASSIGN U3973 ( .B(clk), .A(\g.we_clk [28801]));
Q_ASSIGN U3974 ( .B(clk), .A(\g.we_clk [28800]));
Q_ASSIGN U3975 ( .B(clk), .A(\g.we_clk [28799]));
Q_ASSIGN U3976 ( .B(clk), .A(\g.we_clk [28798]));
Q_ASSIGN U3977 ( .B(clk), .A(\g.we_clk [28797]));
Q_ASSIGN U3978 ( .B(clk), .A(\g.we_clk [28796]));
Q_ASSIGN U3979 ( .B(clk), .A(\g.we_clk [28795]));
Q_ASSIGN U3980 ( .B(clk), .A(\g.we_clk [28794]));
Q_ASSIGN U3981 ( .B(clk), .A(\g.we_clk [28793]));
Q_ASSIGN U3982 ( .B(clk), .A(\g.we_clk [28792]));
Q_ASSIGN U3983 ( .B(clk), .A(\g.we_clk [28791]));
Q_ASSIGN U3984 ( .B(clk), .A(\g.we_clk [28790]));
Q_ASSIGN U3985 ( .B(clk), .A(\g.we_clk [28789]));
Q_ASSIGN U3986 ( .B(clk), .A(\g.we_clk [28788]));
Q_ASSIGN U3987 ( .B(clk), .A(\g.we_clk [28787]));
Q_ASSIGN U3988 ( .B(clk), .A(\g.we_clk [28786]));
Q_ASSIGN U3989 ( .B(clk), .A(\g.we_clk [28785]));
Q_ASSIGN U3990 ( .B(clk), .A(\g.we_clk [28784]));
Q_ASSIGN U3991 ( .B(clk), .A(\g.we_clk [28783]));
Q_ASSIGN U3992 ( .B(clk), .A(\g.we_clk [28782]));
Q_ASSIGN U3993 ( .B(clk), .A(\g.we_clk [28781]));
Q_ASSIGN U3994 ( .B(clk), .A(\g.we_clk [28780]));
Q_ASSIGN U3995 ( .B(clk), .A(\g.we_clk [28779]));
Q_ASSIGN U3996 ( .B(clk), .A(\g.we_clk [28778]));
Q_ASSIGN U3997 ( .B(clk), .A(\g.we_clk [28777]));
Q_ASSIGN U3998 ( .B(clk), .A(\g.we_clk [28776]));
Q_ASSIGN U3999 ( .B(clk), .A(\g.we_clk [28775]));
Q_ASSIGN U4000 ( .B(clk), .A(\g.we_clk [28774]));
Q_ASSIGN U4001 ( .B(clk), .A(\g.we_clk [28773]));
Q_ASSIGN U4002 ( .B(clk), .A(\g.we_clk [28772]));
Q_ASSIGN U4003 ( .B(clk), .A(\g.we_clk [28771]));
Q_ASSIGN U4004 ( .B(clk), .A(\g.we_clk [28770]));
Q_ASSIGN U4005 ( .B(clk), .A(\g.we_clk [28769]));
Q_ASSIGN U4006 ( .B(clk), .A(\g.we_clk [28768]));
Q_ASSIGN U4007 ( .B(clk), .A(\g.we_clk [28767]));
Q_ASSIGN U4008 ( .B(clk), .A(\g.we_clk [28766]));
Q_ASSIGN U4009 ( .B(clk), .A(\g.we_clk [28765]));
Q_ASSIGN U4010 ( .B(clk), .A(\g.we_clk [28764]));
Q_ASSIGN U4011 ( .B(clk), .A(\g.we_clk [28763]));
Q_ASSIGN U4012 ( .B(clk), .A(\g.we_clk [28762]));
Q_ASSIGN U4013 ( .B(clk), .A(\g.we_clk [28761]));
Q_ASSIGN U4014 ( .B(clk), .A(\g.we_clk [28760]));
Q_ASSIGN U4015 ( .B(clk), .A(\g.we_clk [28759]));
Q_ASSIGN U4016 ( .B(clk), .A(\g.we_clk [28758]));
Q_ASSIGN U4017 ( .B(clk), .A(\g.we_clk [28757]));
Q_ASSIGN U4018 ( .B(clk), .A(\g.we_clk [28756]));
Q_ASSIGN U4019 ( .B(clk), .A(\g.we_clk [28755]));
Q_ASSIGN U4020 ( .B(clk), .A(\g.we_clk [28754]));
Q_ASSIGN U4021 ( .B(clk), .A(\g.we_clk [28753]));
Q_ASSIGN U4022 ( .B(clk), .A(\g.we_clk [28752]));
Q_ASSIGN U4023 ( .B(clk), .A(\g.we_clk [28751]));
Q_ASSIGN U4024 ( .B(clk), .A(\g.we_clk [28750]));
Q_ASSIGN U4025 ( .B(clk), .A(\g.we_clk [28749]));
Q_ASSIGN U4026 ( .B(clk), .A(\g.we_clk [28748]));
Q_ASSIGN U4027 ( .B(clk), .A(\g.we_clk [28747]));
Q_ASSIGN U4028 ( .B(clk), .A(\g.we_clk [28746]));
Q_ASSIGN U4029 ( .B(clk), .A(\g.we_clk [28745]));
Q_ASSIGN U4030 ( .B(clk), .A(\g.we_clk [28744]));
Q_ASSIGN U4031 ( .B(clk), .A(\g.we_clk [28743]));
Q_ASSIGN U4032 ( .B(clk), .A(\g.we_clk [28742]));
Q_ASSIGN U4033 ( .B(clk), .A(\g.we_clk [28741]));
Q_ASSIGN U4034 ( .B(clk), .A(\g.we_clk [28740]));
Q_ASSIGN U4035 ( .B(clk), .A(\g.we_clk [28739]));
Q_ASSIGN U4036 ( .B(clk), .A(\g.we_clk [28738]));
Q_ASSIGN U4037 ( .B(clk), .A(\g.we_clk [28737]));
Q_ASSIGN U4038 ( .B(clk), .A(\g.we_clk [28736]));
Q_ASSIGN U4039 ( .B(clk), .A(\g.we_clk [28735]));
Q_ASSIGN U4040 ( .B(clk), .A(\g.we_clk [28734]));
Q_ASSIGN U4041 ( .B(clk), .A(\g.we_clk [28733]));
Q_ASSIGN U4042 ( .B(clk), .A(\g.we_clk [28732]));
Q_ASSIGN U4043 ( .B(clk), .A(\g.we_clk [28731]));
Q_ASSIGN U4044 ( .B(clk), .A(\g.we_clk [28730]));
Q_ASSIGN U4045 ( .B(clk), .A(\g.we_clk [28729]));
Q_ASSIGN U4046 ( .B(clk), .A(\g.we_clk [28728]));
Q_ASSIGN U4047 ( .B(clk), .A(\g.we_clk [28727]));
Q_ASSIGN U4048 ( .B(clk), .A(\g.we_clk [28726]));
Q_ASSIGN U4049 ( .B(clk), .A(\g.we_clk [28725]));
Q_ASSIGN U4050 ( .B(clk), .A(\g.we_clk [28724]));
Q_ASSIGN U4051 ( .B(clk), .A(\g.we_clk [28723]));
Q_ASSIGN U4052 ( .B(clk), .A(\g.we_clk [28722]));
Q_ASSIGN U4053 ( .B(clk), .A(\g.we_clk [28721]));
Q_ASSIGN U4054 ( .B(clk), .A(\g.we_clk [28720]));
Q_ASSIGN U4055 ( .B(clk), .A(\g.we_clk [28719]));
Q_ASSIGN U4056 ( .B(clk), .A(\g.we_clk [28718]));
Q_ASSIGN U4057 ( .B(clk), .A(\g.we_clk [28717]));
Q_ASSIGN U4058 ( .B(clk), .A(\g.we_clk [28716]));
Q_ASSIGN U4059 ( .B(clk), .A(\g.we_clk [28715]));
Q_ASSIGN U4060 ( .B(clk), .A(\g.we_clk [28714]));
Q_ASSIGN U4061 ( .B(clk), .A(\g.we_clk [28713]));
Q_ASSIGN U4062 ( .B(clk), .A(\g.we_clk [28712]));
Q_ASSIGN U4063 ( .B(clk), .A(\g.we_clk [28711]));
Q_ASSIGN U4064 ( .B(clk), .A(\g.we_clk [28710]));
Q_ASSIGN U4065 ( .B(clk), .A(\g.we_clk [28709]));
Q_ASSIGN U4066 ( .B(clk), .A(\g.we_clk [28708]));
Q_ASSIGN U4067 ( .B(clk), .A(\g.we_clk [28707]));
Q_ASSIGN U4068 ( .B(clk), .A(\g.we_clk [28706]));
Q_ASSIGN U4069 ( .B(clk), .A(\g.we_clk [28705]));
Q_ASSIGN U4070 ( .B(clk), .A(\g.we_clk [28704]));
Q_ASSIGN U4071 ( .B(clk), .A(\g.we_clk [28703]));
Q_ASSIGN U4072 ( .B(clk), .A(\g.we_clk [28702]));
Q_ASSIGN U4073 ( .B(clk), .A(\g.we_clk [28701]));
Q_ASSIGN U4074 ( .B(clk), .A(\g.we_clk [28700]));
Q_ASSIGN U4075 ( .B(clk), .A(\g.we_clk [28699]));
Q_ASSIGN U4076 ( .B(clk), .A(\g.we_clk [28698]));
Q_ASSIGN U4077 ( .B(clk), .A(\g.we_clk [28697]));
Q_ASSIGN U4078 ( .B(clk), .A(\g.we_clk [28696]));
Q_ASSIGN U4079 ( .B(clk), .A(\g.we_clk [28695]));
Q_ASSIGN U4080 ( .B(clk), .A(\g.we_clk [28694]));
Q_ASSIGN U4081 ( .B(clk), .A(\g.we_clk [28693]));
Q_ASSIGN U4082 ( .B(clk), .A(\g.we_clk [28692]));
Q_ASSIGN U4083 ( .B(clk), .A(\g.we_clk [28691]));
Q_ASSIGN U4084 ( .B(clk), .A(\g.we_clk [28690]));
Q_ASSIGN U4085 ( .B(clk), .A(\g.we_clk [28689]));
Q_ASSIGN U4086 ( .B(clk), .A(\g.we_clk [28688]));
Q_ASSIGN U4087 ( .B(clk), .A(\g.we_clk [28687]));
Q_ASSIGN U4088 ( .B(clk), .A(\g.we_clk [28686]));
Q_ASSIGN U4089 ( .B(clk), .A(\g.we_clk [28685]));
Q_ASSIGN U4090 ( .B(clk), .A(\g.we_clk [28684]));
Q_ASSIGN U4091 ( .B(clk), .A(\g.we_clk [28683]));
Q_ASSIGN U4092 ( .B(clk), .A(\g.we_clk [28682]));
Q_ASSIGN U4093 ( .B(clk), .A(\g.we_clk [28681]));
Q_ASSIGN U4094 ( .B(clk), .A(\g.we_clk [28680]));
Q_ASSIGN U4095 ( .B(clk), .A(\g.we_clk [28679]));
Q_ASSIGN U4096 ( .B(clk), .A(\g.we_clk [28678]));
Q_ASSIGN U4097 ( .B(clk), .A(\g.we_clk [28677]));
Q_ASSIGN U4098 ( .B(clk), .A(\g.we_clk [28676]));
Q_ASSIGN U4099 ( .B(clk), .A(\g.we_clk [28675]));
Q_ASSIGN U4100 ( .B(clk), .A(\g.we_clk [28674]));
Q_ASSIGN U4101 ( .B(clk), .A(\g.we_clk [28673]));
Q_ASSIGN U4102 ( .B(clk), .A(\g.we_clk [28672]));
Q_ASSIGN U4103 ( .B(clk), .A(\g.we_clk [28671]));
Q_ASSIGN U4104 ( .B(clk), .A(\g.we_clk [28670]));
Q_ASSIGN U4105 ( .B(clk), .A(\g.we_clk [28669]));
Q_ASSIGN U4106 ( .B(clk), .A(\g.we_clk [28668]));
Q_ASSIGN U4107 ( .B(clk), .A(\g.we_clk [28667]));
Q_ASSIGN U4108 ( .B(clk), .A(\g.we_clk [28666]));
Q_ASSIGN U4109 ( .B(clk), .A(\g.we_clk [28665]));
Q_ASSIGN U4110 ( .B(clk), .A(\g.we_clk [28664]));
Q_ASSIGN U4111 ( .B(clk), .A(\g.we_clk [28663]));
Q_ASSIGN U4112 ( .B(clk), .A(\g.we_clk [28662]));
Q_ASSIGN U4113 ( .B(clk), .A(\g.we_clk [28661]));
Q_ASSIGN U4114 ( .B(clk), .A(\g.we_clk [28660]));
Q_ASSIGN U4115 ( .B(clk), .A(\g.we_clk [28659]));
Q_ASSIGN U4116 ( .B(clk), .A(\g.we_clk [28658]));
Q_ASSIGN U4117 ( .B(clk), .A(\g.we_clk [28657]));
Q_ASSIGN U4118 ( .B(clk), .A(\g.we_clk [28656]));
Q_ASSIGN U4119 ( .B(clk), .A(\g.we_clk [28655]));
Q_ASSIGN U4120 ( .B(clk), .A(\g.we_clk [28654]));
Q_ASSIGN U4121 ( .B(clk), .A(\g.we_clk [28653]));
Q_ASSIGN U4122 ( .B(clk), .A(\g.we_clk [28652]));
Q_ASSIGN U4123 ( .B(clk), .A(\g.we_clk [28651]));
Q_ASSIGN U4124 ( .B(clk), .A(\g.we_clk [28650]));
Q_ASSIGN U4125 ( .B(clk), .A(\g.we_clk [28649]));
Q_ASSIGN U4126 ( .B(clk), .A(\g.we_clk [28648]));
Q_ASSIGN U4127 ( .B(clk), .A(\g.we_clk [28647]));
Q_ASSIGN U4128 ( .B(clk), .A(\g.we_clk [28646]));
Q_ASSIGN U4129 ( .B(clk), .A(\g.we_clk [28645]));
Q_ASSIGN U4130 ( .B(clk), .A(\g.we_clk [28644]));
Q_ASSIGN U4131 ( .B(clk), .A(\g.we_clk [28643]));
Q_ASSIGN U4132 ( .B(clk), .A(\g.we_clk [28642]));
Q_ASSIGN U4133 ( .B(clk), .A(\g.we_clk [28641]));
Q_ASSIGN U4134 ( .B(clk), .A(\g.we_clk [28640]));
Q_ASSIGN U4135 ( .B(clk), .A(\g.we_clk [28639]));
Q_ASSIGN U4136 ( .B(clk), .A(\g.we_clk [28638]));
Q_ASSIGN U4137 ( .B(clk), .A(\g.we_clk [28637]));
Q_ASSIGN U4138 ( .B(clk), .A(\g.we_clk [28636]));
Q_ASSIGN U4139 ( .B(clk), .A(\g.we_clk [28635]));
Q_ASSIGN U4140 ( .B(clk), .A(\g.we_clk [28634]));
Q_ASSIGN U4141 ( .B(clk), .A(\g.we_clk [28633]));
Q_ASSIGN U4142 ( .B(clk), .A(\g.we_clk [28632]));
Q_ASSIGN U4143 ( .B(clk), .A(\g.we_clk [28631]));
Q_ASSIGN U4144 ( .B(clk), .A(\g.we_clk [28630]));
Q_ASSIGN U4145 ( .B(clk), .A(\g.we_clk [28629]));
Q_ASSIGN U4146 ( .B(clk), .A(\g.we_clk [28628]));
Q_ASSIGN U4147 ( .B(clk), .A(\g.we_clk [28627]));
Q_ASSIGN U4148 ( .B(clk), .A(\g.we_clk [28626]));
Q_ASSIGN U4149 ( .B(clk), .A(\g.we_clk [28625]));
Q_ASSIGN U4150 ( .B(clk), .A(\g.we_clk [28624]));
Q_ASSIGN U4151 ( .B(clk), .A(\g.we_clk [28623]));
Q_ASSIGN U4152 ( .B(clk), .A(\g.we_clk [28622]));
Q_ASSIGN U4153 ( .B(clk), .A(\g.we_clk [28621]));
Q_ASSIGN U4154 ( .B(clk), .A(\g.we_clk [28620]));
Q_ASSIGN U4155 ( .B(clk), .A(\g.we_clk [28619]));
Q_ASSIGN U4156 ( .B(clk), .A(\g.we_clk [28618]));
Q_ASSIGN U4157 ( .B(clk), .A(\g.we_clk [28617]));
Q_ASSIGN U4158 ( .B(clk), .A(\g.we_clk [28616]));
Q_ASSIGN U4159 ( .B(clk), .A(\g.we_clk [28615]));
Q_ASSIGN U4160 ( .B(clk), .A(\g.we_clk [28614]));
Q_ASSIGN U4161 ( .B(clk), .A(\g.we_clk [28613]));
Q_ASSIGN U4162 ( .B(clk), .A(\g.we_clk [28612]));
Q_ASSIGN U4163 ( .B(clk), .A(\g.we_clk [28611]));
Q_ASSIGN U4164 ( .B(clk), .A(\g.we_clk [28610]));
Q_ASSIGN U4165 ( .B(clk), .A(\g.we_clk [28609]));
Q_ASSIGN U4166 ( .B(clk), .A(\g.we_clk [28608]));
Q_ASSIGN U4167 ( .B(clk), .A(\g.we_clk [28607]));
Q_ASSIGN U4168 ( .B(clk), .A(\g.we_clk [28606]));
Q_ASSIGN U4169 ( .B(clk), .A(\g.we_clk [28605]));
Q_ASSIGN U4170 ( .B(clk), .A(\g.we_clk [28604]));
Q_ASSIGN U4171 ( .B(clk), .A(\g.we_clk [28603]));
Q_ASSIGN U4172 ( .B(clk), .A(\g.we_clk [28602]));
Q_ASSIGN U4173 ( .B(clk), .A(\g.we_clk [28601]));
Q_ASSIGN U4174 ( .B(clk), .A(\g.we_clk [28600]));
Q_ASSIGN U4175 ( .B(clk), .A(\g.we_clk [28599]));
Q_ASSIGN U4176 ( .B(clk), .A(\g.we_clk [28598]));
Q_ASSIGN U4177 ( .B(clk), .A(\g.we_clk [28597]));
Q_ASSIGN U4178 ( .B(clk), .A(\g.we_clk [28596]));
Q_ASSIGN U4179 ( .B(clk), .A(\g.we_clk [28595]));
Q_ASSIGN U4180 ( .B(clk), .A(\g.we_clk [28594]));
Q_ASSIGN U4181 ( .B(clk), .A(\g.we_clk [28593]));
Q_ASSIGN U4182 ( .B(clk), .A(\g.we_clk [28592]));
Q_ASSIGN U4183 ( .B(clk), .A(\g.we_clk [28591]));
Q_ASSIGN U4184 ( .B(clk), .A(\g.we_clk [28590]));
Q_ASSIGN U4185 ( .B(clk), .A(\g.we_clk [28589]));
Q_ASSIGN U4186 ( .B(clk), .A(\g.we_clk [28588]));
Q_ASSIGN U4187 ( .B(clk), .A(\g.we_clk [28587]));
Q_ASSIGN U4188 ( .B(clk), .A(\g.we_clk [28586]));
Q_ASSIGN U4189 ( .B(clk), .A(\g.we_clk [28585]));
Q_ASSIGN U4190 ( .B(clk), .A(\g.we_clk [28584]));
Q_ASSIGN U4191 ( .B(clk), .A(\g.we_clk [28583]));
Q_ASSIGN U4192 ( .B(clk), .A(\g.we_clk [28582]));
Q_ASSIGN U4193 ( .B(clk), .A(\g.we_clk [28581]));
Q_ASSIGN U4194 ( .B(clk), .A(\g.we_clk [28580]));
Q_ASSIGN U4195 ( .B(clk), .A(\g.we_clk [28579]));
Q_ASSIGN U4196 ( .B(clk), .A(\g.we_clk [28578]));
Q_ASSIGN U4197 ( .B(clk), .A(\g.we_clk [28577]));
Q_ASSIGN U4198 ( .B(clk), .A(\g.we_clk [28576]));
Q_ASSIGN U4199 ( .B(clk), .A(\g.we_clk [28575]));
Q_ASSIGN U4200 ( .B(clk), .A(\g.we_clk [28574]));
Q_ASSIGN U4201 ( .B(clk), .A(\g.we_clk [28573]));
Q_ASSIGN U4202 ( .B(clk), .A(\g.we_clk [28572]));
Q_ASSIGN U4203 ( .B(clk), .A(\g.we_clk [28571]));
Q_ASSIGN U4204 ( .B(clk), .A(\g.we_clk [28570]));
Q_ASSIGN U4205 ( .B(clk), .A(\g.we_clk [28569]));
Q_ASSIGN U4206 ( .B(clk), .A(\g.we_clk [28568]));
Q_ASSIGN U4207 ( .B(clk), .A(\g.we_clk [28567]));
Q_ASSIGN U4208 ( .B(clk), .A(\g.we_clk [28566]));
Q_ASSIGN U4209 ( .B(clk), .A(\g.we_clk [28565]));
Q_ASSIGN U4210 ( .B(clk), .A(\g.we_clk [28564]));
Q_ASSIGN U4211 ( .B(clk), .A(\g.we_clk [28563]));
Q_ASSIGN U4212 ( .B(clk), .A(\g.we_clk [28562]));
Q_ASSIGN U4213 ( .B(clk), .A(\g.we_clk [28561]));
Q_ASSIGN U4214 ( .B(clk), .A(\g.we_clk [28560]));
Q_ASSIGN U4215 ( .B(clk), .A(\g.we_clk [28559]));
Q_ASSIGN U4216 ( .B(clk), .A(\g.we_clk [28558]));
Q_ASSIGN U4217 ( .B(clk), .A(\g.we_clk [28557]));
Q_ASSIGN U4218 ( .B(clk), .A(\g.we_clk [28556]));
Q_ASSIGN U4219 ( .B(clk), .A(\g.we_clk [28555]));
Q_ASSIGN U4220 ( .B(clk), .A(\g.we_clk [28554]));
Q_ASSIGN U4221 ( .B(clk), .A(\g.we_clk [28553]));
Q_ASSIGN U4222 ( .B(clk), .A(\g.we_clk [28552]));
Q_ASSIGN U4223 ( .B(clk), .A(\g.we_clk [28551]));
Q_ASSIGN U4224 ( .B(clk), .A(\g.we_clk [28550]));
Q_ASSIGN U4225 ( .B(clk), .A(\g.we_clk [28549]));
Q_ASSIGN U4226 ( .B(clk), .A(\g.we_clk [28548]));
Q_ASSIGN U4227 ( .B(clk), .A(\g.we_clk [28547]));
Q_ASSIGN U4228 ( .B(clk), .A(\g.we_clk [28546]));
Q_ASSIGN U4229 ( .B(clk), .A(\g.we_clk [28545]));
Q_ASSIGN U4230 ( .B(clk), .A(\g.we_clk [28544]));
Q_ASSIGN U4231 ( .B(clk), .A(\g.we_clk [28543]));
Q_ASSIGN U4232 ( .B(clk), .A(\g.we_clk [28542]));
Q_ASSIGN U4233 ( .B(clk), .A(\g.we_clk [28541]));
Q_ASSIGN U4234 ( .B(clk), .A(\g.we_clk [28540]));
Q_ASSIGN U4235 ( .B(clk), .A(\g.we_clk [28539]));
Q_ASSIGN U4236 ( .B(clk), .A(\g.we_clk [28538]));
Q_ASSIGN U4237 ( .B(clk), .A(\g.we_clk [28537]));
Q_ASSIGN U4238 ( .B(clk), .A(\g.we_clk [28536]));
Q_ASSIGN U4239 ( .B(clk), .A(\g.we_clk [28535]));
Q_ASSIGN U4240 ( .B(clk), .A(\g.we_clk [28534]));
Q_ASSIGN U4241 ( .B(clk), .A(\g.we_clk [28533]));
Q_ASSIGN U4242 ( .B(clk), .A(\g.we_clk [28532]));
Q_ASSIGN U4243 ( .B(clk), .A(\g.we_clk [28531]));
Q_ASSIGN U4244 ( .B(clk), .A(\g.we_clk [28530]));
Q_ASSIGN U4245 ( .B(clk), .A(\g.we_clk [28529]));
Q_ASSIGN U4246 ( .B(clk), .A(\g.we_clk [28528]));
Q_ASSIGN U4247 ( .B(clk), .A(\g.we_clk [28527]));
Q_ASSIGN U4248 ( .B(clk), .A(\g.we_clk [28526]));
Q_ASSIGN U4249 ( .B(clk), .A(\g.we_clk [28525]));
Q_ASSIGN U4250 ( .B(clk), .A(\g.we_clk [28524]));
Q_ASSIGN U4251 ( .B(clk), .A(\g.we_clk [28523]));
Q_ASSIGN U4252 ( .B(clk), .A(\g.we_clk [28522]));
Q_ASSIGN U4253 ( .B(clk), .A(\g.we_clk [28521]));
Q_ASSIGN U4254 ( .B(clk), .A(\g.we_clk [28520]));
Q_ASSIGN U4255 ( .B(clk), .A(\g.we_clk [28519]));
Q_ASSIGN U4256 ( .B(clk), .A(\g.we_clk [28518]));
Q_ASSIGN U4257 ( .B(clk), .A(\g.we_clk [28517]));
Q_ASSIGN U4258 ( .B(clk), .A(\g.we_clk [28516]));
Q_ASSIGN U4259 ( .B(clk), .A(\g.we_clk [28515]));
Q_ASSIGN U4260 ( .B(clk), .A(\g.we_clk [28514]));
Q_ASSIGN U4261 ( .B(clk), .A(\g.we_clk [28513]));
Q_ASSIGN U4262 ( .B(clk), .A(\g.we_clk [28512]));
Q_ASSIGN U4263 ( .B(clk), .A(\g.we_clk [28511]));
Q_ASSIGN U4264 ( .B(clk), .A(\g.we_clk [28510]));
Q_ASSIGN U4265 ( .B(clk), .A(\g.we_clk [28509]));
Q_ASSIGN U4266 ( .B(clk), .A(\g.we_clk [28508]));
Q_ASSIGN U4267 ( .B(clk), .A(\g.we_clk [28507]));
Q_ASSIGN U4268 ( .B(clk), .A(\g.we_clk [28506]));
Q_ASSIGN U4269 ( .B(clk), .A(\g.we_clk [28505]));
Q_ASSIGN U4270 ( .B(clk), .A(\g.we_clk [28504]));
Q_ASSIGN U4271 ( .B(clk), .A(\g.we_clk [28503]));
Q_ASSIGN U4272 ( .B(clk), .A(\g.we_clk [28502]));
Q_ASSIGN U4273 ( .B(clk), .A(\g.we_clk [28501]));
Q_ASSIGN U4274 ( .B(clk), .A(\g.we_clk [28500]));
Q_ASSIGN U4275 ( .B(clk), .A(\g.we_clk [28499]));
Q_ASSIGN U4276 ( .B(clk), .A(\g.we_clk [28498]));
Q_ASSIGN U4277 ( .B(clk), .A(\g.we_clk [28497]));
Q_ASSIGN U4278 ( .B(clk), .A(\g.we_clk [28496]));
Q_ASSIGN U4279 ( .B(clk), .A(\g.we_clk [28495]));
Q_ASSIGN U4280 ( .B(clk), .A(\g.we_clk [28494]));
Q_ASSIGN U4281 ( .B(clk), .A(\g.we_clk [28493]));
Q_ASSIGN U4282 ( .B(clk), .A(\g.we_clk [28492]));
Q_ASSIGN U4283 ( .B(clk), .A(\g.we_clk [28491]));
Q_ASSIGN U4284 ( .B(clk), .A(\g.we_clk [28490]));
Q_ASSIGN U4285 ( .B(clk), .A(\g.we_clk [28489]));
Q_ASSIGN U4286 ( .B(clk), .A(\g.we_clk [28488]));
Q_ASSIGN U4287 ( .B(clk), .A(\g.we_clk [28487]));
Q_ASSIGN U4288 ( .B(clk), .A(\g.we_clk [28486]));
Q_ASSIGN U4289 ( .B(clk), .A(\g.we_clk [28485]));
Q_ASSIGN U4290 ( .B(clk), .A(\g.we_clk [28484]));
Q_ASSIGN U4291 ( .B(clk), .A(\g.we_clk [28483]));
Q_ASSIGN U4292 ( .B(clk), .A(\g.we_clk [28482]));
Q_ASSIGN U4293 ( .B(clk), .A(\g.we_clk [28481]));
Q_ASSIGN U4294 ( .B(clk), .A(\g.we_clk [28480]));
Q_ASSIGN U4295 ( .B(clk), .A(\g.we_clk [28479]));
Q_ASSIGN U4296 ( .B(clk), .A(\g.we_clk [28478]));
Q_ASSIGN U4297 ( .B(clk), .A(\g.we_clk [28477]));
Q_ASSIGN U4298 ( .B(clk), .A(\g.we_clk [28476]));
Q_ASSIGN U4299 ( .B(clk), .A(\g.we_clk [28475]));
Q_ASSIGN U4300 ( .B(clk), .A(\g.we_clk [28474]));
Q_ASSIGN U4301 ( .B(clk), .A(\g.we_clk [28473]));
Q_ASSIGN U4302 ( .B(clk), .A(\g.we_clk [28472]));
Q_ASSIGN U4303 ( .B(clk), .A(\g.we_clk [28471]));
Q_ASSIGN U4304 ( .B(clk), .A(\g.we_clk [28470]));
Q_ASSIGN U4305 ( .B(clk), .A(\g.we_clk [28469]));
Q_ASSIGN U4306 ( .B(clk), .A(\g.we_clk [28468]));
Q_ASSIGN U4307 ( .B(clk), .A(\g.we_clk [28467]));
Q_ASSIGN U4308 ( .B(clk), .A(\g.we_clk [28466]));
Q_ASSIGN U4309 ( .B(clk), .A(\g.we_clk [28465]));
Q_ASSIGN U4310 ( .B(clk), .A(\g.we_clk [28464]));
Q_ASSIGN U4311 ( .B(clk), .A(\g.we_clk [28463]));
Q_ASSIGN U4312 ( .B(clk), .A(\g.we_clk [28462]));
Q_ASSIGN U4313 ( .B(clk), .A(\g.we_clk [28461]));
Q_ASSIGN U4314 ( .B(clk), .A(\g.we_clk [28460]));
Q_ASSIGN U4315 ( .B(clk), .A(\g.we_clk [28459]));
Q_ASSIGN U4316 ( .B(clk), .A(\g.we_clk [28458]));
Q_ASSIGN U4317 ( .B(clk), .A(\g.we_clk [28457]));
Q_ASSIGN U4318 ( .B(clk), .A(\g.we_clk [28456]));
Q_ASSIGN U4319 ( .B(clk), .A(\g.we_clk [28455]));
Q_ASSIGN U4320 ( .B(clk), .A(\g.we_clk [28454]));
Q_ASSIGN U4321 ( .B(clk), .A(\g.we_clk [28453]));
Q_ASSIGN U4322 ( .B(clk), .A(\g.we_clk [28452]));
Q_ASSIGN U4323 ( .B(clk), .A(\g.we_clk [28451]));
Q_ASSIGN U4324 ( .B(clk), .A(\g.we_clk [28450]));
Q_ASSIGN U4325 ( .B(clk), .A(\g.we_clk [28449]));
Q_ASSIGN U4326 ( .B(clk), .A(\g.we_clk [28448]));
Q_ASSIGN U4327 ( .B(clk), .A(\g.we_clk [28447]));
Q_ASSIGN U4328 ( .B(clk), .A(\g.we_clk [28446]));
Q_ASSIGN U4329 ( .B(clk), .A(\g.we_clk [28445]));
Q_ASSIGN U4330 ( .B(clk), .A(\g.we_clk [28444]));
Q_ASSIGN U4331 ( .B(clk), .A(\g.we_clk [28443]));
Q_ASSIGN U4332 ( .B(clk), .A(\g.we_clk [28442]));
Q_ASSIGN U4333 ( .B(clk), .A(\g.we_clk [28441]));
Q_ASSIGN U4334 ( .B(clk), .A(\g.we_clk [28440]));
Q_ASSIGN U4335 ( .B(clk), .A(\g.we_clk [28439]));
Q_ASSIGN U4336 ( .B(clk), .A(\g.we_clk [28438]));
Q_ASSIGN U4337 ( .B(clk), .A(\g.we_clk [28437]));
Q_ASSIGN U4338 ( .B(clk), .A(\g.we_clk [28436]));
Q_ASSIGN U4339 ( .B(clk), .A(\g.we_clk [28435]));
Q_ASSIGN U4340 ( .B(clk), .A(\g.we_clk [28434]));
Q_ASSIGN U4341 ( .B(clk), .A(\g.we_clk [28433]));
Q_ASSIGN U4342 ( .B(clk), .A(\g.we_clk [28432]));
Q_ASSIGN U4343 ( .B(clk), .A(\g.we_clk [28431]));
Q_ASSIGN U4344 ( .B(clk), .A(\g.we_clk [28430]));
Q_ASSIGN U4345 ( .B(clk), .A(\g.we_clk [28429]));
Q_ASSIGN U4346 ( .B(clk), .A(\g.we_clk [28428]));
Q_ASSIGN U4347 ( .B(clk), .A(\g.we_clk [28427]));
Q_ASSIGN U4348 ( .B(clk), .A(\g.we_clk [28426]));
Q_ASSIGN U4349 ( .B(clk), .A(\g.we_clk [28425]));
Q_ASSIGN U4350 ( .B(clk), .A(\g.we_clk [28424]));
Q_ASSIGN U4351 ( .B(clk), .A(\g.we_clk [28423]));
Q_ASSIGN U4352 ( .B(clk), .A(\g.we_clk [28422]));
Q_ASSIGN U4353 ( .B(clk), .A(\g.we_clk [28421]));
Q_ASSIGN U4354 ( .B(clk), .A(\g.we_clk [28420]));
Q_ASSIGN U4355 ( .B(clk), .A(\g.we_clk [28419]));
Q_ASSIGN U4356 ( .B(clk), .A(\g.we_clk [28418]));
Q_ASSIGN U4357 ( .B(clk), .A(\g.we_clk [28417]));
Q_ASSIGN U4358 ( .B(clk), .A(\g.we_clk [28416]));
Q_ASSIGN U4359 ( .B(clk), .A(\g.we_clk [28415]));
Q_ASSIGN U4360 ( .B(clk), .A(\g.we_clk [28414]));
Q_ASSIGN U4361 ( .B(clk), .A(\g.we_clk [28413]));
Q_ASSIGN U4362 ( .B(clk), .A(\g.we_clk [28412]));
Q_ASSIGN U4363 ( .B(clk), .A(\g.we_clk [28411]));
Q_ASSIGN U4364 ( .B(clk), .A(\g.we_clk [28410]));
Q_ASSIGN U4365 ( .B(clk), .A(\g.we_clk [28409]));
Q_ASSIGN U4366 ( .B(clk), .A(\g.we_clk [28408]));
Q_ASSIGN U4367 ( .B(clk), .A(\g.we_clk [28407]));
Q_ASSIGN U4368 ( .B(clk), .A(\g.we_clk [28406]));
Q_ASSIGN U4369 ( .B(clk), .A(\g.we_clk [28405]));
Q_ASSIGN U4370 ( .B(clk), .A(\g.we_clk [28404]));
Q_ASSIGN U4371 ( .B(clk), .A(\g.we_clk [28403]));
Q_ASSIGN U4372 ( .B(clk), .A(\g.we_clk [28402]));
Q_ASSIGN U4373 ( .B(clk), .A(\g.we_clk [28401]));
Q_ASSIGN U4374 ( .B(clk), .A(\g.we_clk [28400]));
Q_ASSIGN U4375 ( .B(clk), .A(\g.we_clk [28399]));
Q_ASSIGN U4376 ( .B(clk), .A(\g.we_clk [28398]));
Q_ASSIGN U4377 ( .B(clk), .A(\g.we_clk [28397]));
Q_ASSIGN U4378 ( .B(clk), .A(\g.we_clk [28396]));
Q_ASSIGN U4379 ( .B(clk), .A(\g.we_clk [28395]));
Q_ASSIGN U4380 ( .B(clk), .A(\g.we_clk [28394]));
Q_ASSIGN U4381 ( .B(clk), .A(\g.we_clk [28393]));
Q_ASSIGN U4382 ( .B(clk), .A(\g.we_clk [28392]));
Q_ASSIGN U4383 ( .B(clk), .A(\g.we_clk [28391]));
Q_ASSIGN U4384 ( .B(clk), .A(\g.we_clk [28390]));
Q_ASSIGN U4385 ( .B(clk), .A(\g.we_clk [28389]));
Q_ASSIGN U4386 ( .B(clk), .A(\g.we_clk [28388]));
Q_ASSIGN U4387 ( .B(clk), .A(\g.we_clk [28387]));
Q_ASSIGN U4388 ( .B(clk), .A(\g.we_clk [28386]));
Q_ASSIGN U4389 ( .B(clk), .A(\g.we_clk [28385]));
Q_ASSIGN U4390 ( .B(clk), .A(\g.we_clk [28384]));
Q_ASSIGN U4391 ( .B(clk), .A(\g.we_clk [28383]));
Q_ASSIGN U4392 ( .B(clk), .A(\g.we_clk [28382]));
Q_ASSIGN U4393 ( .B(clk), .A(\g.we_clk [28381]));
Q_ASSIGN U4394 ( .B(clk), .A(\g.we_clk [28380]));
Q_ASSIGN U4395 ( .B(clk), .A(\g.we_clk [28379]));
Q_ASSIGN U4396 ( .B(clk), .A(\g.we_clk [28378]));
Q_ASSIGN U4397 ( .B(clk), .A(\g.we_clk [28377]));
Q_ASSIGN U4398 ( .B(clk), .A(\g.we_clk [28376]));
Q_ASSIGN U4399 ( .B(clk), .A(\g.we_clk [28375]));
Q_ASSIGN U4400 ( .B(clk), .A(\g.we_clk [28374]));
Q_ASSIGN U4401 ( .B(clk), .A(\g.we_clk [28373]));
Q_ASSIGN U4402 ( .B(clk), .A(\g.we_clk [28372]));
Q_ASSIGN U4403 ( .B(clk), .A(\g.we_clk [28371]));
Q_ASSIGN U4404 ( .B(clk), .A(\g.we_clk [28370]));
Q_ASSIGN U4405 ( .B(clk), .A(\g.we_clk [28369]));
Q_ASSIGN U4406 ( .B(clk), .A(\g.we_clk [28368]));
Q_ASSIGN U4407 ( .B(clk), .A(\g.we_clk [28367]));
Q_ASSIGN U4408 ( .B(clk), .A(\g.we_clk [28366]));
Q_ASSIGN U4409 ( .B(clk), .A(\g.we_clk [28365]));
Q_ASSIGN U4410 ( .B(clk), .A(\g.we_clk [28364]));
Q_ASSIGN U4411 ( .B(clk), .A(\g.we_clk [28363]));
Q_ASSIGN U4412 ( .B(clk), .A(\g.we_clk [28362]));
Q_ASSIGN U4413 ( .B(clk), .A(\g.we_clk [28361]));
Q_ASSIGN U4414 ( .B(clk), .A(\g.we_clk [28360]));
Q_ASSIGN U4415 ( .B(clk), .A(\g.we_clk [28359]));
Q_ASSIGN U4416 ( .B(clk), .A(\g.we_clk [28358]));
Q_ASSIGN U4417 ( .B(clk), .A(\g.we_clk [28357]));
Q_ASSIGN U4418 ( .B(clk), .A(\g.we_clk [28356]));
Q_ASSIGN U4419 ( .B(clk), .A(\g.we_clk [28355]));
Q_ASSIGN U4420 ( .B(clk), .A(\g.we_clk [28354]));
Q_ASSIGN U4421 ( .B(clk), .A(\g.we_clk [28353]));
Q_ASSIGN U4422 ( .B(clk), .A(\g.we_clk [28352]));
Q_ASSIGN U4423 ( .B(clk), .A(\g.we_clk [28351]));
Q_ASSIGN U4424 ( .B(clk), .A(\g.we_clk [28350]));
Q_ASSIGN U4425 ( .B(clk), .A(\g.we_clk [28349]));
Q_ASSIGN U4426 ( .B(clk), .A(\g.we_clk [28348]));
Q_ASSIGN U4427 ( .B(clk), .A(\g.we_clk [28347]));
Q_ASSIGN U4428 ( .B(clk), .A(\g.we_clk [28346]));
Q_ASSIGN U4429 ( .B(clk), .A(\g.we_clk [28345]));
Q_ASSIGN U4430 ( .B(clk), .A(\g.we_clk [28344]));
Q_ASSIGN U4431 ( .B(clk), .A(\g.we_clk [28343]));
Q_ASSIGN U4432 ( .B(clk), .A(\g.we_clk [28342]));
Q_ASSIGN U4433 ( .B(clk), .A(\g.we_clk [28341]));
Q_ASSIGN U4434 ( .B(clk), .A(\g.we_clk [28340]));
Q_ASSIGN U4435 ( .B(clk), .A(\g.we_clk [28339]));
Q_ASSIGN U4436 ( .B(clk), .A(\g.we_clk [28338]));
Q_ASSIGN U4437 ( .B(clk), .A(\g.we_clk [28337]));
Q_ASSIGN U4438 ( .B(clk), .A(\g.we_clk [28336]));
Q_ASSIGN U4439 ( .B(clk), .A(\g.we_clk [28335]));
Q_ASSIGN U4440 ( .B(clk), .A(\g.we_clk [28334]));
Q_ASSIGN U4441 ( .B(clk), .A(\g.we_clk [28333]));
Q_ASSIGN U4442 ( .B(clk), .A(\g.we_clk [28332]));
Q_ASSIGN U4443 ( .B(clk), .A(\g.we_clk [28331]));
Q_ASSIGN U4444 ( .B(clk), .A(\g.we_clk [28330]));
Q_ASSIGN U4445 ( .B(clk), .A(\g.we_clk [28329]));
Q_ASSIGN U4446 ( .B(clk), .A(\g.we_clk [28328]));
Q_ASSIGN U4447 ( .B(clk), .A(\g.we_clk [28327]));
Q_ASSIGN U4448 ( .B(clk), .A(\g.we_clk [28326]));
Q_ASSIGN U4449 ( .B(clk), .A(\g.we_clk [28325]));
Q_ASSIGN U4450 ( .B(clk), .A(\g.we_clk [28324]));
Q_ASSIGN U4451 ( .B(clk), .A(\g.we_clk [28323]));
Q_ASSIGN U4452 ( .B(clk), .A(\g.we_clk [28322]));
Q_ASSIGN U4453 ( .B(clk), .A(\g.we_clk [28321]));
Q_ASSIGN U4454 ( .B(clk), .A(\g.we_clk [28320]));
Q_ASSIGN U4455 ( .B(clk), .A(\g.we_clk [28319]));
Q_ASSIGN U4456 ( .B(clk), .A(\g.we_clk [28318]));
Q_ASSIGN U4457 ( .B(clk), .A(\g.we_clk [28317]));
Q_ASSIGN U4458 ( .B(clk), .A(\g.we_clk [28316]));
Q_ASSIGN U4459 ( .B(clk), .A(\g.we_clk [28315]));
Q_ASSIGN U4460 ( .B(clk), .A(\g.we_clk [28314]));
Q_ASSIGN U4461 ( .B(clk), .A(\g.we_clk [28313]));
Q_ASSIGN U4462 ( .B(clk), .A(\g.we_clk [28312]));
Q_ASSIGN U4463 ( .B(clk), .A(\g.we_clk [28311]));
Q_ASSIGN U4464 ( .B(clk), .A(\g.we_clk [28310]));
Q_ASSIGN U4465 ( .B(clk), .A(\g.we_clk [28309]));
Q_ASSIGN U4466 ( .B(clk), .A(\g.we_clk [28308]));
Q_ASSIGN U4467 ( .B(clk), .A(\g.we_clk [28307]));
Q_ASSIGN U4468 ( .B(clk), .A(\g.we_clk [28306]));
Q_ASSIGN U4469 ( .B(clk), .A(\g.we_clk [28305]));
Q_ASSIGN U4470 ( .B(clk), .A(\g.we_clk [28304]));
Q_ASSIGN U4471 ( .B(clk), .A(\g.we_clk [28303]));
Q_ASSIGN U4472 ( .B(clk), .A(\g.we_clk [28302]));
Q_ASSIGN U4473 ( .B(clk), .A(\g.we_clk [28301]));
Q_ASSIGN U4474 ( .B(clk), .A(\g.we_clk [28300]));
Q_ASSIGN U4475 ( .B(clk), .A(\g.we_clk [28299]));
Q_ASSIGN U4476 ( .B(clk), .A(\g.we_clk [28298]));
Q_ASSIGN U4477 ( .B(clk), .A(\g.we_clk [28297]));
Q_ASSIGN U4478 ( .B(clk), .A(\g.we_clk [28296]));
Q_ASSIGN U4479 ( .B(clk), .A(\g.we_clk [28295]));
Q_ASSIGN U4480 ( .B(clk), .A(\g.we_clk [28294]));
Q_ASSIGN U4481 ( .B(clk), .A(\g.we_clk [28293]));
Q_ASSIGN U4482 ( .B(clk), .A(\g.we_clk [28292]));
Q_ASSIGN U4483 ( .B(clk), .A(\g.we_clk [28291]));
Q_ASSIGN U4484 ( .B(clk), .A(\g.we_clk [28290]));
Q_ASSIGN U4485 ( .B(clk), .A(\g.we_clk [28289]));
Q_ASSIGN U4486 ( .B(clk), .A(\g.we_clk [28288]));
Q_ASSIGN U4487 ( .B(clk), .A(\g.we_clk [28287]));
Q_ASSIGN U4488 ( .B(clk), .A(\g.we_clk [28286]));
Q_ASSIGN U4489 ( .B(clk), .A(\g.we_clk [28285]));
Q_ASSIGN U4490 ( .B(clk), .A(\g.we_clk [28284]));
Q_ASSIGN U4491 ( .B(clk), .A(\g.we_clk [28283]));
Q_ASSIGN U4492 ( .B(clk), .A(\g.we_clk [28282]));
Q_ASSIGN U4493 ( .B(clk), .A(\g.we_clk [28281]));
Q_ASSIGN U4494 ( .B(clk), .A(\g.we_clk [28280]));
Q_ASSIGN U4495 ( .B(clk), .A(\g.we_clk [28279]));
Q_ASSIGN U4496 ( .B(clk), .A(\g.we_clk [28278]));
Q_ASSIGN U4497 ( .B(clk), .A(\g.we_clk [28277]));
Q_ASSIGN U4498 ( .B(clk), .A(\g.we_clk [28276]));
Q_ASSIGN U4499 ( .B(clk), .A(\g.we_clk [28275]));
Q_ASSIGN U4500 ( .B(clk), .A(\g.we_clk [28274]));
Q_ASSIGN U4501 ( .B(clk), .A(\g.we_clk [28273]));
Q_ASSIGN U4502 ( .B(clk), .A(\g.we_clk [28272]));
Q_ASSIGN U4503 ( .B(clk), .A(\g.we_clk [28271]));
Q_ASSIGN U4504 ( .B(clk), .A(\g.we_clk [28270]));
Q_ASSIGN U4505 ( .B(clk), .A(\g.we_clk [28269]));
Q_ASSIGN U4506 ( .B(clk), .A(\g.we_clk [28268]));
Q_ASSIGN U4507 ( .B(clk), .A(\g.we_clk [28267]));
Q_ASSIGN U4508 ( .B(clk), .A(\g.we_clk [28266]));
Q_ASSIGN U4509 ( .B(clk), .A(\g.we_clk [28265]));
Q_ASSIGN U4510 ( .B(clk), .A(\g.we_clk [28264]));
Q_ASSIGN U4511 ( .B(clk), .A(\g.we_clk [28263]));
Q_ASSIGN U4512 ( .B(clk), .A(\g.we_clk [28262]));
Q_ASSIGN U4513 ( .B(clk), .A(\g.we_clk [28261]));
Q_ASSIGN U4514 ( .B(clk), .A(\g.we_clk [28260]));
Q_ASSIGN U4515 ( .B(clk), .A(\g.we_clk [28259]));
Q_ASSIGN U4516 ( .B(clk), .A(\g.we_clk [28258]));
Q_ASSIGN U4517 ( .B(clk), .A(\g.we_clk [28257]));
Q_ASSIGN U4518 ( .B(clk), .A(\g.we_clk [28256]));
Q_ASSIGN U4519 ( .B(clk), .A(\g.we_clk [28255]));
Q_ASSIGN U4520 ( .B(clk), .A(\g.we_clk [28254]));
Q_ASSIGN U4521 ( .B(clk), .A(\g.we_clk [28253]));
Q_ASSIGN U4522 ( .B(clk), .A(\g.we_clk [28252]));
Q_ASSIGN U4523 ( .B(clk), .A(\g.we_clk [28251]));
Q_ASSIGN U4524 ( .B(clk), .A(\g.we_clk [28250]));
Q_ASSIGN U4525 ( .B(clk), .A(\g.we_clk [28249]));
Q_ASSIGN U4526 ( .B(clk), .A(\g.we_clk [28248]));
Q_ASSIGN U4527 ( .B(clk), .A(\g.we_clk [28247]));
Q_ASSIGN U4528 ( .B(clk), .A(\g.we_clk [28246]));
Q_ASSIGN U4529 ( .B(clk), .A(\g.we_clk [28245]));
Q_ASSIGN U4530 ( .B(clk), .A(\g.we_clk [28244]));
Q_ASSIGN U4531 ( .B(clk), .A(\g.we_clk [28243]));
Q_ASSIGN U4532 ( .B(clk), .A(\g.we_clk [28242]));
Q_ASSIGN U4533 ( .B(clk), .A(\g.we_clk [28241]));
Q_ASSIGN U4534 ( .B(clk), .A(\g.we_clk [28240]));
Q_ASSIGN U4535 ( .B(clk), .A(\g.we_clk [28239]));
Q_ASSIGN U4536 ( .B(clk), .A(\g.we_clk [28238]));
Q_ASSIGN U4537 ( .B(clk), .A(\g.we_clk [28237]));
Q_ASSIGN U4538 ( .B(clk), .A(\g.we_clk [28236]));
Q_ASSIGN U4539 ( .B(clk), .A(\g.we_clk [28235]));
Q_ASSIGN U4540 ( .B(clk), .A(\g.we_clk [28234]));
Q_ASSIGN U4541 ( .B(clk), .A(\g.we_clk [28233]));
Q_ASSIGN U4542 ( .B(clk), .A(\g.we_clk [28232]));
Q_ASSIGN U4543 ( .B(clk), .A(\g.we_clk [28231]));
Q_ASSIGN U4544 ( .B(clk), .A(\g.we_clk [28230]));
Q_ASSIGN U4545 ( .B(clk), .A(\g.we_clk [28229]));
Q_ASSIGN U4546 ( .B(clk), .A(\g.we_clk [28228]));
Q_ASSIGN U4547 ( .B(clk), .A(\g.we_clk [28227]));
Q_ASSIGN U4548 ( .B(clk), .A(\g.we_clk [28226]));
Q_ASSIGN U4549 ( .B(clk), .A(\g.we_clk [28225]));
Q_ASSIGN U4550 ( .B(clk), .A(\g.we_clk [28224]));
Q_ASSIGN U4551 ( .B(clk), .A(\g.we_clk [28223]));
Q_ASSIGN U4552 ( .B(clk), .A(\g.we_clk [28222]));
Q_ASSIGN U4553 ( .B(clk), .A(\g.we_clk [28221]));
Q_ASSIGN U4554 ( .B(clk), .A(\g.we_clk [28220]));
Q_ASSIGN U4555 ( .B(clk), .A(\g.we_clk [28219]));
Q_ASSIGN U4556 ( .B(clk), .A(\g.we_clk [28218]));
Q_ASSIGN U4557 ( .B(clk), .A(\g.we_clk [28217]));
Q_ASSIGN U4558 ( .B(clk), .A(\g.we_clk [28216]));
Q_ASSIGN U4559 ( .B(clk), .A(\g.we_clk [28215]));
Q_ASSIGN U4560 ( .B(clk), .A(\g.we_clk [28214]));
Q_ASSIGN U4561 ( .B(clk), .A(\g.we_clk [28213]));
Q_ASSIGN U4562 ( .B(clk), .A(\g.we_clk [28212]));
Q_ASSIGN U4563 ( .B(clk), .A(\g.we_clk [28211]));
Q_ASSIGN U4564 ( .B(clk), .A(\g.we_clk [28210]));
Q_ASSIGN U4565 ( .B(clk), .A(\g.we_clk [28209]));
Q_ASSIGN U4566 ( .B(clk), .A(\g.we_clk [28208]));
Q_ASSIGN U4567 ( .B(clk), .A(\g.we_clk [28207]));
Q_ASSIGN U4568 ( .B(clk), .A(\g.we_clk [28206]));
Q_ASSIGN U4569 ( .B(clk), .A(\g.we_clk [28205]));
Q_ASSIGN U4570 ( .B(clk), .A(\g.we_clk [28204]));
Q_ASSIGN U4571 ( .B(clk), .A(\g.we_clk [28203]));
Q_ASSIGN U4572 ( .B(clk), .A(\g.we_clk [28202]));
Q_ASSIGN U4573 ( .B(clk), .A(\g.we_clk [28201]));
Q_ASSIGN U4574 ( .B(clk), .A(\g.we_clk [28200]));
Q_ASSIGN U4575 ( .B(clk), .A(\g.we_clk [28199]));
Q_ASSIGN U4576 ( .B(clk), .A(\g.we_clk [28198]));
Q_ASSIGN U4577 ( .B(clk), .A(\g.we_clk [28197]));
Q_ASSIGN U4578 ( .B(clk), .A(\g.we_clk [28196]));
Q_ASSIGN U4579 ( .B(clk), .A(\g.we_clk [28195]));
Q_ASSIGN U4580 ( .B(clk), .A(\g.we_clk [28194]));
Q_ASSIGN U4581 ( .B(clk), .A(\g.we_clk [28193]));
Q_ASSIGN U4582 ( .B(clk), .A(\g.we_clk [28192]));
Q_ASSIGN U4583 ( .B(clk), .A(\g.we_clk [28191]));
Q_ASSIGN U4584 ( .B(clk), .A(\g.we_clk [28190]));
Q_ASSIGN U4585 ( .B(clk), .A(\g.we_clk [28189]));
Q_ASSIGN U4586 ( .B(clk), .A(\g.we_clk [28188]));
Q_ASSIGN U4587 ( .B(clk), .A(\g.we_clk [28187]));
Q_ASSIGN U4588 ( .B(clk), .A(\g.we_clk [28186]));
Q_ASSIGN U4589 ( .B(clk), .A(\g.we_clk [28185]));
Q_ASSIGN U4590 ( .B(clk), .A(\g.we_clk [28184]));
Q_ASSIGN U4591 ( .B(clk), .A(\g.we_clk [28183]));
Q_ASSIGN U4592 ( .B(clk), .A(\g.we_clk [28182]));
Q_ASSIGN U4593 ( .B(clk), .A(\g.we_clk [28181]));
Q_ASSIGN U4594 ( .B(clk), .A(\g.we_clk [28180]));
Q_ASSIGN U4595 ( .B(clk), .A(\g.we_clk [28179]));
Q_ASSIGN U4596 ( .B(clk), .A(\g.we_clk [28178]));
Q_ASSIGN U4597 ( .B(clk), .A(\g.we_clk [28177]));
Q_ASSIGN U4598 ( .B(clk), .A(\g.we_clk [28176]));
Q_ASSIGN U4599 ( .B(clk), .A(\g.we_clk [28175]));
Q_ASSIGN U4600 ( .B(clk), .A(\g.we_clk [28174]));
Q_ASSIGN U4601 ( .B(clk), .A(\g.we_clk [28173]));
Q_ASSIGN U4602 ( .B(clk), .A(\g.we_clk [28172]));
Q_ASSIGN U4603 ( .B(clk), .A(\g.we_clk [28171]));
Q_ASSIGN U4604 ( .B(clk), .A(\g.we_clk [28170]));
Q_ASSIGN U4605 ( .B(clk), .A(\g.we_clk [28169]));
Q_ASSIGN U4606 ( .B(clk), .A(\g.we_clk [28168]));
Q_ASSIGN U4607 ( .B(clk), .A(\g.we_clk [28167]));
Q_ASSIGN U4608 ( .B(clk), .A(\g.we_clk [28166]));
Q_ASSIGN U4609 ( .B(clk), .A(\g.we_clk [28165]));
Q_ASSIGN U4610 ( .B(clk), .A(\g.we_clk [28164]));
Q_ASSIGN U4611 ( .B(clk), .A(\g.we_clk [28163]));
Q_ASSIGN U4612 ( .B(clk), .A(\g.we_clk [28162]));
Q_ASSIGN U4613 ( .B(clk), .A(\g.we_clk [28161]));
Q_ASSIGN U4614 ( .B(clk), .A(\g.we_clk [28160]));
Q_ASSIGN U4615 ( .B(clk), .A(\g.we_clk [28159]));
Q_ASSIGN U4616 ( .B(clk), .A(\g.we_clk [28158]));
Q_ASSIGN U4617 ( .B(clk), .A(\g.we_clk [28157]));
Q_ASSIGN U4618 ( .B(clk), .A(\g.we_clk [28156]));
Q_ASSIGN U4619 ( .B(clk), .A(\g.we_clk [28155]));
Q_ASSIGN U4620 ( .B(clk), .A(\g.we_clk [28154]));
Q_ASSIGN U4621 ( .B(clk), .A(\g.we_clk [28153]));
Q_ASSIGN U4622 ( .B(clk), .A(\g.we_clk [28152]));
Q_ASSIGN U4623 ( .B(clk), .A(\g.we_clk [28151]));
Q_ASSIGN U4624 ( .B(clk), .A(\g.we_clk [28150]));
Q_ASSIGN U4625 ( .B(clk), .A(\g.we_clk [28149]));
Q_ASSIGN U4626 ( .B(clk), .A(\g.we_clk [28148]));
Q_ASSIGN U4627 ( .B(clk), .A(\g.we_clk [28147]));
Q_ASSIGN U4628 ( .B(clk), .A(\g.we_clk [28146]));
Q_ASSIGN U4629 ( .B(clk), .A(\g.we_clk [28145]));
Q_ASSIGN U4630 ( .B(clk), .A(\g.we_clk [28144]));
Q_ASSIGN U4631 ( .B(clk), .A(\g.we_clk [28143]));
Q_ASSIGN U4632 ( .B(clk), .A(\g.we_clk [28142]));
Q_ASSIGN U4633 ( .B(clk), .A(\g.we_clk [28141]));
Q_ASSIGN U4634 ( .B(clk), .A(\g.we_clk [28140]));
Q_ASSIGN U4635 ( .B(clk), .A(\g.we_clk [28139]));
Q_ASSIGN U4636 ( .B(clk), .A(\g.we_clk [28138]));
Q_ASSIGN U4637 ( .B(clk), .A(\g.we_clk [28137]));
Q_ASSIGN U4638 ( .B(clk), .A(\g.we_clk [28136]));
Q_ASSIGN U4639 ( .B(clk), .A(\g.we_clk [28135]));
Q_ASSIGN U4640 ( .B(clk), .A(\g.we_clk [28134]));
Q_ASSIGN U4641 ( .B(clk), .A(\g.we_clk [28133]));
Q_ASSIGN U4642 ( .B(clk), .A(\g.we_clk [28132]));
Q_ASSIGN U4643 ( .B(clk), .A(\g.we_clk [28131]));
Q_ASSIGN U4644 ( .B(clk), .A(\g.we_clk [28130]));
Q_ASSIGN U4645 ( .B(clk), .A(\g.we_clk [28129]));
Q_ASSIGN U4646 ( .B(clk), .A(\g.we_clk [28128]));
Q_ASSIGN U4647 ( .B(clk), .A(\g.we_clk [28127]));
Q_ASSIGN U4648 ( .B(clk), .A(\g.we_clk [28126]));
Q_ASSIGN U4649 ( .B(clk), .A(\g.we_clk [28125]));
Q_ASSIGN U4650 ( .B(clk), .A(\g.we_clk [28124]));
Q_ASSIGN U4651 ( .B(clk), .A(\g.we_clk [28123]));
Q_ASSIGN U4652 ( .B(clk), .A(\g.we_clk [28122]));
Q_ASSIGN U4653 ( .B(clk), .A(\g.we_clk [28121]));
Q_ASSIGN U4654 ( .B(clk), .A(\g.we_clk [28120]));
Q_ASSIGN U4655 ( .B(clk), .A(\g.we_clk [28119]));
Q_ASSIGN U4656 ( .B(clk), .A(\g.we_clk [28118]));
Q_ASSIGN U4657 ( .B(clk), .A(\g.we_clk [28117]));
Q_ASSIGN U4658 ( .B(clk), .A(\g.we_clk [28116]));
Q_ASSIGN U4659 ( .B(clk), .A(\g.we_clk [28115]));
Q_ASSIGN U4660 ( .B(clk), .A(\g.we_clk [28114]));
Q_ASSIGN U4661 ( .B(clk), .A(\g.we_clk [28113]));
Q_ASSIGN U4662 ( .B(clk), .A(\g.we_clk [28112]));
Q_ASSIGN U4663 ( .B(clk), .A(\g.we_clk [28111]));
Q_ASSIGN U4664 ( .B(clk), .A(\g.we_clk [28110]));
Q_ASSIGN U4665 ( .B(clk), .A(\g.we_clk [28109]));
Q_ASSIGN U4666 ( .B(clk), .A(\g.we_clk [28108]));
Q_ASSIGN U4667 ( .B(clk), .A(\g.we_clk [28107]));
Q_ASSIGN U4668 ( .B(clk), .A(\g.we_clk [28106]));
Q_ASSIGN U4669 ( .B(clk), .A(\g.we_clk [28105]));
Q_ASSIGN U4670 ( .B(clk), .A(\g.we_clk [28104]));
Q_ASSIGN U4671 ( .B(clk), .A(\g.we_clk [28103]));
Q_ASSIGN U4672 ( .B(clk), .A(\g.we_clk [28102]));
Q_ASSIGN U4673 ( .B(clk), .A(\g.we_clk [28101]));
Q_ASSIGN U4674 ( .B(clk), .A(\g.we_clk [28100]));
Q_ASSIGN U4675 ( .B(clk), .A(\g.we_clk [28099]));
Q_ASSIGN U4676 ( .B(clk), .A(\g.we_clk [28098]));
Q_ASSIGN U4677 ( .B(clk), .A(\g.we_clk [28097]));
Q_ASSIGN U4678 ( .B(clk), .A(\g.we_clk [28096]));
Q_ASSIGN U4679 ( .B(clk), .A(\g.we_clk [28095]));
Q_ASSIGN U4680 ( .B(clk), .A(\g.we_clk [28094]));
Q_ASSIGN U4681 ( .B(clk), .A(\g.we_clk [28093]));
Q_ASSIGN U4682 ( .B(clk), .A(\g.we_clk [28092]));
Q_ASSIGN U4683 ( .B(clk), .A(\g.we_clk [28091]));
Q_ASSIGN U4684 ( .B(clk), .A(\g.we_clk [28090]));
Q_ASSIGN U4685 ( .B(clk), .A(\g.we_clk [28089]));
Q_ASSIGN U4686 ( .B(clk), .A(\g.we_clk [28088]));
Q_ASSIGN U4687 ( .B(clk), .A(\g.we_clk [28087]));
Q_ASSIGN U4688 ( .B(clk), .A(\g.we_clk [28086]));
Q_ASSIGN U4689 ( .B(clk), .A(\g.we_clk [28085]));
Q_ASSIGN U4690 ( .B(clk), .A(\g.we_clk [28084]));
Q_ASSIGN U4691 ( .B(clk), .A(\g.we_clk [28083]));
Q_ASSIGN U4692 ( .B(clk), .A(\g.we_clk [28082]));
Q_ASSIGN U4693 ( .B(clk), .A(\g.we_clk [28081]));
Q_ASSIGN U4694 ( .B(clk), .A(\g.we_clk [28080]));
Q_ASSIGN U4695 ( .B(clk), .A(\g.we_clk [28079]));
Q_ASSIGN U4696 ( .B(clk), .A(\g.we_clk [28078]));
Q_ASSIGN U4697 ( .B(clk), .A(\g.we_clk [28077]));
Q_ASSIGN U4698 ( .B(clk), .A(\g.we_clk [28076]));
Q_ASSIGN U4699 ( .B(clk), .A(\g.we_clk [28075]));
Q_ASSIGN U4700 ( .B(clk), .A(\g.we_clk [28074]));
Q_ASSIGN U4701 ( .B(clk), .A(\g.we_clk [28073]));
Q_ASSIGN U4702 ( .B(clk), .A(\g.we_clk [28072]));
Q_ASSIGN U4703 ( .B(clk), .A(\g.we_clk [28071]));
Q_ASSIGN U4704 ( .B(clk), .A(\g.we_clk [28070]));
Q_ASSIGN U4705 ( .B(clk), .A(\g.we_clk [28069]));
Q_ASSIGN U4706 ( .B(clk), .A(\g.we_clk [28068]));
Q_ASSIGN U4707 ( .B(clk), .A(\g.we_clk [28067]));
Q_ASSIGN U4708 ( .B(clk), .A(\g.we_clk [28066]));
Q_ASSIGN U4709 ( .B(clk), .A(\g.we_clk [28065]));
Q_ASSIGN U4710 ( .B(clk), .A(\g.we_clk [28064]));
Q_ASSIGN U4711 ( .B(clk), .A(\g.we_clk [28063]));
Q_ASSIGN U4712 ( .B(clk), .A(\g.we_clk [28062]));
Q_ASSIGN U4713 ( .B(clk), .A(\g.we_clk [28061]));
Q_ASSIGN U4714 ( .B(clk), .A(\g.we_clk [28060]));
Q_ASSIGN U4715 ( .B(clk), .A(\g.we_clk [28059]));
Q_ASSIGN U4716 ( .B(clk), .A(\g.we_clk [28058]));
Q_ASSIGN U4717 ( .B(clk), .A(\g.we_clk [28057]));
Q_ASSIGN U4718 ( .B(clk), .A(\g.we_clk [28056]));
Q_ASSIGN U4719 ( .B(clk), .A(\g.we_clk [28055]));
Q_ASSIGN U4720 ( .B(clk), .A(\g.we_clk [28054]));
Q_ASSIGN U4721 ( .B(clk), .A(\g.we_clk [28053]));
Q_ASSIGN U4722 ( .B(clk), .A(\g.we_clk [28052]));
Q_ASSIGN U4723 ( .B(clk), .A(\g.we_clk [28051]));
Q_ASSIGN U4724 ( .B(clk), .A(\g.we_clk [28050]));
Q_ASSIGN U4725 ( .B(clk), .A(\g.we_clk [28049]));
Q_ASSIGN U4726 ( .B(clk), .A(\g.we_clk [28048]));
Q_ASSIGN U4727 ( .B(clk), .A(\g.we_clk [28047]));
Q_ASSIGN U4728 ( .B(clk), .A(\g.we_clk [28046]));
Q_ASSIGN U4729 ( .B(clk), .A(\g.we_clk [28045]));
Q_ASSIGN U4730 ( .B(clk), .A(\g.we_clk [28044]));
Q_ASSIGN U4731 ( .B(clk), .A(\g.we_clk [28043]));
Q_ASSIGN U4732 ( .B(clk), .A(\g.we_clk [28042]));
Q_ASSIGN U4733 ( .B(clk), .A(\g.we_clk [28041]));
Q_ASSIGN U4734 ( .B(clk), .A(\g.we_clk [28040]));
Q_ASSIGN U4735 ( .B(clk), .A(\g.we_clk [28039]));
Q_ASSIGN U4736 ( .B(clk), .A(\g.we_clk [28038]));
Q_ASSIGN U4737 ( .B(clk), .A(\g.we_clk [28037]));
Q_ASSIGN U4738 ( .B(clk), .A(\g.we_clk [28036]));
Q_ASSIGN U4739 ( .B(clk), .A(\g.we_clk [28035]));
Q_ASSIGN U4740 ( .B(clk), .A(\g.we_clk [28034]));
Q_ASSIGN U4741 ( .B(clk), .A(\g.we_clk [28033]));
Q_ASSIGN U4742 ( .B(clk), .A(\g.we_clk [28032]));
Q_ASSIGN U4743 ( .B(clk), .A(\g.we_clk [28031]));
Q_ASSIGN U4744 ( .B(clk), .A(\g.we_clk [28030]));
Q_ASSIGN U4745 ( .B(clk), .A(\g.we_clk [28029]));
Q_ASSIGN U4746 ( .B(clk), .A(\g.we_clk [28028]));
Q_ASSIGN U4747 ( .B(clk), .A(\g.we_clk [28027]));
Q_ASSIGN U4748 ( .B(clk), .A(\g.we_clk [28026]));
Q_ASSIGN U4749 ( .B(clk), .A(\g.we_clk [28025]));
Q_ASSIGN U4750 ( .B(clk), .A(\g.we_clk [28024]));
Q_ASSIGN U4751 ( .B(clk), .A(\g.we_clk [28023]));
Q_ASSIGN U4752 ( .B(clk), .A(\g.we_clk [28022]));
Q_ASSIGN U4753 ( .B(clk), .A(\g.we_clk [28021]));
Q_ASSIGN U4754 ( .B(clk), .A(\g.we_clk [28020]));
Q_ASSIGN U4755 ( .B(clk), .A(\g.we_clk [28019]));
Q_ASSIGN U4756 ( .B(clk), .A(\g.we_clk [28018]));
Q_ASSIGN U4757 ( .B(clk), .A(\g.we_clk [28017]));
Q_ASSIGN U4758 ( .B(clk), .A(\g.we_clk [28016]));
Q_ASSIGN U4759 ( .B(clk), .A(\g.we_clk [28015]));
Q_ASSIGN U4760 ( .B(clk), .A(\g.we_clk [28014]));
Q_ASSIGN U4761 ( .B(clk), .A(\g.we_clk [28013]));
Q_ASSIGN U4762 ( .B(clk), .A(\g.we_clk [28012]));
Q_ASSIGN U4763 ( .B(clk), .A(\g.we_clk [28011]));
Q_ASSIGN U4764 ( .B(clk), .A(\g.we_clk [28010]));
Q_ASSIGN U4765 ( .B(clk), .A(\g.we_clk [28009]));
Q_ASSIGN U4766 ( .B(clk), .A(\g.we_clk [28008]));
Q_ASSIGN U4767 ( .B(clk), .A(\g.we_clk [28007]));
Q_ASSIGN U4768 ( .B(clk), .A(\g.we_clk [28006]));
Q_ASSIGN U4769 ( .B(clk), .A(\g.we_clk [28005]));
Q_ASSIGN U4770 ( .B(clk), .A(\g.we_clk [28004]));
Q_ASSIGN U4771 ( .B(clk), .A(\g.we_clk [28003]));
Q_ASSIGN U4772 ( .B(clk), .A(\g.we_clk [28002]));
Q_ASSIGN U4773 ( .B(clk), .A(\g.we_clk [28001]));
Q_ASSIGN U4774 ( .B(clk), .A(\g.we_clk [28000]));
Q_ASSIGN U4775 ( .B(clk), .A(\g.we_clk [27999]));
Q_ASSIGN U4776 ( .B(clk), .A(\g.we_clk [27998]));
Q_ASSIGN U4777 ( .B(clk), .A(\g.we_clk [27997]));
Q_ASSIGN U4778 ( .B(clk), .A(\g.we_clk [27996]));
Q_ASSIGN U4779 ( .B(clk), .A(\g.we_clk [27995]));
Q_ASSIGN U4780 ( .B(clk), .A(\g.we_clk [27994]));
Q_ASSIGN U4781 ( .B(clk), .A(\g.we_clk [27993]));
Q_ASSIGN U4782 ( .B(clk), .A(\g.we_clk [27992]));
Q_ASSIGN U4783 ( .B(clk), .A(\g.we_clk [27991]));
Q_ASSIGN U4784 ( .B(clk), .A(\g.we_clk [27990]));
Q_ASSIGN U4785 ( .B(clk), .A(\g.we_clk [27989]));
Q_ASSIGN U4786 ( .B(clk), .A(\g.we_clk [27988]));
Q_ASSIGN U4787 ( .B(clk), .A(\g.we_clk [27987]));
Q_ASSIGN U4788 ( .B(clk), .A(\g.we_clk [27986]));
Q_ASSIGN U4789 ( .B(clk), .A(\g.we_clk [27985]));
Q_ASSIGN U4790 ( .B(clk), .A(\g.we_clk [27984]));
Q_ASSIGN U4791 ( .B(clk), .A(\g.we_clk [27983]));
Q_ASSIGN U4792 ( .B(clk), .A(\g.we_clk [27982]));
Q_ASSIGN U4793 ( .B(clk), .A(\g.we_clk [27981]));
Q_ASSIGN U4794 ( .B(clk), .A(\g.we_clk [27980]));
Q_ASSIGN U4795 ( .B(clk), .A(\g.we_clk [27979]));
Q_ASSIGN U4796 ( .B(clk), .A(\g.we_clk [27978]));
Q_ASSIGN U4797 ( .B(clk), .A(\g.we_clk [27977]));
Q_ASSIGN U4798 ( .B(clk), .A(\g.we_clk [27976]));
Q_ASSIGN U4799 ( .B(clk), .A(\g.we_clk [27975]));
Q_ASSIGN U4800 ( .B(clk), .A(\g.we_clk [27974]));
Q_ASSIGN U4801 ( .B(clk), .A(\g.we_clk [27973]));
Q_ASSIGN U4802 ( .B(clk), .A(\g.we_clk [27972]));
Q_ASSIGN U4803 ( .B(clk), .A(\g.we_clk [27971]));
Q_ASSIGN U4804 ( .B(clk), .A(\g.we_clk [27970]));
Q_ASSIGN U4805 ( .B(clk), .A(\g.we_clk [27969]));
Q_ASSIGN U4806 ( .B(clk), .A(\g.we_clk [27968]));
Q_ASSIGN U4807 ( .B(clk), .A(\g.we_clk [27967]));
Q_ASSIGN U4808 ( .B(clk), .A(\g.we_clk [27966]));
Q_ASSIGN U4809 ( .B(clk), .A(\g.we_clk [27965]));
Q_ASSIGN U4810 ( .B(clk), .A(\g.we_clk [27964]));
Q_ASSIGN U4811 ( .B(clk), .A(\g.we_clk [27963]));
Q_ASSIGN U4812 ( .B(clk), .A(\g.we_clk [27962]));
Q_ASSIGN U4813 ( .B(clk), .A(\g.we_clk [27961]));
Q_ASSIGN U4814 ( .B(clk), .A(\g.we_clk [27960]));
Q_ASSIGN U4815 ( .B(clk), .A(\g.we_clk [27959]));
Q_ASSIGN U4816 ( .B(clk), .A(\g.we_clk [27958]));
Q_ASSIGN U4817 ( .B(clk), .A(\g.we_clk [27957]));
Q_ASSIGN U4818 ( .B(clk), .A(\g.we_clk [27956]));
Q_ASSIGN U4819 ( .B(clk), .A(\g.we_clk [27955]));
Q_ASSIGN U4820 ( .B(clk), .A(\g.we_clk [27954]));
Q_ASSIGN U4821 ( .B(clk), .A(\g.we_clk [27953]));
Q_ASSIGN U4822 ( .B(clk), .A(\g.we_clk [27952]));
Q_ASSIGN U4823 ( .B(clk), .A(\g.we_clk [27951]));
Q_ASSIGN U4824 ( .B(clk), .A(\g.we_clk [27950]));
Q_ASSIGN U4825 ( .B(clk), .A(\g.we_clk [27949]));
Q_ASSIGN U4826 ( .B(clk), .A(\g.we_clk [27948]));
Q_ASSIGN U4827 ( .B(clk), .A(\g.we_clk [27947]));
Q_ASSIGN U4828 ( .B(clk), .A(\g.we_clk [27946]));
Q_ASSIGN U4829 ( .B(clk), .A(\g.we_clk [27945]));
Q_ASSIGN U4830 ( .B(clk), .A(\g.we_clk [27944]));
Q_ASSIGN U4831 ( .B(clk), .A(\g.we_clk [27943]));
Q_ASSIGN U4832 ( .B(clk), .A(\g.we_clk [27942]));
Q_ASSIGN U4833 ( .B(clk), .A(\g.we_clk [27941]));
Q_ASSIGN U4834 ( .B(clk), .A(\g.we_clk [27940]));
Q_ASSIGN U4835 ( .B(clk), .A(\g.we_clk [27939]));
Q_ASSIGN U4836 ( .B(clk), .A(\g.we_clk [27938]));
Q_ASSIGN U4837 ( .B(clk), .A(\g.we_clk [27937]));
Q_ASSIGN U4838 ( .B(clk), .A(\g.we_clk [27936]));
Q_ASSIGN U4839 ( .B(clk), .A(\g.we_clk [27935]));
Q_ASSIGN U4840 ( .B(clk), .A(\g.we_clk [27934]));
Q_ASSIGN U4841 ( .B(clk), .A(\g.we_clk [27933]));
Q_ASSIGN U4842 ( .B(clk), .A(\g.we_clk [27932]));
Q_ASSIGN U4843 ( .B(clk), .A(\g.we_clk [27931]));
Q_ASSIGN U4844 ( .B(clk), .A(\g.we_clk [27930]));
Q_ASSIGN U4845 ( .B(clk), .A(\g.we_clk [27929]));
Q_ASSIGN U4846 ( .B(clk), .A(\g.we_clk [27928]));
Q_ASSIGN U4847 ( .B(clk), .A(\g.we_clk [27927]));
Q_ASSIGN U4848 ( .B(clk), .A(\g.we_clk [27926]));
Q_ASSIGN U4849 ( .B(clk), .A(\g.we_clk [27925]));
Q_ASSIGN U4850 ( .B(clk), .A(\g.we_clk [27924]));
Q_ASSIGN U4851 ( .B(clk), .A(\g.we_clk [27923]));
Q_ASSIGN U4852 ( .B(clk), .A(\g.we_clk [27922]));
Q_ASSIGN U4853 ( .B(clk), .A(\g.we_clk [27921]));
Q_ASSIGN U4854 ( .B(clk), .A(\g.we_clk [27920]));
Q_ASSIGN U4855 ( .B(clk), .A(\g.we_clk [27919]));
Q_ASSIGN U4856 ( .B(clk), .A(\g.we_clk [27918]));
Q_ASSIGN U4857 ( .B(clk), .A(\g.we_clk [27917]));
Q_ASSIGN U4858 ( .B(clk), .A(\g.we_clk [27916]));
Q_ASSIGN U4859 ( .B(clk), .A(\g.we_clk [27915]));
Q_ASSIGN U4860 ( .B(clk), .A(\g.we_clk [27914]));
Q_ASSIGN U4861 ( .B(clk), .A(\g.we_clk [27913]));
Q_ASSIGN U4862 ( .B(clk), .A(\g.we_clk [27912]));
Q_ASSIGN U4863 ( .B(clk), .A(\g.we_clk [27911]));
Q_ASSIGN U4864 ( .B(clk), .A(\g.we_clk [27910]));
Q_ASSIGN U4865 ( .B(clk), .A(\g.we_clk [27909]));
Q_ASSIGN U4866 ( .B(clk), .A(\g.we_clk [27908]));
Q_ASSIGN U4867 ( .B(clk), .A(\g.we_clk [27907]));
Q_ASSIGN U4868 ( .B(clk), .A(\g.we_clk [27906]));
Q_ASSIGN U4869 ( .B(clk), .A(\g.we_clk [27905]));
Q_ASSIGN U4870 ( .B(clk), .A(\g.we_clk [27904]));
Q_ASSIGN U4871 ( .B(clk), .A(\g.we_clk [27903]));
Q_ASSIGN U4872 ( .B(clk), .A(\g.we_clk [27902]));
Q_ASSIGN U4873 ( .B(clk), .A(\g.we_clk [27901]));
Q_ASSIGN U4874 ( .B(clk), .A(\g.we_clk [27900]));
Q_ASSIGN U4875 ( .B(clk), .A(\g.we_clk [27899]));
Q_ASSIGN U4876 ( .B(clk), .A(\g.we_clk [27898]));
Q_ASSIGN U4877 ( .B(clk), .A(\g.we_clk [27897]));
Q_ASSIGN U4878 ( .B(clk), .A(\g.we_clk [27896]));
Q_ASSIGN U4879 ( .B(clk), .A(\g.we_clk [27895]));
Q_ASSIGN U4880 ( .B(clk), .A(\g.we_clk [27894]));
Q_ASSIGN U4881 ( .B(clk), .A(\g.we_clk [27893]));
Q_ASSIGN U4882 ( .B(clk), .A(\g.we_clk [27892]));
Q_ASSIGN U4883 ( .B(clk), .A(\g.we_clk [27891]));
Q_ASSIGN U4884 ( .B(clk), .A(\g.we_clk [27890]));
Q_ASSIGN U4885 ( .B(clk), .A(\g.we_clk [27889]));
Q_ASSIGN U4886 ( .B(clk), .A(\g.we_clk [27888]));
Q_ASSIGN U4887 ( .B(clk), .A(\g.we_clk [27887]));
Q_ASSIGN U4888 ( .B(clk), .A(\g.we_clk [27886]));
Q_ASSIGN U4889 ( .B(clk), .A(\g.we_clk [27885]));
Q_ASSIGN U4890 ( .B(clk), .A(\g.we_clk [27884]));
Q_ASSIGN U4891 ( .B(clk), .A(\g.we_clk [27883]));
Q_ASSIGN U4892 ( .B(clk), .A(\g.we_clk [27882]));
Q_ASSIGN U4893 ( .B(clk), .A(\g.we_clk [27881]));
Q_ASSIGN U4894 ( .B(clk), .A(\g.we_clk [27880]));
Q_ASSIGN U4895 ( .B(clk), .A(\g.we_clk [27879]));
Q_ASSIGN U4896 ( .B(clk), .A(\g.we_clk [27878]));
Q_ASSIGN U4897 ( .B(clk), .A(\g.we_clk [27877]));
Q_ASSIGN U4898 ( .B(clk), .A(\g.we_clk [27876]));
Q_ASSIGN U4899 ( .B(clk), .A(\g.we_clk [27875]));
Q_ASSIGN U4900 ( .B(clk), .A(\g.we_clk [27874]));
Q_ASSIGN U4901 ( .B(clk), .A(\g.we_clk [27873]));
Q_ASSIGN U4902 ( .B(clk), .A(\g.we_clk [27872]));
Q_ASSIGN U4903 ( .B(clk), .A(\g.we_clk [27871]));
Q_ASSIGN U4904 ( .B(clk), .A(\g.we_clk [27870]));
Q_ASSIGN U4905 ( .B(clk), .A(\g.we_clk [27869]));
Q_ASSIGN U4906 ( .B(clk), .A(\g.we_clk [27868]));
Q_ASSIGN U4907 ( .B(clk), .A(\g.we_clk [27867]));
Q_ASSIGN U4908 ( .B(clk), .A(\g.we_clk [27866]));
Q_ASSIGN U4909 ( .B(clk), .A(\g.we_clk [27865]));
Q_ASSIGN U4910 ( .B(clk), .A(\g.we_clk [27864]));
Q_ASSIGN U4911 ( .B(clk), .A(\g.we_clk [27863]));
Q_ASSIGN U4912 ( .B(clk), .A(\g.we_clk [27862]));
Q_ASSIGN U4913 ( .B(clk), .A(\g.we_clk [27861]));
Q_ASSIGN U4914 ( .B(clk), .A(\g.we_clk [27860]));
Q_ASSIGN U4915 ( .B(clk), .A(\g.we_clk [27859]));
Q_ASSIGN U4916 ( .B(clk), .A(\g.we_clk [27858]));
Q_ASSIGN U4917 ( .B(clk), .A(\g.we_clk [27857]));
Q_ASSIGN U4918 ( .B(clk), .A(\g.we_clk [27856]));
Q_ASSIGN U4919 ( .B(clk), .A(\g.we_clk [27855]));
Q_ASSIGN U4920 ( .B(clk), .A(\g.we_clk [27854]));
Q_ASSIGN U4921 ( .B(clk), .A(\g.we_clk [27853]));
Q_ASSIGN U4922 ( .B(clk), .A(\g.we_clk [27852]));
Q_ASSIGN U4923 ( .B(clk), .A(\g.we_clk [27851]));
Q_ASSIGN U4924 ( .B(clk), .A(\g.we_clk [27850]));
Q_ASSIGN U4925 ( .B(clk), .A(\g.we_clk [27849]));
Q_ASSIGN U4926 ( .B(clk), .A(\g.we_clk [27848]));
Q_ASSIGN U4927 ( .B(clk), .A(\g.we_clk [27847]));
Q_ASSIGN U4928 ( .B(clk), .A(\g.we_clk [27846]));
Q_ASSIGN U4929 ( .B(clk), .A(\g.we_clk [27845]));
Q_ASSIGN U4930 ( .B(clk), .A(\g.we_clk [27844]));
Q_ASSIGN U4931 ( .B(clk), .A(\g.we_clk [27843]));
Q_ASSIGN U4932 ( .B(clk), .A(\g.we_clk [27842]));
Q_ASSIGN U4933 ( .B(clk), .A(\g.we_clk [27841]));
Q_ASSIGN U4934 ( .B(clk), .A(\g.we_clk [27840]));
Q_ASSIGN U4935 ( .B(clk), .A(\g.we_clk [27839]));
Q_ASSIGN U4936 ( .B(clk), .A(\g.we_clk [27838]));
Q_ASSIGN U4937 ( .B(clk), .A(\g.we_clk [27837]));
Q_ASSIGN U4938 ( .B(clk), .A(\g.we_clk [27836]));
Q_ASSIGN U4939 ( .B(clk), .A(\g.we_clk [27835]));
Q_ASSIGN U4940 ( .B(clk), .A(\g.we_clk [27834]));
Q_ASSIGN U4941 ( .B(clk), .A(\g.we_clk [27833]));
Q_ASSIGN U4942 ( .B(clk), .A(\g.we_clk [27832]));
Q_ASSIGN U4943 ( .B(clk), .A(\g.we_clk [27831]));
Q_ASSIGN U4944 ( .B(clk), .A(\g.we_clk [27830]));
Q_ASSIGN U4945 ( .B(clk), .A(\g.we_clk [27829]));
Q_ASSIGN U4946 ( .B(clk), .A(\g.we_clk [27828]));
Q_ASSIGN U4947 ( .B(clk), .A(\g.we_clk [27827]));
Q_ASSIGN U4948 ( .B(clk), .A(\g.we_clk [27826]));
Q_ASSIGN U4949 ( .B(clk), .A(\g.we_clk [27825]));
Q_ASSIGN U4950 ( .B(clk), .A(\g.we_clk [27824]));
Q_ASSIGN U4951 ( .B(clk), .A(\g.we_clk [27823]));
Q_ASSIGN U4952 ( .B(clk), .A(\g.we_clk [27822]));
Q_ASSIGN U4953 ( .B(clk), .A(\g.we_clk [27821]));
Q_ASSIGN U4954 ( .B(clk), .A(\g.we_clk [27820]));
Q_ASSIGN U4955 ( .B(clk), .A(\g.we_clk [27819]));
Q_ASSIGN U4956 ( .B(clk), .A(\g.we_clk [27818]));
Q_ASSIGN U4957 ( .B(clk), .A(\g.we_clk [27817]));
Q_ASSIGN U4958 ( .B(clk), .A(\g.we_clk [27816]));
Q_ASSIGN U4959 ( .B(clk), .A(\g.we_clk [27815]));
Q_ASSIGN U4960 ( .B(clk), .A(\g.we_clk [27814]));
Q_ASSIGN U4961 ( .B(clk), .A(\g.we_clk [27813]));
Q_ASSIGN U4962 ( .B(clk), .A(\g.we_clk [27812]));
Q_ASSIGN U4963 ( .B(clk), .A(\g.we_clk [27811]));
Q_ASSIGN U4964 ( .B(clk), .A(\g.we_clk [27810]));
Q_ASSIGN U4965 ( .B(clk), .A(\g.we_clk [27809]));
Q_ASSIGN U4966 ( .B(clk), .A(\g.we_clk [27808]));
Q_ASSIGN U4967 ( .B(clk), .A(\g.we_clk [27807]));
Q_ASSIGN U4968 ( .B(clk), .A(\g.we_clk [27806]));
Q_ASSIGN U4969 ( .B(clk), .A(\g.we_clk [27805]));
Q_ASSIGN U4970 ( .B(clk), .A(\g.we_clk [27804]));
Q_ASSIGN U4971 ( .B(clk), .A(\g.we_clk [27803]));
Q_ASSIGN U4972 ( .B(clk), .A(\g.we_clk [27802]));
Q_ASSIGN U4973 ( .B(clk), .A(\g.we_clk [27801]));
Q_ASSIGN U4974 ( .B(clk), .A(\g.we_clk [27800]));
Q_ASSIGN U4975 ( .B(clk), .A(\g.we_clk [27799]));
Q_ASSIGN U4976 ( .B(clk), .A(\g.we_clk [27798]));
Q_ASSIGN U4977 ( .B(clk), .A(\g.we_clk [27797]));
Q_ASSIGN U4978 ( .B(clk), .A(\g.we_clk [27796]));
Q_ASSIGN U4979 ( .B(clk), .A(\g.we_clk [27795]));
Q_ASSIGN U4980 ( .B(clk), .A(\g.we_clk [27794]));
Q_ASSIGN U4981 ( .B(clk), .A(\g.we_clk [27793]));
Q_ASSIGN U4982 ( .B(clk), .A(\g.we_clk [27792]));
Q_ASSIGN U4983 ( .B(clk), .A(\g.we_clk [27791]));
Q_ASSIGN U4984 ( .B(clk), .A(\g.we_clk [27790]));
Q_ASSIGN U4985 ( .B(clk), .A(\g.we_clk [27789]));
Q_ASSIGN U4986 ( .B(clk), .A(\g.we_clk [27788]));
Q_ASSIGN U4987 ( .B(clk), .A(\g.we_clk [27787]));
Q_ASSIGN U4988 ( .B(clk), .A(\g.we_clk [27786]));
Q_ASSIGN U4989 ( .B(clk), .A(\g.we_clk [27785]));
Q_ASSIGN U4990 ( .B(clk), .A(\g.we_clk [27784]));
Q_ASSIGN U4991 ( .B(clk), .A(\g.we_clk [27783]));
Q_ASSIGN U4992 ( .B(clk), .A(\g.we_clk [27782]));
Q_ASSIGN U4993 ( .B(clk), .A(\g.we_clk [27781]));
Q_ASSIGN U4994 ( .B(clk), .A(\g.we_clk [27780]));
Q_ASSIGN U4995 ( .B(clk), .A(\g.we_clk [27779]));
Q_ASSIGN U4996 ( .B(clk), .A(\g.we_clk [27778]));
Q_ASSIGN U4997 ( .B(clk), .A(\g.we_clk [27777]));
Q_ASSIGN U4998 ( .B(clk), .A(\g.we_clk [27776]));
Q_ASSIGN U4999 ( .B(clk), .A(\g.we_clk [27775]));
Q_ASSIGN U5000 ( .B(clk), .A(\g.we_clk [27774]));
Q_ASSIGN U5001 ( .B(clk), .A(\g.we_clk [27773]));
Q_ASSIGN U5002 ( .B(clk), .A(\g.we_clk [27772]));
Q_ASSIGN U5003 ( .B(clk), .A(\g.we_clk [27771]));
Q_ASSIGN U5004 ( .B(clk), .A(\g.we_clk [27770]));
Q_ASSIGN U5005 ( .B(clk), .A(\g.we_clk [27769]));
Q_ASSIGN U5006 ( .B(clk), .A(\g.we_clk [27768]));
Q_ASSIGN U5007 ( .B(clk), .A(\g.we_clk [27767]));
Q_ASSIGN U5008 ( .B(clk), .A(\g.we_clk [27766]));
Q_ASSIGN U5009 ( .B(clk), .A(\g.we_clk [27765]));
Q_ASSIGN U5010 ( .B(clk), .A(\g.we_clk [27764]));
Q_ASSIGN U5011 ( .B(clk), .A(\g.we_clk [27763]));
Q_ASSIGN U5012 ( .B(clk), .A(\g.we_clk [27762]));
Q_ASSIGN U5013 ( .B(clk), .A(\g.we_clk [27761]));
Q_ASSIGN U5014 ( .B(clk), .A(\g.we_clk [27760]));
Q_ASSIGN U5015 ( .B(clk), .A(\g.we_clk [27759]));
Q_ASSIGN U5016 ( .B(clk), .A(\g.we_clk [27758]));
Q_ASSIGN U5017 ( .B(clk), .A(\g.we_clk [27757]));
Q_ASSIGN U5018 ( .B(clk), .A(\g.we_clk [27756]));
Q_ASSIGN U5019 ( .B(clk), .A(\g.we_clk [27755]));
Q_ASSIGN U5020 ( .B(clk), .A(\g.we_clk [27754]));
Q_ASSIGN U5021 ( .B(clk), .A(\g.we_clk [27753]));
Q_ASSIGN U5022 ( .B(clk), .A(\g.we_clk [27752]));
Q_ASSIGN U5023 ( .B(clk), .A(\g.we_clk [27751]));
Q_ASSIGN U5024 ( .B(clk), .A(\g.we_clk [27750]));
Q_ASSIGN U5025 ( .B(clk), .A(\g.we_clk [27749]));
Q_ASSIGN U5026 ( .B(clk), .A(\g.we_clk [27748]));
Q_ASSIGN U5027 ( .B(clk), .A(\g.we_clk [27747]));
Q_ASSIGN U5028 ( .B(clk), .A(\g.we_clk [27746]));
Q_ASSIGN U5029 ( .B(clk), .A(\g.we_clk [27745]));
Q_ASSIGN U5030 ( .B(clk), .A(\g.we_clk [27744]));
Q_ASSIGN U5031 ( .B(clk), .A(\g.we_clk [27743]));
Q_ASSIGN U5032 ( .B(clk), .A(\g.we_clk [27742]));
Q_ASSIGN U5033 ( .B(clk), .A(\g.we_clk [27741]));
Q_ASSIGN U5034 ( .B(clk), .A(\g.we_clk [27740]));
Q_ASSIGN U5035 ( .B(clk), .A(\g.we_clk [27739]));
Q_ASSIGN U5036 ( .B(clk), .A(\g.we_clk [27738]));
Q_ASSIGN U5037 ( .B(clk), .A(\g.we_clk [27737]));
Q_ASSIGN U5038 ( .B(clk), .A(\g.we_clk [27736]));
Q_ASSIGN U5039 ( .B(clk), .A(\g.we_clk [27735]));
Q_ASSIGN U5040 ( .B(clk), .A(\g.we_clk [27734]));
Q_ASSIGN U5041 ( .B(clk), .A(\g.we_clk [27733]));
Q_ASSIGN U5042 ( .B(clk), .A(\g.we_clk [27732]));
Q_ASSIGN U5043 ( .B(clk), .A(\g.we_clk [27731]));
Q_ASSIGN U5044 ( .B(clk), .A(\g.we_clk [27730]));
Q_ASSIGN U5045 ( .B(clk), .A(\g.we_clk [27729]));
Q_ASSIGN U5046 ( .B(clk), .A(\g.we_clk [27728]));
Q_ASSIGN U5047 ( .B(clk), .A(\g.we_clk [27727]));
Q_ASSIGN U5048 ( .B(clk), .A(\g.we_clk [27726]));
Q_ASSIGN U5049 ( .B(clk), .A(\g.we_clk [27725]));
Q_ASSIGN U5050 ( .B(clk), .A(\g.we_clk [27724]));
Q_ASSIGN U5051 ( .B(clk), .A(\g.we_clk [27723]));
Q_ASSIGN U5052 ( .B(clk), .A(\g.we_clk [27722]));
Q_ASSIGN U5053 ( .B(clk), .A(\g.we_clk [27721]));
Q_ASSIGN U5054 ( .B(clk), .A(\g.we_clk [27720]));
Q_ASSIGN U5055 ( .B(clk), .A(\g.we_clk [27719]));
Q_ASSIGN U5056 ( .B(clk), .A(\g.we_clk [27718]));
Q_ASSIGN U5057 ( .B(clk), .A(\g.we_clk [27717]));
Q_ASSIGN U5058 ( .B(clk), .A(\g.we_clk [27716]));
Q_ASSIGN U5059 ( .B(clk), .A(\g.we_clk [27715]));
Q_ASSIGN U5060 ( .B(clk), .A(\g.we_clk [27714]));
Q_ASSIGN U5061 ( .B(clk), .A(\g.we_clk [27713]));
Q_ASSIGN U5062 ( .B(clk), .A(\g.we_clk [27712]));
Q_ASSIGN U5063 ( .B(clk), .A(\g.we_clk [27711]));
Q_ASSIGN U5064 ( .B(clk), .A(\g.we_clk [27710]));
Q_ASSIGN U5065 ( .B(clk), .A(\g.we_clk [27709]));
Q_ASSIGN U5066 ( .B(clk), .A(\g.we_clk [27708]));
Q_ASSIGN U5067 ( .B(clk), .A(\g.we_clk [27707]));
Q_ASSIGN U5068 ( .B(clk), .A(\g.we_clk [27706]));
Q_ASSIGN U5069 ( .B(clk), .A(\g.we_clk [27705]));
Q_ASSIGN U5070 ( .B(clk), .A(\g.we_clk [27704]));
Q_ASSIGN U5071 ( .B(clk), .A(\g.we_clk [27703]));
Q_ASSIGN U5072 ( .B(clk), .A(\g.we_clk [27702]));
Q_ASSIGN U5073 ( .B(clk), .A(\g.we_clk [27701]));
Q_ASSIGN U5074 ( .B(clk), .A(\g.we_clk [27700]));
Q_ASSIGN U5075 ( .B(clk), .A(\g.we_clk [27699]));
Q_ASSIGN U5076 ( .B(clk), .A(\g.we_clk [27698]));
Q_ASSIGN U5077 ( .B(clk), .A(\g.we_clk [27697]));
Q_ASSIGN U5078 ( .B(clk), .A(\g.we_clk [27696]));
Q_ASSIGN U5079 ( .B(clk), .A(\g.we_clk [27695]));
Q_ASSIGN U5080 ( .B(clk), .A(\g.we_clk [27694]));
Q_ASSIGN U5081 ( .B(clk), .A(\g.we_clk [27693]));
Q_ASSIGN U5082 ( .B(clk), .A(\g.we_clk [27692]));
Q_ASSIGN U5083 ( .B(clk), .A(\g.we_clk [27691]));
Q_ASSIGN U5084 ( .B(clk), .A(\g.we_clk [27690]));
Q_ASSIGN U5085 ( .B(clk), .A(\g.we_clk [27689]));
Q_ASSIGN U5086 ( .B(clk), .A(\g.we_clk [27688]));
Q_ASSIGN U5087 ( .B(clk), .A(\g.we_clk [27687]));
Q_ASSIGN U5088 ( .B(clk), .A(\g.we_clk [27686]));
Q_ASSIGN U5089 ( .B(clk), .A(\g.we_clk [27685]));
Q_ASSIGN U5090 ( .B(clk), .A(\g.we_clk [27684]));
Q_ASSIGN U5091 ( .B(clk), .A(\g.we_clk [27683]));
Q_ASSIGN U5092 ( .B(clk), .A(\g.we_clk [27682]));
Q_ASSIGN U5093 ( .B(clk), .A(\g.we_clk [27681]));
Q_ASSIGN U5094 ( .B(clk), .A(\g.we_clk [27680]));
Q_ASSIGN U5095 ( .B(clk), .A(\g.we_clk [27679]));
Q_ASSIGN U5096 ( .B(clk), .A(\g.we_clk [27678]));
Q_ASSIGN U5097 ( .B(clk), .A(\g.we_clk [27677]));
Q_ASSIGN U5098 ( .B(clk), .A(\g.we_clk [27676]));
Q_ASSIGN U5099 ( .B(clk), .A(\g.we_clk [27675]));
Q_ASSIGN U5100 ( .B(clk), .A(\g.we_clk [27674]));
Q_ASSIGN U5101 ( .B(clk), .A(\g.we_clk [27673]));
Q_ASSIGN U5102 ( .B(clk), .A(\g.we_clk [27672]));
Q_ASSIGN U5103 ( .B(clk), .A(\g.we_clk [27671]));
Q_ASSIGN U5104 ( .B(clk), .A(\g.we_clk [27670]));
Q_ASSIGN U5105 ( .B(clk), .A(\g.we_clk [27669]));
Q_ASSIGN U5106 ( .B(clk), .A(\g.we_clk [27668]));
Q_ASSIGN U5107 ( .B(clk), .A(\g.we_clk [27667]));
Q_ASSIGN U5108 ( .B(clk), .A(\g.we_clk [27666]));
Q_ASSIGN U5109 ( .B(clk), .A(\g.we_clk [27665]));
Q_ASSIGN U5110 ( .B(clk), .A(\g.we_clk [27664]));
Q_ASSIGN U5111 ( .B(clk), .A(\g.we_clk [27663]));
Q_ASSIGN U5112 ( .B(clk), .A(\g.we_clk [27662]));
Q_ASSIGN U5113 ( .B(clk), .A(\g.we_clk [27661]));
Q_ASSIGN U5114 ( .B(clk), .A(\g.we_clk [27660]));
Q_ASSIGN U5115 ( .B(clk), .A(\g.we_clk [27659]));
Q_ASSIGN U5116 ( .B(clk), .A(\g.we_clk [27658]));
Q_ASSIGN U5117 ( .B(clk), .A(\g.we_clk [27657]));
Q_ASSIGN U5118 ( .B(clk), .A(\g.we_clk [27656]));
Q_ASSIGN U5119 ( .B(clk), .A(\g.we_clk [27655]));
Q_ASSIGN U5120 ( .B(clk), .A(\g.we_clk [27654]));
Q_ASSIGN U5121 ( .B(clk), .A(\g.we_clk [27653]));
Q_ASSIGN U5122 ( .B(clk), .A(\g.we_clk [27652]));
Q_ASSIGN U5123 ( .B(clk), .A(\g.we_clk [27651]));
Q_ASSIGN U5124 ( .B(clk), .A(\g.we_clk [27650]));
Q_ASSIGN U5125 ( .B(clk), .A(\g.we_clk [27649]));
Q_ASSIGN U5126 ( .B(clk), .A(\g.we_clk [27648]));
Q_ASSIGN U5127 ( .B(clk), .A(\g.we_clk [27647]));
Q_ASSIGN U5128 ( .B(clk), .A(\g.we_clk [27646]));
Q_ASSIGN U5129 ( .B(clk), .A(\g.we_clk [27645]));
Q_ASSIGN U5130 ( .B(clk), .A(\g.we_clk [27644]));
Q_ASSIGN U5131 ( .B(clk), .A(\g.we_clk [27643]));
Q_ASSIGN U5132 ( .B(clk), .A(\g.we_clk [27642]));
Q_ASSIGN U5133 ( .B(clk), .A(\g.we_clk [27641]));
Q_ASSIGN U5134 ( .B(clk), .A(\g.we_clk [27640]));
Q_ASSIGN U5135 ( .B(clk), .A(\g.we_clk [27639]));
Q_ASSIGN U5136 ( .B(clk), .A(\g.we_clk [27638]));
Q_ASSIGN U5137 ( .B(clk), .A(\g.we_clk [27637]));
Q_ASSIGN U5138 ( .B(clk), .A(\g.we_clk [27636]));
Q_ASSIGN U5139 ( .B(clk), .A(\g.we_clk [27635]));
Q_ASSIGN U5140 ( .B(clk), .A(\g.we_clk [27634]));
Q_ASSIGN U5141 ( .B(clk), .A(\g.we_clk [27633]));
Q_ASSIGN U5142 ( .B(clk), .A(\g.we_clk [27632]));
Q_ASSIGN U5143 ( .B(clk), .A(\g.we_clk [27631]));
Q_ASSIGN U5144 ( .B(clk), .A(\g.we_clk [27630]));
Q_ASSIGN U5145 ( .B(clk), .A(\g.we_clk [27629]));
Q_ASSIGN U5146 ( .B(clk), .A(\g.we_clk [27628]));
Q_ASSIGN U5147 ( .B(clk), .A(\g.we_clk [27627]));
Q_ASSIGN U5148 ( .B(clk), .A(\g.we_clk [27626]));
Q_ASSIGN U5149 ( .B(clk), .A(\g.we_clk [27625]));
Q_ASSIGN U5150 ( .B(clk), .A(\g.we_clk [27624]));
Q_ASSIGN U5151 ( .B(clk), .A(\g.we_clk [27623]));
Q_ASSIGN U5152 ( .B(clk), .A(\g.we_clk [27622]));
Q_ASSIGN U5153 ( .B(clk), .A(\g.we_clk [27621]));
Q_ASSIGN U5154 ( .B(clk), .A(\g.we_clk [27620]));
Q_ASSIGN U5155 ( .B(clk), .A(\g.we_clk [27619]));
Q_ASSIGN U5156 ( .B(clk), .A(\g.we_clk [27618]));
Q_ASSIGN U5157 ( .B(clk), .A(\g.we_clk [27617]));
Q_ASSIGN U5158 ( .B(clk), .A(\g.we_clk [27616]));
Q_ASSIGN U5159 ( .B(clk), .A(\g.we_clk [27615]));
Q_ASSIGN U5160 ( .B(clk), .A(\g.we_clk [27614]));
Q_ASSIGN U5161 ( .B(clk), .A(\g.we_clk [27613]));
Q_ASSIGN U5162 ( .B(clk), .A(\g.we_clk [27612]));
Q_ASSIGN U5163 ( .B(clk), .A(\g.we_clk [27611]));
Q_ASSIGN U5164 ( .B(clk), .A(\g.we_clk [27610]));
Q_ASSIGN U5165 ( .B(clk), .A(\g.we_clk [27609]));
Q_ASSIGN U5166 ( .B(clk), .A(\g.we_clk [27608]));
Q_ASSIGN U5167 ( .B(clk), .A(\g.we_clk [27607]));
Q_ASSIGN U5168 ( .B(clk), .A(\g.we_clk [27606]));
Q_ASSIGN U5169 ( .B(clk), .A(\g.we_clk [27605]));
Q_ASSIGN U5170 ( .B(clk), .A(\g.we_clk [27604]));
Q_ASSIGN U5171 ( .B(clk), .A(\g.we_clk [27603]));
Q_ASSIGN U5172 ( .B(clk), .A(\g.we_clk [27602]));
Q_ASSIGN U5173 ( .B(clk), .A(\g.we_clk [27601]));
Q_ASSIGN U5174 ( .B(clk), .A(\g.we_clk [27600]));
Q_ASSIGN U5175 ( .B(clk), .A(\g.we_clk [27599]));
Q_ASSIGN U5176 ( .B(clk), .A(\g.we_clk [27598]));
Q_ASSIGN U5177 ( .B(clk), .A(\g.we_clk [27597]));
Q_ASSIGN U5178 ( .B(clk), .A(\g.we_clk [27596]));
Q_ASSIGN U5179 ( .B(clk), .A(\g.we_clk [27595]));
Q_ASSIGN U5180 ( .B(clk), .A(\g.we_clk [27594]));
Q_ASSIGN U5181 ( .B(clk), .A(\g.we_clk [27593]));
Q_ASSIGN U5182 ( .B(clk), .A(\g.we_clk [27592]));
Q_ASSIGN U5183 ( .B(clk), .A(\g.we_clk [27591]));
Q_ASSIGN U5184 ( .B(clk), .A(\g.we_clk [27590]));
Q_ASSIGN U5185 ( .B(clk), .A(\g.we_clk [27589]));
Q_ASSIGN U5186 ( .B(clk), .A(\g.we_clk [27588]));
Q_ASSIGN U5187 ( .B(clk), .A(\g.we_clk [27587]));
Q_ASSIGN U5188 ( .B(clk), .A(\g.we_clk [27586]));
Q_ASSIGN U5189 ( .B(clk), .A(\g.we_clk [27585]));
Q_ASSIGN U5190 ( .B(clk), .A(\g.we_clk [27584]));
Q_ASSIGN U5191 ( .B(clk), .A(\g.we_clk [27583]));
Q_ASSIGN U5192 ( .B(clk), .A(\g.we_clk [27582]));
Q_ASSIGN U5193 ( .B(clk), .A(\g.we_clk [27581]));
Q_ASSIGN U5194 ( .B(clk), .A(\g.we_clk [27580]));
Q_ASSIGN U5195 ( .B(clk), .A(\g.we_clk [27579]));
Q_ASSIGN U5196 ( .B(clk), .A(\g.we_clk [27578]));
Q_ASSIGN U5197 ( .B(clk), .A(\g.we_clk [27577]));
Q_ASSIGN U5198 ( .B(clk), .A(\g.we_clk [27576]));
Q_ASSIGN U5199 ( .B(clk), .A(\g.we_clk [27575]));
Q_ASSIGN U5200 ( .B(clk), .A(\g.we_clk [27574]));
Q_ASSIGN U5201 ( .B(clk), .A(\g.we_clk [27573]));
Q_ASSIGN U5202 ( .B(clk), .A(\g.we_clk [27572]));
Q_ASSIGN U5203 ( .B(clk), .A(\g.we_clk [27571]));
Q_ASSIGN U5204 ( .B(clk), .A(\g.we_clk [27570]));
Q_ASSIGN U5205 ( .B(clk), .A(\g.we_clk [27569]));
Q_ASSIGN U5206 ( .B(clk), .A(\g.we_clk [27568]));
Q_ASSIGN U5207 ( .B(clk), .A(\g.we_clk [27567]));
Q_ASSIGN U5208 ( .B(clk), .A(\g.we_clk [27566]));
Q_ASSIGN U5209 ( .B(clk), .A(\g.we_clk [27565]));
Q_ASSIGN U5210 ( .B(clk), .A(\g.we_clk [27564]));
Q_ASSIGN U5211 ( .B(clk), .A(\g.we_clk [27563]));
Q_ASSIGN U5212 ( .B(clk), .A(\g.we_clk [27562]));
Q_ASSIGN U5213 ( .B(clk), .A(\g.we_clk [27561]));
Q_ASSIGN U5214 ( .B(clk), .A(\g.we_clk [27560]));
Q_ASSIGN U5215 ( .B(clk), .A(\g.we_clk [27559]));
Q_ASSIGN U5216 ( .B(clk), .A(\g.we_clk [27558]));
Q_ASSIGN U5217 ( .B(clk), .A(\g.we_clk [27557]));
Q_ASSIGN U5218 ( .B(clk), .A(\g.we_clk [27556]));
Q_ASSIGN U5219 ( .B(clk), .A(\g.we_clk [27555]));
Q_ASSIGN U5220 ( .B(clk), .A(\g.we_clk [27554]));
Q_ASSIGN U5221 ( .B(clk), .A(\g.we_clk [27553]));
Q_ASSIGN U5222 ( .B(clk), .A(\g.we_clk [27552]));
Q_ASSIGN U5223 ( .B(clk), .A(\g.we_clk [27551]));
Q_ASSIGN U5224 ( .B(clk), .A(\g.we_clk [27550]));
Q_ASSIGN U5225 ( .B(clk), .A(\g.we_clk [27549]));
Q_ASSIGN U5226 ( .B(clk), .A(\g.we_clk [27548]));
Q_ASSIGN U5227 ( .B(clk), .A(\g.we_clk [27547]));
Q_ASSIGN U5228 ( .B(clk), .A(\g.we_clk [27546]));
Q_ASSIGN U5229 ( .B(clk), .A(\g.we_clk [27545]));
Q_ASSIGN U5230 ( .B(clk), .A(\g.we_clk [27544]));
Q_ASSIGN U5231 ( .B(clk), .A(\g.we_clk [27543]));
Q_ASSIGN U5232 ( .B(clk), .A(\g.we_clk [27542]));
Q_ASSIGN U5233 ( .B(clk), .A(\g.we_clk [27541]));
Q_ASSIGN U5234 ( .B(clk), .A(\g.we_clk [27540]));
Q_ASSIGN U5235 ( .B(clk), .A(\g.we_clk [27539]));
Q_ASSIGN U5236 ( .B(clk), .A(\g.we_clk [27538]));
Q_ASSIGN U5237 ( .B(clk), .A(\g.we_clk [27537]));
Q_ASSIGN U5238 ( .B(clk), .A(\g.we_clk [27536]));
Q_ASSIGN U5239 ( .B(clk), .A(\g.we_clk [27535]));
Q_ASSIGN U5240 ( .B(clk), .A(\g.we_clk [27534]));
Q_ASSIGN U5241 ( .B(clk), .A(\g.we_clk [27533]));
Q_ASSIGN U5242 ( .B(clk), .A(\g.we_clk [27532]));
Q_ASSIGN U5243 ( .B(clk), .A(\g.we_clk [27531]));
Q_ASSIGN U5244 ( .B(clk), .A(\g.we_clk [27530]));
Q_ASSIGN U5245 ( .B(clk), .A(\g.we_clk [27529]));
Q_ASSIGN U5246 ( .B(clk), .A(\g.we_clk [27528]));
Q_ASSIGN U5247 ( .B(clk), .A(\g.we_clk [27527]));
Q_ASSIGN U5248 ( .B(clk), .A(\g.we_clk [27526]));
Q_ASSIGN U5249 ( .B(clk), .A(\g.we_clk [27525]));
Q_ASSIGN U5250 ( .B(clk), .A(\g.we_clk [27524]));
Q_ASSIGN U5251 ( .B(clk), .A(\g.we_clk [27523]));
Q_ASSIGN U5252 ( .B(clk), .A(\g.we_clk [27522]));
Q_ASSIGN U5253 ( .B(clk), .A(\g.we_clk [27521]));
Q_ASSIGN U5254 ( .B(clk), .A(\g.we_clk [27520]));
Q_ASSIGN U5255 ( .B(clk), .A(\g.we_clk [27519]));
Q_ASSIGN U5256 ( .B(clk), .A(\g.we_clk [27518]));
Q_ASSIGN U5257 ( .B(clk), .A(\g.we_clk [27517]));
Q_ASSIGN U5258 ( .B(clk), .A(\g.we_clk [27516]));
Q_ASSIGN U5259 ( .B(clk), .A(\g.we_clk [27515]));
Q_ASSIGN U5260 ( .B(clk), .A(\g.we_clk [27514]));
Q_ASSIGN U5261 ( .B(clk), .A(\g.we_clk [27513]));
Q_ASSIGN U5262 ( .B(clk), .A(\g.we_clk [27512]));
Q_ASSIGN U5263 ( .B(clk), .A(\g.we_clk [27511]));
Q_ASSIGN U5264 ( .B(clk), .A(\g.we_clk [27510]));
Q_ASSIGN U5265 ( .B(clk), .A(\g.we_clk [27509]));
Q_ASSIGN U5266 ( .B(clk), .A(\g.we_clk [27508]));
Q_ASSIGN U5267 ( .B(clk), .A(\g.we_clk [27507]));
Q_ASSIGN U5268 ( .B(clk), .A(\g.we_clk [27506]));
Q_ASSIGN U5269 ( .B(clk), .A(\g.we_clk [27505]));
Q_ASSIGN U5270 ( .B(clk), .A(\g.we_clk [27504]));
Q_ASSIGN U5271 ( .B(clk), .A(\g.we_clk [27503]));
Q_ASSIGN U5272 ( .B(clk), .A(\g.we_clk [27502]));
Q_ASSIGN U5273 ( .B(clk), .A(\g.we_clk [27501]));
Q_ASSIGN U5274 ( .B(clk), .A(\g.we_clk [27500]));
Q_ASSIGN U5275 ( .B(clk), .A(\g.we_clk [27499]));
Q_ASSIGN U5276 ( .B(clk), .A(\g.we_clk [27498]));
Q_ASSIGN U5277 ( .B(clk), .A(\g.we_clk [27497]));
Q_ASSIGN U5278 ( .B(clk), .A(\g.we_clk [27496]));
Q_ASSIGN U5279 ( .B(clk), .A(\g.we_clk [27495]));
Q_ASSIGN U5280 ( .B(clk), .A(\g.we_clk [27494]));
Q_ASSIGN U5281 ( .B(clk), .A(\g.we_clk [27493]));
Q_ASSIGN U5282 ( .B(clk), .A(\g.we_clk [27492]));
Q_ASSIGN U5283 ( .B(clk), .A(\g.we_clk [27491]));
Q_ASSIGN U5284 ( .B(clk), .A(\g.we_clk [27490]));
Q_ASSIGN U5285 ( .B(clk), .A(\g.we_clk [27489]));
Q_ASSIGN U5286 ( .B(clk), .A(\g.we_clk [27488]));
Q_ASSIGN U5287 ( .B(clk), .A(\g.we_clk [27487]));
Q_ASSIGN U5288 ( .B(clk), .A(\g.we_clk [27486]));
Q_ASSIGN U5289 ( .B(clk), .A(\g.we_clk [27485]));
Q_ASSIGN U5290 ( .B(clk), .A(\g.we_clk [27484]));
Q_ASSIGN U5291 ( .B(clk), .A(\g.we_clk [27483]));
Q_ASSIGN U5292 ( .B(clk), .A(\g.we_clk [27482]));
Q_ASSIGN U5293 ( .B(clk), .A(\g.we_clk [27481]));
Q_ASSIGN U5294 ( .B(clk), .A(\g.we_clk [27480]));
Q_ASSIGN U5295 ( .B(clk), .A(\g.we_clk [27479]));
Q_ASSIGN U5296 ( .B(clk), .A(\g.we_clk [27478]));
Q_ASSIGN U5297 ( .B(clk), .A(\g.we_clk [27477]));
Q_ASSIGN U5298 ( .B(clk), .A(\g.we_clk [27476]));
Q_ASSIGN U5299 ( .B(clk), .A(\g.we_clk [27475]));
Q_ASSIGN U5300 ( .B(clk), .A(\g.we_clk [27474]));
Q_ASSIGN U5301 ( .B(clk), .A(\g.we_clk [27473]));
Q_ASSIGN U5302 ( .B(clk), .A(\g.we_clk [27472]));
Q_ASSIGN U5303 ( .B(clk), .A(\g.we_clk [27471]));
Q_ASSIGN U5304 ( .B(clk), .A(\g.we_clk [27470]));
Q_ASSIGN U5305 ( .B(clk), .A(\g.we_clk [27469]));
Q_ASSIGN U5306 ( .B(clk), .A(\g.we_clk [27468]));
Q_ASSIGN U5307 ( .B(clk), .A(\g.we_clk [27467]));
Q_ASSIGN U5308 ( .B(clk), .A(\g.we_clk [27466]));
Q_ASSIGN U5309 ( .B(clk), .A(\g.we_clk [27465]));
Q_ASSIGN U5310 ( .B(clk), .A(\g.we_clk [27464]));
Q_ASSIGN U5311 ( .B(clk), .A(\g.we_clk [27463]));
Q_ASSIGN U5312 ( .B(clk), .A(\g.we_clk [27462]));
Q_ASSIGN U5313 ( .B(clk), .A(\g.we_clk [27461]));
Q_ASSIGN U5314 ( .B(clk), .A(\g.we_clk [27460]));
Q_ASSIGN U5315 ( .B(clk), .A(\g.we_clk [27459]));
Q_ASSIGN U5316 ( .B(clk), .A(\g.we_clk [27458]));
Q_ASSIGN U5317 ( .B(clk), .A(\g.we_clk [27457]));
Q_ASSIGN U5318 ( .B(clk), .A(\g.we_clk [27456]));
Q_ASSIGN U5319 ( .B(clk), .A(\g.we_clk [27455]));
Q_ASSIGN U5320 ( .B(clk), .A(\g.we_clk [27454]));
Q_ASSIGN U5321 ( .B(clk), .A(\g.we_clk [27453]));
Q_ASSIGN U5322 ( .B(clk), .A(\g.we_clk [27452]));
Q_ASSIGN U5323 ( .B(clk), .A(\g.we_clk [27451]));
Q_ASSIGN U5324 ( .B(clk), .A(\g.we_clk [27450]));
Q_ASSIGN U5325 ( .B(clk), .A(\g.we_clk [27449]));
Q_ASSIGN U5326 ( .B(clk), .A(\g.we_clk [27448]));
Q_ASSIGN U5327 ( .B(clk), .A(\g.we_clk [27447]));
Q_ASSIGN U5328 ( .B(clk), .A(\g.we_clk [27446]));
Q_ASSIGN U5329 ( .B(clk), .A(\g.we_clk [27445]));
Q_ASSIGN U5330 ( .B(clk), .A(\g.we_clk [27444]));
Q_ASSIGN U5331 ( .B(clk), .A(\g.we_clk [27443]));
Q_ASSIGN U5332 ( .B(clk), .A(\g.we_clk [27442]));
Q_ASSIGN U5333 ( .B(clk), .A(\g.we_clk [27441]));
Q_ASSIGN U5334 ( .B(clk), .A(\g.we_clk [27440]));
Q_ASSIGN U5335 ( .B(clk), .A(\g.we_clk [27439]));
Q_ASSIGN U5336 ( .B(clk), .A(\g.we_clk [27438]));
Q_ASSIGN U5337 ( .B(clk), .A(\g.we_clk [27437]));
Q_ASSIGN U5338 ( .B(clk), .A(\g.we_clk [27436]));
Q_ASSIGN U5339 ( .B(clk), .A(\g.we_clk [27435]));
Q_ASSIGN U5340 ( .B(clk), .A(\g.we_clk [27434]));
Q_ASSIGN U5341 ( .B(clk), .A(\g.we_clk [27433]));
Q_ASSIGN U5342 ( .B(clk), .A(\g.we_clk [27432]));
Q_ASSIGN U5343 ( .B(clk), .A(\g.we_clk [27431]));
Q_ASSIGN U5344 ( .B(clk), .A(\g.we_clk [27430]));
Q_ASSIGN U5345 ( .B(clk), .A(\g.we_clk [27429]));
Q_ASSIGN U5346 ( .B(clk), .A(\g.we_clk [27428]));
Q_ASSIGN U5347 ( .B(clk), .A(\g.we_clk [27427]));
Q_ASSIGN U5348 ( .B(clk), .A(\g.we_clk [27426]));
Q_ASSIGN U5349 ( .B(clk), .A(\g.we_clk [27425]));
Q_ASSIGN U5350 ( .B(clk), .A(\g.we_clk [27424]));
Q_ASSIGN U5351 ( .B(clk), .A(\g.we_clk [27423]));
Q_ASSIGN U5352 ( .B(clk), .A(\g.we_clk [27422]));
Q_ASSIGN U5353 ( .B(clk), .A(\g.we_clk [27421]));
Q_ASSIGN U5354 ( .B(clk), .A(\g.we_clk [27420]));
Q_ASSIGN U5355 ( .B(clk), .A(\g.we_clk [27419]));
Q_ASSIGN U5356 ( .B(clk), .A(\g.we_clk [27418]));
Q_ASSIGN U5357 ( .B(clk), .A(\g.we_clk [27417]));
Q_ASSIGN U5358 ( .B(clk), .A(\g.we_clk [27416]));
Q_ASSIGN U5359 ( .B(clk), .A(\g.we_clk [27415]));
Q_ASSIGN U5360 ( .B(clk), .A(\g.we_clk [27414]));
Q_ASSIGN U5361 ( .B(clk), .A(\g.we_clk [27413]));
Q_ASSIGN U5362 ( .B(clk), .A(\g.we_clk [27412]));
Q_ASSIGN U5363 ( .B(clk), .A(\g.we_clk [27411]));
Q_ASSIGN U5364 ( .B(clk), .A(\g.we_clk [27410]));
Q_ASSIGN U5365 ( .B(clk), .A(\g.we_clk [27409]));
Q_ASSIGN U5366 ( .B(clk), .A(\g.we_clk [27408]));
Q_ASSIGN U5367 ( .B(clk), .A(\g.we_clk [27407]));
Q_ASSIGN U5368 ( .B(clk), .A(\g.we_clk [27406]));
Q_ASSIGN U5369 ( .B(clk), .A(\g.we_clk [27405]));
Q_ASSIGN U5370 ( .B(clk), .A(\g.we_clk [27404]));
Q_ASSIGN U5371 ( .B(clk), .A(\g.we_clk [27403]));
Q_ASSIGN U5372 ( .B(clk), .A(\g.we_clk [27402]));
Q_ASSIGN U5373 ( .B(clk), .A(\g.we_clk [27401]));
Q_ASSIGN U5374 ( .B(clk), .A(\g.we_clk [27400]));
Q_ASSIGN U5375 ( .B(clk), .A(\g.we_clk [27399]));
Q_ASSIGN U5376 ( .B(clk), .A(\g.we_clk [27398]));
Q_ASSIGN U5377 ( .B(clk), .A(\g.we_clk [27397]));
Q_ASSIGN U5378 ( .B(clk), .A(\g.we_clk [27396]));
Q_ASSIGN U5379 ( .B(clk), .A(\g.we_clk [27395]));
Q_ASSIGN U5380 ( .B(clk), .A(\g.we_clk [27394]));
Q_ASSIGN U5381 ( .B(clk), .A(\g.we_clk [27393]));
Q_ASSIGN U5382 ( .B(clk), .A(\g.we_clk [27392]));
Q_ASSIGN U5383 ( .B(clk), .A(\g.we_clk [27391]));
Q_ASSIGN U5384 ( .B(clk), .A(\g.we_clk [27390]));
Q_ASSIGN U5385 ( .B(clk), .A(\g.we_clk [27389]));
Q_ASSIGN U5386 ( .B(clk), .A(\g.we_clk [27388]));
Q_ASSIGN U5387 ( .B(clk), .A(\g.we_clk [27387]));
Q_ASSIGN U5388 ( .B(clk), .A(\g.we_clk [27386]));
Q_ASSIGN U5389 ( .B(clk), .A(\g.we_clk [27385]));
Q_ASSIGN U5390 ( .B(clk), .A(\g.we_clk [27384]));
Q_ASSIGN U5391 ( .B(clk), .A(\g.we_clk [27383]));
Q_ASSIGN U5392 ( .B(clk), .A(\g.we_clk [27382]));
Q_ASSIGN U5393 ( .B(clk), .A(\g.we_clk [27381]));
Q_ASSIGN U5394 ( .B(clk), .A(\g.we_clk [27380]));
Q_ASSIGN U5395 ( .B(clk), .A(\g.we_clk [27379]));
Q_ASSIGN U5396 ( .B(clk), .A(\g.we_clk [27378]));
Q_ASSIGN U5397 ( .B(clk), .A(\g.we_clk [27377]));
Q_ASSIGN U5398 ( .B(clk), .A(\g.we_clk [27376]));
Q_ASSIGN U5399 ( .B(clk), .A(\g.we_clk [27375]));
Q_ASSIGN U5400 ( .B(clk), .A(\g.we_clk [27374]));
Q_ASSIGN U5401 ( .B(clk), .A(\g.we_clk [27373]));
Q_ASSIGN U5402 ( .B(clk), .A(\g.we_clk [27372]));
Q_ASSIGN U5403 ( .B(clk), .A(\g.we_clk [27371]));
Q_ASSIGN U5404 ( .B(clk), .A(\g.we_clk [27370]));
Q_ASSIGN U5405 ( .B(clk), .A(\g.we_clk [27369]));
Q_ASSIGN U5406 ( .B(clk), .A(\g.we_clk [27368]));
Q_ASSIGN U5407 ( .B(clk), .A(\g.we_clk [27367]));
Q_ASSIGN U5408 ( .B(clk), .A(\g.we_clk [27366]));
Q_ASSIGN U5409 ( .B(clk), .A(\g.we_clk [27365]));
Q_ASSIGN U5410 ( .B(clk), .A(\g.we_clk [27364]));
Q_ASSIGN U5411 ( .B(clk), .A(\g.we_clk [27363]));
Q_ASSIGN U5412 ( .B(clk), .A(\g.we_clk [27362]));
Q_ASSIGN U5413 ( .B(clk), .A(\g.we_clk [27361]));
Q_ASSIGN U5414 ( .B(clk), .A(\g.we_clk [27360]));
Q_ASSIGN U5415 ( .B(clk), .A(\g.we_clk [27359]));
Q_ASSIGN U5416 ( .B(clk), .A(\g.we_clk [27358]));
Q_ASSIGN U5417 ( .B(clk), .A(\g.we_clk [27357]));
Q_ASSIGN U5418 ( .B(clk), .A(\g.we_clk [27356]));
Q_ASSIGN U5419 ( .B(clk), .A(\g.we_clk [27355]));
Q_ASSIGN U5420 ( .B(clk), .A(\g.we_clk [27354]));
Q_ASSIGN U5421 ( .B(clk), .A(\g.we_clk [27353]));
Q_ASSIGN U5422 ( .B(clk), .A(\g.we_clk [27352]));
Q_ASSIGN U5423 ( .B(clk), .A(\g.we_clk [27351]));
Q_ASSIGN U5424 ( .B(clk), .A(\g.we_clk [27350]));
Q_ASSIGN U5425 ( .B(clk), .A(\g.we_clk [27349]));
Q_ASSIGN U5426 ( .B(clk), .A(\g.we_clk [27348]));
Q_ASSIGN U5427 ( .B(clk), .A(\g.we_clk [27347]));
Q_ASSIGN U5428 ( .B(clk), .A(\g.we_clk [27346]));
Q_ASSIGN U5429 ( .B(clk), .A(\g.we_clk [27345]));
Q_ASSIGN U5430 ( .B(clk), .A(\g.we_clk [27344]));
Q_ASSIGN U5431 ( .B(clk), .A(\g.we_clk [27343]));
Q_ASSIGN U5432 ( .B(clk), .A(\g.we_clk [27342]));
Q_ASSIGN U5433 ( .B(clk), .A(\g.we_clk [27341]));
Q_ASSIGN U5434 ( .B(clk), .A(\g.we_clk [27340]));
Q_ASSIGN U5435 ( .B(clk), .A(\g.we_clk [27339]));
Q_ASSIGN U5436 ( .B(clk), .A(\g.we_clk [27338]));
Q_ASSIGN U5437 ( .B(clk), .A(\g.we_clk [27337]));
Q_ASSIGN U5438 ( .B(clk), .A(\g.we_clk [27336]));
Q_ASSIGN U5439 ( .B(clk), .A(\g.we_clk [27335]));
Q_ASSIGN U5440 ( .B(clk), .A(\g.we_clk [27334]));
Q_ASSIGN U5441 ( .B(clk), .A(\g.we_clk [27333]));
Q_ASSIGN U5442 ( .B(clk), .A(\g.we_clk [27332]));
Q_ASSIGN U5443 ( .B(clk), .A(\g.we_clk [27331]));
Q_ASSIGN U5444 ( .B(clk), .A(\g.we_clk [27330]));
Q_ASSIGN U5445 ( .B(clk), .A(\g.we_clk [27329]));
Q_ASSIGN U5446 ( .B(clk), .A(\g.we_clk [27328]));
Q_ASSIGN U5447 ( .B(clk), .A(\g.we_clk [27327]));
Q_ASSIGN U5448 ( .B(clk), .A(\g.we_clk [27326]));
Q_ASSIGN U5449 ( .B(clk), .A(\g.we_clk [27325]));
Q_ASSIGN U5450 ( .B(clk), .A(\g.we_clk [27324]));
Q_ASSIGN U5451 ( .B(clk), .A(\g.we_clk [27323]));
Q_ASSIGN U5452 ( .B(clk), .A(\g.we_clk [27322]));
Q_ASSIGN U5453 ( .B(clk), .A(\g.we_clk [27321]));
Q_ASSIGN U5454 ( .B(clk), .A(\g.we_clk [27320]));
Q_ASSIGN U5455 ( .B(clk), .A(\g.we_clk [27319]));
Q_ASSIGN U5456 ( .B(clk), .A(\g.we_clk [27318]));
Q_ASSIGN U5457 ( .B(clk), .A(\g.we_clk [27317]));
Q_ASSIGN U5458 ( .B(clk), .A(\g.we_clk [27316]));
Q_ASSIGN U5459 ( .B(clk), .A(\g.we_clk [27315]));
Q_ASSIGN U5460 ( .B(clk), .A(\g.we_clk [27314]));
Q_ASSIGN U5461 ( .B(clk), .A(\g.we_clk [27313]));
Q_ASSIGN U5462 ( .B(clk), .A(\g.we_clk [27312]));
Q_ASSIGN U5463 ( .B(clk), .A(\g.we_clk [27311]));
Q_ASSIGN U5464 ( .B(clk), .A(\g.we_clk [27310]));
Q_ASSIGN U5465 ( .B(clk), .A(\g.we_clk [27309]));
Q_ASSIGN U5466 ( .B(clk), .A(\g.we_clk [27308]));
Q_ASSIGN U5467 ( .B(clk), .A(\g.we_clk [27307]));
Q_ASSIGN U5468 ( .B(clk), .A(\g.we_clk [27306]));
Q_ASSIGN U5469 ( .B(clk), .A(\g.we_clk [27305]));
Q_ASSIGN U5470 ( .B(clk), .A(\g.we_clk [27304]));
Q_ASSIGN U5471 ( .B(clk), .A(\g.we_clk [27303]));
Q_ASSIGN U5472 ( .B(clk), .A(\g.we_clk [27302]));
Q_ASSIGN U5473 ( .B(clk), .A(\g.we_clk [27301]));
Q_ASSIGN U5474 ( .B(clk), .A(\g.we_clk [27300]));
Q_ASSIGN U5475 ( .B(clk), .A(\g.we_clk [27299]));
Q_ASSIGN U5476 ( .B(clk), .A(\g.we_clk [27298]));
Q_ASSIGN U5477 ( .B(clk), .A(\g.we_clk [27297]));
Q_ASSIGN U5478 ( .B(clk), .A(\g.we_clk [27296]));
Q_ASSIGN U5479 ( .B(clk), .A(\g.we_clk [27295]));
Q_ASSIGN U5480 ( .B(clk), .A(\g.we_clk [27294]));
Q_ASSIGN U5481 ( .B(clk), .A(\g.we_clk [27293]));
Q_ASSIGN U5482 ( .B(clk), .A(\g.we_clk [27292]));
Q_ASSIGN U5483 ( .B(clk), .A(\g.we_clk [27291]));
Q_ASSIGN U5484 ( .B(clk), .A(\g.we_clk [27290]));
Q_ASSIGN U5485 ( .B(clk), .A(\g.we_clk [27289]));
Q_ASSIGN U5486 ( .B(clk), .A(\g.we_clk [27288]));
Q_ASSIGN U5487 ( .B(clk), .A(\g.we_clk [27287]));
Q_ASSIGN U5488 ( .B(clk), .A(\g.we_clk [27286]));
Q_ASSIGN U5489 ( .B(clk), .A(\g.we_clk [27285]));
Q_ASSIGN U5490 ( .B(clk), .A(\g.we_clk [27284]));
Q_ASSIGN U5491 ( .B(clk), .A(\g.we_clk [27283]));
Q_ASSIGN U5492 ( .B(clk), .A(\g.we_clk [27282]));
Q_ASSIGN U5493 ( .B(clk), .A(\g.we_clk [27281]));
Q_ASSIGN U5494 ( .B(clk), .A(\g.we_clk [27280]));
Q_ASSIGN U5495 ( .B(clk), .A(\g.we_clk [27279]));
Q_ASSIGN U5496 ( .B(clk), .A(\g.we_clk [27278]));
Q_ASSIGN U5497 ( .B(clk), .A(\g.we_clk [27277]));
Q_ASSIGN U5498 ( .B(clk), .A(\g.we_clk [27276]));
Q_ASSIGN U5499 ( .B(clk), .A(\g.we_clk [27275]));
Q_ASSIGN U5500 ( .B(clk), .A(\g.we_clk [27274]));
Q_ASSIGN U5501 ( .B(clk), .A(\g.we_clk [27273]));
Q_ASSIGN U5502 ( .B(clk), .A(\g.we_clk [27272]));
Q_ASSIGN U5503 ( .B(clk), .A(\g.we_clk [27271]));
Q_ASSIGN U5504 ( .B(clk), .A(\g.we_clk [27270]));
Q_ASSIGN U5505 ( .B(clk), .A(\g.we_clk [27269]));
Q_ASSIGN U5506 ( .B(clk), .A(\g.we_clk [27268]));
Q_ASSIGN U5507 ( .B(clk), .A(\g.we_clk [27267]));
Q_ASSIGN U5508 ( .B(clk), .A(\g.we_clk [27266]));
Q_ASSIGN U5509 ( .B(clk), .A(\g.we_clk [27265]));
Q_ASSIGN U5510 ( .B(clk), .A(\g.we_clk [27264]));
Q_ASSIGN U5511 ( .B(clk), .A(\g.we_clk [27263]));
Q_ASSIGN U5512 ( .B(clk), .A(\g.we_clk [27262]));
Q_ASSIGN U5513 ( .B(clk), .A(\g.we_clk [27261]));
Q_ASSIGN U5514 ( .B(clk), .A(\g.we_clk [27260]));
Q_ASSIGN U5515 ( .B(clk), .A(\g.we_clk [27259]));
Q_ASSIGN U5516 ( .B(clk), .A(\g.we_clk [27258]));
Q_ASSIGN U5517 ( .B(clk), .A(\g.we_clk [27257]));
Q_ASSIGN U5518 ( .B(clk), .A(\g.we_clk [27256]));
Q_ASSIGN U5519 ( .B(clk), .A(\g.we_clk [27255]));
Q_ASSIGN U5520 ( .B(clk), .A(\g.we_clk [27254]));
Q_ASSIGN U5521 ( .B(clk), .A(\g.we_clk [27253]));
Q_ASSIGN U5522 ( .B(clk), .A(\g.we_clk [27252]));
Q_ASSIGN U5523 ( .B(clk), .A(\g.we_clk [27251]));
Q_ASSIGN U5524 ( .B(clk), .A(\g.we_clk [27250]));
Q_ASSIGN U5525 ( .B(clk), .A(\g.we_clk [27249]));
Q_ASSIGN U5526 ( .B(clk), .A(\g.we_clk [27248]));
Q_ASSIGN U5527 ( .B(clk), .A(\g.we_clk [27247]));
Q_ASSIGN U5528 ( .B(clk), .A(\g.we_clk [27246]));
Q_ASSIGN U5529 ( .B(clk), .A(\g.we_clk [27245]));
Q_ASSIGN U5530 ( .B(clk), .A(\g.we_clk [27244]));
Q_ASSIGN U5531 ( .B(clk), .A(\g.we_clk [27243]));
Q_ASSIGN U5532 ( .B(clk), .A(\g.we_clk [27242]));
Q_ASSIGN U5533 ( .B(clk), .A(\g.we_clk [27241]));
Q_ASSIGN U5534 ( .B(clk), .A(\g.we_clk [27240]));
Q_ASSIGN U5535 ( .B(clk), .A(\g.we_clk [27239]));
Q_ASSIGN U5536 ( .B(clk), .A(\g.we_clk [27238]));
Q_ASSIGN U5537 ( .B(clk), .A(\g.we_clk [27237]));
Q_ASSIGN U5538 ( .B(clk), .A(\g.we_clk [27236]));
Q_ASSIGN U5539 ( .B(clk), .A(\g.we_clk [27235]));
Q_ASSIGN U5540 ( .B(clk), .A(\g.we_clk [27234]));
Q_ASSIGN U5541 ( .B(clk), .A(\g.we_clk [27233]));
Q_ASSIGN U5542 ( .B(clk), .A(\g.we_clk [27232]));
Q_ASSIGN U5543 ( .B(clk), .A(\g.we_clk [27231]));
Q_ASSIGN U5544 ( .B(clk), .A(\g.we_clk [27230]));
Q_ASSIGN U5545 ( .B(clk), .A(\g.we_clk [27229]));
Q_ASSIGN U5546 ( .B(clk), .A(\g.we_clk [27228]));
Q_ASSIGN U5547 ( .B(clk), .A(\g.we_clk [27227]));
Q_ASSIGN U5548 ( .B(clk), .A(\g.we_clk [27226]));
Q_ASSIGN U5549 ( .B(clk), .A(\g.we_clk [27225]));
Q_ASSIGN U5550 ( .B(clk), .A(\g.we_clk [27224]));
Q_ASSIGN U5551 ( .B(clk), .A(\g.we_clk [27223]));
Q_ASSIGN U5552 ( .B(clk), .A(\g.we_clk [27222]));
Q_ASSIGN U5553 ( .B(clk), .A(\g.we_clk [27221]));
Q_ASSIGN U5554 ( .B(clk), .A(\g.we_clk [27220]));
Q_ASSIGN U5555 ( .B(clk), .A(\g.we_clk [27219]));
Q_ASSIGN U5556 ( .B(clk), .A(\g.we_clk [27218]));
Q_ASSIGN U5557 ( .B(clk), .A(\g.we_clk [27217]));
Q_ASSIGN U5558 ( .B(clk), .A(\g.we_clk [27216]));
Q_ASSIGN U5559 ( .B(clk), .A(\g.we_clk [27215]));
Q_ASSIGN U5560 ( .B(clk), .A(\g.we_clk [27214]));
Q_ASSIGN U5561 ( .B(clk), .A(\g.we_clk [27213]));
Q_ASSIGN U5562 ( .B(clk), .A(\g.we_clk [27212]));
Q_ASSIGN U5563 ( .B(clk), .A(\g.we_clk [27211]));
Q_ASSIGN U5564 ( .B(clk), .A(\g.we_clk [27210]));
Q_ASSIGN U5565 ( .B(clk), .A(\g.we_clk [27209]));
Q_ASSIGN U5566 ( .B(clk), .A(\g.we_clk [27208]));
Q_ASSIGN U5567 ( .B(clk), .A(\g.we_clk [27207]));
Q_ASSIGN U5568 ( .B(clk), .A(\g.we_clk [27206]));
Q_ASSIGN U5569 ( .B(clk), .A(\g.we_clk [27205]));
Q_ASSIGN U5570 ( .B(clk), .A(\g.we_clk [27204]));
Q_ASSIGN U5571 ( .B(clk), .A(\g.we_clk [27203]));
Q_ASSIGN U5572 ( .B(clk), .A(\g.we_clk [27202]));
Q_ASSIGN U5573 ( .B(clk), .A(\g.we_clk [27201]));
Q_ASSIGN U5574 ( .B(clk), .A(\g.we_clk [27200]));
Q_ASSIGN U5575 ( .B(clk), .A(\g.we_clk [27199]));
Q_ASSIGN U5576 ( .B(clk), .A(\g.we_clk [27198]));
Q_ASSIGN U5577 ( .B(clk), .A(\g.we_clk [27197]));
Q_ASSIGN U5578 ( .B(clk), .A(\g.we_clk [27196]));
Q_ASSIGN U5579 ( .B(clk), .A(\g.we_clk [27195]));
Q_ASSIGN U5580 ( .B(clk), .A(\g.we_clk [27194]));
Q_ASSIGN U5581 ( .B(clk), .A(\g.we_clk [27193]));
Q_ASSIGN U5582 ( .B(clk), .A(\g.we_clk [27192]));
Q_ASSIGN U5583 ( .B(clk), .A(\g.we_clk [27191]));
Q_ASSIGN U5584 ( .B(clk), .A(\g.we_clk [27190]));
Q_ASSIGN U5585 ( .B(clk), .A(\g.we_clk [27189]));
Q_ASSIGN U5586 ( .B(clk), .A(\g.we_clk [27188]));
Q_ASSIGN U5587 ( .B(clk), .A(\g.we_clk [27187]));
Q_ASSIGN U5588 ( .B(clk), .A(\g.we_clk [27186]));
Q_ASSIGN U5589 ( .B(clk), .A(\g.we_clk [27185]));
Q_ASSIGN U5590 ( .B(clk), .A(\g.we_clk [27184]));
Q_ASSIGN U5591 ( .B(clk), .A(\g.we_clk [27183]));
Q_ASSIGN U5592 ( .B(clk), .A(\g.we_clk [27182]));
Q_ASSIGN U5593 ( .B(clk), .A(\g.we_clk [27181]));
Q_ASSIGN U5594 ( .B(clk), .A(\g.we_clk [27180]));
Q_ASSIGN U5595 ( .B(clk), .A(\g.we_clk [27179]));
Q_ASSIGN U5596 ( .B(clk), .A(\g.we_clk [27178]));
Q_ASSIGN U5597 ( .B(clk), .A(\g.we_clk [27177]));
Q_ASSIGN U5598 ( .B(clk), .A(\g.we_clk [27176]));
Q_ASSIGN U5599 ( .B(clk), .A(\g.we_clk [27175]));
Q_ASSIGN U5600 ( .B(clk), .A(\g.we_clk [27174]));
Q_ASSIGN U5601 ( .B(clk), .A(\g.we_clk [27173]));
Q_ASSIGN U5602 ( .B(clk), .A(\g.we_clk [27172]));
Q_ASSIGN U5603 ( .B(clk), .A(\g.we_clk [27171]));
Q_ASSIGN U5604 ( .B(clk), .A(\g.we_clk [27170]));
Q_ASSIGN U5605 ( .B(clk), .A(\g.we_clk [27169]));
Q_ASSIGN U5606 ( .B(clk), .A(\g.we_clk [27168]));
Q_ASSIGN U5607 ( .B(clk), .A(\g.we_clk [27167]));
Q_ASSIGN U5608 ( .B(clk), .A(\g.we_clk [27166]));
Q_ASSIGN U5609 ( .B(clk), .A(\g.we_clk [27165]));
Q_ASSIGN U5610 ( .B(clk), .A(\g.we_clk [27164]));
Q_ASSIGN U5611 ( .B(clk), .A(\g.we_clk [27163]));
Q_ASSIGN U5612 ( .B(clk), .A(\g.we_clk [27162]));
Q_ASSIGN U5613 ( .B(clk), .A(\g.we_clk [27161]));
Q_ASSIGN U5614 ( .B(clk), .A(\g.we_clk [27160]));
Q_ASSIGN U5615 ( .B(clk), .A(\g.we_clk [27159]));
Q_ASSIGN U5616 ( .B(clk), .A(\g.we_clk [27158]));
Q_ASSIGN U5617 ( .B(clk), .A(\g.we_clk [27157]));
Q_ASSIGN U5618 ( .B(clk), .A(\g.we_clk [27156]));
Q_ASSIGN U5619 ( .B(clk), .A(\g.we_clk [27155]));
Q_ASSIGN U5620 ( .B(clk), .A(\g.we_clk [27154]));
Q_ASSIGN U5621 ( .B(clk), .A(\g.we_clk [27153]));
Q_ASSIGN U5622 ( .B(clk), .A(\g.we_clk [27152]));
Q_ASSIGN U5623 ( .B(clk), .A(\g.we_clk [27151]));
Q_ASSIGN U5624 ( .B(clk), .A(\g.we_clk [27150]));
Q_ASSIGN U5625 ( .B(clk), .A(\g.we_clk [27149]));
Q_ASSIGN U5626 ( .B(clk), .A(\g.we_clk [27148]));
Q_ASSIGN U5627 ( .B(clk), .A(\g.we_clk [27147]));
Q_ASSIGN U5628 ( .B(clk), .A(\g.we_clk [27146]));
Q_ASSIGN U5629 ( .B(clk), .A(\g.we_clk [27145]));
Q_ASSIGN U5630 ( .B(clk), .A(\g.we_clk [27144]));
Q_ASSIGN U5631 ( .B(clk), .A(\g.we_clk [27143]));
Q_ASSIGN U5632 ( .B(clk), .A(\g.we_clk [27142]));
Q_ASSIGN U5633 ( .B(clk), .A(\g.we_clk [27141]));
Q_ASSIGN U5634 ( .B(clk), .A(\g.we_clk [27140]));
Q_ASSIGN U5635 ( .B(clk), .A(\g.we_clk [27139]));
Q_ASSIGN U5636 ( .B(clk), .A(\g.we_clk [27138]));
Q_ASSIGN U5637 ( .B(clk), .A(\g.we_clk [27137]));
Q_ASSIGN U5638 ( .B(clk), .A(\g.we_clk [27136]));
Q_ASSIGN U5639 ( .B(clk), .A(\g.we_clk [27135]));
Q_ASSIGN U5640 ( .B(clk), .A(\g.we_clk [27134]));
Q_ASSIGN U5641 ( .B(clk), .A(\g.we_clk [27133]));
Q_ASSIGN U5642 ( .B(clk), .A(\g.we_clk [27132]));
Q_ASSIGN U5643 ( .B(clk), .A(\g.we_clk [27131]));
Q_ASSIGN U5644 ( .B(clk), .A(\g.we_clk [27130]));
Q_ASSIGN U5645 ( .B(clk), .A(\g.we_clk [27129]));
Q_ASSIGN U5646 ( .B(clk), .A(\g.we_clk [27128]));
Q_ASSIGN U5647 ( .B(clk), .A(\g.we_clk [27127]));
Q_ASSIGN U5648 ( .B(clk), .A(\g.we_clk [27126]));
Q_ASSIGN U5649 ( .B(clk), .A(\g.we_clk [27125]));
Q_ASSIGN U5650 ( .B(clk), .A(\g.we_clk [27124]));
Q_ASSIGN U5651 ( .B(clk), .A(\g.we_clk [27123]));
Q_ASSIGN U5652 ( .B(clk), .A(\g.we_clk [27122]));
Q_ASSIGN U5653 ( .B(clk), .A(\g.we_clk [27121]));
Q_ASSIGN U5654 ( .B(clk), .A(\g.we_clk [27120]));
Q_ASSIGN U5655 ( .B(clk), .A(\g.we_clk [27119]));
Q_ASSIGN U5656 ( .B(clk), .A(\g.we_clk [27118]));
Q_ASSIGN U5657 ( .B(clk), .A(\g.we_clk [27117]));
Q_ASSIGN U5658 ( .B(clk), .A(\g.we_clk [27116]));
Q_ASSIGN U5659 ( .B(clk), .A(\g.we_clk [27115]));
Q_ASSIGN U5660 ( .B(clk), .A(\g.we_clk [27114]));
Q_ASSIGN U5661 ( .B(clk), .A(\g.we_clk [27113]));
Q_ASSIGN U5662 ( .B(clk), .A(\g.we_clk [27112]));
Q_ASSIGN U5663 ( .B(clk), .A(\g.we_clk [27111]));
Q_ASSIGN U5664 ( .B(clk), .A(\g.we_clk [27110]));
Q_ASSIGN U5665 ( .B(clk), .A(\g.we_clk [27109]));
Q_ASSIGN U5666 ( .B(clk), .A(\g.we_clk [27108]));
Q_ASSIGN U5667 ( .B(clk), .A(\g.we_clk [27107]));
Q_ASSIGN U5668 ( .B(clk), .A(\g.we_clk [27106]));
Q_ASSIGN U5669 ( .B(clk), .A(\g.we_clk [27105]));
Q_ASSIGN U5670 ( .B(clk), .A(\g.we_clk [27104]));
Q_ASSIGN U5671 ( .B(clk), .A(\g.we_clk [27103]));
Q_ASSIGN U5672 ( .B(clk), .A(\g.we_clk [27102]));
Q_ASSIGN U5673 ( .B(clk), .A(\g.we_clk [27101]));
Q_ASSIGN U5674 ( .B(clk), .A(\g.we_clk [27100]));
Q_ASSIGN U5675 ( .B(clk), .A(\g.we_clk [27099]));
Q_ASSIGN U5676 ( .B(clk), .A(\g.we_clk [27098]));
Q_ASSIGN U5677 ( .B(clk), .A(\g.we_clk [27097]));
Q_ASSIGN U5678 ( .B(clk), .A(\g.we_clk [27096]));
Q_ASSIGN U5679 ( .B(clk), .A(\g.we_clk [27095]));
Q_ASSIGN U5680 ( .B(clk), .A(\g.we_clk [27094]));
Q_ASSIGN U5681 ( .B(clk), .A(\g.we_clk [27093]));
Q_ASSIGN U5682 ( .B(clk), .A(\g.we_clk [27092]));
Q_ASSIGN U5683 ( .B(clk), .A(\g.we_clk [27091]));
Q_ASSIGN U5684 ( .B(clk), .A(\g.we_clk [27090]));
Q_ASSIGN U5685 ( .B(clk), .A(\g.we_clk [27089]));
Q_ASSIGN U5686 ( .B(clk), .A(\g.we_clk [27088]));
Q_ASSIGN U5687 ( .B(clk), .A(\g.we_clk [27087]));
Q_ASSIGN U5688 ( .B(clk), .A(\g.we_clk [27086]));
Q_ASSIGN U5689 ( .B(clk), .A(\g.we_clk [27085]));
Q_ASSIGN U5690 ( .B(clk), .A(\g.we_clk [27084]));
Q_ASSIGN U5691 ( .B(clk), .A(\g.we_clk [27083]));
Q_ASSIGN U5692 ( .B(clk), .A(\g.we_clk [27082]));
Q_ASSIGN U5693 ( .B(clk), .A(\g.we_clk [27081]));
Q_ASSIGN U5694 ( .B(clk), .A(\g.we_clk [27080]));
Q_ASSIGN U5695 ( .B(clk), .A(\g.we_clk [27079]));
Q_ASSIGN U5696 ( .B(clk), .A(\g.we_clk [27078]));
Q_ASSIGN U5697 ( .B(clk), .A(\g.we_clk [27077]));
Q_ASSIGN U5698 ( .B(clk), .A(\g.we_clk [27076]));
Q_ASSIGN U5699 ( .B(clk), .A(\g.we_clk [27075]));
Q_ASSIGN U5700 ( .B(clk), .A(\g.we_clk [27074]));
Q_ASSIGN U5701 ( .B(clk), .A(\g.we_clk [27073]));
Q_ASSIGN U5702 ( .B(clk), .A(\g.we_clk [27072]));
Q_ASSIGN U5703 ( .B(clk), .A(\g.we_clk [27071]));
Q_ASSIGN U5704 ( .B(clk), .A(\g.we_clk [27070]));
Q_ASSIGN U5705 ( .B(clk), .A(\g.we_clk [27069]));
Q_ASSIGN U5706 ( .B(clk), .A(\g.we_clk [27068]));
Q_ASSIGN U5707 ( .B(clk), .A(\g.we_clk [27067]));
Q_ASSIGN U5708 ( .B(clk), .A(\g.we_clk [27066]));
Q_ASSIGN U5709 ( .B(clk), .A(\g.we_clk [27065]));
Q_ASSIGN U5710 ( .B(clk), .A(\g.we_clk [27064]));
Q_ASSIGN U5711 ( .B(clk), .A(\g.we_clk [27063]));
Q_ASSIGN U5712 ( .B(clk), .A(\g.we_clk [27062]));
Q_ASSIGN U5713 ( .B(clk), .A(\g.we_clk [27061]));
Q_ASSIGN U5714 ( .B(clk), .A(\g.we_clk [27060]));
Q_ASSIGN U5715 ( .B(clk), .A(\g.we_clk [27059]));
Q_ASSIGN U5716 ( .B(clk), .A(\g.we_clk [27058]));
Q_ASSIGN U5717 ( .B(clk), .A(\g.we_clk [27057]));
Q_ASSIGN U5718 ( .B(clk), .A(\g.we_clk [27056]));
Q_ASSIGN U5719 ( .B(clk), .A(\g.we_clk [27055]));
Q_ASSIGN U5720 ( .B(clk), .A(\g.we_clk [27054]));
Q_ASSIGN U5721 ( .B(clk), .A(\g.we_clk [27053]));
Q_ASSIGN U5722 ( .B(clk), .A(\g.we_clk [27052]));
Q_ASSIGN U5723 ( .B(clk), .A(\g.we_clk [27051]));
Q_ASSIGN U5724 ( .B(clk), .A(\g.we_clk [27050]));
Q_ASSIGN U5725 ( .B(clk), .A(\g.we_clk [27049]));
Q_ASSIGN U5726 ( .B(clk), .A(\g.we_clk [27048]));
Q_ASSIGN U5727 ( .B(clk), .A(\g.we_clk [27047]));
Q_ASSIGN U5728 ( .B(clk), .A(\g.we_clk [27046]));
Q_ASSIGN U5729 ( .B(clk), .A(\g.we_clk [27045]));
Q_ASSIGN U5730 ( .B(clk), .A(\g.we_clk [27044]));
Q_ASSIGN U5731 ( .B(clk), .A(\g.we_clk [27043]));
Q_ASSIGN U5732 ( .B(clk), .A(\g.we_clk [27042]));
Q_ASSIGN U5733 ( .B(clk), .A(\g.we_clk [27041]));
Q_ASSIGN U5734 ( .B(clk), .A(\g.we_clk [27040]));
Q_ASSIGN U5735 ( .B(clk), .A(\g.we_clk [27039]));
Q_ASSIGN U5736 ( .B(clk), .A(\g.we_clk [27038]));
Q_ASSIGN U5737 ( .B(clk), .A(\g.we_clk [27037]));
Q_ASSIGN U5738 ( .B(clk), .A(\g.we_clk [27036]));
Q_ASSIGN U5739 ( .B(clk), .A(\g.we_clk [27035]));
Q_ASSIGN U5740 ( .B(clk), .A(\g.we_clk [27034]));
Q_ASSIGN U5741 ( .B(clk), .A(\g.we_clk [27033]));
Q_ASSIGN U5742 ( .B(clk), .A(\g.we_clk [27032]));
Q_ASSIGN U5743 ( .B(clk), .A(\g.we_clk [27031]));
Q_ASSIGN U5744 ( .B(clk), .A(\g.we_clk [27030]));
Q_ASSIGN U5745 ( .B(clk), .A(\g.we_clk [27029]));
Q_ASSIGN U5746 ( .B(clk), .A(\g.we_clk [27028]));
Q_ASSIGN U5747 ( .B(clk), .A(\g.we_clk [27027]));
Q_ASSIGN U5748 ( .B(clk), .A(\g.we_clk [27026]));
Q_ASSIGN U5749 ( .B(clk), .A(\g.we_clk [27025]));
Q_ASSIGN U5750 ( .B(clk), .A(\g.we_clk [27024]));
Q_ASSIGN U5751 ( .B(clk), .A(\g.we_clk [27023]));
Q_ASSIGN U5752 ( .B(clk), .A(\g.we_clk [27022]));
Q_ASSIGN U5753 ( .B(clk), .A(\g.we_clk [27021]));
Q_ASSIGN U5754 ( .B(clk), .A(\g.we_clk [27020]));
Q_ASSIGN U5755 ( .B(clk), .A(\g.we_clk [27019]));
Q_ASSIGN U5756 ( .B(clk), .A(\g.we_clk [27018]));
Q_ASSIGN U5757 ( .B(clk), .A(\g.we_clk [27017]));
Q_ASSIGN U5758 ( .B(clk), .A(\g.we_clk [27016]));
Q_ASSIGN U5759 ( .B(clk), .A(\g.we_clk [27015]));
Q_ASSIGN U5760 ( .B(clk), .A(\g.we_clk [27014]));
Q_ASSIGN U5761 ( .B(clk), .A(\g.we_clk [27013]));
Q_ASSIGN U5762 ( .B(clk), .A(\g.we_clk [27012]));
Q_ASSIGN U5763 ( .B(clk), .A(\g.we_clk [27011]));
Q_ASSIGN U5764 ( .B(clk), .A(\g.we_clk [27010]));
Q_ASSIGN U5765 ( .B(clk), .A(\g.we_clk [27009]));
Q_ASSIGN U5766 ( .B(clk), .A(\g.we_clk [27008]));
Q_ASSIGN U5767 ( .B(clk), .A(\g.we_clk [27007]));
Q_ASSIGN U5768 ( .B(clk), .A(\g.we_clk [27006]));
Q_ASSIGN U5769 ( .B(clk), .A(\g.we_clk [27005]));
Q_ASSIGN U5770 ( .B(clk), .A(\g.we_clk [27004]));
Q_ASSIGN U5771 ( .B(clk), .A(\g.we_clk [27003]));
Q_ASSIGN U5772 ( .B(clk), .A(\g.we_clk [27002]));
Q_ASSIGN U5773 ( .B(clk), .A(\g.we_clk [27001]));
Q_ASSIGN U5774 ( .B(clk), .A(\g.we_clk [27000]));
Q_ASSIGN U5775 ( .B(clk), .A(\g.we_clk [26999]));
Q_ASSIGN U5776 ( .B(clk), .A(\g.we_clk [26998]));
Q_ASSIGN U5777 ( .B(clk), .A(\g.we_clk [26997]));
Q_ASSIGN U5778 ( .B(clk), .A(\g.we_clk [26996]));
Q_ASSIGN U5779 ( .B(clk), .A(\g.we_clk [26995]));
Q_ASSIGN U5780 ( .B(clk), .A(\g.we_clk [26994]));
Q_ASSIGN U5781 ( .B(clk), .A(\g.we_clk [26993]));
Q_ASSIGN U5782 ( .B(clk), .A(\g.we_clk [26992]));
Q_ASSIGN U5783 ( .B(clk), .A(\g.we_clk [26991]));
Q_ASSIGN U5784 ( .B(clk), .A(\g.we_clk [26990]));
Q_ASSIGN U5785 ( .B(clk), .A(\g.we_clk [26989]));
Q_ASSIGN U5786 ( .B(clk), .A(\g.we_clk [26988]));
Q_ASSIGN U5787 ( .B(clk), .A(\g.we_clk [26987]));
Q_ASSIGN U5788 ( .B(clk), .A(\g.we_clk [26986]));
Q_ASSIGN U5789 ( .B(clk), .A(\g.we_clk [26985]));
Q_ASSIGN U5790 ( .B(clk), .A(\g.we_clk [26984]));
Q_ASSIGN U5791 ( .B(clk), .A(\g.we_clk [26983]));
Q_ASSIGN U5792 ( .B(clk), .A(\g.we_clk [26982]));
Q_ASSIGN U5793 ( .B(clk), .A(\g.we_clk [26981]));
Q_ASSIGN U5794 ( .B(clk), .A(\g.we_clk [26980]));
Q_ASSIGN U5795 ( .B(clk), .A(\g.we_clk [26979]));
Q_ASSIGN U5796 ( .B(clk), .A(\g.we_clk [26978]));
Q_ASSIGN U5797 ( .B(clk), .A(\g.we_clk [26977]));
Q_ASSIGN U5798 ( .B(clk), .A(\g.we_clk [26976]));
Q_ASSIGN U5799 ( .B(clk), .A(\g.we_clk [26975]));
Q_ASSIGN U5800 ( .B(clk), .A(\g.we_clk [26974]));
Q_ASSIGN U5801 ( .B(clk), .A(\g.we_clk [26973]));
Q_ASSIGN U5802 ( .B(clk), .A(\g.we_clk [26972]));
Q_ASSIGN U5803 ( .B(clk), .A(\g.we_clk [26971]));
Q_ASSIGN U5804 ( .B(clk), .A(\g.we_clk [26970]));
Q_ASSIGN U5805 ( .B(clk), .A(\g.we_clk [26969]));
Q_ASSIGN U5806 ( .B(clk), .A(\g.we_clk [26968]));
Q_ASSIGN U5807 ( .B(clk), .A(\g.we_clk [26967]));
Q_ASSIGN U5808 ( .B(clk), .A(\g.we_clk [26966]));
Q_ASSIGN U5809 ( .B(clk), .A(\g.we_clk [26965]));
Q_ASSIGN U5810 ( .B(clk), .A(\g.we_clk [26964]));
Q_ASSIGN U5811 ( .B(clk), .A(\g.we_clk [26963]));
Q_ASSIGN U5812 ( .B(clk), .A(\g.we_clk [26962]));
Q_ASSIGN U5813 ( .B(clk), .A(\g.we_clk [26961]));
Q_ASSIGN U5814 ( .B(clk), .A(\g.we_clk [26960]));
Q_ASSIGN U5815 ( .B(clk), .A(\g.we_clk [26959]));
Q_ASSIGN U5816 ( .B(clk), .A(\g.we_clk [26958]));
Q_ASSIGN U5817 ( .B(clk), .A(\g.we_clk [26957]));
Q_ASSIGN U5818 ( .B(clk), .A(\g.we_clk [26956]));
Q_ASSIGN U5819 ( .B(clk), .A(\g.we_clk [26955]));
Q_ASSIGN U5820 ( .B(clk), .A(\g.we_clk [26954]));
Q_ASSIGN U5821 ( .B(clk), .A(\g.we_clk [26953]));
Q_ASSIGN U5822 ( .B(clk), .A(\g.we_clk [26952]));
Q_ASSIGN U5823 ( .B(clk), .A(\g.we_clk [26951]));
Q_ASSIGN U5824 ( .B(clk), .A(\g.we_clk [26950]));
Q_ASSIGN U5825 ( .B(clk), .A(\g.we_clk [26949]));
Q_ASSIGN U5826 ( .B(clk), .A(\g.we_clk [26948]));
Q_ASSIGN U5827 ( .B(clk), .A(\g.we_clk [26947]));
Q_ASSIGN U5828 ( .B(clk), .A(\g.we_clk [26946]));
Q_ASSIGN U5829 ( .B(clk), .A(\g.we_clk [26945]));
Q_ASSIGN U5830 ( .B(clk), .A(\g.we_clk [26944]));
Q_ASSIGN U5831 ( .B(clk), .A(\g.we_clk [26943]));
Q_ASSIGN U5832 ( .B(clk), .A(\g.we_clk [26942]));
Q_ASSIGN U5833 ( .B(clk), .A(\g.we_clk [26941]));
Q_ASSIGN U5834 ( .B(clk), .A(\g.we_clk [26940]));
Q_ASSIGN U5835 ( .B(clk), .A(\g.we_clk [26939]));
Q_ASSIGN U5836 ( .B(clk), .A(\g.we_clk [26938]));
Q_ASSIGN U5837 ( .B(clk), .A(\g.we_clk [26937]));
Q_ASSIGN U5838 ( .B(clk), .A(\g.we_clk [26936]));
Q_ASSIGN U5839 ( .B(clk), .A(\g.we_clk [26935]));
Q_ASSIGN U5840 ( .B(clk), .A(\g.we_clk [26934]));
Q_ASSIGN U5841 ( .B(clk), .A(\g.we_clk [26933]));
Q_ASSIGN U5842 ( .B(clk), .A(\g.we_clk [26932]));
Q_ASSIGN U5843 ( .B(clk), .A(\g.we_clk [26931]));
Q_ASSIGN U5844 ( .B(clk), .A(\g.we_clk [26930]));
Q_ASSIGN U5845 ( .B(clk), .A(\g.we_clk [26929]));
Q_ASSIGN U5846 ( .B(clk), .A(\g.we_clk [26928]));
Q_ASSIGN U5847 ( .B(clk), .A(\g.we_clk [26927]));
Q_ASSIGN U5848 ( .B(clk), .A(\g.we_clk [26926]));
Q_ASSIGN U5849 ( .B(clk), .A(\g.we_clk [26925]));
Q_ASSIGN U5850 ( .B(clk), .A(\g.we_clk [26924]));
Q_ASSIGN U5851 ( .B(clk), .A(\g.we_clk [26923]));
Q_ASSIGN U5852 ( .B(clk), .A(\g.we_clk [26922]));
Q_ASSIGN U5853 ( .B(clk), .A(\g.we_clk [26921]));
Q_ASSIGN U5854 ( .B(clk), .A(\g.we_clk [26920]));
Q_ASSIGN U5855 ( .B(clk), .A(\g.we_clk [26919]));
Q_ASSIGN U5856 ( .B(clk), .A(\g.we_clk [26918]));
Q_ASSIGN U5857 ( .B(clk), .A(\g.we_clk [26917]));
Q_ASSIGN U5858 ( .B(clk), .A(\g.we_clk [26916]));
Q_ASSIGN U5859 ( .B(clk), .A(\g.we_clk [26915]));
Q_ASSIGN U5860 ( .B(clk), .A(\g.we_clk [26914]));
Q_ASSIGN U5861 ( .B(clk), .A(\g.we_clk [26913]));
Q_ASSIGN U5862 ( .B(clk), .A(\g.we_clk [26912]));
Q_ASSIGN U5863 ( .B(clk), .A(\g.we_clk [26911]));
Q_ASSIGN U5864 ( .B(clk), .A(\g.we_clk [26910]));
Q_ASSIGN U5865 ( .B(clk), .A(\g.we_clk [26909]));
Q_ASSIGN U5866 ( .B(clk), .A(\g.we_clk [26908]));
Q_ASSIGN U5867 ( .B(clk), .A(\g.we_clk [26907]));
Q_ASSIGN U5868 ( .B(clk), .A(\g.we_clk [26906]));
Q_ASSIGN U5869 ( .B(clk), .A(\g.we_clk [26905]));
Q_ASSIGN U5870 ( .B(clk), .A(\g.we_clk [26904]));
Q_ASSIGN U5871 ( .B(clk), .A(\g.we_clk [26903]));
Q_ASSIGN U5872 ( .B(clk), .A(\g.we_clk [26902]));
Q_ASSIGN U5873 ( .B(clk), .A(\g.we_clk [26901]));
Q_ASSIGN U5874 ( .B(clk), .A(\g.we_clk [26900]));
Q_ASSIGN U5875 ( .B(clk), .A(\g.we_clk [26899]));
Q_ASSIGN U5876 ( .B(clk), .A(\g.we_clk [26898]));
Q_ASSIGN U5877 ( .B(clk), .A(\g.we_clk [26897]));
Q_ASSIGN U5878 ( .B(clk), .A(\g.we_clk [26896]));
Q_ASSIGN U5879 ( .B(clk), .A(\g.we_clk [26895]));
Q_ASSIGN U5880 ( .B(clk), .A(\g.we_clk [26894]));
Q_ASSIGN U5881 ( .B(clk), .A(\g.we_clk [26893]));
Q_ASSIGN U5882 ( .B(clk), .A(\g.we_clk [26892]));
Q_ASSIGN U5883 ( .B(clk), .A(\g.we_clk [26891]));
Q_ASSIGN U5884 ( .B(clk), .A(\g.we_clk [26890]));
Q_ASSIGN U5885 ( .B(clk), .A(\g.we_clk [26889]));
Q_ASSIGN U5886 ( .B(clk), .A(\g.we_clk [26888]));
Q_ASSIGN U5887 ( .B(clk), .A(\g.we_clk [26887]));
Q_ASSIGN U5888 ( .B(clk), .A(\g.we_clk [26886]));
Q_ASSIGN U5889 ( .B(clk), .A(\g.we_clk [26885]));
Q_ASSIGN U5890 ( .B(clk), .A(\g.we_clk [26884]));
Q_ASSIGN U5891 ( .B(clk), .A(\g.we_clk [26883]));
Q_ASSIGN U5892 ( .B(clk), .A(\g.we_clk [26882]));
Q_ASSIGN U5893 ( .B(clk), .A(\g.we_clk [26881]));
Q_ASSIGN U5894 ( .B(clk), .A(\g.we_clk [26880]));
Q_ASSIGN U5895 ( .B(clk), .A(\g.we_clk [26879]));
Q_ASSIGN U5896 ( .B(clk), .A(\g.we_clk [26878]));
Q_ASSIGN U5897 ( .B(clk), .A(\g.we_clk [26877]));
Q_ASSIGN U5898 ( .B(clk), .A(\g.we_clk [26876]));
Q_ASSIGN U5899 ( .B(clk), .A(\g.we_clk [26875]));
Q_ASSIGN U5900 ( .B(clk), .A(\g.we_clk [26874]));
Q_ASSIGN U5901 ( .B(clk), .A(\g.we_clk [26873]));
Q_ASSIGN U5902 ( .B(clk), .A(\g.we_clk [26872]));
Q_ASSIGN U5903 ( .B(clk), .A(\g.we_clk [26871]));
Q_ASSIGN U5904 ( .B(clk), .A(\g.we_clk [26870]));
Q_ASSIGN U5905 ( .B(clk), .A(\g.we_clk [26869]));
Q_ASSIGN U5906 ( .B(clk), .A(\g.we_clk [26868]));
Q_ASSIGN U5907 ( .B(clk), .A(\g.we_clk [26867]));
Q_ASSIGN U5908 ( .B(clk), .A(\g.we_clk [26866]));
Q_ASSIGN U5909 ( .B(clk), .A(\g.we_clk [26865]));
Q_ASSIGN U5910 ( .B(clk), .A(\g.we_clk [26864]));
Q_ASSIGN U5911 ( .B(clk), .A(\g.we_clk [26863]));
Q_ASSIGN U5912 ( .B(clk), .A(\g.we_clk [26862]));
Q_ASSIGN U5913 ( .B(clk), .A(\g.we_clk [26861]));
Q_ASSIGN U5914 ( .B(clk), .A(\g.we_clk [26860]));
Q_ASSIGN U5915 ( .B(clk), .A(\g.we_clk [26859]));
Q_ASSIGN U5916 ( .B(clk), .A(\g.we_clk [26858]));
Q_ASSIGN U5917 ( .B(clk), .A(\g.we_clk [26857]));
Q_ASSIGN U5918 ( .B(clk), .A(\g.we_clk [26856]));
Q_ASSIGN U5919 ( .B(clk), .A(\g.we_clk [26855]));
Q_ASSIGN U5920 ( .B(clk), .A(\g.we_clk [26854]));
Q_ASSIGN U5921 ( .B(clk), .A(\g.we_clk [26853]));
Q_ASSIGN U5922 ( .B(clk), .A(\g.we_clk [26852]));
Q_ASSIGN U5923 ( .B(clk), .A(\g.we_clk [26851]));
Q_ASSIGN U5924 ( .B(clk), .A(\g.we_clk [26850]));
Q_ASSIGN U5925 ( .B(clk), .A(\g.we_clk [26849]));
Q_ASSIGN U5926 ( .B(clk), .A(\g.we_clk [26848]));
Q_ASSIGN U5927 ( .B(clk), .A(\g.we_clk [26847]));
Q_ASSIGN U5928 ( .B(clk), .A(\g.we_clk [26846]));
Q_ASSIGN U5929 ( .B(clk), .A(\g.we_clk [26845]));
Q_ASSIGN U5930 ( .B(clk), .A(\g.we_clk [26844]));
Q_ASSIGN U5931 ( .B(clk), .A(\g.we_clk [26843]));
Q_ASSIGN U5932 ( .B(clk), .A(\g.we_clk [26842]));
Q_ASSIGN U5933 ( .B(clk), .A(\g.we_clk [26841]));
Q_ASSIGN U5934 ( .B(clk), .A(\g.we_clk [26840]));
Q_ASSIGN U5935 ( .B(clk), .A(\g.we_clk [26839]));
Q_ASSIGN U5936 ( .B(clk), .A(\g.we_clk [26838]));
Q_ASSIGN U5937 ( .B(clk), .A(\g.we_clk [26837]));
Q_ASSIGN U5938 ( .B(clk), .A(\g.we_clk [26836]));
Q_ASSIGN U5939 ( .B(clk), .A(\g.we_clk [26835]));
Q_ASSIGN U5940 ( .B(clk), .A(\g.we_clk [26834]));
Q_ASSIGN U5941 ( .B(clk), .A(\g.we_clk [26833]));
Q_ASSIGN U5942 ( .B(clk), .A(\g.we_clk [26832]));
Q_ASSIGN U5943 ( .B(clk), .A(\g.we_clk [26831]));
Q_ASSIGN U5944 ( .B(clk), .A(\g.we_clk [26830]));
Q_ASSIGN U5945 ( .B(clk), .A(\g.we_clk [26829]));
Q_ASSIGN U5946 ( .B(clk), .A(\g.we_clk [26828]));
Q_ASSIGN U5947 ( .B(clk), .A(\g.we_clk [26827]));
Q_ASSIGN U5948 ( .B(clk), .A(\g.we_clk [26826]));
Q_ASSIGN U5949 ( .B(clk), .A(\g.we_clk [26825]));
Q_ASSIGN U5950 ( .B(clk), .A(\g.we_clk [26824]));
Q_ASSIGN U5951 ( .B(clk), .A(\g.we_clk [26823]));
Q_ASSIGN U5952 ( .B(clk), .A(\g.we_clk [26822]));
Q_ASSIGN U5953 ( .B(clk), .A(\g.we_clk [26821]));
Q_ASSIGN U5954 ( .B(clk), .A(\g.we_clk [26820]));
Q_ASSIGN U5955 ( .B(clk), .A(\g.we_clk [26819]));
Q_ASSIGN U5956 ( .B(clk), .A(\g.we_clk [26818]));
Q_ASSIGN U5957 ( .B(clk), .A(\g.we_clk [26817]));
Q_ASSIGN U5958 ( .B(clk), .A(\g.we_clk [26816]));
Q_ASSIGN U5959 ( .B(clk), .A(\g.we_clk [26815]));
Q_ASSIGN U5960 ( .B(clk), .A(\g.we_clk [26814]));
Q_ASSIGN U5961 ( .B(clk), .A(\g.we_clk [26813]));
Q_ASSIGN U5962 ( .B(clk), .A(\g.we_clk [26812]));
Q_ASSIGN U5963 ( .B(clk), .A(\g.we_clk [26811]));
Q_ASSIGN U5964 ( .B(clk), .A(\g.we_clk [26810]));
Q_ASSIGN U5965 ( .B(clk), .A(\g.we_clk [26809]));
Q_ASSIGN U5966 ( .B(clk), .A(\g.we_clk [26808]));
Q_ASSIGN U5967 ( .B(clk), .A(\g.we_clk [26807]));
Q_ASSIGN U5968 ( .B(clk), .A(\g.we_clk [26806]));
Q_ASSIGN U5969 ( .B(clk), .A(\g.we_clk [26805]));
Q_ASSIGN U5970 ( .B(clk), .A(\g.we_clk [26804]));
Q_ASSIGN U5971 ( .B(clk), .A(\g.we_clk [26803]));
Q_ASSIGN U5972 ( .B(clk), .A(\g.we_clk [26802]));
Q_ASSIGN U5973 ( .B(clk), .A(\g.we_clk [26801]));
Q_ASSIGN U5974 ( .B(clk), .A(\g.we_clk [26800]));
Q_ASSIGN U5975 ( .B(clk), .A(\g.we_clk [26799]));
Q_ASSIGN U5976 ( .B(clk), .A(\g.we_clk [26798]));
Q_ASSIGN U5977 ( .B(clk), .A(\g.we_clk [26797]));
Q_ASSIGN U5978 ( .B(clk), .A(\g.we_clk [26796]));
Q_ASSIGN U5979 ( .B(clk), .A(\g.we_clk [26795]));
Q_ASSIGN U5980 ( .B(clk), .A(\g.we_clk [26794]));
Q_ASSIGN U5981 ( .B(clk), .A(\g.we_clk [26793]));
Q_ASSIGN U5982 ( .B(clk), .A(\g.we_clk [26792]));
Q_ASSIGN U5983 ( .B(clk), .A(\g.we_clk [26791]));
Q_ASSIGN U5984 ( .B(clk), .A(\g.we_clk [26790]));
Q_ASSIGN U5985 ( .B(clk), .A(\g.we_clk [26789]));
Q_ASSIGN U5986 ( .B(clk), .A(\g.we_clk [26788]));
Q_ASSIGN U5987 ( .B(clk), .A(\g.we_clk [26787]));
Q_ASSIGN U5988 ( .B(clk), .A(\g.we_clk [26786]));
Q_ASSIGN U5989 ( .B(clk), .A(\g.we_clk [26785]));
Q_ASSIGN U5990 ( .B(clk), .A(\g.we_clk [26784]));
Q_ASSIGN U5991 ( .B(clk), .A(\g.we_clk [26783]));
Q_ASSIGN U5992 ( .B(clk), .A(\g.we_clk [26782]));
Q_ASSIGN U5993 ( .B(clk), .A(\g.we_clk [26781]));
Q_ASSIGN U5994 ( .B(clk), .A(\g.we_clk [26780]));
Q_ASSIGN U5995 ( .B(clk), .A(\g.we_clk [26779]));
Q_ASSIGN U5996 ( .B(clk), .A(\g.we_clk [26778]));
Q_ASSIGN U5997 ( .B(clk), .A(\g.we_clk [26777]));
Q_ASSIGN U5998 ( .B(clk), .A(\g.we_clk [26776]));
Q_ASSIGN U5999 ( .B(clk), .A(\g.we_clk [26775]));
Q_ASSIGN U6000 ( .B(clk), .A(\g.we_clk [26774]));
Q_ASSIGN U6001 ( .B(clk), .A(\g.we_clk [26773]));
Q_ASSIGN U6002 ( .B(clk), .A(\g.we_clk [26772]));
Q_ASSIGN U6003 ( .B(clk), .A(\g.we_clk [26771]));
Q_ASSIGN U6004 ( .B(clk), .A(\g.we_clk [26770]));
Q_ASSIGN U6005 ( .B(clk), .A(\g.we_clk [26769]));
Q_ASSIGN U6006 ( .B(clk), .A(\g.we_clk [26768]));
Q_ASSIGN U6007 ( .B(clk), .A(\g.we_clk [26767]));
Q_ASSIGN U6008 ( .B(clk), .A(\g.we_clk [26766]));
Q_ASSIGN U6009 ( .B(clk), .A(\g.we_clk [26765]));
Q_ASSIGN U6010 ( .B(clk), .A(\g.we_clk [26764]));
Q_ASSIGN U6011 ( .B(clk), .A(\g.we_clk [26763]));
Q_ASSIGN U6012 ( .B(clk), .A(\g.we_clk [26762]));
Q_ASSIGN U6013 ( .B(clk), .A(\g.we_clk [26761]));
Q_ASSIGN U6014 ( .B(clk), .A(\g.we_clk [26760]));
Q_ASSIGN U6015 ( .B(clk), .A(\g.we_clk [26759]));
Q_ASSIGN U6016 ( .B(clk), .A(\g.we_clk [26758]));
Q_ASSIGN U6017 ( .B(clk), .A(\g.we_clk [26757]));
Q_ASSIGN U6018 ( .B(clk), .A(\g.we_clk [26756]));
Q_ASSIGN U6019 ( .B(clk), .A(\g.we_clk [26755]));
Q_ASSIGN U6020 ( .B(clk), .A(\g.we_clk [26754]));
Q_ASSIGN U6021 ( .B(clk), .A(\g.we_clk [26753]));
Q_ASSIGN U6022 ( .B(clk), .A(\g.we_clk [26752]));
Q_ASSIGN U6023 ( .B(clk), .A(\g.we_clk [26751]));
Q_ASSIGN U6024 ( .B(clk), .A(\g.we_clk [26750]));
Q_ASSIGN U6025 ( .B(clk), .A(\g.we_clk [26749]));
Q_ASSIGN U6026 ( .B(clk), .A(\g.we_clk [26748]));
Q_ASSIGN U6027 ( .B(clk), .A(\g.we_clk [26747]));
Q_ASSIGN U6028 ( .B(clk), .A(\g.we_clk [26746]));
Q_ASSIGN U6029 ( .B(clk), .A(\g.we_clk [26745]));
Q_ASSIGN U6030 ( .B(clk), .A(\g.we_clk [26744]));
Q_ASSIGN U6031 ( .B(clk), .A(\g.we_clk [26743]));
Q_ASSIGN U6032 ( .B(clk), .A(\g.we_clk [26742]));
Q_ASSIGN U6033 ( .B(clk), .A(\g.we_clk [26741]));
Q_ASSIGN U6034 ( .B(clk), .A(\g.we_clk [26740]));
Q_ASSIGN U6035 ( .B(clk), .A(\g.we_clk [26739]));
Q_ASSIGN U6036 ( .B(clk), .A(\g.we_clk [26738]));
Q_ASSIGN U6037 ( .B(clk), .A(\g.we_clk [26737]));
Q_ASSIGN U6038 ( .B(clk), .A(\g.we_clk [26736]));
Q_ASSIGN U6039 ( .B(clk), .A(\g.we_clk [26735]));
Q_ASSIGN U6040 ( .B(clk), .A(\g.we_clk [26734]));
Q_ASSIGN U6041 ( .B(clk), .A(\g.we_clk [26733]));
Q_ASSIGN U6042 ( .B(clk), .A(\g.we_clk [26732]));
Q_ASSIGN U6043 ( .B(clk), .A(\g.we_clk [26731]));
Q_ASSIGN U6044 ( .B(clk), .A(\g.we_clk [26730]));
Q_ASSIGN U6045 ( .B(clk), .A(\g.we_clk [26729]));
Q_ASSIGN U6046 ( .B(clk), .A(\g.we_clk [26728]));
Q_ASSIGN U6047 ( .B(clk), .A(\g.we_clk [26727]));
Q_ASSIGN U6048 ( .B(clk), .A(\g.we_clk [26726]));
Q_ASSIGN U6049 ( .B(clk), .A(\g.we_clk [26725]));
Q_ASSIGN U6050 ( .B(clk), .A(\g.we_clk [26724]));
Q_ASSIGN U6051 ( .B(clk), .A(\g.we_clk [26723]));
Q_ASSIGN U6052 ( .B(clk), .A(\g.we_clk [26722]));
Q_ASSIGN U6053 ( .B(clk), .A(\g.we_clk [26721]));
Q_ASSIGN U6054 ( .B(clk), .A(\g.we_clk [26720]));
Q_ASSIGN U6055 ( .B(clk), .A(\g.we_clk [26719]));
Q_ASSIGN U6056 ( .B(clk), .A(\g.we_clk [26718]));
Q_ASSIGN U6057 ( .B(clk), .A(\g.we_clk [26717]));
Q_ASSIGN U6058 ( .B(clk), .A(\g.we_clk [26716]));
Q_ASSIGN U6059 ( .B(clk), .A(\g.we_clk [26715]));
Q_ASSIGN U6060 ( .B(clk), .A(\g.we_clk [26714]));
Q_ASSIGN U6061 ( .B(clk), .A(\g.we_clk [26713]));
Q_ASSIGN U6062 ( .B(clk), .A(\g.we_clk [26712]));
Q_ASSIGN U6063 ( .B(clk), .A(\g.we_clk [26711]));
Q_ASSIGN U6064 ( .B(clk), .A(\g.we_clk [26710]));
Q_ASSIGN U6065 ( .B(clk), .A(\g.we_clk [26709]));
Q_ASSIGN U6066 ( .B(clk), .A(\g.we_clk [26708]));
Q_ASSIGN U6067 ( .B(clk), .A(\g.we_clk [26707]));
Q_ASSIGN U6068 ( .B(clk), .A(\g.we_clk [26706]));
Q_ASSIGN U6069 ( .B(clk), .A(\g.we_clk [26705]));
Q_ASSIGN U6070 ( .B(clk), .A(\g.we_clk [26704]));
Q_ASSIGN U6071 ( .B(clk), .A(\g.we_clk [26703]));
Q_ASSIGN U6072 ( .B(clk), .A(\g.we_clk [26702]));
Q_ASSIGN U6073 ( .B(clk), .A(\g.we_clk [26701]));
Q_ASSIGN U6074 ( .B(clk), .A(\g.we_clk [26700]));
Q_ASSIGN U6075 ( .B(clk), .A(\g.we_clk [26699]));
Q_ASSIGN U6076 ( .B(clk), .A(\g.we_clk [26698]));
Q_ASSIGN U6077 ( .B(clk), .A(\g.we_clk [26697]));
Q_ASSIGN U6078 ( .B(clk), .A(\g.we_clk [26696]));
Q_ASSIGN U6079 ( .B(clk), .A(\g.we_clk [26695]));
Q_ASSIGN U6080 ( .B(clk), .A(\g.we_clk [26694]));
Q_ASSIGN U6081 ( .B(clk), .A(\g.we_clk [26693]));
Q_ASSIGN U6082 ( .B(clk), .A(\g.we_clk [26692]));
Q_ASSIGN U6083 ( .B(clk), .A(\g.we_clk [26691]));
Q_ASSIGN U6084 ( .B(clk), .A(\g.we_clk [26690]));
Q_ASSIGN U6085 ( .B(clk), .A(\g.we_clk [26689]));
Q_ASSIGN U6086 ( .B(clk), .A(\g.we_clk [26688]));
Q_ASSIGN U6087 ( .B(clk), .A(\g.we_clk [26687]));
Q_ASSIGN U6088 ( .B(clk), .A(\g.we_clk [26686]));
Q_ASSIGN U6089 ( .B(clk), .A(\g.we_clk [26685]));
Q_ASSIGN U6090 ( .B(clk), .A(\g.we_clk [26684]));
Q_ASSIGN U6091 ( .B(clk), .A(\g.we_clk [26683]));
Q_ASSIGN U6092 ( .B(clk), .A(\g.we_clk [26682]));
Q_ASSIGN U6093 ( .B(clk), .A(\g.we_clk [26681]));
Q_ASSIGN U6094 ( .B(clk), .A(\g.we_clk [26680]));
Q_ASSIGN U6095 ( .B(clk), .A(\g.we_clk [26679]));
Q_ASSIGN U6096 ( .B(clk), .A(\g.we_clk [26678]));
Q_ASSIGN U6097 ( .B(clk), .A(\g.we_clk [26677]));
Q_ASSIGN U6098 ( .B(clk), .A(\g.we_clk [26676]));
Q_ASSIGN U6099 ( .B(clk), .A(\g.we_clk [26675]));
Q_ASSIGN U6100 ( .B(clk), .A(\g.we_clk [26674]));
Q_ASSIGN U6101 ( .B(clk), .A(\g.we_clk [26673]));
Q_ASSIGN U6102 ( .B(clk), .A(\g.we_clk [26672]));
Q_ASSIGN U6103 ( .B(clk), .A(\g.we_clk [26671]));
Q_ASSIGN U6104 ( .B(clk), .A(\g.we_clk [26670]));
Q_ASSIGN U6105 ( .B(clk), .A(\g.we_clk [26669]));
Q_ASSIGN U6106 ( .B(clk), .A(\g.we_clk [26668]));
Q_ASSIGN U6107 ( .B(clk), .A(\g.we_clk [26667]));
Q_ASSIGN U6108 ( .B(clk), .A(\g.we_clk [26666]));
Q_ASSIGN U6109 ( .B(clk), .A(\g.we_clk [26665]));
Q_ASSIGN U6110 ( .B(clk), .A(\g.we_clk [26664]));
Q_ASSIGN U6111 ( .B(clk), .A(\g.we_clk [26663]));
Q_ASSIGN U6112 ( .B(clk), .A(\g.we_clk [26662]));
Q_ASSIGN U6113 ( .B(clk), .A(\g.we_clk [26661]));
Q_ASSIGN U6114 ( .B(clk), .A(\g.we_clk [26660]));
Q_ASSIGN U6115 ( .B(clk), .A(\g.we_clk [26659]));
Q_ASSIGN U6116 ( .B(clk), .A(\g.we_clk [26658]));
Q_ASSIGN U6117 ( .B(clk), .A(\g.we_clk [26657]));
Q_ASSIGN U6118 ( .B(clk), .A(\g.we_clk [26656]));
Q_ASSIGN U6119 ( .B(clk), .A(\g.we_clk [26655]));
Q_ASSIGN U6120 ( .B(clk), .A(\g.we_clk [26654]));
Q_ASSIGN U6121 ( .B(clk), .A(\g.we_clk [26653]));
Q_ASSIGN U6122 ( .B(clk), .A(\g.we_clk [26652]));
Q_ASSIGN U6123 ( .B(clk), .A(\g.we_clk [26651]));
Q_ASSIGN U6124 ( .B(clk), .A(\g.we_clk [26650]));
Q_ASSIGN U6125 ( .B(clk), .A(\g.we_clk [26649]));
Q_ASSIGN U6126 ( .B(clk), .A(\g.we_clk [26648]));
Q_ASSIGN U6127 ( .B(clk), .A(\g.we_clk [26647]));
Q_ASSIGN U6128 ( .B(clk), .A(\g.we_clk [26646]));
Q_ASSIGN U6129 ( .B(clk), .A(\g.we_clk [26645]));
Q_ASSIGN U6130 ( .B(clk), .A(\g.we_clk [26644]));
Q_ASSIGN U6131 ( .B(clk), .A(\g.we_clk [26643]));
Q_ASSIGN U6132 ( .B(clk), .A(\g.we_clk [26642]));
Q_ASSIGN U6133 ( .B(clk), .A(\g.we_clk [26641]));
Q_ASSIGN U6134 ( .B(clk), .A(\g.we_clk [26640]));
Q_ASSIGN U6135 ( .B(clk), .A(\g.we_clk [26639]));
Q_ASSIGN U6136 ( .B(clk), .A(\g.we_clk [26638]));
Q_ASSIGN U6137 ( .B(clk), .A(\g.we_clk [26637]));
Q_ASSIGN U6138 ( .B(clk), .A(\g.we_clk [26636]));
Q_ASSIGN U6139 ( .B(clk), .A(\g.we_clk [26635]));
Q_ASSIGN U6140 ( .B(clk), .A(\g.we_clk [26634]));
Q_ASSIGN U6141 ( .B(clk), .A(\g.we_clk [26633]));
Q_ASSIGN U6142 ( .B(clk), .A(\g.we_clk [26632]));
Q_ASSIGN U6143 ( .B(clk), .A(\g.we_clk [26631]));
Q_ASSIGN U6144 ( .B(clk), .A(\g.we_clk [26630]));
Q_ASSIGN U6145 ( .B(clk), .A(\g.we_clk [26629]));
Q_ASSIGN U6146 ( .B(clk), .A(\g.we_clk [26628]));
Q_ASSIGN U6147 ( .B(clk), .A(\g.we_clk [26627]));
Q_ASSIGN U6148 ( .B(clk), .A(\g.we_clk [26626]));
Q_ASSIGN U6149 ( .B(clk), .A(\g.we_clk [26625]));
Q_ASSIGN U6150 ( .B(clk), .A(\g.we_clk [26624]));
Q_ASSIGN U6151 ( .B(clk), .A(\g.we_clk [26623]));
Q_ASSIGN U6152 ( .B(clk), .A(\g.we_clk [26622]));
Q_ASSIGN U6153 ( .B(clk), .A(\g.we_clk [26621]));
Q_ASSIGN U6154 ( .B(clk), .A(\g.we_clk [26620]));
Q_ASSIGN U6155 ( .B(clk), .A(\g.we_clk [26619]));
Q_ASSIGN U6156 ( .B(clk), .A(\g.we_clk [26618]));
Q_ASSIGN U6157 ( .B(clk), .A(\g.we_clk [26617]));
Q_ASSIGN U6158 ( .B(clk), .A(\g.we_clk [26616]));
Q_ASSIGN U6159 ( .B(clk), .A(\g.we_clk [26615]));
Q_ASSIGN U6160 ( .B(clk), .A(\g.we_clk [26614]));
Q_ASSIGN U6161 ( .B(clk), .A(\g.we_clk [26613]));
Q_ASSIGN U6162 ( .B(clk), .A(\g.we_clk [26612]));
Q_ASSIGN U6163 ( .B(clk), .A(\g.we_clk [26611]));
Q_ASSIGN U6164 ( .B(clk), .A(\g.we_clk [26610]));
Q_ASSIGN U6165 ( .B(clk), .A(\g.we_clk [26609]));
Q_ASSIGN U6166 ( .B(clk), .A(\g.we_clk [26608]));
Q_ASSIGN U6167 ( .B(clk), .A(\g.we_clk [26607]));
Q_ASSIGN U6168 ( .B(clk), .A(\g.we_clk [26606]));
Q_ASSIGN U6169 ( .B(clk), .A(\g.we_clk [26605]));
Q_ASSIGN U6170 ( .B(clk), .A(\g.we_clk [26604]));
Q_ASSIGN U6171 ( .B(clk), .A(\g.we_clk [26603]));
Q_ASSIGN U6172 ( .B(clk), .A(\g.we_clk [26602]));
Q_ASSIGN U6173 ( .B(clk), .A(\g.we_clk [26601]));
Q_ASSIGN U6174 ( .B(clk), .A(\g.we_clk [26600]));
Q_ASSIGN U6175 ( .B(clk), .A(\g.we_clk [26599]));
Q_ASSIGN U6176 ( .B(clk), .A(\g.we_clk [26598]));
Q_ASSIGN U6177 ( .B(clk), .A(\g.we_clk [26597]));
Q_ASSIGN U6178 ( .B(clk), .A(\g.we_clk [26596]));
Q_ASSIGN U6179 ( .B(clk), .A(\g.we_clk [26595]));
Q_ASSIGN U6180 ( .B(clk), .A(\g.we_clk [26594]));
Q_ASSIGN U6181 ( .B(clk), .A(\g.we_clk [26593]));
Q_ASSIGN U6182 ( .B(clk), .A(\g.we_clk [26592]));
Q_ASSIGN U6183 ( .B(clk), .A(\g.we_clk [26591]));
Q_ASSIGN U6184 ( .B(clk), .A(\g.we_clk [26590]));
Q_ASSIGN U6185 ( .B(clk), .A(\g.we_clk [26589]));
Q_ASSIGN U6186 ( .B(clk), .A(\g.we_clk [26588]));
Q_ASSIGN U6187 ( .B(clk), .A(\g.we_clk [26587]));
Q_ASSIGN U6188 ( .B(clk), .A(\g.we_clk [26586]));
Q_ASSIGN U6189 ( .B(clk), .A(\g.we_clk [26585]));
Q_ASSIGN U6190 ( .B(clk), .A(\g.we_clk [26584]));
Q_ASSIGN U6191 ( .B(clk), .A(\g.we_clk [26583]));
Q_ASSIGN U6192 ( .B(clk), .A(\g.we_clk [26582]));
Q_ASSIGN U6193 ( .B(clk), .A(\g.we_clk [26581]));
Q_ASSIGN U6194 ( .B(clk), .A(\g.we_clk [26580]));
Q_ASSIGN U6195 ( .B(clk), .A(\g.we_clk [26579]));
Q_ASSIGN U6196 ( .B(clk), .A(\g.we_clk [26578]));
Q_ASSIGN U6197 ( .B(clk), .A(\g.we_clk [26577]));
Q_ASSIGN U6198 ( .B(clk), .A(\g.we_clk [26576]));
Q_ASSIGN U6199 ( .B(clk), .A(\g.we_clk [26575]));
Q_ASSIGN U6200 ( .B(clk), .A(\g.we_clk [26574]));
Q_ASSIGN U6201 ( .B(clk), .A(\g.we_clk [26573]));
Q_ASSIGN U6202 ( .B(clk), .A(\g.we_clk [26572]));
Q_ASSIGN U6203 ( .B(clk), .A(\g.we_clk [26571]));
Q_ASSIGN U6204 ( .B(clk), .A(\g.we_clk [26570]));
Q_ASSIGN U6205 ( .B(clk), .A(\g.we_clk [26569]));
Q_ASSIGN U6206 ( .B(clk), .A(\g.we_clk [26568]));
Q_ASSIGN U6207 ( .B(clk), .A(\g.we_clk [26567]));
Q_ASSIGN U6208 ( .B(clk), .A(\g.we_clk [26566]));
Q_ASSIGN U6209 ( .B(clk), .A(\g.we_clk [26565]));
Q_ASSIGN U6210 ( .B(clk), .A(\g.we_clk [26564]));
Q_ASSIGN U6211 ( .B(clk), .A(\g.we_clk [26563]));
Q_ASSIGN U6212 ( .B(clk), .A(\g.we_clk [26562]));
Q_ASSIGN U6213 ( .B(clk), .A(\g.we_clk [26561]));
Q_ASSIGN U6214 ( .B(clk), .A(\g.we_clk [26560]));
Q_ASSIGN U6215 ( .B(clk), .A(\g.we_clk [26559]));
Q_ASSIGN U6216 ( .B(clk), .A(\g.we_clk [26558]));
Q_ASSIGN U6217 ( .B(clk), .A(\g.we_clk [26557]));
Q_ASSIGN U6218 ( .B(clk), .A(\g.we_clk [26556]));
Q_ASSIGN U6219 ( .B(clk), .A(\g.we_clk [26555]));
Q_ASSIGN U6220 ( .B(clk), .A(\g.we_clk [26554]));
Q_ASSIGN U6221 ( .B(clk), .A(\g.we_clk [26553]));
Q_ASSIGN U6222 ( .B(clk), .A(\g.we_clk [26552]));
Q_ASSIGN U6223 ( .B(clk), .A(\g.we_clk [26551]));
Q_ASSIGN U6224 ( .B(clk), .A(\g.we_clk [26550]));
Q_ASSIGN U6225 ( .B(clk), .A(\g.we_clk [26549]));
Q_ASSIGN U6226 ( .B(clk), .A(\g.we_clk [26548]));
Q_ASSIGN U6227 ( .B(clk), .A(\g.we_clk [26547]));
Q_ASSIGN U6228 ( .B(clk), .A(\g.we_clk [26546]));
Q_ASSIGN U6229 ( .B(clk), .A(\g.we_clk [26545]));
Q_ASSIGN U6230 ( .B(clk), .A(\g.we_clk [26544]));
Q_ASSIGN U6231 ( .B(clk), .A(\g.we_clk [26543]));
Q_ASSIGN U6232 ( .B(clk), .A(\g.we_clk [26542]));
Q_ASSIGN U6233 ( .B(clk), .A(\g.we_clk [26541]));
Q_ASSIGN U6234 ( .B(clk), .A(\g.we_clk [26540]));
Q_ASSIGN U6235 ( .B(clk), .A(\g.we_clk [26539]));
Q_ASSIGN U6236 ( .B(clk), .A(\g.we_clk [26538]));
Q_ASSIGN U6237 ( .B(clk), .A(\g.we_clk [26537]));
Q_ASSIGN U6238 ( .B(clk), .A(\g.we_clk [26536]));
Q_ASSIGN U6239 ( .B(clk), .A(\g.we_clk [26535]));
Q_ASSIGN U6240 ( .B(clk), .A(\g.we_clk [26534]));
Q_ASSIGN U6241 ( .B(clk), .A(\g.we_clk [26533]));
Q_ASSIGN U6242 ( .B(clk), .A(\g.we_clk [26532]));
Q_ASSIGN U6243 ( .B(clk), .A(\g.we_clk [26531]));
Q_ASSIGN U6244 ( .B(clk), .A(\g.we_clk [26530]));
Q_ASSIGN U6245 ( .B(clk), .A(\g.we_clk [26529]));
Q_ASSIGN U6246 ( .B(clk), .A(\g.we_clk [26528]));
Q_ASSIGN U6247 ( .B(clk), .A(\g.we_clk [26527]));
Q_ASSIGN U6248 ( .B(clk), .A(\g.we_clk [26526]));
Q_ASSIGN U6249 ( .B(clk), .A(\g.we_clk [26525]));
Q_ASSIGN U6250 ( .B(clk), .A(\g.we_clk [26524]));
Q_ASSIGN U6251 ( .B(clk), .A(\g.we_clk [26523]));
Q_ASSIGN U6252 ( .B(clk), .A(\g.we_clk [26522]));
Q_ASSIGN U6253 ( .B(clk), .A(\g.we_clk [26521]));
Q_ASSIGN U6254 ( .B(clk), .A(\g.we_clk [26520]));
Q_ASSIGN U6255 ( .B(clk), .A(\g.we_clk [26519]));
Q_ASSIGN U6256 ( .B(clk), .A(\g.we_clk [26518]));
Q_ASSIGN U6257 ( .B(clk), .A(\g.we_clk [26517]));
Q_ASSIGN U6258 ( .B(clk), .A(\g.we_clk [26516]));
Q_ASSIGN U6259 ( .B(clk), .A(\g.we_clk [26515]));
Q_ASSIGN U6260 ( .B(clk), .A(\g.we_clk [26514]));
Q_ASSIGN U6261 ( .B(clk), .A(\g.we_clk [26513]));
Q_ASSIGN U6262 ( .B(clk), .A(\g.we_clk [26512]));
Q_ASSIGN U6263 ( .B(clk), .A(\g.we_clk [26511]));
Q_ASSIGN U6264 ( .B(clk), .A(\g.we_clk [26510]));
Q_ASSIGN U6265 ( .B(clk), .A(\g.we_clk [26509]));
Q_ASSIGN U6266 ( .B(clk), .A(\g.we_clk [26508]));
Q_ASSIGN U6267 ( .B(clk), .A(\g.we_clk [26507]));
Q_ASSIGN U6268 ( .B(clk), .A(\g.we_clk [26506]));
Q_ASSIGN U6269 ( .B(clk), .A(\g.we_clk [26505]));
Q_ASSIGN U6270 ( .B(clk), .A(\g.we_clk [26504]));
Q_ASSIGN U6271 ( .B(clk), .A(\g.we_clk [26503]));
Q_ASSIGN U6272 ( .B(clk), .A(\g.we_clk [26502]));
Q_ASSIGN U6273 ( .B(clk), .A(\g.we_clk [26501]));
Q_ASSIGN U6274 ( .B(clk), .A(\g.we_clk [26500]));
Q_ASSIGN U6275 ( .B(clk), .A(\g.we_clk [26499]));
Q_ASSIGN U6276 ( .B(clk), .A(\g.we_clk [26498]));
Q_ASSIGN U6277 ( .B(clk), .A(\g.we_clk [26497]));
Q_ASSIGN U6278 ( .B(clk), .A(\g.we_clk [26496]));
Q_ASSIGN U6279 ( .B(clk), .A(\g.we_clk [26495]));
Q_ASSIGN U6280 ( .B(clk), .A(\g.we_clk [26494]));
Q_ASSIGN U6281 ( .B(clk), .A(\g.we_clk [26493]));
Q_ASSIGN U6282 ( .B(clk), .A(\g.we_clk [26492]));
Q_ASSIGN U6283 ( .B(clk), .A(\g.we_clk [26491]));
Q_ASSIGN U6284 ( .B(clk), .A(\g.we_clk [26490]));
Q_ASSIGN U6285 ( .B(clk), .A(\g.we_clk [26489]));
Q_ASSIGN U6286 ( .B(clk), .A(\g.we_clk [26488]));
Q_ASSIGN U6287 ( .B(clk), .A(\g.we_clk [26487]));
Q_ASSIGN U6288 ( .B(clk), .A(\g.we_clk [26486]));
Q_ASSIGN U6289 ( .B(clk), .A(\g.we_clk [26485]));
Q_ASSIGN U6290 ( .B(clk), .A(\g.we_clk [26484]));
Q_ASSIGN U6291 ( .B(clk), .A(\g.we_clk [26483]));
Q_ASSIGN U6292 ( .B(clk), .A(\g.we_clk [26482]));
Q_ASSIGN U6293 ( .B(clk), .A(\g.we_clk [26481]));
Q_ASSIGN U6294 ( .B(clk), .A(\g.we_clk [26480]));
Q_ASSIGN U6295 ( .B(clk), .A(\g.we_clk [26479]));
Q_ASSIGN U6296 ( .B(clk), .A(\g.we_clk [26478]));
Q_ASSIGN U6297 ( .B(clk), .A(\g.we_clk [26477]));
Q_ASSIGN U6298 ( .B(clk), .A(\g.we_clk [26476]));
Q_ASSIGN U6299 ( .B(clk), .A(\g.we_clk [26475]));
Q_ASSIGN U6300 ( .B(clk), .A(\g.we_clk [26474]));
Q_ASSIGN U6301 ( .B(clk), .A(\g.we_clk [26473]));
Q_ASSIGN U6302 ( .B(clk), .A(\g.we_clk [26472]));
Q_ASSIGN U6303 ( .B(clk), .A(\g.we_clk [26471]));
Q_ASSIGN U6304 ( .B(clk), .A(\g.we_clk [26470]));
Q_ASSIGN U6305 ( .B(clk), .A(\g.we_clk [26469]));
Q_ASSIGN U6306 ( .B(clk), .A(\g.we_clk [26468]));
Q_ASSIGN U6307 ( .B(clk), .A(\g.we_clk [26467]));
Q_ASSIGN U6308 ( .B(clk), .A(\g.we_clk [26466]));
Q_ASSIGN U6309 ( .B(clk), .A(\g.we_clk [26465]));
Q_ASSIGN U6310 ( .B(clk), .A(\g.we_clk [26464]));
Q_ASSIGN U6311 ( .B(clk), .A(\g.we_clk [26463]));
Q_ASSIGN U6312 ( .B(clk), .A(\g.we_clk [26462]));
Q_ASSIGN U6313 ( .B(clk), .A(\g.we_clk [26461]));
Q_ASSIGN U6314 ( .B(clk), .A(\g.we_clk [26460]));
Q_ASSIGN U6315 ( .B(clk), .A(\g.we_clk [26459]));
Q_ASSIGN U6316 ( .B(clk), .A(\g.we_clk [26458]));
Q_ASSIGN U6317 ( .B(clk), .A(\g.we_clk [26457]));
Q_ASSIGN U6318 ( .B(clk), .A(\g.we_clk [26456]));
Q_ASSIGN U6319 ( .B(clk), .A(\g.we_clk [26455]));
Q_ASSIGN U6320 ( .B(clk), .A(\g.we_clk [26454]));
Q_ASSIGN U6321 ( .B(clk), .A(\g.we_clk [26453]));
Q_ASSIGN U6322 ( .B(clk), .A(\g.we_clk [26452]));
Q_ASSIGN U6323 ( .B(clk), .A(\g.we_clk [26451]));
Q_ASSIGN U6324 ( .B(clk), .A(\g.we_clk [26450]));
Q_ASSIGN U6325 ( .B(clk), .A(\g.we_clk [26449]));
Q_ASSIGN U6326 ( .B(clk), .A(\g.we_clk [26448]));
Q_ASSIGN U6327 ( .B(clk), .A(\g.we_clk [26447]));
Q_ASSIGN U6328 ( .B(clk), .A(\g.we_clk [26446]));
Q_ASSIGN U6329 ( .B(clk), .A(\g.we_clk [26445]));
Q_ASSIGN U6330 ( .B(clk), .A(\g.we_clk [26444]));
Q_ASSIGN U6331 ( .B(clk), .A(\g.we_clk [26443]));
Q_ASSIGN U6332 ( .B(clk), .A(\g.we_clk [26442]));
Q_ASSIGN U6333 ( .B(clk), .A(\g.we_clk [26441]));
Q_ASSIGN U6334 ( .B(clk), .A(\g.we_clk [26440]));
Q_ASSIGN U6335 ( .B(clk), .A(\g.we_clk [26439]));
Q_ASSIGN U6336 ( .B(clk), .A(\g.we_clk [26438]));
Q_ASSIGN U6337 ( .B(clk), .A(\g.we_clk [26437]));
Q_ASSIGN U6338 ( .B(clk), .A(\g.we_clk [26436]));
Q_ASSIGN U6339 ( .B(clk), .A(\g.we_clk [26435]));
Q_ASSIGN U6340 ( .B(clk), .A(\g.we_clk [26434]));
Q_ASSIGN U6341 ( .B(clk), .A(\g.we_clk [26433]));
Q_ASSIGN U6342 ( .B(clk), .A(\g.we_clk [26432]));
Q_ASSIGN U6343 ( .B(clk), .A(\g.we_clk [26431]));
Q_ASSIGN U6344 ( .B(clk), .A(\g.we_clk [26430]));
Q_ASSIGN U6345 ( .B(clk), .A(\g.we_clk [26429]));
Q_ASSIGN U6346 ( .B(clk), .A(\g.we_clk [26428]));
Q_ASSIGN U6347 ( .B(clk), .A(\g.we_clk [26427]));
Q_ASSIGN U6348 ( .B(clk), .A(\g.we_clk [26426]));
Q_ASSIGN U6349 ( .B(clk), .A(\g.we_clk [26425]));
Q_ASSIGN U6350 ( .B(clk), .A(\g.we_clk [26424]));
Q_ASSIGN U6351 ( .B(clk), .A(\g.we_clk [26423]));
Q_ASSIGN U6352 ( .B(clk), .A(\g.we_clk [26422]));
Q_ASSIGN U6353 ( .B(clk), .A(\g.we_clk [26421]));
Q_ASSIGN U6354 ( .B(clk), .A(\g.we_clk [26420]));
Q_ASSIGN U6355 ( .B(clk), .A(\g.we_clk [26419]));
Q_ASSIGN U6356 ( .B(clk), .A(\g.we_clk [26418]));
Q_ASSIGN U6357 ( .B(clk), .A(\g.we_clk [26417]));
Q_ASSIGN U6358 ( .B(clk), .A(\g.we_clk [26416]));
Q_ASSIGN U6359 ( .B(clk), .A(\g.we_clk [26415]));
Q_ASSIGN U6360 ( .B(clk), .A(\g.we_clk [26414]));
Q_ASSIGN U6361 ( .B(clk), .A(\g.we_clk [26413]));
Q_ASSIGN U6362 ( .B(clk), .A(\g.we_clk [26412]));
Q_ASSIGN U6363 ( .B(clk), .A(\g.we_clk [26411]));
Q_ASSIGN U6364 ( .B(clk), .A(\g.we_clk [26410]));
Q_ASSIGN U6365 ( .B(clk), .A(\g.we_clk [26409]));
Q_ASSIGN U6366 ( .B(clk), .A(\g.we_clk [26408]));
Q_ASSIGN U6367 ( .B(clk), .A(\g.we_clk [26407]));
Q_ASSIGN U6368 ( .B(clk), .A(\g.we_clk [26406]));
Q_ASSIGN U6369 ( .B(clk), .A(\g.we_clk [26405]));
Q_ASSIGN U6370 ( .B(clk), .A(\g.we_clk [26404]));
Q_ASSIGN U6371 ( .B(clk), .A(\g.we_clk [26403]));
Q_ASSIGN U6372 ( .B(clk), .A(\g.we_clk [26402]));
Q_ASSIGN U6373 ( .B(clk), .A(\g.we_clk [26401]));
Q_ASSIGN U6374 ( .B(clk), .A(\g.we_clk [26400]));
Q_ASSIGN U6375 ( .B(clk), .A(\g.we_clk [26399]));
Q_ASSIGN U6376 ( .B(clk), .A(\g.we_clk [26398]));
Q_ASSIGN U6377 ( .B(clk), .A(\g.we_clk [26397]));
Q_ASSIGN U6378 ( .B(clk), .A(\g.we_clk [26396]));
Q_ASSIGN U6379 ( .B(clk), .A(\g.we_clk [26395]));
Q_ASSIGN U6380 ( .B(clk), .A(\g.we_clk [26394]));
Q_ASSIGN U6381 ( .B(clk), .A(\g.we_clk [26393]));
Q_ASSIGN U6382 ( .B(clk), .A(\g.we_clk [26392]));
Q_ASSIGN U6383 ( .B(clk), .A(\g.we_clk [26391]));
Q_ASSIGN U6384 ( .B(clk), .A(\g.we_clk [26390]));
Q_ASSIGN U6385 ( .B(clk), .A(\g.we_clk [26389]));
Q_ASSIGN U6386 ( .B(clk), .A(\g.we_clk [26388]));
Q_ASSIGN U6387 ( .B(clk), .A(\g.we_clk [26387]));
Q_ASSIGN U6388 ( .B(clk), .A(\g.we_clk [26386]));
Q_ASSIGN U6389 ( .B(clk), .A(\g.we_clk [26385]));
Q_ASSIGN U6390 ( .B(clk), .A(\g.we_clk [26384]));
Q_ASSIGN U6391 ( .B(clk), .A(\g.we_clk [26383]));
Q_ASSIGN U6392 ( .B(clk), .A(\g.we_clk [26382]));
Q_ASSIGN U6393 ( .B(clk), .A(\g.we_clk [26381]));
Q_ASSIGN U6394 ( .B(clk), .A(\g.we_clk [26380]));
Q_ASSIGN U6395 ( .B(clk), .A(\g.we_clk [26379]));
Q_ASSIGN U6396 ( .B(clk), .A(\g.we_clk [26378]));
Q_ASSIGN U6397 ( .B(clk), .A(\g.we_clk [26377]));
Q_ASSIGN U6398 ( .B(clk), .A(\g.we_clk [26376]));
Q_ASSIGN U6399 ( .B(clk), .A(\g.we_clk [26375]));
Q_ASSIGN U6400 ( .B(clk), .A(\g.we_clk [26374]));
Q_ASSIGN U6401 ( .B(clk), .A(\g.we_clk [26373]));
Q_ASSIGN U6402 ( .B(clk), .A(\g.we_clk [26372]));
Q_ASSIGN U6403 ( .B(clk), .A(\g.we_clk [26371]));
Q_ASSIGN U6404 ( .B(clk), .A(\g.we_clk [26370]));
Q_ASSIGN U6405 ( .B(clk), .A(\g.we_clk [26369]));
Q_ASSIGN U6406 ( .B(clk), .A(\g.we_clk [26368]));
Q_ASSIGN U6407 ( .B(clk), .A(\g.we_clk [26367]));
Q_ASSIGN U6408 ( .B(clk), .A(\g.we_clk [26366]));
Q_ASSIGN U6409 ( .B(clk), .A(\g.we_clk [26365]));
Q_ASSIGN U6410 ( .B(clk), .A(\g.we_clk [26364]));
Q_ASSIGN U6411 ( .B(clk), .A(\g.we_clk [26363]));
Q_ASSIGN U6412 ( .B(clk), .A(\g.we_clk [26362]));
Q_ASSIGN U6413 ( .B(clk), .A(\g.we_clk [26361]));
Q_ASSIGN U6414 ( .B(clk), .A(\g.we_clk [26360]));
Q_ASSIGN U6415 ( .B(clk), .A(\g.we_clk [26359]));
Q_ASSIGN U6416 ( .B(clk), .A(\g.we_clk [26358]));
Q_ASSIGN U6417 ( .B(clk), .A(\g.we_clk [26357]));
Q_ASSIGN U6418 ( .B(clk), .A(\g.we_clk [26356]));
Q_ASSIGN U6419 ( .B(clk), .A(\g.we_clk [26355]));
Q_ASSIGN U6420 ( .B(clk), .A(\g.we_clk [26354]));
Q_ASSIGN U6421 ( .B(clk), .A(\g.we_clk [26353]));
Q_ASSIGN U6422 ( .B(clk), .A(\g.we_clk [26352]));
Q_ASSIGN U6423 ( .B(clk), .A(\g.we_clk [26351]));
Q_ASSIGN U6424 ( .B(clk), .A(\g.we_clk [26350]));
Q_ASSIGN U6425 ( .B(clk), .A(\g.we_clk [26349]));
Q_ASSIGN U6426 ( .B(clk), .A(\g.we_clk [26348]));
Q_ASSIGN U6427 ( .B(clk), .A(\g.we_clk [26347]));
Q_ASSIGN U6428 ( .B(clk), .A(\g.we_clk [26346]));
Q_ASSIGN U6429 ( .B(clk), .A(\g.we_clk [26345]));
Q_ASSIGN U6430 ( .B(clk), .A(\g.we_clk [26344]));
Q_ASSIGN U6431 ( .B(clk), .A(\g.we_clk [26343]));
Q_ASSIGN U6432 ( .B(clk), .A(\g.we_clk [26342]));
Q_ASSIGN U6433 ( .B(clk), .A(\g.we_clk [26341]));
Q_ASSIGN U6434 ( .B(clk), .A(\g.we_clk [26340]));
Q_ASSIGN U6435 ( .B(clk), .A(\g.we_clk [26339]));
Q_ASSIGN U6436 ( .B(clk), .A(\g.we_clk [26338]));
Q_ASSIGN U6437 ( .B(clk), .A(\g.we_clk [26337]));
Q_ASSIGN U6438 ( .B(clk), .A(\g.we_clk [26336]));
Q_ASSIGN U6439 ( .B(clk), .A(\g.we_clk [26335]));
Q_ASSIGN U6440 ( .B(clk), .A(\g.we_clk [26334]));
Q_ASSIGN U6441 ( .B(clk), .A(\g.we_clk [26333]));
Q_ASSIGN U6442 ( .B(clk), .A(\g.we_clk [26332]));
Q_ASSIGN U6443 ( .B(clk), .A(\g.we_clk [26331]));
Q_ASSIGN U6444 ( .B(clk), .A(\g.we_clk [26330]));
Q_ASSIGN U6445 ( .B(clk), .A(\g.we_clk [26329]));
Q_ASSIGN U6446 ( .B(clk), .A(\g.we_clk [26328]));
Q_ASSIGN U6447 ( .B(clk), .A(\g.we_clk [26327]));
Q_ASSIGN U6448 ( .B(clk), .A(\g.we_clk [26326]));
Q_ASSIGN U6449 ( .B(clk), .A(\g.we_clk [26325]));
Q_ASSIGN U6450 ( .B(clk), .A(\g.we_clk [26324]));
Q_ASSIGN U6451 ( .B(clk), .A(\g.we_clk [26323]));
Q_ASSIGN U6452 ( .B(clk), .A(\g.we_clk [26322]));
Q_ASSIGN U6453 ( .B(clk), .A(\g.we_clk [26321]));
Q_ASSIGN U6454 ( .B(clk), .A(\g.we_clk [26320]));
Q_ASSIGN U6455 ( .B(clk), .A(\g.we_clk [26319]));
Q_ASSIGN U6456 ( .B(clk), .A(\g.we_clk [26318]));
Q_ASSIGN U6457 ( .B(clk), .A(\g.we_clk [26317]));
Q_ASSIGN U6458 ( .B(clk), .A(\g.we_clk [26316]));
Q_ASSIGN U6459 ( .B(clk), .A(\g.we_clk [26315]));
Q_ASSIGN U6460 ( .B(clk), .A(\g.we_clk [26314]));
Q_ASSIGN U6461 ( .B(clk), .A(\g.we_clk [26313]));
Q_ASSIGN U6462 ( .B(clk), .A(\g.we_clk [26312]));
Q_ASSIGN U6463 ( .B(clk), .A(\g.we_clk [26311]));
Q_ASSIGN U6464 ( .B(clk), .A(\g.we_clk [26310]));
Q_ASSIGN U6465 ( .B(clk), .A(\g.we_clk [26309]));
Q_ASSIGN U6466 ( .B(clk), .A(\g.we_clk [26308]));
Q_ASSIGN U6467 ( .B(clk), .A(\g.we_clk [26307]));
Q_ASSIGN U6468 ( .B(clk), .A(\g.we_clk [26306]));
Q_ASSIGN U6469 ( .B(clk), .A(\g.we_clk [26305]));
Q_ASSIGN U6470 ( .B(clk), .A(\g.we_clk [26304]));
Q_ASSIGN U6471 ( .B(clk), .A(\g.we_clk [26303]));
Q_ASSIGN U6472 ( .B(clk), .A(\g.we_clk [26302]));
Q_ASSIGN U6473 ( .B(clk), .A(\g.we_clk [26301]));
Q_ASSIGN U6474 ( .B(clk), .A(\g.we_clk [26300]));
Q_ASSIGN U6475 ( .B(clk), .A(\g.we_clk [26299]));
Q_ASSIGN U6476 ( .B(clk), .A(\g.we_clk [26298]));
Q_ASSIGN U6477 ( .B(clk), .A(\g.we_clk [26297]));
Q_ASSIGN U6478 ( .B(clk), .A(\g.we_clk [26296]));
Q_ASSIGN U6479 ( .B(clk), .A(\g.we_clk [26295]));
Q_ASSIGN U6480 ( .B(clk), .A(\g.we_clk [26294]));
Q_ASSIGN U6481 ( .B(clk), .A(\g.we_clk [26293]));
Q_ASSIGN U6482 ( .B(clk), .A(\g.we_clk [26292]));
Q_ASSIGN U6483 ( .B(clk), .A(\g.we_clk [26291]));
Q_ASSIGN U6484 ( .B(clk), .A(\g.we_clk [26290]));
Q_ASSIGN U6485 ( .B(clk), .A(\g.we_clk [26289]));
Q_ASSIGN U6486 ( .B(clk), .A(\g.we_clk [26288]));
Q_ASSIGN U6487 ( .B(clk), .A(\g.we_clk [26287]));
Q_ASSIGN U6488 ( .B(clk), .A(\g.we_clk [26286]));
Q_ASSIGN U6489 ( .B(clk), .A(\g.we_clk [26285]));
Q_ASSIGN U6490 ( .B(clk), .A(\g.we_clk [26284]));
Q_ASSIGN U6491 ( .B(clk), .A(\g.we_clk [26283]));
Q_ASSIGN U6492 ( .B(clk), .A(\g.we_clk [26282]));
Q_ASSIGN U6493 ( .B(clk), .A(\g.we_clk [26281]));
Q_ASSIGN U6494 ( .B(clk), .A(\g.we_clk [26280]));
Q_ASSIGN U6495 ( .B(clk), .A(\g.we_clk [26279]));
Q_ASSIGN U6496 ( .B(clk), .A(\g.we_clk [26278]));
Q_ASSIGN U6497 ( .B(clk), .A(\g.we_clk [26277]));
Q_ASSIGN U6498 ( .B(clk), .A(\g.we_clk [26276]));
Q_ASSIGN U6499 ( .B(clk), .A(\g.we_clk [26275]));
Q_ASSIGN U6500 ( .B(clk), .A(\g.we_clk [26274]));
Q_ASSIGN U6501 ( .B(clk), .A(\g.we_clk [26273]));
Q_ASSIGN U6502 ( .B(clk), .A(\g.we_clk [26272]));
Q_ASSIGN U6503 ( .B(clk), .A(\g.we_clk [26271]));
Q_ASSIGN U6504 ( .B(clk), .A(\g.we_clk [26270]));
Q_ASSIGN U6505 ( .B(clk), .A(\g.we_clk [26269]));
Q_ASSIGN U6506 ( .B(clk), .A(\g.we_clk [26268]));
Q_ASSIGN U6507 ( .B(clk), .A(\g.we_clk [26267]));
Q_ASSIGN U6508 ( .B(clk), .A(\g.we_clk [26266]));
Q_ASSIGN U6509 ( .B(clk), .A(\g.we_clk [26265]));
Q_ASSIGN U6510 ( .B(clk), .A(\g.we_clk [26264]));
Q_ASSIGN U6511 ( .B(clk), .A(\g.we_clk [26263]));
Q_ASSIGN U6512 ( .B(clk), .A(\g.we_clk [26262]));
Q_ASSIGN U6513 ( .B(clk), .A(\g.we_clk [26261]));
Q_ASSIGN U6514 ( .B(clk), .A(\g.we_clk [26260]));
Q_ASSIGN U6515 ( .B(clk), .A(\g.we_clk [26259]));
Q_ASSIGN U6516 ( .B(clk), .A(\g.we_clk [26258]));
Q_ASSIGN U6517 ( .B(clk), .A(\g.we_clk [26257]));
Q_ASSIGN U6518 ( .B(clk), .A(\g.we_clk [26256]));
Q_ASSIGN U6519 ( .B(clk), .A(\g.we_clk [26255]));
Q_ASSIGN U6520 ( .B(clk), .A(\g.we_clk [26254]));
Q_ASSIGN U6521 ( .B(clk), .A(\g.we_clk [26253]));
Q_ASSIGN U6522 ( .B(clk), .A(\g.we_clk [26252]));
Q_ASSIGN U6523 ( .B(clk), .A(\g.we_clk [26251]));
Q_ASSIGN U6524 ( .B(clk), .A(\g.we_clk [26250]));
Q_ASSIGN U6525 ( .B(clk), .A(\g.we_clk [26249]));
Q_ASSIGN U6526 ( .B(clk), .A(\g.we_clk [26248]));
Q_ASSIGN U6527 ( .B(clk), .A(\g.we_clk [26247]));
Q_ASSIGN U6528 ( .B(clk), .A(\g.we_clk [26246]));
Q_ASSIGN U6529 ( .B(clk), .A(\g.we_clk [26245]));
Q_ASSIGN U6530 ( .B(clk), .A(\g.we_clk [26244]));
Q_ASSIGN U6531 ( .B(clk), .A(\g.we_clk [26243]));
Q_ASSIGN U6532 ( .B(clk), .A(\g.we_clk [26242]));
Q_ASSIGN U6533 ( .B(clk), .A(\g.we_clk [26241]));
Q_ASSIGN U6534 ( .B(clk), .A(\g.we_clk [26240]));
Q_ASSIGN U6535 ( .B(clk), .A(\g.we_clk [26239]));
Q_ASSIGN U6536 ( .B(clk), .A(\g.we_clk [26238]));
Q_ASSIGN U6537 ( .B(clk), .A(\g.we_clk [26237]));
Q_ASSIGN U6538 ( .B(clk), .A(\g.we_clk [26236]));
Q_ASSIGN U6539 ( .B(clk), .A(\g.we_clk [26235]));
Q_ASSIGN U6540 ( .B(clk), .A(\g.we_clk [26234]));
Q_ASSIGN U6541 ( .B(clk), .A(\g.we_clk [26233]));
Q_ASSIGN U6542 ( .B(clk), .A(\g.we_clk [26232]));
Q_ASSIGN U6543 ( .B(clk), .A(\g.we_clk [26231]));
Q_ASSIGN U6544 ( .B(clk), .A(\g.we_clk [26230]));
Q_ASSIGN U6545 ( .B(clk), .A(\g.we_clk [26229]));
Q_ASSIGN U6546 ( .B(clk), .A(\g.we_clk [26228]));
Q_ASSIGN U6547 ( .B(clk), .A(\g.we_clk [26227]));
Q_ASSIGN U6548 ( .B(clk), .A(\g.we_clk [26226]));
Q_ASSIGN U6549 ( .B(clk), .A(\g.we_clk [26225]));
Q_ASSIGN U6550 ( .B(clk), .A(\g.we_clk [26224]));
Q_ASSIGN U6551 ( .B(clk), .A(\g.we_clk [26223]));
Q_ASSIGN U6552 ( .B(clk), .A(\g.we_clk [26222]));
Q_ASSIGN U6553 ( .B(clk), .A(\g.we_clk [26221]));
Q_ASSIGN U6554 ( .B(clk), .A(\g.we_clk [26220]));
Q_ASSIGN U6555 ( .B(clk), .A(\g.we_clk [26219]));
Q_ASSIGN U6556 ( .B(clk), .A(\g.we_clk [26218]));
Q_ASSIGN U6557 ( .B(clk), .A(\g.we_clk [26217]));
Q_ASSIGN U6558 ( .B(clk), .A(\g.we_clk [26216]));
Q_ASSIGN U6559 ( .B(clk), .A(\g.we_clk [26215]));
Q_ASSIGN U6560 ( .B(clk), .A(\g.we_clk [26214]));
Q_ASSIGN U6561 ( .B(clk), .A(\g.we_clk [26213]));
Q_ASSIGN U6562 ( .B(clk), .A(\g.we_clk [26212]));
Q_ASSIGN U6563 ( .B(clk), .A(\g.we_clk [26211]));
Q_ASSIGN U6564 ( .B(clk), .A(\g.we_clk [26210]));
Q_ASSIGN U6565 ( .B(clk), .A(\g.we_clk [26209]));
Q_ASSIGN U6566 ( .B(clk), .A(\g.we_clk [26208]));
Q_ASSIGN U6567 ( .B(clk), .A(\g.we_clk [26207]));
Q_ASSIGN U6568 ( .B(clk), .A(\g.we_clk [26206]));
Q_ASSIGN U6569 ( .B(clk), .A(\g.we_clk [26205]));
Q_ASSIGN U6570 ( .B(clk), .A(\g.we_clk [26204]));
Q_ASSIGN U6571 ( .B(clk), .A(\g.we_clk [26203]));
Q_ASSIGN U6572 ( .B(clk), .A(\g.we_clk [26202]));
Q_ASSIGN U6573 ( .B(clk), .A(\g.we_clk [26201]));
Q_ASSIGN U6574 ( .B(clk), .A(\g.we_clk [26200]));
Q_ASSIGN U6575 ( .B(clk), .A(\g.we_clk [26199]));
Q_ASSIGN U6576 ( .B(clk), .A(\g.we_clk [26198]));
Q_ASSIGN U6577 ( .B(clk), .A(\g.we_clk [26197]));
Q_ASSIGN U6578 ( .B(clk), .A(\g.we_clk [26196]));
Q_ASSIGN U6579 ( .B(clk), .A(\g.we_clk [26195]));
Q_ASSIGN U6580 ( .B(clk), .A(\g.we_clk [26194]));
Q_ASSIGN U6581 ( .B(clk), .A(\g.we_clk [26193]));
Q_ASSIGN U6582 ( .B(clk), .A(\g.we_clk [26192]));
Q_ASSIGN U6583 ( .B(clk), .A(\g.we_clk [26191]));
Q_ASSIGN U6584 ( .B(clk), .A(\g.we_clk [26190]));
Q_ASSIGN U6585 ( .B(clk), .A(\g.we_clk [26189]));
Q_ASSIGN U6586 ( .B(clk), .A(\g.we_clk [26188]));
Q_ASSIGN U6587 ( .B(clk), .A(\g.we_clk [26187]));
Q_ASSIGN U6588 ( .B(clk), .A(\g.we_clk [26186]));
Q_ASSIGN U6589 ( .B(clk), .A(\g.we_clk [26185]));
Q_ASSIGN U6590 ( .B(clk), .A(\g.we_clk [26184]));
Q_ASSIGN U6591 ( .B(clk), .A(\g.we_clk [26183]));
Q_ASSIGN U6592 ( .B(clk), .A(\g.we_clk [26182]));
Q_ASSIGN U6593 ( .B(clk), .A(\g.we_clk [26181]));
Q_ASSIGN U6594 ( .B(clk), .A(\g.we_clk [26180]));
Q_ASSIGN U6595 ( .B(clk), .A(\g.we_clk [26179]));
Q_ASSIGN U6596 ( .B(clk), .A(\g.we_clk [26178]));
Q_ASSIGN U6597 ( .B(clk), .A(\g.we_clk [26177]));
Q_ASSIGN U6598 ( .B(clk), .A(\g.we_clk [26176]));
Q_ASSIGN U6599 ( .B(clk), .A(\g.we_clk [26175]));
Q_ASSIGN U6600 ( .B(clk), .A(\g.we_clk [26174]));
Q_ASSIGN U6601 ( .B(clk), .A(\g.we_clk [26173]));
Q_ASSIGN U6602 ( .B(clk), .A(\g.we_clk [26172]));
Q_ASSIGN U6603 ( .B(clk), .A(\g.we_clk [26171]));
Q_ASSIGN U6604 ( .B(clk), .A(\g.we_clk [26170]));
Q_ASSIGN U6605 ( .B(clk), .A(\g.we_clk [26169]));
Q_ASSIGN U6606 ( .B(clk), .A(\g.we_clk [26168]));
Q_ASSIGN U6607 ( .B(clk), .A(\g.we_clk [26167]));
Q_ASSIGN U6608 ( .B(clk), .A(\g.we_clk [26166]));
Q_ASSIGN U6609 ( .B(clk), .A(\g.we_clk [26165]));
Q_ASSIGN U6610 ( .B(clk), .A(\g.we_clk [26164]));
Q_ASSIGN U6611 ( .B(clk), .A(\g.we_clk [26163]));
Q_ASSIGN U6612 ( .B(clk), .A(\g.we_clk [26162]));
Q_ASSIGN U6613 ( .B(clk), .A(\g.we_clk [26161]));
Q_ASSIGN U6614 ( .B(clk), .A(\g.we_clk [26160]));
Q_ASSIGN U6615 ( .B(clk), .A(\g.we_clk [26159]));
Q_ASSIGN U6616 ( .B(clk), .A(\g.we_clk [26158]));
Q_ASSIGN U6617 ( .B(clk), .A(\g.we_clk [26157]));
Q_ASSIGN U6618 ( .B(clk), .A(\g.we_clk [26156]));
Q_ASSIGN U6619 ( .B(clk), .A(\g.we_clk [26155]));
Q_ASSIGN U6620 ( .B(clk), .A(\g.we_clk [26154]));
Q_ASSIGN U6621 ( .B(clk), .A(\g.we_clk [26153]));
Q_ASSIGN U6622 ( .B(clk), .A(\g.we_clk [26152]));
Q_ASSIGN U6623 ( .B(clk), .A(\g.we_clk [26151]));
Q_ASSIGN U6624 ( .B(clk), .A(\g.we_clk [26150]));
Q_ASSIGN U6625 ( .B(clk), .A(\g.we_clk [26149]));
Q_ASSIGN U6626 ( .B(clk), .A(\g.we_clk [26148]));
Q_ASSIGN U6627 ( .B(clk), .A(\g.we_clk [26147]));
Q_ASSIGN U6628 ( .B(clk), .A(\g.we_clk [26146]));
Q_ASSIGN U6629 ( .B(clk), .A(\g.we_clk [26145]));
Q_ASSIGN U6630 ( .B(clk), .A(\g.we_clk [26144]));
Q_ASSIGN U6631 ( .B(clk), .A(\g.we_clk [26143]));
Q_ASSIGN U6632 ( .B(clk), .A(\g.we_clk [26142]));
Q_ASSIGN U6633 ( .B(clk), .A(\g.we_clk [26141]));
Q_ASSIGN U6634 ( .B(clk), .A(\g.we_clk [26140]));
Q_ASSIGN U6635 ( .B(clk), .A(\g.we_clk [26139]));
Q_ASSIGN U6636 ( .B(clk), .A(\g.we_clk [26138]));
Q_ASSIGN U6637 ( .B(clk), .A(\g.we_clk [26137]));
Q_ASSIGN U6638 ( .B(clk), .A(\g.we_clk [26136]));
Q_ASSIGN U6639 ( .B(clk), .A(\g.we_clk [26135]));
Q_ASSIGN U6640 ( .B(clk), .A(\g.we_clk [26134]));
Q_ASSIGN U6641 ( .B(clk), .A(\g.we_clk [26133]));
Q_ASSIGN U6642 ( .B(clk), .A(\g.we_clk [26132]));
Q_ASSIGN U6643 ( .B(clk), .A(\g.we_clk [26131]));
Q_ASSIGN U6644 ( .B(clk), .A(\g.we_clk [26130]));
Q_ASSIGN U6645 ( .B(clk), .A(\g.we_clk [26129]));
Q_ASSIGN U6646 ( .B(clk), .A(\g.we_clk [26128]));
Q_ASSIGN U6647 ( .B(clk), .A(\g.we_clk [26127]));
Q_ASSIGN U6648 ( .B(clk), .A(\g.we_clk [26126]));
Q_ASSIGN U6649 ( .B(clk), .A(\g.we_clk [26125]));
Q_ASSIGN U6650 ( .B(clk), .A(\g.we_clk [26124]));
Q_ASSIGN U6651 ( .B(clk), .A(\g.we_clk [26123]));
Q_ASSIGN U6652 ( .B(clk), .A(\g.we_clk [26122]));
Q_ASSIGN U6653 ( .B(clk), .A(\g.we_clk [26121]));
Q_ASSIGN U6654 ( .B(clk), .A(\g.we_clk [26120]));
Q_ASSIGN U6655 ( .B(clk), .A(\g.we_clk [26119]));
Q_ASSIGN U6656 ( .B(clk), .A(\g.we_clk [26118]));
Q_ASSIGN U6657 ( .B(clk), .A(\g.we_clk [26117]));
Q_ASSIGN U6658 ( .B(clk), .A(\g.we_clk [26116]));
Q_ASSIGN U6659 ( .B(clk), .A(\g.we_clk [26115]));
Q_ASSIGN U6660 ( .B(clk), .A(\g.we_clk [26114]));
Q_ASSIGN U6661 ( .B(clk), .A(\g.we_clk [26113]));
Q_ASSIGN U6662 ( .B(clk), .A(\g.we_clk [26112]));
Q_ASSIGN U6663 ( .B(clk), .A(\g.we_clk [26111]));
Q_ASSIGN U6664 ( .B(clk), .A(\g.we_clk [26110]));
Q_ASSIGN U6665 ( .B(clk), .A(\g.we_clk [26109]));
Q_ASSIGN U6666 ( .B(clk), .A(\g.we_clk [26108]));
Q_ASSIGN U6667 ( .B(clk), .A(\g.we_clk [26107]));
Q_ASSIGN U6668 ( .B(clk), .A(\g.we_clk [26106]));
Q_ASSIGN U6669 ( .B(clk), .A(\g.we_clk [26105]));
Q_ASSIGN U6670 ( .B(clk), .A(\g.we_clk [26104]));
Q_ASSIGN U6671 ( .B(clk), .A(\g.we_clk [26103]));
Q_ASSIGN U6672 ( .B(clk), .A(\g.we_clk [26102]));
Q_ASSIGN U6673 ( .B(clk), .A(\g.we_clk [26101]));
Q_ASSIGN U6674 ( .B(clk), .A(\g.we_clk [26100]));
Q_ASSIGN U6675 ( .B(clk), .A(\g.we_clk [26099]));
Q_ASSIGN U6676 ( .B(clk), .A(\g.we_clk [26098]));
Q_ASSIGN U6677 ( .B(clk), .A(\g.we_clk [26097]));
Q_ASSIGN U6678 ( .B(clk), .A(\g.we_clk [26096]));
Q_ASSIGN U6679 ( .B(clk), .A(\g.we_clk [26095]));
Q_ASSIGN U6680 ( .B(clk), .A(\g.we_clk [26094]));
Q_ASSIGN U6681 ( .B(clk), .A(\g.we_clk [26093]));
Q_ASSIGN U6682 ( .B(clk), .A(\g.we_clk [26092]));
Q_ASSIGN U6683 ( .B(clk), .A(\g.we_clk [26091]));
Q_ASSIGN U6684 ( .B(clk), .A(\g.we_clk [26090]));
Q_ASSIGN U6685 ( .B(clk), .A(\g.we_clk [26089]));
Q_ASSIGN U6686 ( .B(clk), .A(\g.we_clk [26088]));
Q_ASSIGN U6687 ( .B(clk), .A(\g.we_clk [26087]));
Q_ASSIGN U6688 ( .B(clk), .A(\g.we_clk [26086]));
Q_ASSIGN U6689 ( .B(clk), .A(\g.we_clk [26085]));
Q_ASSIGN U6690 ( .B(clk), .A(\g.we_clk [26084]));
Q_ASSIGN U6691 ( .B(clk), .A(\g.we_clk [26083]));
Q_ASSIGN U6692 ( .B(clk), .A(\g.we_clk [26082]));
Q_ASSIGN U6693 ( .B(clk), .A(\g.we_clk [26081]));
Q_ASSIGN U6694 ( .B(clk), .A(\g.we_clk [26080]));
Q_ASSIGN U6695 ( .B(clk), .A(\g.we_clk [26079]));
Q_ASSIGN U6696 ( .B(clk), .A(\g.we_clk [26078]));
Q_ASSIGN U6697 ( .B(clk), .A(\g.we_clk [26077]));
Q_ASSIGN U6698 ( .B(clk), .A(\g.we_clk [26076]));
Q_ASSIGN U6699 ( .B(clk), .A(\g.we_clk [26075]));
Q_ASSIGN U6700 ( .B(clk), .A(\g.we_clk [26074]));
Q_ASSIGN U6701 ( .B(clk), .A(\g.we_clk [26073]));
Q_ASSIGN U6702 ( .B(clk), .A(\g.we_clk [26072]));
Q_ASSIGN U6703 ( .B(clk), .A(\g.we_clk [26071]));
Q_ASSIGN U6704 ( .B(clk), .A(\g.we_clk [26070]));
Q_ASSIGN U6705 ( .B(clk), .A(\g.we_clk [26069]));
Q_ASSIGN U6706 ( .B(clk), .A(\g.we_clk [26068]));
Q_ASSIGN U6707 ( .B(clk), .A(\g.we_clk [26067]));
Q_ASSIGN U6708 ( .B(clk), .A(\g.we_clk [26066]));
Q_ASSIGN U6709 ( .B(clk), .A(\g.we_clk [26065]));
Q_ASSIGN U6710 ( .B(clk), .A(\g.we_clk [26064]));
Q_ASSIGN U6711 ( .B(clk), .A(\g.we_clk [26063]));
Q_ASSIGN U6712 ( .B(clk), .A(\g.we_clk [26062]));
Q_ASSIGN U6713 ( .B(clk), .A(\g.we_clk [26061]));
Q_ASSIGN U6714 ( .B(clk), .A(\g.we_clk [26060]));
Q_ASSIGN U6715 ( .B(clk), .A(\g.we_clk [26059]));
Q_ASSIGN U6716 ( .B(clk), .A(\g.we_clk [26058]));
Q_ASSIGN U6717 ( .B(clk), .A(\g.we_clk [26057]));
Q_ASSIGN U6718 ( .B(clk), .A(\g.we_clk [26056]));
Q_ASSIGN U6719 ( .B(clk), .A(\g.we_clk [26055]));
Q_ASSIGN U6720 ( .B(clk), .A(\g.we_clk [26054]));
Q_ASSIGN U6721 ( .B(clk), .A(\g.we_clk [26053]));
Q_ASSIGN U6722 ( .B(clk), .A(\g.we_clk [26052]));
Q_ASSIGN U6723 ( .B(clk), .A(\g.we_clk [26051]));
Q_ASSIGN U6724 ( .B(clk), .A(\g.we_clk [26050]));
Q_ASSIGN U6725 ( .B(clk), .A(\g.we_clk [26049]));
Q_ASSIGN U6726 ( .B(clk), .A(\g.we_clk [26048]));
Q_ASSIGN U6727 ( .B(clk), .A(\g.we_clk [26047]));
Q_ASSIGN U6728 ( .B(clk), .A(\g.we_clk [26046]));
Q_ASSIGN U6729 ( .B(clk), .A(\g.we_clk [26045]));
Q_ASSIGN U6730 ( .B(clk), .A(\g.we_clk [26044]));
Q_ASSIGN U6731 ( .B(clk), .A(\g.we_clk [26043]));
Q_ASSIGN U6732 ( .B(clk), .A(\g.we_clk [26042]));
Q_ASSIGN U6733 ( .B(clk), .A(\g.we_clk [26041]));
Q_ASSIGN U6734 ( .B(clk), .A(\g.we_clk [26040]));
Q_ASSIGN U6735 ( .B(clk), .A(\g.we_clk [26039]));
Q_ASSIGN U6736 ( .B(clk), .A(\g.we_clk [26038]));
Q_ASSIGN U6737 ( .B(clk), .A(\g.we_clk [26037]));
Q_ASSIGN U6738 ( .B(clk), .A(\g.we_clk [26036]));
Q_ASSIGN U6739 ( .B(clk), .A(\g.we_clk [26035]));
Q_ASSIGN U6740 ( .B(clk), .A(\g.we_clk [26034]));
Q_ASSIGN U6741 ( .B(clk), .A(\g.we_clk [26033]));
Q_ASSIGN U6742 ( .B(clk), .A(\g.we_clk [26032]));
Q_ASSIGN U6743 ( .B(clk), .A(\g.we_clk [26031]));
Q_ASSIGN U6744 ( .B(clk), .A(\g.we_clk [26030]));
Q_ASSIGN U6745 ( .B(clk), .A(\g.we_clk [26029]));
Q_ASSIGN U6746 ( .B(clk), .A(\g.we_clk [26028]));
Q_ASSIGN U6747 ( .B(clk), .A(\g.we_clk [26027]));
Q_ASSIGN U6748 ( .B(clk), .A(\g.we_clk [26026]));
Q_ASSIGN U6749 ( .B(clk), .A(\g.we_clk [26025]));
Q_ASSIGN U6750 ( .B(clk), .A(\g.we_clk [26024]));
Q_ASSIGN U6751 ( .B(clk), .A(\g.we_clk [26023]));
Q_ASSIGN U6752 ( .B(clk), .A(\g.we_clk [26022]));
Q_ASSIGN U6753 ( .B(clk), .A(\g.we_clk [26021]));
Q_ASSIGN U6754 ( .B(clk), .A(\g.we_clk [26020]));
Q_ASSIGN U6755 ( .B(clk), .A(\g.we_clk [26019]));
Q_ASSIGN U6756 ( .B(clk), .A(\g.we_clk [26018]));
Q_ASSIGN U6757 ( .B(clk), .A(\g.we_clk [26017]));
Q_ASSIGN U6758 ( .B(clk), .A(\g.we_clk [26016]));
Q_ASSIGN U6759 ( .B(clk), .A(\g.we_clk [26015]));
Q_ASSIGN U6760 ( .B(clk), .A(\g.we_clk [26014]));
Q_ASSIGN U6761 ( .B(clk), .A(\g.we_clk [26013]));
Q_ASSIGN U6762 ( .B(clk), .A(\g.we_clk [26012]));
Q_ASSIGN U6763 ( .B(clk), .A(\g.we_clk [26011]));
Q_ASSIGN U6764 ( .B(clk), .A(\g.we_clk [26010]));
Q_ASSIGN U6765 ( .B(clk), .A(\g.we_clk [26009]));
Q_ASSIGN U6766 ( .B(clk), .A(\g.we_clk [26008]));
Q_ASSIGN U6767 ( .B(clk), .A(\g.we_clk [26007]));
Q_ASSIGN U6768 ( .B(clk), .A(\g.we_clk [26006]));
Q_ASSIGN U6769 ( .B(clk), .A(\g.we_clk [26005]));
Q_ASSIGN U6770 ( .B(clk), .A(\g.we_clk [26004]));
Q_ASSIGN U6771 ( .B(clk), .A(\g.we_clk [26003]));
Q_ASSIGN U6772 ( .B(clk), .A(\g.we_clk [26002]));
Q_ASSIGN U6773 ( .B(clk), .A(\g.we_clk [26001]));
Q_ASSIGN U6774 ( .B(clk), .A(\g.we_clk [26000]));
Q_ASSIGN U6775 ( .B(clk), .A(\g.we_clk [25999]));
Q_ASSIGN U6776 ( .B(clk), .A(\g.we_clk [25998]));
Q_ASSIGN U6777 ( .B(clk), .A(\g.we_clk [25997]));
Q_ASSIGN U6778 ( .B(clk), .A(\g.we_clk [25996]));
Q_ASSIGN U6779 ( .B(clk), .A(\g.we_clk [25995]));
Q_ASSIGN U6780 ( .B(clk), .A(\g.we_clk [25994]));
Q_ASSIGN U6781 ( .B(clk), .A(\g.we_clk [25993]));
Q_ASSIGN U6782 ( .B(clk), .A(\g.we_clk [25992]));
Q_ASSIGN U6783 ( .B(clk), .A(\g.we_clk [25991]));
Q_ASSIGN U6784 ( .B(clk), .A(\g.we_clk [25990]));
Q_ASSIGN U6785 ( .B(clk), .A(\g.we_clk [25989]));
Q_ASSIGN U6786 ( .B(clk), .A(\g.we_clk [25988]));
Q_ASSIGN U6787 ( .B(clk), .A(\g.we_clk [25987]));
Q_ASSIGN U6788 ( .B(clk), .A(\g.we_clk [25986]));
Q_ASSIGN U6789 ( .B(clk), .A(\g.we_clk [25985]));
Q_ASSIGN U6790 ( .B(clk), .A(\g.we_clk [25984]));
Q_ASSIGN U6791 ( .B(clk), .A(\g.we_clk [25983]));
Q_ASSIGN U6792 ( .B(clk), .A(\g.we_clk [25982]));
Q_ASSIGN U6793 ( .B(clk), .A(\g.we_clk [25981]));
Q_ASSIGN U6794 ( .B(clk), .A(\g.we_clk [25980]));
Q_ASSIGN U6795 ( .B(clk), .A(\g.we_clk [25979]));
Q_ASSIGN U6796 ( .B(clk), .A(\g.we_clk [25978]));
Q_ASSIGN U6797 ( .B(clk), .A(\g.we_clk [25977]));
Q_ASSIGN U6798 ( .B(clk), .A(\g.we_clk [25976]));
Q_ASSIGN U6799 ( .B(clk), .A(\g.we_clk [25975]));
Q_ASSIGN U6800 ( .B(clk), .A(\g.we_clk [25974]));
Q_ASSIGN U6801 ( .B(clk), .A(\g.we_clk [25973]));
Q_ASSIGN U6802 ( .B(clk), .A(\g.we_clk [25972]));
Q_ASSIGN U6803 ( .B(clk), .A(\g.we_clk [25971]));
Q_ASSIGN U6804 ( .B(clk), .A(\g.we_clk [25970]));
Q_ASSIGN U6805 ( .B(clk), .A(\g.we_clk [25969]));
Q_ASSIGN U6806 ( .B(clk), .A(\g.we_clk [25968]));
Q_ASSIGN U6807 ( .B(clk), .A(\g.we_clk [25967]));
Q_ASSIGN U6808 ( .B(clk), .A(\g.we_clk [25966]));
Q_ASSIGN U6809 ( .B(clk), .A(\g.we_clk [25965]));
Q_ASSIGN U6810 ( .B(clk), .A(\g.we_clk [25964]));
Q_ASSIGN U6811 ( .B(clk), .A(\g.we_clk [25963]));
Q_ASSIGN U6812 ( .B(clk), .A(\g.we_clk [25962]));
Q_ASSIGN U6813 ( .B(clk), .A(\g.we_clk [25961]));
Q_ASSIGN U6814 ( .B(clk), .A(\g.we_clk [25960]));
Q_ASSIGN U6815 ( .B(clk), .A(\g.we_clk [25959]));
Q_ASSIGN U6816 ( .B(clk), .A(\g.we_clk [25958]));
Q_ASSIGN U6817 ( .B(clk), .A(\g.we_clk [25957]));
Q_ASSIGN U6818 ( .B(clk), .A(\g.we_clk [25956]));
Q_ASSIGN U6819 ( .B(clk), .A(\g.we_clk [25955]));
Q_ASSIGN U6820 ( .B(clk), .A(\g.we_clk [25954]));
Q_ASSIGN U6821 ( .B(clk), .A(\g.we_clk [25953]));
Q_ASSIGN U6822 ( .B(clk), .A(\g.we_clk [25952]));
Q_ASSIGN U6823 ( .B(clk), .A(\g.we_clk [25951]));
Q_ASSIGN U6824 ( .B(clk), .A(\g.we_clk [25950]));
Q_ASSIGN U6825 ( .B(clk), .A(\g.we_clk [25949]));
Q_ASSIGN U6826 ( .B(clk), .A(\g.we_clk [25948]));
Q_ASSIGN U6827 ( .B(clk), .A(\g.we_clk [25947]));
Q_ASSIGN U6828 ( .B(clk), .A(\g.we_clk [25946]));
Q_ASSIGN U6829 ( .B(clk), .A(\g.we_clk [25945]));
Q_ASSIGN U6830 ( .B(clk), .A(\g.we_clk [25944]));
Q_ASSIGN U6831 ( .B(clk), .A(\g.we_clk [25943]));
Q_ASSIGN U6832 ( .B(clk), .A(\g.we_clk [25942]));
Q_ASSIGN U6833 ( .B(clk), .A(\g.we_clk [25941]));
Q_ASSIGN U6834 ( .B(clk), .A(\g.we_clk [25940]));
Q_ASSIGN U6835 ( .B(clk), .A(\g.we_clk [25939]));
Q_ASSIGN U6836 ( .B(clk), .A(\g.we_clk [25938]));
Q_ASSIGN U6837 ( .B(clk), .A(\g.we_clk [25937]));
Q_ASSIGN U6838 ( .B(clk), .A(\g.we_clk [25936]));
Q_ASSIGN U6839 ( .B(clk), .A(\g.we_clk [25935]));
Q_ASSIGN U6840 ( .B(clk), .A(\g.we_clk [25934]));
Q_ASSIGN U6841 ( .B(clk), .A(\g.we_clk [25933]));
Q_ASSIGN U6842 ( .B(clk), .A(\g.we_clk [25932]));
Q_ASSIGN U6843 ( .B(clk), .A(\g.we_clk [25931]));
Q_ASSIGN U6844 ( .B(clk), .A(\g.we_clk [25930]));
Q_ASSIGN U6845 ( .B(clk), .A(\g.we_clk [25929]));
Q_ASSIGN U6846 ( .B(clk), .A(\g.we_clk [25928]));
Q_ASSIGN U6847 ( .B(clk), .A(\g.we_clk [25927]));
Q_ASSIGN U6848 ( .B(clk), .A(\g.we_clk [25926]));
Q_ASSIGN U6849 ( .B(clk), .A(\g.we_clk [25925]));
Q_ASSIGN U6850 ( .B(clk), .A(\g.we_clk [25924]));
Q_ASSIGN U6851 ( .B(clk), .A(\g.we_clk [25923]));
Q_ASSIGN U6852 ( .B(clk), .A(\g.we_clk [25922]));
Q_ASSIGN U6853 ( .B(clk), .A(\g.we_clk [25921]));
Q_ASSIGN U6854 ( .B(clk), .A(\g.we_clk [25920]));
Q_ASSIGN U6855 ( .B(clk), .A(\g.we_clk [25919]));
Q_ASSIGN U6856 ( .B(clk), .A(\g.we_clk [25918]));
Q_ASSIGN U6857 ( .B(clk), .A(\g.we_clk [25917]));
Q_ASSIGN U6858 ( .B(clk), .A(\g.we_clk [25916]));
Q_ASSIGN U6859 ( .B(clk), .A(\g.we_clk [25915]));
Q_ASSIGN U6860 ( .B(clk), .A(\g.we_clk [25914]));
Q_ASSIGN U6861 ( .B(clk), .A(\g.we_clk [25913]));
Q_ASSIGN U6862 ( .B(clk), .A(\g.we_clk [25912]));
Q_ASSIGN U6863 ( .B(clk), .A(\g.we_clk [25911]));
Q_ASSIGN U6864 ( .B(clk), .A(\g.we_clk [25910]));
Q_ASSIGN U6865 ( .B(clk), .A(\g.we_clk [25909]));
Q_ASSIGN U6866 ( .B(clk), .A(\g.we_clk [25908]));
Q_ASSIGN U6867 ( .B(clk), .A(\g.we_clk [25907]));
Q_ASSIGN U6868 ( .B(clk), .A(\g.we_clk [25906]));
Q_ASSIGN U6869 ( .B(clk), .A(\g.we_clk [25905]));
Q_ASSIGN U6870 ( .B(clk), .A(\g.we_clk [25904]));
Q_ASSIGN U6871 ( .B(clk), .A(\g.we_clk [25903]));
Q_ASSIGN U6872 ( .B(clk), .A(\g.we_clk [25902]));
Q_ASSIGN U6873 ( .B(clk), .A(\g.we_clk [25901]));
Q_ASSIGN U6874 ( .B(clk), .A(\g.we_clk [25900]));
Q_ASSIGN U6875 ( .B(clk), .A(\g.we_clk [25899]));
Q_ASSIGN U6876 ( .B(clk), .A(\g.we_clk [25898]));
Q_ASSIGN U6877 ( .B(clk), .A(\g.we_clk [25897]));
Q_ASSIGN U6878 ( .B(clk), .A(\g.we_clk [25896]));
Q_ASSIGN U6879 ( .B(clk), .A(\g.we_clk [25895]));
Q_ASSIGN U6880 ( .B(clk), .A(\g.we_clk [25894]));
Q_ASSIGN U6881 ( .B(clk), .A(\g.we_clk [25893]));
Q_ASSIGN U6882 ( .B(clk), .A(\g.we_clk [25892]));
Q_ASSIGN U6883 ( .B(clk), .A(\g.we_clk [25891]));
Q_ASSIGN U6884 ( .B(clk), .A(\g.we_clk [25890]));
Q_ASSIGN U6885 ( .B(clk), .A(\g.we_clk [25889]));
Q_ASSIGN U6886 ( .B(clk), .A(\g.we_clk [25888]));
Q_ASSIGN U6887 ( .B(clk), .A(\g.we_clk [25887]));
Q_ASSIGN U6888 ( .B(clk), .A(\g.we_clk [25886]));
Q_ASSIGN U6889 ( .B(clk), .A(\g.we_clk [25885]));
Q_ASSIGN U6890 ( .B(clk), .A(\g.we_clk [25884]));
Q_ASSIGN U6891 ( .B(clk), .A(\g.we_clk [25883]));
Q_ASSIGN U6892 ( .B(clk), .A(\g.we_clk [25882]));
Q_ASSIGN U6893 ( .B(clk), .A(\g.we_clk [25881]));
Q_ASSIGN U6894 ( .B(clk), .A(\g.we_clk [25880]));
Q_ASSIGN U6895 ( .B(clk), .A(\g.we_clk [25879]));
Q_ASSIGN U6896 ( .B(clk), .A(\g.we_clk [25878]));
Q_ASSIGN U6897 ( .B(clk), .A(\g.we_clk [25877]));
Q_ASSIGN U6898 ( .B(clk), .A(\g.we_clk [25876]));
Q_ASSIGN U6899 ( .B(clk), .A(\g.we_clk [25875]));
Q_ASSIGN U6900 ( .B(clk), .A(\g.we_clk [25874]));
Q_ASSIGN U6901 ( .B(clk), .A(\g.we_clk [25873]));
Q_ASSIGN U6902 ( .B(clk), .A(\g.we_clk [25872]));
Q_ASSIGN U6903 ( .B(clk), .A(\g.we_clk [25871]));
Q_ASSIGN U6904 ( .B(clk), .A(\g.we_clk [25870]));
Q_ASSIGN U6905 ( .B(clk), .A(\g.we_clk [25869]));
Q_ASSIGN U6906 ( .B(clk), .A(\g.we_clk [25868]));
Q_ASSIGN U6907 ( .B(clk), .A(\g.we_clk [25867]));
Q_ASSIGN U6908 ( .B(clk), .A(\g.we_clk [25866]));
Q_ASSIGN U6909 ( .B(clk), .A(\g.we_clk [25865]));
Q_ASSIGN U6910 ( .B(clk), .A(\g.we_clk [25864]));
Q_ASSIGN U6911 ( .B(clk), .A(\g.we_clk [25863]));
Q_ASSIGN U6912 ( .B(clk), .A(\g.we_clk [25862]));
Q_ASSIGN U6913 ( .B(clk), .A(\g.we_clk [25861]));
Q_ASSIGN U6914 ( .B(clk), .A(\g.we_clk [25860]));
Q_ASSIGN U6915 ( .B(clk), .A(\g.we_clk [25859]));
Q_ASSIGN U6916 ( .B(clk), .A(\g.we_clk [25858]));
Q_ASSIGN U6917 ( .B(clk), .A(\g.we_clk [25857]));
Q_ASSIGN U6918 ( .B(clk), .A(\g.we_clk [25856]));
Q_ASSIGN U6919 ( .B(clk), .A(\g.we_clk [25855]));
Q_ASSIGN U6920 ( .B(clk), .A(\g.we_clk [25854]));
Q_ASSIGN U6921 ( .B(clk), .A(\g.we_clk [25853]));
Q_ASSIGN U6922 ( .B(clk), .A(\g.we_clk [25852]));
Q_ASSIGN U6923 ( .B(clk), .A(\g.we_clk [25851]));
Q_ASSIGN U6924 ( .B(clk), .A(\g.we_clk [25850]));
Q_ASSIGN U6925 ( .B(clk), .A(\g.we_clk [25849]));
Q_ASSIGN U6926 ( .B(clk), .A(\g.we_clk [25848]));
Q_ASSIGN U6927 ( .B(clk), .A(\g.we_clk [25847]));
Q_ASSIGN U6928 ( .B(clk), .A(\g.we_clk [25846]));
Q_ASSIGN U6929 ( .B(clk), .A(\g.we_clk [25845]));
Q_ASSIGN U6930 ( .B(clk), .A(\g.we_clk [25844]));
Q_ASSIGN U6931 ( .B(clk), .A(\g.we_clk [25843]));
Q_ASSIGN U6932 ( .B(clk), .A(\g.we_clk [25842]));
Q_ASSIGN U6933 ( .B(clk), .A(\g.we_clk [25841]));
Q_ASSIGN U6934 ( .B(clk), .A(\g.we_clk [25840]));
Q_ASSIGN U6935 ( .B(clk), .A(\g.we_clk [25839]));
Q_ASSIGN U6936 ( .B(clk), .A(\g.we_clk [25838]));
Q_ASSIGN U6937 ( .B(clk), .A(\g.we_clk [25837]));
Q_ASSIGN U6938 ( .B(clk), .A(\g.we_clk [25836]));
Q_ASSIGN U6939 ( .B(clk), .A(\g.we_clk [25835]));
Q_ASSIGN U6940 ( .B(clk), .A(\g.we_clk [25834]));
Q_ASSIGN U6941 ( .B(clk), .A(\g.we_clk [25833]));
Q_ASSIGN U6942 ( .B(clk), .A(\g.we_clk [25832]));
Q_ASSIGN U6943 ( .B(clk), .A(\g.we_clk [25831]));
Q_ASSIGN U6944 ( .B(clk), .A(\g.we_clk [25830]));
Q_ASSIGN U6945 ( .B(clk), .A(\g.we_clk [25829]));
Q_ASSIGN U6946 ( .B(clk), .A(\g.we_clk [25828]));
Q_ASSIGN U6947 ( .B(clk), .A(\g.we_clk [25827]));
Q_ASSIGN U6948 ( .B(clk), .A(\g.we_clk [25826]));
Q_ASSIGN U6949 ( .B(clk), .A(\g.we_clk [25825]));
Q_ASSIGN U6950 ( .B(clk), .A(\g.we_clk [25824]));
Q_ASSIGN U6951 ( .B(clk), .A(\g.we_clk [25823]));
Q_ASSIGN U6952 ( .B(clk), .A(\g.we_clk [25822]));
Q_ASSIGN U6953 ( .B(clk), .A(\g.we_clk [25821]));
Q_ASSIGN U6954 ( .B(clk), .A(\g.we_clk [25820]));
Q_ASSIGN U6955 ( .B(clk), .A(\g.we_clk [25819]));
Q_ASSIGN U6956 ( .B(clk), .A(\g.we_clk [25818]));
Q_ASSIGN U6957 ( .B(clk), .A(\g.we_clk [25817]));
Q_ASSIGN U6958 ( .B(clk), .A(\g.we_clk [25816]));
Q_ASSIGN U6959 ( .B(clk), .A(\g.we_clk [25815]));
Q_ASSIGN U6960 ( .B(clk), .A(\g.we_clk [25814]));
Q_ASSIGN U6961 ( .B(clk), .A(\g.we_clk [25813]));
Q_ASSIGN U6962 ( .B(clk), .A(\g.we_clk [25812]));
Q_ASSIGN U6963 ( .B(clk), .A(\g.we_clk [25811]));
Q_ASSIGN U6964 ( .B(clk), .A(\g.we_clk [25810]));
Q_ASSIGN U6965 ( .B(clk), .A(\g.we_clk [25809]));
Q_ASSIGN U6966 ( .B(clk), .A(\g.we_clk [25808]));
Q_ASSIGN U6967 ( .B(clk), .A(\g.we_clk [25807]));
Q_ASSIGN U6968 ( .B(clk), .A(\g.we_clk [25806]));
Q_ASSIGN U6969 ( .B(clk), .A(\g.we_clk [25805]));
Q_ASSIGN U6970 ( .B(clk), .A(\g.we_clk [25804]));
Q_ASSIGN U6971 ( .B(clk), .A(\g.we_clk [25803]));
Q_ASSIGN U6972 ( .B(clk), .A(\g.we_clk [25802]));
Q_ASSIGN U6973 ( .B(clk), .A(\g.we_clk [25801]));
Q_ASSIGN U6974 ( .B(clk), .A(\g.we_clk [25800]));
Q_ASSIGN U6975 ( .B(clk), .A(\g.we_clk [25799]));
Q_ASSIGN U6976 ( .B(clk), .A(\g.we_clk [25798]));
Q_ASSIGN U6977 ( .B(clk), .A(\g.we_clk [25797]));
Q_ASSIGN U6978 ( .B(clk), .A(\g.we_clk [25796]));
Q_ASSIGN U6979 ( .B(clk), .A(\g.we_clk [25795]));
Q_ASSIGN U6980 ( .B(clk), .A(\g.we_clk [25794]));
Q_ASSIGN U6981 ( .B(clk), .A(\g.we_clk [25793]));
Q_ASSIGN U6982 ( .B(clk), .A(\g.we_clk [25792]));
Q_ASSIGN U6983 ( .B(clk), .A(\g.we_clk [25791]));
Q_ASSIGN U6984 ( .B(clk), .A(\g.we_clk [25790]));
Q_ASSIGN U6985 ( .B(clk), .A(\g.we_clk [25789]));
Q_ASSIGN U6986 ( .B(clk), .A(\g.we_clk [25788]));
Q_ASSIGN U6987 ( .B(clk), .A(\g.we_clk [25787]));
Q_ASSIGN U6988 ( .B(clk), .A(\g.we_clk [25786]));
Q_ASSIGN U6989 ( .B(clk), .A(\g.we_clk [25785]));
Q_ASSIGN U6990 ( .B(clk), .A(\g.we_clk [25784]));
Q_ASSIGN U6991 ( .B(clk), .A(\g.we_clk [25783]));
Q_ASSIGN U6992 ( .B(clk), .A(\g.we_clk [25782]));
Q_ASSIGN U6993 ( .B(clk), .A(\g.we_clk [25781]));
Q_ASSIGN U6994 ( .B(clk), .A(\g.we_clk [25780]));
Q_ASSIGN U6995 ( .B(clk), .A(\g.we_clk [25779]));
Q_ASSIGN U6996 ( .B(clk), .A(\g.we_clk [25778]));
Q_ASSIGN U6997 ( .B(clk), .A(\g.we_clk [25777]));
Q_ASSIGN U6998 ( .B(clk), .A(\g.we_clk [25776]));
Q_ASSIGN U6999 ( .B(clk), .A(\g.we_clk [25775]));
Q_ASSIGN U7000 ( .B(clk), .A(\g.we_clk [25774]));
Q_ASSIGN U7001 ( .B(clk), .A(\g.we_clk [25773]));
Q_ASSIGN U7002 ( .B(clk), .A(\g.we_clk [25772]));
Q_ASSIGN U7003 ( .B(clk), .A(\g.we_clk [25771]));
Q_ASSIGN U7004 ( .B(clk), .A(\g.we_clk [25770]));
Q_ASSIGN U7005 ( .B(clk), .A(\g.we_clk [25769]));
Q_ASSIGN U7006 ( .B(clk), .A(\g.we_clk [25768]));
Q_ASSIGN U7007 ( .B(clk), .A(\g.we_clk [25767]));
Q_ASSIGN U7008 ( .B(clk), .A(\g.we_clk [25766]));
Q_ASSIGN U7009 ( .B(clk), .A(\g.we_clk [25765]));
Q_ASSIGN U7010 ( .B(clk), .A(\g.we_clk [25764]));
Q_ASSIGN U7011 ( .B(clk), .A(\g.we_clk [25763]));
Q_ASSIGN U7012 ( .B(clk), .A(\g.we_clk [25762]));
Q_ASSIGN U7013 ( .B(clk), .A(\g.we_clk [25761]));
Q_ASSIGN U7014 ( .B(clk), .A(\g.we_clk [25760]));
Q_ASSIGN U7015 ( .B(clk), .A(\g.we_clk [25759]));
Q_ASSIGN U7016 ( .B(clk), .A(\g.we_clk [25758]));
Q_ASSIGN U7017 ( .B(clk), .A(\g.we_clk [25757]));
Q_ASSIGN U7018 ( .B(clk), .A(\g.we_clk [25756]));
Q_ASSIGN U7019 ( .B(clk), .A(\g.we_clk [25755]));
Q_ASSIGN U7020 ( .B(clk), .A(\g.we_clk [25754]));
Q_ASSIGN U7021 ( .B(clk), .A(\g.we_clk [25753]));
Q_ASSIGN U7022 ( .B(clk), .A(\g.we_clk [25752]));
Q_ASSIGN U7023 ( .B(clk), .A(\g.we_clk [25751]));
Q_ASSIGN U7024 ( .B(clk), .A(\g.we_clk [25750]));
Q_ASSIGN U7025 ( .B(clk), .A(\g.we_clk [25749]));
Q_ASSIGN U7026 ( .B(clk), .A(\g.we_clk [25748]));
Q_ASSIGN U7027 ( .B(clk), .A(\g.we_clk [25747]));
Q_ASSIGN U7028 ( .B(clk), .A(\g.we_clk [25746]));
Q_ASSIGN U7029 ( .B(clk), .A(\g.we_clk [25745]));
Q_ASSIGN U7030 ( .B(clk), .A(\g.we_clk [25744]));
Q_ASSIGN U7031 ( .B(clk), .A(\g.we_clk [25743]));
Q_ASSIGN U7032 ( .B(clk), .A(\g.we_clk [25742]));
Q_ASSIGN U7033 ( .B(clk), .A(\g.we_clk [25741]));
Q_ASSIGN U7034 ( .B(clk), .A(\g.we_clk [25740]));
Q_ASSIGN U7035 ( .B(clk), .A(\g.we_clk [25739]));
Q_ASSIGN U7036 ( .B(clk), .A(\g.we_clk [25738]));
Q_ASSIGN U7037 ( .B(clk), .A(\g.we_clk [25737]));
Q_ASSIGN U7038 ( .B(clk), .A(\g.we_clk [25736]));
Q_ASSIGN U7039 ( .B(clk), .A(\g.we_clk [25735]));
Q_ASSIGN U7040 ( .B(clk), .A(\g.we_clk [25734]));
Q_ASSIGN U7041 ( .B(clk), .A(\g.we_clk [25733]));
Q_ASSIGN U7042 ( .B(clk), .A(\g.we_clk [25732]));
Q_ASSIGN U7043 ( .B(clk), .A(\g.we_clk [25731]));
Q_ASSIGN U7044 ( .B(clk), .A(\g.we_clk [25730]));
Q_ASSIGN U7045 ( .B(clk), .A(\g.we_clk [25729]));
Q_ASSIGN U7046 ( .B(clk), .A(\g.we_clk [25728]));
Q_ASSIGN U7047 ( .B(clk), .A(\g.we_clk [25727]));
Q_ASSIGN U7048 ( .B(clk), .A(\g.we_clk [25726]));
Q_ASSIGN U7049 ( .B(clk), .A(\g.we_clk [25725]));
Q_ASSIGN U7050 ( .B(clk), .A(\g.we_clk [25724]));
Q_ASSIGN U7051 ( .B(clk), .A(\g.we_clk [25723]));
Q_ASSIGN U7052 ( .B(clk), .A(\g.we_clk [25722]));
Q_ASSIGN U7053 ( .B(clk), .A(\g.we_clk [25721]));
Q_ASSIGN U7054 ( .B(clk), .A(\g.we_clk [25720]));
Q_ASSIGN U7055 ( .B(clk), .A(\g.we_clk [25719]));
Q_ASSIGN U7056 ( .B(clk), .A(\g.we_clk [25718]));
Q_ASSIGN U7057 ( .B(clk), .A(\g.we_clk [25717]));
Q_ASSIGN U7058 ( .B(clk), .A(\g.we_clk [25716]));
Q_ASSIGN U7059 ( .B(clk), .A(\g.we_clk [25715]));
Q_ASSIGN U7060 ( .B(clk), .A(\g.we_clk [25714]));
Q_ASSIGN U7061 ( .B(clk), .A(\g.we_clk [25713]));
Q_ASSIGN U7062 ( .B(clk), .A(\g.we_clk [25712]));
Q_ASSIGN U7063 ( .B(clk), .A(\g.we_clk [25711]));
Q_ASSIGN U7064 ( .B(clk), .A(\g.we_clk [25710]));
Q_ASSIGN U7065 ( .B(clk), .A(\g.we_clk [25709]));
Q_ASSIGN U7066 ( .B(clk), .A(\g.we_clk [25708]));
Q_ASSIGN U7067 ( .B(clk), .A(\g.we_clk [25707]));
Q_ASSIGN U7068 ( .B(clk), .A(\g.we_clk [25706]));
Q_ASSIGN U7069 ( .B(clk), .A(\g.we_clk [25705]));
Q_ASSIGN U7070 ( .B(clk), .A(\g.we_clk [25704]));
Q_ASSIGN U7071 ( .B(clk), .A(\g.we_clk [25703]));
Q_ASSIGN U7072 ( .B(clk), .A(\g.we_clk [25702]));
Q_ASSIGN U7073 ( .B(clk), .A(\g.we_clk [25701]));
Q_ASSIGN U7074 ( .B(clk), .A(\g.we_clk [25700]));
Q_ASSIGN U7075 ( .B(clk), .A(\g.we_clk [25699]));
Q_ASSIGN U7076 ( .B(clk), .A(\g.we_clk [25698]));
Q_ASSIGN U7077 ( .B(clk), .A(\g.we_clk [25697]));
Q_ASSIGN U7078 ( .B(clk), .A(\g.we_clk [25696]));
Q_ASSIGN U7079 ( .B(clk), .A(\g.we_clk [25695]));
Q_ASSIGN U7080 ( .B(clk), .A(\g.we_clk [25694]));
Q_ASSIGN U7081 ( .B(clk), .A(\g.we_clk [25693]));
Q_ASSIGN U7082 ( .B(clk), .A(\g.we_clk [25692]));
Q_ASSIGN U7083 ( .B(clk), .A(\g.we_clk [25691]));
Q_ASSIGN U7084 ( .B(clk), .A(\g.we_clk [25690]));
Q_ASSIGN U7085 ( .B(clk), .A(\g.we_clk [25689]));
Q_ASSIGN U7086 ( .B(clk), .A(\g.we_clk [25688]));
Q_ASSIGN U7087 ( .B(clk), .A(\g.we_clk [25687]));
Q_ASSIGN U7088 ( .B(clk), .A(\g.we_clk [25686]));
Q_ASSIGN U7089 ( .B(clk), .A(\g.we_clk [25685]));
Q_ASSIGN U7090 ( .B(clk), .A(\g.we_clk [25684]));
Q_ASSIGN U7091 ( .B(clk), .A(\g.we_clk [25683]));
Q_ASSIGN U7092 ( .B(clk), .A(\g.we_clk [25682]));
Q_ASSIGN U7093 ( .B(clk), .A(\g.we_clk [25681]));
Q_ASSIGN U7094 ( .B(clk), .A(\g.we_clk [25680]));
Q_ASSIGN U7095 ( .B(clk), .A(\g.we_clk [25679]));
Q_ASSIGN U7096 ( .B(clk), .A(\g.we_clk [25678]));
Q_ASSIGN U7097 ( .B(clk), .A(\g.we_clk [25677]));
Q_ASSIGN U7098 ( .B(clk), .A(\g.we_clk [25676]));
Q_ASSIGN U7099 ( .B(clk), .A(\g.we_clk [25675]));
Q_ASSIGN U7100 ( .B(clk), .A(\g.we_clk [25674]));
Q_ASSIGN U7101 ( .B(clk), .A(\g.we_clk [25673]));
Q_ASSIGN U7102 ( .B(clk), .A(\g.we_clk [25672]));
Q_ASSIGN U7103 ( .B(clk), .A(\g.we_clk [25671]));
Q_ASSIGN U7104 ( .B(clk), .A(\g.we_clk [25670]));
Q_ASSIGN U7105 ( .B(clk), .A(\g.we_clk [25669]));
Q_ASSIGN U7106 ( .B(clk), .A(\g.we_clk [25668]));
Q_ASSIGN U7107 ( .B(clk), .A(\g.we_clk [25667]));
Q_ASSIGN U7108 ( .B(clk), .A(\g.we_clk [25666]));
Q_ASSIGN U7109 ( .B(clk), .A(\g.we_clk [25665]));
Q_ASSIGN U7110 ( .B(clk), .A(\g.we_clk [25664]));
Q_ASSIGN U7111 ( .B(clk), .A(\g.we_clk [25663]));
Q_ASSIGN U7112 ( .B(clk), .A(\g.we_clk [25662]));
Q_ASSIGN U7113 ( .B(clk), .A(\g.we_clk [25661]));
Q_ASSIGN U7114 ( .B(clk), .A(\g.we_clk [25660]));
Q_ASSIGN U7115 ( .B(clk), .A(\g.we_clk [25659]));
Q_ASSIGN U7116 ( .B(clk), .A(\g.we_clk [25658]));
Q_ASSIGN U7117 ( .B(clk), .A(\g.we_clk [25657]));
Q_ASSIGN U7118 ( .B(clk), .A(\g.we_clk [25656]));
Q_ASSIGN U7119 ( .B(clk), .A(\g.we_clk [25655]));
Q_ASSIGN U7120 ( .B(clk), .A(\g.we_clk [25654]));
Q_ASSIGN U7121 ( .B(clk), .A(\g.we_clk [25653]));
Q_ASSIGN U7122 ( .B(clk), .A(\g.we_clk [25652]));
Q_ASSIGN U7123 ( .B(clk), .A(\g.we_clk [25651]));
Q_ASSIGN U7124 ( .B(clk), .A(\g.we_clk [25650]));
Q_ASSIGN U7125 ( .B(clk), .A(\g.we_clk [25649]));
Q_ASSIGN U7126 ( .B(clk), .A(\g.we_clk [25648]));
Q_ASSIGN U7127 ( .B(clk), .A(\g.we_clk [25647]));
Q_ASSIGN U7128 ( .B(clk), .A(\g.we_clk [25646]));
Q_ASSIGN U7129 ( .B(clk), .A(\g.we_clk [25645]));
Q_ASSIGN U7130 ( .B(clk), .A(\g.we_clk [25644]));
Q_ASSIGN U7131 ( .B(clk), .A(\g.we_clk [25643]));
Q_ASSIGN U7132 ( .B(clk), .A(\g.we_clk [25642]));
Q_ASSIGN U7133 ( .B(clk), .A(\g.we_clk [25641]));
Q_ASSIGN U7134 ( .B(clk), .A(\g.we_clk [25640]));
Q_ASSIGN U7135 ( .B(clk), .A(\g.we_clk [25639]));
Q_ASSIGN U7136 ( .B(clk), .A(\g.we_clk [25638]));
Q_ASSIGN U7137 ( .B(clk), .A(\g.we_clk [25637]));
Q_ASSIGN U7138 ( .B(clk), .A(\g.we_clk [25636]));
Q_ASSIGN U7139 ( .B(clk), .A(\g.we_clk [25635]));
Q_ASSIGN U7140 ( .B(clk), .A(\g.we_clk [25634]));
Q_ASSIGN U7141 ( .B(clk), .A(\g.we_clk [25633]));
Q_ASSIGN U7142 ( .B(clk), .A(\g.we_clk [25632]));
Q_ASSIGN U7143 ( .B(clk), .A(\g.we_clk [25631]));
Q_ASSIGN U7144 ( .B(clk), .A(\g.we_clk [25630]));
Q_ASSIGN U7145 ( .B(clk), .A(\g.we_clk [25629]));
Q_ASSIGN U7146 ( .B(clk), .A(\g.we_clk [25628]));
Q_ASSIGN U7147 ( .B(clk), .A(\g.we_clk [25627]));
Q_ASSIGN U7148 ( .B(clk), .A(\g.we_clk [25626]));
Q_ASSIGN U7149 ( .B(clk), .A(\g.we_clk [25625]));
Q_ASSIGN U7150 ( .B(clk), .A(\g.we_clk [25624]));
Q_ASSIGN U7151 ( .B(clk), .A(\g.we_clk [25623]));
Q_ASSIGN U7152 ( .B(clk), .A(\g.we_clk [25622]));
Q_ASSIGN U7153 ( .B(clk), .A(\g.we_clk [25621]));
Q_ASSIGN U7154 ( .B(clk), .A(\g.we_clk [25620]));
Q_ASSIGN U7155 ( .B(clk), .A(\g.we_clk [25619]));
Q_ASSIGN U7156 ( .B(clk), .A(\g.we_clk [25618]));
Q_ASSIGN U7157 ( .B(clk), .A(\g.we_clk [25617]));
Q_ASSIGN U7158 ( .B(clk), .A(\g.we_clk [25616]));
Q_ASSIGN U7159 ( .B(clk), .A(\g.we_clk [25615]));
Q_ASSIGN U7160 ( .B(clk), .A(\g.we_clk [25614]));
Q_ASSIGN U7161 ( .B(clk), .A(\g.we_clk [25613]));
Q_ASSIGN U7162 ( .B(clk), .A(\g.we_clk [25612]));
Q_ASSIGN U7163 ( .B(clk), .A(\g.we_clk [25611]));
Q_ASSIGN U7164 ( .B(clk), .A(\g.we_clk [25610]));
Q_ASSIGN U7165 ( .B(clk), .A(\g.we_clk [25609]));
Q_ASSIGN U7166 ( .B(clk), .A(\g.we_clk [25608]));
Q_ASSIGN U7167 ( .B(clk), .A(\g.we_clk [25607]));
Q_ASSIGN U7168 ( .B(clk), .A(\g.we_clk [25606]));
Q_ASSIGN U7169 ( .B(clk), .A(\g.we_clk [25605]));
Q_ASSIGN U7170 ( .B(clk), .A(\g.we_clk [25604]));
Q_ASSIGN U7171 ( .B(clk), .A(\g.we_clk [25603]));
Q_ASSIGN U7172 ( .B(clk), .A(\g.we_clk [25602]));
Q_ASSIGN U7173 ( .B(clk), .A(\g.we_clk [25601]));
Q_ASSIGN U7174 ( .B(clk), .A(\g.we_clk [25600]));
Q_ASSIGN U7175 ( .B(clk), .A(\g.we_clk [25599]));
Q_ASSIGN U7176 ( .B(clk), .A(\g.we_clk [25598]));
Q_ASSIGN U7177 ( .B(clk), .A(\g.we_clk [25597]));
Q_ASSIGN U7178 ( .B(clk), .A(\g.we_clk [25596]));
Q_ASSIGN U7179 ( .B(clk), .A(\g.we_clk [25595]));
Q_ASSIGN U7180 ( .B(clk), .A(\g.we_clk [25594]));
Q_ASSIGN U7181 ( .B(clk), .A(\g.we_clk [25593]));
Q_ASSIGN U7182 ( .B(clk), .A(\g.we_clk [25592]));
Q_ASSIGN U7183 ( .B(clk), .A(\g.we_clk [25591]));
Q_ASSIGN U7184 ( .B(clk), .A(\g.we_clk [25590]));
Q_ASSIGN U7185 ( .B(clk), .A(\g.we_clk [25589]));
Q_ASSIGN U7186 ( .B(clk), .A(\g.we_clk [25588]));
Q_ASSIGN U7187 ( .B(clk), .A(\g.we_clk [25587]));
Q_ASSIGN U7188 ( .B(clk), .A(\g.we_clk [25586]));
Q_ASSIGN U7189 ( .B(clk), .A(\g.we_clk [25585]));
Q_ASSIGN U7190 ( .B(clk), .A(\g.we_clk [25584]));
Q_ASSIGN U7191 ( .B(clk), .A(\g.we_clk [25583]));
Q_ASSIGN U7192 ( .B(clk), .A(\g.we_clk [25582]));
Q_ASSIGN U7193 ( .B(clk), .A(\g.we_clk [25581]));
Q_ASSIGN U7194 ( .B(clk), .A(\g.we_clk [25580]));
Q_ASSIGN U7195 ( .B(clk), .A(\g.we_clk [25579]));
Q_ASSIGN U7196 ( .B(clk), .A(\g.we_clk [25578]));
Q_ASSIGN U7197 ( .B(clk), .A(\g.we_clk [25577]));
Q_ASSIGN U7198 ( .B(clk), .A(\g.we_clk [25576]));
Q_ASSIGN U7199 ( .B(clk), .A(\g.we_clk [25575]));
Q_ASSIGN U7200 ( .B(clk), .A(\g.we_clk [25574]));
Q_ASSIGN U7201 ( .B(clk), .A(\g.we_clk [25573]));
Q_ASSIGN U7202 ( .B(clk), .A(\g.we_clk [25572]));
Q_ASSIGN U7203 ( .B(clk), .A(\g.we_clk [25571]));
Q_ASSIGN U7204 ( .B(clk), .A(\g.we_clk [25570]));
Q_ASSIGN U7205 ( .B(clk), .A(\g.we_clk [25569]));
Q_ASSIGN U7206 ( .B(clk), .A(\g.we_clk [25568]));
Q_ASSIGN U7207 ( .B(clk), .A(\g.we_clk [25567]));
Q_ASSIGN U7208 ( .B(clk), .A(\g.we_clk [25566]));
Q_ASSIGN U7209 ( .B(clk), .A(\g.we_clk [25565]));
Q_ASSIGN U7210 ( .B(clk), .A(\g.we_clk [25564]));
Q_ASSIGN U7211 ( .B(clk), .A(\g.we_clk [25563]));
Q_ASSIGN U7212 ( .B(clk), .A(\g.we_clk [25562]));
Q_ASSIGN U7213 ( .B(clk), .A(\g.we_clk [25561]));
Q_ASSIGN U7214 ( .B(clk), .A(\g.we_clk [25560]));
Q_ASSIGN U7215 ( .B(clk), .A(\g.we_clk [25559]));
Q_ASSIGN U7216 ( .B(clk), .A(\g.we_clk [25558]));
Q_ASSIGN U7217 ( .B(clk), .A(\g.we_clk [25557]));
Q_ASSIGN U7218 ( .B(clk), .A(\g.we_clk [25556]));
Q_ASSIGN U7219 ( .B(clk), .A(\g.we_clk [25555]));
Q_ASSIGN U7220 ( .B(clk), .A(\g.we_clk [25554]));
Q_ASSIGN U7221 ( .B(clk), .A(\g.we_clk [25553]));
Q_ASSIGN U7222 ( .B(clk), .A(\g.we_clk [25552]));
Q_ASSIGN U7223 ( .B(clk), .A(\g.we_clk [25551]));
Q_ASSIGN U7224 ( .B(clk), .A(\g.we_clk [25550]));
Q_ASSIGN U7225 ( .B(clk), .A(\g.we_clk [25549]));
Q_ASSIGN U7226 ( .B(clk), .A(\g.we_clk [25548]));
Q_ASSIGN U7227 ( .B(clk), .A(\g.we_clk [25547]));
Q_ASSIGN U7228 ( .B(clk), .A(\g.we_clk [25546]));
Q_ASSIGN U7229 ( .B(clk), .A(\g.we_clk [25545]));
Q_ASSIGN U7230 ( .B(clk), .A(\g.we_clk [25544]));
Q_ASSIGN U7231 ( .B(clk), .A(\g.we_clk [25543]));
Q_ASSIGN U7232 ( .B(clk), .A(\g.we_clk [25542]));
Q_ASSIGN U7233 ( .B(clk), .A(\g.we_clk [25541]));
Q_ASSIGN U7234 ( .B(clk), .A(\g.we_clk [25540]));
Q_ASSIGN U7235 ( .B(clk), .A(\g.we_clk [25539]));
Q_ASSIGN U7236 ( .B(clk), .A(\g.we_clk [25538]));
Q_ASSIGN U7237 ( .B(clk), .A(\g.we_clk [25537]));
Q_ASSIGN U7238 ( .B(clk), .A(\g.we_clk [25536]));
Q_ASSIGN U7239 ( .B(clk), .A(\g.we_clk [25535]));
Q_ASSIGN U7240 ( .B(clk), .A(\g.we_clk [25534]));
Q_ASSIGN U7241 ( .B(clk), .A(\g.we_clk [25533]));
Q_ASSIGN U7242 ( .B(clk), .A(\g.we_clk [25532]));
Q_ASSIGN U7243 ( .B(clk), .A(\g.we_clk [25531]));
Q_ASSIGN U7244 ( .B(clk), .A(\g.we_clk [25530]));
Q_ASSIGN U7245 ( .B(clk), .A(\g.we_clk [25529]));
Q_ASSIGN U7246 ( .B(clk), .A(\g.we_clk [25528]));
Q_ASSIGN U7247 ( .B(clk), .A(\g.we_clk [25527]));
Q_ASSIGN U7248 ( .B(clk), .A(\g.we_clk [25526]));
Q_ASSIGN U7249 ( .B(clk), .A(\g.we_clk [25525]));
Q_ASSIGN U7250 ( .B(clk), .A(\g.we_clk [25524]));
Q_ASSIGN U7251 ( .B(clk), .A(\g.we_clk [25523]));
Q_ASSIGN U7252 ( .B(clk), .A(\g.we_clk [25522]));
Q_ASSIGN U7253 ( .B(clk), .A(\g.we_clk [25521]));
Q_ASSIGN U7254 ( .B(clk), .A(\g.we_clk [25520]));
Q_ASSIGN U7255 ( .B(clk), .A(\g.we_clk [25519]));
Q_ASSIGN U7256 ( .B(clk), .A(\g.we_clk [25518]));
Q_ASSIGN U7257 ( .B(clk), .A(\g.we_clk [25517]));
Q_ASSIGN U7258 ( .B(clk), .A(\g.we_clk [25516]));
Q_ASSIGN U7259 ( .B(clk), .A(\g.we_clk [25515]));
Q_ASSIGN U7260 ( .B(clk), .A(\g.we_clk [25514]));
Q_ASSIGN U7261 ( .B(clk), .A(\g.we_clk [25513]));
Q_ASSIGN U7262 ( .B(clk), .A(\g.we_clk [25512]));
Q_ASSIGN U7263 ( .B(clk), .A(\g.we_clk [25511]));
Q_ASSIGN U7264 ( .B(clk), .A(\g.we_clk [25510]));
Q_ASSIGN U7265 ( .B(clk), .A(\g.we_clk [25509]));
Q_ASSIGN U7266 ( .B(clk), .A(\g.we_clk [25508]));
Q_ASSIGN U7267 ( .B(clk), .A(\g.we_clk [25507]));
Q_ASSIGN U7268 ( .B(clk), .A(\g.we_clk [25506]));
Q_ASSIGN U7269 ( .B(clk), .A(\g.we_clk [25505]));
Q_ASSIGN U7270 ( .B(clk), .A(\g.we_clk [25504]));
Q_ASSIGN U7271 ( .B(clk), .A(\g.we_clk [25503]));
Q_ASSIGN U7272 ( .B(clk), .A(\g.we_clk [25502]));
Q_ASSIGN U7273 ( .B(clk), .A(\g.we_clk [25501]));
Q_ASSIGN U7274 ( .B(clk), .A(\g.we_clk [25500]));
Q_ASSIGN U7275 ( .B(clk), .A(\g.we_clk [25499]));
Q_ASSIGN U7276 ( .B(clk), .A(\g.we_clk [25498]));
Q_ASSIGN U7277 ( .B(clk), .A(\g.we_clk [25497]));
Q_ASSIGN U7278 ( .B(clk), .A(\g.we_clk [25496]));
Q_ASSIGN U7279 ( .B(clk), .A(\g.we_clk [25495]));
Q_ASSIGN U7280 ( .B(clk), .A(\g.we_clk [25494]));
Q_ASSIGN U7281 ( .B(clk), .A(\g.we_clk [25493]));
Q_ASSIGN U7282 ( .B(clk), .A(\g.we_clk [25492]));
Q_ASSIGN U7283 ( .B(clk), .A(\g.we_clk [25491]));
Q_ASSIGN U7284 ( .B(clk), .A(\g.we_clk [25490]));
Q_ASSIGN U7285 ( .B(clk), .A(\g.we_clk [25489]));
Q_ASSIGN U7286 ( .B(clk), .A(\g.we_clk [25488]));
Q_ASSIGN U7287 ( .B(clk), .A(\g.we_clk [25487]));
Q_ASSIGN U7288 ( .B(clk), .A(\g.we_clk [25486]));
Q_ASSIGN U7289 ( .B(clk), .A(\g.we_clk [25485]));
Q_ASSIGN U7290 ( .B(clk), .A(\g.we_clk [25484]));
Q_ASSIGN U7291 ( .B(clk), .A(\g.we_clk [25483]));
Q_ASSIGN U7292 ( .B(clk), .A(\g.we_clk [25482]));
Q_ASSIGN U7293 ( .B(clk), .A(\g.we_clk [25481]));
Q_ASSIGN U7294 ( .B(clk), .A(\g.we_clk [25480]));
Q_ASSIGN U7295 ( .B(clk), .A(\g.we_clk [25479]));
Q_ASSIGN U7296 ( .B(clk), .A(\g.we_clk [25478]));
Q_ASSIGN U7297 ( .B(clk), .A(\g.we_clk [25477]));
Q_ASSIGN U7298 ( .B(clk), .A(\g.we_clk [25476]));
Q_ASSIGN U7299 ( .B(clk), .A(\g.we_clk [25475]));
Q_ASSIGN U7300 ( .B(clk), .A(\g.we_clk [25474]));
Q_ASSIGN U7301 ( .B(clk), .A(\g.we_clk [25473]));
Q_ASSIGN U7302 ( .B(clk), .A(\g.we_clk [25472]));
Q_ASSIGN U7303 ( .B(clk), .A(\g.we_clk [25471]));
Q_ASSIGN U7304 ( .B(clk), .A(\g.we_clk [25470]));
Q_ASSIGN U7305 ( .B(clk), .A(\g.we_clk [25469]));
Q_ASSIGN U7306 ( .B(clk), .A(\g.we_clk [25468]));
Q_ASSIGN U7307 ( .B(clk), .A(\g.we_clk [25467]));
Q_ASSIGN U7308 ( .B(clk), .A(\g.we_clk [25466]));
Q_ASSIGN U7309 ( .B(clk), .A(\g.we_clk [25465]));
Q_ASSIGN U7310 ( .B(clk), .A(\g.we_clk [25464]));
Q_ASSIGN U7311 ( .B(clk), .A(\g.we_clk [25463]));
Q_ASSIGN U7312 ( .B(clk), .A(\g.we_clk [25462]));
Q_ASSIGN U7313 ( .B(clk), .A(\g.we_clk [25461]));
Q_ASSIGN U7314 ( .B(clk), .A(\g.we_clk [25460]));
Q_ASSIGN U7315 ( .B(clk), .A(\g.we_clk [25459]));
Q_ASSIGN U7316 ( .B(clk), .A(\g.we_clk [25458]));
Q_ASSIGN U7317 ( .B(clk), .A(\g.we_clk [25457]));
Q_ASSIGN U7318 ( .B(clk), .A(\g.we_clk [25456]));
Q_ASSIGN U7319 ( .B(clk), .A(\g.we_clk [25455]));
Q_ASSIGN U7320 ( .B(clk), .A(\g.we_clk [25454]));
Q_ASSIGN U7321 ( .B(clk), .A(\g.we_clk [25453]));
Q_ASSIGN U7322 ( .B(clk), .A(\g.we_clk [25452]));
Q_ASSIGN U7323 ( .B(clk), .A(\g.we_clk [25451]));
Q_ASSIGN U7324 ( .B(clk), .A(\g.we_clk [25450]));
Q_ASSIGN U7325 ( .B(clk), .A(\g.we_clk [25449]));
Q_ASSIGN U7326 ( .B(clk), .A(\g.we_clk [25448]));
Q_ASSIGN U7327 ( .B(clk), .A(\g.we_clk [25447]));
Q_ASSIGN U7328 ( .B(clk), .A(\g.we_clk [25446]));
Q_ASSIGN U7329 ( .B(clk), .A(\g.we_clk [25445]));
Q_ASSIGN U7330 ( .B(clk), .A(\g.we_clk [25444]));
Q_ASSIGN U7331 ( .B(clk), .A(\g.we_clk [25443]));
Q_ASSIGN U7332 ( .B(clk), .A(\g.we_clk [25442]));
Q_ASSIGN U7333 ( .B(clk), .A(\g.we_clk [25441]));
Q_ASSIGN U7334 ( .B(clk), .A(\g.we_clk [25440]));
Q_ASSIGN U7335 ( .B(clk), .A(\g.we_clk [25439]));
Q_ASSIGN U7336 ( .B(clk), .A(\g.we_clk [25438]));
Q_ASSIGN U7337 ( .B(clk), .A(\g.we_clk [25437]));
Q_ASSIGN U7338 ( .B(clk), .A(\g.we_clk [25436]));
Q_ASSIGN U7339 ( .B(clk), .A(\g.we_clk [25435]));
Q_ASSIGN U7340 ( .B(clk), .A(\g.we_clk [25434]));
Q_ASSIGN U7341 ( .B(clk), .A(\g.we_clk [25433]));
Q_ASSIGN U7342 ( .B(clk), .A(\g.we_clk [25432]));
Q_ASSIGN U7343 ( .B(clk), .A(\g.we_clk [25431]));
Q_ASSIGN U7344 ( .B(clk), .A(\g.we_clk [25430]));
Q_ASSIGN U7345 ( .B(clk), .A(\g.we_clk [25429]));
Q_ASSIGN U7346 ( .B(clk), .A(\g.we_clk [25428]));
Q_ASSIGN U7347 ( .B(clk), .A(\g.we_clk [25427]));
Q_ASSIGN U7348 ( .B(clk), .A(\g.we_clk [25426]));
Q_ASSIGN U7349 ( .B(clk), .A(\g.we_clk [25425]));
Q_ASSIGN U7350 ( .B(clk), .A(\g.we_clk [25424]));
Q_ASSIGN U7351 ( .B(clk), .A(\g.we_clk [25423]));
Q_ASSIGN U7352 ( .B(clk), .A(\g.we_clk [25422]));
Q_ASSIGN U7353 ( .B(clk), .A(\g.we_clk [25421]));
Q_ASSIGN U7354 ( .B(clk), .A(\g.we_clk [25420]));
Q_ASSIGN U7355 ( .B(clk), .A(\g.we_clk [25419]));
Q_ASSIGN U7356 ( .B(clk), .A(\g.we_clk [25418]));
Q_ASSIGN U7357 ( .B(clk), .A(\g.we_clk [25417]));
Q_ASSIGN U7358 ( .B(clk), .A(\g.we_clk [25416]));
Q_ASSIGN U7359 ( .B(clk), .A(\g.we_clk [25415]));
Q_ASSIGN U7360 ( .B(clk), .A(\g.we_clk [25414]));
Q_ASSIGN U7361 ( .B(clk), .A(\g.we_clk [25413]));
Q_ASSIGN U7362 ( .B(clk), .A(\g.we_clk [25412]));
Q_ASSIGN U7363 ( .B(clk), .A(\g.we_clk [25411]));
Q_ASSIGN U7364 ( .B(clk), .A(\g.we_clk [25410]));
Q_ASSIGN U7365 ( .B(clk), .A(\g.we_clk [25409]));
Q_ASSIGN U7366 ( .B(clk), .A(\g.we_clk [25408]));
Q_ASSIGN U7367 ( .B(clk), .A(\g.we_clk [25407]));
Q_ASSIGN U7368 ( .B(clk), .A(\g.we_clk [25406]));
Q_ASSIGN U7369 ( .B(clk), .A(\g.we_clk [25405]));
Q_ASSIGN U7370 ( .B(clk), .A(\g.we_clk [25404]));
Q_ASSIGN U7371 ( .B(clk), .A(\g.we_clk [25403]));
Q_ASSIGN U7372 ( .B(clk), .A(\g.we_clk [25402]));
Q_ASSIGN U7373 ( .B(clk), .A(\g.we_clk [25401]));
Q_ASSIGN U7374 ( .B(clk), .A(\g.we_clk [25400]));
Q_ASSIGN U7375 ( .B(clk), .A(\g.we_clk [25399]));
Q_ASSIGN U7376 ( .B(clk), .A(\g.we_clk [25398]));
Q_ASSIGN U7377 ( .B(clk), .A(\g.we_clk [25397]));
Q_ASSIGN U7378 ( .B(clk), .A(\g.we_clk [25396]));
Q_ASSIGN U7379 ( .B(clk), .A(\g.we_clk [25395]));
Q_ASSIGN U7380 ( .B(clk), .A(\g.we_clk [25394]));
Q_ASSIGN U7381 ( .B(clk), .A(\g.we_clk [25393]));
Q_ASSIGN U7382 ( .B(clk), .A(\g.we_clk [25392]));
Q_ASSIGN U7383 ( .B(clk), .A(\g.we_clk [25391]));
Q_ASSIGN U7384 ( .B(clk), .A(\g.we_clk [25390]));
Q_ASSIGN U7385 ( .B(clk), .A(\g.we_clk [25389]));
Q_ASSIGN U7386 ( .B(clk), .A(\g.we_clk [25388]));
Q_ASSIGN U7387 ( .B(clk), .A(\g.we_clk [25387]));
Q_ASSIGN U7388 ( .B(clk), .A(\g.we_clk [25386]));
Q_ASSIGN U7389 ( .B(clk), .A(\g.we_clk [25385]));
Q_ASSIGN U7390 ( .B(clk), .A(\g.we_clk [25384]));
Q_ASSIGN U7391 ( .B(clk), .A(\g.we_clk [25383]));
Q_ASSIGN U7392 ( .B(clk), .A(\g.we_clk [25382]));
Q_ASSIGN U7393 ( .B(clk), .A(\g.we_clk [25381]));
Q_ASSIGN U7394 ( .B(clk), .A(\g.we_clk [25380]));
Q_ASSIGN U7395 ( .B(clk), .A(\g.we_clk [25379]));
Q_ASSIGN U7396 ( .B(clk), .A(\g.we_clk [25378]));
Q_ASSIGN U7397 ( .B(clk), .A(\g.we_clk [25377]));
Q_ASSIGN U7398 ( .B(clk), .A(\g.we_clk [25376]));
Q_ASSIGN U7399 ( .B(clk), .A(\g.we_clk [25375]));
Q_ASSIGN U7400 ( .B(clk), .A(\g.we_clk [25374]));
Q_ASSIGN U7401 ( .B(clk), .A(\g.we_clk [25373]));
Q_ASSIGN U7402 ( .B(clk), .A(\g.we_clk [25372]));
Q_ASSIGN U7403 ( .B(clk), .A(\g.we_clk [25371]));
Q_ASSIGN U7404 ( .B(clk), .A(\g.we_clk [25370]));
Q_ASSIGN U7405 ( .B(clk), .A(\g.we_clk [25369]));
Q_ASSIGN U7406 ( .B(clk), .A(\g.we_clk [25368]));
Q_ASSIGN U7407 ( .B(clk), .A(\g.we_clk [25367]));
Q_ASSIGN U7408 ( .B(clk), .A(\g.we_clk [25366]));
Q_ASSIGN U7409 ( .B(clk), .A(\g.we_clk [25365]));
Q_ASSIGN U7410 ( .B(clk), .A(\g.we_clk [25364]));
Q_ASSIGN U7411 ( .B(clk), .A(\g.we_clk [25363]));
Q_ASSIGN U7412 ( .B(clk), .A(\g.we_clk [25362]));
Q_ASSIGN U7413 ( .B(clk), .A(\g.we_clk [25361]));
Q_ASSIGN U7414 ( .B(clk), .A(\g.we_clk [25360]));
Q_ASSIGN U7415 ( .B(clk), .A(\g.we_clk [25359]));
Q_ASSIGN U7416 ( .B(clk), .A(\g.we_clk [25358]));
Q_ASSIGN U7417 ( .B(clk), .A(\g.we_clk [25357]));
Q_ASSIGN U7418 ( .B(clk), .A(\g.we_clk [25356]));
Q_ASSIGN U7419 ( .B(clk), .A(\g.we_clk [25355]));
Q_ASSIGN U7420 ( .B(clk), .A(\g.we_clk [25354]));
Q_ASSIGN U7421 ( .B(clk), .A(\g.we_clk [25353]));
Q_ASSIGN U7422 ( .B(clk), .A(\g.we_clk [25352]));
Q_ASSIGN U7423 ( .B(clk), .A(\g.we_clk [25351]));
Q_ASSIGN U7424 ( .B(clk), .A(\g.we_clk [25350]));
Q_ASSIGN U7425 ( .B(clk), .A(\g.we_clk [25349]));
Q_ASSIGN U7426 ( .B(clk), .A(\g.we_clk [25348]));
Q_ASSIGN U7427 ( .B(clk), .A(\g.we_clk [25347]));
Q_ASSIGN U7428 ( .B(clk), .A(\g.we_clk [25346]));
Q_ASSIGN U7429 ( .B(clk), .A(\g.we_clk [25345]));
Q_ASSIGN U7430 ( .B(clk), .A(\g.we_clk [25344]));
Q_ASSIGN U7431 ( .B(clk), .A(\g.we_clk [25343]));
Q_ASSIGN U7432 ( .B(clk), .A(\g.we_clk [25342]));
Q_ASSIGN U7433 ( .B(clk), .A(\g.we_clk [25341]));
Q_ASSIGN U7434 ( .B(clk), .A(\g.we_clk [25340]));
Q_ASSIGN U7435 ( .B(clk), .A(\g.we_clk [25339]));
Q_ASSIGN U7436 ( .B(clk), .A(\g.we_clk [25338]));
Q_ASSIGN U7437 ( .B(clk), .A(\g.we_clk [25337]));
Q_ASSIGN U7438 ( .B(clk), .A(\g.we_clk [25336]));
Q_ASSIGN U7439 ( .B(clk), .A(\g.we_clk [25335]));
Q_ASSIGN U7440 ( .B(clk), .A(\g.we_clk [25334]));
Q_ASSIGN U7441 ( .B(clk), .A(\g.we_clk [25333]));
Q_ASSIGN U7442 ( .B(clk), .A(\g.we_clk [25332]));
Q_ASSIGN U7443 ( .B(clk), .A(\g.we_clk [25331]));
Q_ASSIGN U7444 ( .B(clk), .A(\g.we_clk [25330]));
Q_ASSIGN U7445 ( .B(clk), .A(\g.we_clk [25329]));
Q_ASSIGN U7446 ( .B(clk), .A(\g.we_clk [25328]));
Q_ASSIGN U7447 ( .B(clk), .A(\g.we_clk [25327]));
Q_ASSIGN U7448 ( .B(clk), .A(\g.we_clk [25326]));
Q_ASSIGN U7449 ( .B(clk), .A(\g.we_clk [25325]));
Q_ASSIGN U7450 ( .B(clk), .A(\g.we_clk [25324]));
Q_ASSIGN U7451 ( .B(clk), .A(\g.we_clk [25323]));
Q_ASSIGN U7452 ( .B(clk), .A(\g.we_clk [25322]));
Q_ASSIGN U7453 ( .B(clk), .A(\g.we_clk [25321]));
Q_ASSIGN U7454 ( .B(clk), .A(\g.we_clk [25320]));
Q_ASSIGN U7455 ( .B(clk), .A(\g.we_clk [25319]));
Q_ASSIGN U7456 ( .B(clk), .A(\g.we_clk [25318]));
Q_ASSIGN U7457 ( .B(clk), .A(\g.we_clk [25317]));
Q_ASSIGN U7458 ( .B(clk), .A(\g.we_clk [25316]));
Q_ASSIGN U7459 ( .B(clk), .A(\g.we_clk [25315]));
Q_ASSIGN U7460 ( .B(clk), .A(\g.we_clk [25314]));
Q_ASSIGN U7461 ( .B(clk), .A(\g.we_clk [25313]));
Q_ASSIGN U7462 ( .B(clk), .A(\g.we_clk [25312]));
Q_ASSIGN U7463 ( .B(clk), .A(\g.we_clk [25311]));
Q_ASSIGN U7464 ( .B(clk), .A(\g.we_clk [25310]));
Q_ASSIGN U7465 ( .B(clk), .A(\g.we_clk [25309]));
Q_ASSIGN U7466 ( .B(clk), .A(\g.we_clk [25308]));
Q_ASSIGN U7467 ( .B(clk), .A(\g.we_clk [25307]));
Q_ASSIGN U7468 ( .B(clk), .A(\g.we_clk [25306]));
Q_ASSIGN U7469 ( .B(clk), .A(\g.we_clk [25305]));
Q_ASSIGN U7470 ( .B(clk), .A(\g.we_clk [25304]));
Q_ASSIGN U7471 ( .B(clk), .A(\g.we_clk [25303]));
Q_ASSIGN U7472 ( .B(clk), .A(\g.we_clk [25302]));
Q_ASSIGN U7473 ( .B(clk), .A(\g.we_clk [25301]));
Q_ASSIGN U7474 ( .B(clk), .A(\g.we_clk [25300]));
Q_ASSIGN U7475 ( .B(clk), .A(\g.we_clk [25299]));
Q_ASSIGN U7476 ( .B(clk), .A(\g.we_clk [25298]));
Q_ASSIGN U7477 ( .B(clk), .A(\g.we_clk [25297]));
Q_ASSIGN U7478 ( .B(clk), .A(\g.we_clk [25296]));
Q_ASSIGN U7479 ( .B(clk), .A(\g.we_clk [25295]));
Q_ASSIGN U7480 ( .B(clk), .A(\g.we_clk [25294]));
Q_ASSIGN U7481 ( .B(clk), .A(\g.we_clk [25293]));
Q_ASSIGN U7482 ( .B(clk), .A(\g.we_clk [25292]));
Q_ASSIGN U7483 ( .B(clk), .A(\g.we_clk [25291]));
Q_ASSIGN U7484 ( .B(clk), .A(\g.we_clk [25290]));
Q_ASSIGN U7485 ( .B(clk), .A(\g.we_clk [25289]));
Q_ASSIGN U7486 ( .B(clk), .A(\g.we_clk [25288]));
Q_ASSIGN U7487 ( .B(clk), .A(\g.we_clk [25287]));
Q_ASSIGN U7488 ( .B(clk), .A(\g.we_clk [25286]));
Q_ASSIGN U7489 ( .B(clk), .A(\g.we_clk [25285]));
Q_ASSIGN U7490 ( .B(clk), .A(\g.we_clk [25284]));
Q_ASSIGN U7491 ( .B(clk), .A(\g.we_clk [25283]));
Q_ASSIGN U7492 ( .B(clk), .A(\g.we_clk [25282]));
Q_ASSIGN U7493 ( .B(clk), .A(\g.we_clk [25281]));
Q_ASSIGN U7494 ( .B(clk), .A(\g.we_clk [25280]));
Q_ASSIGN U7495 ( .B(clk), .A(\g.we_clk [25279]));
Q_ASSIGN U7496 ( .B(clk), .A(\g.we_clk [25278]));
Q_ASSIGN U7497 ( .B(clk), .A(\g.we_clk [25277]));
Q_ASSIGN U7498 ( .B(clk), .A(\g.we_clk [25276]));
Q_ASSIGN U7499 ( .B(clk), .A(\g.we_clk [25275]));
Q_ASSIGN U7500 ( .B(clk), .A(\g.we_clk [25274]));
Q_ASSIGN U7501 ( .B(clk), .A(\g.we_clk [25273]));
Q_ASSIGN U7502 ( .B(clk), .A(\g.we_clk [25272]));
Q_ASSIGN U7503 ( .B(clk), .A(\g.we_clk [25271]));
Q_ASSIGN U7504 ( .B(clk), .A(\g.we_clk [25270]));
Q_ASSIGN U7505 ( .B(clk), .A(\g.we_clk [25269]));
Q_ASSIGN U7506 ( .B(clk), .A(\g.we_clk [25268]));
Q_ASSIGN U7507 ( .B(clk), .A(\g.we_clk [25267]));
Q_ASSIGN U7508 ( .B(clk), .A(\g.we_clk [25266]));
Q_ASSIGN U7509 ( .B(clk), .A(\g.we_clk [25265]));
Q_ASSIGN U7510 ( .B(clk), .A(\g.we_clk [25264]));
Q_ASSIGN U7511 ( .B(clk), .A(\g.we_clk [25263]));
Q_ASSIGN U7512 ( .B(clk), .A(\g.we_clk [25262]));
Q_ASSIGN U7513 ( .B(clk), .A(\g.we_clk [25261]));
Q_ASSIGN U7514 ( .B(clk), .A(\g.we_clk [25260]));
Q_ASSIGN U7515 ( .B(clk), .A(\g.we_clk [25259]));
Q_ASSIGN U7516 ( .B(clk), .A(\g.we_clk [25258]));
Q_ASSIGN U7517 ( .B(clk), .A(\g.we_clk [25257]));
Q_ASSIGN U7518 ( .B(clk), .A(\g.we_clk [25256]));
Q_ASSIGN U7519 ( .B(clk), .A(\g.we_clk [25255]));
Q_ASSIGN U7520 ( .B(clk), .A(\g.we_clk [25254]));
Q_ASSIGN U7521 ( .B(clk), .A(\g.we_clk [25253]));
Q_ASSIGN U7522 ( .B(clk), .A(\g.we_clk [25252]));
Q_ASSIGN U7523 ( .B(clk), .A(\g.we_clk [25251]));
Q_ASSIGN U7524 ( .B(clk), .A(\g.we_clk [25250]));
Q_ASSIGN U7525 ( .B(clk), .A(\g.we_clk [25249]));
Q_ASSIGN U7526 ( .B(clk), .A(\g.we_clk [25248]));
Q_ASSIGN U7527 ( .B(clk), .A(\g.we_clk [25247]));
Q_ASSIGN U7528 ( .B(clk), .A(\g.we_clk [25246]));
Q_ASSIGN U7529 ( .B(clk), .A(\g.we_clk [25245]));
Q_ASSIGN U7530 ( .B(clk), .A(\g.we_clk [25244]));
Q_ASSIGN U7531 ( .B(clk), .A(\g.we_clk [25243]));
Q_ASSIGN U7532 ( .B(clk), .A(\g.we_clk [25242]));
Q_ASSIGN U7533 ( .B(clk), .A(\g.we_clk [25241]));
Q_ASSIGN U7534 ( .B(clk), .A(\g.we_clk [25240]));
Q_ASSIGN U7535 ( .B(clk), .A(\g.we_clk [25239]));
Q_ASSIGN U7536 ( .B(clk), .A(\g.we_clk [25238]));
Q_ASSIGN U7537 ( .B(clk), .A(\g.we_clk [25237]));
Q_ASSIGN U7538 ( .B(clk), .A(\g.we_clk [25236]));
Q_ASSIGN U7539 ( .B(clk), .A(\g.we_clk [25235]));
Q_ASSIGN U7540 ( .B(clk), .A(\g.we_clk [25234]));
Q_ASSIGN U7541 ( .B(clk), .A(\g.we_clk [25233]));
Q_ASSIGN U7542 ( .B(clk), .A(\g.we_clk [25232]));
Q_ASSIGN U7543 ( .B(clk), .A(\g.we_clk [25231]));
Q_ASSIGN U7544 ( .B(clk), .A(\g.we_clk [25230]));
Q_ASSIGN U7545 ( .B(clk), .A(\g.we_clk [25229]));
Q_ASSIGN U7546 ( .B(clk), .A(\g.we_clk [25228]));
Q_ASSIGN U7547 ( .B(clk), .A(\g.we_clk [25227]));
Q_ASSIGN U7548 ( .B(clk), .A(\g.we_clk [25226]));
Q_ASSIGN U7549 ( .B(clk), .A(\g.we_clk [25225]));
Q_ASSIGN U7550 ( .B(clk), .A(\g.we_clk [25224]));
Q_ASSIGN U7551 ( .B(clk), .A(\g.we_clk [25223]));
Q_ASSIGN U7552 ( .B(clk), .A(\g.we_clk [25222]));
Q_ASSIGN U7553 ( .B(clk), .A(\g.we_clk [25221]));
Q_ASSIGN U7554 ( .B(clk), .A(\g.we_clk [25220]));
Q_ASSIGN U7555 ( .B(clk), .A(\g.we_clk [25219]));
Q_ASSIGN U7556 ( .B(clk), .A(\g.we_clk [25218]));
Q_ASSIGN U7557 ( .B(clk), .A(\g.we_clk [25217]));
Q_ASSIGN U7558 ( .B(clk), .A(\g.we_clk [25216]));
Q_ASSIGN U7559 ( .B(clk), .A(\g.we_clk [25215]));
Q_ASSIGN U7560 ( .B(clk), .A(\g.we_clk [25214]));
Q_ASSIGN U7561 ( .B(clk), .A(\g.we_clk [25213]));
Q_ASSIGN U7562 ( .B(clk), .A(\g.we_clk [25212]));
Q_ASSIGN U7563 ( .B(clk), .A(\g.we_clk [25211]));
Q_ASSIGN U7564 ( .B(clk), .A(\g.we_clk [25210]));
Q_ASSIGN U7565 ( .B(clk), .A(\g.we_clk [25209]));
Q_ASSIGN U7566 ( .B(clk), .A(\g.we_clk [25208]));
Q_ASSIGN U7567 ( .B(clk), .A(\g.we_clk [25207]));
Q_ASSIGN U7568 ( .B(clk), .A(\g.we_clk [25206]));
Q_ASSIGN U7569 ( .B(clk), .A(\g.we_clk [25205]));
Q_ASSIGN U7570 ( .B(clk), .A(\g.we_clk [25204]));
Q_ASSIGN U7571 ( .B(clk), .A(\g.we_clk [25203]));
Q_ASSIGN U7572 ( .B(clk), .A(\g.we_clk [25202]));
Q_ASSIGN U7573 ( .B(clk), .A(\g.we_clk [25201]));
Q_ASSIGN U7574 ( .B(clk), .A(\g.we_clk [25200]));
Q_ASSIGN U7575 ( .B(clk), .A(\g.we_clk [25199]));
Q_ASSIGN U7576 ( .B(clk), .A(\g.we_clk [25198]));
Q_ASSIGN U7577 ( .B(clk), .A(\g.we_clk [25197]));
Q_ASSIGN U7578 ( .B(clk), .A(\g.we_clk [25196]));
Q_ASSIGN U7579 ( .B(clk), .A(\g.we_clk [25195]));
Q_ASSIGN U7580 ( .B(clk), .A(\g.we_clk [25194]));
Q_ASSIGN U7581 ( .B(clk), .A(\g.we_clk [25193]));
Q_ASSIGN U7582 ( .B(clk), .A(\g.we_clk [25192]));
Q_ASSIGN U7583 ( .B(clk), .A(\g.we_clk [25191]));
Q_ASSIGN U7584 ( .B(clk), .A(\g.we_clk [25190]));
Q_ASSIGN U7585 ( .B(clk), .A(\g.we_clk [25189]));
Q_ASSIGN U7586 ( .B(clk), .A(\g.we_clk [25188]));
Q_ASSIGN U7587 ( .B(clk), .A(\g.we_clk [25187]));
Q_ASSIGN U7588 ( .B(clk), .A(\g.we_clk [25186]));
Q_ASSIGN U7589 ( .B(clk), .A(\g.we_clk [25185]));
Q_ASSIGN U7590 ( .B(clk), .A(\g.we_clk [25184]));
Q_ASSIGN U7591 ( .B(clk), .A(\g.we_clk [25183]));
Q_ASSIGN U7592 ( .B(clk), .A(\g.we_clk [25182]));
Q_ASSIGN U7593 ( .B(clk), .A(\g.we_clk [25181]));
Q_ASSIGN U7594 ( .B(clk), .A(\g.we_clk [25180]));
Q_ASSIGN U7595 ( .B(clk), .A(\g.we_clk [25179]));
Q_ASSIGN U7596 ( .B(clk), .A(\g.we_clk [25178]));
Q_ASSIGN U7597 ( .B(clk), .A(\g.we_clk [25177]));
Q_ASSIGN U7598 ( .B(clk), .A(\g.we_clk [25176]));
Q_ASSIGN U7599 ( .B(clk), .A(\g.we_clk [25175]));
Q_ASSIGN U7600 ( .B(clk), .A(\g.we_clk [25174]));
Q_ASSIGN U7601 ( .B(clk), .A(\g.we_clk [25173]));
Q_ASSIGN U7602 ( .B(clk), .A(\g.we_clk [25172]));
Q_ASSIGN U7603 ( .B(clk), .A(\g.we_clk [25171]));
Q_ASSIGN U7604 ( .B(clk), .A(\g.we_clk [25170]));
Q_ASSIGN U7605 ( .B(clk), .A(\g.we_clk [25169]));
Q_ASSIGN U7606 ( .B(clk), .A(\g.we_clk [25168]));
Q_ASSIGN U7607 ( .B(clk), .A(\g.we_clk [25167]));
Q_ASSIGN U7608 ( .B(clk), .A(\g.we_clk [25166]));
Q_ASSIGN U7609 ( .B(clk), .A(\g.we_clk [25165]));
Q_ASSIGN U7610 ( .B(clk), .A(\g.we_clk [25164]));
Q_ASSIGN U7611 ( .B(clk), .A(\g.we_clk [25163]));
Q_ASSIGN U7612 ( .B(clk), .A(\g.we_clk [25162]));
Q_ASSIGN U7613 ( .B(clk), .A(\g.we_clk [25161]));
Q_ASSIGN U7614 ( .B(clk), .A(\g.we_clk [25160]));
Q_ASSIGN U7615 ( .B(clk), .A(\g.we_clk [25159]));
Q_ASSIGN U7616 ( .B(clk), .A(\g.we_clk [25158]));
Q_ASSIGN U7617 ( .B(clk), .A(\g.we_clk [25157]));
Q_ASSIGN U7618 ( .B(clk), .A(\g.we_clk [25156]));
Q_ASSIGN U7619 ( .B(clk), .A(\g.we_clk [25155]));
Q_ASSIGN U7620 ( .B(clk), .A(\g.we_clk [25154]));
Q_ASSIGN U7621 ( .B(clk), .A(\g.we_clk [25153]));
Q_ASSIGN U7622 ( .B(clk), .A(\g.we_clk [25152]));
Q_ASSIGN U7623 ( .B(clk), .A(\g.we_clk [25151]));
Q_ASSIGN U7624 ( .B(clk), .A(\g.we_clk [25150]));
Q_ASSIGN U7625 ( .B(clk), .A(\g.we_clk [25149]));
Q_ASSIGN U7626 ( .B(clk), .A(\g.we_clk [25148]));
Q_ASSIGN U7627 ( .B(clk), .A(\g.we_clk [25147]));
Q_ASSIGN U7628 ( .B(clk), .A(\g.we_clk [25146]));
Q_ASSIGN U7629 ( .B(clk), .A(\g.we_clk [25145]));
Q_ASSIGN U7630 ( .B(clk), .A(\g.we_clk [25144]));
Q_ASSIGN U7631 ( .B(clk), .A(\g.we_clk [25143]));
Q_ASSIGN U7632 ( .B(clk), .A(\g.we_clk [25142]));
Q_ASSIGN U7633 ( .B(clk), .A(\g.we_clk [25141]));
Q_ASSIGN U7634 ( .B(clk), .A(\g.we_clk [25140]));
Q_ASSIGN U7635 ( .B(clk), .A(\g.we_clk [25139]));
Q_ASSIGN U7636 ( .B(clk), .A(\g.we_clk [25138]));
Q_ASSIGN U7637 ( .B(clk), .A(\g.we_clk [25137]));
Q_ASSIGN U7638 ( .B(clk), .A(\g.we_clk [25136]));
Q_ASSIGN U7639 ( .B(clk), .A(\g.we_clk [25135]));
Q_ASSIGN U7640 ( .B(clk), .A(\g.we_clk [25134]));
Q_ASSIGN U7641 ( .B(clk), .A(\g.we_clk [25133]));
Q_ASSIGN U7642 ( .B(clk), .A(\g.we_clk [25132]));
Q_ASSIGN U7643 ( .B(clk), .A(\g.we_clk [25131]));
Q_ASSIGN U7644 ( .B(clk), .A(\g.we_clk [25130]));
Q_ASSIGN U7645 ( .B(clk), .A(\g.we_clk [25129]));
Q_ASSIGN U7646 ( .B(clk), .A(\g.we_clk [25128]));
Q_ASSIGN U7647 ( .B(clk), .A(\g.we_clk [25127]));
Q_ASSIGN U7648 ( .B(clk), .A(\g.we_clk [25126]));
Q_ASSIGN U7649 ( .B(clk), .A(\g.we_clk [25125]));
Q_ASSIGN U7650 ( .B(clk), .A(\g.we_clk [25124]));
Q_ASSIGN U7651 ( .B(clk), .A(\g.we_clk [25123]));
Q_ASSIGN U7652 ( .B(clk), .A(\g.we_clk [25122]));
Q_ASSIGN U7653 ( .B(clk), .A(\g.we_clk [25121]));
Q_ASSIGN U7654 ( .B(clk), .A(\g.we_clk [25120]));
Q_ASSIGN U7655 ( .B(clk), .A(\g.we_clk [25119]));
Q_ASSIGN U7656 ( .B(clk), .A(\g.we_clk [25118]));
Q_ASSIGN U7657 ( .B(clk), .A(\g.we_clk [25117]));
Q_ASSIGN U7658 ( .B(clk), .A(\g.we_clk [25116]));
Q_ASSIGN U7659 ( .B(clk), .A(\g.we_clk [25115]));
Q_ASSIGN U7660 ( .B(clk), .A(\g.we_clk [25114]));
Q_ASSIGN U7661 ( .B(clk), .A(\g.we_clk [25113]));
Q_ASSIGN U7662 ( .B(clk), .A(\g.we_clk [25112]));
Q_ASSIGN U7663 ( .B(clk), .A(\g.we_clk [25111]));
Q_ASSIGN U7664 ( .B(clk), .A(\g.we_clk [25110]));
Q_ASSIGN U7665 ( .B(clk), .A(\g.we_clk [25109]));
Q_ASSIGN U7666 ( .B(clk), .A(\g.we_clk [25108]));
Q_ASSIGN U7667 ( .B(clk), .A(\g.we_clk [25107]));
Q_ASSIGN U7668 ( .B(clk), .A(\g.we_clk [25106]));
Q_ASSIGN U7669 ( .B(clk), .A(\g.we_clk [25105]));
Q_ASSIGN U7670 ( .B(clk), .A(\g.we_clk [25104]));
Q_ASSIGN U7671 ( .B(clk), .A(\g.we_clk [25103]));
Q_ASSIGN U7672 ( .B(clk), .A(\g.we_clk [25102]));
Q_ASSIGN U7673 ( .B(clk), .A(\g.we_clk [25101]));
Q_ASSIGN U7674 ( .B(clk), .A(\g.we_clk [25100]));
Q_ASSIGN U7675 ( .B(clk), .A(\g.we_clk [25099]));
Q_ASSIGN U7676 ( .B(clk), .A(\g.we_clk [25098]));
Q_ASSIGN U7677 ( .B(clk), .A(\g.we_clk [25097]));
Q_ASSIGN U7678 ( .B(clk), .A(\g.we_clk [25096]));
Q_ASSIGN U7679 ( .B(clk), .A(\g.we_clk [25095]));
Q_ASSIGN U7680 ( .B(clk), .A(\g.we_clk [25094]));
Q_ASSIGN U7681 ( .B(clk), .A(\g.we_clk [25093]));
Q_ASSIGN U7682 ( .B(clk), .A(\g.we_clk [25092]));
Q_ASSIGN U7683 ( .B(clk), .A(\g.we_clk [25091]));
Q_ASSIGN U7684 ( .B(clk), .A(\g.we_clk [25090]));
Q_ASSIGN U7685 ( .B(clk), .A(\g.we_clk [25089]));
Q_ASSIGN U7686 ( .B(clk), .A(\g.we_clk [25088]));
Q_ASSIGN U7687 ( .B(clk), .A(\g.we_clk [25087]));
Q_ASSIGN U7688 ( .B(clk), .A(\g.we_clk [25086]));
Q_ASSIGN U7689 ( .B(clk), .A(\g.we_clk [25085]));
Q_ASSIGN U7690 ( .B(clk), .A(\g.we_clk [25084]));
Q_ASSIGN U7691 ( .B(clk), .A(\g.we_clk [25083]));
Q_ASSIGN U7692 ( .B(clk), .A(\g.we_clk [25082]));
Q_ASSIGN U7693 ( .B(clk), .A(\g.we_clk [25081]));
Q_ASSIGN U7694 ( .B(clk), .A(\g.we_clk [25080]));
Q_ASSIGN U7695 ( .B(clk), .A(\g.we_clk [25079]));
Q_ASSIGN U7696 ( .B(clk), .A(\g.we_clk [25078]));
Q_ASSIGN U7697 ( .B(clk), .A(\g.we_clk [25077]));
Q_ASSIGN U7698 ( .B(clk), .A(\g.we_clk [25076]));
Q_ASSIGN U7699 ( .B(clk), .A(\g.we_clk [25075]));
Q_ASSIGN U7700 ( .B(clk), .A(\g.we_clk [25074]));
Q_ASSIGN U7701 ( .B(clk), .A(\g.we_clk [25073]));
Q_ASSIGN U7702 ( .B(clk), .A(\g.we_clk [25072]));
Q_ASSIGN U7703 ( .B(clk), .A(\g.we_clk [25071]));
Q_ASSIGN U7704 ( .B(clk), .A(\g.we_clk [25070]));
Q_ASSIGN U7705 ( .B(clk), .A(\g.we_clk [25069]));
Q_ASSIGN U7706 ( .B(clk), .A(\g.we_clk [25068]));
Q_ASSIGN U7707 ( .B(clk), .A(\g.we_clk [25067]));
Q_ASSIGN U7708 ( .B(clk), .A(\g.we_clk [25066]));
Q_ASSIGN U7709 ( .B(clk), .A(\g.we_clk [25065]));
Q_ASSIGN U7710 ( .B(clk), .A(\g.we_clk [25064]));
Q_ASSIGN U7711 ( .B(clk), .A(\g.we_clk [25063]));
Q_ASSIGN U7712 ( .B(clk), .A(\g.we_clk [25062]));
Q_ASSIGN U7713 ( .B(clk), .A(\g.we_clk [25061]));
Q_ASSIGN U7714 ( .B(clk), .A(\g.we_clk [25060]));
Q_ASSIGN U7715 ( .B(clk), .A(\g.we_clk [25059]));
Q_ASSIGN U7716 ( .B(clk), .A(\g.we_clk [25058]));
Q_ASSIGN U7717 ( .B(clk), .A(\g.we_clk [25057]));
Q_ASSIGN U7718 ( .B(clk), .A(\g.we_clk [25056]));
Q_ASSIGN U7719 ( .B(clk), .A(\g.we_clk [25055]));
Q_ASSIGN U7720 ( .B(clk), .A(\g.we_clk [25054]));
Q_ASSIGN U7721 ( .B(clk), .A(\g.we_clk [25053]));
Q_ASSIGN U7722 ( .B(clk), .A(\g.we_clk [25052]));
Q_ASSIGN U7723 ( .B(clk), .A(\g.we_clk [25051]));
Q_ASSIGN U7724 ( .B(clk), .A(\g.we_clk [25050]));
Q_ASSIGN U7725 ( .B(clk), .A(\g.we_clk [25049]));
Q_ASSIGN U7726 ( .B(clk), .A(\g.we_clk [25048]));
Q_ASSIGN U7727 ( .B(clk), .A(\g.we_clk [25047]));
Q_ASSIGN U7728 ( .B(clk), .A(\g.we_clk [25046]));
Q_ASSIGN U7729 ( .B(clk), .A(\g.we_clk [25045]));
Q_ASSIGN U7730 ( .B(clk), .A(\g.we_clk [25044]));
Q_ASSIGN U7731 ( .B(clk), .A(\g.we_clk [25043]));
Q_ASSIGN U7732 ( .B(clk), .A(\g.we_clk [25042]));
Q_ASSIGN U7733 ( .B(clk), .A(\g.we_clk [25041]));
Q_ASSIGN U7734 ( .B(clk), .A(\g.we_clk [25040]));
Q_ASSIGN U7735 ( .B(clk), .A(\g.we_clk [25039]));
Q_ASSIGN U7736 ( .B(clk), .A(\g.we_clk [25038]));
Q_ASSIGN U7737 ( .B(clk), .A(\g.we_clk [25037]));
Q_ASSIGN U7738 ( .B(clk), .A(\g.we_clk [25036]));
Q_ASSIGN U7739 ( .B(clk), .A(\g.we_clk [25035]));
Q_ASSIGN U7740 ( .B(clk), .A(\g.we_clk [25034]));
Q_ASSIGN U7741 ( .B(clk), .A(\g.we_clk [25033]));
Q_ASSIGN U7742 ( .B(clk), .A(\g.we_clk [25032]));
Q_ASSIGN U7743 ( .B(clk), .A(\g.we_clk [25031]));
Q_ASSIGN U7744 ( .B(clk), .A(\g.we_clk [25030]));
Q_ASSIGN U7745 ( .B(clk), .A(\g.we_clk [25029]));
Q_ASSIGN U7746 ( .B(clk), .A(\g.we_clk [25028]));
Q_ASSIGN U7747 ( .B(clk), .A(\g.we_clk [25027]));
Q_ASSIGN U7748 ( .B(clk), .A(\g.we_clk [25026]));
Q_ASSIGN U7749 ( .B(clk), .A(\g.we_clk [25025]));
Q_ASSIGN U7750 ( .B(clk), .A(\g.we_clk [25024]));
Q_ASSIGN U7751 ( .B(clk), .A(\g.we_clk [25023]));
Q_ASSIGN U7752 ( .B(clk), .A(\g.we_clk [25022]));
Q_ASSIGN U7753 ( .B(clk), .A(\g.we_clk [25021]));
Q_ASSIGN U7754 ( .B(clk), .A(\g.we_clk [25020]));
Q_ASSIGN U7755 ( .B(clk), .A(\g.we_clk [25019]));
Q_ASSIGN U7756 ( .B(clk), .A(\g.we_clk [25018]));
Q_ASSIGN U7757 ( .B(clk), .A(\g.we_clk [25017]));
Q_ASSIGN U7758 ( .B(clk), .A(\g.we_clk [25016]));
Q_ASSIGN U7759 ( .B(clk), .A(\g.we_clk [25015]));
Q_ASSIGN U7760 ( .B(clk), .A(\g.we_clk [25014]));
Q_ASSIGN U7761 ( .B(clk), .A(\g.we_clk [25013]));
Q_ASSIGN U7762 ( .B(clk), .A(\g.we_clk [25012]));
Q_ASSIGN U7763 ( .B(clk), .A(\g.we_clk [25011]));
Q_ASSIGN U7764 ( .B(clk), .A(\g.we_clk [25010]));
Q_ASSIGN U7765 ( .B(clk), .A(\g.we_clk [25009]));
Q_ASSIGN U7766 ( .B(clk), .A(\g.we_clk [25008]));
Q_ASSIGN U7767 ( .B(clk), .A(\g.we_clk [25007]));
Q_ASSIGN U7768 ( .B(clk), .A(\g.we_clk [25006]));
Q_ASSIGN U7769 ( .B(clk), .A(\g.we_clk [25005]));
Q_ASSIGN U7770 ( .B(clk), .A(\g.we_clk [25004]));
Q_ASSIGN U7771 ( .B(clk), .A(\g.we_clk [25003]));
Q_ASSIGN U7772 ( .B(clk), .A(\g.we_clk [25002]));
Q_ASSIGN U7773 ( .B(clk), .A(\g.we_clk [25001]));
Q_ASSIGN U7774 ( .B(clk), .A(\g.we_clk [25000]));
Q_ASSIGN U7775 ( .B(clk), .A(\g.we_clk [24999]));
Q_ASSIGN U7776 ( .B(clk), .A(\g.we_clk [24998]));
Q_ASSIGN U7777 ( .B(clk), .A(\g.we_clk [24997]));
Q_ASSIGN U7778 ( .B(clk), .A(\g.we_clk [24996]));
Q_ASSIGN U7779 ( .B(clk), .A(\g.we_clk [24995]));
Q_ASSIGN U7780 ( .B(clk), .A(\g.we_clk [24994]));
Q_ASSIGN U7781 ( .B(clk), .A(\g.we_clk [24993]));
Q_ASSIGN U7782 ( .B(clk), .A(\g.we_clk [24992]));
Q_ASSIGN U7783 ( .B(clk), .A(\g.we_clk [24991]));
Q_ASSIGN U7784 ( .B(clk), .A(\g.we_clk [24990]));
Q_ASSIGN U7785 ( .B(clk), .A(\g.we_clk [24989]));
Q_ASSIGN U7786 ( .B(clk), .A(\g.we_clk [24988]));
Q_ASSIGN U7787 ( .B(clk), .A(\g.we_clk [24987]));
Q_ASSIGN U7788 ( .B(clk), .A(\g.we_clk [24986]));
Q_ASSIGN U7789 ( .B(clk), .A(\g.we_clk [24985]));
Q_ASSIGN U7790 ( .B(clk), .A(\g.we_clk [24984]));
Q_ASSIGN U7791 ( .B(clk), .A(\g.we_clk [24983]));
Q_ASSIGN U7792 ( .B(clk), .A(\g.we_clk [24982]));
Q_ASSIGN U7793 ( .B(clk), .A(\g.we_clk [24981]));
Q_ASSIGN U7794 ( .B(clk), .A(\g.we_clk [24980]));
Q_ASSIGN U7795 ( .B(clk), .A(\g.we_clk [24979]));
Q_ASSIGN U7796 ( .B(clk), .A(\g.we_clk [24978]));
Q_ASSIGN U7797 ( .B(clk), .A(\g.we_clk [24977]));
Q_ASSIGN U7798 ( .B(clk), .A(\g.we_clk [24976]));
Q_ASSIGN U7799 ( .B(clk), .A(\g.we_clk [24975]));
Q_ASSIGN U7800 ( .B(clk), .A(\g.we_clk [24974]));
Q_ASSIGN U7801 ( .B(clk), .A(\g.we_clk [24973]));
Q_ASSIGN U7802 ( .B(clk), .A(\g.we_clk [24972]));
Q_ASSIGN U7803 ( .B(clk), .A(\g.we_clk [24971]));
Q_ASSIGN U7804 ( .B(clk), .A(\g.we_clk [24970]));
Q_ASSIGN U7805 ( .B(clk), .A(\g.we_clk [24969]));
Q_ASSIGN U7806 ( .B(clk), .A(\g.we_clk [24968]));
Q_ASSIGN U7807 ( .B(clk), .A(\g.we_clk [24967]));
Q_ASSIGN U7808 ( .B(clk), .A(\g.we_clk [24966]));
Q_ASSIGN U7809 ( .B(clk), .A(\g.we_clk [24965]));
Q_ASSIGN U7810 ( .B(clk), .A(\g.we_clk [24964]));
Q_ASSIGN U7811 ( .B(clk), .A(\g.we_clk [24963]));
Q_ASSIGN U7812 ( .B(clk), .A(\g.we_clk [24962]));
Q_ASSIGN U7813 ( .B(clk), .A(\g.we_clk [24961]));
Q_ASSIGN U7814 ( .B(clk), .A(\g.we_clk [24960]));
Q_ASSIGN U7815 ( .B(clk), .A(\g.we_clk [24959]));
Q_ASSIGN U7816 ( .B(clk), .A(\g.we_clk [24958]));
Q_ASSIGN U7817 ( .B(clk), .A(\g.we_clk [24957]));
Q_ASSIGN U7818 ( .B(clk), .A(\g.we_clk [24956]));
Q_ASSIGN U7819 ( .B(clk), .A(\g.we_clk [24955]));
Q_ASSIGN U7820 ( .B(clk), .A(\g.we_clk [24954]));
Q_ASSIGN U7821 ( .B(clk), .A(\g.we_clk [24953]));
Q_ASSIGN U7822 ( .B(clk), .A(\g.we_clk [24952]));
Q_ASSIGN U7823 ( .B(clk), .A(\g.we_clk [24951]));
Q_ASSIGN U7824 ( .B(clk), .A(\g.we_clk [24950]));
Q_ASSIGN U7825 ( .B(clk), .A(\g.we_clk [24949]));
Q_ASSIGN U7826 ( .B(clk), .A(\g.we_clk [24948]));
Q_ASSIGN U7827 ( .B(clk), .A(\g.we_clk [24947]));
Q_ASSIGN U7828 ( .B(clk), .A(\g.we_clk [24946]));
Q_ASSIGN U7829 ( .B(clk), .A(\g.we_clk [24945]));
Q_ASSIGN U7830 ( .B(clk), .A(\g.we_clk [24944]));
Q_ASSIGN U7831 ( .B(clk), .A(\g.we_clk [24943]));
Q_ASSIGN U7832 ( .B(clk), .A(\g.we_clk [24942]));
Q_ASSIGN U7833 ( .B(clk), .A(\g.we_clk [24941]));
Q_ASSIGN U7834 ( .B(clk), .A(\g.we_clk [24940]));
Q_ASSIGN U7835 ( .B(clk), .A(\g.we_clk [24939]));
Q_ASSIGN U7836 ( .B(clk), .A(\g.we_clk [24938]));
Q_ASSIGN U7837 ( .B(clk), .A(\g.we_clk [24937]));
Q_ASSIGN U7838 ( .B(clk), .A(\g.we_clk [24936]));
Q_ASSIGN U7839 ( .B(clk), .A(\g.we_clk [24935]));
Q_ASSIGN U7840 ( .B(clk), .A(\g.we_clk [24934]));
Q_ASSIGN U7841 ( .B(clk), .A(\g.we_clk [24933]));
Q_ASSIGN U7842 ( .B(clk), .A(\g.we_clk [24932]));
Q_ASSIGN U7843 ( .B(clk), .A(\g.we_clk [24931]));
Q_ASSIGN U7844 ( .B(clk), .A(\g.we_clk [24930]));
Q_ASSIGN U7845 ( .B(clk), .A(\g.we_clk [24929]));
Q_ASSIGN U7846 ( .B(clk), .A(\g.we_clk [24928]));
Q_ASSIGN U7847 ( .B(clk), .A(\g.we_clk [24927]));
Q_ASSIGN U7848 ( .B(clk), .A(\g.we_clk [24926]));
Q_ASSIGN U7849 ( .B(clk), .A(\g.we_clk [24925]));
Q_ASSIGN U7850 ( .B(clk), .A(\g.we_clk [24924]));
Q_ASSIGN U7851 ( .B(clk), .A(\g.we_clk [24923]));
Q_ASSIGN U7852 ( .B(clk), .A(\g.we_clk [24922]));
Q_ASSIGN U7853 ( .B(clk), .A(\g.we_clk [24921]));
Q_ASSIGN U7854 ( .B(clk), .A(\g.we_clk [24920]));
Q_ASSIGN U7855 ( .B(clk), .A(\g.we_clk [24919]));
Q_ASSIGN U7856 ( .B(clk), .A(\g.we_clk [24918]));
Q_ASSIGN U7857 ( .B(clk), .A(\g.we_clk [24917]));
Q_ASSIGN U7858 ( .B(clk), .A(\g.we_clk [24916]));
Q_ASSIGN U7859 ( .B(clk), .A(\g.we_clk [24915]));
Q_ASSIGN U7860 ( .B(clk), .A(\g.we_clk [24914]));
Q_ASSIGN U7861 ( .B(clk), .A(\g.we_clk [24913]));
Q_ASSIGN U7862 ( .B(clk), .A(\g.we_clk [24912]));
Q_ASSIGN U7863 ( .B(clk), .A(\g.we_clk [24911]));
Q_ASSIGN U7864 ( .B(clk), .A(\g.we_clk [24910]));
Q_ASSIGN U7865 ( .B(clk), .A(\g.we_clk [24909]));
Q_ASSIGN U7866 ( .B(clk), .A(\g.we_clk [24908]));
Q_ASSIGN U7867 ( .B(clk), .A(\g.we_clk [24907]));
Q_ASSIGN U7868 ( .B(clk), .A(\g.we_clk [24906]));
Q_ASSIGN U7869 ( .B(clk), .A(\g.we_clk [24905]));
Q_ASSIGN U7870 ( .B(clk), .A(\g.we_clk [24904]));
Q_ASSIGN U7871 ( .B(clk), .A(\g.we_clk [24903]));
Q_ASSIGN U7872 ( .B(clk), .A(\g.we_clk [24902]));
Q_ASSIGN U7873 ( .B(clk), .A(\g.we_clk [24901]));
Q_ASSIGN U7874 ( .B(clk), .A(\g.we_clk [24900]));
Q_ASSIGN U7875 ( .B(clk), .A(\g.we_clk [24899]));
Q_ASSIGN U7876 ( .B(clk), .A(\g.we_clk [24898]));
Q_ASSIGN U7877 ( .B(clk), .A(\g.we_clk [24897]));
Q_ASSIGN U7878 ( .B(clk), .A(\g.we_clk [24896]));
Q_ASSIGN U7879 ( .B(clk), .A(\g.we_clk [24895]));
Q_ASSIGN U7880 ( .B(clk), .A(\g.we_clk [24894]));
Q_ASSIGN U7881 ( .B(clk), .A(\g.we_clk [24893]));
Q_ASSIGN U7882 ( .B(clk), .A(\g.we_clk [24892]));
Q_ASSIGN U7883 ( .B(clk), .A(\g.we_clk [24891]));
Q_ASSIGN U7884 ( .B(clk), .A(\g.we_clk [24890]));
Q_ASSIGN U7885 ( .B(clk), .A(\g.we_clk [24889]));
Q_ASSIGN U7886 ( .B(clk), .A(\g.we_clk [24888]));
Q_ASSIGN U7887 ( .B(clk), .A(\g.we_clk [24887]));
Q_ASSIGN U7888 ( .B(clk), .A(\g.we_clk [24886]));
Q_ASSIGN U7889 ( .B(clk), .A(\g.we_clk [24885]));
Q_ASSIGN U7890 ( .B(clk), .A(\g.we_clk [24884]));
Q_ASSIGN U7891 ( .B(clk), .A(\g.we_clk [24883]));
Q_ASSIGN U7892 ( .B(clk), .A(\g.we_clk [24882]));
Q_ASSIGN U7893 ( .B(clk), .A(\g.we_clk [24881]));
Q_ASSIGN U7894 ( .B(clk), .A(\g.we_clk [24880]));
Q_ASSIGN U7895 ( .B(clk), .A(\g.we_clk [24879]));
Q_ASSIGN U7896 ( .B(clk), .A(\g.we_clk [24878]));
Q_ASSIGN U7897 ( .B(clk), .A(\g.we_clk [24877]));
Q_ASSIGN U7898 ( .B(clk), .A(\g.we_clk [24876]));
Q_ASSIGN U7899 ( .B(clk), .A(\g.we_clk [24875]));
Q_ASSIGN U7900 ( .B(clk), .A(\g.we_clk [24874]));
Q_ASSIGN U7901 ( .B(clk), .A(\g.we_clk [24873]));
Q_ASSIGN U7902 ( .B(clk), .A(\g.we_clk [24872]));
Q_ASSIGN U7903 ( .B(clk), .A(\g.we_clk [24871]));
Q_ASSIGN U7904 ( .B(clk), .A(\g.we_clk [24870]));
Q_ASSIGN U7905 ( .B(clk), .A(\g.we_clk [24869]));
Q_ASSIGN U7906 ( .B(clk), .A(\g.we_clk [24868]));
Q_ASSIGN U7907 ( .B(clk), .A(\g.we_clk [24867]));
Q_ASSIGN U7908 ( .B(clk), .A(\g.we_clk [24866]));
Q_ASSIGN U7909 ( .B(clk), .A(\g.we_clk [24865]));
Q_ASSIGN U7910 ( .B(clk), .A(\g.we_clk [24864]));
Q_ASSIGN U7911 ( .B(clk), .A(\g.we_clk [24863]));
Q_ASSIGN U7912 ( .B(clk), .A(\g.we_clk [24862]));
Q_ASSIGN U7913 ( .B(clk), .A(\g.we_clk [24861]));
Q_ASSIGN U7914 ( .B(clk), .A(\g.we_clk [24860]));
Q_ASSIGN U7915 ( .B(clk), .A(\g.we_clk [24859]));
Q_ASSIGN U7916 ( .B(clk), .A(\g.we_clk [24858]));
Q_ASSIGN U7917 ( .B(clk), .A(\g.we_clk [24857]));
Q_ASSIGN U7918 ( .B(clk), .A(\g.we_clk [24856]));
Q_ASSIGN U7919 ( .B(clk), .A(\g.we_clk [24855]));
Q_ASSIGN U7920 ( .B(clk), .A(\g.we_clk [24854]));
Q_ASSIGN U7921 ( .B(clk), .A(\g.we_clk [24853]));
Q_ASSIGN U7922 ( .B(clk), .A(\g.we_clk [24852]));
Q_ASSIGN U7923 ( .B(clk), .A(\g.we_clk [24851]));
Q_ASSIGN U7924 ( .B(clk), .A(\g.we_clk [24850]));
Q_ASSIGN U7925 ( .B(clk), .A(\g.we_clk [24849]));
Q_ASSIGN U7926 ( .B(clk), .A(\g.we_clk [24848]));
Q_ASSIGN U7927 ( .B(clk), .A(\g.we_clk [24847]));
Q_ASSIGN U7928 ( .B(clk), .A(\g.we_clk [24846]));
Q_ASSIGN U7929 ( .B(clk), .A(\g.we_clk [24845]));
Q_ASSIGN U7930 ( .B(clk), .A(\g.we_clk [24844]));
Q_ASSIGN U7931 ( .B(clk), .A(\g.we_clk [24843]));
Q_ASSIGN U7932 ( .B(clk), .A(\g.we_clk [24842]));
Q_ASSIGN U7933 ( .B(clk), .A(\g.we_clk [24841]));
Q_ASSIGN U7934 ( .B(clk), .A(\g.we_clk [24840]));
Q_ASSIGN U7935 ( .B(clk), .A(\g.we_clk [24839]));
Q_ASSIGN U7936 ( .B(clk), .A(\g.we_clk [24838]));
Q_ASSIGN U7937 ( .B(clk), .A(\g.we_clk [24837]));
Q_ASSIGN U7938 ( .B(clk), .A(\g.we_clk [24836]));
Q_ASSIGN U7939 ( .B(clk), .A(\g.we_clk [24835]));
Q_ASSIGN U7940 ( .B(clk), .A(\g.we_clk [24834]));
Q_ASSIGN U7941 ( .B(clk), .A(\g.we_clk [24833]));
Q_ASSIGN U7942 ( .B(clk), .A(\g.we_clk [24832]));
Q_ASSIGN U7943 ( .B(clk), .A(\g.we_clk [24831]));
Q_ASSIGN U7944 ( .B(clk), .A(\g.we_clk [24830]));
Q_ASSIGN U7945 ( .B(clk), .A(\g.we_clk [24829]));
Q_ASSIGN U7946 ( .B(clk), .A(\g.we_clk [24828]));
Q_ASSIGN U7947 ( .B(clk), .A(\g.we_clk [24827]));
Q_ASSIGN U7948 ( .B(clk), .A(\g.we_clk [24826]));
Q_ASSIGN U7949 ( .B(clk), .A(\g.we_clk [24825]));
Q_ASSIGN U7950 ( .B(clk), .A(\g.we_clk [24824]));
Q_ASSIGN U7951 ( .B(clk), .A(\g.we_clk [24823]));
Q_ASSIGN U7952 ( .B(clk), .A(\g.we_clk [24822]));
Q_ASSIGN U7953 ( .B(clk), .A(\g.we_clk [24821]));
Q_ASSIGN U7954 ( .B(clk), .A(\g.we_clk [24820]));
Q_ASSIGN U7955 ( .B(clk), .A(\g.we_clk [24819]));
Q_ASSIGN U7956 ( .B(clk), .A(\g.we_clk [24818]));
Q_ASSIGN U7957 ( .B(clk), .A(\g.we_clk [24817]));
Q_ASSIGN U7958 ( .B(clk), .A(\g.we_clk [24816]));
Q_ASSIGN U7959 ( .B(clk), .A(\g.we_clk [24815]));
Q_ASSIGN U7960 ( .B(clk), .A(\g.we_clk [24814]));
Q_ASSIGN U7961 ( .B(clk), .A(\g.we_clk [24813]));
Q_ASSIGN U7962 ( .B(clk), .A(\g.we_clk [24812]));
Q_ASSIGN U7963 ( .B(clk), .A(\g.we_clk [24811]));
Q_ASSIGN U7964 ( .B(clk), .A(\g.we_clk [24810]));
Q_ASSIGN U7965 ( .B(clk), .A(\g.we_clk [24809]));
Q_ASSIGN U7966 ( .B(clk), .A(\g.we_clk [24808]));
Q_ASSIGN U7967 ( .B(clk), .A(\g.we_clk [24807]));
Q_ASSIGN U7968 ( .B(clk), .A(\g.we_clk [24806]));
Q_ASSIGN U7969 ( .B(clk), .A(\g.we_clk [24805]));
Q_ASSIGN U7970 ( .B(clk), .A(\g.we_clk [24804]));
Q_ASSIGN U7971 ( .B(clk), .A(\g.we_clk [24803]));
Q_ASSIGN U7972 ( .B(clk), .A(\g.we_clk [24802]));
Q_ASSIGN U7973 ( .B(clk), .A(\g.we_clk [24801]));
Q_ASSIGN U7974 ( .B(clk), .A(\g.we_clk [24800]));
Q_ASSIGN U7975 ( .B(clk), .A(\g.we_clk [24799]));
Q_ASSIGN U7976 ( .B(clk), .A(\g.we_clk [24798]));
Q_ASSIGN U7977 ( .B(clk), .A(\g.we_clk [24797]));
Q_ASSIGN U7978 ( .B(clk), .A(\g.we_clk [24796]));
Q_ASSIGN U7979 ( .B(clk), .A(\g.we_clk [24795]));
Q_ASSIGN U7980 ( .B(clk), .A(\g.we_clk [24794]));
Q_ASSIGN U7981 ( .B(clk), .A(\g.we_clk [24793]));
Q_ASSIGN U7982 ( .B(clk), .A(\g.we_clk [24792]));
Q_ASSIGN U7983 ( .B(clk), .A(\g.we_clk [24791]));
Q_ASSIGN U7984 ( .B(clk), .A(\g.we_clk [24790]));
Q_ASSIGN U7985 ( .B(clk), .A(\g.we_clk [24789]));
Q_ASSIGN U7986 ( .B(clk), .A(\g.we_clk [24788]));
Q_ASSIGN U7987 ( .B(clk), .A(\g.we_clk [24787]));
Q_ASSIGN U7988 ( .B(clk), .A(\g.we_clk [24786]));
Q_ASSIGN U7989 ( .B(clk), .A(\g.we_clk [24785]));
Q_ASSIGN U7990 ( .B(clk), .A(\g.we_clk [24784]));
Q_ASSIGN U7991 ( .B(clk), .A(\g.we_clk [24783]));
Q_ASSIGN U7992 ( .B(clk), .A(\g.we_clk [24782]));
Q_ASSIGN U7993 ( .B(clk), .A(\g.we_clk [24781]));
Q_ASSIGN U7994 ( .B(clk), .A(\g.we_clk [24780]));
Q_ASSIGN U7995 ( .B(clk), .A(\g.we_clk [24779]));
Q_ASSIGN U7996 ( .B(clk), .A(\g.we_clk [24778]));
Q_ASSIGN U7997 ( .B(clk), .A(\g.we_clk [24777]));
Q_ASSIGN U7998 ( .B(clk), .A(\g.we_clk [24776]));
Q_ASSIGN U7999 ( .B(clk), .A(\g.we_clk [24775]));
Q_ASSIGN U8000 ( .B(clk), .A(\g.we_clk [24774]));
Q_ASSIGN U8001 ( .B(clk), .A(\g.we_clk [24773]));
Q_ASSIGN U8002 ( .B(clk), .A(\g.we_clk [24772]));
Q_ASSIGN U8003 ( .B(clk), .A(\g.we_clk [24771]));
Q_ASSIGN U8004 ( .B(clk), .A(\g.we_clk [24770]));
Q_ASSIGN U8005 ( .B(clk), .A(\g.we_clk [24769]));
Q_ASSIGN U8006 ( .B(clk), .A(\g.we_clk [24768]));
Q_ASSIGN U8007 ( .B(clk), .A(\g.we_clk [24767]));
Q_ASSIGN U8008 ( .B(clk), .A(\g.we_clk [24766]));
Q_ASSIGN U8009 ( .B(clk), .A(\g.we_clk [24765]));
Q_ASSIGN U8010 ( .B(clk), .A(\g.we_clk [24764]));
Q_ASSIGN U8011 ( .B(clk), .A(\g.we_clk [24763]));
Q_ASSIGN U8012 ( .B(clk), .A(\g.we_clk [24762]));
Q_ASSIGN U8013 ( .B(clk), .A(\g.we_clk [24761]));
Q_ASSIGN U8014 ( .B(clk), .A(\g.we_clk [24760]));
Q_ASSIGN U8015 ( .B(clk), .A(\g.we_clk [24759]));
Q_ASSIGN U8016 ( .B(clk), .A(\g.we_clk [24758]));
Q_ASSIGN U8017 ( .B(clk), .A(\g.we_clk [24757]));
Q_ASSIGN U8018 ( .B(clk), .A(\g.we_clk [24756]));
Q_ASSIGN U8019 ( .B(clk), .A(\g.we_clk [24755]));
Q_ASSIGN U8020 ( .B(clk), .A(\g.we_clk [24754]));
Q_ASSIGN U8021 ( .B(clk), .A(\g.we_clk [24753]));
Q_ASSIGN U8022 ( .B(clk), .A(\g.we_clk [24752]));
Q_ASSIGN U8023 ( .B(clk), .A(\g.we_clk [24751]));
Q_ASSIGN U8024 ( .B(clk), .A(\g.we_clk [24750]));
Q_ASSIGN U8025 ( .B(clk), .A(\g.we_clk [24749]));
Q_ASSIGN U8026 ( .B(clk), .A(\g.we_clk [24748]));
Q_ASSIGN U8027 ( .B(clk), .A(\g.we_clk [24747]));
Q_ASSIGN U8028 ( .B(clk), .A(\g.we_clk [24746]));
Q_ASSIGN U8029 ( .B(clk), .A(\g.we_clk [24745]));
Q_ASSIGN U8030 ( .B(clk), .A(\g.we_clk [24744]));
Q_ASSIGN U8031 ( .B(clk), .A(\g.we_clk [24743]));
Q_ASSIGN U8032 ( .B(clk), .A(\g.we_clk [24742]));
Q_ASSIGN U8033 ( .B(clk), .A(\g.we_clk [24741]));
Q_ASSIGN U8034 ( .B(clk), .A(\g.we_clk [24740]));
Q_ASSIGN U8035 ( .B(clk), .A(\g.we_clk [24739]));
Q_ASSIGN U8036 ( .B(clk), .A(\g.we_clk [24738]));
Q_ASSIGN U8037 ( .B(clk), .A(\g.we_clk [24737]));
Q_ASSIGN U8038 ( .B(clk), .A(\g.we_clk [24736]));
Q_ASSIGN U8039 ( .B(clk), .A(\g.we_clk [24735]));
Q_ASSIGN U8040 ( .B(clk), .A(\g.we_clk [24734]));
Q_ASSIGN U8041 ( .B(clk), .A(\g.we_clk [24733]));
Q_ASSIGN U8042 ( .B(clk), .A(\g.we_clk [24732]));
Q_ASSIGN U8043 ( .B(clk), .A(\g.we_clk [24731]));
Q_ASSIGN U8044 ( .B(clk), .A(\g.we_clk [24730]));
Q_ASSIGN U8045 ( .B(clk), .A(\g.we_clk [24729]));
Q_ASSIGN U8046 ( .B(clk), .A(\g.we_clk [24728]));
Q_ASSIGN U8047 ( .B(clk), .A(\g.we_clk [24727]));
Q_ASSIGN U8048 ( .B(clk), .A(\g.we_clk [24726]));
Q_ASSIGN U8049 ( .B(clk), .A(\g.we_clk [24725]));
Q_ASSIGN U8050 ( .B(clk), .A(\g.we_clk [24724]));
Q_ASSIGN U8051 ( .B(clk), .A(\g.we_clk [24723]));
Q_ASSIGN U8052 ( .B(clk), .A(\g.we_clk [24722]));
Q_ASSIGN U8053 ( .B(clk), .A(\g.we_clk [24721]));
Q_ASSIGN U8054 ( .B(clk), .A(\g.we_clk [24720]));
Q_ASSIGN U8055 ( .B(clk), .A(\g.we_clk [24719]));
Q_ASSIGN U8056 ( .B(clk), .A(\g.we_clk [24718]));
Q_ASSIGN U8057 ( .B(clk), .A(\g.we_clk [24717]));
Q_ASSIGN U8058 ( .B(clk), .A(\g.we_clk [24716]));
Q_ASSIGN U8059 ( .B(clk), .A(\g.we_clk [24715]));
Q_ASSIGN U8060 ( .B(clk), .A(\g.we_clk [24714]));
Q_ASSIGN U8061 ( .B(clk), .A(\g.we_clk [24713]));
Q_ASSIGN U8062 ( .B(clk), .A(\g.we_clk [24712]));
Q_ASSIGN U8063 ( .B(clk), .A(\g.we_clk [24711]));
Q_ASSIGN U8064 ( .B(clk), .A(\g.we_clk [24710]));
Q_ASSIGN U8065 ( .B(clk), .A(\g.we_clk [24709]));
Q_ASSIGN U8066 ( .B(clk), .A(\g.we_clk [24708]));
Q_ASSIGN U8067 ( .B(clk), .A(\g.we_clk [24707]));
Q_ASSIGN U8068 ( .B(clk), .A(\g.we_clk [24706]));
Q_ASSIGN U8069 ( .B(clk), .A(\g.we_clk [24705]));
Q_ASSIGN U8070 ( .B(clk), .A(\g.we_clk [24704]));
Q_ASSIGN U8071 ( .B(clk), .A(\g.we_clk [24703]));
Q_ASSIGN U8072 ( .B(clk), .A(\g.we_clk [24702]));
Q_ASSIGN U8073 ( .B(clk), .A(\g.we_clk [24701]));
Q_ASSIGN U8074 ( .B(clk), .A(\g.we_clk [24700]));
Q_ASSIGN U8075 ( .B(clk), .A(\g.we_clk [24699]));
Q_ASSIGN U8076 ( .B(clk), .A(\g.we_clk [24698]));
Q_ASSIGN U8077 ( .B(clk), .A(\g.we_clk [24697]));
Q_ASSIGN U8078 ( .B(clk), .A(\g.we_clk [24696]));
Q_ASSIGN U8079 ( .B(clk), .A(\g.we_clk [24695]));
Q_ASSIGN U8080 ( .B(clk), .A(\g.we_clk [24694]));
Q_ASSIGN U8081 ( .B(clk), .A(\g.we_clk [24693]));
Q_ASSIGN U8082 ( .B(clk), .A(\g.we_clk [24692]));
Q_ASSIGN U8083 ( .B(clk), .A(\g.we_clk [24691]));
Q_ASSIGN U8084 ( .B(clk), .A(\g.we_clk [24690]));
Q_ASSIGN U8085 ( .B(clk), .A(\g.we_clk [24689]));
Q_ASSIGN U8086 ( .B(clk), .A(\g.we_clk [24688]));
Q_ASSIGN U8087 ( .B(clk), .A(\g.we_clk [24687]));
Q_ASSIGN U8088 ( .B(clk), .A(\g.we_clk [24686]));
Q_ASSIGN U8089 ( .B(clk), .A(\g.we_clk [24685]));
Q_ASSIGN U8090 ( .B(clk), .A(\g.we_clk [24684]));
Q_ASSIGN U8091 ( .B(clk), .A(\g.we_clk [24683]));
Q_ASSIGN U8092 ( .B(clk), .A(\g.we_clk [24682]));
Q_ASSIGN U8093 ( .B(clk), .A(\g.we_clk [24681]));
Q_ASSIGN U8094 ( .B(clk), .A(\g.we_clk [24680]));
Q_ASSIGN U8095 ( .B(clk), .A(\g.we_clk [24679]));
Q_ASSIGN U8096 ( .B(clk), .A(\g.we_clk [24678]));
Q_ASSIGN U8097 ( .B(clk), .A(\g.we_clk [24677]));
Q_ASSIGN U8098 ( .B(clk), .A(\g.we_clk [24676]));
Q_ASSIGN U8099 ( .B(clk), .A(\g.we_clk [24675]));
Q_ASSIGN U8100 ( .B(clk), .A(\g.we_clk [24674]));
Q_ASSIGN U8101 ( .B(clk), .A(\g.we_clk [24673]));
Q_ASSIGN U8102 ( .B(clk), .A(\g.we_clk [24672]));
Q_ASSIGN U8103 ( .B(clk), .A(\g.we_clk [24671]));
Q_ASSIGN U8104 ( .B(clk), .A(\g.we_clk [24670]));
Q_ASSIGN U8105 ( .B(clk), .A(\g.we_clk [24669]));
Q_ASSIGN U8106 ( .B(clk), .A(\g.we_clk [24668]));
Q_ASSIGN U8107 ( .B(clk), .A(\g.we_clk [24667]));
Q_ASSIGN U8108 ( .B(clk), .A(\g.we_clk [24666]));
Q_ASSIGN U8109 ( .B(clk), .A(\g.we_clk [24665]));
Q_ASSIGN U8110 ( .B(clk), .A(\g.we_clk [24664]));
Q_ASSIGN U8111 ( .B(clk), .A(\g.we_clk [24663]));
Q_ASSIGN U8112 ( .B(clk), .A(\g.we_clk [24662]));
Q_ASSIGN U8113 ( .B(clk), .A(\g.we_clk [24661]));
Q_ASSIGN U8114 ( .B(clk), .A(\g.we_clk [24660]));
Q_ASSIGN U8115 ( .B(clk), .A(\g.we_clk [24659]));
Q_ASSIGN U8116 ( .B(clk), .A(\g.we_clk [24658]));
Q_ASSIGN U8117 ( .B(clk), .A(\g.we_clk [24657]));
Q_ASSIGN U8118 ( .B(clk), .A(\g.we_clk [24656]));
Q_ASSIGN U8119 ( .B(clk), .A(\g.we_clk [24655]));
Q_ASSIGN U8120 ( .B(clk), .A(\g.we_clk [24654]));
Q_ASSIGN U8121 ( .B(clk), .A(\g.we_clk [24653]));
Q_ASSIGN U8122 ( .B(clk), .A(\g.we_clk [24652]));
Q_ASSIGN U8123 ( .B(clk), .A(\g.we_clk [24651]));
Q_ASSIGN U8124 ( .B(clk), .A(\g.we_clk [24650]));
Q_ASSIGN U8125 ( .B(clk), .A(\g.we_clk [24649]));
Q_ASSIGN U8126 ( .B(clk), .A(\g.we_clk [24648]));
Q_ASSIGN U8127 ( .B(clk), .A(\g.we_clk [24647]));
Q_ASSIGN U8128 ( .B(clk), .A(\g.we_clk [24646]));
Q_ASSIGN U8129 ( .B(clk), .A(\g.we_clk [24645]));
Q_ASSIGN U8130 ( .B(clk), .A(\g.we_clk [24644]));
Q_ASSIGN U8131 ( .B(clk), .A(\g.we_clk [24643]));
Q_ASSIGN U8132 ( .B(clk), .A(\g.we_clk [24642]));
Q_ASSIGN U8133 ( .B(clk), .A(\g.we_clk [24641]));
Q_ASSIGN U8134 ( .B(clk), .A(\g.we_clk [24640]));
Q_ASSIGN U8135 ( .B(clk), .A(\g.we_clk [24639]));
Q_ASSIGN U8136 ( .B(clk), .A(\g.we_clk [24638]));
Q_ASSIGN U8137 ( .B(clk), .A(\g.we_clk [24637]));
Q_ASSIGN U8138 ( .B(clk), .A(\g.we_clk [24636]));
Q_ASSIGN U8139 ( .B(clk), .A(\g.we_clk [24635]));
Q_ASSIGN U8140 ( .B(clk), .A(\g.we_clk [24634]));
Q_ASSIGN U8141 ( .B(clk), .A(\g.we_clk [24633]));
Q_ASSIGN U8142 ( .B(clk), .A(\g.we_clk [24632]));
Q_ASSIGN U8143 ( .B(clk), .A(\g.we_clk [24631]));
Q_ASSIGN U8144 ( .B(clk), .A(\g.we_clk [24630]));
Q_ASSIGN U8145 ( .B(clk), .A(\g.we_clk [24629]));
Q_ASSIGN U8146 ( .B(clk), .A(\g.we_clk [24628]));
Q_ASSIGN U8147 ( .B(clk), .A(\g.we_clk [24627]));
Q_ASSIGN U8148 ( .B(clk), .A(\g.we_clk [24626]));
Q_ASSIGN U8149 ( .B(clk), .A(\g.we_clk [24625]));
Q_ASSIGN U8150 ( .B(clk), .A(\g.we_clk [24624]));
Q_ASSIGN U8151 ( .B(clk), .A(\g.we_clk [24623]));
Q_ASSIGN U8152 ( .B(clk), .A(\g.we_clk [24622]));
Q_ASSIGN U8153 ( .B(clk), .A(\g.we_clk [24621]));
Q_ASSIGN U8154 ( .B(clk), .A(\g.we_clk [24620]));
Q_ASSIGN U8155 ( .B(clk), .A(\g.we_clk [24619]));
Q_ASSIGN U8156 ( .B(clk), .A(\g.we_clk [24618]));
Q_ASSIGN U8157 ( .B(clk), .A(\g.we_clk [24617]));
Q_ASSIGN U8158 ( .B(clk), .A(\g.we_clk [24616]));
Q_ASSIGN U8159 ( .B(clk), .A(\g.we_clk [24615]));
Q_ASSIGN U8160 ( .B(clk), .A(\g.we_clk [24614]));
Q_ASSIGN U8161 ( .B(clk), .A(\g.we_clk [24613]));
Q_ASSIGN U8162 ( .B(clk), .A(\g.we_clk [24612]));
Q_ASSIGN U8163 ( .B(clk), .A(\g.we_clk [24611]));
Q_ASSIGN U8164 ( .B(clk), .A(\g.we_clk [24610]));
Q_ASSIGN U8165 ( .B(clk), .A(\g.we_clk [24609]));
Q_ASSIGN U8166 ( .B(clk), .A(\g.we_clk [24608]));
Q_ASSIGN U8167 ( .B(clk), .A(\g.we_clk [24607]));
Q_ASSIGN U8168 ( .B(clk), .A(\g.we_clk [24606]));
Q_ASSIGN U8169 ( .B(clk), .A(\g.we_clk [24605]));
Q_ASSIGN U8170 ( .B(clk), .A(\g.we_clk [24604]));
Q_ASSIGN U8171 ( .B(clk), .A(\g.we_clk [24603]));
Q_ASSIGN U8172 ( .B(clk), .A(\g.we_clk [24602]));
Q_ASSIGN U8173 ( .B(clk), .A(\g.we_clk [24601]));
Q_ASSIGN U8174 ( .B(clk), .A(\g.we_clk [24600]));
Q_ASSIGN U8175 ( .B(clk), .A(\g.we_clk [24599]));
Q_ASSIGN U8176 ( .B(clk), .A(\g.we_clk [24598]));
Q_ASSIGN U8177 ( .B(clk), .A(\g.we_clk [24597]));
Q_ASSIGN U8178 ( .B(clk), .A(\g.we_clk [24596]));
Q_ASSIGN U8179 ( .B(clk), .A(\g.we_clk [24595]));
Q_ASSIGN U8180 ( .B(clk), .A(\g.we_clk [24594]));
Q_ASSIGN U8181 ( .B(clk), .A(\g.we_clk [24593]));
Q_ASSIGN U8182 ( .B(clk), .A(\g.we_clk [24592]));
Q_ASSIGN U8183 ( .B(clk), .A(\g.we_clk [24591]));
Q_ASSIGN U8184 ( .B(clk), .A(\g.we_clk [24590]));
Q_ASSIGN U8185 ( .B(clk), .A(\g.we_clk [24589]));
Q_ASSIGN U8186 ( .B(clk), .A(\g.we_clk [24588]));
Q_ASSIGN U8187 ( .B(clk), .A(\g.we_clk [24587]));
Q_ASSIGN U8188 ( .B(clk), .A(\g.we_clk [24586]));
Q_ASSIGN U8189 ( .B(clk), .A(\g.we_clk [24585]));
Q_ASSIGN U8190 ( .B(clk), .A(\g.we_clk [24584]));
Q_ASSIGN U8191 ( .B(clk), .A(\g.we_clk [24583]));
Q_ASSIGN U8192 ( .B(clk), .A(\g.we_clk [24582]));
Q_ASSIGN U8193 ( .B(clk), .A(\g.we_clk [24581]));
Q_ASSIGN U8194 ( .B(clk), .A(\g.we_clk [24580]));
Q_ASSIGN U8195 ( .B(clk), .A(\g.we_clk [24579]));
Q_ASSIGN U8196 ( .B(clk), .A(\g.we_clk [24578]));
Q_ASSIGN U8197 ( .B(clk), .A(\g.we_clk [24577]));
Q_ASSIGN U8198 ( .B(clk), .A(\g.we_clk [24576]));
Q_ASSIGN U8199 ( .B(clk), .A(\g.we_clk [24575]));
Q_ASSIGN U8200 ( .B(clk), .A(\g.we_clk [24574]));
Q_ASSIGN U8201 ( .B(clk), .A(\g.we_clk [24573]));
Q_ASSIGN U8202 ( .B(clk), .A(\g.we_clk [24572]));
Q_ASSIGN U8203 ( .B(clk), .A(\g.we_clk [24571]));
Q_ASSIGN U8204 ( .B(clk), .A(\g.we_clk [24570]));
Q_ASSIGN U8205 ( .B(clk), .A(\g.we_clk [24569]));
Q_ASSIGN U8206 ( .B(clk), .A(\g.we_clk [24568]));
Q_ASSIGN U8207 ( .B(clk), .A(\g.we_clk [24567]));
Q_ASSIGN U8208 ( .B(clk), .A(\g.we_clk [24566]));
Q_ASSIGN U8209 ( .B(clk), .A(\g.we_clk [24565]));
Q_ASSIGN U8210 ( .B(clk), .A(\g.we_clk [24564]));
Q_ASSIGN U8211 ( .B(clk), .A(\g.we_clk [24563]));
Q_ASSIGN U8212 ( .B(clk), .A(\g.we_clk [24562]));
Q_ASSIGN U8213 ( .B(clk), .A(\g.we_clk [24561]));
Q_ASSIGN U8214 ( .B(clk), .A(\g.we_clk [24560]));
Q_ASSIGN U8215 ( .B(clk), .A(\g.we_clk [24559]));
Q_ASSIGN U8216 ( .B(clk), .A(\g.we_clk [24558]));
Q_ASSIGN U8217 ( .B(clk), .A(\g.we_clk [24557]));
Q_ASSIGN U8218 ( .B(clk), .A(\g.we_clk [24556]));
Q_ASSIGN U8219 ( .B(clk), .A(\g.we_clk [24555]));
Q_ASSIGN U8220 ( .B(clk), .A(\g.we_clk [24554]));
Q_ASSIGN U8221 ( .B(clk), .A(\g.we_clk [24553]));
Q_ASSIGN U8222 ( .B(clk), .A(\g.we_clk [24552]));
Q_ASSIGN U8223 ( .B(clk), .A(\g.we_clk [24551]));
Q_ASSIGN U8224 ( .B(clk), .A(\g.we_clk [24550]));
Q_ASSIGN U8225 ( .B(clk), .A(\g.we_clk [24549]));
Q_ASSIGN U8226 ( .B(clk), .A(\g.we_clk [24548]));
Q_ASSIGN U8227 ( .B(clk), .A(\g.we_clk [24547]));
Q_ASSIGN U8228 ( .B(clk), .A(\g.we_clk [24546]));
Q_ASSIGN U8229 ( .B(clk), .A(\g.we_clk [24545]));
Q_ASSIGN U8230 ( .B(clk), .A(\g.we_clk [24544]));
Q_ASSIGN U8231 ( .B(clk), .A(\g.we_clk [24543]));
Q_ASSIGN U8232 ( .B(clk), .A(\g.we_clk [24542]));
Q_ASSIGN U8233 ( .B(clk), .A(\g.we_clk [24541]));
Q_ASSIGN U8234 ( .B(clk), .A(\g.we_clk [24540]));
Q_ASSIGN U8235 ( .B(clk), .A(\g.we_clk [24539]));
Q_ASSIGN U8236 ( .B(clk), .A(\g.we_clk [24538]));
Q_ASSIGN U8237 ( .B(clk), .A(\g.we_clk [24537]));
Q_ASSIGN U8238 ( .B(clk), .A(\g.we_clk [24536]));
Q_ASSIGN U8239 ( .B(clk), .A(\g.we_clk [24535]));
Q_ASSIGN U8240 ( .B(clk), .A(\g.we_clk [24534]));
Q_ASSIGN U8241 ( .B(clk), .A(\g.we_clk [24533]));
Q_ASSIGN U8242 ( .B(clk), .A(\g.we_clk [24532]));
Q_ASSIGN U8243 ( .B(clk), .A(\g.we_clk [24531]));
Q_ASSIGN U8244 ( .B(clk), .A(\g.we_clk [24530]));
Q_ASSIGN U8245 ( .B(clk), .A(\g.we_clk [24529]));
Q_ASSIGN U8246 ( .B(clk), .A(\g.we_clk [24528]));
Q_ASSIGN U8247 ( .B(clk), .A(\g.we_clk [24527]));
Q_ASSIGN U8248 ( .B(clk), .A(\g.we_clk [24526]));
Q_ASSIGN U8249 ( .B(clk), .A(\g.we_clk [24525]));
Q_ASSIGN U8250 ( .B(clk), .A(\g.we_clk [24524]));
Q_ASSIGN U8251 ( .B(clk), .A(\g.we_clk [24523]));
Q_ASSIGN U8252 ( .B(clk), .A(\g.we_clk [24522]));
Q_ASSIGN U8253 ( .B(clk), .A(\g.we_clk [24521]));
Q_ASSIGN U8254 ( .B(clk), .A(\g.we_clk [24520]));
Q_ASSIGN U8255 ( .B(clk), .A(\g.we_clk [24519]));
Q_ASSIGN U8256 ( .B(clk), .A(\g.we_clk [24518]));
Q_ASSIGN U8257 ( .B(clk), .A(\g.we_clk [24517]));
Q_ASSIGN U8258 ( .B(clk), .A(\g.we_clk [24516]));
Q_ASSIGN U8259 ( .B(clk), .A(\g.we_clk [24515]));
Q_ASSIGN U8260 ( .B(clk), .A(\g.we_clk [24514]));
Q_ASSIGN U8261 ( .B(clk), .A(\g.we_clk [24513]));
Q_ASSIGN U8262 ( .B(clk), .A(\g.we_clk [24512]));
Q_ASSIGN U8263 ( .B(clk), .A(\g.we_clk [24511]));
Q_ASSIGN U8264 ( .B(clk), .A(\g.we_clk [24510]));
Q_ASSIGN U8265 ( .B(clk), .A(\g.we_clk [24509]));
Q_ASSIGN U8266 ( .B(clk), .A(\g.we_clk [24508]));
Q_ASSIGN U8267 ( .B(clk), .A(\g.we_clk [24507]));
Q_ASSIGN U8268 ( .B(clk), .A(\g.we_clk [24506]));
Q_ASSIGN U8269 ( .B(clk), .A(\g.we_clk [24505]));
Q_ASSIGN U8270 ( .B(clk), .A(\g.we_clk [24504]));
Q_ASSIGN U8271 ( .B(clk), .A(\g.we_clk [24503]));
Q_ASSIGN U8272 ( .B(clk), .A(\g.we_clk [24502]));
Q_ASSIGN U8273 ( .B(clk), .A(\g.we_clk [24501]));
Q_ASSIGN U8274 ( .B(clk), .A(\g.we_clk [24500]));
Q_ASSIGN U8275 ( .B(clk), .A(\g.we_clk [24499]));
Q_ASSIGN U8276 ( .B(clk), .A(\g.we_clk [24498]));
Q_ASSIGN U8277 ( .B(clk), .A(\g.we_clk [24497]));
Q_ASSIGN U8278 ( .B(clk), .A(\g.we_clk [24496]));
Q_ASSIGN U8279 ( .B(clk), .A(\g.we_clk [24495]));
Q_ASSIGN U8280 ( .B(clk), .A(\g.we_clk [24494]));
Q_ASSIGN U8281 ( .B(clk), .A(\g.we_clk [24493]));
Q_ASSIGN U8282 ( .B(clk), .A(\g.we_clk [24492]));
Q_ASSIGN U8283 ( .B(clk), .A(\g.we_clk [24491]));
Q_ASSIGN U8284 ( .B(clk), .A(\g.we_clk [24490]));
Q_ASSIGN U8285 ( .B(clk), .A(\g.we_clk [24489]));
Q_ASSIGN U8286 ( .B(clk), .A(\g.we_clk [24488]));
Q_ASSIGN U8287 ( .B(clk), .A(\g.we_clk [24487]));
Q_ASSIGN U8288 ( .B(clk), .A(\g.we_clk [24486]));
Q_ASSIGN U8289 ( .B(clk), .A(\g.we_clk [24485]));
Q_ASSIGN U8290 ( .B(clk), .A(\g.we_clk [24484]));
Q_ASSIGN U8291 ( .B(clk), .A(\g.we_clk [24483]));
Q_ASSIGN U8292 ( .B(clk), .A(\g.we_clk [24482]));
Q_ASSIGN U8293 ( .B(clk), .A(\g.we_clk [24481]));
Q_ASSIGN U8294 ( .B(clk), .A(\g.we_clk [24480]));
Q_ASSIGN U8295 ( .B(clk), .A(\g.we_clk [24479]));
Q_ASSIGN U8296 ( .B(clk), .A(\g.we_clk [24478]));
Q_ASSIGN U8297 ( .B(clk), .A(\g.we_clk [24477]));
Q_ASSIGN U8298 ( .B(clk), .A(\g.we_clk [24476]));
Q_ASSIGN U8299 ( .B(clk), .A(\g.we_clk [24475]));
Q_ASSIGN U8300 ( .B(clk), .A(\g.we_clk [24474]));
Q_ASSIGN U8301 ( .B(clk), .A(\g.we_clk [24473]));
Q_ASSIGN U8302 ( .B(clk), .A(\g.we_clk [24472]));
Q_ASSIGN U8303 ( .B(clk), .A(\g.we_clk [24471]));
Q_ASSIGN U8304 ( .B(clk), .A(\g.we_clk [24470]));
Q_ASSIGN U8305 ( .B(clk), .A(\g.we_clk [24469]));
Q_ASSIGN U8306 ( .B(clk), .A(\g.we_clk [24468]));
Q_ASSIGN U8307 ( .B(clk), .A(\g.we_clk [24467]));
Q_ASSIGN U8308 ( .B(clk), .A(\g.we_clk [24466]));
Q_ASSIGN U8309 ( .B(clk), .A(\g.we_clk [24465]));
Q_ASSIGN U8310 ( .B(clk), .A(\g.we_clk [24464]));
Q_ASSIGN U8311 ( .B(clk), .A(\g.we_clk [24463]));
Q_ASSIGN U8312 ( .B(clk), .A(\g.we_clk [24462]));
Q_ASSIGN U8313 ( .B(clk), .A(\g.we_clk [24461]));
Q_ASSIGN U8314 ( .B(clk), .A(\g.we_clk [24460]));
Q_ASSIGN U8315 ( .B(clk), .A(\g.we_clk [24459]));
Q_ASSIGN U8316 ( .B(clk), .A(\g.we_clk [24458]));
Q_ASSIGN U8317 ( .B(clk), .A(\g.we_clk [24457]));
Q_ASSIGN U8318 ( .B(clk), .A(\g.we_clk [24456]));
Q_ASSIGN U8319 ( .B(clk), .A(\g.we_clk [24455]));
Q_ASSIGN U8320 ( .B(clk), .A(\g.we_clk [24454]));
Q_ASSIGN U8321 ( .B(clk), .A(\g.we_clk [24453]));
Q_ASSIGN U8322 ( .B(clk), .A(\g.we_clk [24452]));
Q_ASSIGN U8323 ( .B(clk), .A(\g.we_clk [24451]));
Q_ASSIGN U8324 ( .B(clk), .A(\g.we_clk [24450]));
Q_ASSIGN U8325 ( .B(clk), .A(\g.we_clk [24449]));
Q_ASSIGN U8326 ( .B(clk), .A(\g.we_clk [24448]));
Q_ASSIGN U8327 ( .B(clk), .A(\g.we_clk [24447]));
Q_ASSIGN U8328 ( .B(clk), .A(\g.we_clk [24446]));
Q_ASSIGN U8329 ( .B(clk), .A(\g.we_clk [24445]));
Q_ASSIGN U8330 ( .B(clk), .A(\g.we_clk [24444]));
Q_ASSIGN U8331 ( .B(clk), .A(\g.we_clk [24443]));
Q_ASSIGN U8332 ( .B(clk), .A(\g.we_clk [24442]));
Q_ASSIGN U8333 ( .B(clk), .A(\g.we_clk [24441]));
Q_ASSIGN U8334 ( .B(clk), .A(\g.we_clk [24440]));
Q_ASSIGN U8335 ( .B(clk), .A(\g.we_clk [24439]));
Q_ASSIGN U8336 ( .B(clk), .A(\g.we_clk [24438]));
Q_ASSIGN U8337 ( .B(clk), .A(\g.we_clk [24437]));
Q_ASSIGN U8338 ( .B(clk), .A(\g.we_clk [24436]));
Q_ASSIGN U8339 ( .B(clk), .A(\g.we_clk [24435]));
Q_ASSIGN U8340 ( .B(clk), .A(\g.we_clk [24434]));
Q_ASSIGN U8341 ( .B(clk), .A(\g.we_clk [24433]));
Q_ASSIGN U8342 ( .B(clk), .A(\g.we_clk [24432]));
Q_ASSIGN U8343 ( .B(clk), .A(\g.we_clk [24431]));
Q_ASSIGN U8344 ( .B(clk), .A(\g.we_clk [24430]));
Q_ASSIGN U8345 ( .B(clk), .A(\g.we_clk [24429]));
Q_ASSIGN U8346 ( .B(clk), .A(\g.we_clk [24428]));
Q_ASSIGN U8347 ( .B(clk), .A(\g.we_clk [24427]));
Q_ASSIGN U8348 ( .B(clk), .A(\g.we_clk [24426]));
Q_ASSIGN U8349 ( .B(clk), .A(\g.we_clk [24425]));
Q_ASSIGN U8350 ( .B(clk), .A(\g.we_clk [24424]));
Q_ASSIGN U8351 ( .B(clk), .A(\g.we_clk [24423]));
Q_ASSIGN U8352 ( .B(clk), .A(\g.we_clk [24422]));
Q_ASSIGN U8353 ( .B(clk), .A(\g.we_clk [24421]));
Q_ASSIGN U8354 ( .B(clk), .A(\g.we_clk [24420]));
Q_ASSIGN U8355 ( .B(clk), .A(\g.we_clk [24419]));
Q_ASSIGN U8356 ( .B(clk), .A(\g.we_clk [24418]));
Q_ASSIGN U8357 ( .B(clk), .A(\g.we_clk [24417]));
Q_ASSIGN U8358 ( .B(clk), .A(\g.we_clk [24416]));
Q_ASSIGN U8359 ( .B(clk), .A(\g.we_clk [24415]));
Q_ASSIGN U8360 ( .B(clk), .A(\g.we_clk [24414]));
Q_ASSIGN U8361 ( .B(clk), .A(\g.we_clk [24413]));
Q_ASSIGN U8362 ( .B(clk), .A(\g.we_clk [24412]));
Q_ASSIGN U8363 ( .B(clk), .A(\g.we_clk [24411]));
Q_ASSIGN U8364 ( .B(clk), .A(\g.we_clk [24410]));
Q_ASSIGN U8365 ( .B(clk), .A(\g.we_clk [24409]));
Q_ASSIGN U8366 ( .B(clk), .A(\g.we_clk [24408]));
Q_ASSIGN U8367 ( .B(clk), .A(\g.we_clk [24407]));
Q_ASSIGN U8368 ( .B(clk), .A(\g.we_clk [24406]));
Q_ASSIGN U8369 ( .B(clk), .A(\g.we_clk [24405]));
Q_ASSIGN U8370 ( .B(clk), .A(\g.we_clk [24404]));
Q_ASSIGN U8371 ( .B(clk), .A(\g.we_clk [24403]));
Q_ASSIGN U8372 ( .B(clk), .A(\g.we_clk [24402]));
Q_ASSIGN U8373 ( .B(clk), .A(\g.we_clk [24401]));
Q_ASSIGN U8374 ( .B(clk), .A(\g.we_clk [24400]));
Q_ASSIGN U8375 ( .B(clk), .A(\g.we_clk [24399]));
Q_ASSIGN U8376 ( .B(clk), .A(\g.we_clk [24398]));
Q_ASSIGN U8377 ( .B(clk), .A(\g.we_clk [24397]));
Q_ASSIGN U8378 ( .B(clk), .A(\g.we_clk [24396]));
Q_ASSIGN U8379 ( .B(clk), .A(\g.we_clk [24395]));
Q_ASSIGN U8380 ( .B(clk), .A(\g.we_clk [24394]));
Q_ASSIGN U8381 ( .B(clk), .A(\g.we_clk [24393]));
Q_ASSIGN U8382 ( .B(clk), .A(\g.we_clk [24392]));
Q_ASSIGN U8383 ( .B(clk), .A(\g.we_clk [24391]));
Q_ASSIGN U8384 ( .B(clk), .A(\g.we_clk [24390]));
Q_ASSIGN U8385 ( .B(clk), .A(\g.we_clk [24389]));
Q_ASSIGN U8386 ( .B(clk), .A(\g.we_clk [24388]));
Q_ASSIGN U8387 ( .B(clk), .A(\g.we_clk [24387]));
Q_ASSIGN U8388 ( .B(clk), .A(\g.we_clk [24386]));
Q_ASSIGN U8389 ( .B(clk), .A(\g.we_clk [24385]));
Q_ASSIGN U8390 ( .B(clk), .A(\g.we_clk [24384]));
Q_ASSIGN U8391 ( .B(clk), .A(\g.we_clk [24383]));
Q_ASSIGN U8392 ( .B(clk), .A(\g.we_clk [24382]));
Q_ASSIGN U8393 ( .B(clk), .A(\g.we_clk [24381]));
Q_ASSIGN U8394 ( .B(clk), .A(\g.we_clk [24380]));
Q_ASSIGN U8395 ( .B(clk), .A(\g.we_clk [24379]));
Q_ASSIGN U8396 ( .B(clk), .A(\g.we_clk [24378]));
Q_ASSIGN U8397 ( .B(clk), .A(\g.we_clk [24377]));
Q_ASSIGN U8398 ( .B(clk), .A(\g.we_clk [24376]));
Q_ASSIGN U8399 ( .B(clk), .A(\g.we_clk [24375]));
Q_ASSIGN U8400 ( .B(clk), .A(\g.we_clk [24374]));
Q_ASSIGN U8401 ( .B(clk), .A(\g.we_clk [24373]));
Q_ASSIGN U8402 ( .B(clk), .A(\g.we_clk [24372]));
Q_ASSIGN U8403 ( .B(clk), .A(\g.we_clk [24371]));
Q_ASSIGN U8404 ( .B(clk), .A(\g.we_clk [24370]));
Q_ASSIGN U8405 ( .B(clk), .A(\g.we_clk [24369]));
Q_ASSIGN U8406 ( .B(clk), .A(\g.we_clk [24368]));
Q_ASSIGN U8407 ( .B(clk), .A(\g.we_clk [24367]));
Q_ASSIGN U8408 ( .B(clk), .A(\g.we_clk [24366]));
Q_ASSIGN U8409 ( .B(clk), .A(\g.we_clk [24365]));
Q_ASSIGN U8410 ( .B(clk), .A(\g.we_clk [24364]));
Q_ASSIGN U8411 ( .B(clk), .A(\g.we_clk [24363]));
Q_ASSIGN U8412 ( .B(clk), .A(\g.we_clk [24362]));
Q_ASSIGN U8413 ( .B(clk), .A(\g.we_clk [24361]));
Q_ASSIGN U8414 ( .B(clk), .A(\g.we_clk [24360]));
Q_ASSIGN U8415 ( .B(clk), .A(\g.we_clk [24359]));
Q_ASSIGN U8416 ( .B(clk), .A(\g.we_clk [24358]));
Q_ASSIGN U8417 ( .B(clk), .A(\g.we_clk [24357]));
Q_ASSIGN U8418 ( .B(clk), .A(\g.we_clk [24356]));
Q_ASSIGN U8419 ( .B(clk), .A(\g.we_clk [24355]));
Q_ASSIGN U8420 ( .B(clk), .A(\g.we_clk [24354]));
Q_ASSIGN U8421 ( .B(clk), .A(\g.we_clk [24353]));
Q_ASSIGN U8422 ( .B(clk), .A(\g.we_clk [24352]));
Q_ASSIGN U8423 ( .B(clk), .A(\g.we_clk [24351]));
Q_ASSIGN U8424 ( .B(clk), .A(\g.we_clk [24350]));
Q_ASSIGN U8425 ( .B(clk), .A(\g.we_clk [24349]));
Q_ASSIGN U8426 ( .B(clk), .A(\g.we_clk [24348]));
Q_ASSIGN U8427 ( .B(clk), .A(\g.we_clk [24347]));
Q_ASSIGN U8428 ( .B(clk), .A(\g.we_clk [24346]));
Q_ASSIGN U8429 ( .B(clk), .A(\g.we_clk [24345]));
Q_ASSIGN U8430 ( .B(clk), .A(\g.we_clk [24344]));
Q_ASSIGN U8431 ( .B(clk), .A(\g.we_clk [24343]));
Q_ASSIGN U8432 ( .B(clk), .A(\g.we_clk [24342]));
Q_ASSIGN U8433 ( .B(clk), .A(\g.we_clk [24341]));
Q_ASSIGN U8434 ( .B(clk), .A(\g.we_clk [24340]));
Q_ASSIGN U8435 ( .B(clk), .A(\g.we_clk [24339]));
Q_ASSIGN U8436 ( .B(clk), .A(\g.we_clk [24338]));
Q_ASSIGN U8437 ( .B(clk), .A(\g.we_clk [24337]));
Q_ASSIGN U8438 ( .B(clk), .A(\g.we_clk [24336]));
Q_ASSIGN U8439 ( .B(clk), .A(\g.we_clk [24335]));
Q_ASSIGN U8440 ( .B(clk), .A(\g.we_clk [24334]));
Q_ASSIGN U8441 ( .B(clk), .A(\g.we_clk [24333]));
Q_ASSIGN U8442 ( .B(clk), .A(\g.we_clk [24332]));
Q_ASSIGN U8443 ( .B(clk), .A(\g.we_clk [24331]));
Q_ASSIGN U8444 ( .B(clk), .A(\g.we_clk [24330]));
Q_ASSIGN U8445 ( .B(clk), .A(\g.we_clk [24329]));
Q_ASSIGN U8446 ( .B(clk), .A(\g.we_clk [24328]));
Q_ASSIGN U8447 ( .B(clk), .A(\g.we_clk [24327]));
Q_ASSIGN U8448 ( .B(clk), .A(\g.we_clk [24326]));
Q_ASSIGN U8449 ( .B(clk), .A(\g.we_clk [24325]));
Q_ASSIGN U8450 ( .B(clk), .A(\g.we_clk [24324]));
Q_ASSIGN U8451 ( .B(clk), .A(\g.we_clk [24323]));
Q_ASSIGN U8452 ( .B(clk), .A(\g.we_clk [24322]));
Q_ASSIGN U8453 ( .B(clk), .A(\g.we_clk [24321]));
Q_ASSIGN U8454 ( .B(clk), .A(\g.we_clk [24320]));
Q_ASSIGN U8455 ( .B(clk), .A(\g.we_clk [24319]));
Q_ASSIGN U8456 ( .B(clk), .A(\g.we_clk [24318]));
Q_ASSIGN U8457 ( .B(clk), .A(\g.we_clk [24317]));
Q_ASSIGN U8458 ( .B(clk), .A(\g.we_clk [24316]));
Q_ASSIGN U8459 ( .B(clk), .A(\g.we_clk [24315]));
Q_ASSIGN U8460 ( .B(clk), .A(\g.we_clk [24314]));
Q_ASSIGN U8461 ( .B(clk), .A(\g.we_clk [24313]));
Q_ASSIGN U8462 ( .B(clk), .A(\g.we_clk [24312]));
Q_ASSIGN U8463 ( .B(clk), .A(\g.we_clk [24311]));
Q_ASSIGN U8464 ( .B(clk), .A(\g.we_clk [24310]));
Q_ASSIGN U8465 ( .B(clk), .A(\g.we_clk [24309]));
Q_ASSIGN U8466 ( .B(clk), .A(\g.we_clk [24308]));
Q_ASSIGN U8467 ( .B(clk), .A(\g.we_clk [24307]));
Q_ASSIGN U8468 ( .B(clk), .A(\g.we_clk [24306]));
Q_ASSIGN U8469 ( .B(clk), .A(\g.we_clk [24305]));
Q_ASSIGN U8470 ( .B(clk), .A(\g.we_clk [24304]));
Q_ASSIGN U8471 ( .B(clk), .A(\g.we_clk [24303]));
Q_ASSIGN U8472 ( .B(clk), .A(\g.we_clk [24302]));
Q_ASSIGN U8473 ( .B(clk), .A(\g.we_clk [24301]));
Q_ASSIGN U8474 ( .B(clk), .A(\g.we_clk [24300]));
Q_ASSIGN U8475 ( .B(clk), .A(\g.we_clk [24299]));
Q_ASSIGN U8476 ( .B(clk), .A(\g.we_clk [24298]));
Q_ASSIGN U8477 ( .B(clk), .A(\g.we_clk [24297]));
Q_ASSIGN U8478 ( .B(clk), .A(\g.we_clk [24296]));
Q_ASSIGN U8479 ( .B(clk), .A(\g.we_clk [24295]));
Q_ASSIGN U8480 ( .B(clk), .A(\g.we_clk [24294]));
Q_ASSIGN U8481 ( .B(clk), .A(\g.we_clk [24293]));
Q_ASSIGN U8482 ( .B(clk), .A(\g.we_clk [24292]));
Q_ASSIGN U8483 ( .B(clk), .A(\g.we_clk [24291]));
Q_ASSIGN U8484 ( .B(clk), .A(\g.we_clk [24290]));
Q_ASSIGN U8485 ( .B(clk), .A(\g.we_clk [24289]));
Q_ASSIGN U8486 ( .B(clk), .A(\g.we_clk [24288]));
Q_ASSIGN U8487 ( .B(clk), .A(\g.we_clk [24287]));
Q_ASSIGN U8488 ( .B(clk), .A(\g.we_clk [24286]));
Q_ASSIGN U8489 ( .B(clk), .A(\g.we_clk [24285]));
Q_ASSIGN U8490 ( .B(clk), .A(\g.we_clk [24284]));
Q_ASSIGN U8491 ( .B(clk), .A(\g.we_clk [24283]));
Q_ASSIGN U8492 ( .B(clk), .A(\g.we_clk [24282]));
Q_ASSIGN U8493 ( .B(clk), .A(\g.we_clk [24281]));
Q_ASSIGN U8494 ( .B(clk), .A(\g.we_clk [24280]));
Q_ASSIGN U8495 ( .B(clk), .A(\g.we_clk [24279]));
Q_ASSIGN U8496 ( .B(clk), .A(\g.we_clk [24278]));
Q_ASSIGN U8497 ( .B(clk), .A(\g.we_clk [24277]));
Q_ASSIGN U8498 ( .B(clk), .A(\g.we_clk [24276]));
Q_ASSIGN U8499 ( .B(clk), .A(\g.we_clk [24275]));
Q_ASSIGN U8500 ( .B(clk), .A(\g.we_clk [24274]));
Q_ASSIGN U8501 ( .B(clk), .A(\g.we_clk [24273]));
Q_ASSIGN U8502 ( .B(clk), .A(\g.we_clk [24272]));
Q_ASSIGN U8503 ( .B(clk), .A(\g.we_clk [24271]));
Q_ASSIGN U8504 ( .B(clk), .A(\g.we_clk [24270]));
Q_ASSIGN U8505 ( .B(clk), .A(\g.we_clk [24269]));
Q_ASSIGN U8506 ( .B(clk), .A(\g.we_clk [24268]));
Q_ASSIGN U8507 ( .B(clk), .A(\g.we_clk [24267]));
Q_ASSIGN U8508 ( .B(clk), .A(\g.we_clk [24266]));
Q_ASSIGN U8509 ( .B(clk), .A(\g.we_clk [24265]));
Q_ASSIGN U8510 ( .B(clk), .A(\g.we_clk [24264]));
Q_ASSIGN U8511 ( .B(clk), .A(\g.we_clk [24263]));
Q_ASSIGN U8512 ( .B(clk), .A(\g.we_clk [24262]));
Q_ASSIGN U8513 ( .B(clk), .A(\g.we_clk [24261]));
Q_ASSIGN U8514 ( .B(clk), .A(\g.we_clk [24260]));
Q_ASSIGN U8515 ( .B(clk), .A(\g.we_clk [24259]));
Q_ASSIGN U8516 ( .B(clk), .A(\g.we_clk [24258]));
Q_ASSIGN U8517 ( .B(clk), .A(\g.we_clk [24257]));
Q_ASSIGN U8518 ( .B(clk), .A(\g.we_clk [24256]));
Q_ASSIGN U8519 ( .B(clk), .A(\g.we_clk [24255]));
Q_ASSIGN U8520 ( .B(clk), .A(\g.we_clk [24254]));
Q_ASSIGN U8521 ( .B(clk), .A(\g.we_clk [24253]));
Q_ASSIGN U8522 ( .B(clk), .A(\g.we_clk [24252]));
Q_ASSIGN U8523 ( .B(clk), .A(\g.we_clk [24251]));
Q_ASSIGN U8524 ( .B(clk), .A(\g.we_clk [24250]));
Q_ASSIGN U8525 ( .B(clk), .A(\g.we_clk [24249]));
Q_ASSIGN U8526 ( .B(clk), .A(\g.we_clk [24248]));
Q_ASSIGN U8527 ( .B(clk), .A(\g.we_clk [24247]));
Q_ASSIGN U8528 ( .B(clk), .A(\g.we_clk [24246]));
Q_ASSIGN U8529 ( .B(clk), .A(\g.we_clk [24245]));
Q_ASSIGN U8530 ( .B(clk), .A(\g.we_clk [24244]));
Q_ASSIGN U8531 ( .B(clk), .A(\g.we_clk [24243]));
Q_ASSIGN U8532 ( .B(clk), .A(\g.we_clk [24242]));
Q_ASSIGN U8533 ( .B(clk), .A(\g.we_clk [24241]));
Q_ASSIGN U8534 ( .B(clk), .A(\g.we_clk [24240]));
Q_ASSIGN U8535 ( .B(clk), .A(\g.we_clk [24239]));
Q_ASSIGN U8536 ( .B(clk), .A(\g.we_clk [24238]));
Q_ASSIGN U8537 ( .B(clk), .A(\g.we_clk [24237]));
Q_ASSIGN U8538 ( .B(clk), .A(\g.we_clk [24236]));
Q_ASSIGN U8539 ( .B(clk), .A(\g.we_clk [24235]));
Q_ASSIGN U8540 ( .B(clk), .A(\g.we_clk [24234]));
Q_ASSIGN U8541 ( .B(clk), .A(\g.we_clk [24233]));
Q_ASSIGN U8542 ( .B(clk), .A(\g.we_clk [24232]));
Q_ASSIGN U8543 ( .B(clk), .A(\g.we_clk [24231]));
Q_ASSIGN U8544 ( .B(clk), .A(\g.we_clk [24230]));
Q_ASSIGN U8545 ( .B(clk), .A(\g.we_clk [24229]));
Q_ASSIGN U8546 ( .B(clk), .A(\g.we_clk [24228]));
Q_ASSIGN U8547 ( .B(clk), .A(\g.we_clk [24227]));
Q_ASSIGN U8548 ( .B(clk), .A(\g.we_clk [24226]));
Q_ASSIGN U8549 ( .B(clk), .A(\g.we_clk [24225]));
Q_ASSIGN U8550 ( .B(clk), .A(\g.we_clk [24224]));
Q_ASSIGN U8551 ( .B(clk), .A(\g.we_clk [24223]));
Q_ASSIGN U8552 ( .B(clk), .A(\g.we_clk [24222]));
Q_ASSIGN U8553 ( .B(clk), .A(\g.we_clk [24221]));
Q_ASSIGN U8554 ( .B(clk), .A(\g.we_clk [24220]));
Q_ASSIGN U8555 ( .B(clk), .A(\g.we_clk [24219]));
Q_ASSIGN U8556 ( .B(clk), .A(\g.we_clk [24218]));
Q_ASSIGN U8557 ( .B(clk), .A(\g.we_clk [24217]));
Q_ASSIGN U8558 ( .B(clk), .A(\g.we_clk [24216]));
Q_ASSIGN U8559 ( .B(clk), .A(\g.we_clk [24215]));
Q_ASSIGN U8560 ( .B(clk), .A(\g.we_clk [24214]));
Q_ASSIGN U8561 ( .B(clk), .A(\g.we_clk [24213]));
Q_ASSIGN U8562 ( .B(clk), .A(\g.we_clk [24212]));
Q_ASSIGN U8563 ( .B(clk), .A(\g.we_clk [24211]));
Q_ASSIGN U8564 ( .B(clk), .A(\g.we_clk [24210]));
Q_ASSIGN U8565 ( .B(clk), .A(\g.we_clk [24209]));
Q_ASSIGN U8566 ( .B(clk), .A(\g.we_clk [24208]));
Q_ASSIGN U8567 ( .B(clk), .A(\g.we_clk [24207]));
Q_ASSIGN U8568 ( .B(clk), .A(\g.we_clk [24206]));
Q_ASSIGN U8569 ( .B(clk), .A(\g.we_clk [24205]));
Q_ASSIGN U8570 ( .B(clk), .A(\g.we_clk [24204]));
Q_ASSIGN U8571 ( .B(clk), .A(\g.we_clk [24203]));
Q_ASSIGN U8572 ( .B(clk), .A(\g.we_clk [24202]));
Q_ASSIGN U8573 ( .B(clk), .A(\g.we_clk [24201]));
Q_ASSIGN U8574 ( .B(clk), .A(\g.we_clk [24200]));
Q_ASSIGN U8575 ( .B(clk), .A(\g.we_clk [24199]));
Q_ASSIGN U8576 ( .B(clk), .A(\g.we_clk [24198]));
Q_ASSIGN U8577 ( .B(clk), .A(\g.we_clk [24197]));
Q_ASSIGN U8578 ( .B(clk), .A(\g.we_clk [24196]));
Q_ASSIGN U8579 ( .B(clk), .A(\g.we_clk [24195]));
Q_ASSIGN U8580 ( .B(clk), .A(\g.we_clk [24194]));
Q_ASSIGN U8581 ( .B(clk), .A(\g.we_clk [24193]));
Q_ASSIGN U8582 ( .B(clk), .A(\g.we_clk [24192]));
Q_ASSIGN U8583 ( .B(clk), .A(\g.we_clk [24191]));
Q_ASSIGN U8584 ( .B(clk), .A(\g.we_clk [24190]));
Q_ASSIGN U8585 ( .B(clk), .A(\g.we_clk [24189]));
Q_ASSIGN U8586 ( .B(clk), .A(\g.we_clk [24188]));
Q_ASSIGN U8587 ( .B(clk), .A(\g.we_clk [24187]));
Q_ASSIGN U8588 ( .B(clk), .A(\g.we_clk [24186]));
Q_ASSIGN U8589 ( .B(clk), .A(\g.we_clk [24185]));
Q_ASSIGN U8590 ( .B(clk), .A(\g.we_clk [24184]));
Q_ASSIGN U8591 ( .B(clk), .A(\g.we_clk [24183]));
Q_ASSIGN U8592 ( .B(clk), .A(\g.we_clk [24182]));
Q_ASSIGN U8593 ( .B(clk), .A(\g.we_clk [24181]));
Q_ASSIGN U8594 ( .B(clk), .A(\g.we_clk [24180]));
Q_ASSIGN U8595 ( .B(clk), .A(\g.we_clk [24179]));
Q_ASSIGN U8596 ( .B(clk), .A(\g.we_clk [24178]));
Q_ASSIGN U8597 ( .B(clk), .A(\g.we_clk [24177]));
Q_ASSIGN U8598 ( .B(clk), .A(\g.we_clk [24176]));
Q_ASSIGN U8599 ( .B(clk), .A(\g.we_clk [24175]));
Q_ASSIGN U8600 ( .B(clk), .A(\g.we_clk [24174]));
Q_ASSIGN U8601 ( .B(clk), .A(\g.we_clk [24173]));
Q_ASSIGN U8602 ( .B(clk), .A(\g.we_clk [24172]));
Q_ASSIGN U8603 ( .B(clk), .A(\g.we_clk [24171]));
Q_ASSIGN U8604 ( .B(clk), .A(\g.we_clk [24170]));
Q_ASSIGN U8605 ( .B(clk), .A(\g.we_clk [24169]));
Q_ASSIGN U8606 ( .B(clk), .A(\g.we_clk [24168]));
Q_ASSIGN U8607 ( .B(clk), .A(\g.we_clk [24167]));
Q_ASSIGN U8608 ( .B(clk), .A(\g.we_clk [24166]));
Q_ASSIGN U8609 ( .B(clk), .A(\g.we_clk [24165]));
Q_ASSIGN U8610 ( .B(clk), .A(\g.we_clk [24164]));
Q_ASSIGN U8611 ( .B(clk), .A(\g.we_clk [24163]));
Q_ASSIGN U8612 ( .B(clk), .A(\g.we_clk [24162]));
Q_ASSIGN U8613 ( .B(clk), .A(\g.we_clk [24161]));
Q_ASSIGN U8614 ( .B(clk), .A(\g.we_clk [24160]));
Q_ASSIGN U8615 ( .B(clk), .A(\g.we_clk [24159]));
Q_ASSIGN U8616 ( .B(clk), .A(\g.we_clk [24158]));
Q_ASSIGN U8617 ( .B(clk), .A(\g.we_clk [24157]));
Q_ASSIGN U8618 ( .B(clk), .A(\g.we_clk [24156]));
Q_ASSIGN U8619 ( .B(clk), .A(\g.we_clk [24155]));
Q_ASSIGN U8620 ( .B(clk), .A(\g.we_clk [24154]));
Q_ASSIGN U8621 ( .B(clk), .A(\g.we_clk [24153]));
Q_ASSIGN U8622 ( .B(clk), .A(\g.we_clk [24152]));
Q_ASSIGN U8623 ( .B(clk), .A(\g.we_clk [24151]));
Q_ASSIGN U8624 ( .B(clk), .A(\g.we_clk [24150]));
Q_ASSIGN U8625 ( .B(clk), .A(\g.we_clk [24149]));
Q_ASSIGN U8626 ( .B(clk), .A(\g.we_clk [24148]));
Q_ASSIGN U8627 ( .B(clk), .A(\g.we_clk [24147]));
Q_ASSIGN U8628 ( .B(clk), .A(\g.we_clk [24146]));
Q_ASSIGN U8629 ( .B(clk), .A(\g.we_clk [24145]));
Q_ASSIGN U8630 ( .B(clk), .A(\g.we_clk [24144]));
Q_ASSIGN U8631 ( .B(clk), .A(\g.we_clk [24143]));
Q_ASSIGN U8632 ( .B(clk), .A(\g.we_clk [24142]));
Q_ASSIGN U8633 ( .B(clk), .A(\g.we_clk [24141]));
Q_ASSIGN U8634 ( .B(clk), .A(\g.we_clk [24140]));
Q_ASSIGN U8635 ( .B(clk), .A(\g.we_clk [24139]));
Q_ASSIGN U8636 ( .B(clk), .A(\g.we_clk [24138]));
Q_ASSIGN U8637 ( .B(clk), .A(\g.we_clk [24137]));
Q_ASSIGN U8638 ( .B(clk), .A(\g.we_clk [24136]));
Q_ASSIGN U8639 ( .B(clk), .A(\g.we_clk [24135]));
Q_ASSIGN U8640 ( .B(clk), .A(\g.we_clk [24134]));
Q_ASSIGN U8641 ( .B(clk), .A(\g.we_clk [24133]));
Q_ASSIGN U8642 ( .B(clk), .A(\g.we_clk [24132]));
Q_ASSIGN U8643 ( .B(clk), .A(\g.we_clk [24131]));
Q_ASSIGN U8644 ( .B(clk), .A(\g.we_clk [24130]));
Q_ASSIGN U8645 ( .B(clk), .A(\g.we_clk [24129]));
Q_ASSIGN U8646 ( .B(clk), .A(\g.we_clk [24128]));
Q_ASSIGN U8647 ( .B(clk), .A(\g.we_clk [24127]));
Q_ASSIGN U8648 ( .B(clk), .A(\g.we_clk [24126]));
Q_ASSIGN U8649 ( .B(clk), .A(\g.we_clk [24125]));
Q_ASSIGN U8650 ( .B(clk), .A(\g.we_clk [24124]));
Q_ASSIGN U8651 ( .B(clk), .A(\g.we_clk [24123]));
Q_ASSIGN U8652 ( .B(clk), .A(\g.we_clk [24122]));
Q_ASSIGN U8653 ( .B(clk), .A(\g.we_clk [24121]));
Q_ASSIGN U8654 ( .B(clk), .A(\g.we_clk [24120]));
Q_ASSIGN U8655 ( .B(clk), .A(\g.we_clk [24119]));
Q_ASSIGN U8656 ( .B(clk), .A(\g.we_clk [24118]));
Q_ASSIGN U8657 ( .B(clk), .A(\g.we_clk [24117]));
Q_ASSIGN U8658 ( .B(clk), .A(\g.we_clk [24116]));
Q_ASSIGN U8659 ( .B(clk), .A(\g.we_clk [24115]));
Q_ASSIGN U8660 ( .B(clk), .A(\g.we_clk [24114]));
Q_ASSIGN U8661 ( .B(clk), .A(\g.we_clk [24113]));
Q_ASSIGN U8662 ( .B(clk), .A(\g.we_clk [24112]));
Q_ASSIGN U8663 ( .B(clk), .A(\g.we_clk [24111]));
Q_ASSIGN U8664 ( .B(clk), .A(\g.we_clk [24110]));
Q_ASSIGN U8665 ( .B(clk), .A(\g.we_clk [24109]));
Q_ASSIGN U8666 ( .B(clk), .A(\g.we_clk [24108]));
Q_ASSIGN U8667 ( .B(clk), .A(\g.we_clk [24107]));
Q_ASSIGN U8668 ( .B(clk), .A(\g.we_clk [24106]));
Q_ASSIGN U8669 ( .B(clk), .A(\g.we_clk [24105]));
Q_ASSIGN U8670 ( .B(clk), .A(\g.we_clk [24104]));
Q_ASSIGN U8671 ( .B(clk), .A(\g.we_clk [24103]));
Q_ASSIGN U8672 ( .B(clk), .A(\g.we_clk [24102]));
Q_ASSIGN U8673 ( .B(clk), .A(\g.we_clk [24101]));
Q_ASSIGN U8674 ( .B(clk), .A(\g.we_clk [24100]));
Q_ASSIGN U8675 ( .B(clk), .A(\g.we_clk [24099]));
Q_ASSIGN U8676 ( .B(clk), .A(\g.we_clk [24098]));
Q_ASSIGN U8677 ( .B(clk), .A(\g.we_clk [24097]));
Q_ASSIGN U8678 ( .B(clk), .A(\g.we_clk [24096]));
Q_ASSIGN U8679 ( .B(clk), .A(\g.we_clk [24095]));
Q_ASSIGN U8680 ( .B(clk), .A(\g.we_clk [24094]));
Q_ASSIGN U8681 ( .B(clk), .A(\g.we_clk [24093]));
Q_ASSIGN U8682 ( .B(clk), .A(\g.we_clk [24092]));
Q_ASSIGN U8683 ( .B(clk), .A(\g.we_clk [24091]));
Q_ASSIGN U8684 ( .B(clk), .A(\g.we_clk [24090]));
Q_ASSIGN U8685 ( .B(clk), .A(\g.we_clk [24089]));
Q_ASSIGN U8686 ( .B(clk), .A(\g.we_clk [24088]));
Q_ASSIGN U8687 ( .B(clk), .A(\g.we_clk [24087]));
Q_ASSIGN U8688 ( .B(clk), .A(\g.we_clk [24086]));
Q_ASSIGN U8689 ( .B(clk), .A(\g.we_clk [24085]));
Q_ASSIGN U8690 ( .B(clk), .A(\g.we_clk [24084]));
Q_ASSIGN U8691 ( .B(clk), .A(\g.we_clk [24083]));
Q_ASSIGN U8692 ( .B(clk), .A(\g.we_clk [24082]));
Q_ASSIGN U8693 ( .B(clk), .A(\g.we_clk [24081]));
Q_ASSIGN U8694 ( .B(clk), .A(\g.we_clk [24080]));
Q_ASSIGN U8695 ( .B(clk), .A(\g.we_clk [24079]));
Q_ASSIGN U8696 ( .B(clk), .A(\g.we_clk [24078]));
Q_ASSIGN U8697 ( .B(clk), .A(\g.we_clk [24077]));
Q_ASSIGN U8698 ( .B(clk), .A(\g.we_clk [24076]));
Q_ASSIGN U8699 ( .B(clk), .A(\g.we_clk [24075]));
Q_ASSIGN U8700 ( .B(clk), .A(\g.we_clk [24074]));
Q_ASSIGN U8701 ( .B(clk), .A(\g.we_clk [24073]));
Q_ASSIGN U8702 ( .B(clk), .A(\g.we_clk [24072]));
Q_ASSIGN U8703 ( .B(clk), .A(\g.we_clk [24071]));
Q_ASSIGN U8704 ( .B(clk), .A(\g.we_clk [24070]));
Q_ASSIGN U8705 ( .B(clk), .A(\g.we_clk [24069]));
Q_ASSIGN U8706 ( .B(clk), .A(\g.we_clk [24068]));
Q_ASSIGN U8707 ( .B(clk), .A(\g.we_clk [24067]));
Q_ASSIGN U8708 ( .B(clk), .A(\g.we_clk [24066]));
Q_ASSIGN U8709 ( .B(clk), .A(\g.we_clk [24065]));
Q_ASSIGN U8710 ( .B(clk), .A(\g.we_clk [24064]));
Q_ASSIGN U8711 ( .B(clk), .A(\g.we_clk [24063]));
Q_ASSIGN U8712 ( .B(clk), .A(\g.we_clk [24062]));
Q_ASSIGN U8713 ( .B(clk), .A(\g.we_clk [24061]));
Q_ASSIGN U8714 ( .B(clk), .A(\g.we_clk [24060]));
Q_ASSIGN U8715 ( .B(clk), .A(\g.we_clk [24059]));
Q_ASSIGN U8716 ( .B(clk), .A(\g.we_clk [24058]));
Q_ASSIGN U8717 ( .B(clk), .A(\g.we_clk [24057]));
Q_ASSIGN U8718 ( .B(clk), .A(\g.we_clk [24056]));
Q_ASSIGN U8719 ( .B(clk), .A(\g.we_clk [24055]));
Q_ASSIGN U8720 ( .B(clk), .A(\g.we_clk [24054]));
Q_ASSIGN U8721 ( .B(clk), .A(\g.we_clk [24053]));
Q_ASSIGN U8722 ( .B(clk), .A(\g.we_clk [24052]));
Q_ASSIGN U8723 ( .B(clk), .A(\g.we_clk [24051]));
Q_ASSIGN U8724 ( .B(clk), .A(\g.we_clk [24050]));
Q_ASSIGN U8725 ( .B(clk), .A(\g.we_clk [24049]));
Q_ASSIGN U8726 ( .B(clk), .A(\g.we_clk [24048]));
Q_ASSIGN U8727 ( .B(clk), .A(\g.we_clk [24047]));
Q_ASSIGN U8728 ( .B(clk), .A(\g.we_clk [24046]));
Q_ASSIGN U8729 ( .B(clk), .A(\g.we_clk [24045]));
Q_ASSIGN U8730 ( .B(clk), .A(\g.we_clk [24044]));
Q_ASSIGN U8731 ( .B(clk), .A(\g.we_clk [24043]));
Q_ASSIGN U8732 ( .B(clk), .A(\g.we_clk [24042]));
Q_ASSIGN U8733 ( .B(clk), .A(\g.we_clk [24041]));
Q_ASSIGN U8734 ( .B(clk), .A(\g.we_clk [24040]));
Q_ASSIGN U8735 ( .B(clk), .A(\g.we_clk [24039]));
Q_ASSIGN U8736 ( .B(clk), .A(\g.we_clk [24038]));
Q_ASSIGN U8737 ( .B(clk), .A(\g.we_clk [24037]));
Q_ASSIGN U8738 ( .B(clk), .A(\g.we_clk [24036]));
Q_ASSIGN U8739 ( .B(clk), .A(\g.we_clk [24035]));
Q_ASSIGN U8740 ( .B(clk), .A(\g.we_clk [24034]));
Q_ASSIGN U8741 ( .B(clk), .A(\g.we_clk [24033]));
Q_ASSIGN U8742 ( .B(clk), .A(\g.we_clk [24032]));
Q_ASSIGN U8743 ( .B(clk), .A(\g.we_clk [24031]));
Q_ASSIGN U8744 ( .B(clk), .A(\g.we_clk [24030]));
Q_ASSIGN U8745 ( .B(clk), .A(\g.we_clk [24029]));
Q_ASSIGN U8746 ( .B(clk), .A(\g.we_clk [24028]));
Q_ASSIGN U8747 ( .B(clk), .A(\g.we_clk [24027]));
Q_ASSIGN U8748 ( .B(clk), .A(\g.we_clk [24026]));
Q_ASSIGN U8749 ( .B(clk), .A(\g.we_clk [24025]));
Q_ASSIGN U8750 ( .B(clk), .A(\g.we_clk [24024]));
Q_ASSIGN U8751 ( .B(clk), .A(\g.we_clk [24023]));
Q_ASSIGN U8752 ( .B(clk), .A(\g.we_clk [24022]));
Q_ASSIGN U8753 ( .B(clk), .A(\g.we_clk [24021]));
Q_ASSIGN U8754 ( .B(clk), .A(\g.we_clk [24020]));
Q_ASSIGN U8755 ( .B(clk), .A(\g.we_clk [24019]));
Q_ASSIGN U8756 ( .B(clk), .A(\g.we_clk [24018]));
Q_ASSIGN U8757 ( .B(clk), .A(\g.we_clk [24017]));
Q_ASSIGN U8758 ( .B(clk), .A(\g.we_clk [24016]));
Q_ASSIGN U8759 ( .B(clk), .A(\g.we_clk [24015]));
Q_ASSIGN U8760 ( .B(clk), .A(\g.we_clk [24014]));
Q_ASSIGN U8761 ( .B(clk), .A(\g.we_clk [24013]));
Q_ASSIGN U8762 ( .B(clk), .A(\g.we_clk [24012]));
Q_ASSIGN U8763 ( .B(clk), .A(\g.we_clk [24011]));
Q_ASSIGN U8764 ( .B(clk), .A(\g.we_clk [24010]));
Q_ASSIGN U8765 ( .B(clk), .A(\g.we_clk [24009]));
Q_ASSIGN U8766 ( .B(clk), .A(\g.we_clk [24008]));
Q_ASSIGN U8767 ( .B(clk), .A(\g.we_clk [24007]));
Q_ASSIGN U8768 ( .B(clk), .A(\g.we_clk [24006]));
Q_ASSIGN U8769 ( .B(clk), .A(\g.we_clk [24005]));
Q_ASSIGN U8770 ( .B(clk), .A(\g.we_clk [24004]));
Q_ASSIGN U8771 ( .B(clk), .A(\g.we_clk [24003]));
Q_ASSIGN U8772 ( .B(clk), .A(\g.we_clk [24002]));
Q_ASSIGN U8773 ( .B(clk), .A(\g.we_clk [24001]));
Q_ASSIGN U8774 ( .B(clk), .A(\g.we_clk [24000]));
Q_ASSIGN U8775 ( .B(clk), .A(\g.we_clk [23999]));
Q_ASSIGN U8776 ( .B(clk), .A(\g.we_clk [23998]));
Q_ASSIGN U8777 ( .B(clk), .A(\g.we_clk [23997]));
Q_ASSIGN U8778 ( .B(clk), .A(\g.we_clk [23996]));
Q_ASSIGN U8779 ( .B(clk), .A(\g.we_clk [23995]));
Q_ASSIGN U8780 ( .B(clk), .A(\g.we_clk [23994]));
Q_ASSIGN U8781 ( .B(clk), .A(\g.we_clk [23993]));
Q_ASSIGN U8782 ( .B(clk), .A(\g.we_clk [23992]));
Q_ASSIGN U8783 ( .B(clk), .A(\g.we_clk [23991]));
Q_ASSIGN U8784 ( .B(clk), .A(\g.we_clk [23990]));
Q_ASSIGN U8785 ( .B(clk), .A(\g.we_clk [23989]));
Q_ASSIGN U8786 ( .B(clk), .A(\g.we_clk [23988]));
Q_ASSIGN U8787 ( .B(clk), .A(\g.we_clk [23987]));
Q_ASSIGN U8788 ( .B(clk), .A(\g.we_clk [23986]));
Q_ASSIGN U8789 ( .B(clk), .A(\g.we_clk [23985]));
Q_ASSIGN U8790 ( .B(clk), .A(\g.we_clk [23984]));
Q_ASSIGN U8791 ( .B(clk), .A(\g.we_clk [23983]));
Q_ASSIGN U8792 ( .B(clk), .A(\g.we_clk [23982]));
Q_ASSIGN U8793 ( .B(clk), .A(\g.we_clk [23981]));
Q_ASSIGN U8794 ( .B(clk), .A(\g.we_clk [23980]));
Q_ASSIGN U8795 ( .B(clk), .A(\g.we_clk [23979]));
Q_ASSIGN U8796 ( .B(clk), .A(\g.we_clk [23978]));
Q_ASSIGN U8797 ( .B(clk), .A(\g.we_clk [23977]));
Q_ASSIGN U8798 ( .B(clk), .A(\g.we_clk [23976]));
Q_ASSIGN U8799 ( .B(clk), .A(\g.we_clk [23975]));
Q_ASSIGN U8800 ( .B(clk), .A(\g.we_clk [23974]));
Q_ASSIGN U8801 ( .B(clk), .A(\g.we_clk [23973]));
Q_ASSIGN U8802 ( .B(clk), .A(\g.we_clk [23972]));
Q_ASSIGN U8803 ( .B(clk), .A(\g.we_clk [23971]));
Q_ASSIGN U8804 ( .B(clk), .A(\g.we_clk [23970]));
Q_ASSIGN U8805 ( .B(clk), .A(\g.we_clk [23969]));
Q_ASSIGN U8806 ( .B(clk), .A(\g.we_clk [23968]));
Q_ASSIGN U8807 ( .B(clk), .A(\g.we_clk [23967]));
Q_ASSIGN U8808 ( .B(clk), .A(\g.we_clk [23966]));
Q_ASSIGN U8809 ( .B(clk), .A(\g.we_clk [23965]));
Q_ASSIGN U8810 ( .B(clk), .A(\g.we_clk [23964]));
Q_ASSIGN U8811 ( .B(clk), .A(\g.we_clk [23963]));
Q_ASSIGN U8812 ( .B(clk), .A(\g.we_clk [23962]));
Q_ASSIGN U8813 ( .B(clk), .A(\g.we_clk [23961]));
Q_ASSIGN U8814 ( .B(clk), .A(\g.we_clk [23960]));
Q_ASSIGN U8815 ( .B(clk), .A(\g.we_clk [23959]));
Q_ASSIGN U8816 ( .B(clk), .A(\g.we_clk [23958]));
Q_ASSIGN U8817 ( .B(clk), .A(\g.we_clk [23957]));
Q_ASSIGN U8818 ( .B(clk), .A(\g.we_clk [23956]));
Q_ASSIGN U8819 ( .B(clk), .A(\g.we_clk [23955]));
Q_ASSIGN U8820 ( .B(clk), .A(\g.we_clk [23954]));
Q_ASSIGN U8821 ( .B(clk), .A(\g.we_clk [23953]));
Q_ASSIGN U8822 ( .B(clk), .A(\g.we_clk [23952]));
Q_ASSIGN U8823 ( .B(clk), .A(\g.we_clk [23951]));
Q_ASSIGN U8824 ( .B(clk), .A(\g.we_clk [23950]));
Q_ASSIGN U8825 ( .B(clk), .A(\g.we_clk [23949]));
Q_ASSIGN U8826 ( .B(clk), .A(\g.we_clk [23948]));
Q_ASSIGN U8827 ( .B(clk), .A(\g.we_clk [23947]));
Q_ASSIGN U8828 ( .B(clk), .A(\g.we_clk [23946]));
Q_ASSIGN U8829 ( .B(clk), .A(\g.we_clk [23945]));
Q_ASSIGN U8830 ( .B(clk), .A(\g.we_clk [23944]));
Q_ASSIGN U8831 ( .B(clk), .A(\g.we_clk [23943]));
Q_ASSIGN U8832 ( .B(clk), .A(\g.we_clk [23942]));
Q_ASSIGN U8833 ( .B(clk), .A(\g.we_clk [23941]));
Q_ASSIGN U8834 ( .B(clk), .A(\g.we_clk [23940]));
Q_ASSIGN U8835 ( .B(clk), .A(\g.we_clk [23939]));
Q_ASSIGN U8836 ( .B(clk), .A(\g.we_clk [23938]));
Q_ASSIGN U8837 ( .B(clk), .A(\g.we_clk [23937]));
Q_ASSIGN U8838 ( .B(clk), .A(\g.we_clk [23936]));
Q_ASSIGN U8839 ( .B(clk), .A(\g.we_clk [23935]));
Q_ASSIGN U8840 ( .B(clk), .A(\g.we_clk [23934]));
Q_ASSIGN U8841 ( .B(clk), .A(\g.we_clk [23933]));
Q_ASSIGN U8842 ( .B(clk), .A(\g.we_clk [23932]));
Q_ASSIGN U8843 ( .B(clk), .A(\g.we_clk [23931]));
Q_ASSIGN U8844 ( .B(clk), .A(\g.we_clk [23930]));
Q_ASSIGN U8845 ( .B(clk), .A(\g.we_clk [23929]));
Q_ASSIGN U8846 ( .B(clk), .A(\g.we_clk [23928]));
Q_ASSIGN U8847 ( .B(clk), .A(\g.we_clk [23927]));
Q_ASSIGN U8848 ( .B(clk), .A(\g.we_clk [23926]));
Q_ASSIGN U8849 ( .B(clk), .A(\g.we_clk [23925]));
Q_ASSIGN U8850 ( .B(clk), .A(\g.we_clk [23924]));
Q_ASSIGN U8851 ( .B(clk), .A(\g.we_clk [23923]));
Q_ASSIGN U8852 ( .B(clk), .A(\g.we_clk [23922]));
Q_ASSIGN U8853 ( .B(clk), .A(\g.we_clk [23921]));
Q_ASSIGN U8854 ( .B(clk), .A(\g.we_clk [23920]));
Q_ASSIGN U8855 ( .B(clk), .A(\g.we_clk [23919]));
Q_ASSIGN U8856 ( .B(clk), .A(\g.we_clk [23918]));
Q_ASSIGN U8857 ( .B(clk), .A(\g.we_clk [23917]));
Q_ASSIGN U8858 ( .B(clk), .A(\g.we_clk [23916]));
Q_ASSIGN U8859 ( .B(clk), .A(\g.we_clk [23915]));
Q_ASSIGN U8860 ( .B(clk), .A(\g.we_clk [23914]));
Q_ASSIGN U8861 ( .B(clk), .A(\g.we_clk [23913]));
Q_ASSIGN U8862 ( .B(clk), .A(\g.we_clk [23912]));
Q_ASSIGN U8863 ( .B(clk), .A(\g.we_clk [23911]));
Q_ASSIGN U8864 ( .B(clk), .A(\g.we_clk [23910]));
Q_ASSIGN U8865 ( .B(clk), .A(\g.we_clk [23909]));
Q_ASSIGN U8866 ( .B(clk), .A(\g.we_clk [23908]));
Q_ASSIGN U8867 ( .B(clk), .A(\g.we_clk [23907]));
Q_ASSIGN U8868 ( .B(clk), .A(\g.we_clk [23906]));
Q_ASSIGN U8869 ( .B(clk), .A(\g.we_clk [23905]));
Q_ASSIGN U8870 ( .B(clk), .A(\g.we_clk [23904]));
Q_ASSIGN U8871 ( .B(clk), .A(\g.we_clk [23903]));
Q_ASSIGN U8872 ( .B(clk), .A(\g.we_clk [23902]));
Q_ASSIGN U8873 ( .B(clk), .A(\g.we_clk [23901]));
Q_ASSIGN U8874 ( .B(clk), .A(\g.we_clk [23900]));
Q_ASSIGN U8875 ( .B(clk), .A(\g.we_clk [23899]));
Q_ASSIGN U8876 ( .B(clk), .A(\g.we_clk [23898]));
Q_ASSIGN U8877 ( .B(clk), .A(\g.we_clk [23897]));
Q_ASSIGN U8878 ( .B(clk), .A(\g.we_clk [23896]));
Q_ASSIGN U8879 ( .B(clk), .A(\g.we_clk [23895]));
Q_ASSIGN U8880 ( .B(clk), .A(\g.we_clk [23894]));
Q_ASSIGN U8881 ( .B(clk), .A(\g.we_clk [23893]));
Q_ASSIGN U8882 ( .B(clk), .A(\g.we_clk [23892]));
Q_ASSIGN U8883 ( .B(clk), .A(\g.we_clk [23891]));
Q_ASSIGN U8884 ( .B(clk), .A(\g.we_clk [23890]));
Q_ASSIGN U8885 ( .B(clk), .A(\g.we_clk [23889]));
Q_ASSIGN U8886 ( .B(clk), .A(\g.we_clk [23888]));
Q_ASSIGN U8887 ( .B(clk), .A(\g.we_clk [23887]));
Q_ASSIGN U8888 ( .B(clk), .A(\g.we_clk [23886]));
Q_ASSIGN U8889 ( .B(clk), .A(\g.we_clk [23885]));
Q_ASSIGN U8890 ( .B(clk), .A(\g.we_clk [23884]));
Q_ASSIGN U8891 ( .B(clk), .A(\g.we_clk [23883]));
Q_ASSIGN U8892 ( .B(clk), .A(\g.we_clk [23882]));
Q_ASSIGN U8893 ( .B(clk), .A(\g.we_clk [23881]));
Q_ASSIGN U8894 ( .B(clk), .A(\g.we_clk [23880]));
Q_ASSIGN U8895 ( .B(clk), .A(\g.we_clk [23879]));
Q_ASSIGN U8896 ( .B(clk), .A(\g.we_clk [23878]));
Q_ASSIGN U8897 ( .B(clk), .A(\g.we_clk [23877]));
Q_ASSIGN U8898 ( .B(clk), .A(\g.we_clk [23876]));
Q_ASSIGN U8899 ( .B(clk), .A(\g.we_clk [23875]));
Q_ASSIGN U8900 ( .B(clk), .A(\g.we_clk [23874]));
Q_ASSIGN U8901 ( .B(clk), .A(\g.we_clk [23873]));
Q_ASSIGN U8902 ( .B(clk), .A(\g.we_clk [23872]));
Q_ASSIGN U8903 ( .B(clk), .A(\g.we_clk [23871]));
Q_ASSIGN U8904 ( .B(clk), .A(\g.we_clk [23870]));
Q_ASSIGN U8905 ( .B(clk), .A(\g.we_clk [23869]));
Q_ASSIGN U8906 ( .B(clk), .A(\g.we_clk [23868]));
Q_ASSIGN U8907 ( .B(clk), .A(\g.we_clk [23867]));
Q_ASSIGN U8908 ( .B(clk), .A(\g.we_clk [23866]));
Q_ASSIGN U8909 ( .B(clk), .A(\g.we_clk [23865]));
Q_ASSIGN U8910 ( .B(clk), .A(\g.we_clk [23864]));
Q_ASSIGN U8911 ( .B(clk), .A(\g.we_clk [23863]));
Q_ASSIGN U8912 ( .B(clk), .A(\g.we_clk [23862]));
Q_ASSIGN U8913 ( .B(clk), .A(\g.we_clk [23861]));
Q_ASSIGN U8914 ( .B(clk), .A(\g.we_clk [23860]));
Q_ASSIGN U8915 ( .B(clk), .A(\g.we_clk [23859]));
Q_ASSIGN U8916 ( .B(clk), .A(\g.we_clk [23858]));
Q_ASSIGN U8917 ( .B(clk), .A(\g.we_clk [23857]));
Q_ASSIGN U8918 ( .B(clk), .A(\g.we_clk [23856]));
Q_ASSIGN U8919 ( .B(clk), .A(\g.we_clk [23855]));
Q_ASSIGN U8920 ( .B(clk), .A(\g.we_clk [23854]));
Q_ASSIGN U8921 ( .B(clk), .A(\g.we_clk [23853]));
Q_ASSIGN U8922 ( .B(clk), .A(\g.we_clk [23852]));
Q_ASSIGN U8923 ( .B(clk), .A(\g.we_clk [23851]));
Q_ASSIGN U8924 ( .B(clk), .A(\g.we_clk [23850]));
Q_ASSIGN U8925 ( .B(clk), .A(\g.we_clk [23849]));
Q_ASSIGN U8926 ( .B(clk), .A(\g.we_clk [23848]));
Q_ASSIGN U8927 ( .B(clk), .A(\g.we_clk [23847]));
Q_ASSIGN U8928 ( .B(clk), .A(\g.we_clk [23846]));
Q_ASSIGN U8929 ( .B(clk), .A(\g.we_clk [23845]));
Q_ASSIGN U8930 ( .B(clk), .A(\g.we_clk [23844]));
Q_ASSIGN U8931 ( .B(clk), .A(\g.we_clk [23843]));
Q_ASSIGN U8932 ( .B(clk), .A(\g.we_clk [23842]));
Q_ASSIGN U8933 ( .B(clk), .A(\g.we_clk [23841]));
Q_ASSIGN U8934 ( .B(clk), .A(\g.we_clk [23840]));
Q_ASSIGN U8935 ( .B(clk), .A(\g.we_clk [23839]));
Q_ASSIGN U8936 ( .B(clk), .A(\g.we_clk [23838]));
Q_ASSIGN U8937 ( .B(clk), .A(\g.we_clk [23837]));
Q_ASSIGN U8938 ( .B(clk), .A(\g.we_clk [23836]));
Q_ASSIGN U8939 ( .B(clk), .A(\g.we_clk [23835]));
Q_ASSIGN U8940 ( .B(clk), .A(\g.we_clk [23834]));
Q_ASSIGN U8941 ( .B(clk), .A(\g.we_clk [23833]));
Q_ASSIGN U8942 ( .B(clk), .A(\g.we_clk [23832]));
Q_ASSIGN U8943 ( .B(clk), .A(\g.we_clk [23831]));
Q_ASSIGN U8944 ( .B(clk), .A(\g.we_clk [23830]));
Q_ASSIGN U8945 ( .B(clk), .A(\g.we_clk [23829]));
Q_ASSIGN U8946 ( .B(clk), .A(\g.we_clk [23828]));
Q_ASSIGN U8947 ( .B(clk), .A(\g.we_clk [23827]));
Q_ASSIGN U8948 ( .B(clk), .A(\g.we_clk [23826]));
Q_ASSIGN U8949 ( .B(clk), .A(\g.we_clk [23825]));
Q_ASSIGN U8950 ( .B(clk), .A(\g.we_clk [23824]));
Q_ASSIGN U8951 ( .B(clk), .A(\g.we_clk [23823]));
Q_ASSIGN U8952 ( .B(clk), .A(\g.we_clk [23822]));
Q_ASSIGN U8953 ( .B(clk), .A(\g.we_clk [23821]));
Q_ASSIGN U8954 ( .B(clk), .A(\g.we_clk [23820]));
Q_ASSIGN U8955 ( .B(clk), .A(\g.we_clk [23819]));
Q_ASSIGN U8956 ( .B(clk), .A(\g.we_clk [23818]));
Q_ASSIGN U8957 ( .B(clk), .A(\g.we_clk [23817]));
Q_ASSIGN U8958 ( .B(clk), .A(\g.we_clk [23816]));
Q_ASSIGN U8959 ( .B(clk), .A(\g.we_clk [23815]));
Q_ASSIGN U8960 ( .B(clk), .A(\g.we_clk [23814]));
Q_ASSIGN U8961 ( .B(clk), .A(\g.we_clk [23813]));
Q_ASSIGN U8962 ( .B(clk), .A(\g.we_clk [23812]));
Q_ASSIGN U8963 ( .B(clk), .A(\g.we_clk [23811]));
Q_ASSIGN U8964 ( .B(clk), .A(\g.we_clk [23810]));
Q_ASSIGN U8965 ( .B(clk), .A(\g.we_clk [23809]));
Q_ASSIGN U8966 ( .B(clk), .A(\g.we_clk [23808]));
Q_ASSIGN U8967 ( .B(clk), .A(\g.we_clk [23807]));
Q_ASSIGN U8968 ( .B(clk), .A(\g.we_clk [23806]));
Q_ASSIGN U8969 ( .B(clk), .A(\g.we_clk [23805]));
Q_ASSIGN U8970 ( .B(clk), .A(\g.we_clk [23804]));
Q_ASSIGN U8971 ( .B(clk), .A(\g.we_clk [23803]));
Q_ASSIGN U8972 ( .B(clk), .A(\g.we_clk [23802]));
Q_ASSIGN U8973 ( .B(clk), .A(\g.we_clk [23801]));
Q_ASSIGN U8974 ( .B(clk), .A(\g.we_clk [23800]));
Q_ASSIGN U8975 ( .B(clk), .A(\g.we_clk [23799]));
Q_ASSIGN U8976 ( .B(clk), .A(\g.we_clk [23798]));
Q_ASSIGN U8977 ( .B(clk), .A(\g.we_clk [23797]));
Q_ASSIGN U8978 ( .B(clk), .A(\g.we_clk [23796]));
Q_ASSIGN U8979 ( .B(clk), .A(\g.we_clk [23795]));
Q_ASSIGN U8980 ( .B(clk), .A(\g.we_clk [23794]));
Q_ASSIGN U8981 ( .B(clk), .A(\g.we_clk [23793]));
Q_ASSIGN U8982 ( .B(clk), .A(\g.we_clk [23792]));
Q_ASSIGN U8983 ( .B(clk), .A(\g.we_clk [23791]));
Q_ASSIGN U8984 ( .B(clk), .A(\g.we_clk [23790]));
Q_ASSIGN U8985 ( .B(clk), .A(\g.we_clk [23789]));
Q_ASSIGN U8986 ( .B(clk), .A(\g.we_clk [23788]));
Q_ASSIGN U8987 ( .B(clk), .A(\g.we_clk [23787]));
Q_ASSIGN U8988 ( .B(clk), .A(\g.we_clk [23786]));
Q_ASSIGN U8989 ( .B(clk), .A(\g.we_clk [23785]));
Q_ASSIGN U8990 ( .B(clk), .A(\g.we_clk [23784]));
Q_ASSIGN U8991 ( .B(clk), .A(\g.we_clk [23783]));
Q_ASSIGN U8992 ( .B(clk), .A(\g.we_clk [23782]));
Q_ASSIGN U8993 ( .B(clk), .A(\g.we_clk [23781]));
Q_ASSIGN U8994 ( .B(clk), .A(\g.we_clk [23780]));
Q_ASSIGN U8995 ( .B(clk), .A(\g.we_clk [23779]));
Q_ASSIGN U8996 ( .B(clk), .A(\g.we_clk [23778]));
Q_ASSIGN U8997 ( .B(clk), .A(\g.we_clk [23777]));
Q_ASSIGN U8998 ( .B(clk), .A(\g.we_clk [23776]));
Q_ASSIGN U8999 ( .B(clk), .A(\g.we_clk [23775]));
Q_ASSIGN U9000 ( .B(clk), .A(\g.we_clk [23774]));
Q_ASSIGN U9001 ( .B(clk), .A(\g.we_clk [23773]));
Q_ASSIGN U9002 ( .B(clk), .A(\g.we_clk [23772]));
Q_ASSIGN U9003 ( .B(clk), .A(\g.we_clk [23771]));
Q_ASSIGN U9004 ( .B(clk), .A(\g.we_clk [23770]));
Q_ASSIGN U9005 ( .B(clk), .A(\g.we_clk [23769]));
Q_ASSIGN U9006 ( .B(clk), .A(\g.we_clk [23768]));
Q_ASSIGN U9007 ( .B(clk), .A(\g.we_clk [23767]));
Q_ASSIGN U9008 ( .B(clk), .A(\g.we_clk [23766]));
Q_ASSIGN U9009 ( .B(clk), .A(\g.we_clk [23765]));
Q_ASSIGN U9010 ( .B(clk), .A(\g.we_clk [23764]));
Q_ASSIGN U9011 ( .B(clk), .A(\g.we_clk [23763]));
Q_ASSIGN U9012 ( .B(clk), .A(\g.we_clk [23762]));
Q_ASSIGN U9013 ( .B(clk), .A(\g.we_clk [23761]));
Q_ASSIGN U9014 ( .B(clk), .A(\g.we_clk [23760]));
Q_ASSIGN U9015 ( .B(clk), .A(\g.we_clk [23759]));
Q_ASSIGN U9016 ( .B(clk), .A(\g.we_clk [23758]));
Q_ASSIGN U9017 ( .B(clk), .A(\g.we_clk [23757]));
Q_ASSIGN U9018 ( .B(clk), .A(\g.we_clk [23756]));
Q_ASSIGN U9019 ( .B(clk), .A(\g.we_clk [23755]));
Q_ASSIGN U9020 ( .B(clk), .A(\g.we_clk [23754]));
Q_ASSIGN U9021 ( .B(clk), .A(\g.we_clk [23753]));
Q_ASSIGN U9022 ( .B(clk), .A(\g.we_clk [23752]));
Q_ASSIGN U9023 ( .B(clk), .A(\g.we_clk [23751]));
Q_ASSIGN U9024 ( .B(clk), .A(\g.we_clk [23750]));
Q_ASSIGN U9025 ( .B(clk), .A(\g.we_clk [23749]));
Q_ASSIGN U9026 ( .B(clk), .A(\g.we_clk [23748]));
Q_ASSIGN U9027 ( .B(clk), .A(\g.we_clk [23747]));
Q_ASSIGN U9028 ( .B(clk), .A(\g.we_clk [23746]));
Q_ASSIGN U9029 ( .B(clk), .A(\g.we_clk [23745]));
Q_ASSIGN U9030 ( .B(clk), .A(\g.we_clk [23744]));
Q_ASSIGN U9031 ( .B(clk), .A(\g.we_clk [23743]));
Q_ASSIGN U9032 ( .B(clk), .A(\g.we_clk [23742]));
Q_ASSIGN U9033 ( .B(clk), .A(\g.we_clk [23741]));
Q_ASSIGN U9034 ( .B(clk), .A(\g.we_clk [23740]));
Q_ASSIGN U9035 ( .B(clk), .A(\g.we_clk [23739]));
Q_ASSIGN U9036 ( .B(clk), .A(\g.we_clk [23738]));
Q_ASSIGN U9037 ( .B(clk), .A(\g.we_clk [23737]));
Q_ASSIGN U9038 ( .B(clk), .A(\g.we_clk [23736]));
Q_ASSIGN U9039 ( .B(clk), .A(\g.we_clk [23735]));
Q_ASSIGN U9040 ( .B(clk), .A(\g.we_clk [23734]));
Q_ASSIGN U9041 ( .B(clk), .A(\g.we_clk [23733]));
Q_ASSIGN U9042 ( .B(clk), .A(\g.we_clk [23732]));
Q_ASSIGN U9043 ( .B(clk), .A(\g.we_clk [23731]));
Q_ASSIGN U9044 ( .B(clk), .A(\g.we_clk [23730]));
Q_ASSIGN U9045 ( .B(clk), .A(\g.we_clk [23729]));
Q_ASSIGN U9046 ( .B(clk), .A(\g.we_clk [23728]));
Q_ASSIGN U9047 ( .B(clk), .A(\g.we_clk [23727]));
Q_ASSIGN U9048 ( .B(clk), .A(\g.we_clk [23726]));
Q_ASSIGN U9049 ( .B(clk), .A(\g.we_clk [23725]));
Q_ASSIGN U9050 ( .B(clk), .A(\g.we_clk [23724]));
Q_ASSIGN U9051 ( .B(clk), .A(\g.we_clk [23723]));
Q_ASSIGN U9052 ( .B(clk), .A(\g.we_clk [23722]));
Q_ASSIGN U9053 ( .B(clk), .A(\g.we_clk [23721]));
Q_ASSIGN U9054 ( .B(clk), .A(\g.we_clk [23720]));
Q_ASSIGN U9055 ( .B(clk), .A(\g.we_clk [23719]));
Q_ASSIGN U9056 ( .B(clk), .A(\g.we_clk [23718]));
Q_ASSIGN U9057 ( .B(clk), .A(\g.we_clk [23717]));
Q_ASSIGN U9058 ( .B(clk), .A(\g.we_clk [23716]));
Q_ASSIGN U9059 ( .B(clk), .A(\g.we_clk [23715]));
Q_ASSIGN U9060 ( .B(clk), .A(\g.we_clk [23714]));
Q_ASSIGN U9061 ( .B(clk), .A(\g.we_clk [23713]));
Q_ASSIGN U9062 ( .B(clk), .A(\g.we_clk [23712]));
Q_ASSIGN U9063 ( .B(clk), .A(\g.we_clk [23711]));
Q_ASSIGN U9064 ( .B(clk), .A(\g.we_clk [23710]));
Q_ASSIGN U9065 ( .B(clk), .A(\g.we_clk [23709]));
Q_ASSIGN U9066 ( .B(clk), .A(\g.we_clk [23708]));
Q_ASSIGN U9067 ( .B(clk), .A(\g.we_clk [23707]));
Q_ASSIGN U9068 ( .B(clk), .A(\g.we_clk [23706]));
Q_ASSIGN U9069 ( .B(clk), .A(\g.we_clk [23705]));
Q_ASSIGN U9070 ( .B(clk), .A(\g.we_clk [23704]));
Q_ASSIGN U9071 ( .B(clk), .A(\g.we_clk [23703]));
Q_ASSIGN U9072 ( .B(clk), .A(\g.we_clk [23702]));
Q_ASSIGN U9073 ( .B(clk), .A(\g.we_clk [23701]));
Q_ASSIGN U9074 ( .B(clk), .A(\g.we_clk [23700]));
Q_ASSIGN U9075 ( .B(clk), .A(\g.we_clk [23699]));
Q_ASSIGN U9076 ( .B(clk), .A(\g.we_clk [23698]));
Q_ASSIGN U9077 ( .B(clk), .A(\g.we_clk [23697]));
Q_ASSIGN U9078 ( .B(clk), .A(\g.we_clk [23696]));
Q_ASSIGN U9079 ( .B(clk), .A(\g.we_clk [23695]));
Q_ASSIGN U9080 ( .B(clk), .A(\g.we_clk [23694]));
Q_ASSIGN U9081 ( .B(clk), .A(\g.we_clk [23693]));
Q_ASSIGN U9082 ( .B(clk), .A(\g.we_clk [23692]));
Q_ASSIGN U9083 ( .B(clk), .A(\g.we_clk [23691]));
Q_ASSIGN U9084 ( .B(clk), .A(\g.we_clk [23690]));
Q_ASSIGN U9085 ( .B(clk), .A(\g.we_clk [23689]));
Q_ASSIGN U9086 ( .B(clk), .A(\g.we_clk [23688]));
Q_ASSIGN U9087 ( .B(clk), .A(\g.we_clk [23687]));
Q_ASSIGN U9088 ( .B(clk), .A(\g.we_clk [23686]));
Q_ASSIGN U9089 ( .B(clk), .A(\g.we_clk [23685]));
Q_ASSIGN U9090 ( .B(clk), .A(\g.we_clk [23684]));
Q_ASSIGN U9091 ( .B(clk), .A(\g.we_clk [23683]));
Q_ASSIGN U9092 ( .B(clk), .A(\g.we_clk [23682]));
Q_ASSIGN U9093 ( .B(clk), .A(\g.we_clk [23681]));
Q_ASSIGN U9094 ( .B(clk), .A(\g.we_clk [23680]));
Q_ASSIGN U9095 ( .B(clk), .A(\g.we_clk [23679]));
Q_ASSIGN U9096 ( .B(clk), .A(\g.we_clk [23678]));
Q_ASSIGN U9097 ( .B(clk), .A(\g.we_clk [23677]));
Q_ASSIGN U9098 ( .B(clk), .A(\g.we_clk [23676]));
Q_ASSIGN U9099 ( .B(clk), .A(\g.we_clk [23675]));
Q_ASSIGN U9100 ( .B(clk), .A(\g.we_clk [23674]));
Q_ASSIGN U9101 ( .B(clk), .A(\g.we_clk [23673]));
Q_ASSIGN U9102 ( .B(clk), .A(\g.we_clk [23672]));
Q_ASSIGN U9103 ( .B(clk), .A(\g.we_clk [23671]));
Q_ASSIGN U9104 ( .B(clk), .A(\g.we_clk [23670]));
Q_ASSIGN U9105 ( .B(clk), .A(\g.we_clk [23669]));
Q_ASSIGN U9106 ( .B(clk), .A(\g.we_clk [23668]));
Q_ASSIGN U9107 ( .B(clk), .A(\g.we_clk [23667]));
Q_ASSIGN U9108 ( .B(clk), .A(\g.we_clk [23666]));
Q_ASSIGN U9109 ( .B(clk), .A(\g.we_clk [23665]));
Q_ASSIGN U9110 ( .B(clk), .A(\g.we_clk [23664]));
Q_ASSIGN U9111 ( .B(clk), .A(\g.we_clk [23663]));
Q_ASSIGN U9112 ( .B(clk), .A(\g.we_clk [23662]));
Q_ASSIGN U9113 ( .B(clk), .A(\g.we_clk [23661]));
Q_ASSIGN U9114 ( .B(clk), .A(\g.we_clk [23660]));
Q_ASSIGN U9115 ( .B(clk), .A(\g.we_clk [23659]));
Q_ASSIGN U9116 ( .B(clk), .A(\g.we_clk [23658]));
Q_ASSIGN U9117 ( .B(clk), .A(\g.we_clk [23657]));
Q_ASSIGN U9118 ( .B(clk), .A(\g.we_clk [23656]));
Q_ASSIGN U9119 ( .B(clk), .A(\g.we_clk [23655]));
Q_ASSIGN U9120 ( .B(clk), .A(\g.we_clk [23654]));
Q_ASSIGN U9121 ( .B(clk), .A(\g.we_clk [23653]));
Q_ASSIGN U9122 ( .B(clk), .A(\g.we_clk [23652]));
Q_ASSIGN U9123 ( .B(clk), .A(\g.we_clk [23651]));
Q_ASSIGN U9124 ( .B(clk), .A(\g.we_clk [23650]));
Q_ASSIGN U9125 ( .B(clk), .A(\g.we_clk [23649]));
Q_ASSIGN U9126 ( .B(clk), .A(\g.we_clk [23648]));
Q_ASSIGN U9127 ( .B(clk), .A(\g.we_clk [23647]));
Q_ASSIGN U9128 ( .B(clk), .A(\g.we_clk [23646]));
Q_ASSIGN U9129 ( .B(clk), .A(\g.we_clk [23645]));
Q_ASSIGN U9130 ( .B(clk), .A(\g.we_clk [23644]));
Q_ASSIGN U9131 ( .B(clk), .A(\g.we_clk [23643]));
Q_ASSIGN U9132 ( .B(clk), .A(\g.we_clk [23642]));
Q_ASSIGN U9133 ( .B(clk), .A(\g.we_clk [23641]));
Q_ASSIGN U9134 ( .B(clk), .A(\g.we_clk [23640]));
Q_ASSIGN U9135 ( .B(clk), .A(\g.we_clk [23639]));
Q_ASSIGN U9136 ( .B(clk), .A(\g.we_clk [23638]));
Q_ASSIGN U9137 ( .B(clk), .A(\g.we_clk [23637]));
Q_ASSIGN U9138 ( .B(clk), .A(\g.we_clk [23636]));
Q_ASSIGN U9139 ( .B(clk), .A(\g.we_clk [23635]));
Q_ASSIGN U9140 ( .B(clk), .A(\g.we_clk [23634]));
Q_ASSIGN U9141 ( .B(clk), .A(\g.we_clk [23633]));
Q_ASSIGN U9142 ( .B(clk), .A(\g.we_clk [23632]));
Q_ASSIGN U9143 ( .B(clk), .A(\g.we_clk [23631]));
Q_ASSIGN U9144 ( .B(clk), .A(\g.we_clk [23630]));
Q_ASSIGN U9145 ( .B(clk), .A(\g.we_clk [23629]));
Q_ASSIGN U9146 ( .B(clk), .A(\g.we_clk [23628]));
Q_ASSIGN U9147 ( .B(clk), .A(\g.we_clk [23627]));
Q_ASSIGN U9148 ( .B(clk), .A(\g.we_clk [23626]));
Q_ASSIGN U9149 ( .B(clk), .A(\g.we_clk [23625]));
Q_ASSIGN U9150 ( .B(clk), .A(\g.we_clk [23624]));
Q_ASSIGN U9151 ( .B(clk), .A(\g.we_clk [23623]));
Q_ASSIGN U9152 ( .B(clk), .A(\g.we_clk [23622]));
Q_ASSIGN U9153 ( .B(clk), .A(\g.we_clk [23621]));
Q_ASSIGN U9154 ( .B(clk), .A(\g.we_clk [23620]));
Q_ASSIGN U9155 ( .B(clk), .A(\g.we_clk [23619]));
Q_ASSIGN U9156 ( .B(clk), .A(\g.we_clk [23618]));
Q_ASSIGN U9157 ( .B(clk), .A(\g.we_clk [23617]));
Q_ASSIGN U9158 ( .B(clk), .A(\g.we_clk [23616]));
Q_ASSIGN U9159 ( .B(clk), .A(\g.we_clk [23615]));
Q_ASSIGN U9160 ( .B(clk), .A(\g.we_clk [23614]));
Q_ASSIGN U9161 ( .B(clk), .A(\g.we_clk [23613]));
Q_ASSIGN U9162 ( .B(clk), .A(\g.we_clk [23612]));
Q_ASSIGN U9163 ( .B(clk), .A(\g.we_clk [23611]));
Q_ASSIGN U9164 ( .B(clk), .A(\g.we_clk [23610]));
Q_ASSIGN U9165 ( .B(clk), .A(\g.we_clk [23609]));
Q_ASSIGN U9166 ( .B(clk), .A(\g.we_clk [23608]));
Q_ASSIGN U9167 ( .B(clk), .A(\g.we_clk [23607]));
Q_ASSIGN U9168 ( .B(clk), .A(\g.we_clk [23606]));
Q_ASSIGN U9169 ( .B(clk), .A(\g.we_clk [23605]));
Q_ASSIGN U9170 ( .B(clk), .A(\g.we_clk [23604]));
Q_ASSIGN U9171 ( .B(clk), .A(\g.we_clk [23603]));
Q_ASSIGN U9172 ( .B(clk), .A(\g.we_clk [23602]));
Q_ASSIGN U9173 ( .B(clk), .A(\g.we_clk [23601]));
Q_ASSIGN U9174 ( .B(clk), .A(\g.we_clk [23600]));
Q_ASSIGN U9175 ( .B(clk), .A(\g.we_clk [23599]));
Q_ASSIGN U9176 ( .B(clk), .A(\g.we_clk [23598]));
Q_ASSIGN U9177 ( .B(clk), .A(\g.we_clk [23597]));
Q_ASSIGN U9178 ( .B(clk), .A(\g.we_clk [23596]));
Q_ASSIGN U9179 ( .B(clk), .A(\g.we_clk [23595]));
Q_ASSIGN U9180 ( .B(clk), .A(\g.we_clk [23594]));
Q_ASSIGN U9181 ( .B(clk), .A(\g.we_clk [23593]));
Q_ASSIGN U9182 ( .B(clk), .A(\g.we_clk [23592]));
Q_ASSIGN U9183 ( .B(clk), .A(\g.we_clk [23591]));
Q_ASSIGN U9184 ( .B(clk), .A(\g.we_clk [23590]));
Q_ASSIGN U9185 ( .B(clk), .A(\g.we_clk [23589]));
Q_ASSIGN U9186 ( .B(clk), .A(\g.we_clk [23588]));
Q_ASSIGN U9187 ( .B(clk), .A(\g.we_clk [23587]));
Q_ASSIGN U9188 ( .B(clk), .A(\g.we_clk [23586]));
Q_ASSIGN U9189 ( .B(clk), .A(\g.we_clk [23585]));
Q_ASSIGN U9190 ( .B(clk), .A(\g.we_clk [23584]));
Q_ASSIGN U9191 ( .B(clk), .A(\g.we_clk [23583]));
Q_ASSIGN U9192 ( .B(clk), .A(\g.we_clk [23582]));
Q_ASSIGN U9193 ( .B(clk), .A(\g.we_clk [23581]));
Q_ASSIGN U9194 ( .B(clk), .A(\g.we_clk [23580]));
Q_ASSIGN U9195 ( .B(clk), .A(\g.we_clk [23579]));
Q_ASSIGN U9196 ( .B(clk), .A(\g.we_clk [23578]));
Q_ASSIGN U9197 ( .B(clk), .A(\g.we_clk [23577]));
Q_ASSIGN U9198 ( .B(clk), .A(\g.we_clk [23576]));
Q_ASSIGN U9199 ( .B(clk), .A(\g.we_clk [23575]));
Q_ASSIGN U9200 ( .B(clk), .A(\g.we_clk [23574]));
Q_ASSIGN U9201 ( .B(clk), .A(\g.we_clk [23573]));
Q_ASSIGN U9202 ( .B(clk), .A(\g.we_clk [23572]));
Q_ASSIGN U9203 ( .B(clk), .A(\g.we_clk [23571]));
Q_ASSIGN U9204 ( .B(clk), .A(\g.we_clk [23570]));
Q_ASSIGN U9205 ( .B(clk), .A(\g.we_clk [23569]));
Q_ASSIGN U9206 ( .B(clk), .A(\g.we_clk [23568]));
Q_ASSIGN U9207 ( .B(clk), .A(\g.we_clk [23567]));
Q_ASSIGN U9208 ( .B(clk), .A(\g.we_clk [23566]));
Q_ASSIGN U9209 ( .B(clk), .A(\g.we_clk [23565]));
Q_ASSIGN U9210 ( .B(clk), .A(\g.we_clk [23564]));
Q_ASSIGN U9211 ( .B(clk), .A(\g.we_clk [23563]));
Q_ASSIGN U9212 ( .B(clk), .A(\g.we_clk [23562]));
Q_ASSIGN U9213 ( .B(clk), .A(\g.we_clk [23561]));
Q_ASSIGN U9214 ( .B(clk), .A(\g.we_clk [23560]));
Q_ASSIGN U9215 ( .B(clk), .A(\g.we_clk [23559]));
Q_ASSIGN U9216 ( .B(clk), .A(\g.we_clk [23558]));
Q_ASSIGN U9217 ( .B(clk), .A(\g.we_clk [23557]));
Q_ASSIGN U9218 ( .B(clk), .A(\g.we_clk [23556]));
Q_ASSIGN U9219 ( .B(clk), .A(\g.we_clk [23555]));
Q_ASSIGN U9220 ( .B(clk), .A(\g.we_clk [23554]));
Q_ASSIGN U9221 ( .B(clk), .A(\g.we_clk [23553]));
Q_ASSIGN U9222 ( .B(clk), .A(\g.we_clk [23552]));
Q_ASSIGN U9223 ( .B(clk), .A(\g.we_clk [23551]));
Q_ASSIGN U9224 ( .B(clk), .A(\g.we_clk [23550]));
Q_ASSIGN U9225 ( .B(clk), .A(\g.we_clk [23549]));
Q_ASSIGN U9226 ( .B(clk), .A(\g.we_clk [23548]));
Q_ASSIGN U9227 ( .B(clk), .A(\g.we_clk [23547]));
Q_ASSIGN U9228 ( .B(clk), .A(\g.we_clk [23546]));
Q_ASSIGN U9229 ( .B(clk), .A(\g.we_clk [23545]));
Q_ASSIGN U9230 ( .B(clk), .A(\g.we_clk [23544]));
Q_ASSIGN U9231 ( .B(clk), .A(\g.we_clk [23543]));
Q_ASSIGN U9232 ( .B(clk), .A(\g.we_clk [23542]));
Q_ASSIGN U9233 ( .B(clk), .A(\g.we_clk [23541]));
Q_ASSIGN U9234 ( .B(clk), .A(\g.we_clk [23540]));
Q_ASSIGN U9235 ( .B(clk), .A(\g.we_clk [23539]));
Q_ASSIGN U9236 ( .B(clk), .A(\g.we_clk [23538]));
Q_ASSIGN U9237 ( .B(clk), .A(\g.we_clk [23537]));
Q_ASSIGN U9238 ( .B(clk), .A(\g.we_clk [23536]));
Q_ASSIGN U9239 ( .B(clk), .A(\g.we_clk [23535]));
Q_ASSIGN U9240 ( .B(clk), .A(\g.we_clk [23534]));
Q_ASSIGN U9241 ( .B(clk), .A(\g.we_clk [23533]));
Q_ASSIGN U9242 ( .B(clk), .A(\g.we_clk [23532]));
Q_ASSIGN U9243 ( .B(clk), .A(\g.we_clk [23531]));
Q_ASSIGN U9244 ( .B(clk), .A(\g.we_clk [23530]));
Q_ASSIGN U9245 ( .B(clk), .A(\g.we_clk [23529]));
Q_ASSIGN U9246 ( .B(clk), .A(\g.we_clk [23528]));
Q_ASSIGN U9247 ( .B(clk), .A(\g.we_clk [23527]));
Q_ASSIGN U9248 ( .B(clk), .A(\g.we_clk [23526]));
Q_ASSIGN U9249 ( .B(clk), .A(\g.we_clk [23525]));
Q_ASSIGN U9250 ( .B(clk), .A(\g.we_clk [23524]));
Q_ASSIGN U9251 ( .B(clk), .A(\g.we_clk [23523]));
Q_ASSIGN U9252 ( .B(clk), .A(\g.we_clk [23522]));
Q_ASSIGN U9253 ( .B(clk), .A(\g.we_clk [23521]));
Q_ASSIGN U9254 ( .B(clk), .A(\g.we_clk [23520]));
Q_ASSIGN U9255 ( .B(clk), .A(\g.we_clk [23519]));
Q_ASSIGN U9256 ( .B(clk), .A(\g.we_clk [23518]));
Q_ASSIGN U9257 ( .B(clk), .A(\g.we_clk [23517]));
Q_ASSIGN U9258 ( .B(clk), .A(\g.we_clk [23516]));
Q_ASSIGN U9259 ( .B(clk), .A(\g.we_clk [23515]));
Q_ASSIGN U9260 ( .B(clk), .A(\g.we_clk [23514]));
Q_ASSIGN U9261 ( .B(clk), .A(\g.we_clk [23513]));
Q_ASSIGN U9262 ( .B(clk), .A(\g.we_clk [23512]));
Q_ASSIGN U9263 ( .B(clk), .A(\g.we_clk [23511]));
Q_ASSIGN U9264 ( .B(clk), .A(\g.we_clk [23510]));
Q_ASSIGN U9265 ( .B(clk), .A(\g.we_clk [23509]));
Q_ASSIGN U9266 ( .B(clk), .A(\g.we_clk [23508]));
Q_ASSIGN U9267 ( .B(clk), .A(\g.we_clk [23507]));
Q_ASSIGN U9268 ( .B(clk), .A(\g.we_clk [23506]));
Q_ASSIGN U9269 ( .B(clk), .A(\g.we_clk [23505]));
Q_ASSIGN U9270 ( .B(clk), .A(\g.we_clk [23504]));
Q_ASSIGN U9271 ( .B(clk), .A(\g.we_clk [23503]));
Q_ASSIGN U9272 ( .B(clk), .A(\g.we_clk [23502]));
Q_ASSIGN U9273 ( .B(clk), .A(\g.we_clk [23501]));
Q_ASSIGN U9274 ( .B(clk), .A(\g.we_clk [23500]));
Q_ASSIGN U9275 ( .B(clk), .A(\g.we_clk [23499]));
Q_ASSIGN U9276 ( .B(clk), .A(\g.we_clk [23498]));
Q_ASSIGN U9277 ( .B(clk), .A(\g.we_clk [23497]));
Q_ASSIGN U9278 ( .B(clk), .A(\g.we_clk [23496]));
Q_ASSIGN U9279 ( .B(clk), .A(\g.we_clk [23495]));
Q_ASSIGN U9280 ( .B(clk), .A(\g.we_clk [23494]));
Q_ASSIGN U9281 ( .B(clk), .A(\g.we_clk [23493]));
Q_ASSIGN U9282 ( .B(clk), .A(\g.we_clk [23492]));
Q_ASSIGN U9283 ( .B(clk), .A(\g.we_clk [23491]));
Q_ASSIGN U9284 ( .B(clk), .A(\g.we_clk [23490]));
Q_ASSIGN U9285 ( .B(clk), .A(\g.we_clk [23489]));
Q_ASSIGN U9286 ( .B(clk), .A(\g.we_clk [23488]));
Q_ASSIGN U9287 ( .B(clk), .A(\g.we_clk [23487]));
Q_ASSIGN U9288 ( .B(clk), .A(\g.we_clk [23486]));
Q_ASSIGN U9289 ( .B(clk), .A(\g.we_clk [23485]));
Q_ASSIGN U9290 ( .B(clk), .A(\g.we_clk [23484]));
Q_ASSIGN U9291 ( .B(clk), .A(\g.we_clk [23483]));
Q_ASSIGN U9292 ( .B(clk), .A(\g.we_clk [23482]));
Q_ASSIGN U9293 ( .B(clk), .A(\g.we_clk [23481]));
Q_ASSIGN U9294 ( .B(clk), .A(\g.we_clk [23480]));
Q_ASSIGN U9295 ( .B(clk), .A(\g.we_clk [23479]));
Q_ASSIGN U9296 ( .B(clk), .A(\g.we_clk [23478]));
Q_ASSIGN U9297 ( .B(clk), .A(\g.we_clk [23477]));
Q_ASSIGN U9298 ( .B(clk), .A(\g.we_clk [23476]));
Q_ASSIGN U9299 ( .B(clk), .A(\g.we_clk [23475]));
Q_ASSIGN U9300 ( .B(clk), .A(\g.we_clk [23474]));
Q_ASSIGN U9301 ( .B(clk), .A(\g.we_clk [23473]));
Q_ASSIGN U9302 ( .B(clk), .A(\g.we_clk [23472]));
Q_ASSIGN U9303 ( .B(clk), .A(\g.we_clk [23471]));
Q_ASSIGN U9304 ( .B(clk), .A(\g.we_clk [23470]));
Q_ASSIGN U9305 ( .B(clk), .A(\g.we_clk [23469]));
Q_ASSIGN U9306 ( .B(clk), .A(\g.we_clk [23468]));
Q_ASSIGN U9307 ( .B(clk), .A(\g.we_clk [23467]));
Q_ASSIGN U9308 ( .B(clk), .A(\g.we_clk [23466]));
Q_ASSIGN U9309 ( .B(clk), .A(\g.we_clk [23465]));
Q_ASSIGN U9310 ( .B(clk), .A(\g.we_clk [23464]));
Q_ASSIGN U9311 ( .B(clk), .A(\g.we_clk [23463]));
Q_ASSIGN U9312 ( .B(clk), .A(\g.we_clk [23462]));
Q_ASSIGN U9313 ( .B(clk), .A(\g.we_clk [23461]));
Q_ASSIGN U9314 ( .B(clk), .A(\g.we_clk [23460]));
Q_ASSIGN U9315 ( .B(clk), .A(\g.we_clk [23459]));
Q_ASSIGN U9316 ( .B(clk), .A(\g.we_clk [23458]));
Q_ASSIGN U9317 ( .B(clk), .A(\g.we_clk [23457]));
Q_ASSIGN U9318 ( .B(clk), .A(\g.we_clk [23456]));
Q_ASSIGN U9319 ( .B(clk), .A(\g.we_clk [23455]));
Q_ASSIGN U9320 ( .B(clk), .A(\g.we_clk [23454]));
Q_ASSIGN U9321 ( .B(clk), .A(\g.we_clk [23453]));
Q_ASSIGN U9322 ( .B(clk), .A(\g.we_clk [23452]));
Q_ASSIGN U9323 ( .B(clk), .A(\g.we_clk [23451]));
Q_ASSIGN U9324 ( .B(clk), .A(\g.we_clk [23450]));
Q_ASSIGN U9325 ( .B(clk), .A(\g.we_clk [23449]));
Q_ASSIGN U9326 ( .B(clk), .A(\g.we_clk [23448]));
Q_ASSIGN U9327 ( .B(clk), .A(\g.we_clk [23447]));
Q_ASSIGN U9328 ( .B(clk), .A(\g.we_clk [23446]));
Q_ASSIGN U9329 ( .B(clk), .A(\g.we_clk [23445]));
Q_ASSIGN U9330 ( .B(clk), .A(\g.we_clk [23444]));
Q_ASSIGN U9331 ( .B(clk), .A(\g.we_clk [23443]));
Q_ASSIGN U9332 ( .B(clk), .A(\g.we_clk [23442]));
Q_ASSIGN U9333 ( .B(clk), .A(\g.we_clk [23441]));
Q_ASSIGN U9334 ( .B(clk), .A(\g.we_clk [23440]));
Q_ASSIGN U9335 ( .B(clk), .A(\g.we_clk [23439]));
Q_ASSIGN U9336 ( .B(clk), .A(\g.we_clk [23438]));
Q_ASSIGN U9337 ( .B(clk), .A(\g.we_clk [23437]));
Q_ASSIGN U9338 ( .B(clk), .A(\g.we_clk [23436]));
Q_ASSIGN U9339 ( .B(clk), .A(\g.we_clk [23435]));
Q_ASSIGN U9340 ( .B(clk), .A(\g.we_clk [23434]));
Q_ASSIGN U9341 ( .B(clk), .A(\g.we_clk [23433]));
Q_ASSIGN U9342 ( .B(clk), .A(\g.we_clk [23432]));
Q_ASSIGN U9343 ( .B(clk), .A(\g.we_clk [23431]));
Q_ASSIGN U9344 ( .B(clk), .A(\g.we_clk [23430]));
Q_ASSIGN U9345 ( .B(clk), .A(\g.we_clk [23429]));
Q_ASSIGN U9346 ( .B(clk), .A(\g.we_clk [23428]));
Q_ASSIGN U9347 ( .B(clk), .A(\g.we_clk [23427]));
Q_ASSIGN U9348 ( .B(clk), .A(\g.we_clk [23426]));
Q_ASSIGN U9349 ( .B(clk), .A(\g.we_clk [23425]));
Q_ASSIGN U9350 ( .B(clk), .A(\g.we_clk [23424]));
Q_ASSIGN U9351 ( .B(clk), .A(\g.we_clk [23423]));
Q_ASSIGN U9352 ( .B(clk), .A(\g.we_clk [23422]));
Q_ASSIGN U9353 ( .B(clk), .A(\g.we_clk [23421]));
Q_ASSIGN U9354 ( .B(clk), .A(\g.we_clk [23420]));
Q_ASSIGN U9355 ( .B(clk), .A(\g.we_clk [23419]));
Q_ASSIGN U9356 ( .B(clk), .A(\g.we_clk [23418]));
Q_ASSIGN U9357 ( .B(clk), .A(\g.we_clk [23417]));
Q_ASSIGN U9358 ( .B(clk), .A(\g.we_clk [23416]));
Q_ASSIGN U9359 ( .B(clk), .A(\g.we_clk [23415]));
Q_ASSIGN U9360 ( .B(clk), .A(\g.we_clk [23414]));
Q_ASSIGN U9361 ( .B(clk), .A(\g.we_clk [23413]));
Q_ASSIGN U9362 ( .B(clk), .A(\g.we_clk [23412]));
Q_ASSIGN U9363 ( .B(clk), .A(\g.we_clk [23411]));
Q_ASSIGN U9364 ( .B(clk), .A(\g.we_clk [23410]));
Q_ASSIGN U9365 ( .B(clk), .A(\g.we_clk [23409]));
Q_ASSIGN U9366 ( .B(clk), .A(\g.we_clk [23408]));
Q_ASSIGN U9367 ( .B(clk), .A(\g.we_clk [23407]));
Q_ASSIGN U9368 ( .B(clk), .A(\g.we_clk [23406]));
Q_ASSIGN U9369 ( .B(clk), .A(\g.we_clk [23405]));
Q_ASSIGN U9370 ( .B(clk), .A(\g.we_clk [23404]));
Q_ASSIGN U9371 ( .B(clk), .A(\g.we_clk [23403]));
Q_ASSIGN U9372 ( .B(clk), .A(\g.we_clk [23402]));
Q_ASSIGN U9373 ( .B(clk), .A(\g.we_clk [23401]));
Q_ASSIGN U9374 ( .B(clk), .A(\g.we_clk [23400]));
Q_ASSIGN U9375 ( .B(clk), .A(\g.we_clk [23399]));
Q_ASSIGN U9376 ( .B(clk), .A(\g.we_clk [23398]));
Q_ASSIGN U9377 ( .B(clk), .A(\g.we_clk [23397]));
Q_ASSIGN U9378 ( .B(clk), .A(\g.we_clk [23396]));
Q_ASSIGN U9379 ( .B(clk), .A(\g.we_clk [23395]));
Q_ASSIGN U9380 ( .B(clk), .A(\g.we_clk [23394]));
Q_ASSIGN U9381 ( .B(clk), .A(\g.we_clk [23393]));
Q_ASSIGN U9382 ( .B(clk), .A(\g.we_clk [23392]));
Q_ASSIGN U9383 ( .B(clk), .A(\g.we_clk [23391]));
Q_ASSIGN U9384 ( .B(clk), .A(\g.we_clk [23390]));
Q_ASSIGN U9385 ( .B(clk), .A(\g.we_clk [23389]));
Q_ASSIGN U9386 ( .B(clk), .A(\g.we_clk [23388]));
Q_ASSIGN U9387 ( .B(clk), .A(\g.we_clk [23387]));
Q_ASSIGN U9388 ( .B(clk), .A(\g.we_clk [23386]));
Q_ASSIGN U9389 ( .B(clk), .A(\g.we_clk [23385]));
Q_ASSIGN U9390 ( .B(clk), .A(\g.we_clk [23384]));
Q_ASSIGN U9391 ( .B(clk), .A(\g.we_clk [23383]));
Q_ASSIGN U9392 ( .B(clk), .A(\g.we_clk [23382]));
Q_ASSIGN U9393 ( .B(clk), .A(\g.we_clk [23381]));
Q_ASSIGN U9394 ( .B(clk), .A(\g.we_clk [23380]));
Q_ASSIGN U9395 ( .B(clk), .A(\g.we_clk [23379]));
Q_ASSIGN U9396 ( .B(clk), .A(\g.we_clk [23378]));
Q_ASSIGN U9397 ( .B(clk), .A(\g.we_clk [23377]));
Q_ASSIGN U9398 ( .B(clk), .A(\g.we_clk [23376]));
Q_ASSIGN U9399 ( .B(clk), .A(\g.we_clk [23375]));
Q_ASSIGN U9400 ( .B(clk), .A(\g.we_clk [23374]));
Q_ASSIGN U9401 ( .B(clk), .A(\g.we_clk [23373]));
Q_ASSIGN U9402 ( .B(clk), .A(\g.we_clk [23372]));
Q_ASSIGN U9403 ( .B(clk), .A(\g.we_clk [23371]));
Q_ASSIGN U9404 ( .B(clk), .A(\g.we_clk [23370]));
Q_ASSIGN U9405 ( .B(clk), .A(\g.we_clk [23369]));
Q_ASSIGN U9406 ( .B(clk), .A(\g.we_clk [23368]));
Q_ASSIGN U9407 ( .B(clk), .A(\g.we_clk [23367]));
Q_ASSIGN U9408 ( .B(clk), .A(\g.we_clk [23366]));
Q_ASSIGN U9409 ( .B(clk), .A(\g.we_clk [23365]));
Q_ASSIGN U9410 ( .B(clk), .A(\g.we_clk [23364]));
Q_ASSIGN U9411 ( .B(clk), .A(\g.we_clk [23363]));
Q_ASSIGN U9412 ( .B(clk), .A(\g.we_clk [23362]));
Q_ASSIGN U9413 ( .B(clk), .A(\g.we_clk [23361]));
Q_ASSIGN U9414 ( .B(clk), .A(\g.we_clk [23360]));
Q_ASSIGN U9415 ( .B(clk), .A(\g.we_clk [23359]));
Q_ASSIGN U9416 ( .B(clk), .A(\g.we_clk [23358]));
Q_ASSIGN U9417 ( .B(clk), .A(\g.we_clk [23357]));
Q_ASSIGN U9418 ( .B(clk), .A(\g.we_clk [23356]));
Q_ASSIGN U9419 ( .B(clk), .A(\g.we_clk [23355]));
Q_ASSIGN U9420 ( .B(clk), .A(\g.we_clk [23354]));
Q_ASSIGN U9421 ( .B(clk), .A(\g.we_clk [23353]));
Q_ASSIGN U9422 ( .B(clk), .A(\g.we_clk [23352]));
Q_ASSIGN U9423 ( .B(clk), .A(\g.we_clk [23351]));
Q_ASSIGN U9424 ( .B(clk), .A(\g.we_clk [23350]));
Q_ASSIGN U9425 ( .B(clk), .A(\g.we_clk [23349]));
Q_ASSIGN U9426 ( .B(clk), .A(\g.we_clk [23348]));
Q_ASSIGN U9427 ( .B(clk), .A(\g.we_clk [23347]));
Q_ASSIGN U9428 ( .B(clk), .A(\g.we_clk [23346]));
Q_ASSIGN U9429 ( .B(clk), .A(\g.we_clk [23345]));
Q_ASSIGN U9430 ( .B(clk), .A(\g.we_clk [23344]));
Q_ASSIGN U9431 ( .B(clk), .A(\g.we_clk [23343]));
Q_ASSIGN U9432 ( .B(clk), .A(\g.we_clk [23342]));
Q_ASSIGN U9433 ( .B(clk), .A(\g.we_clk [23341]));
Q_ASSIGN U9434 ( .B(clk), .A(\g.we_clk [23340]));
Q_ASSIGN U9435 ( .B(clk), .A(\g.we_clk [23339]));
Q_ASSIGN U9436 ( .B(clk), .A(\g.we_clk [23338]));
Q_ASSIGN U9437 ( .B(clk), .A(\g.we_clk [23337]));
Q_ASSIGN U9438 ( .B(clk), .A(\g.we_clk [23336]));
Q_ASSIGN U9439 ( .B(clk), .A(\g.we_clk [23335]));
Q_ASSIGN U9440 ( .B(clk), .A(\g.we_clk [23334]));
Q_ASSIGN U9441 ( .B(clk), .A(\g.we_clk [23333]));
Q_ASSIGN U9442 ( .B(clk), .A(\g.we_clk [23332]));
Q_ASSIGN U9443 ( .B(clk), .A(\g.we_clk [23331]));
Q_ASSIGN U9444 ( .B(clk), .A(\g.we_clk [23330]));
Q_ASSIGN U9445 ( .B(clk), .A(\g.we_clk [23329]));
Q_ASSIGN U9446 ( .B(clk), .A(\g.we_clk [23328]));
Q_ASSIGN U9447 ( .B(clk), .A(\g.we_clk [23327]));
Q_ASSIGN U9448 ( .B(clk), .A(\g.we_clk [23326]));
Q_ASSIGN U9449 ( .B(clk), .A(\g.we_clk [23325]));
Q_ASSIGN U9450 ( .B(clk), .A(\g.we_clk [23324]));
Q_ASSIGN U9451 ( .B(clk), .A(\g.we_clk [23323]));
Q_ASSIGN U9452 ( .B(clk), .A(\g.we_clk [23322]));
Q_ASSIGN U9453 ( .B(clk), .A(\g.we_clk [23321]));
Q_ASSIGN U9454 ( .B(clk), .A(\g.we_clk [23320]));
Q_ASSIGN U9455 ( .B(clk), .A(\g.we_clk [23319]));
Q_ASSIGN U9456 ( .B(clk), .A(\g.we_clk [23318]));
Q_ASSIGN U9457 ( .B(clk), .A(\g.we_clk [23317]));
Q_ASSIGN U9458 ( .B(clk), .A(\g.we_clk [23316]));
Q_ASSIGN U9459 ( .B(clk), .A(\g.we_clk [23315]));
Q_ASSIGN U9460 ( .B(clk), .A(\g.we_clk [23314]));
Q_ASSIGN U9461 ( .B(clk), .A(\g.we_clk [23313]));
Q_ASSIGN U9462 ( .B(clk), .A(\g.we_clk [23312]));
Q_ASSIGN U9463 ( .B(clk), .A(\g.we_clk [23311]));
Q_ASSIGN U9464 ( .B(clk), .A(\g.we_clk [23310]));
Q_ASSIGN U9465 ( .B(clk), .A(\g.we_clk [23309]));
Q_ASSIGN U9466 ( .B(clk), .A(\g.we_clk [23308]));
Q_ASSIGN U9467 ( .B(clk), .A(\g.we_clk [23307]));
Q_ASSIGN U9468 ( .B(clk), .A(\g.we_clk [23306]));
Q_ASSIGN U9469 ( .B(clk), .A(\g.we_clk [23305]));
Q_ASSIGN U9470 ( .B(clk), .A(\g.we_clk [23304]));
Q_ASSIGN U9471 ( .B(clk), .A(\g.we_clk [23303]));
Q_ASSIGN U9472 ( .B(clk), .A(\g.we_clk [23302]));
Q_ASSIGN U9473 ( .B(clk), .A(\g.we_clk [23301]));
Q_ASSIGN U9474 ( .B(clk), .A(\g.we_clk [23300]));
Q_ASSIGN U9475 ( .B(clk), .A(\g.we_clk [23299]));
Q_ASSIGN U9476 ( .B(clk), .A(\g.we_clk [23298]));
Q_ASSIGN U9477 ( .B(clk), .A(\g.we_clk [23297]));
Q_ASSIGN U9478 ( .B(clk), .A(\g.we_clk [23296]));
Q_ASSIGN U9479 ( .B(clk), .A(\g.we_clk [23295]));
Q_ASSIGN U9480 ( .B(clk), .A(\g.we_clk [23294]));
Q_ASSIGN U9481 ( .B(clk), .A(\g.we_clk [23293]));
Q_ASSIGN U9482 ( .B(clk), .A(\g.we_clk [23292]));
Q_ASSIGN U9483 ( .B(clk), .A(\g.we_clk [23291]));
Q_ASSIGN U9484 ( .B(clk), .A(\g.we_clk [23290]));
Q_ASSIGN U9485 ( .B(clk), .A(\g.we_clk [23289]));
Q_ASSIGN U9486 ( .B(clk), .A(\g.we_clk [23288]));
Q_ASSIGN U9487 ( .B(clk), .A(\g.we_clk [23287]));
Q_ASSIGN U9488 ( .B(clk), .A(\g.we_clk [23286]));
Q_ASSIGN U9489 ( .B(clk), .A(\g.we_clk [23285]));
Q_ASSIGN U9490 ( .B(clk), .A(\g.we_clk [23284]));
Q_ASSIGN U9491 ( .B(clk), .A(\g.we_clk [23283]));
Q_ASSIGN U9492 ( .B(clk), .A(\g.we_clk [23282]));
Q_ASSIGN U9493 ( .B(clk), .A(\g.we_clk [23281]));
Q_ASSIGN U9494 ( .B(clk), .A(\g.we_clk [23280]));
Q_ASSIGN U9495 ( .B(clk), .A(\g.we_clk [23279]));
Q_ASSIGN U9496 ( .B(clk), .A(\g.we_clk [23278]));
Q_ASSIGN U9497 ( .B(clk), .A(\g.we_clk [23277]));
Q_ASSIGN U9498 ( .B(clk), .A(\g.we_clk [23276]));
Q_ASSIGN U9499 ( .B(clk), .A(\g.we_clk [23275]));
Q_ASSIGN U9500 ( .B(clk), .A(\g.we_clk [23274]));
Q_ASSIGN U9501 ( .B(clk), .A(\g.we_clk [23273]));
Q_ASSIGN U9502 ( .B(clk), .A(\g.we_clk [23272]));
Q_ASSIGN U9503 ( .B(clk), .A(\g.we_clk [23271]));
Q_ASSIGN U9504 ( .B(clk), .A(\g.we_clk [23270]));
Q_ASSIGN U9505 ( .B(clk), .A(\g.we_clk [23269]));
Q_ASSIGN U9506 ( .B(clk), .A(\g.we_clk [23268]));
Q_ASSIGN U9507 ( .B(clk), .A(\g.we_clk [23267]));
Q_ASSIGN U9508 ( .B(clk), .A(\g.we_clk [23266]));
Q_ASSIGN U9509 ( .B(clk), .A(\g.we_clk [23265]));
Q_ASSIGN U9510 ( .B(clk), .A(\g.we_clk [23264]));
Q_ASSIGN U9511 ( .B(clk), .A(\g.we_clk [23263]));
Q_ASSIGN U9512 ( .B(clk), .A(\g.we_clk [23262]));
Q_ASSIGN U9513 ( .B(clk), .A(\g.we_clk [23261]));
Q_ASSIGN U9514 ( .B(clk), .A(\g.we_clk [23260]));
Q_ASSIGN U9515 ( .B(clk), .A(\g.we_clk [23259]));
Q_ASSIGN U9516 ( .B(clk), .A(\g.we_clk [23258]));
Q_ASSIGN U9517 ( .B(clk), .A(\g.we_clk [23257]));
Q_ASSIGN U9518 ( .B(clk), .A(\g.we_clk [23256]));
Q_ASSIGN U9519 ( .B(clk), .A(\g.we_clk [23255]));
Q_ASSIGN U9520 ( .B(clk), .A(\g.we_clk [23254]));
Q_ASSIGN U9521 ( .B(clk), .A(\g.we_clk [23253]));
Q_ASSIGN U9522 ( .B(clk), .A(\g.we_clk [23252]));
Q_ASSIGN U9523 ( .B(clk), .A(\g.we_clk [23251]));
Q_ASSIGN U9524 ( .B(clk), .A(\g.we_clk [23250]));
Q_ASSIGN U9525 ( .B(clk), .A(\g.we_clk [23249]));
Q_ASSIGN U9526 ( .B(clk), .A(\g.we_clk [23248]));
Q_ASSIGN U9527 ( .B(clk), .A(\g.we_clk [23247]));
Q_ASSIGN U9528 ( .B(clk), .A(\g.we_clk [23246]));
Q_ASSIGN U9529 ( .B(clk), .A(\g.we_clk [23245]));
Q_ASSIGN U9530 ( .B(clk), .A(\g.we_clk [23244]));
Q_ASSIGN U9531 ( .B(clk), .A(\g.we_clk [23243]));
Q_ASSIGN U9532 ( .B(clk), .A(\g.we_clk [23242]));
Q_ASSIGN U9533 ( .B(clk), .A(\g.we_clk [23241]));
Q_ASSIGN U9534 ( .B(clk), .A(\g.we_clk [23240]));
Q_ASSIGN U9535 ( .B(clk), .A(\g.we_clk [23239]));
Q_ASSIGN U9536 ( .B(clk), .A(\g.we_clk [23238]));
Q_ASSIGN U9537 ( .B(clk), .A(\g.we_clk [23237]));
Q_ASSIGN U9538 ( .B(clk), .A(\g.we_clk [23236]));
Q_ASSIGN U9539 ( .B(clk), .A(\g.we_clk [23235]));
Q_ASSIGN U9540 ( .B(clk), .A(\g.we_clk [23234]));
Q_ASSIGN U9541 ( .B(clk), .A(\g.we_clk [23233]));
Q_ASSIGN U9542 ( .B(clk), .A(\g.we_clk [23232]));
Q_ASSIGN U9543 ( .B(clk), .A(\g.we_clk [23231]));
Q_ASSIGN U9544 ( .B(clk), .A(\g.we_clk [23230]));
Q_ASSIGN U9545 ( .B(clk), .A(\g.we_clk [23229]));
Q_ASSIGN U9546 ( .B(clk), .A(\g.we_clk [23228]));
Q_ASSIGN U9547 ( .B(clk), .A(\g.we_clk [23227]));
Q_ASSIGN U9548 ( .B(clk), .A(\g.we_clk [23226]));
Q_ASSIGN U9549 ( .B(clk), .A(\g.we_clk [23225]));
Q_ASSIGN U9550 ( .B(clk), .A(\g.we_clk [23224]));
Q_ASSIGN U9551 ( .B(clk), .A(\g.we_clk [23223]));
Q_ASSIGN U9552 ( .B(clk), .A(\g.we_clk [23222]));
Q_ASSIGN U9553 ( .B(clk), .A(\g.we_clk [23221]));
Q_ASSIGN U9554 ( .B(clk), .A(\g.we_clk [23220]));
Q_ASSIGN U9555 ( .B(clk), .A(\g.we_clk [23219]));
Q_ASSIGN U9556 ( .B(clk), .A(\g.we_clk [23218]));
Q_ASSIGN U9557 ( .B(clk), .A(\g.we_clk [23217]));
Q_ASSIGN U9558 ( .B(clk), .A(\g.we_clk [23216]));
Q_ASSIGN U9559 ( .B(clk), .A(\g.we_clk [23215]));
Q_ASSIGN U9560 ( .B(clk), .A(\g.we_clk [23214]));
Q_ASSIGN U9561 ( .B(clk), .A(\g.we_clk [23213]));
Q_ASSIGN U9562 ( .B(clk), .A(\g.we_clk [23212]));
Q_ASSIGN U9563 ( .B(clk), .A(\g.we_clk [23211]));
Q_ASSIGN U9564 ( .B(clk), .A(\g.we_clk [23210]));
Q_ASSIGN U9565 ( .B(clk), .A(\g.we_clk [23209]));
Q_ASSIGN U9566 ( .B(clk), .A(\g.we_clk [23208]));
Q_ASSIGN U9567 ( .B(clk), .A(\g.we_clk [23207]));
Q_ASSIGN U9568 ( .B(clk), .A(\g.we_clk [23206]));
Q_ASSIGN U9569 ( .B(clk), .A(\g.we_clk [23205]));
Q_ASSIGN U9570 ( .B(clk), .A(\g.we_clk [23204]));
Q_ASSIGN U9571 ( .B(clk), .A(\g.we_clk [23203]));
Q_ASSIGN U9572 ( .B(clk), .A(\g.we_clk [23202]));
Q_ASSIGN U9573 ( .B(clk), .A(\g.we_clk [23201]));
Q_ASSIGN U9574 ( .B(clk), .A(\g.we_clk [23200]));
Q_ASSIGN U9575 ( .B(clk), .A(\g.we_clk [23199]));
Q_ASSIGN U9576 ( .B(clk), .A(\g.we_clk [23198]));
Q_ASSIGN U9577 ( .B(clk), .A(\g.we_clk [23197]));
Q_ASSIGN U9578 ( .B(clk), .A(\g.we_clk [23196]));
Q_ASSIGN U9579 ( .B(clk), .A(\g.we_clk [23195]));
Q_ASSIGN U9580 ( .B(clk), .A(\g.we_clk [23194]));
Q_ASSIGN U9581 ( .B(clk), .A(\g.we_clk [23193]));
Q_ASSIGN U9582 ( .B(clk), .A(\g.we_clk [23192]));
Q_ASSIGN U9583 ( .B(clk), .A(\g.we_clk [23191]));
Q_ASSIGN U9584 ( .B(clk), .A(\g.we_clk [23190]));
Q_ASSIGN U9585 ( .B(clk), .A(\g.we_clk [23189]));
Q_ASSIGN U9586 ( .B(clk), .A(\g.we_clk [23188]));
Q_ASSIGN U9587 ( .B(clk), .A(\g.we_clk [23187]));
Q_ASSIGN U9588 ( .B(clk), .A(\g.we_clk [23186]));
Q_ASSIGN U9589 ( .B(clk), .A(\g.we_clk [23185]));
Q_ASSIGN U9590 ( .B(clk), .A(\g.we_clk [23184]));
Q_ASSIGN U9591 ( .B(clk), .A(\g.we_clk [23183]));
Q_ASSIGN U9592 ( .B(clk), .A(\g.we_clk [23182]));
Q_ASSIGN U9593 ( .B(clk), .A(\g.we_clk [23181]));
Q_ASSIGN U9594 ( .B(clk), .A(\g.we_clk [23180]));
Q_ASSIGN U9595 ( .B(clk), .A(\g.we_clk [23179]));
Q_ASSIGN U9596 ( .B(clk), .A(\g.we_clk [23178]));
Q_ASSIGN U9597 ( .B(clk), .A(\g.we_clk [23177]));
Q_ASSIGN U9598 ( .B(clk), .A(\g.we_clk [23176]));
Q_ASSIGN U9599 ( .B(clk), .A(\g.we_clk [23175]));
Q_ASSIGN U9600 ( .B(clk), .A(\g.we_clk [23174]));
Q_ASSIGN U9601 ( .B(clk), .A(\g.we_clk [23173]));
Q_ASSIGN U9602 ( .B(clk), .A(\g.we_clk [23172]));
Q_ASSIGN U9603 ( .B(clk), .A(\g.we_clk [23171]));
Q_ASSIGN U9604 ( .B(clk), .A(\g.we_clk [23170]));
Q_ASSIGN U9605 ( .B(clk), .A(\g.we_clk [23169]));
Q_ASSIGN U9606 ( .B(clk), .A(\g.we_clk [23168]));
Q_ASSIGN U9607 ( .B(clk), .A(\g.we_clk [23167]));
Q_ASSIGN U9608 ( .B(clk), .A(\g.we_clk [23166]));
Q_ASSIGN U9609 ( .B(clk), .A(\g.we_clk [23165]));
Q_ASSIGN U9610 ( .B(clk), .A(\g.we_clk [23164]));
Q_ASSIGN U9611 ( .B(clk), .A(\g.we_clk [23163]));
Q_ASSIGN U9612 ( .B(clk), .A(\g.we_clk [23162]));
Q_ASSIGN U9613 ( .B(clk), .A(\g.we_clk [23161]));
Q_ASSIGN U9614 ( .B(clk), .A(\g.we_clk [23160]));
Q_ASSIGN U9615 ( .B(clk), .A(\g.we_clk [23159]));
Q_ASSIGN U9616 ( .B(clk), .A(\g.we_clk [23158]));
Q_ASSIGN U9617 ( .B(clk), .A(\g.we_clk [23157]));
Q_ASSIGN U9618 ( .B(clk), .A(\g.we_clk [23156]));
Q_ASSIGN U9619 ( .B(clk), .A(\g.we_clk [23155]));
Q_ASSIGN U9620 ( .B(clk), .A(\g.we_clk [23154]));
Q_ASSIGN U9621 ( .B(clk), .A(\g.we_clk [23153]));
Q_ASSIGN U9622 ( .B(clk), .A(\g.we_clk [23152]));
Q_ASSIGN U9623 ( .B(clk), .A(\g.we_clk [23151]));
Q_ASSIGN U9624 ( .B(clk), .A(\g.we_clk [23150]));
Q_ASSIGN U9625 ( .B(clk), .A(\g.we_clk [23149]));
Q_ASSIGN U9626 ( .B(clk), .A(\g.we_clk [23148]));
Q_ASSIGN U9627 ( .B(clk), .A(\g.we_clk [23147]));
Q_ASSIGN U9628 ( .B(clk), .A(\g.we_clk [23146]));
Q_ASSIGN U9629 ( .B(clk), .A(\g.we_clk [23145]));
Q_ASSIGN U9630 ( .B(clk), .A(\g.we_clk [23144]));
Q_ASSIGN U9631 ( .B(clk), .A(\g.we_clk [23143]));
Q_ASSIGN U9632 ( .B(clk), .A(\g.we_clk [23142]));
Q_ASSIGN U9633 ( .B(clk), .A(\g.we_clk [23141]));
Q_ASSIGN U9634 ( .B(clk), .A(\g.we_clk [23140]));
Q_ASSIGN U9635 ( .B(clk), .A(\g.we_clk [23139]));
Q_ASSIGN U9636 ( .B(clk), .A(\g.we_clk [23138]));
Q_ASSIGN U9637 ( .B(clk), .A(\g.we_clk [23137]));
Q_ASSIGN U9638 ( .B(clk), .A(\g.we_clk [23136]));
Q_ASSIGN U9639 ( .B(clk), .A(\g.we_clk [23135]));
Q_ASSIGN U9640 ( .B(clk), .A(\g.we_clk [23134]));
Q_ASSIGN U9641 ( .B(clk), .A(\g.we_clk [23133]));
Q_ASSIGN U9642 ( .B(clk), .A(\g.we_clk [23132]));
Q_ASSIGN U9643 ( .B(clk), .A(\g.we_clk [23131]));
Q_ASSIGN U9644 ( .B(clk), .A(\g.we_clk [23130]));
Q_ASSIGN U9645 ( .B(clk), .A(\g.we_clk [23129]));
Q_ASSIGN U9646 ( .B(clk), .A(\g.we_clk [23128]));
Q_ASSIGN U9647 ( .B(clk), .A(\g.we_clk [23127]));
Q_ASSIGN U9648 ( .B(clk), .A(\g.we_clk [23126]));
Q_ASSIGN U9649 ( .B(clk), .A(\g.we_clk [23125]));
Q_ASSIGN U9650 ( .B(clk), .A(\g.we_clk [23124]));
Q_ASSIGN U9651 ( .B(clk), .A(\g.we_clk [23123]));
Q_ASSIGN U9652 ( .B(clk), .A(\g.we_clk [23122]));
Q_ASSIGN U9653 ( .B(clk), .A(\g.we_clk [23121]));
Q_ASSIGN U9654 ( .B(clk), .A(\g.we_clk [23120]));
Q_ASSIGN U9655 ( .B(clk), .A(\g.we_clk [23119]));
Q_ASSIGN U9656 ( .B(clk), .A(\g.we_clk [23118]));
Q_ASSIGN U9657 ( .B(clk), .A(\g.we_clk [23117]));
Q_ASSIGN U9658 ( .B(clk), .A(\g.we_clk [23116]));
Q_ASSIGN U9659 ( .B(clk), .A(\g.we_clk [23115]));
Q_ASSIGN U9660 ( .B(clk), .A(\g.we_clk [23114]));
Q_ASSIGN U9661 ( .B(clk), .A(\g.we_clk [23113]));
Q_ASSIGN U9662 ( .B(clk), .A(\g.we_clk [23112]));
Q_ASSIGN U9663 ( .B(clk), .A(\g.we_clk [23111]));
Q_ASSIGN U9664 ( .B(clk), .A(\g.we_clk [23110]));
Q_ASSIGN U9665 ( .B(clk), .A(\g.we_clk [23109]));
Q_ASSIGN U9666 ( .B(clk), .A(\g.we_clk [23108]));
Q_ASSIGN U9667 ( .B(clk), .A(\g.we_clk [23107]));
Q_ASSIGN U9668 ( .B(clk), .A(\g.we_clk [23106]));
Q_ASSIGN U9669 ( .B(clk), .A(\g.we_clk [23105]));
Q_ASSIGN U9670 ( .B(clk), .A(\g.we_clk [23104]));
Q_ASSIGN U9671 ( .B(clk), .A(\g.we_clk [23103]));
Q_ASSIGN U9672 ( .B(clk), .A(\g.we_clk [23102]));
Q_ASSIGN U9673 ( .B(clk), .A(\g.we_clk [23101]));
Q_ASSIGN U9674 ( .B(clk), .A(\g.we_clk [23100]));
Q_ASSIGN U9675 ( .B(clk), .A(\g.we_clk [23099]));
Q_ASSIGN U9676 ( .B(clk), .A(\g.we_clk [23098]));
Q_ASSIGN U9677 ( .B(clk), .A(\g.we_clk [23097]));
Q_ASSIGN U9678 ( .B(clk), .A(\g.we_clk [23096]));
Q_ASSIGN U9679 ( .B(clk), .A(\g.we_clk [23095]));
Q_ASSIGN U9680 ( .B(clk), .A(\g.we_clk [23094]));
Q_ASSIGN U9681 ( .B(clk), .A(\g.we_clk [23093]));
Q_ASSIGN U9682 ( .B(clk), .A(\g.we_clk [23092]));
Q_ASSIGN U9683 ( .B(clk), .A(\g.we_clk [23091]));
Q_ASSIGN U9684 ( .B(clk), .A(\g.we_clk [23090]));
Q_ASSIGN U9685 ( .B(clk), .A(\g.we_clk [23089]));
Q_ASSIGN U9686 ( .B(clk), .A(\g.we_clk [23088]));
Q_ASSIGN U9687 ( .B(clk), .A(\g.we_clk [23087]));
Q_ASSIGN U9688 ( .B(clk), .A(\g.we_clk [23086]));
Q_ASSIGN U9689 ( .B(clk), .A(\g.we_clk [23085]));
Q_ASSIGN U9690 ( .B(clk), .A(\g.we_clk [23084]));
Q_ASSIGN U9691 ( .B(clk), .A(\g.we_clk [23083]));
Q_ASSIGN U9692 ( .B(clk), .A(\g.we_clk [23082]));
Q_ASSIGN U9693 ( .B(clk), .A(\g.we_clk [23081]));
Q_ASSIGN U9694 ( .B(clk), .A(\g.we_clk [23080]));
Q_ASSIGN U9695 ( .B(clk), .A(\g.we_clk [23079]));
Q_ASSIGN U9696 ( .B(clk), .A(\g.we_clk [23078]));
Q_ASSIGN U9697 ( .B(clk), .A(\g.we_clk [23077]));
Q_ASSIGN U9698 ( .B(clk), .A(\g.we_clk [23076]));
Q_ASSIGN U9699 ( .B(clk), .A(\g.we_clk [23075]));
Q_ASSIGN U9700 ( .B(clk), .A(\g.we_clk [23074]));
Q_ASSIGN U9701 ( .B(clk), .A(\g.we_clk [23073]));
Q_ASSIGN U9702 ( .B(clk), .A(\g.we_clk [23072]));
Q_ASSIGN U9703 ( .B(clk), .A(\g.we_clk [23071]));
Q_ASSIGN U9704 ( .B(clk), .A(\g.we_clk [23070]));
Q_ASSIGN U9705 ( .B(clk), .A(\g.we_clk [23069]));
Q_ASSIGN U9706 ( .B(clk), .A(\g.we_clk [23068]));
Q_ASSIGN U9707 ( .B(clk), .A(\g.we_clk [23067]));
Q_ASSIGN U9708 ( .B(clk), .A(\g.we_clk [23066]));
Q_ASSIGN U9709 ( .B(clk), .A(\g.we_clk [23065]));
Q_ASSIGN U9710 ( .B(clk), .A(\g.we_clk [23064]));
Q_ASSIGN U9711 ( .B(clk), .A(\g.we_clk [23063]));
Q_ASSIGN U9712 ( .B(clk), .A(\g.we_clk [23062]));
Q_ASSIGN U9713 ( .B(clk), .A(\g.we_clk [23061]));
Q_ASSIGN U9714 ( .B(clk), .A(\g.we_clk [23060]));
Q_ASSIGN U9715 ( .B(clk), .A(\g.we_clk [23059]));
Q_ASSIGN U9716 ( .B(clk), .A(\g.we_clk [23058]));
Q_ASSIGN U9717 ( .B(clk), .A(\g.we_clk [23057]));
Q_ASSIGN U9718 ( .B(clk), .A(\g.we_clk [23056]));
Q_ASSIGN U9719 ( .B(clk), .A(\g.we_clk [23055]));
Q_ASSIGN U9720 ( .B(clk), .A(\g.we_clk [23054]));
Q_ASSIGN U9721 ( .B(clk), .A(\g.we_clk [23053]));
Q_ASSIGN U9722 ( .B(clk), .A(\g.we_clk [23052]));
Q_ASSIGN U9723 ( .B(clk), .A(\g.we_clk [23051]));
Q_ASSIGN U9724 ( .B(clk), .A(\g.we_clk [23050]));
Q_ASSIGN U9725 ( .B(clk), .A(\g.we_clk [23049]));
Q_ASSIGN U9726 ( .B(clk), .A(\g.we_clk [23048]));
Q_ASSIGN U9727 ( .B(clk), .A(\g.we_clk [23047]));
Q_ASSIGN U9728 ( .B(clk), .A(\g.we_clk [23046]));
Q_ASSIGN U9729 ( .B(clk), .A(\g.we_clk [23045]));
Q_ASSIGN U9730 ( .B(clk), .A(\g.we_clk [23044]));
Q_ASSIGN U9731 ( .B(clk), .A(\g.we_clk [23043]));
Q_ASSIGN U9732 ( .B(clk), .A(\g.we_clk [23042]));
Q_ASSIGN U9733 ( .B(clk), .A(\g.we_clk [23041]));
Q_ASSIGN U9734 ( .B(clk), .A(\g.we_clk [23040]));
Q_ASSIGN U9735 ( .B(clk), .A(\g.we_clk [23039]));
Q_ASSIGN U9736 ( .B(clk), .A(\g.we_clk [23038]));
Q_ASSIGN U9737 ( .B(clk), .A(\g.we_clk [23037]));
Q_ASSIGN U9738 ( .B(clk), .A(\g.we_clk [23036]));
Q_ASSIGN U9739 ( .B(clk), .A(\g.we_clk [23035]));
Q_ASSIGN U9740 ( .B(clk), .A(\g.we_clk [23034]));
Q_ASSIGN U9741 ( .B(clk), .A(\g.we_clk [23033]));
Q_ASSIGN U9742 ( .B(clk), .A(\g.we_clk [23032]));
Q_ASSIGN U9743 ( .B(clk), .A(\g.we_clk [23031]));
Q_ASSIGN U9744 ( .B(clk), .A(\g.we_clk [23030]));
Q_ASSIGN U9745 ( .B(clk), .A(\g.we_clk [23029]));
Q_ASSIGN U9746 ( .B(clk), .A(\g.we_clk [23028]));
Q_ASSIGN U9747 ( .B(clk), .A(\g.we_clk [23027]));
Q_ASSIGN U9748 ( .B(clk), .A(\g.we_clk [23026]));
Q_ASSIGN U9749 ( .B(clk), .A(\g.we_clk [23025]));
Q_ASSIGN U9750 ( .B(clk), .A(\g.we_clk [23024]));
Q_ASSIGN U9751 ( .B(clk), .A(\g.we_clk [23023]));
Q_ASSIGN U9752 ( .B(clk), .A(\g.we_clk [23022]));
Q_ASSIGN U9753 ( .B(clk), .A(\g.we_clk [23021]));
Q_ASSIGN U9754 ( .B(clk), .A(\g.we_clk [23020]));
Q_ASSIGN U9755 ( .B(clk), .A(\g.we_clk [23019]));
Q_ASSIGN U9756 ( .B(clk), .A(\g.we_clk [23018]));
Q_ASSIGN U9757 ( .B(clk), .A(\g.we_clk [23017]));
Q_ASSIGN U9758 ( .B(clk), .A(\g.we_clk [23016]));
Q_ASSIGN U9759 ( .B(clk), .A(\g.we_clk [23015]));
Q_ASSIGN U9760 ( .B(clk), .A(\g.we_clk [23014]));
Q_ASSIGN U9761 ( .B(clk), .A(\g.we_clk [23013]));
Q_ASSIGN U9762 ( .B(clk), .A(\g.we_clk [23012]));
Q_ASSIGN U9763 ( .B(clk), .A(\g.we_clk [23011]));
Q_ASSIGN U9764 ( .B(clk), .A(\g.we_clk [23010]));
Q_ASSIGN U9765 ( .B(clk), .A(\g.we_clk [23009]));
Q_ASSIGN U9766 ( .B(clk), .A(\g.we_clk [23008]));
Q_ASSIGN U9767 ( .B(clk), .A(\g.we_clk [23007]));
Q_ASSIGN U9768 ( .B(clk), .A(\g.we_clk [23006]));
Q_ASSIGN U9769 ( .B(clk), .A(\g.we_clk [23005]));
Q_ASSIGN U9770 ( .B(clk), .A(\g.we_clk [23004]));
Q_ASSIGN U9771 ( .B(clk), .A(\g.we_clk [23003]));
Q_ASSIGN U9772 ( .B(clk), .A(\g.we_clk [23002]));
Q_ASSIGN U9773 ( .B(clk), .A(\g.we_clk [23001]));
Q_ASSIGN U9774 ( .B(clk), .A(\g.we_clk [23000]));
Q_ASSIGN U9775 ( .B(clk), .A(\g.we_clk [22999]));
Q_ASSIGN U9776 ( .B(clk), .A(\g.we_clk [22998]));
Q_ASSIGN U9777 ( .B(clk), .A(\g.we_clk [22997]));
Q_ASSIGN U9778 ( .B(clk), .A(\g.we_clk [22996]));
Q_ASSIGN U9779 ( .B(clk), .A(\g.we_clk [22995]));
Q_ASSIGN U9780 ( .B(clk), .A(\g.we_clk [22994]));
Q_ASSIGN U9781 ( .B(clk), .A(\g.we_clk [22993]));
Q_ASSIGN U9782 ( .B(clk), .A(\g.we_clk [22992]));
Q_ASSIGN U9783 ( .B(clk), .A(\g.we_clk [22991]));
Q_ASSIGN U9784 ( .B(clk), .A(\g.we_clk [22990]));
Q_ASSIGN U9785 ( .B(clk), .A(\g.we_clk [22989]));
Q_ASSIGN U9786 ( .B(clk), .A(\g.we_clk [22988]));
Q_ASSIGN U9787 ( .B(clk), .A(\g.we_clk [22987]));
Q_ASSIGN U9788 ( .B(clk), .A(\g.we_clk [22986]));
Q_ASSIGN U9789 ( .B(clk), .A(\g.we_clk [22985]));
Q_ASSIGN U9790 ( .B(clk), .A(\g.we_clk [22984]));
Q_ASSIGN U9791 ( .B(clk), .A(\g.we_clk [22983]));
Q_ASSIGN U9792 ( .B(clk), .A(\g.we_clk [22982]));
Q_ASSIGN U9793 ( .B(clk), .A(\g.we_clk [22981]));
Q_ASSIGN U9794 ( .B(clk), .A(\g.we_clk [22980]));
Q_ASSIGN U9795 ( .B(clk), .A(\g.we_clk [22979]));
Q_ASSIGN U9796 ( .B(clk), .A(\g.we_clk [22978]));
Q_ASSIGN U9797 ( .B(clk), .A(\g.we_clk [22977]));
Q_ASSIGN U9798 ( .B(clk), .A(\g.we_clk [22976]));
Q_ASSIGN U9799 ( .B(clk), .A(\g.we_clk [22975]));
Q_ASSIGN U9800 ( .B(clk), .A(\g.we_clk [22974]));
Q_ASSIGN U9801 ( .B(clk), .A(\g.we_clk [22973]));
Q_ASSIGN U9802 ( .B(clk), .A(\g.we_clk [22972]));
Q_ASSIGN U9803 ( .B(clk), .A(\g.we_clk [22971]));
Q_ASSIGN U9804 ( .B(clk), .A(\g.we_clk [22970]));
Q_ASSIGN U9805 ( .B(clk), .A(\g.we_clk [22969]));
Q_ASSIGN U9806 ( .B(clk), .A(\g.we_clk [22968]));
Q_ASSIGN U9807 ( .B(clk), .A(\g.we_clk [22967]));
Q_ASSIGN U9808 ( .B(clk), .A(\g.we_clk [22966]));
Q_ASSIGN U9809 ( .B(clk), .A(\g.we_clk [22965]));
Q_ASSIGN U9810 ( .B(clk), .A(\g.we_clk [22964]));
Q_ASSIGN U9811 ( .B(clk), .A(\g.we_clk [22963]));
Q_ASSIGN U9812 ( .B(clk), .A(\g.we_clk [22962]));
Q_ASSIGN U9813 ( .B(clk), .A(\g.we_clk [22961]));
Q_ASSIGN U9814 ( .B(clk), .A(\g.we_clk [22960]));
Q_ASSIGN U9815 ( .B(clk), .A(\g.we_clk [22959]));
Q_ASSIGN U9816 ( .B(clk), .A(\g.we_clk [22958]));
Q_ASSIGN U9817 ( .B(clk), .A(\g.we_clk [22957]));
Q_ASSIGN U9818 ( .B(clk), .A(\g.we_clk [22956]));
Q_ASSIGN U9819 ( .B(clk), .A(\g.we_clk [22955]));
Q_ASSIGN U9820 ( .B(clk), .A(\g.we_clk [22954]));
Q_ASSIGN U9821 ( .B(clk), .A(\g.we_clk [22953]));
Q_ASSIGN U9822 ( .B(clk), .A(\g.we_clk [22952]));
Q_ASSIGN U9823 ( .B(clk), .A(\g.we_clk [22951]));
Q_ASSIGN U9824 ( .B(clk), .A(\g.we_clk [22950]));
Q_ASSIGN U9825 ( .B(clk), .A(\g.we_clk [22949]));
Q_ASSIGN U9826 ( .B(clk), .A(\g.we_clk [22948]));
Q_ASSIGN U9827 ( .B(clk), .A(\g.we_clk [22947]));
Q_ASSIGN U9828 ( .B(clk), .A(\g.we_clk [22946]));
Q_ASSIGN U9829 ( .B(clk), .A(\g.we_clk [22945]));
Q_ASSIGN U9830 ( .B(clk), .A(\g.we_clk [22944]));
Q_ASSIGN U9831 ( .B(clk), .A(\g.we_clk [22943]));
Q_ASSIGN U9832 ( .B(clk), .A(\g.we_clk [22942]));
Q_ASSIGN U9833 ( .B(clk), .A(\g.we_clk [22941]));
Q_ASSIGN U9834 ( .B(clk), .A(\g.we_clk [22940]));
Q_ASSIGN U9835 ( .B(clk), .A(\g.we_clk [22939]));
Q_ASSIGN U9836 ( .B(clk), .A(\g.we_clk [22938]));
Q_ASSIGN U9837 ( .B(clk), .A(\g.we_clk [22937]));
Q_ASSIGN U9838 ( .B(clk), .A(\g.we_clk [22936]));
Q_ASSIGN U9839 ( .B(clk), .A(\g.we_clk [22935]));
Q_ASSIGN U9840 ( .B(clk), .A(\g.we_clk [22934]));
Q_ASSIGN U9841 ( .B(clk), .A(\g.we_clk [22933]));
Q_ASSIGN U9842 ( .B(clk), .A(\g.we_clk [22932]));
Q_ASSIGN U9843 ( .B(clk), .A(\g.we_clk [22931]));
Q_ASSIGN U9844 ( .B(clk), .A(\g.we_clk [22930]));
Q_ASSIGN U9845 ( .B(clk), .A(\g.we_clk [22929]));
Q_ASSIGN U9846 ( .B(clk), .A(\g.we_clk [22928]));
Q_ASSIGN U9847 ( .B(clk), .A(\g.we_clk [22927]));
Q_ASSIGN U9848 ( .B(clk), .A(\g.we_clk [22926]));
Q_ASSIGN U9849 ( .B(clk), .A(\g.we_clk [22925]));
Q_ASSIGN U9850 ( .B(clk), .A(\g.we_clk [22924]));
Q_ASSIGN U9851 ( .B(clk), .A(\g.we_clk [22923]));
Q_ASSIGN U9852 ( .B(clk), .A(\g.we_clk [22922]));
Q_ASSIGN U9853 ( .B(clk), .A(\g.we_clk [22921]));
Q_ASSIGN U9854 ( .B(clk), .A(\g.we_clk [22920]));
Q_ASSIGN U9855 ( .B(clk), .A(\g.we_clk [22919]));
Q_ASSIGN U9856 ( .B(clk), .A(\g.we_clk [22918]));
Q_ASSIGN U9857 ( .B(clk), .A(\g.we_clk [22917]));
Q_ASSIGN U9858 ( .B(clk), .A(\g.we_clk [22916]));
Q_ASSIGN U9859 ( .B(clk), .A(\g.we_clk [22915]));
Q_ASSIGN U9860 ( .B(clk), .A(\g.we_clk [22914]));
Q_ASSIGN U9861 ( .B(clk), .A(\g.we_clk [22913]));
Q_ASSIGN U9862 ( .B(clk), .A(\g.we_clk [22912]));
Q_ASSIGN U9863 ( .B(clk), .A(\g.we_clk [22911]));
Q_ASSIGN U9864 ( .B(clk), .A(\g.we_clk [22910]));
Q_ASSIGN U9865 ( .B(clk), .A(\g.we_clk [22909]));
Q_ASSIGN U9866 ( .B(clk), .A(\g.we_clk [22908]));
Q_ASSIGN U9867 ( .B(clk), .A(\g.we_clk [22907]));
Q_ASSIGN U9868 ( .B(clk), .A(\g.we_clk [22906]));
Q_ASSIGN U9869 ( .B(clk), .A(\g.we_clk [22905]));
Q_ASSIGN U9870 ( .B(clk), .A(\g.we_clk [22904]));
Q_ASSIGN U9871 ( .B(clk), .A(\g.we_clk [22903]));
Q_ASSIGN U9872 ( .B(clk), .A(\g.we_clk [22902]));
Q_ASSIGN U9873 ( .B(clk), .A(\g.we_clk [22901]));
Q_ASSIGN U9874 ( .B(clk), .A(\g.we_clk [22900]));
Q_ASSIGN U9875 ( .B(clk), .A(\g.we_clk [22899]));
Q_ASSIGN U9876 ( .B(clk), .A(\g.we_clk [22898]));
Q_ASSIGN U9877 ( .B(clk), .A(\g.we_clk [22897]));
Q_ASSIGN U9878 ( .B(clk), .A(\g.we_clk [22896]));
Q_ASSIGN U9879 ( .B(clk), .A(\g.we_clk [22895]));
Q_ASSIGN U9880 ( .B(clk), .A(\g.we_clk [22894]));
Q_ASSIGN U9881 ( .B(clk), .A(\g.we_clk [22893]));
Q_ASSIGN U9882 ( .B(clk), .A(\g.we_clk [22892]));
Q_ASSIGN U9883 ( .B(clk), .A(\g.we_clk [22891]));
Q_ASSIGN U9884 ( .B(clk), .A(\g.we_clk [22890]));
Q_ASSIGN U9885 ( .B(clk), .A(\g.we_clk [22889]));
Q_ASSIGN U9886 ( .B(clk), .A(\g.we_clk [22888]));
Q_ASSIGN U9887 ( .B(clk), .A(\g.we_clk [22887]));
Q_ASSIGN U9888 ( .B(clk), .A(\g.we_clk [22886]));
Q_ASSIGN U9889 ( .B(clk), .A(\g.we_clk [22885]));
Q_ASSIGN U9890 ( .B(clk), .A(\g.we_clk [22884]));
Q_ASSIGN U9891 ( .B(clk), .A(\g.we_clk [22883]));
Q_ASSIGN U9892 ( .B(clk), .A(\g.we_clk [22882]));
Q_ASSIGN U9893 ( .B(clk), .A(\g.we_clk [22881]));
Q_ASSIGN U9894 ( .B(clk), .A(\g.we_clk [22880]));
Q_ASSIGN U9895 ( .B(clk), .A(\g.we_clk [22879]));
Q_ASSIGN U9896 ( .B(clk), .A(\g.we_clk [22878]));
Q_ASSIGN U9897 ( .B(clk), .A(\g.we_clk [22877]));
Q_ASSIGN U9898 ( .B(clk), .A(\g.we_clk [22876]));
Q_ASSIGN U9899 ( .B(clk), .A(\g.we_clk [22875]));
Q_ASSIGN U9900 ( .B(clk), .A(\g.we_clk [22874]));
Q_ASSIGN U9901 ( .B(clk), .A(\g.we_clk [22873]));
Q_ASSIGN U9902 ( .B(clk), .A(\g.we_clk [22872]));
Q_ASSIGN U9903 ( .B(clk), .A(\g.we_clk [22871]));
Q_ASSIGN U9904 ( .B(clk), .A(\g.we_clk [22870]));
Q_ASSIGN U9905 ( .B(clk), .A(\g.we_clk [22869]));
Q_ASSIGN U9906 ( .B(clk), .A(\g.we_clk [22868]));
Q_ASSIGN U9907 ( .B(clk), .A(\g.we_clk [22867]));
Q_ASSIGN U9908 ( .B(clk), .A(\g.we_clk [22866]));
Q_ASSIGN U9909 ( .B(clk), .A(\g.we_clk [22865]));
Q_ASSIGN U9910 ( .B(clk), .A(\g.we_clk [22864]));
Q_ASSIGN U9911 ( .B(clk), .A(\g.we_clk [22863]));
Q_ASSIGN U9912 ( .B(clk), .A(\g.we_clk [22862]));
Q_ASSIGN U9913 ( .B(clk), .A(\g.we_clk [22861]));
Q_ASSIGN U9914 ( .B(clk), .A(\g.we_clk [22860]));
Q_ASSIGN U9915 ( .B(clk), .A(\g.we_clk [22859]));
Q_ASSIGN U9916 ( .B(clk), .A(\g.we_clk [22858]));
Q_ASSIGN U9917 ( .B(clk), .A(\g.we_clk [22857]));
Q_ASSIGN U9918 ( .B(clk), .A(\g.we_clk [22856]));
Q_ASSIGN U9919 ( .B(clk), .A(\g.we_clk [22855]));
Q_ASSIGN U9920 ( .B(clk), .A(\g.we_clk [22854]));
Q_ASSIGN U9921 ( .B(clk), .A(\g.we_clk [22853]));
Q_ASSIGN U9922 ( .B(clk), .A(\g.we_clk [22852]));
Q_ASSIGN U9923 ( .B(clk), .A(\g.we_clk [22851]));
Q_ASSIGN U9924 ( .B(clk), .A(\g.we_clk [22850]));
Q_ASSIGN U9925 ( .B(clk), .A(\g.we_clk [22849]));
Q_ASSIGN U9926 ( .B(clk), .A(\g.we_clk [22848]));
Q_ASSIGN U9927 ( .B(clk), .A(\g.we_clk [22847]));
Q_ASSIGN U9928 ( .B(clk), .A(\g.we_clk [22846]));
Q_ASSIGN U9929 ( .B(clk), .A(\g.we_clk [22845]));
Q_ASSIGN U9930 ( .B(clk), .A(\g.we_clk [22844]));
Q_ASSIGN U9931 ( .B(clk), .A(\g.we_clk [22843]));
Q_ASSIGN U9932 ( .B(clk), .A(\g.we_clk [22842]));
Q_ASSIGN U9933 ( .B(clk), .A(\g.we_clk [22841]));
Q_ASSIGN U9934 ( .B(clk), .A(\g.we_clk [22840]));
Q_ASSIGN U9935 ( .B(clk), .A(\g.we_clk [22839]));
Q_ASSIGN U9936 ( .B(clk), .A(\g.we_clk [22838]));
Q_ASSIGN U9937 ( .B(clk), .A(\g.we_clk [22837]));
Q_ASSIGN U9938 ( .B(clk), .A(\g.we_clk [22836]));
Q_ASSIGN U9939 ( .B(clk), .A(\g.we_clk [22835]));
Q_ASSIGN U9940 ( .B(clk), .A(\g.we_clk [22834]));
Q_ASSIGN U9941 ( .B(clk), .A(\g.we_clk [22833]));
Q_ASSIGN U9942 ( .B(clk), .A(\g.we_clk [22832]));
Q_ASSIGN U9943 ( .B(clk), .A(\g.we_clk [22831]));
Q_ASSIGN U9944 ( .B(clk), .A(\g.we_clk [22830]));
Q_ASSIGN U9945 ( .B(clk), .A(\g.we_clk [22829]));
Q_ASSIGN U9946 ( .B(clk), .A(\g.we_clk [22828]));
Q_ASSIGN U9947 ( .B(clk), .A(\g.we_clk [22827]));
Q_ASSIGN U9948 ( .B(clk), .A(\g.we_clk [22826]));
Q_ASSIGN U9949 ( .B(clk), .A(\g.we_clk [22825]));
Q_ASSIGN U9950 ( .B(clk), .A(\g.we_clk [22824]));
Q_ASSIGN U9951 ( .B(clk), .A(\g.we_clk [22823]));
Q_ASSIGN U9952 ( .B(clk), .A(\g.we_clk [22822]));
Q_ASSIGN U9953 ( .B(clk), .A(\g.we_clk [22821]));
Q_ASSIGN U9954 ( .B(clk), .A(\g.we_clk [22820]));
Q_ASSIGN U9955 ( .B(clk), .A(\g.we_clk [22819]));
Q_ASSIGN U9956 ( .B(clk), .A(\g.we_clk [22818]));
Q_ASSIGN U9957 ( .B(clk), .A(\g.we_clk [22817]));
Q_ASSIGN U9958 ( .B(clk), .A(\g.we_clk [22816]));
Q_ASSIGN U9959 ( .B(clk), .A(\g.we_clk [22815]));
Q_ASSIGN U9960 ( .B(clk), .A(\g.we_clk [22814]));
Q_ASSIGN U9961 ( .B(clk), .A(\g.we_clk [22813]));
Q_ASSIGN U9962 ( .B(clk), .A(\g.we_clk [22812]));
Q_ASSIGN U9963 ( .B(clk), .A(\g.we_clk [22811]));
Q_ASSIGN U9964 ( .B(clk), .A(\g.we_clk [22810]));
Q_ASSIGN U9965 ( .B(clk), .A(\g.we_clk [22809]));
Q_ASSIGN U9966 ( .B(clk), .A(\g.we_clk [22808]));
Q_ASSIGN U9967 ( .B(clk), .A(\g.we_clk [22807]));
Q_ASSIGN U9968 ( .B(clk), .A(\g.we_clk [22806]));
Q_ASSIGN U9969 ( .B(clk), .A(\g.we_clk [22805]));
Q_ASSIGN U9970 ( .B(clk), .A(\g.we_clk [22804]));
Q_ASSIGN U9971 ( .B(clk), .A(\g.we_clk [22803]));
Q_ASSIGN U9972 ( .B(clk), .A(\g.we_clk [22802]));
Q_ASSIGN U9973 ( .B(clk), .A(\g.we_clk [22801]));
Q_ASSIGN U9974 ( .B(clk), .A(\g.we_clk [22800]));
Q_ASSIGN U9975 ( .B(clk), .A(\g.we_clk [22799]));
Q_ASSIGN U9976 ( .B(clk), .A(\g.we_clk [22798]));
Q_ASSIGN U9977 ( .B(clk), .A(\g.we_clk [22797]));
Q_ASSIGN U9978 ( .B(clk), .A(\g.we_clk [22796]));
Q_ASSIGN U9979 ( .B(clk), .A(\g.we_clk [22795]));
Q_ASSIGN U9980 ( .B(clk), .A(\g.we_clk [22794]));
Q_ASSIGN U9981 ( .B(clk), .A(\g.we_clk [22793]));
Q_ASSIGN U9982 ( .B(clk), .A(\g.we_clk [22792]));
Q_ASSIGN U9983 ( .B(clk), .A(\g.we_clk [22791]));
Q_ASSIGN U9984 ( .B(clk), .A(\g.we_clk [22790]));
Q_ASSIGN U9985 ( .B(clk), .A(\g.we_clk [22789]));
Q_ASSIGN U9986 ( .B(clk), .A(\g.we_clk [22788]));
Q_ASSIGN U9987 ( .B(clk), .A(\g.we_clk [22787]));
Q_ASSIGN U9988 ( .B(clk), .A(\g.we_clk [22786]));
Q_ASSIGN U9989 ( .B(clk), .A(\g.we_clk [22785]));
Q_ASSIGN U9990 ( .B(clk), .A(\g.we_clk [22784]));
Q_ASSIGN U9991 ( .B(clk), .A(\g.we_clk [22783]));
Q_ASSIGN U9992 ( .B(clk), .A(\g.we_clk [22782]));
Q_ASSIGN U9993 ( .B(clk), .A(\g.we_clk [22781]));
Q_ASSIGN U9994 ( .B(clk), .A(\g.we_clk [22780]));
Q_ASSIGN U9995 ( .B(clk), .A(\g.we_clk [22779]));
Q_ASSIGN U9996 ( .B(clk), .A(\g.we_clk [22778]));
Q_ASSIGN U9997 ( .B(clk), .A(\g.we_clk [22777]));
Q_ASSIGN U9998 ( .B(clk), .A(\g.we_clk [22776]));
Q_ASSIGN U9999 ( .B(clk), .A(\g.we_clk [22775]));
Q_ASSIGN U10000 ( .B(clk), .A(\g.we_clk [22774]));
Q_ASSIGN U10001 ( .B(clk), .A(\g.we_clk [22773]));
Q_ASSIGN U10002 ( .B(clk), .A(\g.we_clk [22772]));
Q_ASSIGN U10003 ( .B(clk), .A(\g.we_clk [22771]));
Q_ASSIGN U10004 ( .B(clk), .A(\g.we_clk [22770]));
Q_ASSIGN U10005 ( .B(clk), .A(\g.we_clk [22769]));
Q_ASSIGN U10006 ( .B(clk), .A(\g.we_clk [22768]));
Q_ASSIGN U10007 ( .B(clk), .A(\g.we_clk [22767]));
Q_ASSIGN U10008 ( .B(clk), .A(\g.we_clk [22766]));
Q_ASSIGN U10009 ( .B(clk), .A(\g.we_clk [22765]));
Q_ASSIGN U10010 ( .B(clk), .A(\g.we_clk [22764]));
Q_ASSIGN U10011 ( .B(clk), .A(\g.we_clk [22763]));
Q_ASSIGN U10012 ( .B(clk), .A(\g.we_clk [22762]));
Q_ASSIGN U10013 ( .B(clk), .A(\g.we_clk [22761]));
Q_ASSIGN U10014 ( .B(clk), .A(\g.we_clk [22760]));
Q_ASSIGN U10015 ( .B(clk), .A(\g.we_clk [22759]));
Q_ASSIGN U10016 ( .B(clk), .A(\g.we_clk [22758]));
Q_ASSIGN U10017 ( .B(clk), .A(\g.we_clk [22757]));
Q_ASSIGN U10018 ( .B(clk), .A(\g.we_clk [22756]));
Q_ASSIGN U10019 ( .B(clk), .A(\g.we_clk [22755]));
Q_ASSIGN U10020 ( .B(clk), .A(\g.we_clk [22754]));
Q_ASSIGN U10021 ( .B(clk), .A(\g.we_clk [22753]));
Q_ASSIGN U10022 ( .B(clk), .A(\g.we_clk [22752]));
Q_ASSIGN U10023 ( .B(clk), .A(\g.we_clk [22751]));
Q_ASSIGN U10024 ( .B(clk), .A(\g.we_clk [22750]));
Q_ASSIGN U10025 ( .B(clk), .A(\g.we_clk [22749]));
Q_ASSIGN U10026 ( .B(clk), .A(\g.we_clk [22748]));
Q_ASSIGN U10027 ( .B(clk), .A(\g.we_clk [22747]));
Q_ASSIGN U10028 ( .B(clk), .A(\g.we_clk [22746]));
Q_ASSIGN U10029 ( .B(clk), .A(\g.we_clk [22745]));
Q_ASSIGN U10030 ( .B(clk), .A(\g.we_clk [22744]));
Q_ASSIGN U10031 ( .B(clk), .A(\g.we_clk [22743]));
Q_ASSIGN U10032 ( .B(clk), .A(\g.we_clk [22742]));
Q_ASSIGN U10033 ( .B(clk), .A(\g.we_clk [22741]));
Q_ASSIGN U10034 ( .B(clk), .A(\g.we_clk [22740]));
Q_ASSIGN U10035 ( .B(clk), .A(\g.we_clk [22739]));
Q_ASSIGN U10036 ( .B(clk), .A(\g.we_clk [22738]));
Q_ASSIGN U10037 ( .B(clk), .A(\g.we_clk [22737]));
Q_ASSIGN U10038 ( .B(clk), .A(\g.we_clk [22736]));
Q_ASSIGN U10039 ( .B(clk), .A(\g.we_clk [22735]));
Q_ASSIGN U10040 ( .B(clk), .A(\g.we_clk [22734]));
Q_ASSIGN U10041 ( .B(clk), .A(\g.we_clk [22733]));
Q_ASSIGN U10042 ( .B(clk), .A(\g.we_clk [22732]));
Q_ASSIGN U10043 ( .B(clk), .A(\g.we_clk [22731]));
Q_ASSIGN U10044 ( .B(clk), .A(\g.we_clk [22730]));
Q_ASSIGN U10045 ( .B(clk), .A(\g.we_clk [22729]));
Q_ASSIGN U10046 ( .B(clk), .A(\g.we_clk [22728]));
Q_ASSIGN U10047 ( .B(clk), .A(\g.we_clk [22727]));
Q_ASSIGN U10048 ( .B(clk), .A(\g.we_clk [22726]));
Q_ASSIGN U10049 ( .B(clk), .A(\g.we_clk [22725]));
Q_ASSIGN U10050 ( .B(clk), .A(\g.we_clk [22724]));
Q_ASSIGN U10051 ( .B(clk), .A(\g.we_clk [22723]));
Q_ASSIGN U10052 ( .B(clk), .A(\g.we_clk [22722]));
Q_ASSIGN U10053 ( .B(clk), .A(\g.we_clk [22721]));
Q_ASSIGN U10054 ( .B(clk), .A(\g.we_clk [22720]));
Q_ASSIGN U10055 ( .B(clk), .A(\g.we_clk [22719]));
Q_ASSIGN U10056 ( .B(clk), .A(\g.we_clk [22718]));
Q_ASSIGN U10057 ( .B(clk), .A(\g.we_clk [22717]));
Q_ASSIGN U10058 ( .B(clk), .A(\g.we_clk [22716]));
Q_ASSIGN U10059 ( .B(clk), .A(\g.we_clk [22715]));
Q_ASSIGN U10060 ( .B(clk), .A(\g.we_clk [22714]));
Q_ASSIGN U10061 ( .B(clk), .A(\g.we_clk [22713]));
Q_ASSIGN U10062 ( .B(clk), .A(\g.we_clk [22712]));
Q_ASSIGN U10063 ( .B(clk), .A(\g.we_clk [22711]));
Q_ASSIGN U10064 ( .B(clk), .A(\g.we_clk [22710]));
Q_ASSIGN U10065 ( .B(clk), .A(\g.we_clk [22709]));
Q_ASSIGN U10066 ( .B(clk), .A(\g.we_clk [22708]));
Q_ASSIGN U10067 ( .B(clk), .A(\g.we_clk [22707]));
Q_ASSIGN U10068 ( .B(clk), .A(\g.we_clk [22706]));
Q_ASSIGN U10069 ( .B(clk), .A(\g.we_clk [22705]));
Q_ASSIGN U10070 ( .B(clk), .A(\g.we_clk [22704]));
Q_ASSIGN U10071 ( .B(clk), .A(\g.we_clk [22703]));
Q_ASSIGN U10072 ( .B(clk), .A(\g.we_clk [22702]));
Q_ASSIGN U10073 ( .B(clk), .A(\g.we_clk [22701]));
Q_ASSIGN U10074 ( .B(clk), .A(\g.we_clk [22700]));
Q_ASSIGN U10075 ( .B(clk), .A(\g.we_clk [22699]));
Q_ASSIGN U10076 ( .B(clk), .A(\g.we_clk [22698]));
Q_ASSIGN U10077 ( .B(clk), .A(\g.we_clk [22697]));
Q_ASSIGN U10078 ( .B(clk), .A(\g.we_clk [22696]));
Q_ASSIGN U10079 ( .B(clk), .A(\g.we_clk [22695]));
Q_ASSIGN U10080 ( .B(clk), .A(\g.we_clk [22694]));
Q_ASSIGN U10081 ( .B(clk), .A(\g.we_clk [22693]));
Q_ASSIGN U10082 ( .B(clk), .A(\g.we_clk [22692]));
Q_ASSIGN U10083 ( .B(clk), .A(\g.we_clk [22691]));
Q_ASSIGN U10084 ( .B(clk), .A(\g.we_clk [22690]));
Q_ASSIGN U10085 ( .B(clk), .A(\g.we_clk [22689]));
Q_ASSIGN U10086 ( .B(clk), .A(\g.we_clk [22688]));
Q_ASSIGN U10087 ( .B(clk), .A(\g.we_clk [22687]));
Q_ASSIGN U10088 ( .B(clk), .A(\g.we_clk [22686]));
Q_ASSIGN U10089 ( .B(clk), .A(\g.we_clk [22685]));
Q_ASSIGN U10090 ( .B(clk), .A(\g.we_clk [22684]));
Q_ASSIGN U10091 ( .B(clk), .A(\g.we_clk [22683]));
Q_ASSIGN U10092 ( .B(clk), .A(\g.we_clk [22682]));
Q_ASSIGN U10093 ( .B(clk), .A(\g.we_clk [22681]));
Q_ASSIGN U10094 ( .B(clk), .A(\g.we_clk [22680]));
Q_ASSIGN U10095 ( .B(clk), .A(\g.we_clk [22679]));
Q_ASSIGN U10096 ( .B(clk), .A(\g.we_clk [22678]));
Q_ASSIGN U10097 ( .B(clk), .A(\g.we_clk [22677]));
Q_ASSIGN U10098 ( .B(clk), .A(\g.we_clk [22676]));
Q_ASSIGN U10099 ( .B(clk), .A(\g.we_clk [22675]));
Q_ASSIGN U10100 ( .B(clk), .A(\g.we_clk [22674]));
Q_ASSIGN U10101 ( .B(clk), .A(\g.we_clk [22673]));
Q_ASSIGN U10102 ( .B(clk), .A(\g.we_clk [22672]));
Q_ASSIGN U10103 ( .B(clk), .A(\g.we_clk [22671]));
Q_ASSIGN U10104 ( .B(clk), .A(\g.we_clk [22670]));
Q_ASSIGN U10105 ( .B(clk), .A(\g.we_clk [22669]));
Q_ASSIGN U10106 ( .B(clk), .A(\g.we_clk [22668]));
Q_ASSIGN U10107 ( .B(clk), .A(\g.we_clk [22667]));
Q_ASSIGN U10108 ( .B(clk), .A(\g.we_clk [22666]));
Q_ASSIGN U10109 ( .B(clk), .A(\g.we_clk [22665]));
Q_ASSIGN U10110 ( .B(clk), .A(\g.we_clk [22664]));
Q_ASSIGN U10111 ( .B(clk), .A(\g.we_clk [22663]));
Q_ASSIGN U10112 ( .B(clk), .A(\g.we_clk [22662]));
Q_ASSIGN U10113 ( .B(clk), .A(\g.we_clk [22661]));
Q_ASSIGN U10114 ( .B(clk), .A(\g.we_clk [22660]));
Q_ASSIGN U10115 ( .B(clk), .A(\g.we_clk [22659]));
Q_ASSIGN U10116 ( .B(clk), .A(\g.we_clk [22658]));
Q_ASSIGN U10117 ( .B(clk), .A(\g.we_clk [22657]));
Q_ASSIGN U10118 ( .B(clk), .A(\g.we_clk [22656]));
Q_ASSIGN U10119 ( .B(clk), .A(\g.we_clk [22655]));
Q_ASSIGN U10120 ( .B(clk), .A(\g.we_clk [22654]));
Q_ASSIGN U10121 ( .B(clk), .A(\g.we_clk [22653]));
Q_ASSIGN U10122 ( .B(clk), .A(\g.we_clk [22652]));
Q_ASSIGN U10123 ( .B(clk), .A(\g.we_clk [22651]));
Q_ASSIGN U10124 ( .B(clk), .A(\g.we_clk [22650]));
Q_ASSIGN U10125 ( .B(clk), .A(\g.we_clk [22649]));
Q_ASSIGN U10126 ( .B(clk), .A(\g.we_clk [22648]));
Q_ASSIGN U10127 ( .B(clk), .A(\g.we_clk [22647]));
Q_ASSIGN U10128 ( .B(clk), .A(\g.we_clk [22646]));
Q_ASSIGN U10129 ( .B(clk), .A(\g.we_clk [22645]));
Q_ASSIGN U10130 ( .B(clk), .A(\g.we_clk [22644]));
Q_ASSIGN U10131 ( .B(clk), .A(\g.we_clk [22643]));
Q_ASSIGN U10132 ( .B(clk), .A(\g.we_clk [22642]));
Q_ASSIGN U10133 ( .B(clk), .A(\g.we_clk [22641]));
Q_ASSIGN U10134 ( .B(clk), .A(\g.we_clk [22640]));
Q_ASSIGN U10135 ( .B(clk), .A(\g.we_clk [22639]));
Q_ASSIGN U10136 ( .B(clk), .A(\g.we_clk [22638]));
Q_ASSIGN U10137 ( .B(clk), .A(\g.we_clk [22637]));
Q_ASSIGN U10138 ( .B(clk), .A(\g.we_clk [22636]));
Q_ASSIGN U10139 ( .B(clk), .A(\g.we_clk [22635]));
Q_ASSIGN U10140 ( .B(clk), .A(\g.we_clk [22634]));
Q_ASSIGN U10141 ( .B(clk), .A(\g.we_clk [22633]));
Q_ASSIGN U10142 ( .B(clk), .A(\g.we_clk [22632]));
Q_ASSIGN U10143 ( .B(clk), .A(\g.we_clk [22631]));
Q_ASSIGN U10144 ( .B(clk), .A(\g.we_clk [22630]));
Q_ASSIGN U10145 ( .B(clk), .A(\g.we_clk [22629]));
Q_ASSIGN U10146 ( .B(clk), .A(\g.we_clk [22628]));
Q_ASSIGN U10147 ( .B(clk), .A(\g.we_clk [22627]));
Q_ASSIGN U10148 ( .B(clk), .A(\g.we_clk [22626]));
Q_ASSIGN U10149 ( .B(clk), .A(\g.we_clk [22625]));
Q_ASSIGN U10150 ( .B(clk), .A(\g.we_clk [22624]));
Q_ASSIGN U10151 ( .B(clk), .A(\g.we_clk [22623]));
Q_ASSIGN U10152 ( .B(clk), .A(\g.we_clk [22622]));
Q_ASSIGN U10153 ( .B(clk), .A(\g.we_clk [22621]));
Q_ASSIGN U10154 ( .B(clk), .A(\g.we_clk [22620]));
Q_ASSIGN U10155 ( .B(clk), .A(\g.we_clk [22619]));
Q_ASSIGN U10156 ( .B(clk), .A(\g.we_clk [22618]));
Q_ASSIGN U10157 ( .B(clk), .A(\g.we_clk [22617]));
Q_ASSIGN U10158 ( .B(clk), .A(\g.we_clk [22616]));
Q_ASSIGN U10159 ( .B(clk), .A(\g.we_clk [22615]));
Q_ASSIGN U10160 ( .B(clk), .A(\g.we_clk [22614]));
Q_ASSIGN U10161 ( .B(clk), .A(\g.we_clk [22613]));
Q_ASSIGN U10162 ( .B(clk), .A(\g.we_clk [22612]));
Q_ASSIGN U10163 ( .B(clk), .A(\g.we_clk [22611]));
Q_ASSIGN U10164 ( .B(clk), .A(\g.we_clk [22610]));
Q_ASSIGN U10165 ( .B(clk), .A(\g.we_clk [22609]));
Q_ASSIGN U10166 ( .B(clk), .A(\g.we_clk [22608]));
Q_ASSIGN U10167 ( .B(clk), .A(\g.we_clk [22607]));
Q_ASSIGN U10168 ( .B(clk), .A(\g.we_clk [22606]));
Q_ASSIGN U10169 ( .B(clk), .A(\g.we_clk [22605]));
Q_ASSIGN U10170 ( .B(clk), .A(\g.we_clk [22604]));
Q_ASSIGN U10171 ( .B(clk), .A(\g.we_clk [22603]));
Q_ASSIGN U10172 ( .B(clk), .A(\g.we_clk [22602]));
Q_ASSIGN U10173 ( .B(clk), .A(\g.we_clk [22601]));
Q_ASSIGN U10174 ( .B(clk), .A(\g.we_clk [22600]));
Q_ASSIGN U10175 ( .B(clk), .A(\g.we_clk [22599]));
Q_ASSIGN U10176 ( .B(clk), .A(\g.we_clk [22598]));
Q_ASSIGN U10177 ( .B(clk), .A(\g.we_clk [22597]));
Q_ASSIGN U10178 ( .B(clk), .A(\g.we_clk [22596]));
Q_ASSIGN U10179 ( .B(clk), .A(\g.we_clk [22595]));
Q_ASSIGN U10180 ( .B(clk), .A(\g.we_clk [22594]));
Q_ASSIGN U10181 ( .B(clk), .A(\g.we_clk [22593]));
Q_ASSIGN U10182 ( .B(clk), .A(\g.we_clk [22592]));
Q_ASSIGN U10183 ( .B(clk), .A(\g.we_clk [22591]));
Q_ASSIGN U10184 ( .B(clk), .A(\g.we_clk [22590]));
Q_ASSIGN U10185 ( .B(clk), .A(\g.we_clk [22589]));
Q_ASSIGN U10186 ( .B(clk), .A(\g.we_clk [22588]));
Q_ASSIGN U10187 ( .B(clk), .A(\g.we_clk [22587]));
Q_ASSIGN U10188 ( .B(clk), .A(\g.we_clk [22586]));
Q_ASSIGN U10189 ( .B(clk), .A(\g.we_clk [22585]));
Q_ASSIGN U10190 ( .B(clk), .A(\g.we_clk [22584]));
Q_ASSIGN U10191 ( .B(clk), .A(\g.we_clk [22583]));
Q_ASSIGN U10192 ( .B(clk), .A(\g.we_clk [22582]));
Q_ASSIGN U10193 ( .B(clk), .A(\g.we_clk [22581]));
Q_ASSIGN U10194 ( .B(clk), .A(\g.we_clk [22580]));
Q_ASSIGN U10195 ( .B(clk), .A(\g.we_clk [22579]));
Q_ASSIGN U10196 ( .B(clk), .A(\g.we_clk [22578]));
Q_ASSIGN U10197 ( .B(clk), .A(\g.we_clk [22577]));
Q_ASSIGN U10198 ( .B(clk), .A(\g.we_clk [22576]));
Q_ASSIGN U10199 ( .B(clk), .A(\g.we_clk [22575]));
Q_ASSIGN U10200 ( .B(clk), .A(\g.we_clk [22574]));
Q_ASSIGN U10201 ( .B(clk), .A(\g.we_clk [22573]));
Q_ASSIGN U10202 ( .B(clk), .A(\g.we_clk [22572]));
Q_ASSIGN U10203 ( .B(clk), .A(\g.we_clk [22571]));
Q_ASSIGN U10204 ( .B(clk), .A(\g.we_clk [22570]));
Q_ASSIGN U10205 ( .B(clk), .A(\g.we_clk [22569]));
Q_ASSIGN U10206 ( .B(clk), .A(\g.we_clk [22568]));
Q_ASSIGN U10207 ( .B(clk), .A(\g.we_clk [22567]));
Q_ASSIGN U10208 ( .B(clk), .A(\g.we_clk [22566]));
Q_ASSIGN U10209 ( .B(clk), .A(\g.we_clk [22565]));
Q_ASSIGN U10210 ( .B(clk), .A(\g.we_clk [22564]));
Q_ASSIGN U10211 ( .B(clk), .A(\g.we_clk [22563]));
Q_ASSIGN U10212 ( .B(clk), .A(\g.we_clk [22562]));
Q_ASSIGN U10213 ( .B(clk), .A(\g.we_clk [22561]));
Q_ASSIGN U10214 ( .B(clk), .A(\g.we_clk [22560]));
Q_ASSIGN U10215 ( .B(clk), .A(\g.we_clk [22559]));
Q_ASSIGN U10216 ( .B(clk), .A(\g.we_clk [22558]));
Q_ASSIGN U10217 ( .B(clk), .A(\g.we_clk [22557]));
Q_ASSIGN U10218 ( .B(clk), .A(\g.we_clk [22556]));
Q_ASSIGN U10219 ( .B(clk), .A(\g.we_clk [22555]));
Q_ASSIGN U10220 ( .B(clk), .A(\g.we_clk [22554]));
Q_ASSIGN U10221 ( .B(clk), .A(\g.we_clk [22553]));
Q_ASSIGN U10222 ( .B(clk), .A(\g.we_clk [22552]));
Q_ASSIGN U10223 ( .B(clk), .A(\g.we_clk [22551]));
Q_ASSIGN U10224 ( .B(clk), .A(\g.we_clk [22550]));
Q_ASSIGN U10225 ( .B(clk), .A(\g.we_clk [22549]));
Q_ASSIGN U10226 ( .B(clk), .A(\g.we_clk [22548]));
Q_ASSIGN U10227 ( .B(clk), .A(\g.we_clk [22547]));
Q_ASSIGN U10228 ( .B(clk), .A(\g.we_clk [22546]));
Q_ASSIGN U10229 ( .B(clk), .A(\g.we_clk [22545]));
Q_ASSIGN U10230 ( .B(clk), .A(\g.we_clk [22544]));
Q_ASSIGN U10231 ( .B(clk), .A(\g.we_clk [22543]));
Q_ASSIGN U10232 ( .B(clk), .A(\g.we_clk [22542]));
Q_ASSIGN U10233 ( .B(clk), .A(\g.we_clk [22541]));
Q_ASSIGN U10234 ( .B(clk), .A(\g.we_clk [22540]));
Q_ASSIGN U10235 ( .B(clk), .A(\g.we_clk [22539]));
Q_ASSIGN U10236 ( .B(clk), .A(\g.we_clk [22538]));
Q_ASSIGN U10237 ( .B(clk), .A(\g.we_clk [22537]));
Q_ASSIGN U10238 ( .B(clk), .A(\g.we_clk [22536]));
Q_ASSIGN U10239 ( .B(clk), .A(\g.we_clk [22535]));
Q_ASSIGN U10240 ( .B(clk), .A(\g.we_clk [22534]));
Q_ASSIGN U10241 ( .B(clk), .A(\g.we_clk [22533]));
Q_ASSIGN U10242 ( .B(clk), .A(\g.we_clk [22532]));
Q_ASSIGN U10243 ( .B(clk), .A(\g.we_clk [22531]));
Q_ASSIGN U10244 ( .B(clk), .A(\g.we_clk [22530]));
Q_ASSIGN U10245 ( .B(clk), .A(\g.we_clk [22529]));
Q_ASSIGN U10246 ( .B(clk), .A(\g.we_clk [22528]));
Q_ASSIGN U10247 ( .B(clk), .A(\g.we_clk [22527]));
Q_ASSIGN U10248 ( .B(clk), .A(\g.we_clk [22526]));
Q_ASSIGN U10249 ( .B(clk), .A(\g.we_clk [22525]));
Q_ASSIGN U10250 ( .B(clk), .A(\g.we_clk [22524]));
Q_ASSIGN U10251 ( .B(clk), .A(\g.we_clk [22523]));
Q_ASSIGN U10252 ( .B(clk), .A(\g.we_clk [22522]));
Q_ASSIGN U10253 ( .B(clk), .A(\g.we_clk [22521]));
Q_ASSIGN U10254 ( .B(clk), .A(\g.we_clk [22520]));
Q_ASSIGN U10255 ( .B(clk), .A(\g.we_clk [22519]));
Q_ASSIGN U10256 ( .B(clk), .A(\g.we_clk [22518]));
Q_ASSIGN U10257 ( .B(clk), .A(\g.we_clk [22517]));
Q_ASSIGN U10258 ( .B(clk), .A(\g.we_clk [22516]));
Q_ASSIGN U10259 ( .B(clk), .A(\g.we_clk [22515]));
Q_ASSIGN U10260 ( .B(clk), .A(\g.we_clk [22514]));
Q_ASSIGN U10261 ( .B(clk), .A(\g.we_clk [22513]));
Q_ASSIGN U10262 ( .B(clk), .A(\g.we_clk [22512]));
Q_ASSIGN U10263 ( .B(clk), .A(\g.we_clk [22511]));
Q_ASSIGN U10264 ( .B(clk), .A(\g.we_clk [22510]));
Q_ASSIGN U10265 ( .B(clk), .A(\g.we_clk [22509]));
Q_ASSIGN U10266 ( .B(clk), .A(\g.we_clk [22508]));
Q_ASSIGN U10267 ( .B(clk), .A(\g.we_clk [22507]));
Q_ASSIGN U10268 ( .B(clk), .A(\g.we_clk [22506]));
Q_ASSIGN U10269 ( .B(clk), .A(\g.we_clk [22505]));
Q_ASSIGN U10270 ( .B(clk), .A(\g.we_clk [22504]));
Q_ASSIGN U10271 ( .B(clk), .A(\g.we_clk [22503]));
Q_ASSIGN U10272 ( .B(clk), .A(\g.we_clk [22502]));
Q_ASSIGN U10273 ( .B(clk), .A(\g.we_clk [22501]));
Q_ASSIGN U10274 ( .B(clk), .A(\g.we_clk [22500]));
Q_ASSIGN U10275 ( .B(clk), .A(\g.we_clk [22499]));
Q_ASSIGN U10276 ( .B(clk), .A(\g.we_clk [22498]));
Q_ASSIGN U10277 ( .B(clk), .A(\g.we_clk [22497]));
Q_ASSIGN U10278 ( .B(clk), .A(\g.we_clk [22496]));
Q_ASSIGN U10279 ( .B(clk), .A(\g.we_clk [22495]));
Q_ASSIGN U10280 ( .B(clk), .A(\g.we_clk [22494]));
Q_ASSIGN U10281 ( .B(clk), .A(\g.we_clk [22493]));
Q_ASSIGN U10282 ( .B(clk), .A(\g.we_clk [22492]));
Q_ASSIGN U10283 ( .B(clk), .A(\g.we_clk [22491]));
Q_ASSIGN U10284 ( .B(clk), .A(\g.we_clk [22490]));
Q_ASSIGN U10285 ( .B(clk), .A(\g.we_clk [22489]));
Q_ASSIGN U10286 ( .B(clk), .A(\g.we_clk [22488]));
Q_ASSIGN U10287 ( .B(clk), .A(\g.we_clk [22487]));
Q_ASSIGN U10288 ( .B(clk), .A(\g.we_clk [22486]));
Q_ASSIGN U10289 ( .B(clk), .A(\g.we_clk [22485]));
Q_ASSIGN U10290 ( .B(clk), .A(\g.we_clk [22484]));
Q_ASSIGN U10291 ( .B(clk), .A(\g.we_clk [22483]));
Q_ASSIGN U10292 ( .B(clk), .A(\g.we_clk [22482]));
Q_ASSIGN U10293 ( .B(clk), .A(\g.we_clk [22481]));
Q_ASSIGN U10294 ( .B(clk), .A(\g.we_clk [22480]));
Q_ASSIGN U10295 ( .B(clk), .A(\g.we_clk [22479]));
Q_ASSIGN U10296 ( .B(clk), .A(\g.we_clk [22478]));
Q_ASSIGN U10297 ( .B(clk), .A(\g.we_clk [22477]));
Q_ASSIGN U10298 ( .B(clk), .A(\g.we_clk [22476]));
Q_ASSIGN U10299 ( .B(clk), .A(\g.we_clk [22475]));
Q_ASSIGN U10300 ( .B(clk), .A(\g.we_clk [22474]));
Q_ASSIGN U10301 ( .B(clk), .A(\g.we_clk [22473]));
Q_ASSIGN U10302 ( .B(clk), .A(\g.we_clk [22472]));
Q_ASSIGN U10303 ( .B(clk), .A(\g.we_clk [22471]));
Q_ASSIGN U10304 ( .B(clk), .A(\g.we_clk [22470]));
Q_ASSIGN U10305 ( .B(clk), .A(\g.we_clk [22469]));
Q_ASSIGN U10306 ( .B(clk), .A(\g.we_clk [22468]));
Q_ASSIGN U10307 ( .B(clk), .A(\g.we_clk [22467]));
Q_ASSIGN U10308 ( .B(clk), .A(\g.we_clk [22466]));
Q_ASSIGN U10309 ( .B(clk), .A(\g.we_clk [22465]));
Q_ASSIGN U10310 ( .B(clk), .A(\g.we_clk [22464]));
Q_ASSIGN U10311 ( .B(clk), .A(\g.we_clk [22463]));
Q_ASSIGN U10312 ( .B(clk), .A(\g.we_clk [22462]));
Q_ASSIGN U10313 ( .B(clk), .A(\g.we_clk [22461]));
Q_ASSIGN U10314 ( .B(clk), .A(\g.we_clk [22460]));
Q_ASSIGN U10315 ( .B(clk), .A(\g.we_clk [22459]));
Q_ASSIGN U10316 ( .B(clk), .A(\g.we_clk [22458]));
Q_ASSIGN U10317 ( .B(clk), .A(\g.we_clk [22457]));
Q_ASSIGN U10318 ( .B(clk), .A(\g.we_clk [22456]));
Q_ASSIGN U10319 ( .B(clk), .A(\g.we_clk [22455]));
Q_ASSIGN U10320 ( .B(clk), .A(\g.we_clk [22454]));
Q_ASSIGN U10321 ( .B(clk), .A(\g.we_clk [22453]));
Q_ASSIGN U10322 ( .B(clk), .A(\g.we_clk [22452]));
Q_ASSIGN U10323 ( .B(clk), .A(\g.we_clk [22451]));
Q_ASSIGN U10324 ( .B(clk), .A(\g.we_clk [22450]));
Q_ASSIGN U10325 ( .B(clk), .A(\g.we_clk [22449]));
Q_ASSIGN U10326 ( .B(clk), .A(\g.we_clk [22448]));
Q_ASSIGN U10327 ( .B(clk), .A(\g.we_clk [22447]));
Q_ASSIGN U10328 ( .B(clk), .A(\g.we_clk [22446]));
Q_ASSIGN U10329 ( .B(clk), .A(\g.we_clk [22445]));
Q_ASSIGN U10330 ( .B(clk), .A(\g.we_clk [22444]));
Q_ASSIGN U10331 ( .B(clk), .A(\g.we_clk [22443]));
Q_ASSIGN U10332 ( .B(clk), .A(\g.we_clk [22442]));
Q_ASSIGN U10333 ( .B(clk), .A(\g.we_clk [22441]));
Q_ASSIGN U10334 ( .B(clk), .A(\g.we_clk [22440]));
Q_ASSIGN U10335 ( .B(clk), .A(\g.we_clk [22439]));
Q_ASSIGN U10336 ( .B(clk), .A(\g.we_clk [22438]));
Q_ASSIGN U10337 ( .B(clk), .A(\g.we_clk [22437]));
Q_ASSIGN U10338 ( .B(clk), .A(\g.we_clk [22436]));
Q_ASSIGN U10339 ( .B(clk), .A(\g.we_clk [22435]));
Q_ASSIGN U10340 ( .B(clk), .A(\g.we_clk [22434]));
Q_ASSIGN U10341 ( .B(clk), .A(\g.we_clk [22433]));
Q_ASSIGN U10342 ( .B(clk), .A(\g.we_clk [22432]));
Q_ASSIGN U10343 ( .B(clk), .A(\g.we_clk [22431]));
Q_ASSIGN U10344 ( .B(clk), .A(\g.we_clk [22430]));
Q_ASSIGN U10345 ( .B(clk), .A(\g.we_clk [22429]));
Q_ASSIGN U10346 ( .B(clk), .A(\g.we_clk [22428]));
Q_ASSIGN U10347 ( .B(clk), .A(\g.we_clk [22427]));
Q_ASSIGN U10348 ( .B(clk), .A(\g.we_clk [22426]));
Q_ASSIGN U10349 ( .B(clk), .A(\g.we_clk [22425]));
Q_ASSIGN U10350 ( .B(clk), .A(\g.we_clk [22424]));
Q_ASSIGN U10351 ( .B(clk), .A(\g.we_clk [22423]));
Q_ASSIGN U10352 ( .B(clk), .A(\g.we_clk [22422]));
Q_ASSIGN U10353 ( .B(clk), .A(\g.we_clk [22421]));
Q_ASSIGN U10354 ( .B(clk), .A(\g.we_clk [22420]));
Q_ASSIGN U10355 ( .B(clk), .A(\g.we_clk [22419]));
Q_ASSIGN U10356 ( .B(clk), .A(\g.we_clk [22418]));
Q_ASSIGN U10357 ( .B(clk), .A(\g.we_clk [22417]));
Q_ASSIGN U10358 ( .B(clk), .A(\g.we_clk [22416]));
Q_ASSIGN U10359 ( .B(clk), .A(\g.we_clk [22415]));
Q_ASSIGN U10360 ( .B(clk), .A(\g.we_clk [22414]));
Q_ASSIGN U10361 ( .B(clk), .A(\g.we_clk [22413]));
Q_ASSIGN U10362 ( .B(clk), .A(\g.we_clk [22412]));
Q_ASSIGN U10363 ( .B(clk), .A(\g.we_clk [22411]));
Q_ASSIGN U10364 ( .B(clk), .A(\g.we_clk [22410]));
Q_ASSIGN U10365 ( .B(clk), .A(\g.we_clk [22409]));
Q_ASSIGN U10366 ( .B(clk), .A(\g.we_clk [22408]));
Q_ASSIGN U10367 ( .B(clk), .A(\g.we_clk [22407]));
Q_ASSIGN U10368 ( .B(clk), .A(\g.we_clk [22406]));
Q_ASSIGN U10369 ( .B(clk), .A(\g.we_clk [22405]));
Q_ASSIGN U10370 ( .B(clk), .A(\g.we_clk [22404]));
Q_ASSIGN U10371 ( .B(clk), .A(\g.we_clk [22403]));
Q_ASSIGN U10372 ( .B(clk), .A(\g.we_clk [22402]));
Q_ASSIGN U10373 ( .B(clk), .A(\g.we_clk [22401]));
Q_ASSIGN U10374 ( .B(clk), .A(\g.we_clk [22400]));
Q_ASSIGN U10375 ( .B(clk), .A(\g.we_clk [22399]));
Q_ASSIGN U10376 ( .B(clk), .A(\g.we_clk [22398]));
Q_ASSIGN U10377 ( .B(clk), .A(\g.we_clk [22397]));
Q_ASSIGN U10378 ( .B(clk), .A(\g.we_clk [22396]));
Q_ASSIGN U10379 ( .B(clk), .A(\g.we_clk [22395]));
Q_ASSIGN U10380 ( .B(clk), .A(\g.we_clk [22394]));
Q_ASSIGN U10381 ( .B(clk), .A(\g.we_clk [22393]));
Q_ASSIGN U10382 ( .B(clk), .A(\g.we_clk [22392]));
Q_ASSIGN U10383 ( .B(clk), .A(\g.we_clk [22391]));
Q_ASSIGN U10384 ( .B(clk), .A(\g.we_clk [22390]));
Q_ASSIGN U10385 ( .B(clk), .A(\g.we_clk [22389]));
Q_ASSIGN U10386 ( .B(clk), .A(\g.we_clk [22388]));
Q_ASSIGN U10387 ( .B(clk), .A(\g.we_clk [22387]));
Q_ASSIGN U10388 ( .B(clk), .A(\g.we_clk [22386]));
Q_ASSIGN U10389 ( .B(clk), .A(\g.we_clk [22385]));
Q_ASSIGN U10390 ( .B(clk), .A(\g.we_clk [22384]));
Q_ASSIGN U10391 ( .B(clk), .A(\g.we_clk [22383]));
Q_ASSIGN U10392 ( .B(clk), .A(\g.we_clk [22382]));
Q_ASSIGN U10393 ( .B(clk), .A(\g.we_clk [22381]));
Q_ASSIGN U10394 ( .B(clk), .A(\g.we_clk [22380]));
Q_ASSIGN U10395 ( .B(clk), .A(\g.we_clk [22379]));
Q_ASSIGN U10396 ( .B(clk), .A(\g.we_clk [22378]));
Q_ASSIGN U10397 ( .B(clk), .A(\g.we_clk [22377]));
Q_ASSIGN U10398 ( .B(clk), .A(\g.we_clk [22376]));
Q_ASSIGN U10399 ( .B(clk), .A(\g.we_clk [22375]));
Q_ASSIGN U10400 ( .B(clk), .A(\g.we_clk [22374]));
Q_ASSIGN U10401 ( .B(clk), .A(\g.we_clk [22373]));
Q_ASSIGN U10402 ( .B(clk), .A(\g.we_clk [22372]));
Q_ASSIGN U10403 ( .B(clk), .A(\g.we_clk [22371]));
Q_ASSIGN U10404 ( .B(clk), .A(\g.we_clk [22370]));
Q_ASSIGN U10405 ( .B(clk), .A(\g.we_clk [22369]));
Q_ASSIGN U10406 ( .B(clk), .A(\g.we_clk [22368]));
Q_ASSIGN U10407 ( .B(clk), .A(\g.we_clk [22367]));
Q_ASSIGN U10408 ( .B(clk), .A(\g.we_clk [22366]));
Q_ASSIGN U10409 ( .B(clk), .A(\g.we_clk [22365]));
Q_ASSIGN U10410 ( .B(clk), .A(\g.we_clk [22364]));
Q_ASSIGN U10411 ( .B(clk), .A(\g.we_clk [22363]));
Q_ASSIGN U10412 ( .B(clk), .A(\g.we_clk [22362]));
Q_ASSIGN U10413 ( .B(clk), .A(\g.we_clk [22361]));
Q_ASSIGN U10414 ( .B(clk), .A(\g.we_clk [22360]));
Q_ASSIGN U10415 ( .B(clk), .A(\g.we_clk [22359]));
Q_ASSIGN U10416 ( .B(clk), .A(\g.we_clk [22358]));
Q_ASSIGN U10417 ( .B(clk), .A(\g.we_clk [22357]));
Q_ASSIGN U10418 ( .B(clk), .A(\g.we_clk [22356]));
Q_ASSIGN U10419 ( .B(clk), .A(\g.we_clk [22355]));
Q_ASSIGN U10420 ( .B(clk), .A(\g.we_clk [22354]));
Q_ASSIGN U10421 ( .B(clk), .A(\g.we_clk [22353]));
Q_ASSIGN U10422 ( .B(clk), .A(\g.we_clk [22352]));
Q_ASSIGN U10423 ( .B(clk), .A(\g.we_clk [22351]));
Q_ASSIGN U10424 ( .B(clk), .A(\g.we_clk [22350]));
Q_ASSIGN U10425 ( .B(clk), .A(\g.we_clk [22349]));
Q_ASSIGN U10426 ( .B(clk), .A(\g.we_clk [22348]));
Q_ASSIGN U10427 ( .B(clk), .A(\g.we_clk [22347]));
Q_ASSIGN U10428 ( .B(clk), .A(\g.we_clk [22346]));
Q_ASSIGN U10429 ( .B(clk), .A(\g.we_clk [22345]));
Q_ASSIGN U10430 ( .B(clk), .A(\g.we_clk [22344]));
Q_ASSIGN U10431 ( .B(clk), .A(\g.we_clk [22343]));
Q_ASSIGN U10432 ( .B(clk), .A(\g.we_clk [22342]));
Q_ASSIGN U10433 ( .B(clk), .A(\g.we_clk [22341]));
Q_ASSIGN U10434 ( .B(clk), .A(\g.we_clk [22340]));
Q_ASSIGN U10435 ( .B(clk), .A(\g.we_clk [22339]));
Q_ASSIGN U10436 ( .B(clk), .A(\g.we_clk [22338]));
Q_ASSIGN U10437 ( .B(clk), .A(\g.we_clk [22337]));
Q_ASSIGN U10438 ( .B(clk), .A(\g.we_clk [22336]));
Q_ASSIGN U10439 ( .B(clk), .A(\g.we_clk [22335]));
Q_ASSIGN U10440 ( .B(clk), .A(\g.we_clk [22334]));
Q_ASSIGN U10441 ( .B(clk), .A(\g.we_clk [22333]));
Q_ASSIGN U10442 ( .B(clk), .A(\g.we_clk [22332]));
Q_ASSIGN U10443 ( .B(clk), .A(\g.we_clk [22331]));
Q_ASSIGN U10444 ( .B(clk), .A(\g.we_clk [22330]));
Q_ASSIGN U10445 ( .B(clk), .A(\g.we_clk [22329]));
Q_ASSIGN U10446 ( .B(clk), .A(\g.we_clk [22328]));
Q_ASSIGN U10447 ( .B(clk), .A(\g.we_clk [22327]));
Q_ASSIGN U10448 ( .B(clk), .A(\g.we_clk [22326]));
Q_ASSIGN U10449 ( .B(clk), .A(\g.we_clk [22325]));
Q_ASSIGN U10450 ( .B(clk), .A(\g.we_clk [22324]));
Q_ASSIGN U10451 ( .B(clk), .A(\g.we_clk [22323]));
Q_ASSIGN U10452 ( .B(clk), .A(\g.we_clk [22322]));
Q_ASSIGN U10453 ( .B(clk), .A(\g.we_clk [22321]));
Q_ASSIGN U10454 ( .B(clk), .A(\g.we_clk [22320]));
Q_ASSIGN U10455 ( .B(clk), .A(\g.we_clk [22319]));
Q_ASSIGN U10456 ( .B(clk), .A(\g.we_clk [22318]));
Q_ASSIGN U10457 ( .B(clk), .A(\g.we_clk [22317]));
Q_ASSIGN U10458 ( .B(clk), .A(\g.we_clk [22316]));
Q_ASSIGN U10459 ( .B(clk), .A(\g.we_clk [22315]));
Q_ASSIGN U10460 ( .B(clk), .A(\g.we_clk [22314]));
Q_ASSIGN U10461 ( .B(clk), .A(\g.we_clk [22313]));
Q_ASSIGN U10462 ( .B(clk), .A(\g.we_clk [22312]));
Q_ASSIGN U10463 ( .B(clk), .A(\g.we_clk [22311]));
Q_ASSIGN U10464 ( .B(clk), .A(\g.we_clk [22310]));
Q_ASSIGN U10465 ( .B(clk), .A(\g.we_clk [22309]));
Q_ASSIGN U10466 ( .B(clk), .A(\g.we_clk [22308]));
Q_ASSIGN U10467 ( .B(clk), .A(\g.we_clk [22307]));
Q_ASSIGN U10468 ( .B(clk), .A(\g.we_clk [22306]));
Q_ASSIGN U10469 ( .B(clk), .A(\g.we_clk [22305]));
Q_ASSIGN U10470 ( .B(clk), .A(\g.we_clk [22304]));
Q_ASSIGN U10471 ( .B(clk), .A(\g.we_clk [22303]));
Q_ASSIGN U10472 ( .B(clk), .A(\g.we_clk [22302]));
Q_ASSIGN U10473 ( .B(clk), .A(\g.we_clk [22301]));
Q_ASSIGN U10474 ( .B(clk), .A(\g.we_clk [22300]));
Q_ASSIGN U10475 ( .B(clk), .A(\g.we_clk [22299]));
Q_ASSIGN U10476 ( .B(clk), .A(\g.we_clk [22298]));
Q_ASSIGN U10477 ( .B(clk), .A(\g.we_clk [22297]));
Q_ASSIGN U10478 ( .B(clk), .A(\g.we_clk [22296]));
Q_ASSIGN U10479 ( .B(clk), .A(\g.we_clk [22295]));
Q_ASSIGN U10480 ( .B(clk), .A(\g.we_clk [22294]));
Q_ASSIGN U10481 ( .B(clk), .A(\g.we_clk [22293]));
Q_ASSIGN U10482 ( .B(clk), .A(\g.we_clk [22292]));
Q_ASSIGN U10483 ( .B(clk), .A(\g.we_clk [22291]));
Q_ASSIGN U10484 ( .B(clk), .A(\g.we_clk [22290]));
Q_ASSIGN U10485 ( .B(clk), .A(\g.we_clk [22289]));
Q_ASSIGN U10486 ( .B(clk), .A(\g.we_clk [22288]));
Q_ASSIGN U10487 ( .B(clk), .A(\g.we_clk [22287]));
Q_ASSIGN U10488 ( .B(clk), .A(\g.we_clk [22286]));
Q_ASSIGN U10489 ( .B(clk), .A(\g.we_clk [22285]));
Q_ASSIGN U10490 ( .B(clk), .A(\g.we_clk [22284]));
Q_ASSIGN U10491 ( .B(clk), .A(\g.we_clk [22283]));
Q_ASSIGN U10492 ( .B(clk), .A(\g.we_clk [22282]));
Q_ASSIGN U10493 ( .B(clk), .A(\g.we_clk [22281]));
Q_ASSIGN U10494 ( .B(clk), .A(\g.we_clk [22280]));
Q_ASSIGN U10495 ( .B(clk), .A(\g.we_clk [22279]));
Q_ASSIGN U10496 ( .B(clk), .A(\g.we_clk [22278]));
Q_ASSIGN U10497 ( .B(clk), .A(\g.we_clk [22277]));
Q_ASSIGN U10498 ( .B(clk), .A(\g.we_clk [22276]));
Q_ASSIGN U10499 ( .B(clk), .A(\g.we_clk [22275]));
Q_ASSIGN U10500 ( .B(clk), .A(\g.we_clk [22274]));
Q_ASSIGN U10501 ( .B(clk), .A(\g.we_clk [22273]));
Q_ASSIGN U10502 ( .B(clk), .A(\g.we_clk [22272]));
Q_ASSIGN U10503 ( .B(clk), .A(\g.we_clk [22271]));
Q_ASSIGN U10504 ( .B(clk), .A(\g.we_clk [22270]));
Q_ASSIGN U10505 ( .B(clk), .A(\g.we_clk [22269]));
Q_ASSIGN U10506 ( .B(clk), .A(\g.we_clk [22268]));
Q_ASSIGN U10507 ( .B(clk), .A(\g.we_clk [22267]));
Q_ASSIGN U10508 ( .B(clk), .A(\g.we_clk [22266]));
Q_ASSIGN U10509 ( .B(clk), .A(\g.we_clk [22265]));
Q_ASSIGN U10510 ( .B(clk), .A(\g.we_clk [22264]));
Q_ASSIGN U10511 ( .B(clk), .A(\g.we_clk [22263]));
Q_ASSIGN U10512 ( .B(clk), .A(\g.we_clk [22262]));
Q_ASSIGN U10513 ( .B(clk), .A(\g.we_clk [22261]));
Q_ASSIGN U10514 ( .B(clk), .A(\g.we_clk [22260]));
Q_ASSIGN U10515 ( .B(clk), .A(\g.we_clk [22259]));
Q_ASSIGN U10516 ( .B(clk), .A(\g.we_clk [22258]));
Q_ASSIGN U10517 ( .B(clk), .A(\g.we_clk [22257]));
Q_ASSIGN U10518 ( .B(clk), .A(\g.we_clk [22256]));
Q_ASSIGN U10519 ( .B(clk), .A(\g.we_clk [22255]));
Q_ASSIGN U10520 ( .B(clk), .A(\g.we_clk [22254]));
Q_ASSIGN U10521 ( .B(clk), .A(\g.we_clk [22253]));
Q_ASSIGN U10522 ( .B(clk), .A(\g.we_clk [22252]));
Q_ASSIGN U10523 ( .B(clk), .A(\g.we_clk [22251]));
Q_ASSIGN U10524 ( .B(clk), .A(\g.we_clk [22250]));
Q_ASSIGN U10525 ( .B(clk), .A(\g.we_clk [22249]));
Q_ASSIGN U10526 ( .B(clk), .A(\g.we_clk [22248]));
Q_ASSIGN U10527 ( .B(clk), .A(\g.we_clk [22247]));
Q_ASSIGN U10528 ( .B(clk), .A(\g.we_clk [22246]));
Q_ASSIGN U10529 ( .B(clk), .A(\g.we_clk [22245]));
Q_ASSIGN U10530 ( .B(clk), .A(\g.we_clk [22244]));
Q_ASSIGN U10531 ( .B(clk), .A(\g.we_clk [22243]));
Q_ASSIGN U10532 ( .B(clk), .A(\g.we_clk [22242]));
Q_ASSIGN U10533 ( .B(clk), .A(\g.we_clk [22241]));
Q_ASSIGN U10534 ( .B(clk), .A(\g.we_clk [22240]));
Q_ASSIGN U10535 ( .B(clk), .A(\g.we_clk [22239]));
Q_ASSIGN U10536 ( .B(clk), .A(\g.we_clk [22238]));
Q_ASSIGN U10537 ( .B(clk), .A(\g.we_clk [22237]));
Q_ASSIGN U10538 ( .B(clk), .A(\g.we_clk [22236]));
Q_ASSIGN U10539 ( .B(clk), .A(\g.we_clk [22235]));
Q_ASSIGN U10540 ( .B(clk), .A(\g.we_clk [22234]));
Q_ASSIGN U10541 ( .B(clk), .A(\g.we_clk [22233]));
Q_ASSIGN U10542 ( .B(clk), .A(\g.we_clk [22232]));
Q_ASSIGN U10543 ( .B(clk), .A(\g.we_clk [22231]));
Q_ASSIGN U10544 ( .B(clk), .A(\g.we_clk [22230]));
Q_ASSIGN U10545 ( .B(clk), .A(\g.we_clk [22229]));
Q_ASSIGN U10546 ( .B(clk), .A(\g.we_clk [22228]));
Q_ASSIGN U10547 ( .B(clk), .A(\g.we_clk [22227]));
Q_ASSIGN U10548 ( .B(clk), .A(\g.we_clk [22226]));
Q_ASSIGN U10549 ( .B(clk), .A(\g.we_clk [22225]));
Q_ASSIGN U10550 ( .B(clk), .A(\g.we_clk [22224]));
Q_ASSIGN U10551 ( .B(clk), .A(\g.we_clk [22223]));
Q_ASSIGN U10552 ( .B(clk), .A(\g.we_clk [22222]));
Q_ASSIGN U10553 ( .B(clk), .A(\g.we_clk [22221]));
Q_ASSIGN U10554 ( .B(clk), .A(\g.we_clk [22220]));
Q_ASSIGN U10555 ( .B(clk), .A(\g.we_clk [22219]));
Q_ASSIGN U10556 ( .B(clk), .A(\g.we_clk [22218]));
Q_ASSIGN U10557 ( .B(clk), .A(\g.we_clk [22217]));
Q_ASSIGN U10558 ( .B(clk), .A(\g.we_clk [22216]));
Q_ASSIGN U10559 ( .B(clk), .A(\g.we_clk [22215]));
Q_ASSIGN U10560 ( .B(clk), .A(\g.we_clk [22214]));
Q_ASSIGN U10561 ( .B(clk), .A(\g.we_clk [22213]));
Q_ASSIGN U10562 ( .B(clk), .A(\g.we_clk [22212]));
Q_ASSIGN U10563 ( .B(clk), .A(\g.we_clk [22211]));
Q_ASSIGN U10564 ( .B(clk), .A(\g.we_clk [22210]));
Q_ASSIGN U10565 ( .B(clk), .A(\g.we_clk [22209]));
Q_ASSIGN U10566 ( .B(clk), .A(\g.we_clk [22208]));
Q_ASSIGN U10567 ( .B(clk), .A(\g.we_clk [22207]));
Q_ASSIGN U10568 ( .B(clk), .A(\g.we_clk [22206]));
Q_ASSIGN U10569 ( .B(clk), .A(\g.we_clk [22205]));
Q_ASSIGN U10570 ( .B(clk), .A(\g.we_clk [22204]));
Q_ASSIGN U10571 ( .B(clk), .A(\g.we_clk [22203]));
Q_ASSIGN U10572 ( .B(clk), .A(\g.we_clk [22202]));
Q_ASSIGN U10573 ( .B(clk), .A(\g.we_clk [22201]));
Q_ASSIGN U10574 ( .B(clk), .A(\g.we_clk [22200]));
Q_ASSIGN U10575 ( .B(clk), .A(\g.we_clk [22199]));
Q_ASSIGN U10576 ( .B(clk), .A(\g.we_clk [22198]));
Q_ASSIGN U10577 ( .B(clk), .A(\g.we_clk [22197]));
Q_ASSIGN U10578 ( .B(clk), .A(\g.we_clk [22196]));
Q_ASSIGN U10579 ( .B(clk), .A(\g.we_clk [22195]));
Q_ASSIGN U10580 ( .B(clk), .A(\g.we_clk [22194]));
Q_ASSIGN U10581 ( .B(clk), .A(\g.we_clk [22193]));
Q_ASSIGN U10582 ( .B(clk), .A(\g.we_clk [22192]));
Q_ASSIGN U10583 ( .B(clk), .A(\g.we_clk [22191]));
Q_ASSIGN U10584 ( .B(clk), .A(\g.we_clk [22190]));
Q_ASSIGN U10585 ( .B(clk), .A(\g.we_clk [22189]));
Q_ASSIGN U10586 ( .B(clk), .A(\g.we_clk [22188]));
Q_ASSIGN U10587 ( .B(clk), .A(\g.we_clk [22187]));
Q_ASSIGN U10588 ( .B(clk), .A(\g.we_clk [22186]));
Q_ASSIGN U10589 ( .B(clk), .A(\g.we_clk [22185]));
Q_ASSIGN U10590 ( .B(clk), .A(\g.we_clk [22184]));
Q_ASSIGN U10591 ( .B(clk), .A(\g.we_clk [22183]));
Q_ASSIGN U10592 ( .B(clk), .A(\g.we_clk [22182]));
Q_ASSIGN U10593 ( .B(clk), .A(\g.we_clk [22181]));
Q_ASSIGN U10594 ( .B(clk), .A(\g.we_clk [22180]));
Q_ASSIGN U10595 ( .B(clk), .A(\g.we_clk [22179]));
Q_ASSIGN U10596 ( .B(clk), .A(\g.we_clk [22178]));
Q_ASSIGN U10597 ( .B(clk), .A(\g.we_clk [22177]));
Q_ASSIGN U10598 ( .B(clk), .A(\g.we_clk [22176]));
Q_ASSIGN U10599 ( .B(clk), .A(\g.we_clk [22175]));
Q_ASSIGN U10600 ( .B(clk), .A(\g.we_clk [22174]));
Q_ASSIGN U10601 ( .B(clk), .A(\g.we_clk [22173]));
Q_ASSIGN U10602 ( .B(clk), .A(\g.we_clk [22172]));
Q_ASSIGN U10603 ( .B(clk), .A(\g.we_clk [22171]));
Q_ASSIGN U10604 ( .B(clk), .A(\g.we_clk [22170]));
Q_ASSIGN U10605 ( .B(clk), .A(\g.we_clk [22169]));
Q_ASSIGN U10606 ( .B(clk), .A(\g.we_clk [22168]));
Q_ASSIGN U10607 ( .B(clk), .A(\g.we_clk [22167]));
Q_ASSIGN U10608 ( .B(clk), .A(\g.we_clk [22166]));
Q_ASSIGN U10609 ( .B(clk), .A(\g.we_clk [22165]));
Q_ASSIGN U10610 ( .B(clk), .A(\g.we_clk [22164]));
Q_ASSIGN U10611 ( .B(clk), .A(\g.we_clk [22163]));
Q_ASSIGN U10612 ( .B(clk), .A(\g.we_clk [22162]));
Q_ASSIGN U10613 ( .B(clk), .A(\g.we_clk [22161]));
Q_ASSIGN U10614 ( .B(clk), .A(\g.we_clk [22160]));
Q_ASSIGN U10615 ( .B(clk), .A(\g.we_clk [22159]));
Q_ASSIGN U10616 ( .B(clk), .A(\g.we_clk [22158]));
Q_ASSIGN U10617 ( .B(clk), .A(\g.we_clk [22157]));
Q_ASSIGN U10618 ( .B(clk), .A(\g.we_clk [22156]));
Q_ASSIGN U10619 ( .B(clk), .A(\g.we_clk [22155]));
Q_ASSIGN U10620 ( .B(clk), .A(\g.we_clk [22154]));
Q_ASSIGN U10621 ( .B(clk), .A(\g.we_clk [22153]));
Q_ASSIGN U10622 ( .B(clk), .A(\g.we_clk [22152]));
Q_ASSIGN U10623 ( .B(clk), .A(\g.we_clk [22151]));
Q_ASSIGN U10624 ( .B(clk), .A(\g.we_clk [22150]));
Q_ASSIGN U10625 ( .B(clk), .A(\g.we_clk [22149]));
Q_ASSIGN U10626 ( .B(clk), .A(\g.we_clk [22148]));
Q_ASSIGN U10627 ( .B(clk), .A(\g.we_clk [22147]));
Q_ASSIGN U10628 ( .B(clk), .A(\g.we_clk [22146]));
Q_ASSIGN U10629 ( .B(clk), .A(\g.we_clk [22145]));
Q_ASSIGN U10630 ( .B(clk), .A(\g.we_clk [22144]));
Q_ASSIGN U10631 ( .B(clk), .A(\g.we_clk [22143]));
Q_ASSIGN U10632 ( .B(clk), .A(\g.we_clk [22142]));
Q_ASSIGN U10633 ( .B(clk), .A(\g.we_clk [22141]));
Q_ASSIGN U10634 ( .B(clk), .A(\g.we_clk [22140]));
Q_ASSIGN U10635 ( .B(clk), .A(\g.we_clk [22139]));
Q_ASSIGN U10636 ( .B(clk), .A(\g.we_clk [22138]));
Q_ASSIGN U10637 ( .B(clk), .A(\g.we_clk [22137]));
Q_ASSIGN U10638 ( .B(clk), .A(\g.we_clk [22136]));
Q_ASSIGN U10639 ( .B(clk), .A(\g.we_clk [22135]));
Q_ASSIGN U10640 ( .B(clk), .A(\g.we_clk [22134]));
Q_ASSIGN U10641 ( .B(clk), .A(\g.we_clk [22133]));
Q_ASSIGN U10642 ( .B(clk), .A(\g.we_clk [22132]));
Q_ASSIGN U10643 ( .B(clk), .A(\g.we_clk [22131]));
Q_ASSIGN U10644 ( .B(clk), .A(\g.we_clk [22130]));
Q_ASSIGN U10645 ( .B(clk), .A(\g.we_clk [22129]));
Q_ASSIGN U10646 ( .B(clk), .A(\g.we_clk [22128]));
Q_ASSIGN U10647 ( .B(clk), .A(\g.we_clk [22127]));
Q_ASSIGN U10648 ( .B(clk), .A(\g.we_clk [22126]));
Q_ASSIGN U10649 ( .B(clk), .A(\g.we_clk [22125]));
Q_ASSIGN U10650 ( .B(clk), .A(\g.we_clk [22124]));
Q_ASSIGN U10651 ( .B(clk), .A(\g.we_clk [22123]));
Q_ASSIGN U10652 ( .B(clk), .A(\g.we_clk [22122]));
Q_ASSIGN U10653 ( .B(clk), .A(\g.we_clk [22121]));
Q_ASSIGN U10654 ( .B(clk), .A(\g.we_clk [22120]));
Q_ASSIGN U10655 ( .B(clk), .A(\g.we_clk [22119]));
Q_ASSIGN U10656 ( .B(clk), .A(\g.we_clk [22118]));
Q_ASSIGN U10657 ( .B(clk), .A(\g.we_clk [22117]));
Q_ASSIGN U10658 ( .B(clk), .A(\g.we_clk [22116]));
Q_ASSIGN U10659 ( .B(clk), .A(\g.we_clk [22115]));
Q_ASSIGN U10660 ( .B(clk), .A(\g.we_clk [22114]));
Q_ASSIGN U10661 ( .B(clk), .A(\g.we_clk [22113]));
Q_ASSIGN U10662 ( .B(clk), .A(\g.we_clk [22112]));
Q_ASSIGN U10663 ( .B(clk), .A(\g.we_clk [22111]));
Q_ASSIGN U10664 ( .B(clk), .A(\g.we_clk [22110]));
Q_ASSIGN U10665 ( .B(clk), .A(\g.we_clk [22109]));
Q_ASSIGN U10666 ( .B(clk), .A(\g.we_clk [22108]));
Q_ASSIGN U10667 ( .B(clk), .A(\g.we_clk [22107]));
Q_ASSIGN U10668 ( .B(clk), .A(\g.we_clk [22106]));
Q_ASSIGN U10669 ( .B(clk), .A(\g.we_clk [22105]));
Q_ASSIGN U10670 ( .B(clk), .A(\g.we_clk [22104]));
Q_ASSIGN U10671 ( .B(clk), .A(\g.we_clk [22103]));
Q_ASSIGN U10672 ( .B(clk), .A(\g.we_clk [22102]));
Q_ASSIGN U10673 ( .B(clk), .A(\g.we_clk [22101]));
Q_ASSIGN U10674 ( .B(clk), .A(\g.we_clk [22100]));
Q_ASSIGN U10675 ( .B(clk), .A(\g.we_clk [22099]));
Q_ASSIGN U10676 ( .B(clk), .A(\g.we_clk [22098]));
Q_ASSIGN U10677 ( .B(clk), .A(\g.we_clk [22097]));
Q_ASSIGN U10678 ( .B(clk), .A(\g.we_clk [22096]));
Q_ASSIGN U10679 ( .B(clk), .A(\g.we_clk [22095]));
Q_ASSIGN U10680 ( .B(clk), .A(\g.we_clk [22094]));
Q_ASSIGN U10681 ( .B(clk), .A(\g.we_clk [22093]));
Q_ASSIGN U10682 ( .B(clk), .A(\g.we_clk [22092]));
Q_ASSIGN U10683 ( .B(clk), .A(\g.we_clk [22091]));
Q_ASSIGN U10684 ( .B(clk), .A(\g.we_clk [22090]));
Q_ASSIGN U10685 ( .B(clk), .A(\g.we_clk [22089]));
Q_ASSIGN U10686 ( .B(clk), .A(\g.we_clk [22088]));
Q_ASSIGN U10687 ( .B(clk), .A(\g.we_clk [22087]));
Q_ASSIGN U10688 ( .B(clk), .A(\g.we_clk [22086]));
Q_ASSIGN U10689 ( .B(clk), .A(\g.we_clk [22085]));
Q_ASSIGN U10690 ( .B(clk), .A(\g.we_clk [22084]));
Q_ASSIGN U10691 ( .B(clk), .A(\g.we_clk [22083]));
Q_ASSIGN U10692 ( .B(clk), .A(\g.we_clk [22082]));
Q_ASSIGN U10693 ( .B(clk), .A(\g.we_clk [22081]));
Q_ASSIGN U10694 ( .B(clk), .A(\g.we_clk [22080]));
Q_ASSIGN U10695 ( .B(clk), .A(\g.we_clk [22079]));
Q_ASSIGN U10696 ( .B(clk), .A(\g.we_clk [22078]));
Q_ASSIGN U10697 ( .B(clk), .A(\g.we_clk [22077]));
Q_ASSIGN U10698 ( .B(clk), .A(\g.we_clk [22076]));
Q_ASSIGN U10699 ( .B(clk), .A(\g.we_clk [22075]));
Q_ASSIGN U10700 ( .B(clk), .A(\g.we_clk [22074]));
Q_ASSIGN U10701 ( .B(clk), .A(\g.we_clk [22073]));
Q_ASSIGN U10702 ( .B(clk), .A(\g.we_clk [22072]));
Q_ASSIGN U10703 ( .B(clk), .A(\g.we_clk [22071]));
Q_ASSIGN U10704 ( .B(clk), .A(\g.we_clk [22070]));
Q_ASSIGN U10705 ( .B(clk), .A(\g.we_clk [22069]));
Q_ASSIGN U10706 ( .B(clk), .A(\g.we_clk [22068]));
Q_ASSIGN U10707 ( .B(clk), .A(\g.we_clk [22067]));
Q_ASSIGN U10708 ( .B(clk), .A(\g.we_clk [22066]));
Q_ASSIGN U10709 ( .B(clk), .A(\g.we_clk [22065]));
Q_ASSIGN U10710 ( .B(clk), .A(\g.we_clk [22064]));
Q_ASSIGN U10711 ( .B(clk), .A(\g.we_clk [22063]));
Q_ASSIGN U10712 ( .B(clk), .A(\g.we_clk [22062]));
Q_ASSIGN U10713 ( .B(clk), .A(\g.we_clk [22061]));
Q_ASSIGN U10714 ( .B(clk), .A(\g.we_clk [22060]));
Q_ASSIGN U10715 ( .B(clk), .A(\g.we_clk [22059]));
Q_ASSIGN U10716 ( .B(clk), .A(\g.we_clk [22058]));
Q_ASSIGN U10717 ( .B(clk), .A(\g.we_clk [22057]));
Q_ASSIGN U10718 ( .B(clk), .A(\g.we_clk [22056]));
Q_ASSIGN U10719 ( .B(clk), .A(\g.we_clk [22055]));
Q_ASSIGN U10720 ( .B(clk), .A(\g.we_clk [22054]));
Q_ASSIGN U10721 ( .B(clk), .A(\g.we_clk [22053]));
Q_ASSIGN U10722 ( .B(clk), .A(\g.we_clk [22052]));
Q_ASSIGN U10723 ( .B(clk), .A(\g.we_clk [22051]));
Q_ASSIGN U10724 ( .B(clk), .A(\g.we_clk [22050]));
Q_ASSIGN U10725 ( .B(clk), .A(\g.we_clk [22049]));
Q_ASSIGN U10726 ( .B(clk), .A(\g.we_clk [22048]));
Q_ASSIGN U10727 ( .B(clk), .A(\g.we_clk [22047]));
Q_ASSIGN U10728 ( .B(clk), .A(\g.we_clk [22046]));
Q_ASSIGN U10729 ( .B(clk), .A(\g.we_clk [22045]));
Q_ASSIGN U10730 ( .B(clk), .A(\g.we_clk [22044]));
Q_ASSIGN U10731 ( .B(clk), .A(\g.we_clk [22043]));
Q_ASSIGN U10732 ( .B(clk), .A(\g.we_clk [22042]));
Q_ASSIGN U10733 ( .B(clk), .A(\g.we_clk [22041]));
Q_ASSIGN U10734 ( .B(clk), .A(\g.we_clk [22040]));
Q_ASSIGN U10735 ( .B(clk), .A(\g.we_clk [22039]));
Q_ASSIGN U10736 ( .B(clk), .A(\g.we_clk [22038]));
Q_ASSIGN U10737 ( .B(clk), .A(\g.we_clk [22037]));
Q_ASSIGN U10738 ( .B(clk), .A(\g.we_clk [22036]));
Q_ASSIGN U10739 ( .B(clk), .A(\g.we_clk [22035]));
Q_ASSIGN U10740 ( .B(clk), .A(\g.we_clk [22034]));
Q_ASSIGN U10741 ( .B(clk), .A(\g.we_clk [22033]));
Q_ASSIGN U10742 ( .B(clk), .A(\g.we_clk [22032]));
Q_ASSIGN U10743 ( .B(clk), .A(\g.we_clk [22031]));
Q_ASSIGN U10744 ( .B(clk), .A(\g.we_clk [22030]));
Q_ASSIGN U10745 ( .B(clk), .A(\g.we_clk [22029]));
Q_ASSIGN U10746 ( .B(clk), .A(\g.we_clk [22028]));
Q_ASSIGN U10747 ( .B(clk), .A(\g.we_clk [22027]));
Q_ASSIGN U10748 ( .B(clk), .A(\g.we_clk [22026]));
Q_ASSIGN U10749 ( .B(clk), .A(\g.we_clk [22025]));
Q_ASSIGN U10750 ( .B(clk), .A(\g.we_clk [22024]));
Q_ASSIGN U10751 ( .B(clk), .A(\g.we_clk [22023]));
Q_ASSIGN U10752 ( .B(clk), .A(\g.we_clk [22022]));
Q_ASSIGN U10753 ( .B(clk), .A(\g.we_clk [22021]));
Q_ASSIGN U10754 ( .B(clk), .A(\g.we_clk [22020]));
Q_ASSIGN U10755 ( .B(clk), .A(\g.we_clk [22019]));
Q_ASSIGN U10756 ( .B(clk), .A(\g.we_clk [22018]));
Q_ASSIGN U10757 ( .B(clk), .A(\g.we_clk [22017]));
Q_ASSIGN U10758 ( .B(clk), .A(\g.we_clk [22016]));
Q_ASSIGN U10759 ( .B(clk), .A(\g.we_clk [22015]));
Q_ASSIGN U10760 ( .B(clk), .A(\g.we_clk [22014]));
Q_ASSIGN U10761 ( .B(clk), .A(\g.we_clk [22013]));
Q_ASSIGN U10762 ( .B(clk), .A(\g.we_clk [22012]));
Q_ASSIGN U10763 ( .B(clk), .A(\g.we_clk [22011]));
Q_ASSIGN U10764 ( .B(clk), .A(\g.we_clk [22010]));
Q_ASSIGN U10765 ( .B(clk), .A(\g.we_clk [22009]));
Q_ASSIGN U10766 ( .B(clk), .A(\g.we_clk [22008]));
Q_ASSIGN U10767 ( .B(clk), .A(\g.we_clk [22007]));
Q_ASSIGN U10768 ( .B(clk), .A(\g.we_clk [22006]));
Q_ASSIGN U10769 ( .B(clk), .A(\g.we_clk [22005]));
Q_ASSIGN U10770 ( .B(clk), .A(\g.we_clk [22004]));
Q_ASSIGN U10771 ( .B(clk), .A(\g.we_clk [22003]));
Q_ASSIGN U10772 ( .B(clk), .A(\g.we_clk [22002]));
Q_ASSIGN U10773 ( .B(clk), .A(\g.we_clk [22001]));
Q_ASSIGN U10774 ( .B(clk), .A(\g.we_clk [22000]));
Q_ASSIGN U10775 ( .B(clk), .A(\g.we_clk [21999]));
Q_ASSIGN U10776 ( .B(clk), .A(\g.we_clk [21998]));
Q_ASSIGN U10777 ( .B(clk), .A(\g.we_clk [21997]));
Q_ASSIGN U10778 ( .B(clk), .A(\g.we_clk [21996]));
Q_ASSIGN U10779 ( .B(clk), .A(\g.we_clk [21995]));
Q_ASSIGN U10780 ( .B(clk), .A(\g.we_clk [21994]));
Q_ASSIGN U10781 ( .B(clk), .A(\g.we_clk [21993]));
Q_ASSIGN U10782 ( .B(clk), .A(\g.we_clk [21992]));
Q_ASSIGN U10783 ( .B(clk), .A(\g.we_clk [21991]));
Q_ASSIGN U10784 ( .B(clk), .A(\g.we_clk [21990]));
Q_ASSIGN U10785 ( .B(clk), .A(\g.we_clk [21989]));
Q_ASSIGN U10786 ( .B(clk), .A(\g.we_clk [21988]));
Q_ASSIGN U10787 ( .B(clk), .A(\g.we_clk [21987]));
Q_ASSIGN U10788 ( .B(clk), .A(\g.we_clk [21986]));
Q_ASSIGN U10789 ( .B(clk), .A(\g.we_clk [21985]));
Q_ASSIGN U10790 ( .B(clk), .A(\g.we_clk [21984]));
Q_ASSIGN U10791 ( .B(clk), .A(\g.we_clk [21983]));
Q_ASSIGN U10792 ( .B(clk), .A(\g.we_clk [21982]));
Q_ASSIGN U10793 ( .B(clk), .A(\g.we_clk [21981]));
Q_ASSIGN U10794 ( .B(clk), .A(\g.we_clk [21980]));
Q_ASSIGN U10795 ( .B(clk), .A(\g.we_clk [21979]));
Q_ASSIGN U10796 ( .B(clk), .A(\g.we_clk [21978]));
Q_ASSIGN U10797 ( .B(clk), .A(\g.we_clk [21977]));
Q_ASSIGN U10798 ( .B(clk), .A(\g.we_clk [21976]));
Q_ASSIGN U10799 ( .B(clk), .A(\g.we_clk [21975]));
Q_ASSIGN U10800 ( .B(clk), .A(\g.we_clk [21974]));
Q_ASSIGN U10801 ( .B(clk), .A(\g.we_clk [21973]));
Q_ASSIGN U10802 ( .B(clk), .A(\g.we_clk [21972]));
Q_ASSIGN U10803 ( .B(clk), .A(\g.we_clk [21971]));
Q_ASSIGN U10804 ( .B(clk), .A(\g.we_clk [21970]));
Q_ASSIGN U10805 ( .B(clk), .A(\g.we_clk [21969]));
Q_ASSIGN U10806 ( .B(clk), .A(\g.we_clk [21968]));
Q_ASSIGN U10807 ( .B(clk), .A(\g.we_clk [21967]));
Q_ASSIGN U10808 ( .B(clk), .A(\g.we_clk [21966]));
Q_ASSIGN U10809 ( .B(clk), .A(\g.we_clk [21965]));
Q_ASSIGN U10810 ( .B(clk), .A(\g.we_clk [21964]));
Q_ASSIGN U10811 ( .B(clk), .A(\g.we_clk [21963]));
Q_ASSIGN U10812 ( .B(clk), .A(\g.we_clk [21962]));
Q_ASSIGN U10813 ( .B(clk), .A(\g.we_clk [21961]));
Q_ASSIGN U10814 ( .B(clk), .A(\g.we_clk [21960]));
Q_ASSIGN U10815 ( .B(clk), .A(\g.we_clk [21959]));
Q_ASSIGN U10816 ( .B(clk), .A(\g.we_clk [21958]));
Q_ASSIGN U10817 ( .B(clk), .A(\g.we_clk [21957]));
Q_ASSIGN U10818 ( .B(clk), .A(\g.we_clk [21956]));
Q_ASSIGN U10819 ( .B(clk), .A(\g.we_clk [21955]));
Q_ASSIGN U10820 ( .B(clk), .A(\g.we_clk [21954]));
Q_ASSIGN U10821 ( .B(clk), .A(\g.we_clk [21953]));
Q_ASSIGN U10822 ( .B(clk), .A(\g.we_clk [21952]));
Q_ASSIGN U10823 ( .B(clk), .A(\g.we_clk [21951]));
Q_ASSIGN U10824 ( .B(clk), .A(\g.we_clk [21950]));
Q_ASSIGN U10825 ( .B(clk), .A(\g.we_clk [21949]));
Q_ASSIGN U10826 ( .B(clk), .A(\g.we_clk [21948]));
Q_ASSIGN U10827 ( .B(clk), .A(\g.we_clk [21947]));
Q_ASSIGN U10828 ( .B(clk), .A(\g.we_clk [21946]));
Q_ASSIGN U10829 ( .B(clk), .A(\g.we_clk [21945]));
Q_ASSIGN U10830 ( .B(clk), .A(\g.we_clk [21944]));
Q_ASSIGN U10831 ( .B(clk), .A(\g.we_clk [21943]));
Q_ASSIGN U10832 ( .B(clk), .A(\g.we_clk [21942]));
Q_ASSIGN U10833 ( .B(clk), .A(\g.we_clk [21941]));
Q_ASSIGN U10834 ( .B(clk), .A(\g.we_clk [21940]));
Q_ASSIGN U10835 ( .B(clk), .A(\g.we_clk [21939]));
Q_ASSIGN U10836 ( .B(clk), .A(\g.we_clk [21938]));
Q_ASSIGN U10837 ( .B(clk), .A(\g.we_clk [21937]));
Q_ASSIGN U10838 ( .B(clk), .A(\g.we_clk [21936]));
Q_ASSIGN U10839 ( .B(clk), .A(\g.we_clk [21935]));
Q_ASSIGN U10840 ( .B(clk), .A(\g.we_clk [21934]));
Q_ASSIGN U10841 ( .B(clk), .A(\g.we_clk [21933]));
Q_ASSIGN U10842 ( .B(clk), .A(\g.we_clk [21932]));
Q_ASSIGN U10843 ( .B(clk), .A(\g.we_clk [21931]));
Q_ASSIGN U10844 ( .B(clk), .A(\g.we_clk [21930]));
Q_ASSIGN U10845 ( .B(clk), .A(\g.we_clk [21929]));
Q_ASSIGN U10846 ( .B(clk), .A(\g.we_clk [21928]));
Q_ASSIGN U10847 ( .B(clk), .A(\g.we_clk [21927]));
Q_ASSIGN U10848 ( .B(clk), .A(\g.we_clk [21926]));
Q_ASSIGN U10849 ( .B(clk), .A(\g.we_clk [21925]));
Q_ASSIGN U10850 ( .B(clk), .A(\g.we_clk [21924]));
Q_ASSIGN U10851 ( .B(clk), .A(\g.we_clk [21923]));
Q_ASSIGN U10852 ( .B(clk), .A(\g.we_clk [21922]));
Q_ASSIGN U10853 ( .B(clk), .A(\g.we_clk [21921]));
Q_ASSIGN U10854 ( .B(clk), .A(\g.we_clk [21920]));
Q_ASSIGN U10855 ( .B(clk), .A(\g.we_clk [21919]));
Q_ASSIGN U10856 ( .B(clk), .A(\g.we_clk [21918]));
Q_ASSIGN U10857 ( .B(clk), .A(\g.we_clk [21917]));
Q_ASSIGN U10858 ( .B(clk), .A(\g.we_clk [21916]));
Q_ASSIGN U10859 ( .B(clk), .A(\g.we_clk [21915]));
Q_ASSIGN U10860 ( .B(clk), .A(\g.we_clk [21914]));
Q_ASSIGN U10861 ( .B(clk), .A(\g.we_clk [21913]));
Q_ASSIGN U10862 ( .B(clk), .A(\g.we_clk [21912]));
Q_ASSIGN U10863 ( .B(clk), .A(\g.we_clk [21911]));
Q_ASSIGN U10864 ( .B(clk), .A(\g.we_clk [21910]));
Q_ASSIGN U10865 ( .B(clk), .A(\g.we_clk [21909]));
Q_ASSIGN U10866 ( .B(clk), .A(\g.we_clk [21908]));
Q_ASSIGN U10867 ( .B(clk), .A(\g.we_clk [21907]));
Q_ASSIGN U10868 ( .B(clk), .A(\g.we_clk [21906]));
Q_ASSIGN U10869 ( .B(clk), .A(\g.we_clk [21905]));
Q_ASSIGN U10870 ( .B(clk), .A(\g.we_clk [21904]));
Q_ASSIGN U10871 ( .B(clk), .A(\g.we_clk [21903]));
Q_ASSIGN U10872 ( .B(clk), .A(\g.we_clk [21902]));
Q_ASSIGN U10873 ( .B(clk), .A(\g.we_clk [21901]));
Q_ASSIGN U10874 ( .B(clk), .A(\g.we_clk [21900]));
Q_ASSIGN U10875 ( .B(clk), .A(\g.we_clk [21899]));
Q_ASSIGN U10876 ( .B(clk), .A(\g.we_clk [21898]));
Q_ASSIGN U10877 ( .B(clk), .A(\g.we_clk [21897]));
Q_ASSIGN U10878 ( .B(clk), .A(\g.we_clk [21896]));
Q_ASSIGN U10879 ( .B(clk), .A(\g.we_clk [21895]));
Q_ASSIGN U10880 ( .B(clk), .A(\g.we_clk [21894]));
Q_ASSIGN U10881 ( .B(clk), .A(\g.we_clk [21893]));
Q_ASSIGN U10882 ( .B(clk), .A(\g.we_clk [21892]));
Q_ASSIGN U10883 ( .B(clk), .A(\g.we_clk [21891]));
Q_ASSIGN U10884 ( .B(clk), .A(\g.we_clk [21890]));
Q_ASSIGN U10885 ( .B(clk), .A(\g.we_clk [21889]));
Q_ASSIGN U10886 ( .B(clk), .A(\g.we_clk [21888]));
Q_ASSIGN U10887 ( .B(clk), .A(\g.we_clk [21887]));
Q_ASSIGN U10888 ( .B(clk), .A(\g.we_clk [21886]));
Q_ASSIGN U10889 ( .B(clk), .A(\g.we_clk [21885]));
Q_ASSIGN U10890 ( .B(clk), .A(\g.we_clk [21884]));
Q_ASSIGN U10891 ( .B(clk), .A(\g.we_clk [21883]));
Q_ASSIGN U10892 ( .B(clk), .A(\g.we_clk [21882]));
Q_ASSIGN U10893 ( .B(clk), .A(\g.we_clk [21881]));
Q_ASSIGN U10894 ( .B(clk), .A(\g.we_clk [21880]));
Q_ASSIGN U10895 ( .B(clk), .A(\g.we_clk [21879]));
Q_ASSIGN U10896 ( .B(clk), .A(\g.we_clk [21878]));
Q_ASSIGN U10897 ( .B(clk), .A(\g.we_clk [21877]));
Q_ASSIGN U10898 ( .B(clk), .A(\g.we_clk [21876]));
Q_ASSIGN U10899 ( .B(clk), .A(\g.we_clk [21875]));
Q_ASSIGN U10900 ( .B(clk), .A(\g.we_clk [21874]));
Q_ASSIGN U10901 ( .B(clk), .A(\g.we_clk [21873]));
Q_ASSIGN U10902 ( .B(clk), .A(\g.we_clk [21872]));
Q_ASSIGN U10903 ( .B(clk), .A(\g.we_clk [21871]));
Q_ASSIGN U10904 ( .B(clk), .A(\g.we_clk [21870]));
Q_ASSIGN U10905 ( .B(clk), .A(\g.we_clk [21869]));
Q_ASSIGN U10906 ( .B(clk), .A(\g.we_clk [21868]));
Q_ASSIGN U10907 ( .B(clk), .A(\g.we_clk [21867]));
Q_ASSIGN U10908 ( .B(clk), .A(\g.we_clk [21866]));
Q_ASSIGN U10909 ( .B(clk), .A(\g.we_clk [21865]));
Q_ASSIGN U10910 ( .B(clk), .A(\g.we_clk [21864]));
Q_ASSIGN U10911 ( .B(clk), .A(\g.we_clk [21863]));
Q_ASSIGN U10912 ( .B(clk), .A(\g.we_clk [21862]));
Q_ASSIGN U10913 ( .B(clk), .A(\g.we_clk [21861]));
Q_ASSIGN U10914 ( .B(clk), .A(\g.we_clk [21860]));
Q_ASSIGN U10915 ( .B(clk), .A(\g.we_clk [21859]));
Q_ASSIGN U10916 ( .B(clk), .A(\g.we_clk [21858]));
Q_ASSIGN U10917 ( .B(clk), .A(\g.we_clk [21857]));
Q_ASSIGN U10918 ( .B(clk), .A(\g.we_clk [21856]));
Q_ASSIGN U10919 ( .B(clk), .A(\g.we_clk [21855]));
Q_ASSIGN U10920 ( .B(clk), .A(\g.we_clk [21854]));
Q_ASSIGN U10921 ( .B(clk), .A(\g.we_clk [21853]));
Q_ASSIGN U10922 ( .B(clk), .A(\g.we_clk [21852]));
Q_ASSIGN U10923 ( .B(clk), .A(\g.we_clk [21851]));
Q_ASSIGN U10924 ( .B(clk), .A(\g.we_clk [21850]));
Q_ASSIGN U10925 ( .B(clk), .A(\g.we_clk [21849]));
Q_ASSIGN U10926 ( .B(clk), .A(\g.we_clk [21848]));
Q_ASSIGN U10927 ( .B(clk), .A(\g.we_clk [21847]));
Q_ASSIGN U10928 ( .B(clk), .A(\g.we_clk [21846]));
Q_ASSIGN U10929 ( .B(clk), .A(\g.we_clk [21845]));
Q_ASSIGN U10930 ( .B(clk), .A(\g.we_clk [21844]));
Q_ASSIGN U10931 ( .B(clk), .A(\g.we_clk [21843]));
Q_ASSIGN U10932 ( .B(clk), .A(\g.we_clk [21842]));
Q_ASSIGN U10933 ( .B(clk), .A(\g.we_clk [21841]));
Q_ASSIGN U10934 ( .B(clk), .A(\g.we_clk [21840]));
Q_ASSIGN U10935 ( .B(clk), .A(\g.we_clk [21839]));
Q_ASSIGN U10936 ( .B(clk), .A(\g.we_clk [21838]));
Q_ASSIGN U10937 ( .B(clk), .A(\g.we_clk [21837]));
Q_ASSIGN U10938 ( .B(clk), .A(\g.we_clk [21836]));
Q_ASSIGN U10939 ( .B(clk), .A(\g.we_clk [21835]));
Q_ASSIGN U10940 ( .B(clk), .A(\g.we_clk [21834]));
Q_ASSIGN U10941 ( .B(clk), .A(\g.we_clk [21833]));
Q_ASSIGN U10942 ( .B(clk), .A(\g.we_clk [21832]));
Q_ASSIGN U10943 ( .B(clk), .A(\g.we_clk [21831]));
Q_ASSIGN U10944 ( .B(clk), .A(\g.we_clk [21830]));
Q_ASSIGN U10945 ( .B(clk), .A(\g.we_clk [21829]));
Q_ASSIGN U10946 ( .B(clk), .A(\g.we_clk [21828]));
Q_ASSIGN U10947 ( .B(clk), .A(\g.we_clk [21827]));
Q_ASSIGN U10948 ( .B(clk), .A(\g.we_clk [21826]));
Q_ASSIGN U10949 ( .B(clk), .A(\g.we_clk [21825]));
Q_ASSIGN U10950 ( .B(clk), .A(\g.we_clk [21824]));
Q_ASSIGN U10951 ( .B(clk), .A(\g.we_clk [21823]));
Q_ASSIGN U10952 ( .B(clk), .A(\g.we_clk [21822]));
Q_ASSIGN U10953 ( .B(clk), .A(\g.we_clk [21821]));
Q_ASSIGN U10954 ( .B(clk), .A(\g.we_clk [21820]));
Q_ASSIGN U10955 ( .B(clk), .A(\g.we_clk [21819]));
Q_ASSIGN U10956 ( .B(clk), .A(\g.we_clk [21818]));
Q_ASSIGN U10957 ( .B(clk), .A(\g.we_clk [21817]));
Q_ASSIGN U10958 ( .B(clk), .A(\g.we_clk [21816]));
Q_ASSIGN U10959 ( .B(clk), .A(\g.we_clk [21815]));
Q_ASSIGN U10960 ( .B(clk), .A(\g.we_clk [21814]));
Q_ASSIGN U10961 ( .B(clk), .A(\g.we_clk [21813]));
Q_ASSIGN U10962 ( .B(clk), .A(\g.we_clk [21812]));
Q_ASSIGN U10963 ( .B(clk), .A(\g.we_clk [21811]));
Q_ASSIGN U10964 ( .B(clk), .A(\g.we_clk [21810]));
Q_ASSIGN U10965 ( .B(clk), .A(\g.we_clk [21809]));
Q_ASSIGN U10966 ( .B(clk), .A(\g.we_clk [21808]));
Q_ASSIGN U10967 ( .B(clk), .A(\g.we_clk [21807]));
Q_ASSIGN U10968 ( .B(clk), .A(\g.we_clk [21806]));
Q_ASSIGN U10969 ( .B(clk), .A(\g.we_clk [21805]));
Q_ASSIGN U10970 ( .B(clk), .A(\g.we_clk [21804]));
Q_ASSIGN U10971 ( .B(clk), .A(\g.we_clk [21803]));
Q_ASSIGN U10972 ( .B(clk), .A(\g.we_clk [21802]));
Q_ASSIGN U10973 ( .B(clk), .A(\g.we_clk [21801]));
Q_ASSIGN U10974 ( .B(clk), .A(\g.we_clk [21800]));
Q_ASSIGN U10975 ( .B(clk), .A(\g.we_clk [21799]));
Q_ASSIGN U10976 ( .B(clk), .A(\g.we_clk [21798]));
Q_ASSIGN U10977 ( .B(clk), .A(\g.we_clk [21797]));
Q_ASSIGN U10978 ( .B(clk), .A(\g.we_clk [21796]));
Q_ASSIGN U10979 ( .B(clk), .A(\g.we_clk [21795]));
Q_ASSIGN U10980 ( .B(clk), .A(\g.we_clk [21794]));
Q_ASSIGN U10981 ( .B(clk), .A(\g.we_clk [21793]));
Q_ASSIGN U10982 ( .B(clk), .A(\g.we_clk [21792]));
Q_ASSIGN U10983 ( .B(clk), .A(\g.we_clk [21791]));
Q_ASSIGN U10984 ( .B(clk), .A(\g.we_clk [21790]));
Q_ASSIGN U10985 ( .B(clk), .A(\g.we_clk [21789]));
Q_ASSIGN U10986 ( .B(clk), .A(\g.we_clk [21788]));
Q_ASSIGN U10987 ( .B(clk), .A(\g.we_clk [21787]));
Q_ASSIGN U10988 ( .B(clk), .A(\g.we_clk [21786]));
Q_ASSIGN U10989 ( .B(clk), .A(\g.we_clk [21785]));
Q_ASSIGN U10990 ( .B(clk), .A(\g.we_clk [21784]));
Q_ASSIGN U10991 ( .B(clk), .A(\g.we_clk [21783]));
Q_ASSIGN U10992 ( .B(clk), .A(\g.we_clk [21782]));
Q_ASSIGN U10993 ( .B(clk), .A(\g.we_clk [21781]));
Q_ASSIGN U10994 ( .B(clk), .A(\g.we_clk [21780]));
Q_ASSIGN U10995 ( .B(clk), .A(\g.we_clk [21779]));
Q_ASSIGN U10996 ( .B(clk), .A(\g.we_clk [21778]));
Q_ASSIGN U10997 ( .B(clk), .A(\g.we_clk [21777]));
Q_ASSIGN U10998 ( .B(clk), .A(\g.we_clk [21776]));
Q_ASSIGN U10999 ( .B(clk), .A(\g.we_clk [21775]));
Q_ASSIGN U11000 ( .B(clk), .A(\g.we_clk [21774]));
Q_ASSIGN U11001 ( .B(clk), .A(\g.we_clk [21773]));
Q_ASSIGN U11002 ( .B(clk), .A(\g.we_clk [21772]));
Q_ASSIGN U11003 ( .B(clk), .A(\g.we_clk [21771]));
Q_ASSIGN U11004 ( .B(clk), .A(\g.we_clk [21770]));
Q_ASSIGN U11005 ( .B(clk), .A(\g.we_clk [21769]));
Q_ASSIGN U11006 ( .B(clk), .A(\g.we_clk [21768]));
Q_ASSIGN U11007 ( .B(clk), .A(\g.we_clk [21767]));
Q_ASSIGN U11008 ( .B(clk), .A(\g.we_clk [21766]));
Q_ASSIGN U11009 ( .B(clk), .A(\g.we_clk [21765]));
Q_ASSIGN U11010 ( .B(clk), .A(\g.we_clk [21764]));
Q_ASSIGN U11011 ( .B(clk), .A(\g.we_clk [21763]));
Q_ASSIGN U11012 ( .B(clk), .A(\g.we_clk [21762]));
Q_ASSIGN U11013 ( .B(clk), .A(\g.we_clk [21761]));
Q_ASSIGN U11014 ( .B(clk), .A(\g.we_clk [21760]));
Q_ASSIGN U11015 ( .B(clk), .A(\g.we_clk [21759]));
Q_ASSIGN U11016 ( .B(clk), .A(\g.we_clk [21758]));
Q_ASSIGN U11017 ( .B(clk), .A(\g.we_clk [21757]));
Q_ASSIGN U11018 ( .B(clk), .A(\g.we_clk [21756]));
Q_ASSIGN U11019 ( .B(clk), .A(\g.we_clk [21755]));
Q_ASSIGN U11020 ( .B(clk), .A(\g.we_clk [21754]));
Q_ASSIGN U11021 ( .B(clk), .A(\g.we_clk [21753]));
Q_ASSIGN U11022 ( .B(clk), .A(\g.we_clk [21752]));
Q_ASSIGN U11023 ( .B(clk), .A(\g.we_clk [21751]));
Q_ASSIGN U11024 ( .B(clk), .A(\g.we_clk [21750]));
Q_ASSIGN U11025 ( .B(clk), .A(\g.we_clk [21749]));
Q_ASSIGN U11026 ( .B(clk), .A(\g.we_clk [21748]));
Q_ASSIGN U11027 ( .B(clk), .A(\g.we_clk [21747]));
Q_ASSIGN U11028 ( .B(clk), .A(\g.we_clk [21746]));
Q_ASSIGN U11029 ( .B(clk), .A(\g.we_clk [21745]));
Q_ASSIGN U11030 ( .B(clk), .A(\g.we_clk [21744]));
Q_ASSIGN U11031 ( .B(clk), .A(\g.we_clk [21743]));
Q_ASSIGN U11032 ( .B(clk), .A(\g.we_clk [21742]));
Q_ASSIGN U11033 ( .B(clk), .A(\g.we_clk [21741]));
Q_ASSIGN U11034 ( .B(clk), .A(\g.we_clk [21740]));
Q_ASSIGN U11035 ( .B(clk), .A(\g.we_clk [21739]));
Q_ASSIGN U11036 ( .B(clk), .A(\g.we_clk [21738]));
Q_ASSIGN U11037 ( .B(clk), .A(\g.we_clk [21737]));
Q_ASSIGN U11038 ( .B(clk), .A(\g.we_clk [21736]));
Q_ASSIGN U11039 ( .B(clk), .A(\g.we_clk [21735]));
Q_ASSIGN U11040 ( .B(clk), .A(\g.we_clk [21734]));
Q_ASSIGN U11041 ( .B(clk), .A(\g.we_clk [21733]));
Q_ASSIGN U11042 ( .B(clk), .A(\g.we_clk [21732]));
Q_ASSIGN U11043 ( .B(clk), .A(\g.we_clk [21731]));
Q_ASSIGN U11044 ( .B(clk), .A(\g.we_clk [21730]));
Q_ASSIGN U11045 ( .B(clk), .A(\g.we_clk [21729]));
Q_ASSIGN U11046 ( .B(clk), .A(\g.we_clk [21728]));
Q_ASSIGN U11047 ( .B(clk), .A(\g.we_clk [21727]));
Q_ASSIGN U11048 ( .B(clk), .A(\g.we_clk [21726]));
Q_ASSIGN U11049 ( .B(clk), .A(\g.we_clk [21725]));
Q_ASSIGN U11050 ( .B(clk), .A(\g.we_clk [21724]));
Q_ASSIGN U11051 ( .B(clk), .A(\g.we_clk [21723]));
Q_ASSIGN U11052 ( .B(clk), .A(\g.we_clk [21722]));
Q_ASSIGN U11053 ( .B(clk), .A(\g.we_clk [21721]));
Q_ASSIGN U11054 ( .B(clk), .A(\g.we_clk [21720]));
Q_ASSIGN U11055 ( .B(clk), .A(\g.we_clk [21719]));
Q_ASSIGN U11056 ( .B(clk), .A(\g.we_clk [21718]));
Q_ASSIGN U11057 ( .B(clk), .A(\g.we_clk [21717]));
Q_ASSIGN U11058 ( .B(clk), .A(\g.we_clk [21716]));
Q_ASSIGN U11059 ( .B(clk), .A(\g.we_clk [21715]));
Q_ASSIGN U11060 ( .B(clk), .A(\g.we_clk [21714]));
Q_ASSIGN U11061 ( .B(clk), .A(\g.we_clk [21713]));
Q_ASSIGN U11062 ( .B(clk), .A(\g.we_clk [21712]));
Q_ASSIGN U11063 ( .B(clk), .A(\g.we_clk [21711]));
Q_ASSIGN U11064 ( .B(clk), .A(\g.we_clk [21710]));
Q_ASSIGN U11065 ( .B(clk), .A(\g.we_clk [21709]));
Q_ASSIGN U11066 ( .B(clk), .A(\g.we_clk [21708]));
Q_ASSIGN U11067 ( .B(clk), .A(\g.we_clk [21707]));
Q_ASSIGN U11068 ( .B(clk), .A(\g.we_clk [21706]));
Q_ASSIGN U11069 ( .B(clk), .A(\g.we_clk [21705]));
Q_ASSIGN U11070 ( .B(clk), .A(\g.we_clk [21704]));
Q_ASSIGN U11071 ( .B(clk), .A(\g.we_clk [21703]));
Q_ASSIGN U11072 ( .B(clk), .A(\g.we_clk [21702]));
Q_ASSIGN U11073 ( .B(clk), .A(\g.we_clk [21701]));
Q_ASSIGN U11074 ( .B(clk), .A(\g.we_clk [21700]));
Q_ASSIGN U11075 ( .B(clk), .A(\g.we_clk [21699]));
Q_ASSIGN U11076 ( .B(clk), .A(\g.we_clk [21698]));
Q_ASSIGN U11077 ( .B(clk), .A(\g.we_clk [21697]));
Q_ASSIGN U11078 ( .B(clk), .A(\g.we_clk [21696]));
Q_ASSIGN U11079 ( .B(clk), .A(\g.we_clk [21695]));
Q_ASSIGN U11080 ( .B(clk), .A(\g.we_clk [21694]));
Q_ASSIGN U11081 ( .B(clk), .A(\g.we_clk [21693]));
Q_ASSIGN U11082 ( .B(clk), .A(\g.we_clk [21692]));
Q_ASSIGN U11083 ( .B(clk), .A(\g.we_clk [21691]));
Q_ASSIGN U11084 ( .B(clk), .A(\g.we_clk [21690]));
Q_ASSIGN U11085 ( .B(clk), .A(\g.we_clk [21689]));
Q_ASSIGN U11086 ( .B(clk), .A(\g.we_clk [21688]));
Q_ASSIGN U11087 ( .B(clk), .A(\g.we_clk [21687]));
Q_ASSIGN U11088 ( .B(clk), .A(\g.we_clk [21686]));
Q_ASSIGN U11089 ( .B(clk), .A(\g.we_clk [21685]));
Q_ASSIGN U11090 ( .B(clk), .A(\g.we_clk [21684]));
Q_ASSIGN U11091 ( .B(clk), .A(\g.we_clk [21683]));
Q_ASSIGN U11092 ( .B(clk), .A(\g.we_clk [21682]));
Q_ASSIGN U11093 ( .B(clk), .A(\g.we_clk [21681]));
Q_ASSIGN U11094 ( .B(clk), .A(\g.we_clk [21680]));
Q_ASSIGN U11095 ( .B(clk), .A(\g.we_clk [21679]));
Q_ASSIGN U11096 ( .B(clk), .A(\g.we_clk [21678]));
Q_ASSIGN U11097 ( .B(clk), .A(\g.we_clk [21677]));
Q_ASSIGN U11098 ( .B(clk), .A(\g.we_clk [21676]));
Q_ASSIGN U11099 ( .B(clk), .A(\g.we_clk [21675]));
Q_ASSIGN U11100 ( .B(clk), .A(\g.we_clk [21674]));
Q_ASSIGN U11101 ( .B(clk), .A(\g.we_clk [21673]));
Q_ASSIGN U11102 ( .B(clk), .A(\g.we_clk [21672]));
Q_ASSIGN U11103 ( .B(clk), .A(\g.we_clk [21671]));
Q_ASSIGN U11104 ( .B(clk), .A(\g.we_clk [21670]));
Q_ASSIGN U11105 ( .B(clk), .A(\g.we_clk [21669]));
Q_ASSIGN U11106 ( .B(clk), .A(\g.we_clk [21668]));
Q_ASSIGN U11107 ( .B(clk), .A(\g.we_clk [21667]));
Q_ASSIGN U11108 ( .B(clk), .A(\g.we_clk [21666]));
Q_ASSIGN U11109 ( .B(clk), .A(\g.we_clk [21665]));
Q_ASSIGN U11110 ( .B(clk), .A(\g.we_clk [21664]));
Q_ASSIGN U11111 ( .B(clk), .A(\g.we_clk [21663]));
Q_ASSIGN U11112 ( .B(clk), .A(\g.we_clk [21662]));
Q_ASSIGN U11113 ( .B(clk), .A(\g.we_clk [21661]));
Q_ASSIGN U11114 ( .B(clk), .A(\g.we_clk [21660]));
Q_ASSIGN U11115 ( .B(clk), .A(\g.we_clk [21659]));
Q_ASSIGN U11116 ( .B(clk), .A(\g.we_clk [21658]));
Q_ASSIGN U11117 ( .B(clk), .A(\g.we_clk [21657]));
Q_ASSIGN U11118 ( .B(clk), .A(\g.we_clk [21656]));
Q_ASSIGN U11119 ( .B(clk), .A(\g.we_clk [21655]));
Q_ASSIGN U11120 ( .B(clk), .A(\g.we_clk [21654]));
Q_ASSIGN U11121 ( .B(clk), .A(\g.we_clk [21653]));
Q_ASSIGN U11122 ( .B(clk), .A(\g.we_clk [21652]));
Q_ASSIGN U11123 ( .B(clk), .A(\g.we_clk [21651]));
Q_ASSIGN U11124 ( .B(clk), .A(\g.we_clk [21650]));
Q_ASSIGN U11125 ( .B(clk), .A(\g.we_clk [21649]));
Q_ASSIGN U11126 ( .B(clk), .A(\g.we_clk [21648]));
Q_ASSIGN U11127 ( .B(clk), .A(\g.we_clk [21647]));
Q_ASSIGN U11128 ( .B(clk), .A(\g.we_clk [21646]));
Q_ASSIGN U11129 ( .B(clk), .A(\g.we_clk [21645]));
Q_ASSIGN U11130 ( .B(clk), .A(\g.we_clk [21644]));
Q_ASSIGN U11131 ( .B(clk), .A(\g.we_clk [21643]));
Q_ASSIGN U11132 ( .B(clk), .A(\g.we_clk [21642]));
Q_ASSIGN U11133 ( .B(clk), .A(\g.we_clk [21641]));
Q_ASSIGN U11134 ( .B(clk), .A(\g.we_clk [21640]));
Q_ASSIGN U11135 ( .B(clk), .A(\g.we_clk [21639]));
Q_ASSIGN U11136 ( .B(clk), .A(\g.we_clk [21638]));
Q_ASSIGN U11137 ( .B(clk), .A(\g.we_clk [21637]));
Q_ASSIGN U11138 ( .B(clk), .A(\g.we_clk [21636]));
Q_ASSIGN U11139 ( .B(clk), .A(\g.we_clk [21635]));
Q_ASSIGN U11140 ( .B(clk), .A(\g.we_clk [21634]));
Q_ASSIGN U11141 ( .B(clk), .A(\g.we_clk [21633]));
Q_ASSIGN U11142 ( .B(clk), .A(\g.we_clk [21632]));
Q_ASSIGN U11143 ( .B(clk), .A(\g.we_clk [21631]));
Q_ASSIGN U11144 ( .B(clk), .A(\g.we_clk [21630]));
Q_ASSIGN U11145 ( .B(clk), .A(\g.we_clk [21629]));
Q_ASSIGN U11146 ( .B(clk), .A(\g.we_clk [21628]));
Q_ASSIGN U11147 ( .B(clk), .A(\g.we_clk [21627]));
Q_ASSIGN U11148 ( .B(clk), .A(\g.we_clk [21626]));
Q_ASSIGN U11149 ( .B(clk), .A(\g.we_clk [21625]));
Q_ASSIGN U11150 ( .B(clk), .A(\g.we_clk [21624]));
Q_ASSIGN U11151 ( .B(clk), .A(\g.we_clk [21623]));
Q_ASSIGN U11152 ( .B(clk), .A(\g.we_clk [21622]));
Q_ASSIGN U11153 ( .B(clk), .A(\g.we_clk [21621]));
Q_ASSIGN U11154 ( .B(clk), .A(\g.we_clk [21620]));
Q_ASSIGN U11155 ( .B(clk), .A(\g.we_clk [21619]));
Q_ASSIGN U11156 ( .B(clk), .A(\g.we_clk [21618]));
Q_ASSIGN U11157 ( .B(clk), .A(\g.we_clk [21617]));
Q_ASSIGN U11158 ( .B(clk), .A(\g.we_clk [21616]));
Q_ASSIGN U11159 ( .B(clk), .A(\g.we_clk [21615]));
Q_ASSIGN U11160 ( .B(clk), .A(\g.we_clk [21614]));
Q_ASSIGN U11161 ( .B(clk), .A(\g.we_clk [21613]));
Q_ASSIGN U11162 ( .B(clk), .A(\g.we_clk [21612]));
Q_ASSIGN U11163 ( .B(clk), .A(\g.we_clk [21611]));
Q_ASSIGN U11164 ( .B(clk), .A(\g.we_clk [21610]));
Q_ASSIGN U11165 ( .B(clk), .A(\g.we_clk [21609]));
Q_ASSIGN U11166 ( .B(clk), .A(\g.we_clk [21608]));
Q_ASSIGN U11167 ( .B(clk), .A(\g.we_clk [21607]));
Q_ASSIGN U11168 ( .B(clk), .A(\g.we_clk [21606]));
Q_ASSIGN U11169 ( .B(clk), .A(\g.we_clk [21605]));
Q_ASSIGN U11170 ( .B(clk), .A(\g.we_clk [21604]));
Q_ASSIGN U11171 ( .B(clk), .A(\g.we_clk [21603]));
Q_ASSIGN U11172 ( .B(clk), .A(\g.we_clk [21602]));
Q_ASSIGN U11173 ( .B(clk), .A(\g.we_clk [21601]));
Q_ASSIGN U11174 ( .B(clk), .A(\g.we_clk [21600]));
Q_ASSIGN U11175 ( .B(clk), .A(\g.we_clk [21599]));
Q_ASSIGN U11176 ( .B(clk), .A(\g.we_clk [21598]));
Q_ASSIGN U11177 ( .B(clk), .A(\g.we_clk [21597]));
Q_ASSIGN U11178 ( .B(clk), .A(\g.we_clk [21596]));
Q_ASSIGN U11179 ( .B(clk), .A(\g.we_clk [21595]));
Q_ASSIGN U11180 ( .B(clk), .A(\g.we_clk [21594]));
Q_ASSIGN U11181 ( .B(clk), .A(\g.we_clk [21593]));
Q_ASSIGN U11182 ( .B(clk), .A(\g.we_clk [21592]));
Q_ASSIGN U11183 ( .B(clk), .A(\g.we_clk [21591]));
Q_ASSIGN U11184 ( .B(clk), .A(\g.we_clk [21590]));
Q_ASSIGN U11185 ( .B(clk), .A(\g.we_clk [21589]));
Q_ASSIGN U11186 ( .B(clk), .A(\g.we_clk [21588]));
Q_ASSIGN U11187 ( .B(clk), .A(\g.we_clk [21587]));
Q_ASSIGN U11188 ( .B(clk), .A(\g.we_clk [21586]));
Q_ASSIGN U11189 ( .B(clk), .A(\g.we_clk [21585]));
Q_ASSIGN U11190 ( .B(clk), .A(\g.we_clk [21584]));
Q_ASSIGN U11191 ( .B(clk), .A(\g.we_clk [21583]));
Q_ASSIGN U11192 ( .B(clk), .A(\g.we_clk [21582]));
Q_ASSIGN U11193 ( .B(clk), .A(\g.we_clk [21581]));
Q_ASSIGN U11194 ( .B(clk), .A(\g.we_clk [21580]));
Q_ASSIGN U11195 ( .B(clk), .A(\g.we_clk [21579]));
Q_ASSIGN U11196 ( .B(clk), .A(\g.we_clk [21578]));
Q_ASSIGN U11197 ( .B(clk), .A(\g.we_clk [21577]));
Q_ASSIGN U11198 ( .B(clk), .A(\g.we_clk [21576]));
Q_ASSIGN U11199 ( .B(clk), .A(\g.we_clk [21575]));
Q_ASSIGN U11200 ( .B(clk), .A(\g.we_clk [21574]));
Q_ASSIGN U11201 ( .B(clk), .A(\g.we_clk [21573]));
Q_ASSIGN U11202 ( .B(clk), .A(\g.we_clk [21572]));
Q_ASSIGN U11203 ( .B(clk), .A(\g.we_clk [21571]));
Q_ASSIGN U11204 ( .B(clk), .A(\g.we_clk [21570]));
Q_ASSIGN U11205 ( .B(clk), .A(\g.we_clk [21569]));
Q_ASSIGN U11206 ( .B(clk), .A(\g.we_clk [21568]));
Q_ASSIGN U11207 ( .B(clk), .A(\g.we_clk [21567]));
Q_ASSIGN U11208 ( .B(clk), .A(\g.we_clk [21566]));
Q_ASSIGN U11209 ( .B(clk), .A(\g.we_clk [21565]));
Q_ASSIGN U11210 ( .B(clk), .A(\g.we_clk [21564]));
Q_ASSIGN U11211 ( .B(clk), .A(\g.we_clk [21563]));
Q_ASSIGN U11212 ( .B(clk), .A(\g.we_clk [21562]));
Q_ASSIGN U11213 ( .B(clk), .A(\g.we_clk [21561]));
Q_ASSIGN U11214 ( .B(clk), .A(\g.we_clk [21560]));
Q_ASSIGN U11215 ( .B(clk), .A(\g.we_clk [21559]));
Q_ASSIGN U11216 ( .B(clk), .A(\g.we_clk [21558]));
Q_ASSIGN U11217 ( .B(clk), .A(\g.we_clk [21557]));
Q_ASSIGN U11218 ( .B(clk), .A(\g.we_clk [21556]));
Q_ASSIGN U11219 ( .B(clk), .A(\g.we_clk [21555]));
Q_ASSIGN U11220 ( .B(clk), .A(\g.we_clk [21554]));
Q_ASSIGN U11221 ( .B(clk), .A(\g.we_clk [21553]));
Q_ASSIGN U11222 ( .B(clk), .A(\g.we_clk [21552]));
Q_ASSIGN U11223 ( .B(clk), .A(\g.we_clk [21551]));
Q_ASSIGN U11224 ( .B(clk), .A(\g.we_clk [21550]));
Q_ASSIGN U11225 ( .B(clk), .A(\g.we_clk [21549]));
Q_ASSIGN U11226 ( .B(clk), .A(\g.we_clk [21548]));
Q_ASSIGN U11227 ( .B(clk), .A(\g.we_clk [21547]));
Q_ASSIGN U11228 ( .B(clk), .A(\g.we_clk [21546]));
Q_ASSIGN U11229 ( .B(clk), .A(\g.we_clk [21545]));
Q_ASSIGN U11230 ( .B(clk), .A(\g.we_clk [21544]));
Q_ASSIGN U11231 ( .B(clk), .A(\g.we_clk [21543]));
Q_ASSIGN U11232 ( .B(clk), .A(\g.we_clk [21542]));
Q_ASSIGN U11233 ( .B(clk), .A(\g.we_clk [21541]));
Q_ASSIGN U11234 ( .B(clk), .A(\g.we_clk [21540]));
Q_ASSIGN U11235 ( .B(clk), .A(\g.we_clk [21539]));
Q_ASSIGN U11236 ( .B(clk), .A(\g.we_clk [21538]));
Q_ASSIGN U11237 ( .B(clk), .A(\g.we_clk [21537]));
Q_ASSIGN U11238 ( .B(clk), .A(\g.we_clk [21536]));
Q_ASSIGN U11239 ( .B(clk), .A(\g.we_clk [21535]));
Q_ASSIGN U11240 ( .B(clk), .A(\g.we_clk [21534]));
Q_ASSIGN U11241 ( .B(clk), .A(\g.we_clk [21533]));
Q_ASSIGN U11242 ( .B(clk), .A(\g.we_clk [21532]));
Q_ASSIGN U11243 ( .B(clk), .A(\g.we_clk [21531]));
Q_ASSIGN U11244 ( .B(clk), .A(\g.we_clk [21530]));
Q_ASSIGN U11245 ( .B(clk), .A(\g.we_clk [21529]));
Q_ASSIGN U11246 ( .B(clk), .A(\g.we_clk [21528]));
Q_ASSIGN U11247 ( .B(clk), .A(\g.we_clk [21527]));
Q_ASSIGN U11248 ( .B(clk), .A(\g.we_clk [21526]));
Q_ASSIGN U11249 ( .B(clk), .A(\g.we_clk [21525]));
Q_ASSIGN U11250 ( .B(clk), .A(\g.we_clk [21524]));
Q_ASSIGN U11251 ( .B(clk), .A(\g.we_clk [21523]));
Q_ASSIGN U11252 ( .B(clk), .A(\g.we_clk [21522]));
Q_ASSIGN U11253 ( .B(clk), .A(\g.we_clk [21521]));
Q_ASSIGN U11254 ( .B(clk), .A(\g.we_clk [21520]));
Q_ASSIGN U11255 ( .B(clk), .A(\g.we_clk [21519]));
Q_ASSIGN U11256 ( .B(clk), .A(\g.we_clk [21518]));
Q_ASSIGN U11257 ( .B(clk), .A(\g.we_clk [21517]));
Q_ASSIGN U11258 ( .B(clk), .A(\g.we_clk [21516]));
Q_ASSIGN U11259 ( .B(clk), .A(\g.we_clk [21515]));
Q_ASSIGN U11260 ( .B(clk), .A(\g.we_clk [21514]));
Q_ASSIGN U11261 ( .B(clk), .A(\g.we_clk [21513]));
Q_ASSIGN U11262 ( .B(clk), .A(\g.we_clk [21512]));
Q_ASSIGN U11263 ( .B(clk), .A(\g.we_clk [21511]));
Q_ASSIGN U11264 ( .B(clk), .A(\g.we_clk [21510]));
Q_ASSIGN U11265 ( .B(clk), .A(\g.we_clk [21509]));
Q_ASSIGN U11266 ( .B(clk), .A(\g.we_clk [21508]));
Q_ASSIGN U11267 ( .B(clk), .A(\g.we_clk [21507]));
Q_ASSIGN U11268 ( .B(clk), .A(\g.we_clk [21506]));
Q_ASSIGN U11269 ( .B(clk), .A(\g.we_clk [21505]));
Q_ASSIGN U11270 ( .B(clk), .A(\g.we_clk [21504]));
Q_ASSIGN U11271 ( .B(clk), .A(\g.we_clk [21503]));
Q_ASSIGN U11272 ( .B(clk), .A(\g.we_clk [21502]));
Q_ASSIGN U11273 ( .B(clk), .A(\g.we_clk [21501]));
Q_ASSIGN U11274 ( .B(clk), .A(\g.we_clk [21500]));
Q_ASSIGN U11275 ( .B(clk), .A(\g.we_clk [21499]));
Q_ASSIGN U11276 ( .B(clk), .A(\g.we_clk [21498]));
Q_ASSIGN U11277 ( .B(clk), .A(\g.we_clk [21497]));
Q_ASSIGN U11278 ( .B(clk), .A(\g.we_clk [21496]));
Q_ASSIGN U11279 ( .B(clk), .A(\g.we_clk [21495]));
Q_ASSIGN U11280 ( .B(clk), .A(\g.we_clk [21494]));
Q_ASSIGN U11281 ( .B(clk), .A(\g.we_clk [21493]));
Q_ASSIGN U11282 ( .B(clk), .A(\g.we_clk [21492]));
Q_ASSIGN U11283 ( .B(clk), .A(\g.we_clk [21491]));
Q_ASSIGN U11284 ( .B(clk), .A(\g.we_clk [21490]));
Q_ASSIGN U11285 ( .B(clk), .A(\g.we_clk [21489]));
Q_ASSIGN U11286 ( .B(clk), .A(\g.we_clk [21488]));
Q_ASSIGN U11287 ( .B(clk), .A(\g.we_clk [21487]));
Q_ASSIGN U11288 ( .B(clk), .A(\g.we_clk [21486]));
Q_ASSIGN U11289 ( .B(clk), .A(\g.we_clk [21485]));
Q_ASSIGN U11290 ( .B(clk), .A(\g.we_clk [21484]));
Q_ASSIGN U11291 ( .B(clk), .A(\g.we_clk [21483]));
Q_ASSIGN U11292 ( .B(clk), .A(\g.we_clk [21482]));
Q_ASSIGN U11293 ( .B(clk), .A(\g.we_clk [21481]));
Q_ASSIGN U11294 ( .B(clk), .A(\g.we_clk [21480]));
Q_ASSIGN U11295 ( .B(clk), .A(\g.we_clk [21479]));
Q_ASSIGN U11296 ( .B(clk), .A(\g.we_clk [21478]));
Q_ASSIGN U11297 ( .B(clk), .A(\g.we_clk [21477]));
Q_ASSIGN U11298 ( .B(clk), .A(\g.we_clk [21476]));
Q_ASSIGN U11299 ( .B(clk), .A(\g.we_clk [21475]));
Q_ASSIGN U11300 ( .B(clk), .A(\g.we_clk [21474]));
Q_ASSIGN U11301 ( .B(clk), .A(\g.we_clk [21473]));
Q_ASSIGN U11302 ( .B(clk), .A(\g.we_clk [21472]));
Q_ASSIGN U11303 ( .B(clk), .A(\g.we_clk [21471]));
Q_ASSIGN U11304 ( .B(clk), .A(\g.we_clk [21470]));
Q_ASSIGN U11305 ( .B(clk), .A(\g.we_clk [21469]));
Q_ASSIGN U11306 ( .B(clk), .A(\g.we_clk [21468]));
Q_ASSIGN U11307 ( .B(clk), .A(\g.we_clk [21467]));
Q_ASSIGN U11308 ( .B(clk), .A(\g.we_clk [21466]));
Q_ASSIGN U11309 ( .B(clk), .A(\g.we_clk [21465]));
Q_ASSIGN U11310 ( .B(clk), .A(\g.we_clk [21464]));
Q_ASSIGN U11311 ( .B(clk), .A(\g.we_clk [21463]));
Q_ASSIGN U11312 ( .B(clk), .A(\g.we_clk [21462]));
Q_ASSIGN U11313 ( .B(clk), .A(\g.we_clk [21461]));
Q_ASSIGN U11314 ( .B(clk), .A(\g.we_clk [21460]));
Q_ASSIGN U11315 ( .B(clk), .A(\g.we_clk [21459]));
Q_ASSIGN U11316 ( .B(clk), .A(\g.we_clk [21458]));
Q_ASSIGN U11317 ( .B(clk), .A(\g.we_clk [21457]));
Q_ASSIGN U11318 ( .B(clk), .A(\g.we_clk [21456]));
Q_ASSIGN U11319 ( .B(clk), .A(\g.we_clk [21455]));
Q_ASSIGN U11320 ( .B(clk), .A(\g.we_clk [21454]));
Q_ASSIGN U11321 ( .B(clk), .A(\g.we_clk [21453]));
Q_ASSIGN U11322 ( .B(clk), .A(\g.we_clk [21452]));
Q_ASSIGN U11323 ( .B(clk), .A(\g.we_clk [21451]));
Q_ASSIGN U11324 ( .B(clk), .A(\g.we_clk [21450]));
Q_ASSIGN U11325 ( .B(clk), .A(\g.we_clk [21449]));
Q_ASSIGN U11326 ( .B(clk), .A(\g.we_clk [21448]));
Q_ASSIGN U11327 ( .B(clk), .A(\g.we_clk [21447]));
Q_ASSIGN U11328 ( .B(clk), .A(\g.we_clk [21446]));
Q_ASSIGN U11329 ( .B(clk), .A(\g.we_clk [21445]));
Q_ASSIGN U11330 ( .B(clk), .A(\g.we_clk [21444]));
Q_ASSIGN U11331 ( .B(clk), .A(\g.we_clk [21443]));
Q_ASSIGN U11332 ( .B(clk), .A(\g.we_clk [21442]));
Q_ASSIGN U11333 ( .B(clk), .A(\g.we_clk [21441]));
Q_ASSIGN U11334 ( .B(clk), .A(\g.we_clk [21440]));
Q_ASSIGN U11335 ( .B(clk), .A(\g.we_clk [21439]));
Q_ASSIGN U11336 ( .B(clk), .A(\g.we_clk [21438]));
Q_ASSIGN U11337 ( .B(clk), .A(\g.we_clk [21437]));
Q_ASSIGN U11338 ( .B(clk), .A(\g.we_clk [21436]));
Q_ASSIGN U11339 ( .B(clk), .A(\g.we_clk [21435]));
Q_ASSIGN U11340 ( .B(clk), .A(\g.we_clk [21434]));
Q_ASSIGN U11341 ( .B(clk), .A(\g.we_clk [21433]));
Q_ASSIGN U11342 ( .B(clk), .A(\g.we_clk [21432]));
Q_ASSIGN U11343 ( .B(clk), .A(\g.we_clk [21431]));
Q_ASSIGN U11344 ( .B(clk), .A(\g.we_clk [21430]));
Q_ASSIGN U11345 ( .B(clk), .A(\g.we_clk [21429]));
Q_ASSIGN U11346 ( .B(clk), .A(\g.we_clk [21428]));
Q_ASSIGN U11347 ( .B(clk), .A(\g.we_clk [21427]));
Q_ASSIGN U11348 ( .B(clk), .A(\g.we_clk [21426]));
Q_ASSIGN U11349 ( .B(clk), .A(\g.we_clk [21425]));
Q_ASSIGN U11350 ( .B(clk), .A(\g.we_clk [21424]));
Q_ASSIGN U11351 ( .B(clk), .A(\g.we_clk [21423]));
Q_ASSIGN U11352 ( .B(clk), .A(\g.we_clk [21422]));
Q_ASSIGN U11353 ( .B(clk), .A(\g.we_clk [21421]));
Q_ASSIGN U11354 ( .B(clk), .A(\g.we_clk [21420]));
Q_ASSIGN U11355 ( .B(clk), .A(\g.we_clk [21419]));
Q_ASSIGN U11356 ( .B(clk), .A(\g.we_clk [21418]));
Q_ASSIGN U11357 ( .B(clk), .A(\g.we_clk [21417]));
Q_ASSIGN U11358 ( .B(clk), .A(\g.we_clk [21416]));
Q_ASSIGN U11359 ( .B(clk), .A(\g.we_clk [21415]));
Q_ASSIGN U11360 ( .B(clk), .A(\g.we_clk [21414]));
Q_ASSIGN U11361 ( .B(clk), .A(\g.we_clk [21413]));
Q_ASSIGN U11362 ( .B(clk), .A(\g.we_clk [21412]));
Q_ASSIGN U11363 ( .B(clk), .A(\g.we_clk [21411]));
Q_ASSIGN U11364 ( .B(clk), .A(\g.we_clk [21410]));
Q_ASSIGN U11365 ( .B(clk), .A(\g.we_clk [21409]));
Q_ASSIGN U11366 ( .B(clk), .A(\g.we_clk [21408]));
Q_ASSIGN U11367 ( .B(clk), .A(\g.we_clk [21407]));
Q_ASSIGN U11368 ( .B(clk), .A(\g.we_clk [21406]));
Q_ASSIGN U11369 ( .B(clk), .A(\g.we_clk [21405]));
Q_ASSIGN U11370 ( .B(clk), .A(\g.we_clk [21404]));
Q_ASSIGN U11371 ( .B(clk), .A(\g.we_clk [21403]));
Q_ASSIGN U11372 ( .B(clk), .A(\g.we_clk [21402]));
Q_ASSIGN U11373 ( .B(clk), .A(\g.we_clk [21401]));
Q_ASSIGN U11374 ( .B(clk), .A(\g.we_clk [21400]));
Q_ASSIGN U11375 ( .B(clk), .A(\g.we_clk [21399]));
Q_ASSIGN U11376 ( .B(clk), .A(\g.we_clk [21398]));
Q_ASSIGN U11377 ( .B(clk), .A(\g.we_clk [21397]));
Q_ASSIGN U11378 ( .B(clk), .A(\g.we_clk [21396]));
Q_ASSIGN U11379 ( .B(clk), .A(\g.we_clk [21395]));
Q_ASSIGN U11380 ( .B(clk), .A(\g.we_clk [21394]));
Q_ASSIGN U11381 ( .B(clk), .A(\g.we_clk [21393]));
Q_ASSIGN U11382 ( .B(clk), .A(\g.we_clk [21392]));
Q_ASSIGN U11383 ( .B(clk), .A(\g.we_clk [21391]));
Q_ASSIGN U11384 ( .B(clk), .A(\g.we_clk [21390]));
Q_ASSIGN U11385 ( .B(clk), .A(\g.we_clk [21389]));
Q_ASSIGN U11386 ( .B(clk), .A(\g.we_clk [21388]));
Q_ASSIGN U11387 ( .B(clk), .A(\g.we_clk [21387]));
Q_ASSIGN U11388 ( .B(clk), .A(\g.we_clk [21386]));
Q_ASSIGN U11389 ( .B(clk), .A(\g.we_clk [21385]));
Q_ASSIGN U11390 ( .B(clk), .A(\g.we_clk [21384]));
Q_ASSIGN U11391 ( .B(clk), .A(\g.we_clk [21383]));
Q_ASSIGN U11392 ( .B(clk), .A(\g.we_clk [21382]));
Q_ASSIGN U11393 ( .B(clk), .A(\g.we_clk [21381]));
Q_ASSIGN U11394 ( .B(clk), .A(\g.we_clk [21380]));
Q_ASSIGN U11395 ( .B(clk), .A(\g.we_clk [21379]));
Q_ASSIGN U11396 ( .B(clk), .A(\g.we_clk [21378]));
Q_ASSIGN U11397 ( .B(clk), .A(\g.we_clk [21377]));
Q_ASSIGN U11398 ( .B(clk), .A(\g.we_clk [21376]));
Q_ASSIGN U11399 ( .B(clk), .A(\g.we_clk [21375]));
Q_ASSIGN U11400 ( .B(clk), .A(\g.we_clk [21374]));
Q_ASSIGN U11401 ( .B(clk), .A(\g.we_clk [21373]));
Q_ASSIGN U11402 ( .B(clk), .A(\g.we_clk [21372]));
Q_ASSIGN U11403 ( .B(clk), .A(\g.we_clk [21371]));
Q_ASSIGN U11404 ( .B(clk), .A(\g.we_clk [21370]));
Q_ASSIGN U11405 ( .B(clk), .A(\g.we_clk [21369]));
Q_ASSIGN U11406 ( .B(clk), .A(\g.we_clk [21368]));
Q_ASSIGN U11407 ( .B(clk), .A(\g.we_clk [21367]));
Q_ASSIGN U11408 ( .B(clk), .A(\g.we_clk [21366]));
Q_ASSIGN U11409 ( .B(clk), .A(\g.we_clk [21365]));
Q_ASSIGN U11410 ( .B(clk), .A(\g.we_clk [21364]));
Q_ASSIGN U11411 ( .B(clk), .A(\g.we_clk [21363]));
Q_ASSIGN U11412 ( .B(clk), .A(\g.we_clk [21362]));
Q_ASSIGN U11413 ( .B(clk), .A(\g.we_clk [21361]));
Q_ASSIGN U11414 ( .B(clk), .A(\g.we_clk [21360]));
Q_ASSIGN U11415 ( .B(clk), .A(\g.we_clk [21359]));
Q_ASSIGN U11416 ( .B(clk), .A(\g.we_clk [21358]));
Q_ASSIGN U11417 ( .B(clk), .A(\g.we_clk [21357]));
Q_ASSIGN U11418 ( .B(clk), .A(\g.we_clk [21356]));
Q_ASSIGN U11419 ( .B(clk), .A(\g.we_clk [21355]));
Q_ASSIGN U11420 ( .B(clk), .A(\g.we_clk [21354]));
Q_ASSIGN U11421 ( .B(clk), .A(\g.we_clk [21353]));
Q_ASSIGN U11422 ( .B(clk), .A(\g.we_clk [21352]));
Q_ASSIGN U11423 ( .B(clk), .A(\g.we_clk [21351]));
Q_ASSIGN U11424 ( .B(clk), .A(\g.we_clk [21350]));
Q_ASSIGN U11425 ( .B(clk), .A(\g.we_clk [21349]));
Q_ASSIGN U11426 ( .B(clk), .A(\g.we_clk [21348]));
Q_ASSIGN U11427 ( .B(clk), .A(\g.we_clk [21347]));
Q_ASSIGN U11428 ( .B(clk), .A(\g.we_clk [21346]));
Q_ASSIGN U11429 ( .B(clk), .A(\g.we_clk [21345]));
Q_ASSIGN U11430 ( .B(clk), .A(\g.we_clk [21344]));
Q_ASSIGN U11431 ( .B(clk), .A(\g.we_clk [21343]));
Q_ASSIGN U11432 ( .B(clk), .A(\g.we_clk [21342]));
Q_ASSIGN U11433 ( .B(clk), .A(\g.we_clk [21341]));
Q_ASSIGN U11434 ( .B(clk), .A(\g.we_clk [21340]));
Q_ASSIGN U11435 ( .B(clk), .A(\g.we_clk [21339]));
Q_ASSIGN U11436 ( .B(clk), .A(\g.we_clk [21338]));
Q_ASSIGN U11437 ( .B(clk), .A(\g.we_clk [21337]));
Q_ASSIGN U11438 ( .B(clk), .A(\g.we_clk [21336]));
Q_ASSIGN U11439 ( .B(clk), .A(\g.we_clk [21335]));
Q_ASSIGN U11440 ( .B(clk), .A(\g.we_clk [21334]));
Q_ASSIGN U11441 ( .B(clk), .A(\g.we_clk [21333]));
Q_ASSIGN U11442 ( .B(clk), .A(\g.we_clk [21332]));
Q_ASSIGN U11443 ( .B(clk), .A(\g.we_clk [21331]));
Q_ASSIGN U11444 ( .B(clk), .A(\g.we_clk [21330]));
Q_ASSIGN U11445 ( .B(clk), .A(\g.we_clk [21329]));
Q_ASSIGN U11446 ( .B(clk), .A(\g.we_clk [21328]));
Q_ASSIGN U11447 ( .B(clk), .A(\g.we_clk [21327]));
Q_ASSIGN U11448 ( .B(clk), .A(\g.we_clk [21326]));
Q_ASSIGN U11449 ( .B(clk), .A(\g.we_clk [21325]));
Q_ASSIGN U11450 ( .B(clk), .A(\g.we_clk [21324]));
Q_ASSIGN U11451 ( .B(clk), .A(\g.we_clk [21323]));
Q_ASSIGN U11452 ( .B(clk), .A(\g.we_clk [21322]));
Q_ASSIGN U11453 ( .B(clk), .A(\g.we_clk [21321]));
Q_ASSIGN U11454 ( .B(clk), .A(\g.we_clk [21320]));
Q_ASSIGN U11455 ( .B(clk), .A(\g.we_clk [21319]));
Q_ASSIGN U11456 ( .B(clk), .A(\g.we_clk [21318]));
Q_ASSIGN U11457 ( .B(clk), .A(\g.we_clk [21317]));
Q_ASSIGN U11458 ( .B(clk), .A(\g.we_clk [21316]));
Q_ASSIGN U11459 ( .B(clk), .A(\g.we_clk [21315]));
Q_ASSIGN U11460 ( .B(clk), .A(\g.we_clk [21314]));
Q_ASSIGN U11461 ( .B(clk), .A(\g.we_clk [21313]));
Q_ASSIGN U11462 ( .B(clk), .A(\g.we_clk [21312]));
Q_ASSIGN U11463 ( .B(clk), .A(\g.we_clk [21311]));
Q_ASSIGN U11464 ( .B(clk), .A(\g.we_clk [21310]));
Q_ASSIGN U11465 ( .B(clk), .A(\g.we_clk [21309]));
Q_ASSIGN U11466 ( .B(clk), .A(\g.we_clk [21308]));
Q_ASSIGN U11467 ( .B(clk), .A(\g.we_clk [21307]));
Q_ASSIGN U11468 ( .B(clk), .A(\g.we_clk [21306]));
Q_ASSIGN U11469 ( .B(clk), .A(\g.we_clk [21305]));
Q_ASSIGN U11470 ( .B(clk), .A(\g.we_clk [21304]));
Q_ASSIGN U11471 ( .B(clk), .A(\g.we_clk [21303]));
Q_ASSIGN U11472 ( .B(clk), .A(\g.we_clk [21302]));
Q_ASSIGN U11473 ( .B(clk), .A(\g.we_clk [21301]));
Q_ASSIGN U11474 ( .B(clk), .A(\g.we_clk [21300]));
Q_ASSIGN U11475 ( .B(clk), .A(\g.we_clk [21299]));
Q_ASSIGN U11476 ( .B(clk), .A(\g.we_clk [21298]));
Q_ASSIGN U11477 ( .B(clk), .A(\g.we_clk [21297]));
Q_ASSIGN U11478 ( .B(clk), .A(\g.we_clk [21296]));
Q_ASSIGN U11479 ( .B(clk), .A(\g.we_clk [21295]));
Q_ASSIGN U11480 ( .B(clk), .A(\g.we_clk [21294]));
Q_ASSIGN U11481 ( .B(clk), .A(\g.we_clk [21293]));
Q_ASSIGN U11482 ( .B(clk), .A(\g.we_clk [21292]));
Q_ASSIGN U11483 ( .B(clk), .A(\g.we_clk [21291]));
Q_ASSIGN U11484 ( .B(clk), .A(\g.we_clk [21290]));
Q_ASSIGN U11485 ( .B(clk), .A(\g.we_clk [21289]));
Q_ASSIGN U11486 ( .B(clk), .A(\g.we_clk [21288]));
Q_ASSIGN U11487 ( .B(clk), .A(\g.we_clk [21287]));
Q_ASSIGN U11488 ( .B(clk), .A(\g.we_clk [21286]));
Q_ASSIGN U11489 ( .B(clk), .A(\g.we_clk [21285]));
Q_ASSIGN U11490 ( .B(clk), .A(\g.we_clk [21284]));
Q_ASSIGN U11491 ( .B(clk), .A(\g.we_clk [21283]));
Q_ASSIGN U11492 ( .B(clk), .A(\g.we_clk [21282]));
Q_ASSIGN U11493 ( .B(clk), .A(\g.we_clk [21281]));
Q_ASSIGN U11494 ( .B(clk), .A(\g.we_clk [21280]));
Q_ASSIGN U11495 ( .B(clk), .A(\g.we_clk [21279]));
Q_ASSIGN U11496 ( .B(clk), .A(\g.we_clk [21278]));
Q_ASSIGN U11497 ( .B(clk), .A(\g.we_clk [21277]));
Q_ASSIGN U11498 ( .B(clk), .A(\g.we_clk [21276]));
Q_ASSIGN U11499 ( .B(clk), .A(\g.we_clk [21275]));
Q_ASSIGN U11500 ( .B(clk), .A(\g.we_clk [21274]));
Q_ASSIGN U11501 ( .B(clk), .A(\g.we_clk [21273]));
Q_ASSIGN U11502 ( .B(clk), .A(\g.we_clk [21272]));
Q_ASSIGN U11503 ( .B(clk), .A(\g.we_clk [21271]));
Q_ASSIGN U11504 ( .B(clk), .A(\g.we_clk [21270]));
Q_ASSIGN U11505 ( .B(clk), .A(\g.we_clk [21269]));
Q_ASSIGN U11506 ( .B(clk), .A(\g.we_clk [21268]));
Q_ASSIGN U11507 ( .B(clk), .A(\g.we_clk [21267]));
Q_ASSIGN U11508 ( .B(clk), .A(\g.we_clk [21266]));
Q_ASSIGN U11509 ( .B(clk), .A(\g.we_clk [21265]));
Q_ASSIGN U11510 ( .B(clk), .A(\g.we_clk [21264]));
Q_ASSIGN U11511 ( .B(clk), .A(\g.we_clk [21263]));
Q_ASSIGN U11512 ( .B(clk), .A(\g.we_clk [21262]));
Q_ASSIGN U11513 ( .B(clk), .A(\g.we_clk [21261]));
Q_ASSIGN U11514 ( .B(clk), .A(\g.we_clk [21260]));
Q_ASSIGN U11515 ( .B(clk), .A(\g.we_clk [21259]));
Q_ASSIGN U11516 ( .B(clk), .A(\g.we_clk [21258]));
Q_ASSIGN U11517 ( .B(clk), .A(\g.we_clk [21257]));
Q_ASSIGN U11518 ( .B(clk), .A(\g.we_clk [21256]));
Q_ASSIGN U11519 ( .B(clk), .A(\g.we_clk [21255]));
Q_ASSIGN U11520 ( .B(clk), .A(\g.we_clk [21254]));
Q_ASSIGN U11521 ( .B(clk), .A(\g.we_clk [21253]));
Q_ASSIGN U11522 ( .B(clk), .A(\g.we_clk [21252]));
Q_ASSIGN U11523 ( .B(clk), .A(\g.we_clk [21251]));
Q_ASSIGN U11524 ( .B(clk), .A(\g.we_clk [21250]));
Q_ASSIGN U11525 ( .B(clk), .A(\g.we_clk [21249]));
Q_ASSIGN U11526 ( .B(clk), .A(\g.we_clk [21248]));
Q_ASSIGN U11527 ( .B(clk), .A(\g.we_clk [21247]));
Q_ASSIGN U11528 ( .B(clk), .A(\g.we_clk [21246]));
Q_ASSIGN U11529 ( .B(clk), .A(\g.we_clk [21245]));
Q_ASSIGN U11530 ( .B(clk), .A(\g.we_clk [21244]));
Q_ASSIGN U11531 ( .B(clk), .A(\g.we_clk [21243]));
Q_ASSIGN U11532 ( .B(clk), .A(\g.we_clk [21242]));
Q_ASSIGN U11533 ( .B(clk), .A(\g.we_clk [21241]));
Q_ASSIGN U11534 ( .B(clk), .A(\g.we_clk [21240]));
Q_ASSIGN U11535 ( .B(clk), .A(\g.we_clk [21239]));
Q_ASSIGN U11536 ( .B(clk), .A(\g.we_clk [21238]));
Q_ASSIGN U11537 ( .B(clk), .A(\g.we_clk [21237]));
Q_ASSIGN U11538 ( .B(clk), .A(\g.we_clk [21236]));
Q_ASSIGN U11539 ( .B(clk), .A(\g.we_clk [21235]));
Q_ASSIGN U11540 ( .B(clk), .A(\g.we_clk [21234]));
Q_ASSIGN U11541 ( .B(clk), .A(\g.we_clk [21233]));
Q_ASSIGN U11542 ( .B(clk), .A(\g.we_clk [21232]));
Q_ASSIGN U11543 ( .B(clk), .A(\g.we_clk [21231]));
Q_ASSIGN U11544 ( .B(clk), .A(\g.we_clk [21230]));
Q_ASSIGN U11545 ( .B(clk), .A(\g.we_clk [21229]));
Q_ASSIGN U11546 ( .B(clk), .A(\g.we_clk [21228]));
Q_ASSIGN U11547 ( .B(clk), .A(\g.we_clk [21227]));
Q_ASSIGN U11548 ( .B(clk), .A(\g.we_clk [21226]));
Q_ASSIGN U11549 ( .B(clk), .A(\g.we_clk [21225]));
Q_ASSIGN U11550 ( .B(clk), .A(\g.we_clk [21224]));
Q_ASSIGN U11551 ( .B(clk), .A(\g.we_clk [21223]));
Q_ASSIGN U11552 ( .B(clk), .A(\g.we_clk [21222]));
Q_ASSIGN U11553 ( .B(clk), .A(\g.we_clk [21221]));
Q_ASSIGN U11554 ( .B(clk), .A(\g.we_clk [21220]));
Q_ASSIGN U11555 ( .B(clk), .A(\g.we_clk [21219]));
Q_ASSIGN U11556 ( .B(clk), .A(\g.we_clk [21218]));
Q_ASSIGN U11557 ( .B(clk), .A(\g.we_clk [21217]));
Q_ASSIGN U11558 ( .B(clk), .A(\g.we_clk [21216]));
Q_ASSIGN U11559 ( .B(clk), .A(\g.we_clk [21215]));
Q_ASSIGN U11560 ( .B(clk), .A(\g.we_clk [21214]));
Q_ASSIGN U11561 ( .B(clk), .A(\g.we_clk [21213]));
Q_ASSIGN U11562 ( .B(clk), .A(\g.we_clk [21212]));
Q_ASSIGN U11563 ( .B(clk), .A(\g.we_clk [21211]));
Q_ASSIGN U11564 ( .B(clk), .A(\g.we_clk [21210]));
Q_ASSIGN U11565 ( .B(clk), .A(\g.we_clk [21209]));
Q_ASSIGN U11566 ( .B(clk), .A(\g.we_clk [21208]));
Q_ASSIGN U11567 ( .B(clk), .A(\g.we_clk [21207]));
Q_ASSIGN U11568 ( .B(clk), .A(\g.we_clk [21206]));
Q_ASSIGN U11569 ( .B(clk), .A(\g.we_clk [21205]));
Q_ASSIGN U11570 ( .B(clk), .A(\g.we_clk [21204]));
Q_ASSIGN U11571 ( .B(clk), .A(\g.we_clk [21203]));
Q_ASSIGN U11572 ( .B(clk), .A(\g.we_clk [21202]));
Q_ASSIGN U11573 ( .B(clk), .A(\g.we_clk [21201]));
Q_ASSIGN U11574 ( .B(clk), .A(\g.we_clk [21200]));
Q_ASSIGN U11575 ( .B(clk), .A(\g.we_clk [21199]));
Q_ASSIGN U11576 ( .B(clk), .A(\g.we_clk [21198]));
Q_ASSIGN U11577 ( .B(clk), .A(\g.we_clk [21197]));
Q_ASSIGN U11578 ( .B(clk), .A(\g.we_clk [21196]));
Q_ASSIGN U11579 ( .B(clk), .A(\g.we_clk [21195]));
Q_ASSIGN U11580 ( .B(clk), .A(\g.we_clk [21194]));
Q_ASSIGN U11581 ( .B(clk), .A(\g.we_clk [21193]));
Q_ASSIGN U11582 ( .B(clk), .A(\g.we_clk [21192]));
Q_ASSIGN U11583 ( .B(clk), .A(\g.we_clk [21191]));
Q_ASSIGN U11584 ( .B(clk), .A(\g.we_clk [21190]));
Q_ASSIGN U11585 ( .B(clk), .A(\g.we_clk [21189]));
Q_ASSIGN U11586 ( .B(clk), .A(\g.we_clk [21188]));
Q_ASSIGN U11587 ( .B(clk), .A(\g.we_clk [21187]));
Q_ASSIGN U11588 ( .B(clk), .A(\g.we_clk [21186]));
Q_ASSIGN U11589 ( .B(clk), .A(\g.we_clk [21185]));
Q_ASSIGN U11590 ( .B(clk), .A(\g.we_clk [21184]));
Q_ASSIGN U11591 ( .B(clk), .A(\g.we_clk [21183]));
Q_ASSIGN U11592 ( .B(clk), .A(\g.we_clk [21182]));
Q_ASSIGN U11593 ( .B(clk), .A(\g.we_clk [21181]));
Q_ASSIGN U11594 ( .B(clk), .A(\g.we_clk [21180]));
Q_ASSIGN U11595 ( .B(clk), .A(\g.we_clk [21179]));
Q_ASSIGN U11596 ( .B(clk), .A(\g.we_clk [21178]));
Q_ASSIGN U11597 ( .B(clk), .A(\g.we_clk [21177]));
Q_ASSIGN U11598 ( .B(clk), .A(\g.we_clk [21176]));
Q_ASSIGN U11599 ( .B(clk), .A(\g.we_clk [21175]));
Q_ASSIGN U11600 ( .B(clk), .A(\g.we_clk [21174]));
Q_ASSIGN U11601 ( .B(clk), .A(\g.we_clk [21173]));
Q_ASSIGN U11602 ( .B(clk), .A(\g.we_clk [21172]));
Q_ASSIGN U11603 ( .B(clk), .A(\g.we_clk [21171]));
Q_ASSIGN U11604 ( .B(clk), .A(\g.we_clk [21170]));
Q_ASSIGN U11605 ( .B(clk), .A(\g.we_clk [21169]));
Q_ASSIGN U11606 ( .B(clk), .A(\g.we_clk [21168]));
Q_ASSIGN U11607 ( .B(clk), .A(\g.we_clk [21167]));
Q_ASSIGN U11608 ( .B(clk), .A(\g.we_clk [21166]));
Q_ASSIGN U11609 ( .B(clk), .A(\g.we_clk [21165]));
Q_ASSIGN U11610 ( .B(clk), .A(\g.we_clk [21164]));
Q_ASSIGN U11611 ( .B(clk), .A(\g.we_clk [21163]));
Q_ASSIGN U11612 ( .B(clk), .A(\g.we_clk [21162]));
Q_ASSIGN U11613 ( .B(clk), .A(\g.we_clk [21161]));
Q_ASSIGN U11614 ( .B(clk), .A(\g.we_clk [21160]));
Q_ASSIGN U11615 ( .B(clk), .A(\g.we_clk [21159]));
Q_ASSIGN U11616 ( .B(clk), .A(\g.we_clk [21158]));
Q_ASSIGN U11617 ( .B(clk), .A(\g.we_clk [21157]));
Q_ASSIGN U11618 ( .B(clk), .A(\g.we_clk [21156]));
Q_ASSIGN U11619 ( .B(clk), .A(\g.we_clk [21155]));
Q_ASSIGN U11620 ( .B(clk), .A(\g.we_clk [21154]));
Q_ASSIGN U11621 ( .B(clk), .A(\g.we_clk [21153]));
Q_ASSIGN U11622 ( .B(clk), .A(\g.we_clk [21152]));
Q_ASSIGN U11623 ( .B(clk), .A(\g.we_clk [21151]));
Q_ASSIGN U11624 ( .B(clk), .A(\g.we_clk [21150]));
Q_ASSIGN U11625 ( .B(clk), .A(\g.we_clk [21149]));
Q_ASSIGN U11626 ( .B(clk), .A(\g.we_clk [21148]));
Q_ASSIGN U11627 ( .B(clk), .A(\g.we_clk [21147]));
Q_ASSIGN U11628 ( .B(clk), .A(\g.we_clk [21146]));
Q_ASSIGN U11629 ( .B(clk), .A(\g.we_clk [21145]));
Q_ASSIGN U11630 ( .B(clk), .A(\g.we_clk [21144]));
Q_ASSIGN U11631 ( .B(clk), .A(\g.we_clk [21143]));
Q_ASSIGN U11632 ( .B(clk), .A(\g.we_clk [21142]));
Q_ASSIGN U11633 ( .B(clk), .A(\g.we_clk [21141]));
Q_ASSIGN U11634 ( .B(clk), .A(\g.we_clk [21140]));
Q_ASSIGN U11635 ( .B(clk), .A(\g.we_clk [21139]));
Q_ASSIGN U11636 ( .B(clk), .A(\g.we_clk [21138]));
Q_ASSIGN U11637 ( .B(clk), .A(\g.we_clk [21137]));
Q_ASSIGN U11638 ( .B(clk), .A(\g.we_clk [21136]));
Q_ASSIGN U11639 ( .B(clk), .A(\g.we_clk [21135]));
Q_ASSIGN U11640 ( .B(clk), .A(\g.we_clk [21134]));
Q_ASSIGN U11641 ( .B(clk), .A(\g.we_clk [21133]));
Q_ASSIGN U11642 ( .B(clk), .A(\g.we_clk [21132]));
Q_ASSIGN U11643 ( .B(clk), .A(\g.we_clk [21131]));
Q_ASSIGN U11644 ( .B(clk), .A(\g.we_clk [21130]));
Q_ASSIGN U11645 ( .B(clk), .A(\g.we_clk [21129]));
Q_ASSIGN U11646 ( .B(clk), .A(\g.we_clk [21128]));
Q_ASSIGN U11647 ( .B(clk), .A(\g.we_clk [21127]));
Q_ASSIGN U11648 ( .B(clk), .A(\g.we_clk [21126]));
Q_ASSIGN U11649 ( .B(clk), .A(\g.we_clk [21125]));
Q_ASSIGN U11650 ( .B(clk), .A(\g.we_clk [21124]));
Q_ASSIGN U11651 ( .B(clk), .A(\g.we_clk [21123]));
Q_ASSIGN U11652 ( .B(clk), .A(\g.we_clk [21122]));
Q_ASSIGN U11653 ( .B(clk), .A(\g.we_clk [21121]));
Q_ASSIGN U11654 ( .B(clk), .A(\g.we_clk [21120]));
Q_ASSIGN U11655 ( .B(clk), .A(\g.we_clk [21119]));
Q_ASSIGN U11656 ( .B(clk), .A(\g.we_clk [21118]));
Q_ASSIGN U11657 ( .B(clk), .A(\g.we_clk [21117]));
Q_ASSIGN U11658 ( .B(clk), .A(\g.we_clk [21116]));
Q_ASSIGN U11659 ( .B(clk), .A(\g.we_clk [21115]));
Q_ASSIGN U11660 ( .B(clk), .A(\g.we_clk [21114]));
Q_ASSIGN U11661 ( .B(clk), .A(\g.we_clk [21113]));
Q_ASSIGN U11662 ( .B(clk), .A(\g.we_clk [21112]));
Q_ASSIGN U11663 ( .B(clk), .A(\g.we_clk [21111]));
Q_ASSIGN U11664 ( .B(clk), .A(\g.we_clk [21110]));
Q_ASSIGN U11665 ( .B(clk), .A(\g.we_clk [21109]));
Q_ASSIGN U11666 ( .B(clk), .A(\g.we_clk [21108]));
Q_ASSIGN U11667 ( .B(clk), .A(\g.we_clk [21107]));
Q_ASSIGN U11668 ( .B(clk), .A(\g.we_clk [21106]));
Q_ASSIGN U11669 ( .B(clk), .A(\g.we_clk [21105]));
Q_ASSIGN U11670 ( .B(clk), .A(\g.we_clk [21104]));
Q_ASSIGN U11671 ( .B(clk), .A(\g.we_clk [21103]));
Q_ASSIGN U11672 ( .B(clk), .A(\g.we_clk [21102]));
Q_ASSIGN U11673 ( .B(clk), .A(\g.we_clk [21101]));
Q_ASSIGN U11674 ( .B(clk), .A(\g.we_clk [21100]));
Q_ASSIGN U11675 ( .B(clk), .A(\g.we_clk [21099]));
Q_ASSIGN U11676 ( .B(clk), .A(\g.we_clk [21098]));
Q_ASSIGN U11677 ( .B(clk), .A(\g.we_clk [21097]));
Q_ASSIGN U11678 ( .B(clk), .A(\g.we_clk [21096]));
Q_ASSIGN U11679 ( .B(clk), .A(\g.we_clk [21095]));
Q_ASSIGN U11680 ( .B(clk), .A(\g.we_clk [21094]));
Q_ASSIGN U11681 ( .B(clk), .A(\g.we_clk [21093]));
Q_ASSIGN U11682 ( .B(clk), .A(\g.we_clk [21092]));
Q_ASSIGN U11683 ( .B(clk), .A(\g.we_clk [21091]));
Q_ASSIGN U11684 ( .B(clk), .A(\g.we_clk [21090]));
Q_ASSIGN U11685 ( .B(clk), .A(\g.we_clk [21089]));
Q_ASSIGN U11686 ( .B(clk), .A(\g.we_clk [21088]));
Q_ASSIGN U11687 ( .B(clk), .A(\g.we_clk [21087]));
Q_ASSIGN U11688 ( .B(clk), .A(\g.we_clk [21086]));
Q_ASSIGN U11689 ( .B(clk), .A(\g.we_clk [21085]));
Q_ASSIGN U11690 ( .B(clk), .A(\g.we_clk [21084]));
Q_ASSIGN U11691 ( .B(clk), .A(\g.we_clk [21083]));
Q_ASSIGN U11692 ( .B(clk), .A(\g.we_clk [21082]));
Q_ASSIGN U11693 ( .B(clk), .A(\g.we_clk [21081]));
Q_ASSIGN U11694 ( .B(clk), .A(\g.we_clk [21080]));
Q_ASSIGN U11695 ( .B(clk), .A(\g.we_clk [21079]));
Q_ASSIGN U11696 ( .B(clk), .A(\g.we_clk [21078]));
Q_ASSIGN U11697 ( .B(clk), .A(\g.we_clk [21077]));
Q_ASSIGN U11698 ( .B(clk), .A(\g.we_clk [21076]));
Q_ASSIGN U11699 ( .B(clk), .A(\g.we_clk [21075]));
Q_ASSIGN U11700 ( .B(clk), .A(\g.we_clk [21074]));
Q_ASSIGN U11701 ( .B(clk), .A(\g.we_clk [21073]));
Q_ASSIGN U11702 ( .B(clk), .A(\g.we_clk [21072]));
Q_ASSIGN U11703 ( .B(clk), .A(\g.we_clk [21071]));
Q_ASSIGN U11704 ( .B(clk), .A(\g.we_clk [21070]));
Q_ASSIGN U11705 ( .B(clk), .A(\g.we_clk [21069]));
Q_ASSIGN U11706 ( .B(clk), .A(\g.we_clk [21068]));
Q_ASSIGN U11707 ( .B(clk), .A(\g.we_clk [21067]));
Q_ASSIGN U11708 ( .B(clk), .A(\g.we_clk [21066]));
Q_ASSIGN U11709 ( .B(clk), .A(\g.we_clk [21065]));
Q_ASSIGN U11710 ( .B(clk), .A(\g.we_clk [21064]));
Q_ASSIGN U11711 ( .B(clk), .A(\g.we_clk [21063]));
Q_ASSIGN U11712 ( .B(clk), .A(\g.we_clk [21062]));
Q_ASSIGN U11713 ( .B(clk), .A(\g.we_clk [21061]));
Q_ASSIGN U11714 ( .B(clk), .A(\g.we_clk [21060]));
Q_ASSIGN U11715 ( .B(clk), .A(\g.we_clk [21059]));
Q_ASSIGN U11716 ( .B(clk), .A(\g.we_clk [21058]));
Q_ASSIGN U11717 ( .B(clk), .A(\g.we_clk [21057]));
Q_ASSIGN U11718 ( .B(clk), .A(\g.we_clk [21056]));
Q_ASSIGN U11719 ( .B(clk), .A(\g.we_clk [21055]));
Q_ASSIGN U11720 ( .B(clk), .A(\g.we_clk [21054]));
Q_ASSIGN U11721 ( .B(clk), .A(\g.we_clk [21053]));
Q_ASSIGN U11722 ( .B(clk), .A(\g.we_clk [21052]));
Q_ASSIGN U11723 ( .B(clk), .A(\g.we_clk [21051]));
Q_ASSIGN U11724 ( .B(clk), .A(\g.we_clk [21050]));
Q_ASSIGN U11725 ( .B(clk), .A(\g.we_clk [21049]));
Q_ASSIGN U11726 ( .B(clk), .A(\g.we_clk [21048]));
Q_ASSIGN U11727 ( .B(clk), .A(\g.we_clk [21047]));
Q_ASSIGN U11728 ( .B(clk), .A(\g.we_clk [21046]));
Q_ASSIGN U11729 ( .B(clk), .A(\g.we_clk [21045]));
Q_ASSIGN U11730 ( .B(clk), .A(\g.we_clk [21044]));
Q_ASSIGN U11731 ( .B(clk), .A(\g.we_clk [21043]));
Q_ASSIGN U11732 ( .B(clk), .A(\g.we_clk [21042]));
Q_ASSIGN U11733 ( .B(clk), .A(\g.we_clk [21041]));
Q_ASSIGN U11734 ( .B(clk), .A(\g.we_clk [21040]));
Q_ASSIGN U11735 ( .B(clk), .A(\g.we_clk [21039]));
Q_ASSIGN U11736 ( .B(clk), .A(\g.we_clk [21038]));
Q_ASSIGN U11737 ( .B(clk), .A(\g.we_clk [21037]));
Q_ASSIGN U11738 ( .B(clk), .A(\g.we_clk [21036]));
Q_ASSIGN U11739 ( .B(clk), .A(\g.we_clk [21035]));
Q_ASSIGN U11740 ( .B(clk), .A(\g.we_clk [21034]));
Q_ASSIGN U11741 ( .B(clk), .A(\g.we_clk [21033]));
Q_ASSIGN U11742 ( .B(clk), .A(\g.we_clk [21032]));
Q_ASSIGN U11743 ( .B(clk), .A(\g.we_clk [21031]));
Q_ASSIGN U11744 ( .B(clk), .A(\g.we_clk [21030]));
Q_ASSIGN U11745 ( .B(clk), .A(\g.we_clk [21029]));
Q_ASSIGN U11746 ( .B(clk), .A(\g.we_clk [21028]));
Q_ASSIGN U11747 ( .B(clk), .A(\g.we_clk [21027]));
Q_ASSIGN U11748 ( .B(clk), .A(\g.we_clk [21026]));
Q_ASSIGN U11749 ( .B(clk), .A(\g.we_clk [21025]));
Q_ASSIGN U11750 ( .B(clk), .A(\g.we_clk [21024]));
Q_ASSIGN U11751 ( .B(clk), .A(\g.we_clk [21023]));
Q_ASSIGN U11752 ( .B(clk), .A(\g.we_clk [21022]));
Q_ASSIGN U11753 ( .B(clk), .A(\g.we_clk [21021]));
Q_ASSIGN U11754 ( .B(clk), .A(\g.we_clk [21020]));
Q_ASSIGN U11755 ( .B(clk), .A(\g.we_clk [21019]));
Q_ASSIGN U11756 ( .B(clk), .A(\g.we_clk [21018]));
Q_ASSIGN U11757 ( .B(clk), .A(\g.we_clk [21017]));
Q_ASSIGN U11758 ( .B(clk), .A(\g.we_clk [21016]));
Q_ASSIGN U11759 ( .B(clk), .A(\g.we_clk [21015]));
Q_ASSIGN U11760 ( .B(clk), .A(\g.we_clk [21014]));
Q_ASSIGN U11761 ( .B(clk), .A(\g.we_clk [21013]));
Q_ASSIGN U11762 ( .B(clk), .A(\g.we_clk [21012]));
Q_ASSIGN U11763 ( .B(clk), .A(\g.we_clk [21011]));
Q_ASSIGN U11764 ( .B(clk), .A(\g.we_clk [21010]));
Q_ASSIGN U11765 ( .B(clk), .A(\g.we_clk [21009]));
Q_ASSIGN U11766 ( .B(clk), .A(\g.we_clk [21008]));
Q_ASSIGN U11767 ( .B(clk), .A(\g.we_clk [21007]));
Q_ASSIGN U11768 ( .B(clk), .A(\g.we_clk [21006]));
Q_ASSIGN U11769 ( .B(clk), .A(\g.we_clk [21005]));
Q_ASSIGN U11770 ( .B(clk), .A(\g.we_clk [21004]));
Q_ASSIGN U11771 ( .B(clk), .A(\g.we_clk [21003]));
Q_ASSIGN U11772 ( .B(clk), .A(\g.we_clk [21002]));
Q_ASSIGN U11773 ( .B(clk), .A(\g.we_clk [21001]));
Q_ASSIGN U11774 ( .B(clk), .A(\g.we_clk [21000]));
Q_ASSIGN U11775 ( .B(clk), .A(\g.we_clk [20999]));
Q_ASSIGN U11776 ( .B(clk), .A(\g.we_clk [20998]));
Q_ASSIGN U11777 ( .B(clk), .A(\g.we_clk [20997]));
Q_ASSIGN U11778 ( .B(clk), .A(\g.we_clk [20996]));
Q_ASSIGN U11779 ( .B(clk), .A(\g.we_clk [20995]));
Q_ASSIGN U11780 ( .B(clk), .A(\g.we_clk [20994]));
Q_ASSIGN U11781 ( .B(clk), .A(\g.we_clk [20993]));
Q_ASSIGN U11782 ( .B(clk), .A(\g.we_clk [20992]));
Q_ASSIGN U11783 ( .B(clk), .A(\g.we_clk [20991]));
Q_ASSIGN U11784 ( .B(clk), .A(\g.we_clk [20990]));
Q_ASSIGN U11785 ( .B(clk), .A(\g.we_clk [20989]));
Q_ASSIGN U11786 ( .B(clk), .A(\g.we_clk [20988]));
Q_ASSIGN U11787 ( .B(clk), .A(\g.we_clk [20987]));
Q_ASSIGN U11788 ( .B(clk), .A(\g.we_clk [20986]));
Q_ASSIGN U11789 ( .B(clk), .A(\g.we_clk [20985]));
Q_ASSIGN U11790 ( .B(clk), .A(\g.we_clk [20984]));
Q_ASSIGN U11791 ( .B(clk), .A(\g.we_clk [20983]));
Q_ASSIGN U11792 ( .B(clk), .A(\g.we_clk [20982]));
Q_ASSIGN U11793 ( .B(clk), .A(\g.we_clk [20981]));
Q_ASSIGN U11794 ( .B(clk), .A(\g.we_clk [20980]));
Q_ASSIGN U11795 ( .B(clk), .A(\g.we_clk [20979]));
Q_ASSIGN U11796 ( .B(clk), .A(\g.we_clk [20978]));
Q_ASSIGN U11797 ( .B(clk), .A(\g.we_clk [20977]));
Q_ASSIGN U11798 ( .B(clk), .A(\g.we_clk [20976]));
Q_ASSIGN U11799 ( .B(clk), .A(\g.we_clk [20975]));
Q_ASSIGN U11800 ( .B(clk), .A(\g.we_clk [20974]));
Q_ASSIGN U11801 ( .B(clk), .A(\g.we_clk [20973]));
Q_ASSIGN U11802 ( .B(clk), .A(\g.we_clk [20972]));
Q_ASSIGN U11803 ( .B(clk), .A(\g.we_clk [20971]));
Q_ASSIGN U11804 ( .B(clk), .A(\g.we_clk [20970]));
Q_ASSIGN U11805 ( .B(clk), .A(\g.we_clk [20969]));
Q_ASSIGN U11806 ( .B(clk), .A(\g.we_clk [20968]));
Q_ASSIGN U11807 ( .B(clk), .A(\g.we_clk [20967]));
Q_ASSIGN U11808 ( .B(clk), .A(\g.we_clk [20966]));
Q_ASSIGN U11809 ( .B(clk), .A(\g.we_clk [20965]));
Q_ASSIGN U11810 ( .B(clk), .A(\g.we_clk [20964]));
Q_ASSIGN U11811 ( .B(clk), .A(\g.we_clk [20963]));
Q_ASSIGN U11812 ( .B(clk), .A(\g.we_clk [20962]));
Q_ASSIGN U11813 ( .B(clk), .A(\g.we_clk [20961]));
Q_ASSIGN U11814 ( .B(clk), .A(\g.we_clk [20960]));
Q_ASSIGN U11815 ( .B(clk), .A(\g.we_clk [20959]));
Q_ASSIGN U11816 ( .B(clk), .A(\g.we_clk [20958]));
Q_ASSIGN U11817 ( .B(clk), .A(\g.we_clk [20957]));
Q_ASSIGN U11818 ( .B(clk), .A(\g.we_clk [20956]));
Q_ASSIGN U11819 ( .B(clk), .A(\g.we_clk [20955]));
Q_ASSIGN U11820 ( .B(clk), .A(\g.we_clk [20954]));
Q_ASSIGN U11821 ( .B(clk), .A(\g.we_clk [20953]));
Q_ASSIGN U11822 ( .B(clk), .A(\g.we_clk [20952]));
Q_ASSIGN U11823 ( .B(clk), .A(\g.we_clk [20951]));
Q_ASSIGN U11824 ( .B(clk), .A(\g.we_clk [20950]));
Q_ASSIGN U11825 ( .B(clk), .A(\g.we_clk [20949]));
Q_ASSIGN U11826 ( .B(clk), .A(\g.we_clk [20948]));
Q_ASSIGN U11827 ( .B(clk), .A(\g.we_clk [20947]));
Q_ASSIGN U11828 ( .B(clk), .A(\g.we_clk [20946]));
Q_ASSIGN U11829 ( .B(clk), .A(\g.we_clk [20945]));
Q_ASSIGN U11830 ( .B(clk), .A(\g.we_clk [20944]));
Q_ASSIGN U11831 ( .B(clk), .A(\g.we_clk [20943]));
Q_ASSIGN U11832 ( .B(clk), .A(\g.we_clk [20942]));
Q_ASSIGN U11833 ( .B(clk), .A(\g.we_clk [20941]));
Q_ASSIGN U11834 ( .B(clk), .A(\g.we_clk [20940]));
Q_ASSIGN U11835 ( .B(clk), .A(\g.we_clk [20939]));
Q_ASSIGN U11836 ( .B(clk), .A(\g.we_clk [20938]));
Q_ASSIGN U11837 ( .B(clk), .A(\g.we_clk [20937]));
Q_ASSIGN U11838 ( .B(clk), .A(\g.we_clk [20936]));
Q_ASSIGN U11839 ( .B(clk), .A(\g.we_clk [20935]));
Q_ASSIGN U11840 ( .B(clk), .A(\g.we_clk [20934]));
Q_ASSIGN U11841 ( .B(clk), .A(\g.we_clk [20933]));
Q_ASSIGN U11842 ( .B(clk), .A(\g.we_clk [20932]));
Q_ASSIGN U11843 ( .B(clk), .A(\g.we_clk [20931]));
Q_ASSIGN U11844 ( .B(clk), .A(\g.we_clk [20930]));
Q_ASSIGN U11845 ( .B(clk), .A(\g.we_clk [20929]));
Q_ASSIGN U11846 ( .B(clk), .A(\g.we_clk [20928]));
Q_ASSIGN U11847 ( .B(clk), .A(\g.we_clk [20927]));
Q_ASSIGN U11848 ( .B(clk), .A(\g.we_clk [20926]));
Q_ASSIGN U11849 ( .B(clk), .A(\g.we_clk [20925]));
Q_ASSIGN U11850 ( .B(clk), .A(\g.we_clk [20924]));
Q_ASSIGN U11851 ( .B(clk), .A(\g.we_clk [20923]));
Q_ASSIGN U11852 ( .B(clk), .A(\g.we_clk [20922]));
Q_ASSIGN U11853 ( .B(clk), .A(\g.we_clk [20921]));
Q_ASSIGN U11854 ( .B(clk), .A(\g.we_clk [20920]));
Q_ASSIGN U11855 ( .B(clk), .A(\g.we_clk [20919]));
Q_ASSIGN U11856 ( .B(clk), .A(\g.we_clk [20918]));
Q_ASSIGN U11857 ( .B(clk), .A(\g.we_clk [20917]));
Q_ASSIGN U11858 ( .B(clk), .A(\g.we_clk [20916]));
Q_ASSIGN U11859 ( .B(clk), .A(\g.we_clk [20915]));
Q_ASSIGN U11860 ( .B(clk), .A(\g.we_clk [20914]));
Q_ASSIGN U11861 ( .B(clk), .A(\g.we_clk [20913]));
Q_ASSIGN U11862 ( .B(clk), .A(\g.we_clk [20912]));
Q_ASSIGN U11863 ( .B(clk), .A(\g.we_clk [20911]));
Q_ASSIGN U11864 ( .B(clk), .A(\g.we_clk [20910]));
Q_ASSIGN U11865 ( .B(clk), .A(\g.we_clk [20909]));
Q_ASSIGN U11866 ( .B(clk), .A(\g.we_clk [20908]));
Q_ASSIGN U11867 ( .B(clk), .A(\g.we_clk [20907]));
Q_ASSIGN U11868 ( .B(clk), .A(\g.we_clk [20906]));
Q_ASSIGN U11869 ( .B(clk), .A(\g.we_clk [20905]));
Q_ASSIGN U11870 ( .B(clk), .A(\g.we_clk [20904]));
Q_ASSIGN U11871 ( .B(clk), .A(\g.we_clk [20903]));
Q_ASSIGN U11872 ( .B(clk), .A(\g.we_clk [20902]));
Q_ASSIGN U11873 ( .B(clk), .A(\g.we_clk [20901]));
Q_ASSIGN U11874 ( .B(clk), .A(\g.we_clk [20900]));
Q_ASSIGN U11875 ( .B(clk), .A(\g.we_clk [20899]));
Q_ASSIGN U11876 ( .B(clk), .A(\g.we_clk [20898]));
Q_ASSIGN U11877 ( .B(clk), .A(\g.we_clk [20897]));
Q_ASSIGN U11878 ( .B(clk), .A(\g.we_clk [20896]));
Q_ASSIGN U11879 ( .B(clk), .A(\g.we_clk [20895]));
Q_ASSIGN U11880 ( .B(clk), .A(\g.we_clk [20894]));
Q_ASSIGN U11881 ( .B(clk), .A(\g.we_clk [20893]));
Q_ASSIGN U11882 ( .B(clk), .A(\g.we_clk [20892]));
Q_ASSIGN U11883 ( .B(clk), .A(\g.we_clk [20891]));
Q_ASSIGN U11884 ( .B(clk), .A(\g.we_clk [20890]));
Q_ASSIGN U11885 ( .B(clk), .A(\g.we_clk [20889]));
Q_ASSIGN U11886 ( .B(clk), .A(\g.we_clk [20888]));
Q_ASSIGN U11887 ( .B(clk), .A(\g.we_clk [20887]));
Q_ASSIGN U11888 ( .B(clk), .A(\g.we_clk [20886]));
Q_ASSIGN U11889 ( .B(clk), .A(\g.we_clk [20885]));
Q_ASSIGN U11890 ( .B(clk), .A(\g.we_clk [20884]));
Q_ASSIGN U11891 ( .B(clk), .A(\g.we_clk [20883]));
Q_ASSIGN U11892 ( .B(clk), .A(\g.we_clk [20882]));
Q_ASSIGN U11893 ( .B(clk), .A(\g.we_clk [20881]));
Q_ASSIGN U11894 ( .B(clk), .A(\g.we_clk [20880]));
Q_ASSIGN U11895 ( .B(clk), .A(\g.we_clk [20879]));
Q_ASSIGN U11896 ( .B(clk), .A(\g.we_clk [20878]));
Q_ASSIGN U11897 ( .B(clk), .A(\g.we_clk [20877]));
Q_ASSIGN U11898 ( .B(clk), .A(\g.we_clk [20876]));
Q_ASSIGN U11899 ( .B(clk), .A(\g.we_clk [20875]));
Q_ASSIGN U11900 ( .B(clk), .A(\g.we_clk [20874]));
Q_ASSIGN U11901 ( .B(clk), .A(\g.we_clk [20873]));
Q_ASSIGN U11902 ( .B(clk), .A(\g.we_clk [20872]));
Q_ASSIGN U11903 ( .B(clk), .A(\g.we_clk [20871]));
Q_ASSIGN U11904 ( .B(clk), .A(\g.we_clk [20870]));
Q_ASSIGN U11905 ( .B(clk), .A(\g.we_clk [20869]));
Q_ASSIGN U11906 ( .B(clk), .A(\g.we_clk [20868]));
Q_ASSIGN U11907 ( .B(clk), .A(\g.we_clk [20867]));
Q_ASSIGN U11908 ( .B(clk), .A(\g.we_clk [20866]));
Q_ASSIGN U11909 ( .B(clk), .A(\g.we_clk [20865]));
Q_ASSIGN U11910 ( .B(clk), .A(\g.we_clk [20864]));
Q_ASSIGN U11911 ( .B(clk), .A(\g.we_clk [20863]));
Q_ASSIGN U11912 ( .B(clk), .A(\g.we_clk [20862]));
Q_ASSIGN U11913 ( .B(clk), .A(\g.we_clk [20861]));
Q_ASSIGN U11914 ( .B(clk), .A(\g.we_clk [20860]));
Q_ASSIGN U11915 ( .B(clk), .A(\g.we_clk [20859]));
Q_ASSIGN U11916 ( .B(clk), .A(\g.we_clk [20858]));
Q_ASSIGN U11917 ( .B(clk), .A(\g.we_clk [20857]));
Q_ASSIGN U11918 ( .B(clk), .A(\g.we_clk [20856]));
Q_ASSIGN U11919 ( .B(clk), .A(\g.we_clk [20855]));
Q_ASSIGN U11920 ( .B(clk), .A(\g.we_clk [20854]));
Q_ASSIGN U11921 ( .B(clk), .A(\g.we_clk [20853]));
Q_ASSIGN U11922 ( .B(clk), .A(\g.we_clk [20852]));
Q_ASSIGN U11923 ( .B(clk), .A(\g.we_clk [20851]));
Q_ASSIGN U11924 ( .B(clk), .A(\g.we_clk [20850]));
Q_ASSIGN U11925 ( .B(clk), .A(\g.we_clk [20849]));
Q_ASSIGN U11926 ( .B(clk), .A(\g.we_clk [20848]));
Q_ASSIGN U11927 ( .B(clk), .A(\g.we_clk [20847]));
Q_ASSIGN U11928 ( .B(clk), .A(\g.we_clk [20846]));
Q_ASSIGN U11929 ( .B(clk), .A(\g.we_clk [20845]));
Q_ASSIGN U11930 ( .B(clk), .A(\g.we_clk [20844]));
Q_ASSIGN U11931 ( .B(clk), .A(\g.we_clk [20843]));
Q_ASSIGN U11932 ( .B(clk), .A(\g.we_clk [20842]));
Q_ASSIGN U11933 ( .B(clk), .A(\g.we_clk [20841]));
Q_ASSIGN U11934 ( .B(clk), .A(\g.we_clk [20840]));
Q_ASSIGN U11935 ( .B(clk), .A(\g.we_clk [20839]));
Q_ASSIGN U11936 ( .B(clk), .A(\g.we_clk [20838]));
Q_ASSIGN U11937 ( .B(clk), .A(\g.we_clk [20837]));
Q_ASSIGN U11938 ( .B(clk), .A(\g.we_clk [20836]));
Q_ASSIGN U11939 ( .B(clk), .A(\g.we_clk [20835]));
Q_ASSIGN U11940 ( .B(clk), .A(\g.we_clk [20834]));
Q_ASSIGN U11941 ( .B(clk), .A(\g.we_clk [20833]));
Q_ASSIGN U11942 ( .B(clk), .A(\g.we_clk [20832]));
Q_ASSIGN U11943 ( .B(clk), .A(\g.we_clk [20831]));
Q_ASSIGN U11944 ( .B(clk), .A(\g.we_clk [20830]));
Q_ASSIGN U11945 ( .B(clk), .A(\g.we_clk [20829]));
Q_ASSIGN U11946 ( .B(clk), .A(\g.we_clk [20828]));
Q_ASSIGN U11947 ( .B(clk), .A(\g.we_clk [20827]));
Q_ASSIGN U11948 ( .B(clk), .A(\g.we_clk [20826]));
Q_ASSIGN U11949 ( .B(clk), .A(\g.we_clk [20825]));
Q_ASSIGN U11950 ( .B(clk), .A(\g.we_clk [20824]));
Q_ASSIGN U11951 ( .B(clk), .A(\g.we_clk [20823]));
Q_ASSIGN U11952 ( .B(clk), .A(\g.we_clk [20822]));
Q_ASSIGN U11953 ( .B(clk), .A(\g.we_clk [20821]));
Q_ASSIGN U11954 ( .B(clk), .A(\g.we_clk [20820]));
Q_ASSIGN U11955 ( .B(clk), .A(\g.we_clk [20819]));
Q_ASSIGN U11956 ( .B(clk), .A(\g.we_clk [20818]));
Q_ASSIGN U11957 ( .B(clk), .A(\g.we_clk [20817]));
Q_ASSIGN U11958 ( .B(clk), .A(\g.we_clk [20816]));
Q_ASSIGN U11959 ( .B(clk), .A(\g.we_clk [20815]));
Q_ASSIGN U11960 ( .B(clk), .A(\g.we_clk [20814]));
Q_ASSIGN U11961 ( .B(clk), .A(\g.we_clk [20813]));
Q_ASSIGN U11962 ( .B(clk), .A(\g.we_clk [20812]));
Q_ASSIGN U11963 ( .B(clk), .A(\g.we_clk [20811]));
Q_ASSIGN U11964 ( .B(clk), .A(\g.we_clk [20810]));
Q_ASSIGN U11965 ( .B(clk), .A(\g.we_clk [20809]));
Q_ASSIGN U11966 ( .B(clk), .A(\g.we_clk [20808]));
Q_ASSIGN U11967 ( .B(clk), .A(\g.we_clk [20807]));
Q_ASSIGN U11968 ( .B(clk), .A(\g.we_clk [20806]));
Q_ASSIGN U11969 ( .B(clk), .A(\g.we_clk [20805]));
Q_ASSIGN U11970 ( .B(clk), .A(\g.we_clk [20804]));
Q_ASSIGN U11971 ( .B(clk), .A(\g.we_clk [20803]));
Q_ASSIGN U11972 ( .B(clk), .A(\g.we_clk [20802]));
Q_ASSIGN U11973 ( .B(clk), .A(\g.we_clk [20801]));
Q_ASSIGN U11974 ( .B(clk), .A(\g.we_clk [20800]));
Q_ASSIGN U11975 ( .B(clk), .A(\g.we_clk [20799]));
Q_ASSIGN U11976 ( .B(clk), .A(\g.we_clk [20798]));
Q_ASSIGN U11977 ( .B(clk), .A(\g.we_clk [20797]));
Q_ASSIGN U11978 ( .B(clk), .A(\g.we_clk [20796]));
Q_ASSIGN U11979 ( .B(clk), .A(\g.we_clk [20795]));
Q_ASSIGN U11980 ( .B(clk), .A(\g.we_clk [20794]));
Q_ASSIGN U11981 ( .B(clk), .A(\g.we_clk [20793]));
Q_ASSIGN U11982 ( .B(clk), .A(\g.we_clk [20792]));
Q_ASSIGN U11983 ( .B(clk), .A(\g.we_clk [20791]));
Q_ASSIGN U11984 ( .B(clk), .A(\g.we_clk [20790]));
Q_ASSIGN U11985 ( .B(clk), .A(\g.we_clk [20789]));
Q_ASSIGN U11986 ( .B(clk), .A(\g.we_clk [20788]));
Q_ASSIGN U11987 ( .B(clk), .A(\g.we_clk [20787]));
Q_ASSIGN U11988 ( .B(clk), .A(\g.we_clk [20786]));
Q_ASSIGN U11989 ( .B(clk), .A(\g.we_clk [20785]));
Q_ASSIGN U11990 ( .B(clk), .A(\g.we_clk [20784]));
Q_ASSIGN U11991 ( .B(clk), .A(\g.we_clk [20783]));
Q_ASSIGN U11992 ( .B(clk), .A(\g.we_clk [20782]));
Q_ASSIGN U11993 ( .B(clk), .A(\g.we_clk [20781]));
Q_ASSIGN U11994 ( .B(clk), .A(\g.we_clk [20780]));
Q_ASSIGN U11995 ( .B(clk), .A(\g.we_clk [20779]));
Q_ASSIGN U11996 ( .B(clk), .A(\g.we_clk [20778]));
Q_ASSIGN U11997 ( .B(clk), .A(\g.we_clk [20777]));
Q_ASSIGN U11998 ( .B(clk), .A(\g.we_clk [20776]));
Q_ASSIGN U11999 ( .B(clk), .A(\g.we_clk [20775]));
Q_ASSIGN U12000 ( .B(clk), .A(\g.we_clk [20774]));
Q_ASSIGN U12001 ( .B(clk), .A(\g.we_clk [20773]));
Q_ASSIGN U12002 ( .B(clk), .A(\g.we_clk [20772]));
Q_ASSIGN U12003 ( .B(clk), .A(\g.we_clk [20771]));
Q_ASSIGN U12004 ( .B(clk), .A(\g.we_clk [20770]));
Q_ASSIGN U12005 ( .B(clk), .A(\g.we_clk [20769]));
Q_ASSIGN U12006 ( .B(clk), .A(\g.we_clk [20768]));
Q_ASSIGN U12007 ( .B(clk), .A(\g.we_clk [20767]));
Q_ASSIGN U12008 ( .B(clk), .A(\g.we_clk [20766]));
Q_ASSIGN U12009 ( .B(clk), .A(\g.we_clk [20765]));
Q_ASSIGN U12010 ( .B(clk), .A(\g.we_clk [20764]));
Q_ASSIGN U12011 ( .B(clk), .A(\g.we_clk [20763]));
Q_ASSIGN U12012 ( .B(clk), .A(\g.we_clk [20762]));
Q_ASSIGN U12013 ( .B(clk), .A(\g.we_clk [20761]));
Q_ASSIGN U12014 ( .B(clk), .A(\g.we_clk [20760]));
Q_ASSIGN U12015 ( .B(clk), .A(\g.we_clk [20759]));
Q_ASSIGN U12016 ( .B(clk), .A(\g.we_clk [20758]));
Q_ASSIGN U12017 ( .B(clk), .A(\g.we_clk [20757]));
Q_ASSIGN U12018 ( .B(clk), .A(\g.we_clk [20756]));
Q_ASSIGN U12019 ( .B(clk), .A(\g.we_clk [20755]));
Q_ASSIGN U12020 ( .B(clk), .A(\g.we_clk [20754]));
Q_ASSIGN U12021 ( .B(clk), .A(\g.we_clk [20753]));
Q_ASSIGN U12022 ( .B(clk), .A(\g.we_clk [20752]));
Q_ASSIGN U12023 ( .B(clk), .A(\g.we_clk [20751]));
Q_ASSIGN U12024 ( .B(clk), .A(\g.we_clk [20750]));
Q_ASSIGN U12025 ( .B(clk), .A(\g.we_clk [20749]));
Q_ASSIGN U12026 ( .B(clk), .A(\g.we_clk [20748]));
Q_ASSIGN U12027 ( .B(clk), .A(\g.we_clk [20747]));
Q_ASSIGN U12028 ( .B(clk), .A(\g.we_clk [20746]));
Q_ASSIGN U12029 ( .B(clk), .A(\g.we_clk [20745]));
Q_ASSIGN U12030 ( .B(clk), .A(\g.we_clk [20744]));
Q_ASSIGN U12031 ( .B(clk), .A(\g.we_clk [20743]));
Q_ASSIGN U12032 ( .B(clk), .A(\g.we_clk [20742]));
Q_ASSIGN U12033 ( .B(clk), .A(\g.we_clk [20741]));
Q_ASSIGN U12034 ( .B(clk), .A(\g.we_clk [20740]));
Q_ASSIGN U12035 ( .B(clk), .A(\g.we_clk [20739]));
Q_ASSIGN U12036 ( .B(clk), .A(\g.we_clk [20738]));
Q_ASSIGN U12037 ( .B(clk), .A(\g.we_clk [20737]));
Q_ASSIGN U12038 ( .B(clk), .A(\g.we_clk [20736]));
Q_ASSIGN U12039 ( .B(clk), .A(\g.we_clk [20735]));
Q_ASSIGN U12040 ( .B(clk), .A(\g.we_clk [20734]));
Q_ASSIGN U12041 ( .B(clk), .A(\g.we_clk [20733]));
Q_ASSIGN U12042 ( .B(clk), .A(\g.we_clk [20732]));
Q_ASSIGN U12043 ( .B(clk), .A(\g.we_clk [20731]));
Q_ASSIGN U12044 ( .B(clk), .A(\g.we_clk [20730]));
Q_ASSIGN U12045 ( .B(clk), .A(\g.we_clk [20729]));
Q_ASSIGN U12046 ( .B(clk), .A(\g.we_clk [20728]));
Q_ASSIGN U12047 ( .B(clk), .A(\g.we_clk [20727]));
Q_ASSIGN U12048 ( .B(clk), .A(\g.we_clk [20726]));
Q_ASSIGN U12049 ( .B(clk), .A(\g.we_clk [20725]));
Q_ASSIGN U12050 ( .B(clk), .A(\g.we_clk [20724]));
Q_ASSIGN U12051 ( .B(clk), .A(\g.we_clk [20723]));
Q_ASSIGN U12052 ( .B(clk), .A(\g.we_clk [20722]));
Q_ASSIGN U12053 ( .B(clk), .A(\g.we_clk [20721]));
Q_ASSIGN U12054 ( .B(clk), .A(\g.we_clk [20720]));
Q_ASSIGN U12055 ( .B(clk), .A(\g.we_clk [20719]));
Q_ASSIGN U12056 ( .B(clk), .A(\g.we_clk [20718]));
Q_ASSIGN U12057 ( .B(clk), .A(\g.we_clk [20717]));
Q_ASSIGN U12058 ( .B(clk), .A(\g.we_clk [20716]));
Q_ASSIGN U12059 ( .B(clk), .A(\g.we_clk [20715]));
Q_ASSIGN U12060 ( .B(clk), .A(\g.we_clk [20714]));
Q_ASSIGN U12061 ( .B(clk), .A(\g.we_clk [20713]));
Q_ASSIGN U12062 ( .B(clk), .A(\g.we_clk [20712]));
Q_ASSIGN U12063 ( .B(clk), .A(\g.we_clk [20711]));
Q_ASSIGN U12064 ( .B(clk), .A(\g.we_clk [20710]));
Q_ASSIGN U12065 ( .B(clk), .A(\g.we_clk [20709]));
Q_ASSIGN U12066 ( .B(clk), .A(\g.we_clk [20708]));
Q_ASSIGN U12067 ( .B(clk), .A(\g.we_clk [20707]));
Q_ASSIGN U12068 ( .B(clk), .A(\g.we_clk [20706]));
Q_ASSIGN U12069 ( .B(clk), .A(\g.we_clk [20705]));
Q_ASSIGN U12070 ( .B(clk), .A(\g.we_clk [20704]));
Q_ASSIGN U12071 ( .B(clk), .A(\g.we_clk [20703]));
Q_ASSIGN U12072 ( .B(clk), .A(\g.we_clk [20702]));
Q_ASSIGN U12073 ( .B(clk), .A(\g.we_clk [20701]));
Q_ASSIGN U12074 ( .B(clk), .A(\g.we_clk [20700]));
Q_ASSIGN U12075 ( .B(clk), .A(\g.we_clk [20699]));
Q_ASSIGN U12076 ( .B(clk), .A(\g.we_clk [20698]));
Q_ASSIGN U12077 ( .B(clk), .A(\g.we_clk [20697]));
Q_ASSIGN U12078 ( .B(clk), .A(\g.we_clk [20696]));
Q_ASSIGN U12079 ( .B(clk), .A(\g.we_clk [20695]));
Q_ASSIGN U12080 ( .B(clk), .A(\g.we_clk [20694]));
Q_ASSIGN U12081 ( .B(clk), .A(\g.we_clk [20693]));
Q_ASSIGN U12082 ( .B(clk), .A(\g.we_clk [20692]));
Q_ASSIGN U12083 ( .B(clk), .A(\g.we_clk [20691]));
Q_ASSIGN U12084 ( .B(clk), .A(\g.we_clk [20690]));
Q_ASSIGN U12085 ( .B(clk), .A(\g.we_clk [20689]));
Q_ASSIGN U12086 ( .B(clk), .A(\g.we_clk [20688]));
Q_ASSIGN U12087 ( .B(clk), .A(\g.we_clk [20687]));
Q_ASSIGN U12088 ( .B(clk), .A(\g.we_clk [20686]));
Q_ASSIGN U12089 ( .B(clk), .A(\g.we_clk [20685]));
Q_ASSIGN U12090 ( .B(clk), .A(\g.we_clk [20684]));
Q_ASSIGN U12091 ( .B(clk), .A(\g.we_clk [20683]));
Q_ASSIGN U12092 ( .B(clk), .A(\g.we_clk [20682]));
Q_ASSIGN U12093 ( .B(clk), .A(\g.we_clk [20681]));
Q_ASSIGN U12094 ( .B(clk), .A(\g.we_clk [20680]));
Q_ASSIGN U12095 ( .B(clk), .A(\g.we_clk [20679]));
Q_ASSIGN U12096 ( .B(clk), .A(\g.we_clk [20678]));
Q_ASSIGN U12097 ( .B(clk), .A(\g.we_clk [20677]));
Q_ASSIGN U12098 ( .B(clk), .A(\g.we_clk [20676]));
Q_ASSIGN U12099 ( .B(clk), .A(\g.we_clk [20675]));
Q_ASSIGN U12100 ( .B(clk), .A(\g.we_clk [20674]));
Q_ASSIGN U12101 ( .B(clk), .A(\g.we_clk [20673]));
Q_ASSIGN U12102 ( .B(clk), .A(\g.we_clk [20672]));
Q_ASSIGN U12103 ( .B(clk), .A(\g.we_clk [20671]));
Q_ASSIGN U12104 ( .B(clk), .A(\g.we_clk [20670]));
Q_ASSIGN U12105 ( .B(clk), .A(\g.we_clk [20669]));
Q_ASSIGN U12106 ( .B(clk), .A(\g.we_clk [20668]));
Q_ASSIGN U12107 ( .B(clk), .A(\g.we_clk [20667]));
Q_ASSIGN U12108 ( .B(clk), .A(\g.we_clk [20666]));
Q_ASSIGN U12109 ( .B(clk), .A(\g.we_clk [20665]));
Q_ASSIGN U12110 ( .B(clk), .A(\g.we_clk [20664]));
Q_ASSIGN U12111 ( .B(clk), .A(\g.we_clk [20663]));
Q_ASSIGN U12112 ( .B(clk), .A(\g.we_clk [20662]));
Q_ASSIGN U12113 ( .B(clk), .A(\g.we_clk [20661]));
Q_ASSIGN U12114 ( .B(clk), .A(\g.we_clk [20660]));
Q_ASSIGN U12115 ( .B(clk), .A(\g.we_clk [20659]));
Q_ASSIGN U12116 ( .B(clk), .A(\g.we_clk [20658]));
Q_ASSIGN U12117 ( .B(clk), .A(\g.we_clk [20657]));
Q_ASSIGN U12118 ( .B(clk), .A(\g.we_clk [20656]));
Q_ASSIGN U12119 ( .B(clk), .A(\g.we_clk [20655]));
Q_ASSIGN U12120 ( .B(clk), .A(\g.we_clk [20654]));
Q_ASSIGN U12121 ( .B(clk), .A(\g.we_clk [20653]));
Q_ASSIGN U12122 ( .B(clk), .A(\g.we_clk [20652]));
Q_ASSIGN U12123 ( .B(clk), .A(\g.we_clk [20651]));
Q_ASSIGN U12124 ( .B(clk), .A(\g.we_clk [20650]));
Q_ASSIGN U12125 ( .B(clk), .A(\g.we_clk [20649]));
Q_ASSIGN U12126 ( .B(clk), .A(\g.we_clk [20648]));
Q_ASSIGN U12127 ( .B(clk), .A(\g.we_clk [20647]));
Q_ASSIGN U12128 ( .B(clk), .A(\g.we_clk [20646]));
Q_ASSIGN U12129 ( .B(clk), .A(\g.we_clk [20645]));
Q_ASSIGN U12130 ( .B(clk), .A(\g.we_clk [20644]));
Q_ASSIGN U12131 ( .B(clk), .A(\g.we_clk [20643]));
Q_ASSIGN U12132 ( .B(clk), .A(\g.we_clk [20642]));
Q_ASSIGN U12133 ( .B(clk), .A(\g.we_clk [20641]));
Q_ASSIGN U12134 ( .B(clk), .A(\g.we_clk [20640]));
Q_ASSIGN U12135 ( .B(clk), .A(\g.we_clk [20639]));
Q_ASSIGN U12136 ( .B(clk), .A(\g.we_clk [20638]));
Q_ASSIGN U12137 ( .B(clk), .A(\g.we_clk [20637]));
Q_ASSIGN U12138 ( .B(clk), .A(\g.we_clk [20636]));
Q_ASSIGN U12139 ( .B(clk), .A(\g.we_clk [20635]));
Q_ASSIGN U12140 ( .B(clk), .A(\g.we_clk [20634]));
Q_ASSIGN U12141 ( .B(clk), .A(\g.we_clk [20633]));
Q_ASSIGN U12142 ( .B(clk), .A(\g.we_clk [20632]));
Q_ASSIGN U12143 ( .B(clk), .A(\g.we_clk [20631]));
Q_ASSIGN U12144 ( .B(clk), .A(\g.we_clk [20630]));
Q_ASSIGN U12145 ( .B(clk), .A(\g.we_clk [20629]));
Q_ASSIGN U12146 ( .B(clk), .A(\g.we_clk [20628]));
Q_ASSIGN U12147 ( .B(clk), .A(\g.we_clk [20627]));
Q_ASSIGN U12148 ( .B(clk), .A(\g.we_clk [20626]));
Q_ASSIGN U12149 ( .B(clk), .A(\g.we_clk [20625]));
Q_ASSIGN U12150 ( .B(clk), .A(\g.we_clk [20624]));
Q_ASSIGN U12151 ( .B(clk), .A(\g.we_clk [20623]));
Q_ASSIGN U12152 ( .B(clk), .A(\g.we_clk [20622]));
Q_ASSIGN U12153 ( .B(clk), .A(\g.we_clk [20621]));
Q_ASSIGN U12154 ( .B(clk), .A(\g.we_clk [20620]));
Q_ASSIGN U12155 ( .B(clk), .A(\g.we_clk [20619]));
Q_ASSIGN U12156 ( .B(clk), .A(\g.we_clk [20618]));
Q_ASSIGN U12157 ( .B(clk), .A(\g.we_clk [20617]));
Q_ASSIGN U12158 ( .B(clk), .A(\g.we_clk [20616]));
Q_ASSIGN U12159 ( .B(clk), .A(\g.we_clk [20615]));
Q_ASSIGN U12160 ( .B(clk), .A(\g.we_clk [20614]));
Q_ASSIGN U12161 ( .B(clk), .A(\g.we_clk [20613]));
Q_ASSIGN U12162 ( .B(clk), .A(\g.we_clk [20612]));
Q_ASSIGN U12163 ( .B(clk), .A(\g.we_clk [20611]));
Q_ASSIGN U12164 ( .B(clk), .A(\g.we_clk [20610]));
Q_ASSIGN U12165 ( .B(clk), .A(\g.we_clk [20609]));
Q_ASSIGN U12166 ( .B(clk), .A(\g.we_clk [20608]));
Q_ASSIGN U12167 ( .B(clk), .A(\g.we_clk [20607]));
Q_ASSIGN U12168 ( .B(clk), .A(\g.we_clk [20606]));
Q_ASSIGN U12169 ( .B(clk), .A(\g.we_clk [20605]));
Q_ASSIGN U12170 ( .B(clk), .A(\g.we_clk [20604]));
Q_ASSIGN U12171 ( .B(clk), .A(\g.we_clk [20603]));
Q_ASSIGN U12172 ( .B(clk), .A(\g.we_clk [20602]));
Q_ASSIGN U12173 ( .B(clk), .A(\g.we_clk [20601]));
Q_ASSIGN U12174 ( .B(clk), .A(\g.we_clk [20600]));
Q_ASSIGN U12175 ( .B(clk), .A(\g.we_clk [20599]));
Q_ASSIGN U12176 ( .B(clk), .A(\g.we_clk [20598]));
Q_ASSIGN U12177 ( .B(clk), .A(\g.we_clk [20597]));
Q_ASSIGN U12178 ( .B(clk), .A(\g.we_clk [20596]));
Q_ASSIGN U12179 ( .B(clk), .A(\g.we_clk [20595]));
Q_ASSIGN U12180 ( .B(clk), .A(\g.we_clk [20594]));
Q_ASSIGN U12181 ( .B(clk), .A(\g.we_clk [20593]));
Q_ASSIGN U12182 ( .B(clk), .A(\g.we_clk [20592]));
Q_ASSIGN U12183 ( .B(clk), .A(\g.we_clk [20591]));
Q_ASSIGN U12184 ( .B(clk), .A(\g.we_clk [20590]));
Q_ASSIGN U12185 ( .B(clk), .A(\g.we_clk [20589]));
Q_ASSIGN U12186 ( .B(clk), .A(\g.we_clk [20588]));
Q_ASSIGN U12187 ( .B(clk), .A(\g.we_clk [20587]));
Q_ASSIGN U12188 ( .B(clk), .A(\g.we_clk [20586]));
Q_ASSIGN U12189 ( .B(clk), .A(\g.we_clk [20585]));
Q_ASSIGN U12190 ( .B(clk), .A(\g.we_clk [20584]));
Q_ASSIGN U12191 ( .B(clk), .A(\g.we_clk [20583]));
Q_ASSIGN U12192 ( .B(clk), .A(\g.we_clk [20582]));
Q_ASSIGN U12193 ( .B(clk), .A(\g.we_clk [20581]));
Q_ASSIGN U12194 ( .B(clk), .A(\g.we_clk [20580]));
Q_ASSIGN U12195 ( .B(clk), .A(\g.we_clk [20579]));
Q_ASSIGN U12196 ( .B(clk), .A(\g.we_clk [20578]));
Q_ASSIGN U12197 ( .B(clk), .A(\g.we_clk [20577]));
Q_ASSIGN U12198 ( .B(clk), .A(\g.we_clk [20576]));
Q_ASSIGN U12199 ( .B(clk), .A(\g.we_clk [20575]));
Q_ASSIGN U12200 ( .B(clk), .A(\g.we_clk [20574]));
Q_ASSIGN U12201 ( .B(clk), .A(\g.we_clk [20573]));
Q_ASSIGN U12202 ( .B(clk), .A(\g.we_clk [20572]));
Q_ASSIGN U12203 ( .B(clk), .A(\g.we_clk [20571]));
Q_ASSIGN U12204 ( .B(clk), .A(\g.we_clk [20570]));
Q_ASSIGN U12205 ( .B(clk), .A(\g.we_clk [20569]));
Q_ASSIGN U12206 ( .B(clk), .A(\g.we_clk [20568]));
Q_ASSIGN U12207 ( .B(clk), .A(\g.we_clk [20567]));
Q_ASSIGN U12208 ( .B(clk), .A(\g.we_clk [20566]));
Q_ASSIGN U12209 ( .B(clk), .A(\g.we_clk [20565]));
Q_ASSIGN U12210 ( .B(clk), .A(\g.we_clk [20564]));
Q_ASSIGN U12211 ( .B(clk), .A(\g.we_clk [20563]));
Q_ASSIGN U12212 ( .B(clk), .A(\g.we_clk [20562]));
Q_ASSIGN U12213 ( .B(clk), .A(\g.we_clk [20561]));
Q_ASSIGN U12214 ( .B(clk), .A(\g.we_clk [20560]));
Q_ASSIGN U12215 ( .B(clk), .A(\g.we_clk [20559]));
Q_ASSIGN U12216 ( .B(clk), .A(\g.we_clk [20558]));
Q_ASSIGN U12217 ( .B(clk), .A(\g.we_clk [20557]));
Q_ASSIGN U12218 ( .B(clk), .A(\g.we_clk [20556]));
Q_ASSIGN U12219 ( .B(clk), .A(\g.we_clk [20555]));
Q_ASSIGN U12220 ( .B(clk), .A(\g.we_clk [20554]));
Q_ASSIGN U12221 ( .B(clk), .A(\g.we_clk [20553]));
Q_ASSIGN U12222 ( .B(clk), .A(\g.we_clk [20552]));
Q_ASSIGN U12223 ( .B(clk), .A(\g.we_clk [20551]));
Q_ASSIGN U12224 ( .B(clk), .A(\g.we_clk [20550]));
Q_ASSIGN U12225 ( .B(clk), .A(\g.we_clk [20549]));
Q_ASSIGN U12226 ( .B(clk), .A(\g.we_clk [20548]));
Q_ASSIGN U12227 ( .B(clk), .A(\g.we_clk [20547]));
Q_ASSIGN U12228 ( .B(clk), .A(\g.we_clk [20546]));
Q_ASSIGN U12229 ( .B(clk), .A(\g.we_clk [20545]));
Q_ASSIGN U12230 ( .B(clk), .A(\g.we_clk [20544]));
Q_ASSIGN U12231 ( .B(clk), .A(\g.we_clk [20543]));
Q_ASSIGN U12232 ( .B(clk), .A(\g.we_clk [20542]));
Q_ASSIGN U12233 ( .B(clk), .A(\g.we_clk [20541]));
Q_ASSIGN U12234 ( .B(clk), .A(\g.we_clk [20540]));
Q_ASSIGN U12235 ( .B(clk), .A(\g.we_clk [20539]));
Q_ASSIGN U12236 ( .B(clk), .A(\g.we_clk [20538]));
Q_ASSIGN U12237 ( .B(clk), .A(\g.we_clk [20537]));
Q_ASSIGN U12238 ( .B(clk), .A(\g.we_clk [20536]));
Q_ASSIGN U12239 ( .B(clk), .A(\g.we_clk [20535]));
Q_ASSIGN U12240 ( .B(clk), .A(\g.we_clk [20534]));
Q_ASSIGN U12241 ( .B(clk), .A(\g.we_clk [20533]));
Q_ASSIGN U12242 ( .B(clk), .A(\g.we_clk [20532]));
Q_ASSIGN U12243 ( .B(clk), .A(\g.we_clk [20531]));
Q_ASSIGN U12244 ( .B(clk), .A(\g.we_clk [20530]));
Q_ASSIGN U12245 ( .B(clk), .A(\g.we_clk [20529]));
Q_ASSIGN U12246 ( .B(clk), .A(\g.we_clk [20528]));
Q_ASSIGN U12247 ( .B(clk), .A(\g.we_clk [20527]));
Q_ASSIGN U12248 ( .B(clk), .A(\g.we_clk [20526]));
Q_ASSIGN U12249 ( .B(clk), .A(\g.we_clk [20525]));
Q_ASSIGN U12250 ( .B(clk), .A(\g.we_clk [20524]));
Q_ASSIGN U12251 ( .B(clk), .A(\g.we_clk [20523]));
Q_ASSIGN U12252 ( .B(clk), .A(\g.we_clk [20522]));
Q_ASSIGN U12253 ( .B(clk), .A(\g.we_clk [20521]));
Q_ASSIGN U12254 ( .B(clk), .A(\g.we_clk [20520]));
Q_ASSIGN U12255 ( .B(clk), .A(\g.we_clk [20519]));
Q_ASSIGN U12256 ( .B(clk), .A(\g.we_clk [20518]));
Q_ASSIGN U12257 ( .B(clk), .A(\g.we_clk [20517]));
Q_ASSIGN U12258 ( .B(clk), .A(\g.we_clk [20516]));
Q_ASSIGN U12259 ( .B(clk), .A(\g.we_clk [20515]));
Q_ASSIGN U12260 ( .B(clk), .A(\g.we_clk [20514]));
Q_ASSIGN U12261 ( .B(clk), .A(\g.we_clk [20513]));
Q_ASSIGN U12262 ( .B(clk), .A(\g.we_clk [20512]));
Q_ASSIGN U12263 ( .B(clk), .A(\g.we_clk [20511]));
Q_ASSIGN U12264 ( .B(clk), .A(\g.we_clk [20510]));
Q_ASSIGN U12265 ( .B(clk), .A(\g.we_clk [20509]));
Q_ASSIGN U12266 ( .B(clk), .A(\g.we_clk [20508]));
Q_ASSIGN U12267 ( .B(clk), .A(\g.we_clk [20507]));
Q_ASSIGN U12268 ( .B(clk), .A(\g.we_clk [20506]));
Q_ASSIGN U12269 ( .B(clk), .A(\g.we_clk [20505]));
Q_ASSIGN U12270 ( .B(clk), .A(\g.we_clk [20504]));
Q_ASSIGN U12271 ( .B(clk), .A(\g.we_clk [20503]));
Q_ASSIGN U12272 ( .B(clk), .A(\g.we_clk [20502]));
Q_ASSIGN U12273 ( .B(clk), .A(\g.we_clk [20501]));
Q_ASSIGN U12274 ( .B(clk), .A(\g.we_clk [20500]));
Q_ASSIGN U12275 ( .B(clk), .A(\g.we_clk [20499]));
Q_ASSIGN U12276 ( .B(clk), .A(\g.we_clk [20498]));
Q_ASSIGN U12277 ( .B(clk), .A(\g.we_clk [20497]));
Q_ASSIGN U12278 ( .B(clk), .A(\g.we_clk [20496]));
Q_ASSIGN U12279 ( .B(clk), .A(\g.we_clk [20495]));
Q_ASSIGN U12280 ( .B(clk), .A(\g.we_clk [20494]));
Q_ASSIGN U12281 ( .B(clk), .A(\g.we_clk [20493]));
Q_ASSIGN U12282 ( .B(clk), .A(\g.we_clk [20492]));
Q_ASSIGN U12283 ( .B(clk), .A(\g.we_clk [20491]));
Q_ASSIGN U12284 ( .B(clk), .A(\g.we_clk [20490]));
Q_ASSIGN U12285 ( .B(clk), .A(\g.we_clk [20489]));
Q_ASSIGN U12286 ( .B(clk), .A(\g.we_clk [20488]));
Q_ASSIGN U12287 ( .B(clk), .A(\g.we_clk [20487]));
Q_ASSIGN U12288 ( .B(clk), .A(\g.we_clk [20486]));
Q_ASSIGN U12289 ( .B(clk), .A(\g.we_clk [20485]));
Q_ASSIGN U12290 ( .B(clk), .A(\g.we_clk [20484]));
Q_ASSIGN U12291 ( .B(clk), .A(\g.we_clk [20483]));
Q_ASSIGN U12292 ( .B(clk), .A(\g.we_clk [20482]));
Q_ASSIGN U12293 ( .B(clk), .A(\g.we_clk [20481]));
Q_ASSIGN U12294 ( .B(clk), .A(\g.we_clk [20480]));
Q_ASSIGN U12295 ( .B(clk), .A(\g.we_clk [20479]));
Q_ASSIGN U12296 ( .B(clk), .A(\g.we_clk [20478]));
Q_ASSIGN U12297 ( .B(clk), .A(\g.we_clk [20477]));
Q_ASSIGN U12298 ( .B(clk), .A(\g.we_clk [20476]));
Q_ASSIGN U12299 ( .B(clk), .A(\g.we_clk [20475]));
Q_ASSIGN U12300 ( .B(clk), .A(\g.we_clk [20474]));
Q_ASSIGN U12301 ( .B(clk), .A(\g.we_clk [20473]));
Q_ASSIGN U12302 ( .B(clk), .A(\g.we_clk [20472]));
Q_ASSIGN U12303 ( .B(clk), .A(\g.we_clk [20471]));
Q_ASSIGN U12304 ( .B(clk), .A(\g.we_clk [20470]));
Q_ASSIGN U12305 ( .B(clk), .A(\g.we_clk [20469]));
Q_ASSIGN U12306 ( .B(clk), .A(\g.we_clk [20468]));
Q_ASSIGN U12307 ( .B(clk), .A(\g.we_clk [20467]));
Q_ASSIGN U12308 ( .B(clk), .A(\g.we_clk [20466]));
Q_ASSIGN U12309 ( .B(clk), .A(\g.we_clk [20465]));
Q_ASSIGN U12310 ( .B(clk), .A(\g.we_clk [20464]));
Q_ASSIGN U12311 ( .B(clk), .A(\g.we_clk [20463]));
Q_ASSIGN U12312 ( .B(clk), .A(\g.we_clk [20462]));
Q_ASSIGN U12313 ( .B(clk), .A(\g.we_clk [20461]));
Q_ASSIGN U12314 ( .B(clk), .A(\g.we_clk [20460]));
Q_ASSIGN U12315 ( .B(clk), .A(\g.we_clk [20459]));
Q_ASSIGN U12316 ( .B(clk), .A(\g.we_clk [20458]));
Q_ASSIGN U12317 ( .B(clk), .A(\g.we_clk [20457]));
Q_ASSIGN U12318 ( .B(clk), .A(\g.we_clk [20456]));
Q_ASSIGN U12319 ( .B(clk), .A(\g.we_clk [20455]));
Q_ASSIGN U12320 ( .B(clk), .A(\g.we_clk [20454]));
Q_ASSIGN U12321 ( .B(clk), .A(\g.we_clk [20453]));
Q_ASSIGN U12322 ( .B(clk), .A(\g.we_clk [20452]));
Q_ASSIGN U12323 ( .B(clk), .A(\g.we_clk [20451]));
Q_ASSIGN U12324 ( .B(clk), .A(\g.we_clk [20450]));
Q_ASSIGN U12325 ( .B(clk), .A(\g.we_clk [20449]));
Q_ASSIGN U12326 ( .B(clk), .A(\g.we_clk [20448]));
Q_ASSIGN U12327 ( .B(clk), .A(\g.we_clk [20447]));
Q_ASSIGN U12328 ( .B(clk), .A(\g.we_clk [20446]));
Q_ASSIGN U12329 ( .B(clk), .A(\g.we_clk [20445]));
Q_ASSIGN U12330 ( .B(clk), .A(\g.we_clk [20444]));
Q_ASSIGN U12331 ( .B(clk), .A(\g.we_clk [20443]));
Q_ASSIGN U12332 ( .B(clk), .A(\g.we_clk [20442]));
Q_ASSIGN U12333 ( .B(clk), .A(\g.we_clk [20441]));
Q_ASSIGN U12334 ( .B(clk), .A(\g.we_clk [20440]));
Q_ASSIGN U12335 ( .B(clk), .A(\g.we_clk [20439]));
Q_ASSIGN U12336 ( .B(clk), .A(\g.we_clk [20438]));
Q_ASSIGN U12337 ( .B(clk), .A(\g.we_clk [20437]));
Q_ASSIGN U12338 ( .B(clk), .A(\g.we_clk [20436]));
Q_ASSIGN U12339 ( .B(clk), .A(\g.we_clk [20435]));
Q_ASSIGN U12340 ( .B(clk), .A(\g.we_clk [20434]));
Q_ASSIGN U12341 ( .B(clk), .A(\g.we_clk [20433]));
Q_ASSIGN U12342 ( .B(clk), .A(\g.we_clk [20432]));
Q_ASSIGN U12343 ( .B(clk), .A(\g.we_clk [20431]));
Q_ASSIGN U12344 ( .B(clk), .A(\g.we_clk [20430]));
Q_ASSIGN U12345 ( .B(clk), .A(\g.we_clk [20429]));
Q_ASSIGN U12346 ( .B(clk), .A(\g.we_clk [20428]));
Q_ASSIGN U12347 ( .B(clk), .A(\g.we_clk [20427]));
Q_ASSIGN U12348 ( .B(clk), .A(\g.we_clk [20426]));
Q_ASSIGN U12349 ( .B(clk), .A(\g.we_clk [20425]));
Q_ASSIGN U12350 ( .B(clk), .A(\g.we_clk [20424]));
Q_ASSIGN U12351 ( .B(clk), .A(\g.we_clk [20423]));
Q_ASSIGN U12352 ( .B(clk), .A(\g.we_clk [20422]));
Q_ASSIGN U12353 ( .B(clk), .A(\g.we_clk [20421]));
Q_ASSIGN U12354 ( .B(clk), .A(\g.we_clk [20420]));
Q_ASSIGN U12355 ( .B(clk), .A(\g.we_clk [20419]));
Q_ASSIGN U12356 ( .B(clk), .A(\g.we_clk [20418]));
Q_ASSIGN U12357 ( .B(clk), .A(\g.we_clk [20417]));
Q_ASSIGN U12358 ( .B(clk), .A(\g.we_clk [20416]));
Q_ASSIGN U12359 ( .B(clk), .A(\g.we_clk [20415]));
Q_ASSIGN U12360 ( .B(clk), .A(\g.we_clk [20414]));
Q_ASSIGN U12361 ( .B(clk), .A(\g.we_clk [20413]));
Q_ASSIGN U12362 ( .B(clk), .A(\g.we_clk [20412]));
Q_ASSIGN U12363 ( .B(clk), .A(\g.we_clk [20411]));
Q_ASSIGN U12364 ( .B(clk), .A(\g.we_clk [20410]));
Q_ASSIGN U12365 ( .B(clk), .A(\g.we_clk [20409]));
Q_ASSIGN U12366 ( .B(clk), .A(\g.we_clk [20408]));
Q_ASSIGN U12367 ( .B(clk), .A(\g.we_clk [20407]));
Q_ASSIGN U12368 ( .B(clk), .A(\g.we_clk [20406]));
Q_ASSIGN U12369 ( .B(clk), .A(\g.we_clk [20405]));
Q_ASSIGN U12370 ( .B(clk), .A(\g.we_clk [20404]));
Q_ASSIGN U12371 ( .B(clk), .A(\g.we_clk [20403]));
Q_ASSIGN U12372 ( .B(clk), .A(\g.we_clk [20402]));
Q_ASSIGN U12373 ( .B(clk), .A(\g.we_clk [20401]));
Q_ASSIGN U12374 ( .B(clk), .A(\g.we_clk [20400]));
Q_ASSIGN U12375 ( .B(clk), .A(\g.we_clk [20399]));
Q_ASSIGN U12376 ( .B(clk), .A(\g.we_clk [20398]));
Q_ASSIGN U12377 ( .B(clk), .A(\g.we_clk [20397]));
Q_ASSIGN U12378 ( .B(clk), .A(\g.we_clk [20396]));
Q_ASSIGN U12379 ( .B(clk), .A(\g.we_clk [20395]));
Q_ASSIGN U12380 ( .B(clk), .A(\g.we_clk [20394]));
Q_ASSIGN U12381 ( .B(clk), .A(\g.we_clk [20393]));
Q_ASSIGN U12382 ( .B(clk), .A(\g.we_clk [20392]));
Q_ASSIGN U12383 ( .B(clk), .A(\g.we_clk [20391]));
Q_ASSIGN U12384 ( .B(clk), .A(\g.we_clk [20390]));
Q_ASSIGN U12385 ( .B(clk), .A(\g.we_clk [20389]));
Q_ASSIGN U12386 ( .B(clk), .A(\g.we_clk [20388]));
Q_ASSIGN U12387 ( .B(clk), .A(\g.we_clk [20387]));
Q_ASSIGN U12388 ( .B(clk), .A(\g.we_clk [20386]));
Q_ASSIGN U12389 ( .B(clk), .A(\g.we_clk [20385]));
Q_ASSIGN U12390 ( .B(clk), .A(\g.we_clk [20384]));
Q_ASSIGN U12391 ( .B(clk), .A(\g.we_clk [20383]));
Q_ASSIGN U12392 ( .B(clk), .A(\g.we_clk [20382]));
Q_ASSIGN U12393 ( .B(clk), .A(\g.we_clk [20381]));
Q_ASSIGN U12394 ( .B(clk), .A(\g.we_clk [20380]));
Q_ASSIGN U12395 ( .B(clk), .A(\g.we_clk [20379]));
Q_ASSIGN U12396 ( .B(clk), .A(\g.we_clk [20378]));
Q_ASSIGN U12397 ( .B(clk), .A(\g.we_clk [20377]));
Q_ASSIGN U12398 ( .B(clk), .A(\g.we_clk [20376]));
Q_ASSIGN U12399 ( .B(clk), .A(\g.we_clk [20375]));
Q_ASSIGN U12400 ( .B(clk), .A(\g.we_clk [20374]));
Q_ASSIGN U12401 ( .B(clk), .A(\g.we_clk [20373]));
Q_ASSIGN U12402 ( .B(clk), .A(\g.we_clk [20372]));
Q_ASSIGN U12403 ( .B(clk), .A(\g.we_clk [20371]));
Q_ASSIGN U12404 ( .B(clk), .A(\g.we_clk [20370]));
Q_ASSIGN U12405 ( .B(clk), .A(\g.we_clk [20369]));
Q_ASSIGN U12406 ( .B(clk), .A(\g.we_clk [20368]));
Q_ASSIGN U12407 ( .B(clk), .A(\g.we_clk [20367]));
Q_ASSIGN U12408 ( .B(clk), .A(\g.we_clk [20366]));
Q_ASSIGN U12409 ( .B(clk), .A(\g.we_clk [20365]));
Q_ASSIGN U12410 ( .B(clk), .A(\g.we_clk [20364]));
Q_ASSIGN U12411 ( .B(clk), .A(\g.we_clk [20363]));
Q_ASSIGN U12412 ( .B(clk), .A(\g.we_clk [20362]));
Q_ASSIGN U12413 ( .B(clk), .A(\g.we_clk [20361]));
Q_ASSIGN U12414 ( .B(clk), .A(\g.we_clk [20360]));
Q_ASSIGN U12415 ( .B(clk), .A(\g.we_clk [20359]));
Q_ASSIGN U12416 ( .B(clk), .A(\g.we_clk [20358]));
Q_ASSIGN U12417 ( .B(clk), .A(\g.we_clk [20357]));
Q_ASSIGN U12418 ( .B(clk), .A(\g.we_clk [20356]));
Q_ASSIGN U12419 ( .B(clk), .A(\g.we_clk [20355]));
Q_ASSIGN U12420 ( .B(clk), .A(\g.we_clk [20354]));
Q_ASSIGN U12421 ( .B(clk), .A(\g.we_clk [20353]));
Q_ASSIGN U12422 ( .B(clk), .A(\g.we_clk [20352]));
Q_ASSIGN U12423 ( .B(clk), .A(\g.we_clk [20351]));
Q_ASSIGN U12424 ( .B(clk), .A(\g.we_clk [20350]));
Q_ASSIGN U12425 ( .B(clk), .A(\g.we_clk [20349]));
Q_ASSIGN U12426 ( .B(clk), .A(\g.we_clk [20348]));
Q_ASSIGN U12427 ( .B(clk), .A(\g.we_clk [20347]));
Q_ASSIGN U12428 ( .B(clk), .A(\g.we_clk [20346]));
Q_ASSIGN U12429 ( .B(clk), .A(\g.we_clk [20345]));
Q_ASSIGN U12430 ( .B(clk), .A(\g.we_clk [20344]));
Q_ASSIGN U12431 ( .B(clk), .A(\g.we_clk [20343]));
Q_ASSIGN U12432 ( .B(clk), .A(\g.we_clk [20342]));
Q_ASSIGN U12433 ( .B(clk), .A(\g.we_clk [20341]));
Q_ASSIGN U12434 ( .B(clk), .A(\g.we_clk [20340]));
Q_ASSIGN U12435 ( .B(clk), .A(\g.we_clk [20339]));
Q_ASSIGN U12436 ( .B(clk), .A(\g.we_clk [20338]));
Q_ASSIGN U12437 ( .B(clk), .A(\g.we_clk [20337]));
Q_ASSIGN U12438 ( .B(clk), .A(\g.we_clk [20336]));
Q_ASSIGN U12439 ( .B(clk), .A(\g.we_clk [20335]));
Q_ASSIGN U12440 ( .B(clk), .A(\g.we_clk [20334]));
Q_ASSIGN U12441 ( .B(clk), .A(\g.we_clk [20333]));
Q_ASSIGN U12442 ( .B(clk), .A(\g.we_clk [20332]));
Q_ASSIGN U12443 ( .B(clk), .A(\g.we_clk [20331]));
Q_ASSIGN U12444 ( .B(clk), .A(\g.we_clk [20330]));
Q_ASSIGN U12445 ( .B(clk), .A(\g.we_clk [20329]));
Q_ASSIGN U12446 ( .B(clk), .A(\g.we_clk [20328]));
Q_ASSIGN U12447 ( .B(clk), .A(\g.we_clk [20327]));
Q_ASSIGN U12448 ( .B(clk), .A(\g.we_clk [20326]));
Q_ASSIGN U12449 ( .B(clk), .A(\g.we_clk [20325]));
Q_ASSIGN U12450 ( .B(clk), .A(\g.we_clk [20324]));
Q_ASSIGN U12451 ( .B(clk), .A(\g.we_clk [20323]));
Q_ASSIGN U12452 ( .B(clk), .A(\g.we_clk [20322]));
Q_ASSIGN U12453 ( .B(clk), .A(\g.we_clk [20321]));
Q_ASSIGN U12454 ( .B(clk), .A(\g.we_clk [20320]));
Q_ASSIGN U12455 ( .B(clk), .A(\g.we_clk [20319]));
Q_ASSIGN U12456 ( .B(clk), .A(\g.we_clk [20318]));
Q_ASSIGN U12457 ( .B(clk), .A(\g.we_clk [20317]));
Q_ASSIGN U12458 ( .B(clk), .A(\g.we_clk [20316]));
Q_ASSIGN U12459 ( .B(clk), .A(\g.we_clk [20315]));
Q_ASSIGN U12460 ( .B(clk), .A(\g.we_clk [20314]));
Q_ASSIGN U12461 ( .B(clk), .A(\g.we_clk [20313]));
Q_ASSIGN U12462 ( .B(clk), .A(\g.we_clk [20312]));
Q_ASSIGN U12463 ( .B(clk), .A(\g.we_clk [20311]));
Q_ASSIGN U12464 ( .B(clk), .A(\g.we_clk [20310]));
Q_ASSIGN U12465 ( .B(clk), .A(\g.we_clk [20309]));
Q_ASSIGN U12466 ( .B(clk), .A(\g.we_clk [20308]));
Q_ASSIGN U12467 ( .B(clk), .A(\g.we_clk [20307]));
Q_ASSIGN U12468 ( .B(clk), .A(\g.we_clk [20306]));
Q_ASSIGN U12469 ( .B(clk), .A(\g.we_clk [20305]));
Q_ASSIGN U12470 ( .B(clk), .A(\g.we_clk [20304]));
Q_ASSIGN U12471 ( .B(clk), .A(\g.we_clk [20303]));
Q_ASSIGN U12472 ( .B(clk), .A(\g.we_clk [20302]));
Q_ASSIGN U12473 ( .B(clk), .A(\g.we_clk [20301]));
Q_ASSIGN U12474 ( .B(clk), .A(\g.we_clk [20300]));
Q_ASSIGN U12475 ( .B(clk), .A(\g.we_clk [20299]));
Q_ASSIGN U12476 ( .B(clk), .A(\g.we_clk [20298]));
Q_ASSIGN U12477 ( .B(clk), .A(\g.we_clk [20297]));
Q_ASSIGN U12478 ( .B(clk), .A(\g.we_clk [20296]));
Q_ASSIGN U12479 ( .B(clk), .A(\g.we_clk [20295]));
Q_ASSIGN U12480 ( .B(clk), .A(\g.we_clk [20294]));
Q_ASSIGN U12481 ( .B(clk), .A(\g.we_clk [20293]));
Q_ASSIGN U12482 ( .B(clk), .A(\g.we_clk [20292]));
Q_ASSIGN U12483 ( .B(clk), .A(\g.we_clk [20291]));
Q_ASSIGN U12484 ( .B(clk), .A(\g.we_clk [20290]));
Q_ASSIGN U12485 ( .B(clk), .A(\g.we_clk [20289]));
Q_ASSIGN U12486 ( .B(clk), .A(\g.we_clk [20288]));
Q_ASSIGN U12487 ( .B(clk), .A(\g.we_clk [20287]));
Q_ASSIGN U12488 ( .B(clk), .A(\g.we_clk [20286]));
Q_ASSIGN U12489 ( .B(clk), .A(\g.we_clk [20285]));
Q_ASSIGN U12490 ( .B(clk), .A(\g.we_clk [20284]));
Q_ASSIGN U12491 ( .B(clk), .A(\g.we_clk [20283]));
Q_ASSIGN U12492 ( .B(clk), .A(\g.we_clk [20282]));
Q_ASSIGN U12493 ( .B(clk), .A(\g.we_clk [20281]));
Q_ASSIGN U12494 ( .B(clk), .A(\g.we_clk [20280]));
Q_ASSIGN U12495 ( .B(clk), .A(\g.we_clk [20279]));
Q_ASSIGN U12496 ( .B(clk), .A(\g.we_clk [20278]));
Q_ASSIGN U12497 ( .B(clk), .A(\g.we_clk [20277]));
Q_ASSIGN U12498 ( .B(clk), .A(\g.we_clk [20276]));
Q_ASSIGN U12499 ( .B(clk), .A(\g.we_clk [20275]));
Q_ASSIGN U12500 ( .B(clk), .A(\g.we_clk [20274]));
Q_ASSIGN U12501 ( .B(clk), .A(\g.we_clk [20273]));
Q_ASSIGN U12502 ( .B(clk), .A(\g.we_clk [20272]));
Q_ASSIGN U12503 ( .B(clk), .A(\g.we_clk [20271]));
Q_ASSIGN U12504 ( .B(clk), .A(\g.we_clk [20270]));
Q_ASSIGN U12505 ( .B(clk), .A(\g.we_clk [20269]));
Q_ASSIGN U12506 ( .B(clk), .A(\g.we_clk [20268]));
Q_ASSIGN U12507 ( .B(clk), .A(\g.we_clk [20267]));
Q_ASSIGN U12508 ( .B(clk), .A(\g.we_clk [20266]));
Q_ASSIGN U12509 ( .B(clk), .A(\g.we_clk [20265]));
Q_ASSIGN U12510 ( .B(clk), .A(\g.we_clk [20264]));
Q_ASSIGN U12511 ( .B(clk), .A(\g.we_clk [20263]));
Q_ASSIGN U12512 ( .B(clk), .A(\g.we_clk [20262]));
Q_ASSIGN U12513 ( .B(clk), .A(\g.we_clk [20261]));
Q_ASSIGN U12514 ( .B(clk), .A(\g.we_clk [20260]));
Q_ASSIGN U12515 ( .B(clk), .A(\g.we_clk [20259]));
Q_ASSIGN U12516 ( .B(clk), .A(\g.we_clk [20258]));
Q_ASSIGN U12517 ( .B(clk), .A(\g.we_clk [20257]));
Q_ASSIGN U12518 ( .B(clk), .A(\g.we_clk [20256]));
Q_ASSIGN U12519 ( .B(clk), .A(\g.we_clk [20255]));
Q_ASSIGN U12520 ( .B(clk), .A(\g.we_clk [20254]));
Q_ASSIGN U12521 ( .B(clk), .A(\g.we_clk [20253]));
Q_ASSIGN U12522 ( .B(clk), .A(\g.we_clk [20252]));
Q_ASSIGN U12523 ( .B(clk), .A(\g.we_clk [20251]));
Q_ASSIGN U12524 ( .B(clk), .A(\g.we_clk [20250]));
Q_ASSIGN U12525 ( .B(clk), .A(\g.we_clk [20249]));
Q_ASSIGN U12526 ( .B(clk), .A(\g.we_clk [20248]));
Q_ASSIGN U12527 ( .B(clk), .A(\g.we_clk [20247]));
Q_ASSIGN U12528 ( .B(clk), .A(\g.we_clk [20246]));
Q_ASSIGN U12529 ( .B(clk), .A(\g.we_clk [20245]));
Q_ASSIGN U12530 ( .B(clk), .A(\g.we_clk [20244]));
Q_ASSIGN U12531 ( .B(clk), .A(\g.we_clk [20243]));
Q_ASSIGN U12532 ( .B(clk), .A(\g.we_clk [20242]));
Q_ASSIGN U12533 ( .B(clk), .A(\g.we_clk [20241]));
Q_ASSIGN U12534 ( .B(clk), .A(\g.we_clk [20240]));
Q_ASSIGN U12535 ( .B(clk), .A(\g.we_clk [20239]));
Q_ASSIGN U12536 ( .B(clk), .A(\g.we_clk [20238]));
Q_ASSIGN U12537 ( .B(clk), .A(\g.we_clk [20237]));
Q_ASSIGN U12538 ( .B(clk), .A(\g.we_clk [20236]));
Q_ASSIGN U12539 ( .B(clk), .A(\g.we_clk [20235]));
Q_ASSIGN U12540 ( .B(clk), .A(\g.we_clk [20234]));
Q_ASSIGN U12541 ( .B(clk), .A(\g.we_clk [20233]));
Q_ASSIGN U12542 ( .B(clk), .A(\g.we_clk [20232]));
Q_ASSIGN U12543 ( .B(clk), .A(\g.we_clk [20231]));
Q_ASSIGN U12544 ( .B(clk), .A(\g.we_clk [20230]));
Q_ASSIGN U12545 ( .B(clk), .A(\g.we_clk [20229]));
Q_ASSIGN U12546 ( .B(clk), .A(\g.we_clk [20228]));
Q_ASSIGN U12547 ( .B(clk), .A(\g.we_clk [20227]));
Q_ASSIGN U12548 ( .B(clk), .A(\g.we_clk [20226]));
Q_ASSIGN U12549 ( .B(clk), .A(\g.we_clk [20225]));
Q_ASSIGN U12550 ( .B(clk), .A(\g.we_clk [20224]));
Q_ASSIGN U12551 ( .B(clk), .A(\g.we_clk [20223]));
Q_ASSIGN U12552 ( .B(clk), .A(\g.we_clk [20222]));
Q_ASSIGN U12553 ( .B(clk), .A(\g.we_clk [20221]));
Q_ASSIGN U12554 ( .B(clk), .A(\g.we_clk [20220]));
Q_ASSIGN U12555 ( .B(clk), .A(\g.we_clk [20219]));
Q_ASSIGN U12556 ( .B(clk), .A(\g.we_clk [20218]));
Q_ASSIGN U12557 ( .B(clk), .A(\g.we_clk [20217]));
Q_ASSIGN U12558 ( .B(clk), .A(\g.we_clk [20216]));
Q_ASSIGN U12559 ( .B(clk), .A(\g.we_clk [20215]));
Q_ASSIGN U12560 ( .B(clk), .A(\g.we_clk [20214]));
Q_ASSIGN U12561 ( .B(clk), .A(\g.we_clk [20213]));
Q_ASSIGN U12562 ( .B(clk), .A(\g.we_clk [20212]));
Q_ASSIGN U12563 ( .B(clk), .A(\g.we_clk [20211]));
Q_ASSIGN U12564 ( .B(clk), .A(\g.we_clk [20210]));
Q_ASSIGN U12565 ( .B(clk), .A(\g.we_clk [20209]));
Q_ASSIGN U12566 ( .B(clk), .A(\g.we_clk [20208]));
Q_ASSIGN U12567 ( .B(clk), .A(\g.we_clk [20207]));
Q_ASSIGN U12568 ( .B(clk), .A(\g.we_clk [20206]));
Q_ASSIGN U12569 ( .B(clk), .A(\g.we_clk [20205]));
Q_ASSIGN U12570 ( .B(clk), .A(\g.we_clk [20204]));
Q_ASSIGN U12571 ( .B(clk), .A(\g.we_clk [20203]));
Q_ASSIGN U12572 ( .B(clk), .A(\g.we_clk [20202]));
Q_ASSIGN U12573 ( .B(clk), .A(\g.we_clk [20201]));
Q_ASSIGN U12574 ( .B(clk), .A(\g.we_clk [20200]));
Q_ASSIGN U12575 ( .B(clk), .A(\g.we_clk [20199]));
Q_ASSIGN U12576 ( .B(clk), .A(\g.we_clk [20198]));
Q_ASSIGN U12577 ( .B(clk), .A(\g.we_clk [20197]));
Q_ASSIGN U12578 ( .B(clk), .A(\g.we_clk [20196]));
Q_ASSIGN U12579 ( .B(clk), .A(\g.we_clk [20195]));
Q_ASSIGN U12580 ( .B(clk), .A(\g.we_clk [20194]));
Q_ASSIGN U12581 ( .B(clk), .A(\g.we_clk [20193]));
Q_ASSIGN U12582 ( .B(clk), .A(\g.we_clk [20192]));
Q_ASSIGN U12583 ( .B(clk), .A(\g.we_clk [20191]));
Q_ASSIGN U12584 ( .B(clk), .A(\g.we_clk [20190]));
Q_ASSIGN U12585 ( .B(clk), .A(\g.we_clk [20189]));
Q_ASSIGN U12586 ( .B(clk), .A(\g.we_clk [20188]));
Q_ASSIGN U12587 ( .B(clk), .A(\g.we_clk [20187]));
Q_ASSIGN U12588 ( .B(clk), .A(\g.we_clk [20186]));
Q_ASSIGN U12589 ( .B(clk), .A(\g.we_clk [20185]));
Q_ASSIGN U12590 ( .B(clk), .A(\g.we_clk [20184]));
Q_ASSIGN U12591 ( .B(clk), .A(\g.we_clk [20183]));
Q_ASSIGN U12592 ( .B(clk), .A(\g.we_clk [20182]));
Q_ASSIGN U12593 ( .B(clk), .A(\g.we_clk [20181]));
Q_ASSIGN U12594 ( .B(clk), .A(\g.we_clk [20180]));
Q_ASSIGN U12595 ( .B(clk), .A(\g.we_clk [20179]));
Q_ASSIGN U12596 ( .B(clk), .A(\g.we_clk [20178]));
Q_ASSIGN U12597 ( .B(clk), .A(\g.we_clk [20177]));
Q_ASSIGN U12598 ( .B(clk), .A(\g.we_clk [20176]));
Q_ASSIGN U12599 ( .B(clk), .A(\g.we_clk [20175]));
Q_ASSIGN U12600 ( .B(clk), .A(\g.we_clk [20174]));
Q_ASSIGN U12601 ( .B(clk), .A(\g.we_clk [20173]));
Q_ASSIGN U12602 ( .B(clk), .A(\g.we_clk [20172]));
Q_ASSIGN U12603 ( .B(clk), .A(\g.we_clk [20171]));
Q_ASSIGN U12604 ( .B(clk), .A(\g.we_clk [20170]));
Q_ASSIGN U12605 ( .B(clk), .A(\g.we_clk [20169]));
Q_ASSIGN U12606 ( .B(clk), .A(\g.we_clk [20168]));
Q_ASSIGN U12607 ( .B(clk), .A(\g.we_clk [20167]));
Q_ASSIGN U12608 ( .B(clk), .A(\g.we_clk [20166]));
Q_ASSIGN U12609 ( .B(clk), .A(\g.we_clk [20165]));
Q_ASSIGN U12610 ( .B(clk), .A(\g.we_clk [20164]));
Q_ASSIGN U12611 ( .B(clk), .A(\g.we_clk [20163]));
Q_ASSIGN U12612 ( .B(clk), .A(\g.we_clk [20162]));
Q_ASSIGN U12613 ( .B(clk), .A(\g.we_clk [20161]));
Q_ASSIGN U12614 ( .B(clk), .A(\g.we_clk [20160]));
Q_ASSIGN U12615 ( .B(clk), .A(\g.we_clk [20159]));
Q_ASSIGN U12616 ( .B(clk), .A(\g.we_clk [20158]));
Q_ASSIGN U12617 ( .B(clk), .A(\g.we_clk [20157]));
Q_ASSIGN U12618 ( .B(clk), .A(\g.we_clk [20156]));
Q_ASSIGN U12619 ( .B(clk), .A(\g.we_clk [20155]));
Q_ASSIGN U12620 ( .B(clk), .A(\g.we_clk [20154]));
Q_ASSIGN U12621 ( .B(clk), .A(\g.we_clk [20153]));
Q_ASSIGN U12622 ( .B(clk), .A(\g.we_clk [20152]));
Q_ASSIGN U12623 ( .B(clk), .A(\g.we_clk [20151]));
Q_ASSIGN U12624 ( .B(clk), .A(\g.we_clk [20150]));
Q_ASSIGN U12625 ( .B(clk), .A(\g.we_clk [20149]));
Q_ASSIGN U12626 ( .B(clk), .A(\g.we_clk [20148]));
Q_ASSIGN U12627 ( .B(clk), .A(\g.we_clk [20147]));
Q_ASSIGN U12628 ( .B(clk), .A(\g.we_clk [20146]));
Q_ASSIGN U12629 ( .B(clk), .A(\g.we_clk [20145]));
Q_ASSIGN U12630 ( .B(clk), .A(\g.we_clk [20144]));
Q_ASSIGN U12631 ( .B(clk), .A(\g.we_clk [20143]));
Q_ASSIGN U12632 ( .B(clk), .A(\g.we_clk [20142]));
Q_ASSIGN U12633 ( .B(clk), .A(\g.we_clk [20141]));
Q_ASSIGN U12634 ( .B(clk), .A(\g.we_clk [20140]));
Q_ASSIGN U12635 ( .B(clk), .A(\g.we_clk [20139]));
Q_ASSIGN U12636 ( .B(clk), .A(\g.we_clk [20138]));
Q_ASSIGN U12637 ( .B(clk), .A(\g.we_clk [20137]));
Q_ASSIGN U12638 ( .B(clk), .A(\g.we_clk [20136]));
Q_ASSIGN U12639 ( .B(clk), .A(\g.we_clk [20135]));
Q_ASSIGN U12640 ( .B(clk), .A(\g.we_clk [20134]));
Q_ASSIGN U12641 ( .B(clk), .A(\g.we_clk [20133]));
Q_ASSIGN U12642 ( .B(clk), .A(\g.we_clk [20132]));
Q_ASSIGN U12643 ( .B(clk), .A(\g.we_clk [20131]));
Q_ASSIGN U12644 ( .B(clk), .A(\g.we_clk [20130]));
Q_ASSIGN U12645 ( .B(clk), .A(\g.we_clk [20129]));
Q_ASSIGN U12646 ( .B(clk), .A(\g.we_clk [20128]));
Q_ASSIGN U12647 ( .B(clk), .A(\g.we_clk [20127]));
Q_ASSIGN U12648 ( .B(clk), .A(\g.we_clk [20126]));
Q_ASSIGN U12649 ( .B(clk), .A(\g.we_clk [20125]));
Q_ASSIGN U12650 ( .B(clk), .A(\g.we_clk [20124]));
Q_ASSIGN U12651 ( .B(clk), .A(\g.we_clk [20123]));
Q_ASSIGN U12652 ( .B(clk), .A(\g.we_clk [20122]));
Q_ASSIGN U12653 ( .B(clk), .A(\g.we_clk [20121]));
Q_ASSIGN U12654 ( .B(clk), .A(\g.we_clk [20120]));
Q_ASSIGN U12655 ( .B(clk), .A(\g.we_clk [20119]));
Q_ASSIGN U12656 ( .B(clk), .A(\g.we_clk [20118]));
Q_ASSIGN U12657 ( .B(clk), .A(\g.we_clk [20117]));
Q_ASSIGN U12658 ( .B(clk), .A(\g.we_clk [20116]));
Q_ASSIGN U12659 ( .B(clk), .A(\g.we_clk [20115]));
Q_ASSIGN U12660 ( .B(clk), .A(\g.we_clk [20114]));
Q_ASSIGN U12661 ( .B(clk), .A(\g.we_clk [20113]));
Q_ASSIGN U12662 ( .B(clk), .A(\g.we_clk [20112]));
Q_ASSIGN U12663 ( .B(clk), .A(\g.we_clk [20111]));
Q_ASSIGN U12664 ( .B(clk), .A(\g.we_clk [20110]));
Q_ASSIGN U12665 ( .B(clk), .A(\g.we_clk [20109]));
Q_ASSIGN U12666 ( .B(clk), .A(\g.we_clk [20108]));
Q_ASSIGN U12667 ( .B(clk), .A(\g.we_clk [20107]));
Q_ASSIGN U12668 ( .B(clk), .A(\g.we_clk [20106]));
Q_ASSIGN U12669 ( .B(clk), .A(\g.we_clk [20105]));
Q_ASSIGN U12670 ( .B(clk), .A(\g.we_clk [20104]));
Q_ASSIGN U12671 ( .B(clk), .A(\g.we_clk [20103]));
Q_ASSIGN U12672 ( .B(clk), .A(\g.we_clk [20102]));
Q_ASSIGN U12673 ( .B(clk), .A(\g.we_clk [20101]));
Q_ASSIGN U12674 ( .B(clk), .A(\g.we_clk [20100]));
Q_ASSIGN U12675 ( .B(clk), .A(\g.we_clk [20099]));
Q_ASSIGN U12676 ( .B(clk), .A(\g.we_clk [20098]));
Q_ASSIGN U12677 ( .B(clk), .A(\g.we_clk [20097]));
Q_ASSIGN U12678 ( .B(clk), .A(\g.we_clk [20096]));
Q_ASSIGN U12679 ( .B(clk), .A(\g.we_clk [20095]));
Q_ASSIGN U12680 ( .B(clk), .A(\g.we_clk [20094]));
Q_ASSIGN U12681 ( .B(clk), .A(\g.we_clk [20093]));
Q_ASSIGN U12682 ( .B(clk), .A(\g.we_clk [20092]));
Q_ASSIGN U12683 ( .B(clk), .A(\g.we_clk [20091]));
Q_ASSIGN U12684 ( .B(clk), .A(\g.we_clk [20090]));
Q_ASSIGN U12685 ( .B(clk), .A(\g.we_clk [20089]));
Q_ASSIGN U12686 ( .B(clk), .A(\g.we_clk [20088]));
Q_ASSIGN U12687 ( .B(clk), .A(\g.we_clk [20087]));
Q_ASSIGN U12688 ( .B(clk), .A(\g.we_clk [20086]));
Q_ASSIGN U12689 ( .B(clk), .A(\g.we_clk [20085]));
Q_ASSIGN U12690 ( .B(clk), .A(\g.we_clk [20084]));
Q_ASSIGN U12691 ( .B(clk), .A(\g.we_clk [20083]));
Q_ASSIGN U12692 ( .B(clk), .A(\g.we_clk [20082]));
Q_ASSIGN U12693 ( .B(clk), .A(\g.we_clk [20081]));
Q_ASSIGN U12694 ( .B(clk), .A(\g.we_clk [20080]));
Q_ASSIGN U12695 ( .B(clk), .A(\g.we_clk [20079]));
Q_ASSIGN U12696 ( .B(clk), .A(\g.we_clk [20078]));
Q_ASSIGN U12697 ( .B(clk), .A(\g.we_clk [20077]));
Q_ASSIGN U12698 ( .B(clk), .A(\g.we_clk [20076]));
Q_ASSIGN U12699 ( .B(clk), .A(\g.we_clk [20075]));
Q_ASSIGN U12700 ( .B(clk), .A(\g.we_clk [20074]));
Q_ASSIGN U12701 ( .B(clk), .A(\g.we_clk [20073]));
Q_ASSIGN U12702 ( .B(clk), .A(\g.we_clk [20072]));
Q_ASSIGN U12703 ( .B(clk), .A(\g.we_clk [20071]));
Q_ASSIGN U12704 ( .B(clk), .A(\g.we_clk [20070]));
Q_ASSIGN U12705 ( .B(clk), .A(\g.we_clk [20069]));
Q_ASSIGN U12706 ( .B(clk), .A(\g.we_clk [20068]));
Q_ASSIGN U12707 ( .B(clk), .A(\g.we_clk [20067]));
Q_ASSIGN U12708 ( .B(clk), .A(\g.we_clk [20066]));
Q_ASSIGN U12709 ( .B(clk), .A(\g.we_clk [20065]));
Q_ASSIGN U12710 ( .B(clk), .A(\g.we_clk [20064]));
Q_ASSIGN U12711 ( .B(clk), .A(\g.we_clk [20063]));
Q_ASSIGN U12712 ( .B(clk), .A(\g.we_clk [20062]));
Q_ASSIGN U12713 ( .B(clk), .A(\g.we_clk [20061]));
Q_ASSIGN U12714 ( .B(clk), .A(\g.we_clk [20060]));
Q_ASSIGN U12715 ( .B(clk), .A(\g.we_clk [20059]));
Q_ASSIGN U12716 ( .B(clk), .A(\g.we_clk [20058]));
Q_ASSIGN U12717 ( .B(clk), .A(\g.we_clk [20057]));
Q_ASSIGN U12718 ( .B(clk), .A(\g.we_clk [20056]));
Q_ASSIGN U12719 ( .B(clk), .A(\g.we_clk [20055]));
Q_ASSIGN U12720 ( .B(clk), .A(\g.we_clk [20054]));
Q_ASSIGN U12721 ( .B(clk), .A(\g.we_clk [20053]));
Q_ASSIGN U12722 ( .B(clk), .A(\g.we_clk [20052]));
Q_ASSIGN U12723 ( .B(clk), .A(\g.we_clk [20051]));
Q_ASSIGN U12724 ( .B(clk), .A(\g.we_clk [20050]));
Q_ASSIGN U12725 ( .B(clk), .A(\g.we_clk [20049]));
Q_ASSIGN U12726 ( .B(clk), .A(\g.we_clk [20048]));
Q_ASSIGN U12727 ( .B(clk), .A(\g.we_clk [20047]));
Q_ASSIGN U12728 ( .B(clk), .A(\g.we_clk [20046]));
Q_ASSIGN U12729 ( .B(clk), .A(\g.we_clk [20045]));
Q_ASSIGN U12730 ( .B(clk), .A(\g.we_clk [20044]));
Q_ASSIGN U12731 ( .B(clk), .A(\g.we_clk [20043]));
Q_ASSIGN U12732 ( .B(clk), .A(\g.we_clk [20042]));
Q_ASSIGN U12733 ( .B(clk), .A(\g.we_clk [20041]));
Q_ASSIGN U12734 ( .B(clk), .A(\g.we_clk [20040]));
Q_ASSIGN U12735 ( .B(clk), .A(\g.we_clk [20039]));
Q_ASSIGN U12736 ( .B(clk), .A(\g.we_clk [20038]));
Q_ASSIGN U12737 ( .B(clk), .A(\g.we_clk [20037]));
Q_ASSIGN U12738 ( .B(clk), .A(\g.we_clk [20036]));
Q_ASSIGN U12739 ( .B(clk), .A(\g.we_clk [20035]));
Q_ASSIGN U12740 ( .B(clk), .A(\g.we_clk [20034]));
Q_ASSIGN U12741 ( .B(clk), .A(\g.we_clk [20033]));
Q_ASSIGN U12742 ( .B(clk), .A(\g.we_clk [20032]));
Q_ASSIGN U12743 ( .B(clk), .A(\g.we_clk [20031]));
Q_ASSIGN U12744 ( .B(clk), .A(\g.we_clk [20030]));
Q_ASSIGN U12745 ( .B(clk), .A(\g.we_clk [20029]));
Q_ASSIGN U12746 ( .B(clk), .A(\g.we_clk [20028]));
Q_ASSIGN U12747 ( .B(clk), .A(\g.we_clk [20027]));
Q_ASSIGN U12748 ( .B(clk), .A(\g.we_clk [20026]));
Q_ASSIGN U12749 ( .B(clk), .A(\g.we_clk [20025]));
Q_ASSIGN U12750 ( .B(clk), .A(\g.we_clk [20024]));
Q_ASSIGN U12751 ( .B(clk), .A(\g.we_clk [20023]));
Q_ASSIGN U12752 ( .B(clk), .A(\g.we_clk [20022]));
Q_ASSIGN U12753 ( .B(clk), .A(\g.we_clk [20021]));
Q_ASSIGN U12754 ( .B(clk), .A(\g.we_clk [20020]));
Q_ASSIGN U12755 ( .B(clk), .A(\g.we_clk [20019]));
Q_ASSIGN U12756 ( .B(clk), .A(\g.we_clk [20018]));
Q_ASSIGN U12757 ( .B(clk), .A(\g.we_clk [20017]));
Q_ASSIGN U12758 ( .B(clk), .A(\g.we_clk [20016]));
Q_ASSIGN U12759 ( .B(clk), .A(\g.we_clk [20015]));
Q_ASSIGN U12760 ( .B(clk), .A(\g.we_clk [20014]));
Q_ASSIGN U12761 ( .B(clk), .A(\g.we_clk [20013]));
Q_ASSIGN U12762 ( .B(clk), .A(\g.we_clk [20012]));
Q_ASSIGN U12763 ( .B(clk), .A(\g.we_clk [20011]));
Q_ASSIGN U12764 ( .B(clk), .A(\g.we_clk [20010]));
Q_ASSIGN U12765 ( .B(clk), .A(\g.we_clk [20009]));
Q_ASSIGN U12766 ( .B(clk), .A(\g.we_clk [20008]));
Q_ASSIGN U12767 ( .B(clk), .A(\g.we_clk [20007]));
Q_ASSIGN U12768 ( .B(clk), .A(\g.we_clk [20006]));
Q_ASSIGN U12769 ( .B(clk), .A(\g.we_clk [20005]));
Q_ASSIGN U12770 ( .B(clk), .A(\g.we_clk [20004]));
Q_ASSIGN U12771 ( .B(clk), .A(\g.we_clk [20003]));
Q_ASSIGN U12772 ( .B(clk), .A(\g.we_clk [20002]));
Q_ASSIGN U12773 ( .B(clk), .A(\g.we_clk [20001]));
Q_ASSIGN U12774 ( .B(clk), .A(\g.we_clk [20000]));
Q_ASSIGN U12775 ( .B(clk), .A(\g.we_clk [19999]));
Q_ASSIGN U12776 ( .B(clk), .A(\g.we_clk [19998]));
Q_ASSIGN U12777 ( .B(clk), .A(\g.we_clk [19997]));
Q_ASSIGN U12778 ( .B(clk), .A(\g.we_clk [19996]));
Q_ASSIGN U12779 ( .B(clk), .A(\g.we_clk [19995]));
Q_ASSIGN U12780 ( .B(clk), .A(\g.we_clk [19994]));
Q_ASSIGN U12781 ( .B(clk), .A(\g.we_clk [19993]));
Q_ASSIGN U12782 ( .B(clk), .A(\g.we_clk [19992]));
Q_ASSIGN U12783 ( .B(clk), .A(\g.we_clk [19991]));
Q_ASSIGN U12784 ( .B(clk), .A(\g.we_clk [19990]));
Q_ASSIGN U12785 ( .B(clk), .A(\g.we_clk [19989]));
Q_ASSIGN U12786 ( .B(clk), .A(\g.we_clk [19988]));
Q_ASSIGN U12787 ( .B(clk), .A(\g.we_clk [19987]));
Q_ASSIGN U12788 ( .B(clk), .A(\g.we_clk [19986]));
Q_ASSIGN U12789 ( .B(clk), .A(\g.we_clk [19985]));
Q_ASSIGN U12790 ( .B(clk), .A(\g.we_clk [19984]));
Q_ASSIGN U12791 ( .B(clk), .A(\g.we_clk [19983]));
Q_ASSIGN U12792 ( .B(clk), .A(\g.we_clk [19982]));
Q_ASSIGN U12793 ( .B(clk), .A(\g.we_clk [19981]));
Q_ASSIGN U12794 ( .B(clk), .A(\g.we_clk [19980]));
Q_ASSIGN U12795 ( .B(clk), .A(\g.we_clk [19979]));
Q_ASSIGN U12796 ( .B(clk), .A(\g.we_clk [19978]));
Q_ASSIGN U12797 ( .B(clk), .A(\g.we_clk [19977]));
Q_ASSIGN U12798 ( .B(clk), .A(\g.we_clk [19976]));
Q_ASSIGN U12799 ( .B(clk), .A(\g.we_clk [19975]));
Q_ASSIGN U12800 ( .B(clk), .A(\g.we_clk [19974]));
Q_ASSIGN U12801 ( .B(clk), .A(\g.we_clk [19973]));
Q_ASSIGN U12802 ( .B(clk), .A(\g.we_clk [19972]));
Q_ASSIGN U12803 ( .B(clk), .A(\g.we_clk [19971]));
Q_ASSIGN U12804 ( .B(clk), .A(\g.we_clk [19970]));
Q_ASSIGN U12805 ( .B(clk), .A(\g.we_clk [19969]));
Q_ASSIGN U12806 ( .B(clk), .A(\g.we_clk [19968]));
Q_ASSIGN U12807 ( .B(clk), .A(\g.we_clk [19967]));
Q_ASSIGN U12808 ( .B(clk), .A(\g.we_clk [19966]));
Q_ASSIGN U12809 ( .B(clk), .A(\g.we_clk [19965]));
Q_ASSIGN U12810 ( .B(clk), .A(\g.we_clk [19964]));
Q_ASSIGN U12811 ( .B(clk), .A(\g.we_clk [19963]));
Q_ASSIGN U12812 ( .B(clk), .A(\g.we_clk [19962]));
Q_ASSIGN U12813 ( .B(clk), .A(\g.we_clk [19961]));
Q_ASSIGN U12814 ( .B(clk), .A(\g.we_clk [19960]));
Q_ASSIGN U12815 ( .B(clk), .A(\g.we_clk [19959]));
Q_ASSIGN U12816 ( .B(clk), .A(\g.we_clk [19958]));
Q_ASSIGN U12817 ( .B(clk), .A(\g.we_clk [19957]));
Q_ASSIGN U12818 ( .B(clk), .A(\g.we_clk [19956]));
Q_ASSIGN U12819 ( .B(clk), .A(\g.we_clk [19955]));
Q_ASSIGN U12820 ( .B(clk), .A(\g.we_clk [19954]));
Q_ASSIGN U12821 ( .B(clk), .A(\g.we_clk [19953]));
Q_ASSIGN U12822 ( .B(clk), .A(\g.we_clk [19952]));
Q_ASSIGN U12823 ( .B(clk), .A(\g.we_clk [19951]));
Q_ASSIGN U12824 ( .B(clk), .A(\g.we_clk [19950]));
Q_ASSIGN U12825 ( .B(clk), .A(\g.we_clk [19949]));
Q_ASSIGN U12826 ( .B(clk), .A(\g.we_clk [19948]));
Q_ASSIGN U12827 ( .B(clk), .A(\g.we_clk [19947]));
Q_ASSIGN U12828 ( .B(clk), .A(\g.we_clk [19946]));
Q_ASSIGN U12829 ( .B(clk), .A(\g.we_clk [19945]));
Q_ASSIGN U12830 ( .B(clk), .A(\g.we_clk [19944]));
Q_ASSIGN U12831 ( .B(clk), .A(\g.we_clk [19943]));
Q_ASSIGN U12832 ( .B(clk), .A(\g.we_clk [19942]));
Q_ASSIGN U12833 ( .B(clk), .A(\g.we_clk [19941]));
Q_ASSIGN U12834 ( .B(clk), .A(\g.we_clk [19940]));
Q_ASSIGN U12835 ( .B(clk), .A(\g.we_clk [19939]));
Q_ASSIGN U12836 ( .B(clk), .A(\g.we_clk [19938]));
Q_ASSIGN U12837 ( .B(clk), .A(\g.we_clk [19937]));
Q_ASSIGN U12838 ( .B(clk), .A(\g.we_clk [19936]));
Q_ASSIGN U12839 ( .B(clk), .A(\g.we_clk [19935]));
Q_ASSIGN U12840 ( .B(clk), .A(\g.we_clk [19934]));
Q_ASSIGN U12841 ( .B(clk), .A(\g.we_clk [19933]));
Q_ASSIGN U12842 ( .B(clk), .A(\g.we_clk [19932]));
Q_ASSIGN U12843 ( .B(clk), .A(\g.we_clk [19931]));
Q_ASSIGN U12844 ( .B(clk), .A(\g.we_clk [19930]));
Q_ASSIGN U12845 ( .B(clk), .A(\g.we_clk [19929]));
Q_ASSIGN U12846 ( .B(clk), .A(\g.we_clk [19928]));
Q_ASSIGN U12847 ( .B(clk), .A(\g.we_clk [19927]));
Q_ASSIGN U12848 ( .B(clk), .A(\g.we_clk [19926]));
Q_ASSIGN U12849 ( .B(clk), .A(\g.we_clk [19925]));
Q_ASSIGN U12850 ( .B(clk), .A(\g.we_clk [19924]));
Q_ASSIGN U12851 ( .B(clk), .A(\g.we_clk [19923]));
Q_ASSIGN U12852 ( .B(clk), .A(\g.we_clk [19922]));
Q_ASSIGN U12853 ( .B(clk), .A(\g.we_clk [19921]));
Q_ASSIGN U12854 ( .B(clk), .A(\g.we_clk [19920]));
Q_ASSIGN U12855 ( .B(clk), .A(\g.we_clk [19919]));
Q_ASSIGN U12856 ( .B(clk), .A(\g.we_clk [19918]));
Q_ASSIGN U12857 ( .B(clk), .A(\g.we_clk [19917]));
Q_ASSIGN U12858 ( .B(clk), .A(\g.we_clk [19916]));
Q_ASSIGN U12859 ( .B(clk), .A(\g.we_clk [19915]));
Q_ASSIGN U12860 ( .B(clk), .A(\g.we_clk [19914]));
Q_ASSIGN U12861 ( .B(clk), .A(\g.we_clk [19913]));
Q_ASSIGN U12862 ( .B(clk), .A(\g.we_clk [19912]));
Q_ASSIGN U12863 ( .B(clk), .A(\g.we_clk [19911]));
Q_ASSIGN U12864 ( .B(clk), .A(\g.we_clk [19910]));
Q_ASSIGN U12865 ( .B(clk), .A(\g.we_clk [19909]));
Q_ASSIGN U12866 ( .B(clk), .A(\g.we_clk [19908]));
Q_ASSIGN U12867 ( .B(clk), .A(\g.we_clk [19907]));
Q_ASSIGN U12868 ( .B(clk), .A(\g.we_clk [19906]));
Q_ASSIGN U12869 ( .B(clk), .A(\g.we_clk [19905]));
Q_ASSIGN U12870 ( .B(clk), .A(\g.we_clk [19904]));
Q_ASSIGN U12871 ( .B(clk), .A(\g.we_clk [19903]));
Q_ASSIGN U12872 ( .B(clk), .A(\g.we_clk [19902]));
Q_ASSIGN U12873 ( .B(clk), .A(\g.we_clk [19901]));
Q_ASSIGN U12874 ( .B(clk), .A(\g.we_clk [19900]));
Q_ASSIGN U12875 ( .B(clk), .A(\g.we_clk [19899]));
Q_ASSIGN U12876 ( .B(clk), .A(\g.we_clk [19898]));
Q_ASSIGN U12877 ( .B(clk), .A(\g.we_clk [19897]));
Q_ASSIGN U12878 ( .B(clk), .A(\g.we_clk [19896]));
Q_ASSIGN U12879 ( .B(clk), .A(\g.we_clk [19895]));
Q_ASSIGN U12880 ( .B(clk), .A(\g.we_clk [19894]));
Q_ASSIGN U12881 ( .B(clk), .A(\g.we_clk [19893]));
Q_ASSIGN U12882 ( .B(clk), .A(\g.we_clk [19892]));
Q_ASSIGN U12883 ( .B(clk), .A(\g.we_clk [19891]));
Q_ASSIGN U12884 ( .B(clk), .A(\g.we_clk [19890]));
Q_ASSIGN U12885 ( .B(clk), .A(\g.we_clk [19889]));
Q_ASSIGN U12886 ( .B(clk), .A(\g.we_clk [19888]));
Q_ASSIGN U12887 ( .B(clk), .A(\g.we_clk [19887]));
Q_ASSIGN U12888 ( .B(clk), .A(\g.we_clk [19886]));
Q_ASSIGN U12889 ( .B(clk), .A(\g.we_clk [19885]));
Q_ASSIGN U12890 ( .B(clk), .A(\g.we_clk [19884]));
Q_ASSIGN U12891 ( .B(clk), .A(\g.we_clk [19883]));
Q_ASSIGN U12892 ( .B(clk), .A(\g.we_clk [19882]));
Q_ASSIGN U12893 ( .B(clk), .A(\g.we_clk [19881]));
Q_ASSIGN U12894 ( .B(clk), .A(\g.we_clk [19880]));
Q_ASSIGN U12895 ( .B(clk), .A(\g.we_clk [19879]));
Q_ASSIGN U12896 ( .B(clk), .A(\g.we_clk [19878]));
Q_ASSIGN U12897 ( .B(clk), .A(\g.we_clk [19877]));
Q_ASSIGN U12898 ( .B(clk), .A(\g.we_clk [19876]));
Q_ASSIGN U12899 ( .B(clk), .A(\g.we_clk [19875]));
Q_ASSIGN U12900 ( .B(clk), .A(\g.we_clk [19874]));
Q_ASSIGN U12901 ( .B(clk), .A(\g.we_clk [19873]));
Q_ASSIGN U12902 ( .B(clk), .A(\g.we_clk [19872]));
Q_ASSIGN U12903 ( .B(clk), .A(\g.we_clk [19871]));
Q_ASSIGN U12904 ( .B(clk), .A(\g.we_clk [19870]));
Q_ASSIGN U12905 ( .B(clk), .A(\g.we_clk [19869]));
Q_ASSIGN U12906 ( .B(clk), .A(\g.we_clk [19868]));
Q_ASSIGN U12907 ( .B(clk), .A(\g.we_clk [19867]));
Q_ASSIGN U12908 ( .B(clk), .A(\g.we_clk [19866]));
Q_ASSIGN U12909 ( .B(clk), .A(\g.we_clk [19865]));
Q_ASSIGN U12910 ( .B(clk), .A(\g.we_clk [19864]));
Q_ASSIGN U12911 ( .B(clk), .A(\g.we_clk [19863]));
Q_ASSIGN U12912 ( .B(clk), .A(\g.we_clk [19862]));
Q_ASSIGN U12913 ( .B(clk), .A(\g.we_clk [19861]));
Q_ASSIGN U12914 ( .B(clk), .A(\g.we_clk [19860]));
Q_ASSIGN U12915 ( .B(clk), .A(\g.we_clk [19859]));
Q_ASSIGN U12916 ( .B(clk), .A(\g.we_clk [19858]));
Q_ASSIGN U12917 ( .B(clk), .A(\g.we_clk [19857]));
Q_ASSIGN U12918 ( .B(clk), .A(\g.we_clk [19856]));
Q_ASSIGN U12919 ( .B(clk), .A(\g.we_clk [19855]));
Q_ASSIGN U12920 ( .B(clk), .A(\g.we_clk [19854]));
Q_ASSIGN U12921 ( .B(clk), .A(\g.we_clk [19853]));
Q_ASSIGN U12922 ( .B(clk), .A(\g.we_clk [19852]));
Q_ASSIGN U12923 ( .B(clk), .A(\g.we_clk [19851]));
Q_ASSIGN U12924 ( .B(clk), .A(\g.we_clk [19850]));
Q_ASSIGN U12925 ( .B(clk), .A(\g.we_clk [19849]));
Q_ASSIGN U12926 ( .B(clk), .A(\g.we_clk [19848]));
Q_ASSIGN U12927 ( .B(clk), .A(\g.we_clk [19847]));
Q_ASSIGN U12928 ( .B(clk), .A(\g.we_clk [19846]));
Q_ASSIGN U12929 ( .B(clk), .A(\g.we_clk [19845]));
Q_ASSIGN U12930 ( .B(clk), .A(\g.we_clk [19844]));
Q_ASSIGN U12931 ( .B(clk), .A(\g.we_clk [19843]));
Q_ASSIGN U12932 ( .B(clk), .A(\g.we_clk [19842]));
Q_ASSIGN U12933 ( .B(clk), .A(\g.we_clk [19841]));
Q_ASSIGN U12934 ( .B(clk), .A(\g.we_clk [19840]));
Q_ASSIGN U12935 ( .B(clk), .A(\g.we_clk [19839]));
Q_ASSIGN U12936 ( .B(clk), .A(\g.we_clk [19838]));
Q_ASSIGN U12937 ( .B(clk), .A(\g.we_clk [19837]));
Q_ASSIGN U12938 ( .B(clk), .A(\g.we_clk [19836]));
Q_ASSIGN U12939 ( .B(clk), .A(\g.we_clk [19835]));
Q_ASSIGN U12940 ( .B(clk), .A(\g.we_clk [19834]));
Q_ASSIGN U12941 ( .B(clk), .A(\g.we_clk [19833]));
Q_ASSIGN U12942 ( .B(clk), .A(\g.we_clk [19832]));
Q_ASSIGN U12943 ( .B(clk), .A(\g.we_clk [19831]));
Q_ASSIGN U12944 ( .B(clk), .A(\g.we_clk [19830]));
Q_ASSIGN U12945 ( .B(clk), .A(\g.we_clk [19829]));
Q_ASSIGN U12946 ( .B(clk), .A(\g.we_clk [19828]));
Q_ASSIGN U12947 ( .B(clk), .A(\g.we_clk [19827]));
Q_ASSIGN U12948 ( .B(clk), .A(\g.we_clk [19826]));
Q_ASSIGN U12949 ( .B(clk), .A(\g.we_clk [19825]));
Q_ASSIGN U12950 ( .B(clk), .A(\g.we_clk [19824]));
Q_ASSIGN U12951 ( .B(clk), .A(\g.we_clk [19823]));
Q_ASSIGN U12952 ( .B(clk), .A(\g.we_clk [19822]));
Q_ASSIGN U12953 ( .B(clk), .A(\g.we_clk [19821]));
Q_ASSIGN U12954 ( .B(clk), .A(\g.we_clk [19820]));
Q_ASSIGN U12955 ( .B(clk), .A(\g.we_clk [19819]));
Q_ASSIGN U12956 ( .B(clk), .A(\g.we_clk [19818]));
Q_ASSIGN U12957 ( .B(clk), .A(\g.we_clk [19817]));
Q_ASSIGN U12958 ( .B(clk), .A(\g.we_clk [19816]));
Q_ASSIGN U12959 ( .B(clk), .A(\g.we_clk [19815]));
Q_ASSIGN U12960 ( .B(clk), .A(\g.we_clk [19814]));
Q_ASSIGN U12961 ( .B(clk), .A(\g.we_clk [19813]));
Q_ASSIGN U12962 ( .B(clk), .A(\g.we_clk [19812]));
Q_ASSIGN U12963 ( .B(clk), .A(\g.we_clk [19811]));
Q_ASSIGN U12964 ( .B(clk), .A(\g.we_clk [19810]));
Q_ASSIGN U12965 ( .B(clk), .A(\g.we_clk [19809]));
Q_ASSIGN U12966 ( .B(clk), .A(\g.we_clk [19808]));
Q_ASSIGN U12967 ( .B(clk), .A(\g.we_clk [19807]));
Q_ASSIGN U12968 ( .B(clk), .A(\g.we_clk [19806]));
Q_ASSIGN U12969 ( .B(clk), .A(\g.we_clk [19805]));
Q_ASSIGN U12970 ( .B(clk), .A(\g.we_clk [19804]));
Q_ASSIGN U12971 ( .B(clk), .A(\g.we_clk [19803]));
Q_ASSIGN U12972 ( .B(clk), .A(\g.we_clk [19802]));
Q_ASSIGN U12973 ( .B(clk), .A(\g.we_clk [19801]));
Q_ASSIGN U12974 ( .B(clk), .A(\g.we_clk [19800]));
Q_ASSIGN U12975 ( .B(clk), .A(\g.we_clk [19799]));
Q_ASSIGN U12976 ( .B(clk), .A(\g.we_clk [19798]));
Q_ASSIGN U12977 ( .B(clk), .A(\g.we_clk [19797]));
Q_ASSIGN U12978 ( .B(clk), .A(\g.we_clk [19796]));
Q_ASSIGN U12979 ( .B(clk), .A(\g.we_clk [19795]));
Q_ASSIGN U12980 ( .B(clk), .A(\g.we_clk [19794]));
Q_ASSIGN U12981 ( .B(clk), .A(\g.we_clk [19793]));
Q_ASSIGN U12982 ( .B(clk), .A(\g.we_clk [19792]));
Q_ASSIGN U12983 ( .B(clk), .A(\g.we_clk [19791]));
Q_ASSIGN U12984 ( .B(clk), .A(\g.we_clk [19790]));
Q_ASSIGN U12985 ( .B(clk), .A(\g.we_clk [19789]));
Q_ASSIGN U12986 ( .B(clk), .A(\g.we_clk [19788]));
Q_ASSIGN U12987 ( .B(clk), .A(\g.we_clk [19787]));
Q_ASSIGN U12988 ( .B(clk), .A(\g.we_clk [19786]));
Q_ASSIGN U12989 ( .B(clk), .A(\g.we_clk [19785]));
Q_ASSIGN U12990 ( .B(clk), .A(\g.we_clk [19784]));
Q_ASSIGN U12991 ( .B(clk), .A(\g.we_clk [19783]));
Q_ASSIGN U12992 ( .B(clk), .A(\g.we_clk [19782]));
Q_ASSIGN U12993 ( .B(clk), .A(\g.we_clk [19781]));
Q_ASSIGN U12994 ( .B(clk), .A(\g.we_clk [19780]));
Q_ASSIGN U12995 ( .B(clk), .A(\g.we_clk [19779]));
Q_ASSIGN U12996 ( .B(clk), .A(\g.we_clk [19778]));
Q_ASSIGN U12997 ( .B(clk), .A(\g.we_clk [19777]));
Q_ASSIGN U12998 ( .B(clk), .A(\g.we_clk [19776]));
Q_ASSIGN U12999 ( .B(clk), .A(\g.we_clk [19775]));
Q_ASSIGN U13000 ( .B(clk), .A(\g.we_clk [19774]));
Q_ASSIGN U13001 ( .B(clk), .A(\g.we_clk [19773]));
Q_ASSIGN U13002 ( .B(clk), .A(\g.we_clk [19772]));
Q_ASSIGN U13003 ( .B(clk), .A(\g.we_clk [19771]));
Q_ASSIGN U13004 ( .B(clk), .A(\g.we_clk [19770]));
Q_ASSIGN U13005 ( .B(clk), .A(\g.we_clk [19769]));
Q_ASSIGN U13006 ( .B(clk), .A(\g.we_clk [19768]));
Q_ASSIGN U13007 ( .B(clk), .A(\g.we_clk [19767]));
Q_ASSIGN U13008 ( .B(clk), .A(\g.we_clk [19766]));
Q_ASSIGN U13009 ( .B(clk), .A(\g.we_clk [19765]));
Q_ASSIGN U13010 ( .B(clk), .A(\g.we_clk [19764]));
Q_ASSIGN U13011 ( .B(clk), .A(\g.we_clk [19763]));
Q_ASSIGN U13012 ( .B(clk), .A(\g.we_clk [19762]));
Q_ASSIGN U13013 ( .B(clk), .A(\g.we_clk [19761]));
Q_ASSIGN U13014 ( .B(clk), .A(\g.we_clk [19760]));
Q_ASSIGN U13015 ( .B(clk), .A(\g.we_clk [19759]));
Q_ASSIGN U13016 ( .B(clk), .A(\g.we_clk [19758]));
Q_ASSIGN U13017 ( .B(clk), .A(\g.we_clk [19757]));
Q_ASSIGN U13018 ( .B(clk), .A(\g.we_clk [19756]));
Q_ASSIGN U13019 ( .B(clk), .A(\g.we_clk [19755]));
Q_ASSIGN U13020 ( .B(clk), .A(\g.we_clk [19754]));
Q_ASSIGN U13021 ( .B(clk), .A(\g.we_clk [19753]));
Q_ASSIGN U13022 ( .B(clk), .A(\g.we_clk [19752]));
Q_ASSIGN U13023 ( .B(clk), .A(\g.we_clk [19751]));
Q_ASSIGN U13024 ( .B(clk), .A(\g.we_clk [19750]));
Q_ASSIGN U13025 ( .B(clk), .A(\g.we_clk [19749]));
Q_ASSIGN U13026 ( .B(clk), .A(\g.we_clk [19748]));
Q_ASSIGN U13027 ( .B(clk), .A(\g.we_clk [19747]));
Q_ASSIGN U13028 ( .B(clk), .A(\g.we_clk [19746]));
Q_ASSIGN U13029 ( .B(clk), .A(\g.we_clk [19745]));
Q_ASSIGN U13030 ( .B(clk), .A(\g.we_clk [19744]));
Q_ASSIGN U13031 ( .B(clk), .A(\g.we_clk [19743]));
Q_ASSIGN U13032 ( .B(clk), .A(\g.we_clk [19742]));
Q_ASSIGN U13033 ( .B(clk), .A(\g.we_clk [19741]));
Q_ASSIGN U13034 ( .B(clk), .A(\g.we_clk [19740]));
Q_ASSIGN U13035 ( .B(clk), .A(\g.we_clk [19739]));
Q_ASSIGN U13036 ( .B(clk), .A(\g.we_clk [19738]));
Q_ASSIGN U13037 ( .B(clk), .A(\g.we_clk [19737]));
Q_ASSIGN U13038 ( .B(clk), .A(\g.we_clk [19736]));
Q_ASSIGN U13039 ( .B(clk), .A(\g.we_clk [19735]));
Q_ASSIGN U13040 ( .B(clk), .A(\g.we_clk [19734]));
Q_ASSIGN U13041 ( .B(clk), .A(\g.we_clk [19733]));
Q_ASSIGN U13042 ( .B(clk), .A(\g.we_clk [19732]));
Q_ASSIGN U13043 ( .B(clk), .A(\g.we_clk [19731]));
Q_ASSIGN U13044 ( .B(clk), .A(\g.we_clk [19730]));
Q_ASSIGN U13045 ( .B(clk), .A(\g.we_clk [19729]));
Q_ASSIGN U13046 ( .B(clk), .A(\g.we_clk [19728]));
Q_ASSIGN U13047 ( .B(clk), .A(\g.we_clk [19727]));
Q_ASSIGN U13048 ( .B(clk), .A(\g.we_clk [19726]));
Q_ASSIGN U13049 ( .B(clk), .A(\g.we_clk [19725]));
Q_ASSIGN U13050 ( .B(clk), .A(\g.we_clk [19724]));
Q_ASSIGN U13051 ( .B(clk), .A(\g.we_clk [19723]));
Q_ASSIGN U13052 ( .B(clk), .A(\g.we_clk [19722]));
Q_ASSIGN U13053 ( .B(clk), .A(\g.we_clk [19721]));
Q_ASSIGN U13054 ( .B(clk), .A(\g.we_clk [19720]));
Q_ASSIGN U13055 ( .B(clk), .A(\g.we_clk [19719]));
Q_ASSIGN U13056 ( .B(clk), .A(\g.we_clk [19718]));
Q_ASSIGN U13057 ( .B(clk), .A(\g.we_clk [19717]));
Q_ASSIGN U13058 ( .B(clk), .A(\g.we_clk [19716]));
Q_ASSIGN U13059 ( .B(clk), .A(\g.we_clk [19715]));
Q_ASSIGN U13060 ( .B(clk), .A(\g.we_clk [19714]));
Q_ASSIGN U13061 ( .B(clk), .A(\g.we_clk [19713]));
Q_ASSIGN U13062 ( .B(clk), .A(\g.we_clk [19712]));
Q_ASSIGN U13063 ( .B(clk), .A(\g.we_clk [19711]));
Q_ASSIGN U13064 ( .B(clk), .A(\g.we_clk [19710]));
Q_ASSIGN U13065 ( .B(clk), .A(\g.we_clk [19709]));
Q_ASSIGN U13066 ( .B(clk), .A(\g.we_clk [19708]));
Q_ASSIGN U13067 ( .B(clk), .A(\g.we_clk [19707]));
Q_ASSIGN U13068 ( .B(clk), .A(\g.we_clk [19706]));
Q_ASSIGN U13069 ( .B(clk), .A(\g.we_clk [19705]));
Q_ASSIGN U13070 ( .B(clk), .A(\g.we_clk [19704]));
Q_ASSIGN U13071 ( .B(clk), .A(\g.we_clk [19703]));
Q_ASSIGN U13072 ( .B(clk), .A(\g.we_clk [19702]));
Q_ASSIGN U13073 ( .B(clk), .A(\g.we_clk [19701]));
Q_ASSIGN U13074 ( .B(clk), .A(\g.we_clk [19700]));
Q_ASSIGN U13075 ( .B(clk), .A(\g.we_clk [19699]));
Q_ASSIGN U13076 ( .B(clk), .A(\g.we_clk [19698]));
Q_ASSIGN U13077 ( .B(clk), .A(\g.we_clk [19697]));
Q_ASSIGN U13078 ( .B(clk), .A(\g.we_clk [19696]));
Q_ASSIGN U13079 ( .B(clk), .A(\g.we_clk [19695]));
Q_ASSIGN U13080 ( .B(clk), .A(\g.we_clk [19694]));
Q_ASSIGN U13081 ( .B(clk), .A(\g.we_clk [19693]));
Q_ASSIGN U13082 ( .B(clk), .A(\g.we_clk [19692]));
Q_ASSIGN U13083 ( .B(clk), .A(\g.we_clk [19691]));
Q_ASSIGN U13084 ( .B(clk), .A(\g.we_clk [19690]));
Q_ASSIGN U13085 ( .B(clk), .A(\g.we_clk [19689]));
Q_ASSIGN U13086 ( .B(clk), .A(\g.we_clk [19688]));
Q_ASSIGN U13087 ( .B(clk), .A(\g.we_clk [19687]));
Q_ASSIGN U13088 ( .B(clk), .A(\g.we_clk [19686]));
Q_ASSIGN U13089 ( .B(clk), .A(\g.we_clk [19685]));
Q_ASSIGN U13090 ( .B(clk), .A(\g.we_clk [19684]));
Q_ASSIGN U13091 ( .B(clk), .A(\g.we_clk [19683]));
Q_ASSIGN U13092 ( .B(clk), .A(\g.we_clk [19682]));
Q_ASSIGN U13093 ( .B(clk), .A(\g.we_clk [19681]));
Q_ASSIGN U13094 ( .B(clk), .A(\g.we_clk [19680]));
Q_ASSIGN U13095 ( .B(clk), .A(\g.we_clk [19679]));
Q_ASSIGN U13096 ( .B(clk), .A(\g.we_clk [19678]));
Q_ASSIGN U13097 ( .B(clk), .A(\g.we_clk [19677]));
Q_ASSIGN U13098 ( .B(clk), .A(\g.we_clk [19676]));
Q_ASSIGN U13099 ( .B(clk), .A(\g.we_clk [19675]));
Q_ASSIGN U13100 ( .B(clk), .A(\g.we_clk [19674]));
Q_ASSIGN U13101 ( .B(clk), .A(\g.we_clk [19673]));
Q_ASSIGN U13102 ( .B(clk), .A(\g.we_clk [19672]));
Q_ASSIGN U13103 ( .B(clk), .A(\g.we_clk [19671]));
Q_ASSIGN U13104 ( .B(clk), .A(\g.we_clk [19670]));
Q_ASSIGN U13105 ( .B(clk), .A(\g.we_clk [19669]));
Q_ASSIGN U13106 ( .B(clk), .A(\g.we_clk [19668]));
Q_ASSIGN U13107 ( .B(clk), .A(\g.we_clk [19667]));
Q_ASSIGN U13108 ( .B(clk), .A(\g.we_clk [19666]));
Q_ASSIGN U13109 ( .B(clk), .A(\g.we_clk [19665]));
Q_ASSIGN U13110 ( .B(clk), .A(\g.we_clk [19664]));
Q_ASSIGN U13111 ( .B(clk), .A(\g.we_clk [19663]));
Q_ASSIGN U13112 ( .B(clk), .A(\g.we_clk [19662]));
Q_ASSIGN U13113 ( .B(clk), .A(\g.we_clk [19661]));
Q_ASSIGN U13114 ( .B(clk), .A(\g.we_clk [19660]));
Q_ASSIGN U13115 ( .B(clk), .A(\g.we_clk [19659]));
Q_ASSIGN U13116 ( .B(clk), .A(\g.we_clk [19658]));
Q_ASSIGN U13117 ( .B(clk), .A(\g.we_clk [19657]));
Q_ASSIGN U13118 ( .B(clk), .A(\g.we_clk [19656]));
Q_ASSIGN U13119 ( .B(clk), .A(\g.we_clk [19655]));
Q_ASSIGN U13120 ( .B(clk), .A(\g.we_clk [19654]));
Q_ASSIGN U13121 ( .B(clk), .A(\g.we_clk [19653]));
Q_ASSIGN U13122 ( .B(clk), .A(\g.we_clk [19652]));
Q_ASSIGN U13123 ( .B(clk), .A(\g.we_clk [19651]));
Q_ASSIGN U13124 ( .B(clk), .A(\g.we_clk [19650]));
Q_ASSIGN U13125 ( .B(clk), .A(\g.we_clk [19649]));
Q_ASSIGN U13126 ( .B(clk), .A(\g.we_clk [19648]));
Q_ASSIGN U13127 ( .B(clk), .A(\g.we_clk [19647]));
Q_ASSIGN U13128 ( .B(clk), .A(\g.we_clk [19646]));
Q_ASSIGN U13129 ( .B(clk), .A(\g.we_clk [19645]));
Q_ASSIGN U13130 ( .B(clk), .A(\g.we_clk [19644]));
Q_ASSIGN U13131 ( .B(clk), .A(\g.we_clk [19643]));
Q_ASSIGN U13132 ( .B(clk), .A(\g.we_clk [19642]));
Q_ASSIGN U13133 ( .B(clk), .A(\g.we_clk [19641]));
Q_ASSIGN U13134 ( .B(clk), .A(\g.we_clk [19640]));
Q_ASSIGN U13135 ( .B(clk), .A(\g.we_clk [19639]));
Q_ASSIGN U13136 ( .B(clk), .A(\g.we_clk [19638]));
Q_ASSIGN U13137 ( .B(clk), .A(\g.we_clk [19637]));
Q_ASSIGN U13138 ( .B(clk), .A(\g.we_clk [19636]));
Q_ASSIGN U13139 ( .B(clk), .A(\g.we_clk [19635]));
Q_ASSIGN U13140 ( .B(clk), .A(\g.we_clk [19634]));
Q_ASSIGN U13141 ( .B(clk), .A(\g.we_clk [19633]));
Q_ASSIGN U13142 ( .B(clk), .A(\g.we_clk [19632]));
Q_ASSIGN U13143 ( .B(clk), .A(\g.we_clk [19631]));
Q_ASSIGN U13144 ( .B(clk), .A(\g.we_clk [19630]));
Q_ASSIGN U13145 ( .B(clk), .A(\g.we_clk [19629]));
Q_ASSIGN U13146 ( .B(clk), .A(\g.we_clk [19628]));
Q_ASSIGN U13147 ( .B(clk), .A(\g.we_clk [19627]));
Q_ASSIGN U13148 ( .B(clk), .A(\g.we_clk [19626]));
Q_ASSIGN U13149 ( .B(clk), .A(\g.we_clk [19625]));
Q_ASSIGN U13150 ( .B(clk), .A(\g.we_clk [19624]));
Q_ASSIGN U13151 ( .B(clk), .A(\g.we_clk [19623]));
Q_ASSIGN U13152 ( .B(clk), .A(\g.we_clk [19622]));
Q_ASSIGN U13153 ( .B(clk), .A(\g.we_clk [19621]));
Q_ASSIGN U13154 ( .B(clk), .A(\g.we_clk [19620]));
Q_ASSIGN U13155 ( .B(clk), .A(\g.we_clk [19619]));
Q_ASSIGN U13156 ( .B(clk), .A(\g.we_clk [19618]));
Q_ASSIGN U13157 ( .B(clk), .A(\g.we_clk [19617]));
Q_ASSIGN U13158 ( .B(clk), .A(\g.we_clk [19616]));
Q_ASSIGN U13159 ( .B(clk), .A(\g.we_clk [19615]));
Q_ASSIGN U13160 ( .B(clk), .A(\g.we_clk [19614]));
Q_ASSIGN U13161 ( .B(clk), .A(\g.we_clk [19613]));
Q_ASSIGN U13162 ( .B(clk), .A(\g.we_clk [19612]));
Q_ASSIGN U13163 ( .B(clk), .A(\g.we_clk [19611]));
Q_ASSIGN U13164 ( .B(clk), .A(\g.we_clk [19610]));
Q_ASSIGN U13165 ( .B(clk), .A(\g.we_clk [19609]));
Q_ASSIGN U13166 ( .B(clk), .A(\g.we_clk [19608]));
Q_ASSIGN U13167 ( .B(clk), .A(\g.we_clk [19607]));
Q_ASSIGN U13168 ( .B(clk), .A(\g.we_clk [19606]));
Q_ASSIGN U13169 ( .B(clk), .A(\g.we_clk [19605]));
Q_ASSIGN U13170 ( .B(clk), .A(\g.we_clk [19604]));
Q_ASSIGN U13171 ( .B(clk), .A(\g.we_clk [19603]));
Q_ASSIGN U13172 ( .B(clk), .A(\g.we_clk [19602]));
Q_ASSIGN U13173 ( .B(clk), .A(\g.we_clk [19601]));
Q_ASSIGN U13174 ( .B(clk), .A(\g.we_clk [19600]));
Q_ASSIGN U13175 ( .B(clk), .A(\g.we_clk [19599]));
Q_ASSIGN U13176 ( .B(clk), .A(\g.we_clk [19598]));
Q_ASSIGN U13177 ( .B(clk), .A(\g.we_clk [19597]));
Q_ASSIGN U13178 ( .B(clk), .A(\g.we_clk [19596]));
Q_ASSIGN U13179 ( .B(clk), .A(\g.we_clk [19595]));
Q_ASSIGN U13180 ( .B(clk), .A(\g.we_clk [19594]));
Q_ASSIGN U13181 ( .B(clk), .A(\g.we_clk [19593]));
Q_ASSIGN U13182 ( .B(clk), .A(\g.we_clk [19592]));
Q_ASSIGN U13183 ( .B(clk), .A(\g.we_clk [19591]));
Q_ASSIGN U13184 ( .B(clk), .A(\g.we_clk [19590]));
Q_ASSIGN U13185 ( .B(clk), .A(\g.we_clk [19589]));
Q_ASSIGN U13186 ( .B(clk), .A(\g.we_clk [19588]));
Q_ASSIGN U13187 ( .B(clk), .A(\g.we_clk [19587]));
Q_ASSIGN U13188 ( .B(clk), .A(\g.we_clk [19586]));
Q_ASSIGN U13189 ( .B(clk), .A(\g.we_clk [19585]));
Q_ASSIGN U13190 ( .B(clk), .A(\g.we_clk [19584]));
Q_ASSIGN U13191 ( .B(clk), .A(\g.we_clk [19583]));
Q_ASSIGN U13192 ( .B(clk), .A(\g.we_clk [19582]));
Q_ASSIGN U13193 ( .B(clk), .A(\g.we_clk [19581]));
Q_ASSIGN U13194 ( .B(clk), .A(\g.we_clk [19580]));
Q_ASSIGN U13195 ( .B(clk), .A(\g.we_clk [19579]));
Q_ASSIGN U13196 ( .B(clk), .A(\g.we_clk [19578]));
Q_ASSIGN U13197 ( .B(clk), .A(\g.we_clk [19577]));
Q_ASSIGN U13198 ( .B(clk), .A(\g.we_clk [19576]));
Q_ASSIGN U13199 ( .B(clk), .A(\g.we_clk [19575]));
Q_ASSIGN U13200 ( .B(clk), .A(\g.we_clk [19574]));
Q_ASSIGN U13201 ( .B(clk), .A(\g.we_clk [19573]));
Q_ASSIGN U13202 ( .B(clk), .A(\g.we_clk [19572]));
Q_ASSIGN U13203 ( .B(clk), .A(\g.we_clk [19571]));
Q_ASSIGN U13204 ( .B(clk), .A(\g.we_clk [19570]));
Q_ASSIGN U13205 ( .B(clk), .A(\g.we_clk [19569]));
Q_ASSIGN U13206 ( .B(clk), .A(\g.we_clk [19568]));
Q_ASSIGN U13207 ( .B(clk), .A(\g.we_clk [19567]));
Q_ASSIGN U13208 ( .B(clk), .A(\g.we_clk [19566]));
Q_ASSIGN U13209 ( .B(clk), .A(\g.we_clk [19565]));
Q_ASSIGN U13210 ( .B(clk), .A(\g.we_clk [19564]));
Q_ASSIGN U13211 ( .B(clk), .A(\g.we_clk [19563]));
Q_ASSIGN U13212 ( .B(clk), .A(\g.we_clk [19562]));
Q_ASSIGN U13213 ( .B(clk), .A(\g.we_clk [19561]));
Q_ASSIGN U13214 ( .B(clk), .A(\g.we_clk [19560]));
Q_ASSIGN U13215 ( .B(clk), .A(\g.we_clk [19559]));
Q_ASSIGN U13216 ( .B(clk), .A(\g.we_clk [19558]));
Q_ASSIGN U13217 ( .B(clk), .A(\g.we_clk [19557]));
Q_ASSIGN U13218 ( .B(clk), .A(\g.we_clk [19556]));
Q_ASSIGN U13219 ( .B(clk), .A(\g.we_clk [19555]));
Q_ASSIGN U13220 ( .B(clk), .A(\g.we_clk [19554]));
Q_ASSIGN U13221 ( .B(clk), .A(\g.we_clk [19553]));
Q_ASSIGN U13222 ( .B(clk), .A(\g.we_clk [19552]));
Q_ASSIGN U13223 ( .B(clk), .A(\g.we_clk [19551]));
Q_ASSIGN U13224 ( .B(clk), .A(\g.we_clk [19550]));
Q_ASSIGN U13225 ( .B(clk), .A(\g.we_clk [19549]));
Q_ASSIGN U13226 ( .B(clk), .A(\g.we_clk [19548]));
Q_ASSIGN U13227 ( .B(clk), .A(\g.we_clk [19547]));
Q_ASSIGN U13228 ( .B(clk), .A(\g.we_clk [19546]));
Q_ASSIGN U13229 ( .B(clk), .A(\g.we_clk [19545]));
Q_ASSIGN U13230 ( .B(clk), .A(\g.we_clk [19544]));
Q_ASSIGN U13231 ( .B(clk), .A(\g.we_clk [19543]));
Q_ASSIGN U13232 ( .B(clk), .A(\g.we_clk [19542]));
Q_ASSIGN U13233 ( .B(clk), .A(\g.we_clk [19541]));
Q_ASSIGN U13234 ( .B(clk), .A(\g.we_clk [19540]));
Q_ASSIGN U13235 ( .B(clk), .A(\g.we_clk [19539]));
Q_ASSIGN U13236 ( .B(clk), .A(\g.we_clk [19538]));
Q_ASSIGN U13237 ( .B(clk), .A(\g.we_clk [19537]));
Q_ASSIGN U13238 ( .B(clk), .A(\g.we_clk [19536]));
Q_ASSIGN U13239 ( .B(clk), .A(\g.we_clk [19535]));
Q_ASSIGN U13240 ( .B(clk), .A(\g.we_clk [19534]));
Q_ASSIGN U13241 ( .B(clk), .A(\g.we_clk [19533]));
Q_ASSIGN U13242 ( .B(clk), .A(\g.we_clk [19532]));
Q_ASSIGN U13243 ( .B(clk), .A(\g.we_clk [19531]));
Q_ASSIGN U13244 ( .B(clk), .A(\g.we_clk [19530]));
Q_ASSIGN U13245 ( .B(clk), .A(\g.we_clk [19529]));
Q_ASSIGN U13246 ( .B(clk), .A(\g.we_clk [19528]));
Q_ASSIGN U13247 ( .B(clk), .A(\g.we_clk [19527]));
Q_ASSIGN U13248 ( .B(clk), .A(\g.we_clk [19526]));
Q_ASSIGN U13249 ( .B(clk), .A(\g.we_clk [19525]));
Q_ASSIGN U13250 ( .B(clk), .A(\g.we_clk [19524]));
Q_ASSIGN U13251 ( .B(clk), .A(\g.we_clk [19523]));
Q_ASSIGN U13252 ( .B(clk), .A(\g.we_clk [19522]));
Q_ASSIGN U13253 ( .B(clk), .A(\g.we_clk [19521]));
Q_ASSIGN U13254 ( .B(clk), .A(\g.we_clk [19520]));
Q_ASSIGN U13255 ( .B(clk), .A(\g.we_clk [19519]));
Q_ASSIGN U13256 ( .B(clk), .A(\g.we_clk [19518]));
Q_ASSIGN U13257 ( .B(clk), .A(\g.we_clk [19517]));
Q_ASSIGN U13258 ( .B(clk), .A(\g.we_clk [19516]));
Q_ASSIGN U13259 ( .B(clk), .A(\g.we_clk [19515]));
Q_ASSIGN U13260 ( .B(clk), .A(\g.we_clk [19514]));
Q_ASSIGN U13261 ( .B(clk), .A(\g.we_clk [19513]));
Q_ASSIGN U13262 ( .B(clk), .A(\g.we_clk [19512]));
Q_ASSIGN U13263 ( .B(clk), .A(\g.we_clk [19511]));
Q_ASSIGN U13264 ( .B(clk), .A(\g.we_clk [19510]));
Q_ASSIGN U13265 ( .B(clk), .A(\g.we_clk [19509]));
Q_ASSIGN U13266 ( .B(clk), .A(\g.we_clk [19508]));
Q_ASSIGN U13267 ( .B(clk), .A(\g.we_clk [19507]));
Q_ASSIGN U13268 ( .B(clk), .A(\g.we_clk [19506]));
Q_ASSIGN U13269 ( .B(clk), .A(\g.we_clk [19505]));
Q_ASSIGN U13270 ( .B(clk), .A(\g.we_clk [19504]));
Q_ASSIGN U13271 ( .B(clk), .A(\g.we_clk [19503]));
Q_ASSIGN U13272 ( .B(clk), .A(\g.we_clk [19502]));
Q_ASSIGN U13273 ( .B(clk), .A(\g.we_clk [19501]));
Q_ASSIGN U13274 ( .B(clk), .A(\g.we_clk [19500]));
Q_ASSIGN U13275 ( .B(clk), .A(\g.we_clk [19499]));
Q_ASSIGN U13276 ( .B(clk), .A(\g.we_clk [19498]));
Q_ASSIGN U13277 ( .B(clk), .A(\g.we_clk [19497]));
Q_ASSIGN U13278 ( .B(clk), .A(\g.we_clk [19496]));
Q_ASSIGN U13279 ( .B(clk), .A(\g.we_clk [19495]));
Q_ASSIGN U13280 ( .B(clk), .A(\g.we_clk [19494]));
Q_ASSIGN U13281 ( .B(clk), .A(\g.we_clk [19493]));
Q_ASSIGN U13282 ( .B(clk), .A(\g.we_clk [19492]));
Q_ASSIGN U13283 ( .B(clk), .A(\g.we_clk [19491]));
Q_ASSIGN U13284 ( .B(clk), .A(\g.we_clk [19490]));
Q_ASSIGN U13285 ( .B(clk), .A(\g.we_clk [19489]));
Q_ASSIGN U13286 ( .B(clk), .A(\g.we_clk [19488]));
Q_ASSIGN U13287 ( .B(clk), .A(\g.we_clk [19487]));
Q_ASSIGN U13288 ( .B(clk), .A(\g.we_clk [19486]));
Q_ASSIGN U13289 ( .B(clk), .A(\g.we_clk [19485]));
Q_ASSIGN U13290 ( .B(clk), .A(\g.we_clk [19484]));
Q_ASSIGN U13291 ( .B(clk), .A(\g.we_clk [19483]));
Q_ASSIGN U13292 ( .B(clk), .A(\g.we_clk [19482]));
Q_ASSIGN U13293 ( .B(clk), .A(\g.we_clk [19481]));
Q_ASSIGN U13294 ( .B(clk), .A(\g.we_clk [19480]));
Q_ASSIGN U13295 ( .B(clk), .A(\g.we_clk [19479]));
Q_ASSIGN U13296 ( .B(clk), .A(\g.we_clk [19478]));
Q_ASSIGN U13297 ( .B(clk), .A(\g.we_clk [19477]));
Q_ASSIGN U13298 ( .B(clk), .A(\g.we_clk [19476]));
Q_ASSIGN U13299 ( .B(clk), .A(\g.we_clk [19475]));
Q_ASSIGN U13300 ( .B(clk), .A(\g.we_clk [19474]));
Q_ASSIGN U13301 ( .B(clk), .A(\g.we_clk [19473]));
Q_ASSIGN U13302 ( .B(clk), .A(\g.we_clk [19472]));
Q_ASSIGN U13303 ( .B(clk), .A(\g.we_clk [19471]));
Q_ASSIGN U13304 ( .B(clk), .A(\g.we_clk [19470]));
Q_ASSIGN U13305 ( .B(clk), .A(\g.we_clk [19469]));
Q_ASSIGN U13306 ( .B(clk), .A(\g.we_clk [19468]));
Q_ASSIGN U13307 ( .B(clk), .A(\g.we_clk [19467]));
Q_ASSIGN U13308 ( .B(clk), .A(\g.we_clk [19466]));
Q_ASSIGN U13309 ( .B(clk), .A(\g.we_clk [19465]));
Q_ASSIGN U13310 ( .B(clk), .A(\g.we_clk [19464]));
Q_ASSIGN U13311 ( .B(clk), .A(\g.we_clk [19463]));
Q_ASSIGN U13312 ( .B(clk), .A(\g.we_clk [19462]));
Q_ASSIGN U13313 ( .B(clk), .A(\g.we_clk [19461]));
Q_ASSIGN U13314 ( .B(clk), .A(\g.we_clk [19460]));
Q_ASSIGN U13315 ( .B(clk), .A(\g.we_clk [19459]));
Q_ASSIGN U13316 ( .B(clk), .A(\g.we_clk [19458]));
Q_ASSIGN U13317 ( .B(clk), .A(\g.we_clk [19457]));
Q_ASSIGN U13318 ( .B(clk), .A(\g.we_clk [19456]));
Q_ASSIGN U13319 ( .B(clk), .A(\g.we_clk [19455]));
Q_ASSIGN U13320 ( .B(clk), .A(\g.we_clk [19454]));
Q_ASSIGN U13321 ( .B(clk), .A(\g.we_clk [19453]));
Q_ASSIGN U13322 ( .B(clk), .A(\g.we_clk [19452]));
Q_ASSIGN U13323 ( .B(clk), .A(\g.we_clk [19451]));
Q_ASSIGN U13324 ( .B(clk), .A(\g.we_clk [19450]));
Q_ASSIGN U13325 ( .B(clk), .A(\g.we_clk [19449]));
Q_ASSIGN U13326 ( .B(clk), .A(\g.we_clk [19448]));
Q_ASSIGN U13327 ( .B(clk), .A(\g.we_clk [19447]));
Q_ASSIGN U13328 ( .B(clk), .A(\g.we_clk [19446]));
Q_ASSIGN U13329 ( .B(clk), .A(\g.we_clk [19445]));
Q_ASSIGN U13330 ( .B(clk), .A(\g.we_clk [19444]));
Q_ASSIGN U13331 ( .B(clk), .A(\g.we_clk [19443]));
Q_ASSIGN U13332 ( .B(clk), .A(\g.we_clk [19442]));
Q_ASSIGN U13333 ( .B(clk), .A(\g.we_clk [19441]));
Q_ASSIGN U13334 ( .B(clk), .A(\g.we_clk [19440]));
Q_ASSIGN U13335 ( .B(clk), .A(\g.we_clk [19439]));
Q_ASSIGN U13336 ( .B(clk), .A(\g.we_clk [19438]));
Q_ASSIGN U13337 ( .B(clk), .A(\g.we_clk [19437]));
Q_ASSIGN U13338 ( .B(clk), .A(\g.we_clk [19436]));
Q_ASSIGN U13339 ( .B(clk), .A(\g.we_clk [19435]));
Q_ASSIGN U13340 ( .B(clk), .A(\g.we_clk [19434]));
Q_ASSIGN U13341 ( .B(clk), .A(\g.we_clk [19433]));
Q_ASSIGN U13342 ( .B(clk), .A(\g.we_clk [19432]));
Q_ASSIGN U13343 ( .B(clk), .A(\g.we_clk [19431]));
Q_ASSIGN U13344 ( .B(clk), .A(\g.we_clk [19430]));
Q_ASSIGN U13345 ( .B(clk), .A(\g.we_clk [19429]));
Q_ASSIGN U13346 ( .B(clk), .A(\g.we_clk [19428]));
Q_ASSIGN U13347 ( .B(clk), .A(\g.we_clk [19427]));
Q_ASSIGN U13348 ( .B(clk), .A(\g.we_clk [19426]));
Q_ASSIGN U13349 ( .B(clk), .A(\g.we_clk [19425]));
Q_ASSIGN U13350 ( .B(clk), .A(\g.we_clk [19424]));
Q_ASSIGN U13351 ( .B(clk), .A(\g.we_clk [19423]));
Q_ASSIGN U13352 ( .B(clk), .A(\g.we_clk [19422]));
Q_ASSIGN U13353 ( .B(clk), .A(\g.we_clk [19421]));
Q_ASSIGN U13354 ( .B(clk), .A(\g.we_clk [19420]));
Q_ASSIGN U13355 ( .B(clk), .A(\g.we_clk [19419]));
Q_ASSIGN U13356 ( .B(clk), .A(\g.we_clk [19418]));
Q_ASSIGN U13357 ( .B(clk), .A(\g.we_clk [19417]));
Q_ASSIGN U13358 ( .B(clk), .A(\g.we_clk [19416]));
Q_ASSIGN U13359 ( .B(clk), .A(\g.we_clk [19415]));
Q_ASSIGN U13360 ( .B(clk), .A(\g.we_clk [19414]));
Q_ASSIGN U13361 ( .B(clk), .A(\g.we_clk [19413]));
Q_ASSIGN U13362 ( .B(clk), .A(\g.we_clk [19412]));
Q_ASSIGN U13363 ( .B(clk), .A(\g.we_clk [19411]));
Q_ASSIGN U13364 ( .B(clk), .A(\g.we_clk [19410]));
Q_ASSIGN U13365 ( .B(clk), .A(\g.we_clk [19409]));
Q_ASSIGN U13366 ( .B(clk), .A(\g.we_clk [19408]));
Q_ASSIGN U13367 ( .B(clk), .A(\g.we_clk [19407]));
Q_ASSIGN U13368 ( .B(clk), .A(\g.we_clk [19406]));
Q_ASSIGN U13369 ( .B(clk), .A(\g.we_clk [19405]));
Q_ASSIGN U13370 ( .B(clk), .A(\g.we_clk [19404]));
Q_ASSIGN U13371 ( .B(clk), .A(\g.we_clk [19403]));
Q_ASSIGN U13372 ( .B(clk), .A(\g.we_clk [19402]));
Q_ASSIGN U13373 ( .B(clk), .A(\g.we_clk [19401]));
Q_ASSIGN U13374 ( .B(clk), .A(\g.we_clk [19400]));
Q_ASSIGN U13375 ( .B(clk), .A(\g.we_clk [19399]));
Q_ASSIGN U13376 ( .B(clk), .A(\g.we_clk [19398]));
Q_ASSIGN U13377 ( .B(clk), .A(\g.we_clk [19397]));
Q_ASSIGN U13378 ( .B(clk), .A(\g.we_clk [19396]));
Q_ASSIGN U13379 ( .B(clk), .A(\g.we_clk [19395]));
Q_ASSIGN U13380 ( .B(clk), .A(\g.we_clk [19394]));
Q_ASSIGN U13381 ( .B(clk), .A(\g.we_clk [19393]));
Q_ASSIGN U13382 ( .B(clk), .A(\g.we_clk [19392]));
Q_ASSIGN U13383 ( .B(clk), .A(\g.we_clk [19391]));
Q_ASSIGN U13384 ( .B(clk), .A(\g.we_clk [19390]));
Q_ASSIGN U13385 ( .B(clk), .A(\g.we_clk [19389]));
Q_ASSIGN U13386 ( .B(clk), .A(\g.we_clk [19388]));
Q_ASSIGN U13387 ( .B(clk), .A(\g.we_clk [19387]));
Q_ASSIGN U13388 ( .B(clk), .A(\g.we_clk [19386]));
Q_ASSIGN U13389 ( .B(clk), .A(\g.we_clk [19385]));
Q_ASSIGN U13390 ( .B(clk), .A(\g.we_clk [19384]));
Q_ASSIGN U13391 ( .B(clk), .A(\g.we_clk [19383]));
Q_ASSIGN U13392 ( .B(clk), .A(\g.we_clk [19382]));
Q_ASSIGN U13393 ( .B(clk), .A(\g.we_clk [19381]));
Q_ASSIGN U13394 ( .B(clk), .A(\g.we_clk [19380]));
Q_ASSIGN U13395 ( .B(clk), .A(\g.we_clk [19379]));
Q_ASSIGN U13396 ( .B(clk), .A(\g.we_clk [19378]));
Q_ASSIGN U13397 ( .B(clk), .A(\g.we_clk [19377]));
Q_ASSIGN U13398 ( .B(clk), .A(\g.we_clk [19376]));
Q_ASSIGN U13399 ( .B(clk), .A(\g.we_clk [19375]));
Q_ASSIGN U13400 ( .B(clk), .A(\g.we_clk [19374]));
Q_ASSIGN U13401 ( .B(clk), .A(\g.we_clk [19373]));
Q_ASSIGN U13402 ( .B(clk), .A(\g.we_clk [19372]));
Q_ASSIGN U13403 ( .B(clk), .A(\g.we_clk [19371]));
Q_ASSIGN U13404 ( .B(clk), .A(\g.we_clk [19370]));
Q_ASSIGN U13405 ( .B(clk), .A(\g.we_clk [19369]));
Q_ASSIGN U13406 ( .B(clk), .A(\g.we_clk [19368]));
Q_ASSIGN U13407 ( .B(clk), .A(\g.we_clk [19367]));
Q_ASSIGN U13408 ( .B(clk), .A(\g.we_clk [19366]));
Q_ASSIGN U13409 ( .B(clk), .A(\g.we_clk [19365]));
Q_ASSIGN U13410 ( .B(clk), .A(\g.we_clk [19364]));
Q_ASSIGN U13411 ( .B(clk), .A(\g.we_clk [19363]));
Q_ASSIGN U13412 ( .B(clk), .A(\g.we_clk [19362]));
Q_ASSIGN U13413 ( .B(clk), .A(\g.we_clk [19361]));
Q_ASSIGN U13414 ( .B(clk), .A(\g.we_clk [19360]));
Q_ASSIGN U13415 ( .B(clk), .A(\g.we_clk [19359]));
Q_ASSIGN U13416 ( .B(clk), .A(\g.we_clk [19358]));
Q_ASSIGN U13417 ( .B(clk), .A(\g.we_clk [19357]));
Q_ASSIGN U13418 ( .B(clk), .A(\g.we_clk [19356]));
Q_ASSIGN U13419 ( .B(clk), .A(\g.we_clk [19355]));
Q_ASSIGN U13420 ( .B(clk), .A(\g.we_clk [19354]));
Q_ASSIGN U13421 ( .B(clk), .A(\g.we_clk [19353]));
Q_ASSIGN U13422 ( .B(clk), .A(\g.we_clk [19352]));
Q_ASSIGN U13423 ( .B(clk), .A(\g.we_clk [19351]));
Q_ASSIGN U13424 ( .B(clk), .A(\g.we_clk [19350]));
Q_ASSIGN U13425 ( .B(clk), .A(\g.we_clk [19349]));
Q_ASSIGN U13426 ( .B(clk), .A(\g.we_clk [19348]));
Q_ASSIGN U13427 ( .B(clk), .A(\g.we_clk [19347]));
Q_ASSIGN U13428 ( .B(clk), .A(\g.we_clk [19346]));
Q_ASSIGN U13429 ( .B(clk), .A(\g.we_clk [19345]));
Q_ASSIGN U13430 ( .B(clk), .A(\g.we_clk [19344]));
Q_ASSIGN U13431 ( .B(clk), .A(\g.we_clk [19343]));
Q_ASSIGN U13432 ( .B(clk), .A(\g.we_clk [19342]));
Q_ASSIGN U13433 ( .B(clk), .A(\g.we_clk [19341]));
Q_ASSIGN U13434 ( .B(clk), .A(\g.we_clk [19340]));
Q_ASSIGN U13435 ( .B(clk), .A(\g.we_clk [19339]));
Q_ASSIGN U13436 ( .B(clk), .A(\g.we_clk [19338]));
Q_ASSIGN U13437 ( .B(clk), .A(\g.we_clk [19337]));
Q_ASSIGN U13438 ( .B(clk), .A(\g.we_clk [19336]));
Q_ASSIGN U13439 ( .B(clk), .A(\g.we_clk [19335]));
Q_ASSIGN U13440 ( .B(clk), .A(\g.we_clk [19334]));
Q_ASSIGN U13441 ( .B(clk), .A(\g.we_clk [19333]));
Q_ASSIGN U13442 ( .B(clk), .A(\g.we_clk [19332]));
Q_ASSIGN U13443 ( .B(clk), .A(\g.we_clk [19331]));
Q_ASSIGN U13444 ( .B(clk), .A(\g.we_clk [19330]));
Q_ASSIGN U13445 ( .B(clk), .A(\g.we_clk [19329]));
Q_ASSIGN U13446 ( .B(clk), .A(\g.we_clk [19328]));
Q_ASSIGN U13447 ( .B(clk), .A(\g.we_clk [19327]));
Q_ASSIGN U13448 ( .B(clk), .A(\g.we_clk [19326]));
Q_ASSIGN U13449 ( .B(clk), .A(\g.we_clk [19325]));
Q_ASSIGN U13450 ( .B(clk), .A(\g.we_clk [19324]));
Q_ASSIGN U13451 ( .B(clk), .A(\g.we_clk [19323]));
Q_ASSIGN U13452 ( .B(clk), .A(\g.we_clk [19322]));
Q_ASSIGN U13453 ( .B(clk), .A(\g.we_clk [19321]));
Q_ASSIGN U13454 ( .B(clk), .A(\g.we_clk [19320]));
Q_ASSIGN U13455 ( .B(clk), .A(\g.we_clk [19319]));
Q_ASSIGN U13456 ( .B(clk), .A(\g.we_clk [19318]));
Q_ASSIGN U13457 ( .B(clk), .A(\g.we_clk [19317]));
Q_ASSIGN U13458 ( .B(clk), .A(\g.we_clk [19316]));
Q_ASSIGN U13459 ( .B(clk), .A(\g.we_clk [19315]));
Q_ASSIGN U13460 ( .B(clk), .A(\g.we_clk [19314]));
Q_ASSIGN U13461 ( .B(clk), .A(\g.we_clk [19313]));
Q_ASSIGN U13462 ( .B(clk), .A(\g.we_clk [19312]));
Q_ASSIGN U13463 ( .B(clk), .A(\g.we_clk [19311]));
Q_ASSIGN U13464 ( .B(clk), .A(\g.we_clk [19310]));
Q_ASSIGN U13465 ( .B(clk), .A(\g.we_clk [19309]));
Q_ASSIGN U13466 ( .B(clk), .A(\g.we_clk [19308]));
Q_ASSIGN U13467 ( .B(clk), .A(\g.we_clk [19307]));
Q_ASSIGN U13468 ( .B(clk), .A(\g.we_clk [19306]));
Q_ASSIGN U13469 ( .B(clk), .A(\g.we_clk [19305]));
Q_ASSIGN U13470 ( .B(clk), .A(\g.we_clk [19304]));
Q_ASSIGN U13471 ( .B(clk), .A(\g.we_clk [19303]));
Q_ASSIGN U13472 ( .B(clk), .A(\g.we_clk [19302]));
Q_ASSIGN U13473 ( .B(clk), .A(\g.we_clk [19301]));
Q_ASSIGN U13474 ( .B(clk), .A(\g.we_clk [19300]));
Q_ASSIGN U13475 ( .B(clk), .A(\g.we_clk [19299]));
Q_ASSIGN U13476 ( .B(clk), .A(\g.we_clk [19298]));
Q_ASSIGN U13477 ( .B(clk), .A(\g.we_clk [19297]));
Q_ASSIGN U13478 ( .B(clk), .A(\g.we_clk [19296]));
Q_ASSIGN U13479 ( .B(clk), .A(\g.we_clk [19295]));
Q_ASSIGN U13480 ( .B(clk), .A(\g.we_clk [19294]));
Q_ASSIGN U13481 ( .B(clk), .A(\g.we_clk [19293]));
Q_ASSIGN U13482 ( .B(clk), .A(\g.we_clk [19292]));
Q_ASSIGN U13483 ( .B(clk), .A(\g.we_clk [19291]));
Q_ASSIGN U13484 ( .B(clk), .A(\g.we_clk [19290]));
Q_ASSIGN U13485 ( .B(clk), .A(\g.we_clk [19289]));
Q_ASSIGN U13486 ( .B(clk), .A(\g.we_clk [19288]));
Q_ASSIGN U13487 ( .B(clk), .A(\g.we_clk [19287]));
Q_ASSIGN U13488 ( .B(clk), .A(\g.we_clk [19286]));
Q_ASSIGN U13489 ( .B(clk), .A(\g.we_clk [19285]));
Q_ASSIGN U13490 ( .B(clk), .A(\g.we_clk [19284]));
Q_ASSIGN U13491 ( .B(clk), .A(\g.we_clk [19283]));
Q_ASSIGN U13492 ( .B(clk), .A(\g.we_clk [19282]));
Q_ASSIGN U13493 ( .B(clk), .A(\g.we_clk [19281]));
Q_ASSIGN U13494 ( .B(clk), .A(\g.we_clk [19280]));
Q_ASSIGN U13495 ( .B(clk), .A(\g.we_clk [19279]));
Q_ASSIGN U13496 ( .B(clk), .A(\g.we_clk [19278]));
Q_ASSIGN U13497 ( .B(clk), .A(\g.we_clk [19277]));
Q_ASSIGN U13498 ( .B(clk), .A(\g.we_clk [19276]));
Q_ASSIGN U13499 ( .B(clk), .A(\g.we_clk [19275]));
Q_ASSIGN U13500 ( .B(clk), .A(\g.we_clk [19274]));
Q_ASSIGN U13501 ( .B(clk), .A(\g.we_clk [19273]));
Q_ASSIGN U13502 ( .B(clk), .A(\g.we_clk [19272]));
Q_ASSIGN U13503 ( .B(clk), .A(\g.we_clk [19271]));
Q_ASSIGN U13504 ( .B(clk), .A(\g.we_clk [19270]));
Q_ASSIGN U13505 ( .B(clk), .A(\g.we_clk [19269]));
Q_ASSIGN U13506 ( .B(clk), .A(\g.we_clk [19268]));
Q_ASSIGN U13507 ( .B(clk), .A(\g.we_clk [19267]));
Q_ASSIGN U13508 ( .B(clk), .A(\g.we_clk [19266]));
Q_ASSIGN U13509 ( .B(clk), .A(\g.we_clk [19265]));
Q_ASSIGN U13510 ( .B(clk), .A(\g.we_clk [19264]));
Q_ASSIGN U13511 ( .B(clk), .A(\g.we_clk [19263]));
Q_ASSIGN U13512 ( .B(clk), .A(\g.we_clk [19262]));
Q_ASSIGN U13513 ( .B(clk), .A(\g.we_clk [19261]));
Q_ASSIGN U13514 ( .B(clk), .A(\g.we_clk [19260]));
Q_ASSIGN U13515 ( .B(clk), .A(\g.we_clk [19259]));
Q_ASSIGN U13516 ( .B(clk), .A(\g.we_clk [19258]));
Q_ASSIGN U13517 ( .B(clk), .A(\g.we_clk [19257]));
Q_ASSIGN U13518 ( .B(clk), .A(\g.we_clk [19256]));
Q_ASSIGN U13519 ( .B(clk), .A(\g.we_clk [19255]));
Q_ASSIGN U13520 ( .B(clk), .A(\g.we_clk [19254]));
Q_ASSIGN U13521 ( .B(clk), .A(\g.we_clk [19253]));
Q_ASSIGN U13522 ( .B(clk), .A(\g.we_clk [19252]));
Q_ASSIGN U13523 ( .B(clk), .A(\g.we_clk [19251]));
Q_ASSIGN U13524 ( .B(clk), .A(\g.we_clk [19250]));
Q_ASSIGN U13525 ( .B(clk), .A(\g.we_clk [19249]));
Q_ASSIGN U13526 ( .B(clk), .A(\g.we_clk [19248]));
Q_ASSIGN U13527 ( .B(clk), .A(\g.we_clk [19247]));
Q_ASSIGN U13528 ( .B(clk), .A(\g.we_clk [19246]));
Q_ASSIGN U13529 ( .B(clk), .A(\g.we_clk [19245]));
Q_ASSIGN U13530 ( .B(clk), .A(\g.we_clk [19244]));
Q_ASSIGN U13531 ( .B(clk), .A(\g.we_clk [19243]));
Q_ASSIGN U13532 ( .B(clk), .A(\g.we_clk [19242]));
Q_ASSIGN U13533 ( .B(clk), .A(\g.we_clk [19241]));
Q_ASSIGN U13534 ( .B(clk), .A(\g.we_clk [19240]));
Q_ASSIGN U13535 ( .B(clk), .A(\g.we_clk [19239]));
Q_ASSIGN U13536 ( .B(clk), .A(\g.we_clk [19238]));
Q_ASSIGN U13537 ( .B(clk), .A(\g.we_clk [19237]));
Q_ASSIGN U13538 ( .B(clk), .A(\g.we_clk [19236]));
Q_ASSIGN U13539 ( .B(clk), .A(\g.we_clk [19235]));
Q_ASSIGN U13540 ( .B(clk), .A(\g.we_clk [19234]));
Q_ASSIGN U13541 ( .B(clk), .A(\g.we_clk [19233]));
Q_ASSIGN U13542 ( .B(clk), .A(\g.we_clk [19232]));
Q_ASSIGN U13543 ( .B(clk), .A(\g.we_clk [19231]));
Q_ASSIGN U13544 ( .B(clk), .A(\g.we_clk [19230]));
Q_ASSIGN U13545 ( .B(clk), .A(\g.we_clk [19229]));
Q_ASSIGN U13546 ( .B(clk), .A(\g.we_clk [19228]));
Q_ASSIGN U13547 ( .B(clk), .A(\g.we_clk [19227]));
Q_ASSIGN U13548 ( .B(clk), .A(\g.we_clk [19226]));
Q_ASSIGN U13549 ( .B(clk), .A(\g.we_clk [19225]));
Q_ASSIGN U13550 ( .B(clk), .A(\g.we_clk [19224]));
Q_ASSIGN U13551 ( .B(clk), .A(\g.we_clk [19223]));
Q_ASSIGN U13552 ( .B(clk), .A(\g.we_clk [19222]));
Q_ASSIGN U13553 ( .B(clk), .A(\g.we_clk [19221]));
Q_ASSIGN U13554 ( .B(clk), .A(\g.we_clk [19220]));
Q_ASSIGN U13555 ( .B(clk), .A(\g.we_clk [19219]));
Q_ASSIGN U13556 ( .B(clk), .A(\g.we_clk [19218]));
Q_ASSIGN U13557 ( .B(clk), .A(\g.we_clk [19217]));
Q_ASSIGN U13558 ( .B(clk), .A(\g.we_clk [19216]));
Q_ASSIGN U13559 ( .B(clk), .A(\g.we_clk [19215]));
Q_ASSIGN U13560 ( .B(clk), .A(\g.we_clk [19214]));
Q_ASSIGN U13561 ( .B(clk), .A(\g.we_clk [19213]));
Q_ASSIGN U13562 ( .B(clk), .A(\g.we_clk [19212]));
Q_ASSIGN U13563 ( .B(clk), .A(\g.we_clk [19211]));
Q_ASSIGN U13564 ( .B(clk), .A(\g.we_clk [19210]));
Q_ASSIGN U13565 ( .B(clk), .A(\g.we_clk [19209]));
Q_ASSIGN U13566 ( .B(clk), .A(\g.we_clk [19208]));
Q_ASSIGN U13567 ( .B(clk), .A(\g.we_clk [19207]));
Q_ASSIGN U13568 ( .B(clk), .A(\g.we_clk [19206]));
Q_ASSIGN U13569 ( .B(clk), .A(\g.we_clk [19205]));
Q_ASSIGN U13570 ( .B(clk), .A(\g.we_clk [19204]));
Q_ASSIGN U13571 ( .B(clk), .A(\g.we_clk [19203]));
Q_ASSIGN U13572 ( .B(clk), .A(\g.we_clk [19202]));
Q_ASSIGN U13573 ( .B(clk), .A(\g.we_clk [19201]));
Q_ASSIGN U13574 ( .B(clk), .A(\g.we_clk [19200]));
Q_ASSIGN U13575 ( .B(clk), .A(\g.we_clk [19199]));
Q_ASSIGN U13576 ( .B(clk), .A(\g.we_clk [19198]));
Q_ASSIGN U13577 ( .B(clk), .A(\g.we_clk [19197]));
Q_ASSIGN U13578 ( .B(clk), .A(\g.we_clk [19196]));
Q_ASSIGN U13579 ( .B(clk), .A(\g.we_clk [19195]));
Q_ASSIGN U13580 ( .B(clk), .A(\g.we_clk [19194]));
Q_ASSIGN U13581 ( .B(clk), .A(\g.we_clk [19193]));
Q_ASSIGN U13582 ( .B(clk), .A(\g.we_clk [19192]));
Q_ASSIGN U13583 ( .B(clk), .A(\g.we_clk [19191]));
Q_ASSIGN U13584 ( .B(clk), .A(\g.we_clk [19190]));
Q_ASSIGN U13585 ( .B(clk), .A(\g.we_clk [19189]));
Q_ASSIGN U13586 ( .B(clk), .A(\g.we_clk [19188]));
Q_ASSIGN U13587 ( .B(clk), .A(\g.we_clk [19187]));
Q_ASSIGN U13588 ( .B(clk), .A(\g.we_clk [19186]));
Q_ASSIGN U13589 ( .B(clk), .A(\g.we_clk [19185]));
Q_ASSIGN U13590 ( .B(clk), .A(\g.we_clk [19184]));
Q_ASSIGN U13591 ( .B(clk), .A(\g.we_clk [19183]));
Q_ASSIGN U13592 ( .B(clk), .A(\g.we_clk [19182]));
Q_ASSIGN U13593 ( .B(clk), .A(\g.we_clk [19181]));
Q_ASSIGN U13594 ( .B(clk), .A(\g.we_clk [19180]));
Q_ASSIGN U13595 ( .B(clk), .A(\g.we_clk [19179]));
Q_ASSIGN U13596 ( .B(clk), .A(\g.we_clk [19178]));
Q_ASSIGN U13597 ( .B(clk), .A(\g.we_clk [19177]));
Q_ASSIGN U13598 ( .B(clk), .A(\g.we_clk [19176]));
Q_ASSIGN U13599 ( .B(clk), .A(\g.we_clk [19175]));
Q_ASSIGN U13600 ( .B(clk), .A(\g.we_clk [19174]));
Q_ASSIGN U13601 ( .B(clk), .A(\g.we_clk [19173]));
Q_ASSIGN U13602 ( .B(clk), .A(\g.we_clk [19172]));
Q_ASSIGN U13603 ( .B(clk), .A(\g.we_clk [19171]));
Q_ASSIGN U13604 ( .B(clk), .A(\g.we_clk [19170]));
Q_ASSIGN U13605 ( .B(clk), .A(\g.we_clk [19169]));
Q_ASSIGN U13606 ( .B(clk), .A(\g.we_clk [19168]));
Q_ASSIGN U13607 ( .B(clk), .A(\g.we_clk [19167]));
Q_ASSIGN U13608 ( .B(clk), .A(\g.we_clk [19166]));
Q_ASSIGN U13609 ( .B(clk), .A(\g.we_clk [19165]));
Q_ASSIGN U13610 ( .B(clk), .A(\g.we_clk [19164]));
Q_ASSIGN U13611 ( .B(clk), .A(\g.we_clk [19163]));
Q_ASSIGN U13612 ( .B(clk), .A(\g.we_clk [19162]));
Q_ASSIGN U13613 ( .B(clk), .A(\g.we_clk [19161]));
Q_ASSIGN U13614 ( .B(clk), .A(\g.we_clk [19160]));
Q_ASSIGN U13615 ( .B(clk), .A(\g.we_clk [19159]));
Q_ASSIGN U13616 ( .B(clk), .A(\g.we_clk [19158]));
Q_ASSIGN U13617 ( .B(clk), .A(\g.we_clk [19157]));
Q_ASSIGN U13618 ( .B(clk), .A(\g.we_clk [19156]));
Q_ASSIGN U13619 ( .B(clk), .A(\g.we_clk [19155]));
Q_ASSIGN U13620 ( .B(clk), .A(\g.we_clk [19154]));
Q_ASSIGN U13621 ( .B(clk), .A(\g.we_clk [19153]));
Q_ASSIGN U13622 ( .B(clk), .A(\g.we_clk [19152]));
Q_ASSIGN U13623 ( .B(clk), .A(\g.we_clk [19151]));
Q_ASSIGN U13624 ( .B(clk), .A(\g.we_clk [19150]));
Q_ASSIGN U13625 ( .B(clk), .A(\g.we_clk [19149]));
Q_ASSIGN U13626 ( .B(clk), .A(\g.we_clk [19148]));
Q_ASSIGN U13627 ( .B(clk), .A(\g.we_clk [19147]));
Q_ASSIGN U13628 ( .B(clk), .A(\g.we_clk [19146]));
Q_ASSIGN U13629 ( .B(clk), .A(\g.we_clk [19145]));
Q_ASSIGN U13630 ( .B(clk), .A(\g.we_clk [19144]));
Q_ASSIGN U13631 ( .B(clk), .A(\g.we_clk [19143]));
Q_ASSIGN U13632 ( .B(clk), .A(\g.we_clk [19142]));
Q_ASSIGN U13633 ( .B(clk), .A(\g.we_clk [19141]));
Q_ASSIGN U13634 ( .B(clk), .A(\g.we_clk [19140]));
Q_ASSIGN U13635 ( .B(clk), .A(\g.we_clk [19139]));
Q_ASSIGN U13636 ( .B(clk), .A(\g.we_clk [19138]));
Q_ASSIGN U13637 ( .B(clk), .A(\g.we_clk [19137]));
Q_ASSIGN U13638 ( .B(clk), .A(\g.we_clk [19136]));
Q_ASSIGN U13639 ( .B(clk), .A(\g.we_clk [19135]));
Q_ASSIGN U13640 ( .B(clk), .A(\g.we_clk [19134]));
Q_ASSIGN U13641 ( .B(clk), .A(\g.we_clk [19133]));
Q_ASSIGN U13642 ( .B(clk), .A(\g.we_clk [19132]));
Q_ASSIGN U13643 ( .B(clk), .A(\g.we_clk [19131]));
Q_ASSIGN U13644 ( .B(clk), .A(\g.we_clk [19130]));
Q_ASSIGN U13645 ( .B(clk), .A(\g.we_clk [19129]));
Q_ASSIGN U13646 ( .B(clk), .A(\g.we_clk [19128]));
Q_ASSIGN U13647 ( .B(clk), .A(\g.we_clk [19127]));
Q_ASSIGN U13648 ( .B(clk), .A(\g.we_clk [19126]));
Q_ASSIGN U13649 ( .B(clk), .A(\g.we_clk [19125]));
Q_ASSIGN U13650 ( .B(clk), .A(\g.we_clk [19124]));
Q_ASSIGN U13651 ( .B(clk), .A(\g.we_clk [19123]));
Q_ASSIGN U13652 ( .B(clk), .A(\g.we_clk [19122]));
Q_ASSIGN U13653 ( .B(clk), .A(\g.we_clk [19121]));
Q_ASSIGN U13654 ( .B(clk), .A(\g.we_clk [19120]));
Q_ASSIGN U13655 ( .B(clk), .A(\g.we_clk [19119]));
Q_ASSIGN U13656 ( .B(clk), .A(\g.we_clk [19118]));
Q_ASSIGN U13657 ( .B(clk), .A(\g.we_clk [19117]));
Q_ASSIGN U13658 ( .B(clk), .A(\g.we_clk [19116]));
Q_ASSIGN U13659 ( .B(clk), .A(\g.we_clk [19115]));
Q_ASSIGN U13660 ( .B(clk), .A(\g.we_clk [19114]));
Q_ASSIGN U13661 ( .B(clk), .A(\g.we_clk [19113]));
Q_ASSIGN U13662 ( .B(clk), .A(\g.we_clk [19112]));
Q_ASSIGN U13663 ( .B(clk), .A(\g.we_clk [19111]));
Q_ASSIGN U13664 ( .B(clk), .A(\g.we_clk [19110]));
Q_ASSIGN U13665 ( .B(clk), .A(\g.we_clk [19109]));
Q_ASSIGN U13666 ( .B(clk), .A(\g.we_clk [19108]));
Q_ASSIGN U13667 ( .B(clk), .A(\g.we_clk [19107]));
Q_ASSIGN U13668 ( .B(clk), .A(\g.we_clk [19106]));
Q_ASSIGN U13669 ( .B(clk), .A(\g.we_clk [19105]));
Q_ASSIGN U13670 ( .B(clk), .A(\g.we_clk [19104]));
Q_ASSIGN U13671 ( .B(clk), .A(\g.we_clk [19103]));
Q_ASSIGN U13672 ( .B(clk), .A(\g.we_clk [19102]));
Q_ASSIGN U13673 ( .B(clk), .A(\g.we_clk [19101]));
Q_ASSIGN U13674 ( .B(clk), .A(\g.we_clk [19100]));
Q_ASSIGN U13675 ( .B(clk), .A(\g.we_clk [19099]));
Q_ASSIGN U13676 ( .B(clk), .A(\g.we_clk [19098]));
Q_ASSIGN U13677 ( .B(clk), .A(\g.we_clk [19097]));
Q_ASSIGN U13678 ( .B(clk), .A(\g.we_clk [19096]));
Q_ASSIGN U13679 ( .B(clk), .A(\g.we_clk [19095]));
Q_ASSIGN U13680 ( .B(clk), .A(\g.we_clk [19094]));
Q_ASSIGN U13681 ( .B(clk), .A(\g.we_clk [19093]));
Q_ASSIGN U13682 ( .B(clk), .A(\g.we_clk [19092]));
Q_ASSIGN U13683 ( .B(clk), .A(\g.we_clk [19091]));
Q_ASSIGN U13684 ( .B(clk), .A(\g.we_clk [19090]));
Q_ASSIGN U13685 ( .B(clk), .A(\g.we_clk [19089]));
Q_ASSIGN U13686 ( .B(clk), .A(\g.we_clk [19088]));
Q_ASSIGN U13687 ( .B(clk), .A(\g.we_clk [19087]));
Q_ASSIGN U13688 ( .B(clk), .A(\g.we_clk [19086]));
Q_ASSIGN U13689 ( .B(clk), .A(\g.we_clk [19085]));
Q_ASSIGN U13690 ( .B(clk), .A(\g.we_clk [19084]));
Q_ASSIGN U13691 ( .B(clk), .A(\g.we_clk [19083]));
Q_ASSIGN U13692 ( .B(clk), .A(\g.we_clk [19082]));
Q_ASSIGN U13693 ( .B(clk), .A(\g.we_clk [19081]));
Q_ASSIGN U13694 ( .B(clk), .A(\g.we_clk [19080]));
Q_ASSIGN U13695 ( .B(clk), .A(\g.we_clk [19079]));
Q_ASSIGN U13696 ( .B(clk), .A(\g.we_clk [19078]));
Q_ASSIGN U13697 ( .B(clk), .A(\g.we_clk [19077]));
Q_ASSIGN U13698 ( .B(clk), .A(\g.we_clk [19076]));
Q_ASSIGN U13699 ( .B(clk), .A(\g.we_clk [19075]));
Q_ASSIGN U13700 ( .B(clk), .A(\g.we_clk [19074]));
Q_ASSIGN U13701 ( .B(clk), .A(\g.we_clk [19073]));
Q_ASSIGN U13702 ( .B(clk), .A(\g.we_clk [19072]));
Q_ASSIGN U13703 ( .B(clk), .A(\g.we_clk [19071]));
Q_ASSIGN U13704 ( .B(clk), .A(\g.we_clk [19070]));
Q_ASSIGN U13705 ( .B(clk), .A(\g.we_clk [19069]));
Q_ASSIGN U13706 ( .B(clk), .A(\g.we_clk [19068]));
Q_ASSIGN U13707 ( .B(clk), .A(\g.we_clk [19067]));
Q_ASSIGN U13708 ( .B(clk), .A(\g.we_clk [19066]));
Q_ASSIGN U13709 ( .B(clk), .A(\g.we_clk [19065]));
Q_ASSIGN U13710 ( .B(clk), .A(\g.we_clk [19064]));
Q_ASSIGN U13711 ( .B(clk), .A(\g.we_clk [19063]));
Q_ASSIGN U13712 ( .B(clk), .A(\g.we_clk [19062]));
Q_ASSIGN U13713 ( .B(clk), .A(\g.we_clk [19061]));
Q_ASSIGN U13714 ( .B(clk), .A(\g.we_clk [19060]));
Q_ASSIGN U13715 ( .B(clk), .A(\g.we_clk [19059]));
Q_ASSIGN U13716 ( .B(clk), .A(\g.we_clk [19058]));
Q_ASSIGN U13717 ( .B(clk), .A(\g.we_clk [19057]));
Q_ASSIGN U13718 ( .B(clk), .A(\g.we_clk [19056]));
Q_ASSIGN U13719 ( .B(clk), .A(\g.we_clk [19055]));
Q_ASSIGN U13720 ( .B(clk), .A(\g.we_clk [19054]));
Q_ASSIGN U13721 ( .B(clk), .A(\g.we_clk [19053]));
Q_ASSIGN U13722 ( .B(clk), .A(\g.we_clk [19052]));
Q_ASSIGN U13723 ( .B(clk), .A(\g.we_clk [19051]));
Q_ASSIGN U13724 ( .B(clk), .A(\g.we_clk [19050]));
Q_ASSIGN U13725 ( .B(clk), .A(\g.we_clk [19049]));
Q_ASSIGN U13726 ( .B(clk), .A(\g.we_clk [19048]));
Q_ASSIGN U13727 ( .B(clk), .A(\g.we_clk [19047]));
Q_ASSIGN U13728 ( .B(clk), .A(\g.we_clk [19046]));
Q_ASSIGN U13729 ( .B(clk), .A(\g.we_clk [19045]));
Q_ASSIGN U13730 ( .B(clk), .A(\g.we_clk [19044]));
Q_ASSIGN U13731 ( .B(clk), .A(\g.we_clk [19043]));
Q_ASSIGN U13732 ( .B(clk), .A(\g.we_clk [19042]));
Q_ASSIGN U13733 ( .B(clk), .A(\g.we_clk [19041]));
Q_ASSIGN U13734 ( .B(clk), .A(\g.we_clk [19040]));
Q_ASSIGN U13735 ( .B(clk), .A(\g.we_clk [19039]));
Q_ASSIGN U13736 ( .B(clk), .A(\g.we_clk [19038]));
Q_ASSIGN U13737 ( .B(clk), .A(\g.we_clk [19037]));
Q_ASSIGN U13738 ( .B(clk), .A(\g.we_clk [19036]));
Q_ASSIGN U13739 ( .B(clk), .A(\g.we_clk [19035]));
Q_ASSIGN U13740 ( .B(clk), .A(\g.we_clk [19034]));
Q_ASSIGN U13741 ( .B(clk), .A(\g.we_clk [19033]));
Q_ASSIGN U13742 ( .B(clk), .A(\g.we_clk [19032]));
Q_ASSIGN U13743 ( .B(clk), .A(\g.we_clk [19031]));
Q_ASSIGN U13744 ( .B(clk), .A(\g.we_clk [19030]));
Q_ASSIGN U13745 ( .B(clk), .A(\g.we_clk [19029]));
Q_ASSIGN U13746 ( .B(clk), .A(\g.we_clk [19028]));
Q_ASSIGN U13747 ( .B(clk), .A(\g.we_clk [19027]));
Q_ASSIGN U13748 ( .B(clk), .A(\g.we_clk [19026]));
Q_ASSIGN U13749 ( .B(clk), .A(\g.we_clk [19025]));
Q_ASSIGN U13750 ( .B(clk), .A(\g.we_clk [19024]));
Q_ASSIGN U13751 ( .B(clk), .A(\g.we_clk [19023]));
Q_ASSIGN U13752 ( .B(clk), .A(\g.we_clk [19022]));
Q_ASSIGN U13753 ( .B(clk), .A(\g.we_clk [19021]));
Q_ASSIGN U13754 ( .B(clk), .A(\g.we_clk [19020]));
Q_ASSIGN U13755 ( .B(clk), .A(\g.we_clk [19019]));
Q_ASSIGN U13756 ( .B(clk), .A(\g.we_clk [19018]));
Q_ASSIGN U13757 ( .B(clk), .A(\g.we_clk [19017]));
Q_ASSIGN U13758 ( .B(clk), .A(\g.we_clk [19016]));
Q_ASSIGN U13759 ( .B(clk), .A(\g.we_clk [19015]));
Q_ASSIGN U13760 ( .B(clk), .A(\g.we_clk [19014]));
Q_ASSIGN U13761 ( .B(clk), .A(\g.we_clk [19013]));
Q_ASSIGN U13762 ( .B(clk), .A(\g.we_clk [19012]));
Q_ASSIGN U13763 ( .B(clk), .A(\g.we_clk [19011]));
Q_ASSIGN U13764 ( .B(clk), .A(\g.we_clk [19010]));
Q_ASSIGN U13765 ( .B(clk), .A(\g.we_clk [19009]));
Q_ASSIGN U13766 ( .B(clk), .A(\g.we_clk [19008]));
Q_ASSIGN U13767 ( .B(clk), .A(\g.we_clk [19007]));
Q_ASSIGN U13768 ( .B(clk), .A(\g.we_clk [19006]));
Q_ASSIGN U13769 ( .B(clk), .A(\g.we_clk [19005]));
Q_ASSIGN U13770 ( .B(clk), .A(\g.we_clk [19004]));
Q_ASSIGN U13771 ( .B(clk), .A(\g.we_clk [19003]));
Q_ASSIGN U13772 ( .B(clk), .A(\g.we_clk [19002]));
Q_ASSIGN U13773 ( .B(clk), .A(\g.we_clk [19001]));
Q_ASSIGN U13774 ( .B(clk), .A(\g.we_clk [19000]));
Q_ASSIGN U13775 ( .B(clk), .A(\g.we_clk [18999]));
Q_ASSIGN U13776 ( .B(clk), .A(\g.we_clk [18998]));
Q_ASSIGN U13777 ( .B(clk), .A(\g.we_clk [18997]));
Q_ASSIGN U13778 ( .B(clk), .A(\g.we_clk [18996]));
Q_ASSIGN U13779 ( .B(clk), .A(\g.we_clk [18995]));
Q_ASSIGN U13780 ( .B(clk), .A(\g.we_clk [18994]));
Q_ASSIGN U13781 ( .B(clk), .A(\g.we_clk [18993]));
Q_ASSIGN U13782 ( .B(clk), .A(\g.we_clk [18992]));
Q_ASSIGN U13783 ( .B(clk), .A(\g.we_clk [18991]));
Q_ASSIGN U13784 ( .B(clk), .A(\g.we_clk [18990]));
Q_ASSIGN U13785 ( .B(clk), .A(\g.we_clk [18989]));
Q_ASSIGN U13786 ( .B(clk), .A(\g.we_clk [18988]));
Q_ASSIGN U13787 ( .B(clk), .A(\g.we_clk [18987]));
Q_ASSIGN U13788 ( .B(clk), .A(\g.we_clk [18986]));
Q_ASSIGN U13789 ( .B(clk), .A(\g.we_clk [18985]));
Q_ASSIGN U13790 ( .B(clk), .A(\g.we_clk [18984]));
Q_ASSIGN U13791 ( .B(clk), .A(\g.we_clk [18983]));
Q_ASSIGN U13792 ( .B(clk), .A(\g.we_clk [18982]));
Q_ASSIGN U13793 ( .B(clk), .A(\g.we_clk [18981]));
Q_ASSIGN U13794 ( .B(clk), .A(\g.we_clk [18980]));
Q_ASSIGN U13795 ( .B(clk), .A(\g.we_clk [18979]));
Q_ASSIGN U13796 ( .B(clk), .A(\g.we_clk [18978]));
Q_ASSIGN U13797 ( .B(clk), .A(\g.we_clk [18977]));
Q_ASSIGN U13798 ( .B(clk), .A(\g.we_clk [18976]));
Q_ASSIGN U13799 ( .B(clk), .A(\g.we_clk [18975]));
Q_ASSIGN U13800 ( .B(clk), .A(\g.we_clk [18974]));
Q_ASSIGN U13801 ( .B(clk), .A(\g.we_clk [18973]));
Q_ASSIGN U13802 ( .B(clk), .A(\g.we_clk [18972]));
Q_ASSIGN U13803 ( .B(clk), .A(\g.we_clk [18971]));
Q_ASSIGN U13804 ( .B(clk), .A(\g.we_clk [18970]));
Q_ASSIGN U13805 ( .B(clk), .A(\g.we_clk [18969]));
Q_ASSIGN U13806 ( .B(clk), .A(\g.we_clk [18968]));
Q_ASSIGN U13807 ( .B(clk), .A(\g.we_clk [18967]));
Q_ASSIGN U13808 ( .B(clk), .A(\g.we_clk [18966]));
Q_ASSIGN U13809 ( .B(clk), .A(\g.we_clk [18965]));
Q_ASSIGN U13810 ( .B(clk), .A(\g.we_clk [18964]));
Q_ASSIGN U13811 ( .B(clk), .A(\g.we_clk [18963]));
Q_ASSIGN U13812 ( .B(clk), .A(\g.we_clk [18962]));
Q_ASSIGN U13813 ( .B(clk), .A(\g.we_clk [18961]));
Q_ASSIGN U13814 ( .B(clk), .A(\g.we_clk [18960]));
Q_ASSIGN U13815 ( .B(clk), .A(\g.we_clk [18959]));
Q_ASSIGN U13816 ( .B(clk), .A(\g.we_clk [18958]));
Q_ASSIGN U13817 ( .B(clk), .A(\g.we_clk [18957]));
Q_ASSIGN U13818 ( .B(clk), .A(\g.we_clk [18956]));
Q_ASSIGN U13819 ( .B(clk), .A(\g.we_clk [18955]));
Q_ASSIGN U13820 ( .B(clk), .A(\g.we_clk [18954]));
Q_ASSIGN U13821 ( .B(clk), .A(\g.we_clk [18953]));
Q_ASSIGN U13822 ( .B(clk), .A(\g.we_clk [18952]));
Q_ASSIGN U13823 ( .B(clk), .A(\g.we_clk [18951]));
Q_ASSIGN U13824 ( .B(clk), .A(\g.we_clk [18950]));
Q_ASSIGN U13825 ( .B(clk), .A(\g.we_clk [18949]));
Q_ASSIGN U13826 ( .B(clk), .A(\g.we_clk [18948]));
Q_ASSIGN U13827 ( .B(clk), .A(\g.we_clk [18947]));
Q_ASSIGN U13828 ( .B(clk), .A(\g.we_clk [18946]));
Q_ASSIGN U13829 ( .B(clk), .A(\g.we_clk [18945]));
Q_ASSIGN U13830 ( .B(clk), .A(\g.we_clk [18944]));
Q_ASSIGN U13831 ( .B(clk), .A(\g.we_clk [18943]));
Q_ASSIGN U13832 ( .B(clk), .A(\g.we_clk [18942]));
Q_ASSIGN U13833 ( .B(clk), .A(\g.we_clk [18941]));
Q_ASSIGN U13834 ( .B(clk), .A(\g.we_clk [18940]));
Q_ASSIGN U13835 ( .B(clk), .A(\g.we_clk [18939]));
Q_ASSIGN U13836 ( .B(clk), .A(\g.we_clk [18938]));
Q_ASSIGN U13837 ( .B(clk), .A(\g.we_clk [18937]));
Q_ASSIGN U13838 ( .B(clk), .A(\g.we_clk [18936]));
Q_ASSIGN U13839 ( .B(clk), .A(\g.we_clk [18935]));
Q_ASSIGN U13840 ( .B(clk), .A(\g.we_clk [18934]));
Q_ASSIGN U13841 ( .B(clk), .A(\g.we_clk [18933]));
Q_ASSIGN U13842 ( .B(clk), .A(\g.we_clk [18932]));
Q_ASSIGN U13843 ( .B(clk), .A(\g.we_clk [18931]));
Q_ASSIGN U13844 ( .B(clk), .A(\g.we_clk [18930]));
Q_ASSIGN U13845 ( .B(clk), .A(\g.we_clk [18929]));
Q_ASSIGN U13846 ( .B(clk), .A(\g.we_clk [18928]));
Q_ASSIGN U13847 ( .B(clk), .A(\g.we_clk [18927]));
Q_ASSIGN U13848 ( .B(clk), .A(\g.we_clk [18926]));
Q_ASSIGN U13849 ( .B(clk), .A(\g.we_clk [18925]));
Q_ASSIGN U13850 ( .B(clk), .A(\g.we_clk [18924]));
Q_ASSIGN U13851 ( .B(clk), .A(\g.we_clk [18923]));
Q_ASSIGN U13852 ( .B(clk), .A(\g.we_clk [18922]));
Q_ASSIGN U13853 ( .B(clk), .A(\g.we_clk [18921]));
Q_ASSIGN U13854 ( .B(clk), .A(\g.we_clk [18920]));
Q_ASSIGN U13855 ( .B(clk), .A(\g.we_clk [18919]));
Q_ASSIGN U13856 ( .B(clk), .A(\g.we_clk [18918]));
Q_ASSIGN U13857 ( .B(clk), .A(\g.we_clk [18917]));
Q_ASSIGN U13858 ( .B(clk), .A(\g.we_clk [18916]));
Q_ASSIGN U13859 ( .B(clk), .A(\g.we_clk [18915]));
Q_ASSIGN U13860 ( .B(clk), .A(\g.we_clk [18914]));
Q_ASSIGN U13861 ( .B(clk), .A(\g.we_clk [18913]));
Q_ASSIGN U13862 ( .B(clk), .A(\g.we_clk [18912]));
Q_ASSIGN U13863 ( .B(clk), .A(\g.we_clk [18911]));
Q_ASSIGN U13864 ( .B(clk), .A(\g.we_clk [18910]));
Q_ASSIGN U13865 ( .B(clk), .A(\g.we_clk [18909]));
Q_ASSIGN U13866 ( .B(clk), .A(\g.we_clk [18908]));
Q_ASSIGN U13867 ( .B(clk), .A(\g.we_clk [18907]));
Q_ASSIGN U13868 ( .B(clk), .A(\g.we_clk [18906]));
Q_ASSIGN U13869 ( .B(clk), .A(\g.we_clk [18905]));
Q_ASSIGN U13870 ( .B(clk), .A(\g.we_clk [18904]));
Q_ASSIGN U13871 ( .B(clk), .A(\g.we_clk [18903]));
Q_ASSIGN U13872 ( .B(clk), .A(\g.we_clk [18902]));
Q_ASSIGN U13873 ( .B(clk), .A(\g.we_clk [18901]));
Q_ASSIGN U13874 ( .B(clk), .A(\g.we_clk [18900]));
Q_ASSIGN U13875 ( .B(clk), .A(\g.we_clk [18899]));
Q_ASSIGN U13876 ( .B(clk), .A(\g.we_clk [18898]));
Q_ASSIGN U13877 ( .B(clk), .A(\g.we_clk [18897]));
Q_ASSIGN U13878 ( .B(clk), .A(\g.we_clk [18896]));
Q_ASSIGN U13879 ( .B(clk), .A(\g.we_clk [18895]));
Q_ASSIGN U13880 ( .B(clk), .A(\g.we_clk [18894]));
Q_ASSIGN U13881 ( .B(clk), .A(\g.we_clk [18893]));
Q_ASSIGN U13882 ( .B(clk), .A(\g.we_clk [18892]));
Q_ASSIGN U13883 ( .B(clk), .A(\g.we_clk [18891]));
Q_ASSIGN U13884 ( .B(clk), .A(\g.we_clk [18890]));
Q_ASSIGN U13885 ( .B(clk), .A(\g.we_clk [18889]));
Q_ASSIGN U13886 ( .B(clk), .A(\g.we_clk [18888]));
Q_ASSIGN U13887 ( .B(clk), .A(\g.we_clk [18887]));
Q_ASSIGN U13888 ( .B(clk), .A(\g.we_clk [18886]));
Q_ASSIGN U13889 ( .B(clk), .A(\g.we_clk [18885]));
Q_ASSIGN U13890 ( .B(clk), .A(\g.we_clk [18884]));
Q_ASSIGN U13891 ( .B(clk), .A(\g.we_clk [18883]));
Q_ASSIGN U13892 ( .B(clk), .A(\g.we_clk [18882]));
Q_ASSIGN U13893 ( .B(clk), .A(\g.we_clk [18881]));
Q_ASSIGN U13894 ( .B(clk), .A(\g.we_clk [18880]));
Q_ASSIGN U13895 ( .B(clk), .A(\g.we_clk [18879]));
Q_ASSIGN U13896 ( .B(clk), .A(\g.we_clk [18878]));
Q_ASSIGN U13897 ( .B(clk), .A(\g.we_clk [18877]));
Q_ASSIGN U13898 ( .B(clk), .A(\g.we_clk [18876]));
Q_ASSIGN U13899 ( .B(clk), .A(\g.we_clk [18875]));
Q_ASSIGN U13900 ( .B(clk), .A(\g.we_clk [18874]));
Q_ASSIGN U13901 ( .B(clk), .A(\g.we_clk [18873]));
Q_ASSIGN U13902 ( .B(clk), .A(\g.we_clk [18872]));
Q_ASSIGN U13903 ( .B(clk), .A(\g.we_clk [18871]));
Q_ASSIGN U13904 ( .B(clk), .A(\g.we_clk [18870]));
Q_ASSIGN U13905 ( .B(clk), .A(\g.we_clk [18869]));
Q_ASSIGN U13906 ( .B(clk), .A(\g.we_clk [18868]));
Q_ASSIGN U13907 ( .B(clk), .A(\g.we_clk [18867]));
Q_ASSIGN U13908 ( .B(clk), .A(\g.we_clk [18866]));
Q_ASSIGN U13909 ( .B(clk), .A(\g.we_clk [18865]));
Q_ASSIGN U13910 ( .B(clk), .A(\g.we_clk [18864]));
Q_ASSIGN U13911 ( .B(clk), .A(\g.we_clk [18863]));
Q_ASSIGN U13912 ( .B(clk), .A(\g.we_clk [18862]));
Q_ASSIGN U13913 ( .B(clk), .A(\g.we_clk [18861]));
Q_ASSIGN U13914 ( .B(clk), .A(\g.we_clk [18860]));
Q_ASSIGN U13915 ( .B(clk), .A(\g.we_clk [18859]));
Q_ASSIGN U13916 ( .B(clk), .A(\g.we_clk [18858]));
Q_ASSIGN U13917 ( .B(clk), .A(\g.we_clk [18857]));
Q_ASSIGN U13918 ( .B(clk), .A(\g.we_clk [18856]));
Q_ASSIGN U13919 ( .B(clk), .A(\g.we_clk [18855]));
Q_ASSIGN U13920 ( .B(clk), .A(\g.we_clk [18854]));
Q_ASSIGN U13921 ( .B(clk), .A(\g.we_clk [18853]));
Q_ASSIGN U13922 ( .B(clk), .A(\g.we_clk [18852]));
Q_ASSIGN U13923 ( .B(clk), .A(\g.we_clk [18851]));
Q_ASSIGN U13924 ( .B(clk), .A(\g.we_clk [18850]));
Q_ASSIGN U13925 ( .B(clk), .A(\g.we_clk [18849]));
Q_ASSIGN U13926 ( .B(clk), .A(\g.we_clk [18848]));
Q_ASSIGN U13927 ( .B(clk), .A(\g.we_clk [18847]));
Q_ASSIGN U13928 ( .B(clk), .A(\g.we_clk [18846]));
Q_ASSIGN U13929 ( .B(clk), .A(\g.we_clk [18845]));
Q_ASSIGN U13930 ( .B(clk), .A(\g.we_clk [18844]));
Q_ASSIGN U13931 ( .B(clk), .A(\g.we_clk [18843]));
Q_ASSIGN U13932 ( .B(clk), .A(\g.we_clk [18842]));
Q_ASSIGN U13933 ( .B(clk), .A(\g.we_clk [18841]));
Q_ASSIGN U13934 ( .B(clk), .A(\g.we_clk [18840]));
Q_ASSIGN U13935 ( .B(clk), .A(\g.we_clk [18839]));
Q_ASSIGN U13936 ( .B(clk), .A(\g.we_clk [18838]));
Q_ASSIGN U13937 ( .B(clk), .A(\g.we_clk [18837]));
Q_ASSIGN U13938 ( .B(clk), .A(\g.we_clk [18836]));
Q_ASSIGN U13939 ( .B(clk), .A(\g.we_clk [18835]));
Q_ASSIGN U13940 ( .B(clk), .A(\g.we_clk [18834]));
Q_ASSIGN U13941 ( .B(clk), .A(\g.we_clk [18833]));
Q_ASSIGN U13942 ( .B(clk), .A(\g.we_clk [18832]));
Q_ASSIGN U13943 ( .B(clk), .A(\g.we_clk [18831]));
Q_ASSIGN U13944 ( .B(clk), .A(\g.we_clk [18830]));
Q_ASSIGN U13945 ( .B(clk), .A(\g.we_clk [18829]));
Q_ASSIGN U13946 ( .B(clk), .A(\g.we_clk [18828]));
Q_ASSIGN U13947 ( .B(clk), .A(\g.we_clk [18827]));
Q_ASSIGN U13948 ( .B(clk), .A(\g.we_clk [18826]));
Q_ASSIGN U13949 ( .B(clk), .A(\g.we_clk [18825]));
Q_ASSIGN U13950 ( .B(clk), .A(\g.we_clk [18824]));
Q_ASSIGN U13951 ( .B(clk), .A(\g.we_clk [18823]));
Q_ASSIGN U13952 ( .B(clk), .A(\g.we_clk [18822]));
Q_ASSIGN U13953 ( .B(clk), .A(\g.we_clk [18821]));
Q_ASSIGN U13954 ( .B(clk), .A(\g.we_clk [18820]));
Q_ASSIGN U13955 ( .B(clk), .A(\g.we_clk [18819]));
Q_ASSIGN U13956 ( .B(clk), .A(\g.we_clk [18818]));
Q_ASSIGN U13957 ( .B(clk), .A(\g.we_clk [18817]));
Q_ASSIGN U13958 ( .B(clk), .A(\g.we_clk [18816]));
Q_ASSIGN U13959 ( .B(clk), .A(\g.we_clk [18815]));
Q_ASSIGN U13960 ( .B(clk), .A(\g.we_clk [18814]));
Q_ASSIGN U13961 ( .B(clk), .A(\g.we_clk [18813]));
Q_ASSIGN U13962 ( .B(clk), .A(\g.we_clk [18812]));
Q_ASSIGN U13963 ( .B(clk), .A(\g.we_clk [18811]));
Q_ASSIGN U13964 ( .B(clk), .A(\g.we_clk [18810]));
Q_ASSIGN U13965 ( .B(clk), .A(\g.we_clk [18809]));
Q_ASSIGN U13966 ( .B(clk), .A(\g.we_clk [18808]));
Q_ASSIGN U13967 ( .B(clk), .A(\g.we_clk [18807]));
Q_ASSIGN U13968 ( .B(clk), .A(\g.we_clk [18806]));
Q_ASSIGN U13969 ( .B(clk), .A(\g.we_clk [18805]));
Q_ASSIGN U13970 ( .B(clk), .A(\g.we_clk [18804]));
Q_ASSIGN U13971 ( .B(clk), .A(\g.we_clk [18803]));
Q_ASSIGN U13972 ( .B(clk), .A(\g.we_clk [18802]));
Q_ASSIGN U13973 ( .B(clk), .A(\g.we_clk [18801]));
Q_ASSIGN U13974 ( .B(clk), .A(\g.we_clk [18800]));
Q_ASSIGN U13975 ( .B(clk), .A(\g.we_clk [18799]));
Q_ASSIGN U13976 ( .B(clk), .A(\g.we_clk [18798]));
Q_ASSIGN U13977 ( .B(clk), .A(\g.we_clk [18797]));
Q_ASSIGN U13978 ( .B(clk), .A(\g.we_clk [18796]));
Q_ASSIGN U13979 ( .B(clk), .A(\g.we_clk [18795]));
Q_ASSIGN U13980 ( .B(clk), .A(\g.we_clk [18794]));
Q_ASSIGN U13981 ( .B(clk), .A(\g.we_clk [18793]));
Q_ASSIGN U13982 ( .B(clk), .A(\g.we_clk [18792]));
Q_ASSIGN U13983 ( .B(clk), .A(\g.we_clk [18791]));
Q_ASSIGN U13984 ( .B(clk), .A(\g.we_clk [18790]));
Q_ASSIGN U13985 ( .B(clk), .A(\g.we_clk [18789]));
Q_ASSIGN U13986 ( .B(clk), .A(\g.we_clk [18788]));
Q_ASSIGN U13987 ( .B(clk), .A(\g.we_clk [18787]));
Q_ASSIGN U13988 ( .B(clk), .A(\g.we_clk [18786]));
Q_ASSIGN U13989 ( .B(clk), .A(\g.we_clk [18785]));
Q_ASSIGN U13990 ( .B(clk), .A(\g.we_clk [18784]));
Q_ASSIGN U13991 ( .B(clk), .A(\g.we_clk [18783]));
Q_ASSIGN U13992 ( .B(clk), .A(\g.we_clk [18782]));
Q_ASSIGN U13993 ( .B(clk), .A(\g.we_clk [18781]));
Q_ASSIGN U13994 ( .B(clk), .A(\g.we_clk [18780]));
Q_ASSIGN U13995 ( .B(clk), .A(\g.we_clk [18779]));
Q_ASSIGN U13996 ( .B(clk), .A(\g.we_clk [18778]));
Q_ASSIGN U13997 ( .B(clk), .A(\g.we_clk [18777]));
Q_ASSIGN U13998 ( .B(clk), .A(\g.we_clk [18776]));
Q_ASSIGN U13999 ( .B(clk), .A(\g.we_clk [18775]));
Q_ASSIGN U14000 ( .B(clk), .A(\g.we_clk [18774]));
Q_ASSIGN U14001 ( .B(clk), .A(\g.we_clk [18773]));
Q_ASSIGN U14002 ( .B(clk), .A(\g.we_clk [18772]));
Q_ASSIGN U14003 ( .B(clk), .A(\g.we_clk [18771]));
Q_ASSIGN U14004 ( .B(clk), .A(\g.we_clk [18770]));
Q_ASSIGN U14005 ( .B(clk), .A(\g.we_clk [18769]));
Q_ASSIGN U14006 ( .B(clk), .A(\g.we_clk [18768]));
Q_ASSIGN U14007 ( .B(clk), .A(\g.we_clk [18767]));
Q_ASSIGN U14008 ( .B(clk), .A(\g.we_clk [18766]));
Q_ASSIGN U14009 ( .B(clk), .A(\g.we_clk [18765]));
Q_ASSIGN U14010 ( .B(clk), .A(\g.we_clk [18764]));
Q_ASSIGN U14011 ( .B(clk), .A(\g.we_clk [18763]));
Q_ASSIGN U14012 ( .B(clk), .A(\g.we_clk [18762]));
Q_ASSIGN U14013 ( .B(clk), .A(\g.we_clk [18761]));
Q_ASSIGN U14014 ( .B(clk), .A(\g.we_clk [18760]));
Q_ASSIGN U14015 ( .B(clk), .A(\g.we_clk [18759]));
Q_ASSIGN U14016 ( .B(clk), .A(\g.we_clk [18758]));
Q_ASSIGN U14017 ( .B(clk), .A(\g.we_clk [18757]));
Q_ASSIGN U14018 ( .B(clk), .A(\g.we_clk [18756]));
Q_ASSIGN U14019 ( .B(clk), .A(\g.we_clk [18755]));
Q_ASSIGN U14020 ( .B(clk), .A(\g.we_clk [18754]));
Q_ASSIGN U14021 ( .B(clk), .A(\g.we_clk [18753]));
Q_ASSIGN U14022 ( .B(clk), .A(\g.we_clk [18752]));
Q_ASSIGN U14023 ( .B(clk), .A(\g.we_clk [18751]));
Q_ASSIGN U14024 ( .B(clk), .A(\g.we_clk [18750]));
Q_ASSIGN U14025 ( .B(clk), .A(\g.we_clk [18749]));
Q_ASSIGN U14026 ( .B(clk), .A(\g.we_clk [18748]));
Q_ASSIGN U14027 ( .B(clk), .A(\g.we_clk [18747]));
Q_ASSIGN U14028 ( .B(clk), .A(\g.we_clk [18746]));
Q_ASSIGN U14029 ( .B(clk), .A(\g.we_clk [18745]));
Q_ASSIGN U14030 ( .B(clk), .A(\g.we_clk [18744]));
Q_ASSIGN U14031 ( .B(clk), .A(\g.we_clk [18743]));
Q_ASSIGN U14032 ( .B(clk), .A(\g.we_clk [18742]));
Q_ASSIGN U14033 ( .B(clk), .A(\g.we_clk [18741]));
Q_ASSIGN U14034 ( .B(clk), .A(\g.we_clk [18740]));
Q_ASSIGN U14035 ( .B(clk), .A(\g.we_clk [18739]));
Q_ASSIGN U14036 ( .B(clk), .A(\g.we_clk [18738]));
Q_ASSIGN U14037 ( .B(clk), .A(\g.we_clk [18737]));
Q_ASSIGN U14038 ( .B(clk), .A(\g.we_clk [18736]));
Q_ASSIGN U14039 ( .B(clk), .A(\g.we_clk [18735]));
Q_ASSIGN U14040 ( .B(clk), .A(\g.we_clk [18734]));
Q_ASSIGN U14041 ( .B(clk), .A(\g.we_clk [18733]));
Q_ASSIGN U14042 ( .B(clk), .A(\g.we_clk [18732]));
Q_ASSIGN U14043 ( .B(clk), .A(\g.we_clk [18731]));
Q_ASSIGN U14044 ( .B(clk), .A(\g.we_clk [18730]));
Q_ASSIGN U14045 ( .B(clk), .A(\g.we_clk [18729]));
Q_ASSIGN U14046 ( .B(clk), .A(\g.we_clk [18728]));
Q_ASSIGN U14047 ( .B(clk), .A(\g.we_clk [18727]));
Q_ASSIGN U14048 ( .B(clk), .A(\g.we_clk [18726]));
Q_ASSIGN U14049 ( .B(clk), .A(\g.we_clk [18725]));
Q_ASSIGN U14050 ( .B(clk), .A(\g.we_clk [18724]));
Q_ASSIGN U14051 ( .B(clk), .A(\g.we_clk [18723]));
Q_ASSIGN U14052 ( .B(clk), .A(\g.we_clk [18722]));
Q_ASSIGN U14053 ( .B(clk), .A(\g.we_clk [18721]));
Q_ASSIGN U14054 ( .B(clk), .A(\g.we_clk [18720]));
Q_ASSIGN U14055 ( .B(clk), .A(\g.we_clk [18719]));
Q_ASSIGN U14056 ( .B(clk), .A(\g.we_clk [18718]));
Q_ASSIGN U14057 ( .B(clk), .A(\g.we_clk [18717]));
Q_ASSIGN U14058 ( .B(clk), .A(\g.we_clk [18716]));
Q_ASSIGN U14059 ( .B(clk), .A(\g.we_clk [18715]));
Q_ASSIGN U14060 ( .B(clk), .A(\g.we_clk [18714]));
Q_ASSIGN U14061 ( .B(clk), .A(\g.we_clk [18713]));
Q_ASSIGN U14062 ( .B(clk), .A(\g.we_clk [18712]));
Q_ASSIGN U14063 ( .B(clk), .A(\g.we_clk [18711]));
Q_ASSIGN U14064 ( .B(clk), .A(\g.we_clk [18710]));
Q_ASSIGN U14065 ( .B(clk), .A(\g.we_clk [18709]));
Q_ASSIGN U14066 ( .B(clk), .A(\g.we_clk [18708]));
Q_ASSIGN U14067 ( .B(clk), .A(\g.we_clk [18707]));
Q_ASSIGN U14068 ( .B(clk), .A(\g.we_clk [18706]));
Q_ASSIGN U14069 ( .B(clk), .A(\g.we_clk [18705]));
Q_ASSIGN U14070 ( .B(clk), .A(\g.we_clk [18704]));
Q_ASSIGN U14071 ( .B(clk), .A(\g.we_clk [18703]));
Q_ASSIGN U14072 ( .B(clk), .A(\g.we_clk [18702]));
Q_ASSIGN U14073 ( .B(clk), .A(\g.we_clk [18701]));
Q_ASSIGN U14074 ( .B(clk), .A(\g.we_clk [18700]));
Q_ASSIGN U14075 ( .B(clk), .A(\g.we_clk [18699]));
Q_ASSIGN U14076 ( .B(clk), .A(\g.we_clk [18698]));
Q_ASSIGN U14077 ( .B(clk), .A(\g.we_clk [18697]));
Q_ASSIGN U14078 ( .B(clk), .A(\g.we_clk [18696]));
Q_ASSIGN U14079 ( .B(clk), .A(\g.we_clk [18695]));
Q_ASSIGN U14080 ( .B(clk), .A(\g.we_clk [18694]));
Q_ASSIGN U14081 ( .B(clk), .A(\g.we_clk [18693]));
Q_ASSIGN U14082 ( .B(clk), .A(\g.we_clk [18692]));
Q_ASSIGN U14083 ( .B(clk), .A(\g.we_clk [18691]));
Q_ASSIGN U14084 ( .B(clk), .A(\g.we_clk [18690]));
Q_ASSIGN U14085 ( .B(clk), .A(\g.we_clk [18689]));
Q_ASSIGN U14086 ( .B(clk), .A(\g.we_clk [18688]));
Q_ASSIGN U14087 ( .B(clk), .A(\g.we_clk [18687]));
Q_ASSIGN U14088 ( .B(clk), .A(\g.we_clk [18686]));
Q_ASSIGN U14089 ( .B(clk), .A(\g.we_clk [18685]));
Q_ASSIGN U14090 ( .B(clk), .A(\g.we_clk [18684]));
Q_ASSIGN U14091 ( .B(clk), .A(\g.we_clk [18683]));
Q_ASSIGN U14092 ( .B(clk), .A(\g.we_clk [18682]));
Q_ASSIGN U14093 ( .B(clk), .A(\g.we_clk [18681]));
Q_ASSIGN U14094 ( .B(clk), .A(\g.we_clk [18680]));
Q_ASSIGN U14095 ( .B(clk), .A(\g.we_clk [18679]));
Q_ASSIGN U14096 ( .B(clk), .A(\g.we_clk [18678]));
Q_ASSIGN U14097 ( .B(clk), .A(\g.we_clk [18677]));
Q_ASSIGN U14098 ( .B(clk), .A(\g.we_clk [18676]));
Q_ASSIGN U14099 ( .B(clk), .A(\g.we_clk [18675]));
Q_ASSIGN U14100 ( .B(clk), .A(\g.we_clk [18674]));
Q_ASSIGN U14101 ( .B(clk), .A(\g.we_clk [18673]));
Q_ASSIGN U14102 ( .B(clk), .A(\g.we_clk [18672]));
Q_ASSIGN U14103 ( .B(clk), .A(\g.we_clk [18671]));
Q_ASSIGN U14104 ( .B(clk), .A(\g.we_clk [18670]));
Q_ASSIGN U14105 ( .B(clk), .A(\g.we_clk [18669]));
Q_ASSIGN U14106 ( .B(clk), .A(\g.we_clk [18668]));
Q_ASSIGN U14107 ( .B(clk), .A(\g.we_clk [18667]));
Q_ASSIGN U14108 ( .B(clk), .A(\g.we_clk [18666]));
Q_ASSIGN U14109 ( .B(clk), .A(\g.we_clk [18665]));
Q_ASSIGN U14110 ( .B(clk), .A(\g.we_clk [18664]));
Q_ASSIGN U14111 ( .B(clk), .A(\g.we_clk [18663]));
Q_ASSIGN U14112 ( .B(clk), .A(\g.we_clk [18662]));
Q_ASSIGN U14113 ( .B(clk), .A(\g.we_clk [18661]));
Q_ASSIGN U14114 ( .B(clk), .A(\g.we_clk [18660]));
Q_ASSIGN U14115 ( .B(clk), .A(\g.we_clk [18659]));
Q_ASSIGN U14116 ( .B(clk), .A(\g.we_clk [18658]));
Q_ASSIGN U14117 ( .B(clk), .A(\g.we_clk [18657]));
Q_ASSIGN U14118 ( .B(clk), .A(\g.we_clk [18656]));
Q_ASSIGN U14119 ( .B(clk), .A(\g.we_clk [18655]));
Q_ASSIGN U14120 ( .B(clk), .A(\g.we_clk [18654]));
Q_ASSIGN U14121 ( .B(clk), .A(\g.we_clk [18653]));
Q_ASSIGN U14122 ( .B(clk), .A(\g.we_clk [18652]));
Q_ASSIGN U14123 ( .B(clk), .A(\g.we_clk [18651]));
Q_ASSIGN U14124 ( .B(clk), .A(\g.we_clk [18650]));
Q_ASSIGN U14125 ( .B(clk), .A(\g.we_clk [18649]));
Q_ASSIGN U14126 ( .B(clk), .A(\g.we_clk [18648]));
Q_ASSIGN U14127 ( .B(clk), .A(\g.we_clk [18647]));
Q_ASSIGN U14128 ( .B(clk), .A(\g.we_clk [18646]));
Q_ASSIGN U14129 ( .B(clk), .A(\g.we_clk [18645]));
Q_ASSIGN U14130 ( .B(clk), .A(\g.we_clk [18644]));
Q_ASSIGN U14131 ( .B(clk), .A(\g.we_clk [18643]));
Q_ASSIGN U14132 ( .B(clk), .A(\g.we_clk [18642]));
Q_ASSIGN U14133 ( .B(clk), .A(\g.we_clk [18641]));
Q_ASSIGN U14134 ( .B(clk), .A(\g.we_clk [18640]));
Q_ASSIGN U14135 ( .B(clk), .A(\g.we_clk [18639]));
Q_ASSIGN U14136 ( .B(clk), .A(\g.we_clk [18638]));
Q_ASSIGN U14137 ( .B(clk), .A(\g.we_clk [18637]));
Q_ASSIGN U14138 ( .B(clk), .A(\g.we_clk [18636]));
Q_ASSIGN U14139 ( .B(clk), .A(\g.we_clk [18635]));
Q_ASSIGN U14140 ( .B(clk), .A(\g.we_clk [18634]));
Q_ASSIGN U14141 ( .B(clk), .A(\g.we_clk [18633]));
Q_ASSIGN U14142 ( .B(clk), .A(\g.we_clk [18632]));
Q_ASSIGN U14143 ( .B(clk), .A(\g.we_clk [18631]));
Q_ASSIGN U14144 ( .B(clk), .A(\g.we_clk [18630]));
Q_ASSIGN U14145 ( .B(clk), .A(\g.we_clk [18629]));
Q_ASSIGN U14146 ( .B(clk), .A(\g.we_clk [18628]));
Q_ASSIGN U14147 ( .B(clk), .A(\g.we_clk [18627]));
Q_ASSIGN U14148 ( .B(clk), .A(\g.we_clk [18626]));
Q_ASSIGN U14149 ( .B(clk), .A(\g.we_clk [18625]));
Q_ASSIGN U14150 ( .B(clk), .A(\g.we_clk [18624]));
Q_ASSIGN U14151 ( .B(clk), .A(\g.we_clk [18623]));
Q_ASSIGN U14152 ( .B(clk), .A(\g.we_clk [18622]));
Q_ASSIGN U14153 ( .B(clk), .A(\g.we_clk [18621]));
Q_ASSIGN U14154 ( .B(clk), .A(\g.we_clk [18620]));
Q_ASSIGN U14155 ( .B(clk), .A(\g.we_clk [18619]));
Q_ASSIGN U14156 ( .B(clk), .A(\g.we_clk [18618]));
Q_ASSIGN U14157 ( .B(clk), .A(\g.we_clk [18617]));
Q_ASSIGN U14158 ( .B(clk), .A(\g.we_clk [18616]));
Q_ASSIGN U14159 ( .B(clk), .A(\g.we_clk [18615]));
Q_ASSIGN U14160 ( .B(clk), .A(\g.we_clk [18614]));
Q_ASSIGN U14161 ( .B(clk), .A(\g.we_clk [18613]));
Q_ASSIGN U14162 ( .B(clk), .A(\g.we_clk [18612]));
Q_ASSIGN U14163 ( .B(clk), .A(\g.we_clk [18611]));
Q_ASSIGN U14164 ( .B(clk), .A(\g.we_clk [18610]));
Q_ASSIGN U14165 ( .B(clk), .A(\g.we_clk [18609]));
Q_ASSIGN U14166 ( .B(clk), .A(\g.we_clk [18608]));
Q_ASSIGN U14167 ( .B(clk), .A(\g.we_clk [18607]));
Q_ASSIGN U14168 ( .B(clk), .A(\g.we_clk [18606]));
Q_ASSIGN U14169 ( .B(clk), .A(\g.we_clk [18605]));
Q_ASSIGN U14170 ( .B(clk), .A(\g.we_clk [18604]));
Q_ASSIGN U14171 ( .B(clk), .A(\g.we_clk [18603]));
Q_ASSIGN U14172 ( .B(clk), .A(\g.we_clk [18602]));
Q_ASSIGN U14173 ( .B(clk), .A(\g.we_clk [18601]));
Q_ASSIGN U14174 ( .B(clk), .A(\g.we_clk [18600]));
Q_ASSIGN U14175 ( .B(clk), .A(\g.we_clk [18599]));
Q_ASSIGN U14176 ( .B(clk), .A(\g.we_clk [18598]));
Q_ASSIGN U14177 ( .B(clk), .A(\g.we_clk [18597]));
Q_ASSIGN U14178 ( .B(clk), .A(\g.we_clk [18596]));
Q_ASSIGN U14179 ( .B(clk), .A(\g.we_clk [18595]));
Q_ASSIGN U14180 ( .B(clk), .A(\g.we_clk [18594]));
Q_ASSIGN U14181 ( .B(clk), .A(\g.we_clk [18593]));
Q_ASSIGN U14182 ( .B(clk), .A(\g.we_clk [18592]));
Q_ASSIGN U14183 ( .B(clk), .A(\g.we_clk [18591]));
Q_ASSIGN U14184 ( .B(clk), .A(\g.we_clk [18590]));
Q_ASSIGN U14185 ( .B(clk), .A(\g.we_clk [18589]));
Q_ASSIGN U14186 ( .B(clk), .A(\g.we_clk [18588]));
Q_ASSIGN U14187 ( .B(clk), .A(\g.we_clk [18587]));
Q_ASSIGN U14188 ( .B(clk), .A(\g.we_clk [18586]));
Q_ASSIGN U14189 ( .B(clk), .A(\g.we_clk [18585]));
Q_ASSIGN U14190 ( .B(clk), .A(\g.we_clk [18584]));
Q_ASSIGN U14191 ( .B(clk), .A(\g.we_clk [18583]));
Q_ASSIGN U14192 ( .B(clk), .A(\g.we_clk [18582]));
Q_ASSIGN U14193 ( .B(clk), .A(\g.we_clk [18581]));
Q_ASSIGN U14194 ( .B(clk), .A(\g.we_clk [18580]));
Q_ASSIGN U14195 ( .B(clk), .A(\g.we_clk [18579]));
Q_ASSIGN U14196 ( .B(clk), .A(\g.we_clk [18578]));
Q_ASSIGN U14197 ( .B(clk), .A(\g.we_clk [18577]));
Q_ASSIGN U14198 ( .B(clk), .A(\g.we_clk [18576]));
Q_ASSIGN U14199 ( .B(clk), .A(\g.we_clk [18575]));
Q_ASSIGN U14200 ( .B(clk), .A(\g.we_clk [18574]));
Q_ASSIGN U14201 ( .B(clk), .A(\g.we_clk [18573]));
Q_ASSIGN U14202 ( .B(clk), .A(\g.we_clk [18572]));
Q_ASSIGN U14203 ( .B(clk), .A(\g.we_clk [18571]));
Q_ASSIGN U14204 ( .B(clk), .A(\g.we_clk [18570]));
Q_ASSIGN U14205 ( .B(clk), .A(\g.we_clk [18569]));
Q_ASSIGN U14206 ( .B(clk), .A(\g.we_clk [18568]));
Q_ASSIGN U14207 ( .B(clk), .A(\g.we_clk [18567]));
Q_ASSIGN U14208 ( .B(clk), .A(\g.we_clk [18566]));
Q_ASSIGN U14209 ( .B(clk), .A(\g.we_clk [18565]));
Q_ASSIGN U14210 ( .B(clk), .A(\g.we_clk [18564]));
Q_ASSIGN U14211 ( .B(clk), .A(\g.we_clk [18563]));
Q_ASSIGN U14212 ( .B(clk), .A(\g.we_clk [18562]));
Q_ASSIGN U14213 ( .B(clk), .A(\g.we_clk [18561]));
Q_ASSIGN U14214 ( .B(clk), .A(\g.we_clk [18560]));
Q_ASSIGN U14215 ( .B(clk), .A(\g.we_clk [18559]));
Q_ASSIGN U14216 ( .B(clk), .A(\g.we_clk [18558]));
Q_ASSIGN U14217 ( .B(clk), .A(\g.we_clk [18557]));
Q_ASSIGN U14218 ( .B(clk), .A(\g.we_clk [18556]));
Q_ASSIGN U14219 ( .B(clk), .A(\g.we_clk [18555]));
Q_ASSIGN U14220 ( .B(clk), .A(\g.we_clk [18554]));
Q_ASSIGN U14221 ( .B(clk), .A(\g.we_clk [18553]));
Q_ASSIGN U14222 ( .B(clk), .A(\g.we_clk [18552]));
Q_ASSIGN U14223 ( .B(clk), .A(\g.we_clk [18551]));
Q_ASSIGN U14224 ( .B(clk), .A(\g.we_clk [18550]));
Q_ASSIGN U14225 ( .B(clk), .A(\g.we_clk [18549]));
Q_ASSIGN U14226 ( .B(clk), .A(\g.we_clk [18548]));
Q_ASSIGN U14227 ( .B(clk), .A(\g.we_clk [18547]));
Q_ASSIGN U14228 ( .B(clk), .A(\g.we_clk [18546]));
Q_ASSIGN U14229 ( .B(clk), .A(\g.we_clk [18545]));
Q_ASSIGN U14230 ( .B(clk), .A(\g.we_clk [18544]));
Q_ASSIGN U14231 ( .B(clk), .A(\g.we_clk [18543]));
Q_ASSIGN U14232 ( .B(clk), .A(\g.we_clk [18542]));
Q_ASSIGN U14233 ( .B(clk), .A(\g.we_clk [18541]));
Q_ASSIGN U14234 ( .B(clk), .A(\g.we_clk [18540]));
Q_ASSIGN U14235 ( .B(clk), .A(\g.we_clk [18539]));
Q_ASSIGN U14236 ( .B(clk), .A(\g.we_clk [18538]));
Q_ASSIGN U14237 ( .B(clk), .A(\g.we_clk [18537]));
Q_ASSIGN U14238 ( .B(clk), .A(\g.we_clk [18536]));
Q_ASSIGN U14239 ( .B(clk), .A(\g.we_clk [18535]));
Q_ASSIGN U14240 ( .B(clk), .A(\g.we_clk [18534]));
Q_ASSIGN U14241 ( .B(clk), .A(\g.we_clk [18533]));
Q_ASSIGN U14242 ( .B(clk), .A(\g.we_clk [18532]));
Q_ASSIGN U14243 ( .B(clk), .A(\g.we_clk [18531]));
Q_ASSIGN U14244 ( .B(clk), .A(\g.we_clk [18530]));
Q_ASSIGN U14245 ( .B(clk), .A(\g.we_clk [18529]));
Q_ASSIGN U14246 ( .B(clk), .A(\g.we_clk [18528]));
Q_ASSIGN U14247 ( .B(clk), .A(\g.we_clk [18527]));
Q_ASSIGN U14248 ( .B(clk), .A(\g.we_clk [18526]));
Q_ASSIGN U14249 ( .B(clk), .A(\g.we_clk [18525]));
Q_ASSIGN U14250 ( .B(clk), .A(\g.we_clk [18524]));
Q_ASSIGN U14251 ( .B(clk), .A(\g.we_clk [18523]));
Q_ASSIGN U14252 ( .B(clk), .A(\g.we_clk [18522]));
Q_ASSIGN U14253 ( .B(clk), .A(\g.we_clk [18521]));
Q_ASSIGN U14254 ( .B(clk), .A(\g.we_clk [18520]));
Q_ASSIGN U14255 ( .B(clk), .A(\g.we_clk [18519]));
Q_ASSIGN U14256 ( .B(clk), .A(\g.we_clk [18518]));
Q_ASSIGN U14257 ( .B(clk), .A(\g.we_clk [18517]));
Q_ASSIGN U14258 ( .B(clk), .A(\g.we_clk [18516]));
Q_ASSIGN U14259 ( .B(clk), .A(\g.we_clk [18515]));
Q_ASSIGN U14260 ( .B(clk), .A(\g.we_clk [18514]));
Q_ASSIGN U14261 ( .B(clk), .A(\g.we_clk [18513]));
Q_ASSIGN U14262 ( .B(clk), .A(\g.we_clk [18512]));
Q_ASSIGN U14263 ( .B(clk), .A(\g.we_clk [18511]));
Q_ASSIGN U14264 ( .B(clk), .A(\g.we_clk [18510]));
Q_ASSIGN U14265 ( .B(clk), .A(\g.we_clk [18509]));
Q_ASSIGN U14266 ( .B(clk), .A(\g.we_clk [18508]));
Q_ASSIGN U14267 ( .B(clk), .A(\g.we_clk [18507]));
Q_ASSIGN U14268 ( .B(clk), .A(\g.we_clk [18506]));
Q_ASSIGN U14269 ( .B(clk), .A(\g.we_clk [18505]));
Q_ASSIGN U14270 ( .B(clk), .A(\g.we_clk [18504]));
Q_ASSIGN U14271 ( .B(clk), .A(\g.we_clk [18503]));
Q_ASSIGN U14272 ( .B(clk), .A(\g.we_clk [18502]));
Q_ASSIGN U14273 ( .B(clk), .A(\g.we_clk [18501]));
Q_ASSIGN U14274 ( .B(clk), .A(\g.we_clk [18500]));
Q_ASSIGN U14275 ( .B(clk), .A(\g.we_clk [18499]));
Q_ASSIGN U14276 ( .B(clk), .A(\g.we_clk [18498]));
Q_ASSIGN U14277 ( .B(clk), .A(\g.we_clk [18497]));
Q_ASSIGN U14278 ( .B(clk), .A(\g.we_clk [18496]));
Q_ASSIGN U14279 ( .B(clk), .A(\g.we_clk [18495]));
Q_ASSIGN U14280 ( .B(clk), .A(\g.we_clk [18494]));
Q_ASSIGN U14281 ( .B(clk), .A(\g.we_clk [18493]));
Q_ASSIGN U14282 ( .B(clk), .A(\g.we_clk [18492]));
Q_ASSIGN U14283 ( .B(clk), .A(\g.we_clk [18491]));
Q_ASSIGN U14284 ( .B(clk), .A(\g.we_clk [18490]));
Q_ASSIGN U14285 ( .B(clk), .A(\g.we_clk [18489]));
Q_ASSIGN U14286 ( .B(clk), .A(\g.we_clk [18488]));
Q_ASSIGN U14287 ( .B(clk), .A(\g.we_clk [18487]));
Q_ASSIGN U14288 ( .B(clk), .A(\g.we_clk [18486]));
Q_ASSIGN U14289 ( .B(clk), .A(\g.we_clk [18485]));
Q_ASSIGN U14290 ( .B(clk), .A(\g.we_clk [18484]));
Q_ASSIGN U14291 ( .B(clk), .A(\g.we_clk [18483]));
Q_ASSIGN U14292 ( .B(clk), .A(\g.we_clk [18482]));
Q_ASSIGN U14293 ( .B(clk), .A(\g.we_clk [18481]));
Q_ASSIGN U14294 ( .B(clk), .A(\g.we_clk [18480]));
Q_ASSIGN U14295 ( .B(clk), .A(\g.we_clk [18479]));
Q_ASSIGN U14296 ( .B(clk), .A(\g.we_clk [18478]));
Q_ASSIGN U14297 ( .B(clk), .A(\g.we_clk [18477]));
Q_ASSIGN U14298 ( .B(clk), .A(\g.we_clk [18476]));
Q_ASSIGN U14299 ( .B(clk), .A(\g.we_clk [18475]));
Q_ASSIGN U14300 ( .B(clk), .A(\g.we_clk [18474]));
Q_ASSIGN U14301 ( .B(clk), .A(\g.we_clk [18473]));
Q_ASSIGN U14302 ( .B(clk), .A(\g.we_clk [18472]));
Q_ASSIGN U14303 ( .B(clk), .A(\g.we_clk [18471]));
Q_ASSIGN U14304 ( .B(clk), .A(\g.we_clk [18470]));
Q_ASSIGN U14305 ( .B(clk), .A(\g.we_clk [18469]));
Q_ASSIGN U14306 ( .B(clk), .A(\g.we_clk [18468]));
Q_ASSIGN U14307 ( .B(clk), .A(\g.we_clk [18467]));
Q_ASSIGN U14308 ( .B(clk), .A(\g.we_clk [18466]));
Q_ASSIGN U14309 ( .B(clk), .A(\g.we_clk [18465]));
Q_ASSIGN U14310 ( .B(clk), .A(\g.we_clk [18464]));
Q_ASSIGN U14311 ( .B(clk), .A(\g.we_clk [18463]));
Q_ASSIGN U14312 ( .B(clk), .A(\g.we_clk [18462]));
Q_ASSIGN U14313 ( .B(clk), .A(\g.we_clk [18461]));
Q_ASSIGN U14314 ( .B(clk), .A(\g.we_clk [18460]));
Q_ASSIGN U14315 ( .B(clk), .A(\g.we_clk [18459]));
Q_ASSIGN U14316 ( .B(clk), .A(\g.we_clk [18458]));
Q_ASSIGN U14317 ( .B(clk), .A(\g.we_clk [18457]));
Q_ASSIGN U14318 ( .B(clk), .A(\g.we_clk [18456]));
Q_ASSIGN U14319 ( .B(clk), .A(\g.we_clk [18455]));
Q_ASSIGN U14320 ( .B(clk), .A(\g.we_clk [18454]));
Q_ASSIGN U14321 ( .B(clk), .A(\g.we_clk [18453]));
Q_ASSIGN U14322 ( .B(clk), .A(\g.we_clk [18452]));
Q_ASSIGN U14323 ( .B(clk), .A(\g.we_clk [18451]));
Q_ASSIGN U14324 ( .B(clk), .A(\g.we_clk [18450]));
Q_ASSIGN U14325 ( .B(clk), .A(\g.we_clk [18449]));
Q_ASSIGN U14326 ( .B(clk), .A(\g.we_clk [18448]));
Q_ASSIGN U14327 ( .B(clk), .A(\g.we_clk [18447]));
Q_ASSIGN U14328 ( .B(clk), .A(\g.we_clk [18446]));
Q_ASSIGN U14329 ( .B(clk), .A(\g.we_clk [18445]));
Q_ASSIGN U14330 ( .B(clk), .A(\g.we_clk [18444]));
Q_ASSIGN U14331 ( .B(clk), .A(\g.we_clk [18443]));
Q_ASSIGN U14332 ( .B(clk), .A(\g.we_clk [18442]));
Q_ASSIGN U14333 ( .B(clk), .A(\g.we_clk [18441]));
Q_ASSIGN U14334 ( .B(clk), .A(\g.we_clk [18440]));
Q_ASSIGN U14335 ( .B(clk), .A(\g.we_clk [18439]));
Q_ASSIGN U14336 ( .B(clk), .A(\g.we_clk [18438]));
Q_ASSIGN U14337 ( .B(clk), .A(\g.we_clk [18437]));
Q_ASSIGN U14338 ( .B(clk), .A(\g.we_clk [18436]));
Q_ASSIGN U14339 ( .B(clk), .A(\g.we_clk [18435]));
Q_ASSIGN U14340 ( .B(clk), .A(\g.we_clk [18434]));
Q_ASSIGN U14341 ( .B(clk), .A(\g.we_clk [18433]));
Q_ASSIGN U14342 ( .B(clk), .A(\g.we_clk [18432]));
Q_ASSIGN U14343 ( .B(clk), .A(\g.we_clk [18431]));
Q_ASSIGN U14344 ( .B(clk), .A(\g.we_clk [18430]));
Q_ASSIGN U14345 ( .B(clk), .A(\g.we_clk [18429]));
Q_ASSIGN U14346 ( .B(clk), .A(\g.we_clk [18428]));
Q_ASSIGN U14347 ( .B(clk), .A(\g.we_clk [18427]));
Q_ASSIGN U14348 ( .B(clk), .A(\g.we_clk [18426]));
Q_ASSIGN U14349 ( .B(clk), .A(\g.we_clk [18425]));
Q_ASSIGN U14350 ( .B(clk), .A(\g.we_clk [18424]));
Q_ASSIGN U14351 ( .B(clk), .A(\g.we_clk [18423]));
Q_ASSIGN U14352 ( .B(clk), .A(\g.we_clk [18422]));
Q_ASSIGN U14353 ( .B(clk), .A(\g.we_clk [18421]));
Q_ASSIGN U14354 ( .B(clk), .A(\g.we_clk [18420]));
Q_ASSIGN U14355 ( .B(clk), .A(\g.we_clk [18419]));
Q_ASSIGN U14356 ( .B(clk), .A(\g.we_clk [18418]));
Q_ASSIGN U14357 ( .B(clk), .A(\g.we_clk [18417]));
Q_ASSIGN U14358 ( .B(clk), .A(\g.we_clk [18416]));
Q_ASSIGN U14359 ( .B(clk), .A(\g.we_clk [18415]));
Q_ASSIGN U14360 ( .B(clk), .A(\g.we_clk [18414]));
Q_ASSIGN U14361 ( .B(clk), .A(\g.we_clk [18413]));
Q_ASSIGN U14362 ( .B(clk), .A(\g.we_clk [18412]));
Q_ASSIGN U14363 ( .B(clk), .A(\g.we_clk [18411]));
Q_ASSIGN U14364 ( .B(clk), .A(\g.we_clk [18410]));
Q_ASSIGN U14365 ( .B(clk), .A(\g.we_clk [18409]));
Q_ASSIGN U14366 ( .B(clk), .A(\g.we_clk [18408]));
Q_ASSIGN U14367 ( .B(clk), .A(\g.we_clk [18407]));
Q_ASSIGN U14368 ( .B(clk), .A(\g.we_clk [18406]));
Q_ASSIGN U14369 ( .B(clk), .A(\g.we_clk [18405]));
Q_ASSIGN U14370 ( .B(clk), .A(\g.we_clk [18404]));
Q_ASSIGN U14371 ( .B(clk), .A(\g.we_clk [18403]));
Q_ASSIGN U14372 ( .B(clk), .A(\g.we_clk [18402]));
Q_ASSIGN U14373 ( .B(clk), .A(\g.we_clk [18401]));
Q_ASSIGN U14374 ( .B(clk), .A(\g.we_clk [18400]));
Q_ASSIGN U14375 ( .B(clk), .A(\g.we_clk [18399]));
Q_ASSIGN U14376 ( .B(clk), .A(\g.we_clk [18398]));
Q_ASSIGN U14377 ( .B(clk), .A(\g.we_clk [18397]));
Q_ASSIGN U14378 ( .B(clk), .A(\g.we_clk [18396]));
Q_ASSIGN U14379 ( .B(clk), .A(\g.we_clk [18395]));
Q_ASSIGN U14380 ( .B(clk), .A(\g.we_clk [18394]));
Q_ASSIGN U14381 ( .B(clk), .A(\g.we_clk [18393]));
Q_ASSIGN U14382 ( .B(clk), .A(\g.we_clk [18392]));
Q_ASSIGN U14383 ( .B(clk), .A(\g.we_clk [18391]));
Q_ASSIGN U14384 ( .B(clk), .A(\g.we_clk [18390]));
Q_ASSIGN U14385 ( .B(clk), .A(\g.we_clk [18389]));
Q_ASSIGN U14386 ( .B(clk), .A(\g.we_clk [18388]));
Q_ASSIGN U14387 ( .B(clk), .A(\g.we_clk [18387]));
Q_ASSIGN U14388 ( .B(clk), .A(\g.we_clk [18386]));
Q_ASSIGN U14389 ( .B(clk), .A(\g.we_clk [18385]));
Q_ASSIGN U14390 ( .B(clk), .A(\g.we_clk [18384]));
Q_ASSIGN U14391 ( .B(clk), .A(\g.we_clk [18383]));
Q_ASSIGN U14392 ( .B(clk), .A(\g.we_clk [18382]));
Q_ASSIGN U14393 ( .B(clk), .A(\g.we_clk [18381]));
Q_ASSIGN U14394 ( .B(clk), .A(\g.we_clk [18380]));
Q_ASSIGN U14395 ( .B(clk), .A(\g.we_clk [18379]));
Q_ASSIGN U14396 ( .B(clk), .A(\g.we_clk [18378]));
Q_ASSIGN U14397 ( .B(clk), .A(\g.we_clk [18377]));
Q_ASSIGN U14398 ( .B(clk), .A(\g.we_clk [18376]));
Q_ASSIGN U14399 ( .B(clk), .A(\g.we_clk [18375]));
Q_ASSIGN U14400 ( .B(clk), .A(\g.we_clk [18374]));
Q_ASSIGN U14401 ( .B(clk), .A(\g.we_clk [18373]));
Q_ASSIGN U14402 ( .B(clk), .A(\g.we_clk [18372]));
Q_ASSIGN U14403 ( .B(clk), .A(\g.we_clk [18371]));
Q_ASSIGN U14404 ( .B(clk), .A(\g.we_clk [18370]));
Q_ASSIGN U14405 ( .B(clk), .A(\g.we_clk [18369]));
Q_ASSIGN U14406 ( .B(clk), .A(\g.we_clk [18368]));
Q_ASSIGN U14407 ( .B(clk), .A(\g.we_clk [18367]));
Q_ASSIGN U14408 ( .B(clk), .A(\g.we_clk [18366]));
Q_ASSIGN U14409 ( .B(clk), .A(\g.we_clk [18365]));
Q_ASSIGN U14410 ( .B(clk), .A(\g.we_clk [18364]));
Q_ASSIGN U14411 ( .B(clk), .A(\g.we_clk [18363]));
Q_ASSIGN U14412 ( .B(clk), .A(\g.we_clk [18362]));
Q_ASSIGN U14413 ( .B(clk), .A(\g.we_clk [18361]));
Q_ASSIGN U14414 ( .B(clk), .A(\g.we_clk [18360]));
Q_ASSIGN U14415 ( .B(clk), .A(\g.we_clk [18359]));
Q_ASSIGN U14416 ( .B(clk), .A(\g.we_clk [18358]));
Q_ASSIGN U14417 ( .B(clk), .A(\g.we_clk [18357]));
Q_ASSIGN U14418 ( .B(clk), .A(\g.we_clk [18356]));
Q_ASSIGN U14419 ( .B(clk), .A(\g.we_clk [18355]));
Q_ASSIGN U14420 ( .B(clk), .A(\g.we_clk [18354]));
Q_ASSIGN U14421 ( .B(clk), .A(\g.we_clk [18353]));
Q_ASSIGN U14422 ( .B(clk), .A(\g.we_clk [18352]));
Q_ASSIGN U14423 ( .B(clk), .A(\g.we_clk [18351]));
Q_ASSIGN U14424 ( .B(clk), .A(\g.we_clk [18350]));
Q_ASSIGN U14425 ( .B(clk), .A(\g.we_clk [18349]));
Q_ASSIGN U14426 ( .B(clk), .A(\g.we_clk [18348]));
Q_ASSIGN U14427 ( .B(clk), .A(\g.we_clk [18347]));
Q_ASSIGN U14428 ( .B(clk), .A(\g.we_clk [18346]));
Q_ASSIGN U14429 ( .B(clk), .A(\g.we_clk [18345]));
Q_ASSIGN U14430 ( .B(clk), .A(\g.we_clk [18344]));
Q_ASSIGN U14431 ( .B(clk), .A(\g.we_clk [18343]));
Q_ASSIGN U14432 ( .B(clk), .A(\g.we_clk [18342]));
Q_ASSIGN U14433 ( .B(clk), .A(\g.we_clk [18341]));
Q_ASSIGN U14434 ( .B(clk), .A(\g.we_clk [18340]));
Q_ASSIGN U14435 ( .B(clk), .A(\g.we_clk [18339]));
Q_ASSIGN U14436 ( .B(clk), .A(\g.we_clk [18338]));
Q_ASSIGN U14437 ( .B(clk), .A(\g.we_clk [18337]));
Q_ASSIGN U14438 ( .B(clk), .A(\g.we_clk [18336]));
Q_ASSIGN U14439 ( .B(clk), .A(\g.we_clk [18335]));
Q_ASSIGN U14440 ( .B(clk), .A(\g.we_clk [18334]));
Q_ASSIGN U14441 ( .B(clk), .A(\g.we_clk [18333]));
Q_ASSIGN U14442 ( .B(clk), .A(\g.we_clk [18332]));
Q_ASSIGN U14443 ( .B(clk), .A(\g.we_clk [18331]));
Q_ASSIGN U14444 ( .B(clk), .A(\g.we_clk [18330]));
Q_ASSIGN U14445 ( .B(clk), .A(\g.we_clk [18329]));
Q_ASSIGN U14446 ( .B(clk), .A(\g.we_clk [18328]));
Q_ASSIGN U14447 ( .B(clk), .A(\g.we_clk [18327]));
Q_ASSIGN U14448 ( .B(clk), .A(\g.we_clk [18326]));
Q_ASSIGN U14449 ( .B(clk), .A(\g.we_clk [18325]));
Q_ASSIGN U14450 ( .B(clk), .A(\g.we_clk [18324]));
Q_ASSIGN U14451 ( .B(clk), .A(\g.we_clk [18323]));
Q_ASSIGN U14452 ( .B(clk), .A(\g.we_clk [18322]));
Q_ASSIGN U14453 ( .B(clk), .A(\g.we_clk [18321]));
Q_ASSIGN U14454 ( .B(clk), .A(\g.we_clk [18320]));
Q_ASSIGN U14455 ( .B(clk), .A(\g.we_clk [18319]));
Q_ASSIGN U14456 ( .B(clk), .A(\g.we_clk [18318]));
Q_ASSIGN U14457 ( .B(clk), .A(\g.we_clk [18317]));
Q_ASSIGN U14458 ( .B(clk), .A(\g.we_clk [18316]));
Q_ASSIGN U14459 ( .B(clk), .A(\g.we_clk [18315]));
Q_ASSIGN U14460 ( .B(clk), .A(\g.we_clk [18314]));
Q_ASSIGN U14461 ( .B(clk), .A(\g.we_clk [18313]));
Q_ASSIGN U14462 ( .B(clk), .A(\g.we_clk [18312]));
Q_ASSIGN U14463 ( .B(clk), .A(\g.we_clk [18311]));
Q_ASSIGN U14464 ( .B(clk), .A(\g.we_clk [18310]));
Q_ASSIGN U14465 ( .B(clk), .A(\g.we_clk [18309]));
Q_ASSIGN U14466 ( .B(clk), .A(\g.we_clk [18308]));
Q_ASSIGN U14467 ( .B(clk), .A(\g.we_clk [18307]));
Q_ASSIGN U14468 ( .B(clk), .A(\g.we_clk [18306]));
Q_ASSIGN U14469 ( .B(clk), .A(\g.we_clk [18305]));
Q_ASSIGN U14470 ( .B(clk), .A(\g.we_clk [18304]));
Q_ASSIGN U14471 ( .B(clk), .A(\g.we_clk [18303]));
Q_ASSIGN U14472 ( .B(clk), .A(\g.we_clk [18302]));
Q_ASSIGN U14473 ( .B(clk), .A(\g.we_clk [18301]));
Q_ASSIGN U14474 ( .B(clk), .A(\g.we_clk [18300]));
Q_ASSIGN U14475 ( .B(clk), .A(\g.we_clk [18299]));
Q_ASSIGN U14476 ( .B(clk), .A(\g.we_clk [18298]));
Q_ASSIGN U14477 ( .B(clk), .A(\g.we_clk [18297]));
Q_ASSIGN U14478 ( .B(clk), .A(\g.we_clk [18296]));
Q_ASSIGN U14479 ( .B(clk), .A(\g.we_clk [18295]));
Q_ASSIGN U14480 ( .B(clk), .A(\g.we_clk [18294]));
Q_ASSIGN U14481 ( .B(clk), .A(\g.we_clk [18293]));
Q_ASSIGN U14482 ( .B(clk), .A(\g.we_clk [18292]));
Q_ASSIGN U14483 ( .B(clk), .A(\g.we_clk [18291]));
Q_ASSIGN U14484 ( .B(clk), .A(\g.we_clk [18290]));
Q_ASSIGN U14485 ( .B(clk), .A(\g.we_clk [18289]));
Q_ASSIGN U14486 ( .B(clk), .A(\g.we_clk [18288]));
Q_ASSIGN U14487 ( .B(clk), .A(\g.we_clk [18287]));
Q_ASSIGN U14488 ( .B(clk), .A(\g.we_clk [18286]));
Q_ASSIGN U14489 ( .B(clk), .A(\g.we_clk [18285]));
Q_ASSIGN U14490 ( .B(clk), .A(\g.we_clk [18284]));
Q_ASSIGN U14491 ( .B(clk), .A(\g.we_clk [18283]));
Q_ASSIGN U14492 ( .B(clk), .A(\g.we_clk [18282]));
Q_ASSIGN U14493 ( .B(clk), .A(\g.we_clk [18281]));
Q_ASSIGN U14494 ( .B(clk), .A(\g.we_clk [18280]));
Q_ASSIGN U14495 ( .B(clk), .A(\g.we_clk [18279]));
Q_ASSIGN U14496 ( .B(clk), .A(\g.we_clk [18278]));
Q_ASSIGN U14497 ( .B(clk), .A(\g.we_clk [18277]));
Q_ASSIGN U14498 ( .B(clk), .A(\g.we_clk [18276]));
Q_ASSIGN U14499 ( .B(clk), .A(\g.we_clk [18275]));
Q_ASSIGN U14500 ( .B(clk), .A(\g.we_clk [18274]));
Q_ASSIGN U14501 ( .B(clk), .A(\g.we_clk [18273]));
Q_ASSIGN U14502 ( .B(clk), .A(\g.we_clk [18272]));
Q_ASSIGN U14503 ( .B(clk), .A(\g.we_clk [18271]));
Q_ASSIGN U14504 ( .B(clk), .A(\g.we_clk [18270]));
Q_ASSIGN U14505 ( .B(clk), .A(\g.we_clk [18269]));
Q_ASSIGN U14506 ( .B(clk), .A(\g.we_clk [18268]));
Q_ASSIGN U14507 ( .B(clk), .A(\g.we_clk [18267]));
Q_ASSIGN U14508 ( .B(clk), .A(\g.we_clk [18266]));
Q_ASSIGN U14509 ( .B(clk), .A(\g.we_clk [18265]));
Q_ASSIGN U14510 ( .B(clk), .A(\g.we_clk [18264]));
Q_ASSIGN U14511 ( .B(clk), .A(\g.we_clk [18263]));
Q_ASSIGN U14512 ( .B(clk), .A(\g.we_clk [18262]));
Q_ASSIGN U14513 ( .B(clk), .A(\g.we_clk [18261]));
Q_ASSIGN U14514 ( .B(clk), .A(\g.we_clk [18260]));
Q_ASSIGN U14515 ( .B(clk), .A(\g.we_clk [18259]));
Q_ASSIGN U14516 ( .B(clk), .A(\g.we_clk [18258]));
Q_ASSIGN U14517 ( .B(clk), .A(\g.we_clk [18257]));
Q_ASSIGN U14518 ( .B(clk), .A(\g.we_clk [18256]));
Q_ASSIGN U14519 ( .B(clk), .A(\g.we_clk [18255]));
Q_ASSIGN U14520 ( .B(clk), .A(\g.we_clk [18254]));
Q_ASSIGN U14521 ( .B(clk), .A(\g.we_clk [18253]));
Q_ASSIGN U14522 ( .B(clk), .A(\g.we_clk [18252]));
Q_ASSIGN U14523 ( .B(clk), .A(\g.we_clk [18251]));
Q_ASSIGN U14524 ( .B(clk), .A(\g.we_clk [18250]));
Q_ASSIGN U14525 ( .B(clk), .A(\g.we_clk [18249]));
Q_ASSIGN U14526 ( .B(clk), .A(\g.we_clk [18248]));
Q_ASSIGN U14527 ( .B(clk), .A(\g.we_clk [18247]));
Q_ASSIGN U14528 ( .B(clk), .A(\g.we_clk [18246]));
Q_ASSIGN U14529 ( .B(clk), .A(\g.we_clk [18245]));
Q_ASSIGN U14530 ( .B(clk), .A(\g.we_clk [18244]));
Q_ASSIGN U14531 ( .B(clk), .A(\g.we_clk [18243]));
Q_ASSIGN U14532 ( .B(clk), .A(\g.we_clk [18242]));
Q_ASSIGN U14533 ( .B(clk), .A(\g.we_clk [18241]));
Q_ASSIGN U14534 ( .B(clk), .A(\g.we_clk [18240]));
Q_ASSIGN U14535 ( .B(clk), .A(\g.we_clk [18239]));
Q_ASSIGN U14536 ( .B(clk), .A(\g.we_clk [18238]));
Q_ASSIGN U14537 ( .B(clk), .A(\g.we_clk [18237]));
Q_ASSIGN U14538 ( .B(clk), .A(\g.we_clk [18236]));
Q_ASSIGN U14539 ( .B(clk), .A(\g.we_clk [18235]));
Q_ASSIGN U14540 ( .B(clk), .A(\g.we_clk [18234]));
Q_ASSIGN U14541 ( .B(clk), .A(\g.we_clk [18233]));
Q_ASSIGN U14542 ( .B(clk), .A(\g.we_clk [18232]));
Q_ASSIGN U14543 ( .B(clk), .A(\g.we_clk [18231]));
Q_ASSIGN U14544 ( .B(clk), .A(\g.we_clk [18230]));
Q_ASSIGN U14545 ( .B(clk), .A(\g.we_clk [18229]));
Q_ASSIGN U14546 ( .B(clk), .A(\g.we_clk [18228]));
Q_ASSIGN U14547 ( .B(clk), .A(\g.we_clk [18227]));
Q_ASSIGN U14548 ( .B(clk), .A(\g.we_clk [18226]));
Q_ASSIGN U14549 ( .B(clk), .A(\g.we_clk [18225]));
Q_ASSIGN U14550 ( .B(clk), .A(\g.we_clk [18224]));
Q_ASSIGN U14551 ( .B(clk), .A(\g.we_clk [18223]));
Q_ASSIGN U14552 ( .B(clk), .A(\g.we_clk [18222]));
Q_ASSIGN U14553 ( .B(clk), .A(\g.we_clk [18221]));
Q_ASSIGN U14554 ( .B(clk), .A(\g.we_clk [18220]));
Q_ASSIGN U14555 ( .B(clk), .A(\g.we_clk [18219]));
Q_ASSIGN U14556 ( .B(clk), .A(\g.we_clk [18218]));
Q_ASSIGN U14557 ( .B(clk), .A(\g.we_clk [18217]));
Q_ASSIGN U14558 ( .B(clk), .A(\g.we_clk [18216]));
Q_ASSIGN U14559 ( .B(clk), .A(\g.we_clk [18215]));
Q_ASSIGN U14560 ( .B(clk), .A(\g.we_clk [18214]));
Q_ASSIGN U14561 ( .B(clk), .A(\g.we_clk [18213]));
Q_ASSIGN U14562 ( .B(clk), .A(\g.we_clk [18212]));
Q_ASSIGN U14563 ( .B(clk), .A(\g.we_clk [18211]));
Q_ASSIGN U14564 ( .B(clk), .A(\g.we_clk [18210]));
Q_ASSIGN U14565 ( .B(clk), .A(\g.we_clk [18209]));
Q_ASSIGN U14566 ( .B(clk), .A(\g.we_clk [18208]));
Q_ASSIGN U14567 ( .B(clk), .A(\g.we_clk [18207]));
Q_ASSIGN U14568 ( .B(clk), .A(\g.we_clk [18206]));
Q_ASSIGN U14569 ( .B(clk), .A(\g.we_clk [18205]));
Q_ASSIGN U14570 ( .B(clk), .A(\g.we_clk [18204]));
Q_ASSIGN U14571 ( .B(clk), .A(\g.we_clk [18203]));
Q_ASSIGN U14572 ( .B(clk), .A(\g.we_clk [18202]));
Q_ASSIGN U14573 ( .B(clk), .A(\g.we_clk [18201]));
Q_ASSIGN U14574 ( .B(clk), .A(\g.we_clk [18200]));
Q_ASSIGN U14575 ( .B(clk), .A(\g.we_clk [18199]));
Q_ASSIGN U14576 ( .B(clk), .A(\g.we_clk [18198]));
Q_ASSIGN U14577 ( .B(clk), .A(\g.we_clk [18197]));
Q_ASSIGN U14578 ( .B(clk), .A(\g.we_clk [18196]));
Q_ASSIGN U14579 ( .B(clk), .A(\g.we_clk [18195]));
Q_ASSIGN U14580 ( .B(clk), .A(\g.we_clk [18194]));
Q_ASSIGN U14581 ( .B(clk), .A(\g.we_clk [18193]));
Q_ASSIGN U14582 ( .B(clk), .A(\g.we_clk [18192]));
Q_ASSIGN U14583 ( .B(clk), .A(\g.we_clk [18191]));
Q_ASSIGN U14584 ( .B(clk), .A(\g.we_clk [18190]));
Q_ASSIGN U14585 ( .B(clk), .A(\g.we_clk [18189]));
Q_ASSIGN U14586 ( .B(clk), .A(\g.we_clk [18188]));
Q_ASSIGN U14587 ( .B(clk), .A(\g.we_clk [18187]));
Q_ASSIGN U14588 ( .B(clk), .A(\g.we_clk [18186]));
Q_ASSIGN U14589 ( .B(clk), .A(\g.we_clk [18185]));
Q_ASSIGN U14590 ( .B(clk), .A(\g.we_clk [18184]));
Q_ASSIGN U14591 ( .B(clk), .A(\g.we_clk [18183]));
Q_ASSIGN U14592 ( .B(clk), .A(\g.we_clk [18182]));
Q_ASSIGN U14593 ( .B(clk), .A(\g.we_clk [18181]));
Q_ASSIGN U14594 ( .B(clk), .A(\g.we_clk [18180]));
Q_ASSIGN U14595 ( .B(clk), .A(\g.we_clk [18179]));
Q_ASSIGN U14596 ( .B(clk), .A(\g.we_clk [18178]));
Q_ASSIGN U14597 ( .B(clk), .A(\g.we_clk [18177]));
Q_ASSIGN U14598 ( .B(clk), .A(\g.we_clk [18176]));
Q_ASSIGN U14599 ( .B(clk), .A(\g.we_clk [18175]));
Q_ASSIGN U14600 ( .B(clk), .A(\g.we_clk [18174]));
Q_ASSIGN U14601 ( .B(clk), .A(\g.we_clk [18173]));
Q_ASSIGN U14602 ( .B(clk), .A(\g.we_clk [18172]));
Q_ASSIGN U14603 ( .B(clk), .A(\g.we_clk [18171]));
Q_ASSIGN U14604 ( .B(clk), .A(\g.we_clk [18170]));
Q_ASSIGN U14605 ( .B(clk), .A(\g.we_clk [18169]));
Q_ASSIGN U14606 ( .B(clk), .A(\g.we_clk [18168]));
Q_ASSIGN U14607 ( .B(clk), .A(\g.we_clk [18167]));
Q_ASSIGN U14608 ( .B(clk), .A(\g.we_clk [18166]));
Q_ASSIGN U14609 ( .B(clk), .A(\g.we_clk [18165]));
Q_ASSIGN U14610 ( .B(clk), .A(\g.we_clk [18164]));
Q_ASSIGN U14611 ( .B(clk), .A(\g.we_clk [18163]));
Q_ASSIGN U14612 ( .B(clk), .A(\g.we_clk [18162]));
Q_ASSIGN U14613 ( .B(clk), .A(\g.we_clk [18161]));
Q_ASSIGN U14614 ( .B(clk), .A(\g.we_clk [18160]));
Q_ASSIGN U14615 ( .B(clk), .A(\g.we_clk [18159]));
Q_ASSIGN U14616 ( .B(clk), .A(\g.we_clk [18158]));
Q_ASSIGN U14617 ( .B(clk), .A(\g.we_clk [18157]));
Q_ASSIGN U14618 ( .B(clk), .A(\g.we_clk [18156]));
Q_ASSIGN U14619 ( .B(clk), .A(\g.we_clk [18155]));
Q_ASSIGN U14620 ( .B(clk), .A(\g.we_clk [18154]));
Q_ASSIGN U14621 ( .B(clk), .A(\g.we_clk [18153]));
Q_ASSIGN U14622 ( .B(clk), .A(\g.we_clk [18152]));
Q_ASSIGN U14623 ( .B(clk), .A(\g.we_clk [18151]));
Q_ASSIGN U14624 ( .B(clk), .A(\g.we_clk [18150]));
Q_ASSIGN U14625 ( .B(clk), .A(\g.we_clk [18149]));
Q_ASSIGN U14626 ( .B(clk), .A(\g.we_clk [18148]));
Q_ASSIGN U14627 ( .B(clk), .A(\g.we_clk [18147]));
Q_ASSIGN U14628 ( .B(clk), .A(\g.we_clk [18146]));
Q_ASSIGN U14629 ( .B(clk), .A(\g.we_clk [18145]));
Q_ASSIGN U14630 ( .B(clk), .A(\g.we_clk [18144]));
Q_ASSIGN U14631 ( .B(clk), .A(\g.we_clk [18143]));
Q_ASSIGN U14632 ( .B(clk), .A(\g.we_clk [18142]));
Q_ASSIGN U14633 ( .B(clk), .A(\g.we_clk [18141]));
Q_ASSIGN U14634 ( .B(clk), .A(\g.we_clk [18140]));
Q_ASSIGN U14635 ( .B(clk), .A(\g.we_clk [18139]));
Q_ASSIGN U14636 ( .B(clk), .A(\g.we_clk [18138]));
Q_ASSIGN U14637 ( .B(clk), .A(\g.we_clk [18137]));
Q_ASSIGN U14638 ( .B(clk), .A(\g.we_clk [18136]));
Q_ASSIGN U14639 ( .B(clk), .A(\g.we_clk [18135]));
Q_ASSIGN U14640 ( .B(clk), .A(\g.we_clk [18134]));
Q_ASSIGN U14641 ( .B(clk), .A(\g.we_clk [18133]));
Q_ASSIGN U14642 ( .B(clk), .A(\g.we_clk [18132]));
Q_ASSIGN U14643 ( .B(clk), .A(\g.we_clk [18131]));
Q_ASSIGN U14644 ( .B(clk), .A(\g.we_clk [18130]));
Q_ASSIGN U14645 ( .B(clk), .A(\g.we_clk [18129]));
Q_ASSIGN U14646 ( .B(clk), .A(\g.we_clk [18128]));
Q_ASSIGN U14647 ( .B(clk), .A(\g.we_clk [18127]));
Q_ASSIGN U14648 ( .B(clk), .A(\g.we_clk [18126]));
Q_ASSIGN U14649 ( .B(clk), .A(\g.we_clk [18125]));
Q_ASSIGN U14650 ( .B(clk), .A(\g.we_clk [18124]));
Q_ASSIGN U14651 ( .B(clk), .A(\g.we_clk [18123]));
Q_ASSIGN U14652 ( .B(clk), .A(\g.we_clk [18122]));
Q_ASSIGN U14653 ( .B(clk), .A(\g.we_clk [18121]));
Q_ASSIGN U14654 ( .B(clk), .A(\g.we_clk [18120]));
Q_ASSIGN U14655 ( .B(clk), .A(\g.we_clk [18119]));
Q_ASSIGN U14656 ( .B(clk), .A(\g.we_clk [18118]));
Q_ASSIGN U14657 ( .B(clk), .A(\g.we_clk [18117]));
Q_ASSIGN U14658 ( .B(clk), .A(\g.we_clk [18116]));
Q_ASSIGN U14659 ( .B(clk), .A(\g.we_clk [18115]));
Q_ASSIGN U14660 ( .B(clk), .A(\g.we_clk [18114]));
Q_ASSIGN U14661 ( .B(clk), .A(\g.we_clk [18113]));
Q_ASSIGN U14662 ( .B(clk), .A(\g.we_clk [18112]));
Q_ASSIGN U14663 ( .B(clk), .A(\g.we_clk [18111]));
Q_ASSIGN U14664 ( .B(clk), .A(\g.we_clk [18110]));
Q_ASSIGN U14665 ( .B(clk), .A(\g.we_clk [18109]));
Q_ASSIGN U14666 ( .B(clk), .A(\g.we_clk [18108]));
Q_ASSIGN U14667 ( .B(clk), .A(\g.we_clk [18107]));
Q_ASSIGN U14668 ( .B(clk), .A(\g.we_clk [18106]));
Q_ASSIGN U14669 ( .B(clk), .A(\g.we_clk [18105]));
Q_ASSIGN U14670 ( .B(clk), .A(\g.we_clk [18104]));
Q_ASSIGN U14671 ( .B(clk), .A(\g.we_clk [18103]));
Q_ASSIGN U14672 ( .B(clk), .A(\g.we_clk [18102]));
Q_ASSIGN U14673 ( .B(clk), .A(\g.we_clk [18101]));
Q_ASSIGN U14674 ( .B(clk), .A(\g.we_clk [18100]));
Q_ASSIGN U14675 ( .B(clk), .A(\g.we_clk [18099]));
Q_ASSIGN U14676 ( .B(clk), .A(\g.we_clk [18098]));
Q_ASSIGN U14677 ( .B(clk), .A(\g.we_clk [18097]));
Q_ASSIGN U14678 ( .B(clk), .A(\g.we_clk [18096]));
Q_ASSIGN U14679 ( .B(clk), .A(\g.we_clk [18095]));
Q_ASSIGN U14680 ( .B(clk), .A(\g.we_clk [18094]));
Q_ASSIGN U14681 ( .B(clk), .A(\g.we_clk [18093]));
Q_ASSIGN U14682 ( .B(clk), .A(\g.we_clk [18092]));
Q_ASSIGN U14683 ( .B(clk), .A(\g.we_clk [18091]));
Q_ASSIGN U14684 ( .B(clk), .A(\g.we_clk [18090]));
Q_ASSIGN U14685 ( .B(clk), .A(\g.we_clk [18089]));
Q_ASSIGN U14686 ( .B(clk), .A(\g.we_clk [18088]));
Q_ASSIGN U14687 ( .B(clk), .A(\g.we_clk [18087]));
Q_ASSIGN U14688 ( .B(clk), .A(\g.we_clk [18086]));
Q_ASSIGN U14689 ( .B(clk), .A(\g.we_clk [18085]));
Q_ASSIGN U14690 ( .B(clk), .A(\g.we_clk [18084]));
Q_ASSIGN U14691 ( .B(clk), .A(\g.we_clk [18083]));
Q_ASSIGN U14692 ( .B(clk), .A(\g.we_clk [18082]));
Q_ASSIGN U14693 ( .B(clk), .A(\g.we_clk [18081]));
Q_ASSIGN U14694 ( .B(clk), .A(\g.we_clk [18080]));
Q_ASSIGN U14695 ( .B(clk), .A(\g.we_clk [18079]));
Q_ASSIGN U14696 ( .B(clk), .A(\g.we_clk [18078]));
Q_ASSIGN U14697 ( .B(clk), .A(\g.we_clk [18077]));
Q_ASSIGN U14698 ( .B(clk), .A(\g.we_clk [18076]));
Q_ASSIGN U14699 ( .B(clk), .A(\g.we_clk [18075]));
Q_ASSIGN U14700 ( .B(clk), .A(\g.we_clk [18074]));
Q_ASSIGN U14701 ( .B(clk), .A(\g.we_clk [18073]));
Q_ASSIGN U14702 ( .B(clk), .A(\g.we_clk [18072]));
Q_ASSIGN U14703 ( .B(clk), .A(\g.we_clk [18071]));
Q_ASSIGN U14704 ( .B(clk), .A(\g.we_clk [18070]));
Q_ASSIGN U14705 ( .B(clk), .A(\g.we_clk [18069]));
Q_ASSIGN U14706 ( .B(clk), .A(\g.we_clk [18068]));
Q_ASSIGN U14707 ( .B(clk), .A(\g.we_clk [18067]));
Q_ASSIGN U14708 ( .B(clk), .A(\g.we_clk [18066]));
Q_ASSIGN U14709 ( .B(clk), .A(\g.we_clk [18065]));
Q_ASSIGN U14710 ( .B(clk), .A(\g.we_clk [18064]));
Q_ASSIGN U14711 ( .B(clk), .A(\g.we_clk [18063]));
Q_ASSIGN U14712 ( .B(clk), .A(\g.we_clk [18062]));
Q_ASSIGN U14713 ( .B(clk), .A(\g.we_clk [18061]));
Q_ASSIGN U14714 ( .B(clk), .A(\g.we_clk [18060]));
Q_ASSIGN U14715 ( .B(clk), .A(\g.we_clk [18059]));
Q_ASSIGN U14716 ( .B(clk), .A(\g.we_clk [18058]));
Q_ASSIGN U14717 ( .B(clk), .A(\g.we_clk [18057]));
Q_ASSIGN U14718 ( .B(clk), .A(\g.we_clk [18056]));
Q_ASSIGN U14719 ( .B(clk), .A(\g.we_clk [18055]));
Q_ASSIGN U14720 ( .B(clk), .A(\g.we_clk [18054]));
Q_ASSIGN U14721 ( .B(clk), .A(\g.we_clk [18053]));
Q_ASSIGN U14722 ( .B(clk), .A(\g.we_clk [18052]));
Q_ASSIGN U14723 ( .B(clk), .A(\g.we_clk [18051]));
Q_ASSIGN U14724 ( .B(clk), .A(\g.we_clk [18050]));
Q_ASSIGN U14725 ( .B(clk), .A(\g.we_clk [18049]));
Q_ASSIGN U14726 ( .B(clk), .A(\g.we_clk [18048]));
Q_ASSIGN U14727 ( .B(clk), .A(\g.we_clk [18047]));
Q_ASSIGN U14728 ( .B(clk), .A(\g.we_clk [18046]));
Q_ASSIGN U14729 ( .B(clk), .A(\g.we_clk [18045]));
Q_ASSIGN U14730 ( .B(clk), .A(\g.we_clk [18044]));
Q_ASSIGN U14731 ( .B(clk), .A(\g.we_clk [18043]));
Q_ASSIGN U14732 ( .B(clk), .A(\g.we_clk [18042]));
Q_ASSIGN U14733 ( .B(clk), .A(\g.we_clk [18041]));
Q_ASSIGN U14734 ( .B(clk), .A(\g.we_clk [18040]));
Q_ASSIGN U14735 ( .B(clk), .A(\g.we_clk [18039]));
Q_ASSIGN U14736 ( .B(clk), .A(\g.we_clk [18038]));
Q_ASSIGN U14737 ( .B(clk), .A(\g.we_clk [18037]));
Q_ASSIGN U14738 ( .B(clk), .A(\g.we_clk [18036]));
Q_ASSIGN U14739 ( .B(clk), .A(\g.we_clk [18035]));
Q_ASSIGN U14740 ( .B(clk), .A(\g.we_clk [18034]));
Q_ASSIGN U14741 ( .B(clk), .A(\g.we_clk [18033]));
Q_ASSIGN U14742 ( .B(clk), .A(\g.we_clk [18032]));
Q_ASSIGN U14743 ( .B(clk), .A(\g.we_clk [18031]));
Q_ASSIGN U14744 ( .B(clk), .A(\g.we_clk [18030]));
Q_ASSIGN U14745 ( .B(clk), .A(\g.we_clk [18029]));
Q_ASSIGN U14746 ( .B(clk), .A(\g.we_clk [18028]));
Q_ASSIGN U14747 ( .B(clk), .A(\g.we_clk [18027]));
Q_ASSIGN U14748 ( .B(clk), .A(\g.we_clk [18026]));
Q_ASSIGN U14749 ( .B(clk), .A(\g.we_clk [18025]));
Q_ASSIGN U14750 ( .B(clk), .A(\g.we_clk [18024]));
Q_ASSIGN U14751 ( .B(clk), .A(\g.we_clk [18023]));
Q_ASSIGN U14752 ( .B(clk), .A(\g.we_clk [18022]));
Q_ASSIGN U14753 ( .B(clk), .A(\g.we_clk [18021]));
Q_ASSIGN U14754 ( .B(clk), .A(\g.we_clk [18020]));
Q_ASSIGN U14755 ( .B(clk), .A(\g.we_clk [18019]));
Q_ASSIGN U14756 ( .B(clk), .A(\g.we_clk [18018]));
Q_ASSIGN U14757 ( .B(clk), .A(\g.we_clk [18017]));
Q_ASSIGN U14758 ( .B(clk), .A(\g.we_clk [18016]));
Q_ASSIGN U14759 ( .B(clk), .A(\g.we_clk [18015]));
Q_ASSIGN U14760 ( .B(clk), .A(\g.we_clk [18014]));
Q_ASSIGN U14761 ( .B(clk), .A(\g.we_clk [18013]));
Q_ASSIGN U14762 ( .B(clk), .A(\g.we_clk [18012]));
Q_ASSIGN U14763 ( .B(clk), .A(\g.we_clk [18011]));
Q_ASSIGN U14764 ( .B(clk), .A(\g.we_clk [18010]));
Q_ASSIGN U14765 ( .B(clk), .A(\g.we_clk [18009]));
Q_ASSIGN U14766 ( .B(clk), .A(\g.we_clk [18008]));
Q_ASSIGN U14767 ( .B(clk), .A(\g.we_clk [18007]));
Q_ASSIGN U14768 ( .B(clk), .A(\g.we_clk [18006]));
Q_ASSIGN U14769 ( .B(clk), .A(\g.we_clk [18005]));
Q_ASSIGN U14770 ( .B(clk), .A(\g.we_clk [18004]));
Q_ASSIGN U14771 ( .B(clk), .A(\g.we_clk [18003]));
Q_ASSIGN U14772 ( .B(clk), .A(\g.we_clk [18002]));
Q_ASSIGN U14773 ( .B(clk), .A(\g.we_clk [18001]));
Q_ASSIGN U14774 ( .B(clk), .A(\g.we_clk [18000]));
Q_ASSIGN U14775 ( .B(clk), .A(\g.we_clk [17999]));
Q_ASSIGN U14776 ( .B(clk), .A(\g.we_clk [17998]));
Q_ASSIGN U14777 ( .B(clk), .A(\g.we_clk [17997]));
Q_ASSIGN U14778 ( .B(clk), .A(\g.we_clk [17996]));
Q_ASSIGN U14779 ( .B(clk), .A(\g.we_clk [17995]));
Q_ASSIGN U14780 ( .B(clk), .A(\g.we_clk [17994]));
Q_ASSIGN U14781 ( .B(clk), .A(\g.we_clk [17993]));
Q_ASSIGN U14782 ( .B(clk), .A(\g.we_clk [17992]));
Q_ASSIGN U14783 ( .B(clk), .A(\g.we_clk [17991]));
Q_ASSIGN U14784 ( .B(clk), .A(\g.we_clk [17990]));
Q_ASSIGN U14785 ( .B(clk), .A(\g.we_clk [17989]));
Q_ASSIGN U14786 ( .B(clk), .A(\g.we_clk [17988]));
Q_ASSIGN U14787 ( .B(clk), .A(\g.we_clk [17987]));
Q_ASSIGN U14788 ( .B(clk), .A(\g.we_clk [17986]));
Q_ASSIGN U14789 ( .B(clk), .A(\g.we_clk [17985]));
Q_ASSIGN U14790 ( .B(clk), .A(\g.we_clk [17984]));
Q_ASSIGN U14791 ( .B(clk), .A(\g.we_clk [17983]));
Q_ASSIGN U14792 ( .B(clk), .A(\g.we_clk [17982]));
Q_ASSIGN U14793 ( .B(clk), .A(\g.we_clk [17981]));
Q_ASSIGN U14794 ( .B(clk), .A(\g.we_clk [17980]));
Q_ASSIGN U14795 ( .B(clk), .A(\g.we_clk [17979]));
Q_ASSIGN U14796 ( .B(clk), .A(\g.we_clk [17978]));
Q_ASSIGN U14797 ( .B(clk), .A(\g.we_clk [17977]));
Q_ASSIGN U14798 ( .B(clk), .A(\g.we_clk [17976]));
Q_ASSIGN U14799 ( .B(clk), .A(\g.we_clk [17975]));
Q_ASSIGN U14800 ( .B(clk), .A(\g.we_clk [17974]));
Q_ASSIGN U14801 ( .B(clk), .A(\g.we_clk [17973]));
Q_ASSIGN U14802 ( .B(clk), .A(\g.we_clk [17972]));
Q_ASSIGN U14803 ( .B(clk), .A(\g.we_clk [17971]));
Q_ASSIGN U14804 ( .B(clk), .A(\g.we_clk [17970]));
Q_ASSIGN U14805 ( .B(clk), .A(\g.we_clk [17969]));
Q_ASSIGN U14806 ( .B(clk), .A(\g.we_clk [17968]));
Q_ASSIGN U14807 ( .B(clk), .A(\g.we_clk [17967]));
Q_ASSIGN U14808 ( .B(clk), .A(\g.we_clk [17966]));
Q_ASSIGN U14809 ( .B(clk), .A(\g.we_clk [17965]));
Q_ASSIGN U14810 ( .B(clk), .A(\g.we_clk [17964]));
Q_ASSIGN U14811 ( .B(clk), .A(\g.we_clk [17963]));
Q_ASSIGN U14812 ( .B(clk), .A(\g.we_clk [17962]));
Q_ASSIGN U14813 ( .B(clk), .A(\g.we_clk [17961]));
Q_ASSIGN U14814 ( .B(clk), .A(\g.we_clk [17960]));
Q_ASSIGN U14815 ( .B(clk), .A(\g.we_clk [17959]));
Q_ASSIGN U14816 ( .B(clk), .A(\g.we_clk [17958]));
Q_ASSIGN U14817 ( .B(clk), .A(\g.we_clk [17957]));
Q_ASSIGN U14818 ( .B(clk), .A(\g.we_clk [17956]));
Q_ASSIGN U14819 ( .B(clk), .A(\g.we_clk [17955]));
Q_ASSIGN U14820 ( .B(clk), .A(\g.we_clk [17954]));
Q_ASSIGN U14821 ( .B(clk), .A(\g.we_clk [17953]));
Q_ASSIGN U14822 ( .B(clk), .A(\g.we_clk [17952]));
Q_ASSIGN U14823 ( .B(clk), .A(\g.we_clk [17951]));
Q_ASSIGN U14824 ( .B(clk), .A(\g.we_clk [17950]));
Q_ASSIGN U14825 ( .B(clk), .A(\g.we_clk [17949]));
Q_ASSIGN U14826 ( .B(clk), .A(\g.we_clk [17948]));
Q_ASSIGN U14827 ( .B(clk), .A(\g.we_clk [17947]));
Q_ASSIGN U14828 ( .B(clk), .A(\g.we_clk [17946]));
Q_ASSIGN U14829 ( .B(clk), .A(\g.we_clk [17945]));
Q_ASSIGN U14830 ( .B(clk), .A(\g.we_clk [17944]));
Q_ASSIGN U14831 ( .B(clk), .A(\g.we_clk [17943]));
Q_ASSIGN U14832 ( .B(clk), .A(\g.we_clk [17942]));
Q_ASSIGN U14833 ( .B(clk), .A(\g.we_clk [17941]));
Q_ASSIGN U14834 ( .B(clk), .A(\g.we_clk [17940]));
Q_ASSIGN U14835 ( .B(clk), .A(\g.we_clk [17939]));
Q_ASSIGN U14836 ( .B(clk), .A(\g.we_clk [17938]));
Q_ASSIGN U14837 ( .B(clk), .A(\g.we_clk [17937]));
Q_ASSIGN U14838 ( .B(clk), .A(\g.we_clk [17936]));
Q_ASSIGN U14839 ( .B(clk), .A(\g.we_clk [17935]));
Q_ASSIGN U14840 ( .B(clk), .A(\g.we_clk [17934]));
Q_ASSIGN U14841 ( .B(clk), .A(\g.we_clk [17933]));
Q_ASSIGN U14842 ( .B(clk), .A(\g.we_clk [17932]));
Q_ASSIGN U14843 ( .B(clk), .A(\g.we_clk [17931]));
Q_ASSIGN U14844 ( .B(clk), .A(\g.we_clk [17930]));
Q_ASSIGN U14845 ( .B(clk), .A(\g.we_clk [17929]));
Q_ASSIGN U14846 ( .B(clk), .A(\g.we_clk [17928]));
Q_ASSIGN U14847 ( .B(clk), .A(\g.we_clk [17927]));
Q_ASSIGN U14848 ( .B(clk), .A(\g.we_clk [17926]));
Q_ASSIGN U14849 ( .B(clk), .A(\g.we_clk [17925]));
Q_ASSIGN U14850 ( .B(clk), .A(\g.we_clk [17924]));
Q_ASSIGN U14851 ( .B(clk), .A(\g.we_clk [17923]));
Q_ASSIGN U14852 ( .B(clk), .A(\g.we_clk [17922]));
Q_ASSIGN U14853 ( .B(clk), .A(\g.we_clk [17921]));
Q_ASSIGN U14854 ( .B(clk), .A(\g.we_clk [17920]));
Q_ASSIGN U14855 ( .B(clk), .A(\g.we_clk [17919]));
Q_ASSIGN U14856 ( .B(clk), .A(\g.we_clk [17918]));
Q_ASSIGN U14857 ( .B(clk), .A(\g.we_clk [17917]));
Q_ASSIGN U14858 ( .B(clk), .A(\g.we_clk [17916]));
Q_ASSIGN U14859 ( .B(clk), .A(\g.we_clk [17915]));
Q_ASSIGN U14860 ( .B(clk), .A(\g.we_clk [17914]));
Q_ASSIGN U14861 ( .B(clk), .A(\g.we_clk [17913]));
Q_ASSIGN U14862 ( .B(clk), .A(\g.we_clk [17912]));
Q_ASSIGN U14863 ( .B(clk), .A(\g.we_clk [17911]));
Q_ASSIGN U14864 ( .B(clk), .A(\g.we_clk [17910]));
Q_ASSIGN U14865 ( .B(clk), .A(\g.we_clk [17909]));
Q_ASSIGN U14866 ( .B(clk), .A(\g.we_clk [17908]));
Q_ASSIGN U14867 ( .B(clk), .A(\g.we_clk [17907]));
Q_ASSIGN U14868 ( .B(clk), .A(\g.we_clk [17906]));
Q_ASSIGN U14869 ( .B(clk), .A(\g.we_clk [17905]));
Q_ASSIGN U14870 ( .B(clk), .A(\g.we_clk [17904]));
Q_ASSIGN U14871 ( .B(clk), .A(\g.we_clk [17903]));
Q_ASSIGN U14872 ( .B(clk), .A(\g.we_clk [17902]));
Q_ASSIGN U14873 ( .B(clk), .A(\g.we_clk [17901]));
Q_ASSIGN U14874 ( .B(clk), .A(\g.we_clk [17900]));
Q_ASSIGN U14875 ( .B(clk), .A(\g.we_clk [17899]));
Q_ASSIGN U14876 ( .B(clk), .A(\g.we_clk [17898]));
Q_ASSIGN U14877 ( .B(clk), .A(\g.we_clk [17897]));
Q_ASSIGN U14878 ( .B(clk), .A(\g.we_clk [17896]));
Q_ASSIGN U14879 ( .B(clk), .A(\g.we_clk [17895]));
Q_ASSIGN U14880 ( .B(clk), .A(\g.we_clk [17894]));
Q_ASSIGN U14881 ( .B(clk), .A(\g.we_clk [17893]));
Q_ASSIGN U14882 ( .B(clk), .A(\g.we_clk [17892]));
Q_ASSIGN U14883 ( .B(clk), .A(\g.we_clk [17891]));
Q_ASSIGN U14884 ( .B(clk), .A(\g.we_clk [17890]));
Q_ASSIGN U14885 ( .B(clk), .A(\g.we_clk [17889]));
Q_ASSIGN U14886 ( .B(clk), .A(\g.we_clk [17888]));
Q_ASSIGN U14887 ( .B(clk), .A(\g.we_clk [17887]));
Q_ASSIGN U14888 ( .B(clk), .A(\g.we_clk [17886]));
Q_ASSIGN U14889 ( .B(clk), .A(\g.we_clk [17885]));
Q_ASSIGN U14890 ( .B(clk), .A(\g.we_clk [17884]));
Q_ASSIGN U14891 ( .B(clk), .A(\g.we_clk [17883]));
Q_ASSIGN U14892 ( .B(clk), .A(\g.we_clk [17882]));
Q_ASSIGN U14893 ( .B(clk), .A(\g.we_clk [17881]));
Q_ASSIGN U14894 ( .B(clk), .A(\g.we_clk [17880]));
Q_ASSIGN U14895 ( .B(clk), .A(\g.we_clk [17879]));
Q_ASSIGN U14896 ( .B(clk), .A(\g.we_clk [17878]));
Q_ASSIGN U14897 ( .B(clk), .A(\g.we_clk [17877]));
Q_ASSIGN U14898 ( .B(clk), .A(\g.we_clk [17876]));
Q_ASSIGN U14899 ( .B(clk), .A(\g.we_clk [17875]));
Q_ASSIGN U14900 ( .B(clk), .A(\g.we_clk [17874]));
Q_ASSIGN U14901 ( .B(clk), .A(\g.we_clk [17873]));
Q_ASSIGN U14902 ( .B(clk), .A(\g.we_clk [17872]));
Q_ASSIGN U14903 ( .B(clk), .A(\g.we_clk [17871]));
Q_ASSIGN U14904 ( .B(clk), .A(\g.we_clk [17870]));
Q_ASSIGN U14905 ( .B(clk), .A(\g.we_clk [17869]));
Q_ASSIGN U14906 ( .B(clk), .A(\g.we_clk [17868]));
Q_ASSIGN U14907 ( .B(clk), .A(\g.we_clk [17867]));
Q_ASSIGN U14908 ( .B(clk), .A(\g.we_clk [17866]));
Q_ASSIGN U14909 ( .B(clk), .A(\g.we_clk [17865]));
Q_ASSIGN U14910 ( .B(clk), .A(\g.we_clk [17864]));
Q_ASSIGN U14911 ( .B(clk), .A(\g.we_clk [17863]));
Q_ASSIGN U14912 ( .B(clk), .A(\g.we_clk [17862]));
Q_ASSIGN U14913 ( .B(clk), .A(\g.we_clk [17861]));
Q_ASSIGN U14914 ( .B(clk), .A(\g.we_clk [17860]));
Q_ASSIGN U14915 ( .B(clk), .A(\g.we_clk [17859]));
Q_ASSIGN U14916 ( .B(clk), .A(\g.we_clk [17858]));
Q_ASSIGN U14917 ( .B(clk), .A(\g.we_clk [17857]));
Q_ASSIGN U14918 ( .B(clk), .A(\g.we_clk [17856]));
Q_ASSIGN U14919 ( .B(clk), .A(\g.we_clk [17855]));
Q_ASSIGN U14920 ( .B(clk), .A(\g.we_clk [17854]));
Q_ASSIGN U14921 ( .B(clk), .A(\g.we_clk [17853]));
Q_ASSIGN U14922 ( .B(clk), .A(\g.we_clk [17852]));
Q_ASSIGN U14923 ( .B(clk), .A(\g.we_clk [17851]));
Q_ASSIGN U14924 ( .B(clk), .A(\g.we_clk [17850]));
Q_ASSIGN U14925 ( .B(clk), .A(\g.we_clk [17849]));
Q_ASSIGN U14926 ( .B(clk), .A(\g.we_clk [17848]));
Q_ASSIGN U14927 ( .B(clk), .A(\g.we_clk [17847]));
Q_ASSIGN U14928 ( .B(clk), .A(\g.we_clk [17846]));
Q_ASSIGN U14929 ( .B(clk), .A(\g.we_clk [17845]));
Q_ASSIGN U14930 ( .B(clk), .A(\g.we_clk [17844]));
Q_ASSIGN U14931 ( .B(clk), .A(\g.we_clk [17843]));
Q_ASSIGN U14932 ( .B(clk), .A(\g.we_clk [17842]));
Q_ASSIGN U14933 ( .B(clk), .A(\g.we_clk [17841]));
Q_ASSIGN U14934 ( .B(clk), .A(\g.we_clk [17840]));
Q_ASSIGN U14935 ( .B(clk), .A(\g.we_clk [17839]));
Q_ASSIGN U14936 ( .B(clk), .A(\g.we_clk [17838]));
Q_ASSIGN U14937 ( .B(clk), .A(\g.we_clk [17837]));
Q_ASSIGN U14938 ( .B(clk), .A(\g.we_clk [17836]));
Q_ASSIGN U14939 ( .B(clk), .A(\g.we_clk [17835]));
Q_ASSIGN U14940 ( .B(clk), .A(\g.we_clk [17834]));
Q_ASSIGN U14941 ( .B(clk), .A(\g.we_clk [17833]));
Q_ASSIGN U14942 ( .B(clk), .A(\g.we_clk [17832]));
Q_ASSIGN U14943 ( .B(clk), .A(\g.we_clk [17831]));
Q_ASSIGN U14944 ( .B(clk), .A(\g.we_clk [17830]));
Q_ASSIGN U14945 ( .B(clk), .A(\g.we_clk [17829]));
Q_ASSIGN U14946 ( .B(clk), .A(\g.we_clk [17828]));
Q_ASSIGN U14947 ( .B(clk), .A(\g.we_clk [17827]));
Q_ASSIGN U14948 ( .B(clk), .A(\g.we_clk [17826]));
Q_ASSIGN U14949 ( .B(clk), .A(\g.we_clk [17825]));
Q_ASSIGN U14950 ( .B(clk), .A(\g.we_clk [17824]));
Q_ASSIGN U14951 ( .B(clk), .A(\g.we_clk [17823]));
Q_ASSIGN U14952 ( .B(clk), .A(\g.we_clk [17822]));
Q_ASSIGN U14953 ( .B(clk), .A(\g.we_clk [17821]));
Q_ASSIGN U14954 ( .B(clk), .A(\g.we_clk [17820]));
Q_ASSIGN U14955 ( .B(clk), .A(\g.we_clk [17819]));
Q_ASSIGN U14956 ( .B(clk), .A(\g.we_clk [17818]));
Q_ASSIGN U14957 ( .B(clk), .A(\g.we_clk [17817]));
Q_ASSIGN U14958 ( .B(clk), .A(\g.we_clk [17816]));
Q_ASSIGN U14959 ( .B(clk), .A(\g.we_clk [17815]));
Q_ASSIGN U14960 ( .B(clk), .A(\g.we_clk [17814]));
Q_ASSIGN U14961 ( .B(clk), .A(\g.we_clk [17813]));
Q_ASSIGN U14962 ( .B(clk), .A(\g.we_clk [17812]));
Q_ASSIGN U14963 ( .B(clk), .A(\g.we_clk [17811]));
Q_ASSIGN U14964 ( .B(clk), .A(\g.we_clk [17810]));
Q_ASSIGN U14965 ( .B(clk), .A(\g.we_clk [17809]));
Q_ASSIGN U14966 ( .B(clk), .A(\g.we_clk [17808]));
Q_ASSIGN U14967 ( .B(clk), .A(\g.we_clk [17807]));
Q_ASSIGN U14968 ( .B(clk), .A(\g.we_clk [17806]));
Q_ASSIGN U14969 ( .B(clk), .A(\g.we_clk [17805]));
Q_ASSIGN U14970 ( .B(clk), .A(\g.we_clk [17804]));
Q_ASSIGN U14971 ( .B(clk), .A(\g.we_clk [17803]));
Q_ASSIGN U14972 ( .B(clk), .A(\g.we_clk [17802]));
Q_ASSIGN U14973 ( .B(clk), .A(\g.we_clk [17801]));
Q_ASSIGN U14974 ( .B(clk), .A(\g.we_clk [17800]));
Q_ASSIGN U14975 ( .B(clk), .A(\g.we_clk [17799]));
Q_ASSIGN U14976 ( .B(clk), .A(\g.we_clk [17798]));
Q_ASSIGN U14977 ( .B(clk), .A(\g.we_clk [17797]));
Q_ASSIGN U14978 ( .B(clk), .A(\g.we_clk [17796]));
Q_ASSIGN U14979 ( .B(clk), .A(\g.we_clk [17795]));
Q_ASSIGN U14980 ( .B(clk), .A(\g.we_clk [17794]));
Q_ASSIGN U14981 ( .B(clk), .A(\g.we_clk [17793]));
Q_ASSIGN U14982 ( .B(clk), .A(\g.we_clk [17792]));
Q_ASSIGN U14983 ( .B(clk), .A(\g.we_clk [17791]));
Q_ASSIGN U14984 ( .B(clk), .A(\g.we_clk [17790]));
Q_ASSIGN U14985 ( .B(clk), .A(\g.we_clk [17789]));
Q_ASSIGN U14986 ( .B(clk), .A(\g.we_clk [17788]));
Q_ASSIGN U14987 ( .B(clk), .A(\g.we_clk [17787]));
Q_ASSIGN U14988 ( .B(clk), .A(\g.we_clk [17786]));
Q_ASSIGN U14989 ( .B(clk), .A(\g.we_clk [17785]));
Q_ASSIGN U14990 ( .B(clk), .A(\g.we_clk [17784]));
Q_ASSIGN U14991 ( .B(clk), .A(\g.we_clk [17783]));
Q_ASSIGN U14992 ( .B(clk), .A(\g.we_clk [17782]));
Q_ASSIGN U14993 ( .B(clk), .A(\g.we_clk [17781]));
Q_ASSIGN U14994 ( .B(clk), .A(\g.we_clk [17780]));
Q_ASSIGN U14995 ( .B(clk), .A(\g.we_clk [17779]));
Q_ASSIGN U14996 ( .B(clk), .A(\g.we_clk [17778]));
Q_ASSIGN U14997 ( .B(clk), .A(\g.we_clk [17777]));
Q_ASSIGN U14998 ( .B(clk), .A(\g.we_clk [17776]));
Q_ASSIGN U14999 ( .B(clk), .A(\g.we_clk [17775]));
Q_ASSIGN U15000 ( .B(clk), .A(\g.we_clk [17774]));
Q_ASSIGN U15001 ( .B(clk), .A(\g.we_clk [17773]));
Q_ASSIGN U15002 ( .B(clk), .A(\g.we_clk [17772]));
Q_ASSIGN U15003 ( .B(clk), .A(\g.we_clk [17771]));
Q_ASSIGN U15004 ( .B(clk), .A(\g.we_clk [17770]));
Q_ASSIGN U15005 ( .B(clk), .A(\g.we_clk [17769]));
Q_ASSIGN U15006 ( .B(clk), .A(\g.we_clk [17768]));
Q_ASSIGN U15007 ( .B(clk), .A(\g.we_clk [17767]));
Q_ASSIGN U15008 ( .B(clk), .A(\g.we_clk [17766]));
Q_ASSIGN U15009 ( .B(clk), .A(\g.we_clk [17765]));
Q_ASSIGN U15010 ( .B(clk), .A(\g.we_clk [17764]));
Q_ASSIGN U15011 ( .B(clk), .A(\g.we_clk [17763]));
Q_ASSIGN U15012 ( .B(clk), .A(\g.we_clk [17762]));
Q_ASSIGN U15013 ( .B(clk), .A(\g.we_clk [17761]));
Q_ASSIGN U15014 ( .B(clk), .A(\g.we_clk [17760]));
Q_ASSIGN U15015 ( .B(clk), .A(\g.we_clk [17759]));
Q_ASSIGN U15016 ( .B(clk), .A(\g.we_clk [17758]));
Q_ASSIGN U15017 ( .B(clk), .A(\g.we_clk [17757]));
Q_ASSIGN U15018 ( .B(clk), .A(\g.we_clk [17756]));
Q_ASSIGN U15019 ( .B(clk), .A(\g.we_clk [17755]));
Q_ASSIGN U15020 ( .B(clk), .A(\g.we_clk [17754]));
Q_ASSIGN U15021 ( .B(clk), .A(\g.we_clk [17753]));
Q_ASSIGN U15022 ( .B(clk), .A(\g.we_clk [17752]));
Q_ASSIGN U15023 ( .B(clk), .A(\g.we_clk [17751]));
Q_ASSIGN U15024 ( .B(clk), .A(\g.we_clk [17750]));
Q_ASSIGN U15025 ( .B(clk), .A(\g.we_clk [17749]));
Q_ASSIGN U15026 ( .B(clk), .A(\g.we_clk [17748]));
Q_ASSIGN U15027 ( .B(clk), .A(\g.we_clk [17747]));
Q_ASSIGN U15028 ( .B(clk), .A(\g.we_clk [17746]));
Q_ASSIGN U15029 ( .B(clk), .A(\g.we_clk [17745]));
Q_ASSIGN U15030 ( .B(clk), .A(\g.we_clk [17744]));
Q_ASSIGN U15031 ( .B(clk), .A(\g.we_clk [17743]));
Q_ASSIGN U15032 ( .B(clk), .A(\g.we_clk [17742]));
Q_ASSIGN U15033 ( .B(clk), .A(\g.we_clk [17741]));
Q_ASSIGN U15034 ( .B(clk), .A(\g.we_clk [17740]));
Q_ASSIGN U15035 ( .B(clk), .A(\g.we_clk [17739]));
Q_ASSIGN U15036 ( .B(clk), .A(\g.we_clk [17738]));
Q_ASSIGN U15037 ( .B(clk), .A(\g.we_clk [17737]));
Q_ASSIGN U15038 ( .B(clk), .A(\g.we_clk [17736]));
Q_ASSIGN U15039 ( .B(clk), .A(\g.we_clk [17735]));
Q_ASSIGN U15040 ( .B(clk), .A(\g.we_clk [17734]));
Q_ASSIGN U15041 ( .B(clk), .A(\g.we_clk [17733]));
Q_ASSIGN U15042 ( .B(clk), .A(\g.we_clk [17732]));
Q_ASSIGN U15043 ( .B(clk), .A(\g.we_clk [17731]));
Q_ASSIGN U15044 ( .B(clk), .A(\g.we_clk [17730]));
Q_ASSIGN U15045 ( .B(clk), .A(\g.we_clk [17729]));
Q_ASSIGN U15046 ( .B(clk), .A(\g.we_clk [17728]));
Q_ASSIGN U15047 ( .B(clk), .A(\g.we_clk [17727]));
Q_ASSIGN U15048 ( .B(clk), .A(\g.we_clk [17726]));
Q_ASSIGN U15049 ( .B(clk), .A(\g.we_clk [17725]));
Q_ASSIGN U15050 ( .B(clk), .A(\g.we_clk [17724]));
Q_ASSIGN U15051 ( .B(clk), .A(\g.we_clk [17723]));
Q_ASSIGN U15052 ( .B(clk), .A(\g.we_clk [17722]));
Q_ASSIGN U15053 ( .B(clk), .A(\g.we_clk [17721]));
Q_ASSIGN U15054 ( .B(clk), .A(\g.we_clk [17720]));
Q_ASSIGN U15055 ( .B(clk), .A(\g.we_clk [17719]));
Q_ASSIGN U15056 ( .B(clk), .A(\g.we_clk [17718]));
Q_ASSIGN U15057 ( .B(clk), .A(\g.we_clk [17717]));
Q_ASSIGN U15058 ( .B(clk), .A(\g.we_clk [17716]));
Q_ASSIGN U15059 ( .B(clk), .A(\g.we_clk [17715]));
Q_ASSIGN U15060 ( .B(clk), .A(\g.we_clk [17714]));
Q_ASSIGN U15061 ( .B(clk), .A(\g.we_clk [17713]));
Q_ASSIGN U15062 ( .B(clk), .A(\g.we_clk [17712]));
Q_ASSIGN U15063 ( .B(clk), .A(\g.we_clk [17711]));
Q_ASSIGN U15064 ( .B(clk), .A(\g.we_clk [17710]));
Q_ASSIGN U15065 ( .B(clk), .A(\g.we_clk [17709]));
Q_ASSIGN U15066 ( .B(clk), .A(\g.we_clk [17708]));
Q_ASSIGN U15067 ( .B(clk), .A(\g.we_clk [17707]));
Q_ASSIGN U15068 ( .B(clk), .A(\g.we_clk [17706]));
Q_ASSIGN U15069 ( .B(clk), .A(\g.we_clk [17705]));
Q_ASSIGN U15070 ( .B(clk), .A(\g.we_clk [17704]));
Q_ASSIGN U15071 ( .B(clk), .A(\g.we_clk [17703]));
Q_ASSIGN U15072 ( .B(clk), .A(\g.we_clk [17702]));
Q_ASSIGN U15073 ( .B(clk), .A(\g.we_clk [17701]));
Q_ASSIGN U15074 ( .B(clk), .A(\g.we_clk [17700]));
Q_ASSIGN U15075 ( .B(clk), .A(\g.we_clk [17699]));
Q_ASSIGN U15076 ( .B(clk), .A(\g.we_clk [17698]));
Q_ASSIGN U15077 ( .B(clk), .A(\g.we_clk [17697]));
Q_ASSIGN U15078 ( .B(clk), .A(\g.we_clk [17696]));
Q_ASSIGN U15079 ( .B(clk), .A(\g.we_clk [17695]));
Q_ASSIGN U15080 ( .B(clk), .A(\g.we_clk [17694]));
Q_ASSIGN U15081 ( .B(clk), .A(\g.we_clk [17693]));
Q_ASSIGN U15082 ( .B(clk), .A(\g.we_clk [17692]));
Q_ASSIGN U15083 ( .B(clk), .A(\g.we_clk [17691]));
Q_ASSIGN U15084 ( .B(clk), .A(\g.we_clk [17690]));
Q_ASSIGN U15085 ( .B(clk), .A(\g.we_clk [17689]));
Q_ASSIGN U15086 ( .B(clk), .A(\g.we_clk [17688]));
Q_ASSIGN U15087 ( .B(clk), .A(\g.we_clk [17687]));
Q_ASSIGN U15088 ( .B(clk), .A(\g.we_clk [17686]));
Q_ASSIGN U15089 ( .B(clk), .A(\g.we_clk [17685]));
Q_ASSIGN U15090 ( .B(clk), .A(\g.we_clk [17684]));
Q_ASSIGN U15091 ( .B(clk), .A(\g.we_clk [17683]));
Q_ASSIGN U15092 ( .B(clk), .A(\g.we_clk [17682]));
Q_ASSIGN U15093 ( .B(clk), .A(\g.we_clk [17681]));
Q_ASSIGN U15094 ( .B(clk), .A(\g.we_clk [17680]));
Q_ASSIGN U15095 ( .B(clk), .A(\g.we_clk [17679]));
Q_ASSIGN U15096 ( .B(clk), .A(\g.we_clk [17678]));
Q_ASSIGN U15097 ( .B(clk), .A(\g.we_clk [17677]));
Q_ASSIGN U15098 ( .B(clk), .A(\g.we_clk [17676]));
Q_ASSIGN U15099 ( .B(clk), .A(\g.we_clk [17675]));
Q_ASSIGN U15100 ( .B(clk), .A(\g.we_clk [17674]));
Q_ASSIGN U15101 ( .B(clk), .A(\g.we_clk [17673]));
Q_ASSIGN U15102 ( .B(clk), .A(\g.we_clk [17672]));
Q_ASSIGN U15103 ( .B(clk), .A(\g.we_clk [17671]));
Q_ASSIGN U15104 ( .B(clk), .A(\g.we_clk [17670]));
Q_ASSIGN U15105 ( .B(clk), .A(\g.we_clk [17669]));
Q_ASSIGN U15106 ( .B(clk), .A(\g.we_clk [17668]));
Q_ASSIGN U15107 ( .B(clk), .A(\g.we_clk [17667]));
Q_ASSIGN U15108 ( .B(clk), .A(\g.we_clk [17666]));
Q_ASSIGN U15109 ( .B(clk), .A(\g.we_clk [17665]));
Q_ASSIGN U15110 ( .B(clk), .A(\g.we_clk [17664]));
Q_ASSIGN U15111 ( .B(clk), .A(\g.we_clk [17663]));
Q_ASSIGN U15112 ( .B(clk), .A(\g.we_clk [17662]));
Q_ASSIGN U15113 ( .B(clk), .A(\g.we_clk [17661]));
Q_ASSIGN U15114 ( .B(clk), .A(\g.we_clk [17660]));
Q_ASSIGN U15115 ( .B(clk), .A(\g.we_clk [17659]));
Q_ASSIGN U15116 ( .B(clk), .A(\g.we_clk [17658]));
Q_ASSIGN U15117 ( .B(clk), .A(\g.we_clk [17657]));
Q_ASSIGN U15118 ( .B(clk), .A(\g.we_clk [17656]));
Q_ASSIGN U15119 ( .B(clk), .A(\g.we_clk [17655]));
Q_ASSIGN U15120 ( .B(clk), .A(\g.we_clk [17654]));
Q_ASSIGN U15121 ( .B(clk), .A(\g.we_clk [17653]));
Q_ASSIGN U15122 ( .B(clk), .A(\g.we_clk [17652]));
Q_ASSIGN U15123 ( .B(clk), .A(\g.we_clk [17651]));
Q_ASSIGN U15124 ( .B(clk), .A(\g.we_clk [17650]));
Q_ASSIGN U15125 ( .B(clk), .A(\g.we_clk [17649]));
Q_ASSIGN U15126 ( .B(clk), .A(\g.we_clk [17648]));
Q_ASSIGN U15127 ( .B(clk), .A(\g.we_clk [17647]));
Q_ASSIGN U15128 ( .B(clk), .A(\g.we_clk [17646]));
Q_ASSIGN U15129 ( .B(clk), .A(\g.we_clk [17645]));
Q_ASSIGN U15130 ( .B(clk), .A(\g.we_clk [17644]));
Q_ASSIGN U15131 ( .B(clk), .A(\g.we_clk [17643]));
Q_ASSIGN U15132 ( .B(clk), .A(\g.we_clk [17642]));
Q_ASSIGN U15133 ( .B(clk), .A(\g.we_clk [17641]));
Q_ASSIGN U15134 ( .B(clk), .A(\g.we_clk [17640]));
Q_ASSIGN U15135 ( .B(clk), .A(\g.we_clk [17639]));
Q_ASSIGN U15136 ( .B(clk), .A(\g.we_clk [17638]));
Q_ASSIGN U15137 ( .B(clk), .A(\g.we_clk [17637]));
Q_ASSIGN U15138 ( .B(clk), .A(\g.we_clk [17636]));
Q_ASSIGN U15139 ( .B(clk), .A(\g.we_clk [17635]));
Q_ASSIGN U15140 ( .B(clk), .A(\g.we_clk [17634]));
Q_ASSIGN U15141 ( .B(clk), .A(\g.we_clk [17633]));
Q_ASSIGN U15142 ( .B(clk), .A(\g.we_clk [17632]));
Q_ASSIGN U15143 ( .B(clk), .A(\g.we_clk [17631]));
Q_ASSIGN U15144 ( .B(clk), .A(\g.we_clk [17630]));
Q_ASSIGN U15145 ( .B(clk), .A(\g.we_clk [17629]));
Q_ASSIGN U15146 ( .B(clk), .A(\g.we_clk [17628]));
Q_ASSIGN U15147 ( .B(clk), .A(\g.we_clk [17627]));
Q_ASSIGN U15148 ( .B(clk), .A(\g.we_clk [17626]));
Q_ASSIGN U15149 ( .B(clk), .A(\g.we_clk [17625]));
Q_ASSIGN U15150 ( .B(clk), .A(\g.we_clk [17624]));
Q_ASSIGN U15151 ( .B(clk), .A(\g.we_clk [17623]));
Q_ASSIGN U15152 ( .B(clk), .A(\g.we_clk [17622]));
Q_ASSIGN U15153 ( .B(clk), .A(\g.we_clk [17621]));
Q_ASSIGN U15154 ( .B(clk), .A(\g.we_clk [17620]));
Q_ASSIGN U15155 ( .B(clk), .A(\g.we_clk [17619]));
Q_ASSIGN U15156 ( .B(clk), .A(\g.we_clk [17618]));
Q_ASSIGN U15157 ( .B(clk), .A(\g.we_clk [17617]));
Q_ASSIGN U15158 ( .B(clk), .A(\g.we_clk [17616]));
Q_ASSIGN U15159 ( .B(clk), .A(\g.we_clk [17615]));
Q_ASSIGN U15160 ( .B(clk), .A(\g.we_clk [17614]));
Q_ASSIGN U15161 ( .B(clk), .A(\g.we_clk [17613]));
Q_ASSIGN U15162 ( .B(clk), .A(\g.we_clk [17612]));
Q_ASSIGN U15163 ( .B(clk), .A(\g.we_clk [17611]));
Q_ASSIGN U15164 ( .B(clk), .A(\g.we_clk [17610]));
Q_ASSIGN U15165 ( .B(clk), .A(\g.we_clk [17609]));
Q_ASSIGN U15166 ( .B(clk), .A(\g.we_clk [17608]));
Q_ASSIGN U15167 ( .B(clk), .A(\g.we_clk [17607]));
Q_ASSIGN U15168 ( .B(clk), .A(\g.we_clk [17606]));
Q_ASSIGN U15169 ( .B(clk), .A(\g.we_clk [17605]));
Q_ASSIGN U15170 ( .B(clk), .A(\g.we_clk [17604]));
Q_ASSIGN U15171 ( .B(clk), .A(\g.we_clk [17603]));
Q_ASSIGN U15172 ( .B(clk), .A(\g.we_clk [17602]));
Q_ASSIGN U15173 ( .B(clk), .A(\g.we_clk [17601]));
Q_ASSIGN U15174 ( .B(clk), .A(\g.we_clk [17600]));
Q_ASSIGN U15175 ( .B(clk), .A(\g.we_clk [17599]));
Q_ASSIGN U15176 ( .B(clk), .A(\g.we_clk [17598]));
Q_ASSIGN U15177 ( .B(clk), .A(\g.we_clk [17597]));
Q_ASSIGN U15178 ( .B(clk), .A(\g.we_clk [17596]));
Q_ASSIGN U15179 ( .B(clk), .A(\g.we_clk [17595]));
Q_ASSIGN U15180 ( .B(clk), .A(\g.we_clk [17594]));
Q_ASSIGN U15181 ( .B(clk), .A(\g.we_clk [17593]));
Q_ASSIGN U15182 ( .B(clk), .A(\g.we_clk [17592]));
Q_ASSIGN U15183 ( .B(clk), .A(\g.we_clk [17591]));
Q_ASSIGN U15184 ( .B(clk), .A(\g.we_clk [17590]));
Q_ASSIGN U15185 ( .B(clk), .A(\g.we_clk [17589]));
Q_ASSIGN U15186 ( .B(clk), .A(\g.we_clk [17588]));
Q_ASSIGN U15187 ( .B(clk), .A(\g.we_clk [17587]));
Q_ASSIGN U15188 ( .B(clk), .A(\g.we_clk [17586]));
Q_ASSIGN U15189 ( .B(clk), .A(\g.we_clk [17585]));
Q_ASSIGN U15190 ( .B(clk), .A(\g.we_clk [17584]));
Q_ASSIGN U15191 ( .B(clk), .A(\g.we_clk [17583]));
Q_ASSIGN U15192 ( .B(clk), .A(\g.we_clk [17582]));
Q_ASSIGN U15193 ( .B(clk), .A(\g.we_clk [17581]));
Q_ASSIGN U15194 ( .B(clk), .A(\g.we_clk [17580]));
Q_ASSIGN U15195 ( .B(clk), .A(\g.we_clk [17579]));
Q_ASSIGN U15196 ( .B(clk), .A(\g.we_clk [17578]));
Q_ASSIGN U15197 ( .B(clk), .A(\g.we_clk [17577]));
Q_ASSIGN U15198 ( .B(clk), .A(\g.we_clk [17576]));
Q_ASSIGN U15199 ( .B(clk), .A(\g.we_clk [17575]));
Q_ASSIGN U15200 ( .B(clk), .A(\g.we_clk [17574]));
Q_ASSIGN U15201 ( .B(clk), .A(\g.we_clk [17573]));
Q_ASSIGN U15202 ( .B(clk), .A(\g.we_clk [17572]));
Q_ASSIGN U15203 ( .B(clk), .A(\g.we_clk [17571]));
Q_ASSIGN U15204 ( .B(clk), .A(\g.we_clk [17570]));
Q_ASSIGN U15205 ( .B(clk), .A(\g.we_clk [17569]));
Q_ASSIGN U15206 ( .B(clk), .A(\g.we_clk [17568]));
Q_ASSIGN U15207 ( .B(clk), .A(\g.we_clk [17567]));
Q_ASSIGN U15208 ( .B(clk), .A(\g.we_clk [17566]));
Q_ASSIGN U15209 ( .B(clk), .A(\g.we_clk [17565]));
Q_ASSIGN U15210 ( .B(clk), .A(\g.we_clk [17564]));
Q_ASSIGN U15211 ( .B(clk), .A(\g.we_clk [17563]));
Q_ASSIGN U15212 ( .B(clk), .A(\g.we_clk [17562]));
Q_ASSIGN U15213 ( .B(clk), .A(\g.we_clk [17561]));
Q_ASSIGN U15214 ( .B(clk), .A(\g.we_clk [17560]));
Q_ASSIGN U15215 ( .B(clk), .A(\g.we_clk [17559]));
Q_ASSIGN U15216 ( .B(clk), .A(\g.we_clk [17558]));
Q_ASSIGN U15217 ( .B(clk), .A(\g.we_clk [17557]));
Q_ASSIGN U15218 ( .B(clk), .A(\g.we_clk [17556]));
Q_ASSIGN U15219 ( .B(clk), .A(\g.we_clk [17555]));
Q_ASSIGN U15220 ( .B(clk), .A(\g.we_clk [17554]));
Q_ASSIGN U15221 ( .B(clk), .A(\g.we_clk [17553]));
Q_ASSIGN U15222 ( .B(clk), .A(\g.we_clk [17552]));
Q_ASSIGN U15223 ( .B(clk), .A(\g.we_clk [17551]));
Q_ASSIGN U15224 ( .B(clk), .A(\g.we_clk [17550]));
Q_ASSIGN U15225 ( .B(clk), .A(\g.we_clk [17549]));
Q_ASSIGN U15226 ( .B(clk), .A(\g.we_clk [17548]));
Q_ASSIGN U15227 ( .B(clk), .A(\g.we_clk [17547]));
Q_ASSIGN U15228 ( .B(clk), .A(\g.we_clk [17546]));
Q_ASSIGN U15229 ( .B(clk), .A(\g.we_clk [17545]));
Q_ASSIGN U15230 ( .B(clk), .A(\g.we_clk [17544]));
Q_ASSIGN U15231 ( .B(clk), .A(\g.we_clk [17543]));
Q_ASSIGN U15232 ( .B(clk), .A(\g.we_clk [17542]));
Q_ASSIGN U15233 ( .B(clk), .A(\g.we_clk [17541]));
Q_ASSIGN U15234 ( .B(clk), .A(\g.we_clk [17540]));
Q_ASSIGN U15235 ( .B(clk), .A(\g.we_clk [17539]));
Q_ASSIGN U15236 ( .B(clk), .A(\g.we_clk [17538]));
Q_ASSIGN U15237 ( .B(clk), .A(\g.we_clk [17537]));
Q_ASSIGN U15238 ( .B(clk), .A(\g.we_clk [17536]));
Q_ASSIGN U15239 ( .B(clk), .A(\g.we_clk [17535]));
Q_ASSIGN U15240 ( .B(clk), .A(\g.we_clk [17534]));
Q_ASSIGN U15241 ( .B(clk), .A(\g.we_clk [17533]));
Q_ASSIGN U15242 ( .B(clk), .A(\g.we_clk [17532]));
Q_ASSIGN U15243 ( .B(clk), .A(\g.we_clk [17531]));
Q_ASSIGN U15244 ( .B(clk), .A(\g.we_clk [17530]));
Q_ASSIGN U15245 ( .B(clk), .A(\g.we_clk [17529]));
Q_ASSIGN U15246 ( .B(clk), .A(\g.we_clk [17528]));
Q_ASSIGN U15247 ( .B(clk), .A(\g.we_clk [17527]));
Q_ASSIGN U15248 ( .B(clk), .A(\g.we_clk [17526]));
Q_ASSIGN U15249 ( .B(clk), .A(\g.we_clk [17525]));
Q_ASSIGN U15250 ( .B(clk), .A(\g.we_clk [17524]));
Q_ASSIGN U15251 ( .B(clk), .A(\g.we_clk [17523]));
Q_ASSIGN U15252 ( .B(clk), .A(\g.we_clk [17522]));
Q_ASSIGN U15253 ( .B(clk), .A(\g.we_clk [17521]));
Q_ASSIGN U15254 ( .B(clk), .A(\g.we_clk [17520]));
Q_ASSIGN U15255 ( .B(clk), .A(\g.we_clk [17519]));
Q_ASSIGN U15256 ( .B(clk), .A(\g.we_clk [17518]));
Q_ASSIGN U15257 ( .B(clk), .A(\g.we_clk [17517]));
Q_ASSIGN U15258 ( .B(clk), .A(\g.we_clk [17516]));
Q_ASSIGN U15259 ( .B(clk), .A(\g.we_clk [17515]));
Q_ASSIGN U15260 ( .B(clk), .A(\g.we_clk [17514]));
Q_ASSIGN U15261 ( .B(clk), .A(\g.we_clk [17513]));
Q_ASSIGN U15262 ( .B(clk), .A(\g.we_clk [17512]));
Q_ASSIGN U15263 ( .B(clk), .A(\g.we_clk [17511]));
Q_ASSIGN U15264 ( .B(clk), .A(\g.we_clk [17510]));
Q_ASSIGN U15265 ( .B(clk), .A(\g.we_clk [17509]));
Q_ASSIGN U15266 ( .B(clk), .A(\g.we_clk [17508]));
Q_ASSIGN U15267 ( .B(clk), .A(\g.we_clk [17507]));
Q_ASSIGN U15268 ( .B(clk), .A(\g.we_clk [17506]));
Q_ASSIGN U15269 ( .B(clk), .A(\g.we_clk [17505]));
Q_ASSIGN U15270 ( .B(clk), .A(\g.we_clk [17504]));
Q_ASSIGN U15271 ( .B(clk), .A(\g.we_clk [17503]));
Q_ASSIGN U15272 ( .B(clk), .A(\g.we_clk [17502]));
Q_ASSIGN U15273 ( .B(clk), .A(\g.we_clk [17501]));
Q_ASSIGN U15274 ( .B(clk), .A(\g.we_clk [17500]));
Q_ASSIGN U15275 ( .B(clk), .A(\g.we_clk [17499]));
Q_ASSIGN U15276 ( .B(clk), .A(\g.we_clk [17498]));
Q_ASSIGN U15277 ( .B(clk), .A(\g.we_clk [17497]));
Q_ASSIGN U15278 ( .B(clk), .A(\g.we_clk [17496]));
Q_ASSIGN U15279 ( .B(clk), .A(\g.we_clk [17495]));
Q_ASSIGN U15280 ( .B(clk), .A(\g.we_clk [17494]));
Q_ASSIGN U15281 ( .B(clk), .A(\g.we_clk [17493]));
Q_ASSIGN U15282 ( .B(clk), .A(\g.we_clk [17492]));
Q_ASSIGN U15283 ( .B(clk), .A(\g.we_clk [17491]));
Q_ASSIGN U15284 ( .B(clk), .A(\g.we_clk [17490]));
Q_ASSIGN U15285 ( .B(clk), .A(\g.we_clk [17489]));
Q_ASSIGN U15286 ( .B(clk), .A(\g.we_clk [17488]));
Q_ASSIGN U15287 ( .B(clk), .A(\g.we_clk [17487]));
Q_ASSIGN U15288 ( .B(clk), .A(\g.we_clk [17486]));
Q_ASSIGN U15289 ( .B(clk), .A(\g.we_clk [17485]));
Q_ASSIGN U15290 ( .B(clk), .A(\g.we_clk [17484]));
Q_ASSIGN U15291 ( .B(clk), .A(\g.we_clk [17483]));
Q_ASSIGN U15292 ( .B(clk), .A(\g.we_clk [17482]));
Q_ASSIGN U15293 ( .B(clk), .A(\g.we_clk [17481]));
Q_ASSIGN U15294 ( .B(clk), .A(\g.we_clk [17480]));
Q_ASSIGN U15295 ( .B(clk), .A(\g.we_clk [17479]));
Q_ASSIGN U15296 ( .B(clk), .A(\g.we_clk [17478]));
Q_ASSIGN U15297 ( .B(clk), .A(\g.we_clk [17477]));
Q_ASSIGN U15298 ( .B(clk), .A(\g.we_clk [17476]));
Q_ASSIGN U15299 ( .B(clk), .A(\g.we_clk [17475]));
Q_ASSIGN U15300 ( .B(clk), .A(\g.we_clk [17474]));
Q_ASSIGN U15301 ( .B(clk), .A(\g.we_clk [17473]));
Q_ASSIGN U15302 ( .B(clk), .A(\g.we_clk [17472]));
Q_ASSIGN U15303 ( .B(clk), .A(\g.we_clk [17471]));
Q_ASSIGN U15304 ( .B(clk), .A(\g.we_clk [17470]));
Q_ASSIGN U15305 ( .B(clk), .A(\g.we_clk [17469]));
Q_ASSIGN U15306 ( .B(clk), .A(\g.we_clk [17468]));
Q_ASSIGN U15307 ( .B(clk), .A(\g.we_clk [17467]));
Q_ASSIGN U15308 ( .B(clk), .A(\g.we_clk [17466]));
Q_ASSIGN U15309 ( .B(clk), .A(\g.we_clk [17465]));
Q_ASSIGN U15310 ( .B(clk), .A(\g.we_clk [17464]));
Q_ASSIGN U15311 ( .B(clk), .A(\g.we_clk [17463]));
Q_ASSIGN U15312 ( .B(clk), .A(\g.we_clk [17462]));
Q_ASSIGN U15313 ( .B(clk), .A(\g.we_clk [17461]));
Q_ASSIGN U15314 ( .B(clk), .A(\g.we_clk [17460]));
Q_ASSIGN U15315 ( .B(clk), .A(\g.we_clk [17459]));
Q_ASSIGN U15316 ( .B(clk), .A(\g.we_clk [17458]));
Q_ASSIGN U15317 ( .B(clk), .A(\g.we_clk [17457]));
Q_ASSIGN U15318 ( .B(clk), .A(\g.we_clk [17456]));
Q_ASSIGN U15319 ( .B(clk), .A(\g.we_clk [17455]));
Q_ASSIGN U15320 ( .B(clk), .A(\g.we_clk [17454]));
Q_ASSIGN U15321 ( .B(clk), .A(\g.we_clk [17453]));
Q_ASSIGN U15322 ( .B(clk), .A(\g.we_clk [17452]));
Q_ASSIGN U15323 ( .B(clk), .A(\g.we_clk [17451]));
Q_ASSIGN U15324 ( .B(clk), .A(\g.we_clk [17450]));
Q_ASSIGN U15325 ( .B(clk), .A(\g.we_clk [17449]));
Q_ASSIGN U15326 ( .B(clk), .A(\g.we_clk [17448]));
Q_ASSIGN U15327 ( .B(clk), .A(\g.we_clk [17447]));
Q_ASSIGN U15328 ( .B(clk), .A(\g.we_clk [17446]));
Q_ASSIGN U15329 ( .B(clk), .A(\g.we_clk [17445]));
Q_ASSIGN U15330 ( .B(clk), .A(\g.we_clk [17444]));
Q_ASSIGN U15331 ( .B(clk), .A(\g.we_clk [17443]));
Q_ASSIGN U15332 ( .B(clk), .A(\g.we_clk [17442]));
Q_ASSIGN U15333 ( .B(clk), .A(\g.we_clk [17441]));
Q_ASSIGN U15334 ( .B(clk), .A(\g.we_clk [17440]));
Q_ASSIGN U15335 ( .B(clk), .A(\g.we_clk [17439]));
Q_ASSIGN U15336 ( .B(clk), .A(\g.we_clk [17438]));
Q_ASSIGN U15337 ( .B(clk), .A(\g.we_clk [17437]));
Q_ASSIGN U15338 ( .B(clk), .A(\g.we_clk [17436]));
Q_ASSIGN U15339 ( .B(clk), .A(\g.we_clk [17435]));
Q_ASSIGN U15340 ( .B(clk), .A(\g.we_clk [17434]));
Q_ASSIGN U15341 ( .B(clk), .A(\g.we_clk [17433]));
Q_ASSIGN U15342 ( .B(clk), .A(\g.we_clk [17432]));
Q_ASSIGN U15343 ( .B(clk), .A(\g.we_clk [17431]));
Q_ASSIGN U15344 ( .B(clk), .A(\g.we_clk [17430]));
Q_ASSIGN U15345 ( .B(clk), .A(\g.we_clk [17429]));
Q_ASSIGN U15346 ( .B(clk), .A(\g.we_clk [17428]));
Q_ASSIGN U15347 ( .B(clk), .A(\g.we_clk [17427]));
Q_ASSIGN U15348 ( .B(clk), .A(\g.we_clk [17426]));
Q_ASSIGN U15349 ( .B(clk), .A(\g.we_clk [17425]));
Q_ASSIGN U15350 ( .B(clk), .A(\g.we_clk [17424]));
Q_ASSIGN U15351 ( .B(clk), .A(\g.we_clk [17423]));
Q_ASSIGN U15352 ( .B(clk), .A(\g.we_clk [17422]));
Q_ASSIGN U15353 ( .B(clk), .A(\g.we_clk [17421]));
Q_ASSIGN U15354 ( .B(clk), .A(\g.we_clk [17420]));
Q_ASSIGN U15355 ( .B(clk), .A(\g.we_clk [17419]));
Q_ASSIGN U15356 ( .B(clk), .A(\g.we_clk [17418]));
Q_ASSIGN U15357 ( .B(clk), .A(\g.we_clk [17417]));
Q_ASSIGN U15358 ( .B(clk), .A(\g.we_clk [17416]));
Q_ASSIGN U15359 ( .B(clk), .A(\g.we_clk [17415]));
Q_ASSIGN U15360 ( .B(clk), .A(\g.we_clk [17414]));
Q_ASSIGN U15361 ( .B(clk), .A(\g.we_clk [17413]));
Q_ASSIGN U15362 ( .B(clk), .A(\g.we_clk [17412]));
Q_ASSIGN U15363 ( .B(clk), .A(\g.we_clk [17411]));
Q_ASSIGN U15364 ( .B(clk), .A(\g.we_clk [17410]));
Q_ASSIGN U15365 ( .B(clk), .A(\g.we_clk [17409]));
Q_ASSIGN U15366 ( .B(clk), .A(\g.we_clk [17408]));
Q_ASSIGN U15367 ( .B(clk), .A(\g.we_clk [17407]));
Q_ASSIGN U15368 ( .B(clk), .A(\g.we_clk [17406]));
Q_ASSIGN U15369 ( .B(clk), .A(\g.we_clk [17405]));
Q_ASSIGN U15370 ( .B(clk), .A(\g.we_clk [17404]));
Q_ASSIGN U15371 ( .B(clk), .A(\g.we_clk [17403]));
Q_ASSIGN U15372 ( .B(clk), .A(\g.we_clk [17402]));
Q_ASSIGN U15373 ( .B(clk), .A(\g.we_clk [17401]));
Q_ASSIGN U15374 ( .B(clk), .A(\g.we_clk [17400]));
Q_ASSIGN U15375 ( .B(clk), .A(\g.we_clk [17399]));
Q_ASSIGN U15376 ( .B(clk), .A(\g.we_clk [17398]));
Q_ASSIGN U15377 ( .B(clk), .A(\g.we_clk [17397]));
Q_ASSIGN U15378 ( .B(clk), .A(\g.we_clk [17396]));
Q_ASSIGN U15379 ( .B(clk), .A(\g.we_clk [17395]));
Q_ASSIGN U15380 ( .B(clk), .A(\g.we_clk [17394]));
Q_ASSIGN U15381 ( .B(clk), .A(\g.we_clk [17393]));
Q_ASSIGN U15382 ( .B(clk), .A(\g.we_clk [17392]));
Q_ASSIGN U15383 ( .B(clk), .A(\g.we_clk [17391]));
Q_ASSIGN U15384 ( .B(clk), .A(\g.we_clk [17390]));
Q_ASSIGN U15385 ( .B(clk), .A(\g.we_clk [17389]));
Q_ASSIGN U15386 ( .B(clk), .A(\g.we_clk [17388]));
Q_ASSIGN U15387 ( .B(clk), .A(\g.we_clk [17387]));
Q_ASSIGN U15388 ( .B(clk), .A(\g.we_clk [17386]));
Q_ASSIGN U15389 ( .B(clk), .A(\g.we_clk [17385]));
Q_ASSIGN U15390 ( .B(clk), .A(\g.we_clk [17384]));
Q_ASSIGN U15391 ( .B(clk), .A(\g.we_clk [17383]));
Q_ASSIGN U15392 ( .B(clk), .A(\g.we_clk [17382]));
Q_ASSIGN U15393 ( .B(clk), .A(\g.we_clk [17381]));
Q_ASSIGN U15394 ( .B(clk), .A(\g.we_clk [17380]));
Q_ASSIGN U15395 ( .B(clk), .A(\g.we_clk [17379]));
Q_ASSIGN U15396 ( .B(clk), .A(\g.we_clk [17378]));
Q_ASSIGN U15397 ( .B(clk), .A(\g.we_clk [17377]));
Q_ASSIGN U15398 ( .B(clk), .A(\g.we_clk [17376]));
Q_ASSIGN U15399 ( .B(clk), .A(\g.we_clk [17375]));
Q_ASSIGN U15400 ( .B(clk), .A(\g.we_clk [17374]));
Q_ASSIGN U15401 ( .B(clk), .A(\g.we_clk [17373]));
Q_ASSIGN U15402 ( .B(clk), .A(\g.we_clk [17372]));
Q_ASSIGN U15403 ( .B(clk), .A(\g.we_clk [17371]));
Q_ASSIGN U15404 ( .B(clk), .A(\g.we_clk [17370]));
Q_ASSIGN U15405 ( .B(clk), .A(\g.we_clk [17369]));
Q_ASSIGN U15406 ( .B(clk), .A(\g.we_clk [17368]));
Q_ASSIGN U15407 ( .B(clk), .A(\g.we_clk [17367]));
Q_ASSIGN U15408 ( .B(clk), .A(\g.we_clk [17366]));
Q_ASSIGN U15409 ( .B(clk), .A(\g.we_clk [17365]));
Q_ASSIGN U15410 ( .B(clk), .A(\g.we_clk [17364]));
Q_ASSIGN U15411 ( .B(clk), .A(\g.we_clk [17363]));
Q_ASSIGN U15412 ( .B(clk), .A(\g.we_clk [17362]));
Q_ASSIGN U15413 ( .B(clk), .A(\g.we_clk [17361]));
Q_ASSIGN U15414 ( .B(clk), .A(\g.we_clk [17360]));
Q_ASSIGN U15415 ( .B(clk), .A(\g.we_clk [17359]));
Q_ASSIGN U15416 ( .B(clk), .A(\g.we_clk [17358]));
Q_ASSIGN U15417 ( .B(clk), .A(\g.we_clk [17357]));
Q_ASSIGN U15418 ( .B(clk), .A(\g.we_clk [17356]));
Q_ASSIGN U15419 ( .B(clk), .A(\g.we_clk [17355]));
Q_ASSIGN U15420 ( .B(clk), .A(\g.we_clk [17354]));
Q_ASSIGN U15421 ( .B(clk), .A(\g.we_clk [17353]));
Q_ASSIGN U15422 ( .B(clk), .A(\g.we_clk [17352]));
Q_ASSIGN U15423 ( .B(clk), .A(\g.we_clk [17351]));
Q_ASSIGN U15424 ( .B(clk), .A(\g.we_clk [17350]));
Q_ASSIGN U15425 ( .B(clk), .A(\g.we_clk [17349]));
Q_ASSIGN U15426 ( .B(clk), .A(\g.we_clk [17348]));
Q_ASSIGN U15427 ( .B(clk), .A(\g.we_clk [17347]));
Q_ASSIGN U15428 ( .B(clk), .A(\g.we_clk [17346]));
Q_ASSIGN U15429 ( .B(clk), .A(\g.we_clk [17345]));
Q_ASSIGN U15430 ( .B(clk), .A(\g.we_clk [17344]));
Q_ASSIGN U15431 ( .B(clk), .A(\g.we_clk [17343]));
Q_ASSIGN U15432 ( .B(clk), .A(\g.we_clk [17342]));
Q_ASSIGN U15433 ( .B(clk), .A(\g.we_clk [17341]));
Q_ASSIGN U15434 ( .B(clk), .A(\g.we_clk [17340]));
Q_ASSIGN U15435 ( .B(clk), .A(\g.we_clk [17339]));
Q_ASSIGN U15436 ( .B(clk), .A(\g.we_clk [17338]));
Q_ASSIGN U15437 ( .B(clk), .A(\g.we_clk [17337]));
Q_ASSIGN U15438 ( .B(clk), .A(\g.we_clk [17336]));
Q_ASSIGN U15439 ( .B(clk), .A(\g.we_clk [17335]));
Q_ASSIGN U15440 ( .B(clk), .A(\g.we_clk [17334]));
Q_ASSIGN U15441 ( .B(clk), .A(\g.we_clk [17333]));
Q_ASSIGN U15442 ( .B(clk), .A(\g.we_clk [17332]));
Q_ASSIGN U15443 ( .B(clk), .A(\g.we_clk [17331]));
Q_ASSIGN U15444 ( .B(clk), .A(\g.we_clk [17330]));
Q_ASSIGN U15445 ( .B(clk), .A(\g.we_clk [17329]));
Q_ASSIGN U15446 ( .B(clk), .A(\g.we_clk [17328]));
Q_ASSIGN U15447 ( .B(clk), .A(\g.we_clk [17327]));
Q_ASSIGN U15448 ( .B(clk), .A(\g.we_clk [17326]));
Q_ASSIGN U15449 ( .B(clk), .A(\g.we_clk [17325]));
Q_ASSIGN U15450 ( .B(clk), .A(\g.we_clk [17324]));
Q_ASSIGN U15451 ( .B(clk), .A(\g.we_clk [17323]));
Q_ASSIGN U15452 ( .B(clk), .A(\g.we_clk [17322]));
Q_ASSIGN U15453 ( .B(clk), .A(\g.we_clk [17321]));
Q_ASSIGN U15454 ( .B(clk), .A(\g.we_clk [17320]));
Q_ASSIGN U15455 ( .B(clk), .A(\g.we_clk [17319]));
Q_ASSIGN U15456 ( .B(clk), .A(\g.we_clk [17318]));
Q_ASSIGN U15457 ( .B(clk), .A(\g.we_clk [17317]));
Q_ASSIGN U15458 ( .B(clk), .A(\g.we_clk [17316]));
Q_ASSIGN U15459 ( .B(clk), .A(\g.we_clk [17315]));
Q_ASSIGN U15460 ( .B(clk), .A(\g.we_clk [17314]));
Q_ASSIGN U15461 ( .B(clk), .A(\g.we_clk [17313]));
Q_ASSIGN U15462 ( .B(clk), .A(\g.we_clk [17312]));
Q_ASSIGN U15463 ( .B(clk), .A(\g.we_clk [17311]));
Q_ASSIGN U15464 ( .B(clk), .A(\g.we_clk [17310]));
Q_ASSIGN U15465 ( .B(clk), .A(\g.we_clk [17309]));
Q_ASSIGN U15466 ( .B(clk), .A(\g.we_clk [17308]));
Q_ASSIGN U15467 ( .B(clk), .A(\g.we_clk [17307]));
Q_ASSIGN U15468 ( .B(clk), .A(\g.we_clk [17306]));
Q_ASSIGN U15469 ( .B(clk), .A(\g.we_clk [17305]));
Q_ASSIGN U15470 ( .B(clk), .A(\g.we_clk [17304]));
Q_ASSIGN U15471 ( .B(clk), .A(\g.we_clk [17303]));
Q_ASSIGN U15472 ( .B(clk), .A(\g.we_clk [17302]));
Q_ASSIGN U15473 ( .B(clk), .A(\g.we_clk [17301]));
Q_ASSIGN U15474 ( .B(clk), .A(\g.we_clk [17300]));
Q_ASSIGN U15475 ( .B(clk), .A(\g.we_clk [17299]));
Q_ASSIGN U15476 ( .B(clk), .A(\g.we_clk [17298]));
Q_ASSIGN U15477 ( .B(clk), .A(\g.we_clk [17297]));
Q_ASSIGN U15478 ( .B(clk), .A(\g.we_clk [17296]));
Q_ASSIGN U15479 ( .B(clk), .A(\g.we_clk [17295]));
Q_ASSIGN U15480 ( .B(clk), .A(\g.we_clk [17294]));
Q_ASSIGN U15481 ( .B(clk), .A(\g.we_clk [17293]));
Q_ASSIGN U15482 ( .B(clk), .A(\g.we_clk [17292]));
Q_ASSIGN U15483 ( .B(clk), .A(\g.we_clk [17291]));
Q_ASSIGN U15484 ( .B(clk), .A(\g.we_clk [17290]));
Q_ASSIGN U15485 ( .B(clk), .A(\g.we_clk [17289]));
Q_ASSIGN U15486 ( .B(clk), .A(\g.we_clk [17288]));
Q_ASSIGN U15487 ( .B(clk), .A(\g.we_clk [17287]));
Q_ASSIGN U15488 ( .B(clk), .A(\g.we_clk [17286]));
Q_ASSIGN U15489 ( .B(clk), .A(\g.we_clk [17285]));
Q_ASSIGN U15490 ( .B(clk), .A(\g.we_clk [17284]));
Q_ASSIGN U15491 ( .B(clk), .A(\g.we_clk [17283]));
Q_ASSIGN U15492 ( .B(clk), .A(\g.we_clk [17282]));
Q_ASSIGN U15493 ( .B(clk), .A(\g.we_clk [17281]));
Q_ASSIGN U15494 ( .B(clk), .A(\g.we_clk [17280]));
Q_ASSIGN U15495 ( .B(clk), .A(\g.we_clk [17279]));
Q_ASSIGN U15496 ( .B(clk), .A(\g.we_clk [17278]));
Q_ASSIGN U15497 ( .B(clk), .A(\g.we_clk [17277]));
Q_ASSIGN U15498 ( .B(clk), .A(\g.we_clk [17276]));
Q_ASSIGN U15499 ( .B(clk), .A(\g.we_clk [17275]));
Q_ASSIGN U15500 ( .B(clk), .A(\g.we_clk [17274]));
Q_ASSIGN U15501 ( .B(clk), .A(\g.we_clk [17273]));
Q_ASSIGN U15502 ( .B(clk), .A(\g.we_clk [17272]));
Q_ASSIGN U15503 ( .B(clk), .A(\g.we_clk [17271]));
Q_ASSIGN U15504 ( .B(clk), .A(\g.we_clk [17270]));
Q_ASSIGN U15505 ( .B(clk), .A(\g.we_clk [17269]));
Q_ASSIGN U15506 ( .B(clk), .A(\g.we_clk [17268]));
Q_ASSIGN U15507 ( .B(clk), .A(\g.we_clk [17267]));
Q_ASSIGN U15508 ( .B(clk), .A(\g.we_clk [17266]));
Q_ASSIGN U15509 ( .B(clk), .A(\g.we_clk [17265]));
Q_ASSIGN U15510 ( .B(clk), .A(\g.we_clk [17264]));
Q_ASSIGN U15511 ( .B(clk), .A(\g.we_clk [17263]));
Q_ASSIGN U15512 ( .B(clk), .A(\g.we_clk [17262]));
Q_ASSIGN U15513 ( .B(clk), .A(\g.we_clk [17261]));
Q_ASSIGN U15514 ( .B(clk), .A(\g.we_clk [17260]));
Q_ASSIGN U15515 ( .B(clk), .A(\g.we_clk [17259]));
Q_ASSIGN U15516 ( .B(clk), .A(\g.we_clk [17258]));
Q_ASSIGN U15517 ( .B(clk), .A(\g.we_clk [17257]));
Q_ASSIGN U15518 ( .B(clk), .A(\g.we_clk [17256]));
Q_ASSIGN U15519 ( .B(clk), .A(\g.we_clk [17255]));
Q_ASSIGN U15520 ( .B(clk), .A(\g.we_clk [17254]));
Q_ASSIGN U15521 ( .B(clk), .A(\g.we_clk [17253]));
Q_ASSIGN U15522 ( .B(clk), .A(\g.we_clk [17252]));
Q_ASSIGN U15523 ( .B(clk), .A(\g.we_clk [17251]));
Q_ASSIGN U15524 ( .B(clk), .A(\g.we_clk [17250]));
Q_ASSIGN U15525 ( .B(clk), .A(\g.we_clk [17249]));
Q_ASSIGN U15526 ( .B(clk), .A(\g.we_clk [17248]));
Q_ASSIGN U15527 ( .B(clk), .A(\g.we_clk [17247]));
Q_ASSIGN U15528 ( .B(clk), .A(\g.we_clk [17246]));
Q_ASSIGN U15529 ( .B(clk), .A(\g.we_clk [17245]));
Q_ASSIGN U15530 ( .B(clk), .A(\g.we_clk [17244]));
Q_ASSIGN U15531 ( .B(clk), .A(\g.we_clk [17243]));
Q_ASSIGN U15532 ( .B(clk), .A(\g.we_clk [17242]));
Q_ASSIGN U15533 ( .B(clk), .A(\g.we_clk [17241]));
Q_ASSIGN U15534 ( .B(clk), .A(\g.we_clk [17240]));
Q_ASSIGN U15535 ( .B(clk), .A(\g.we_clk [17239]));
Q_ASSIGN U15536 ( .B(clk), .A(\g.we_clk [17238]));
Q_ASSIGN U15537 ( .B(clk), .A(\g.we_clk [17237]));
Q_ASSIGN U15538 ( .B(clk), .A(\g.we_clk [17236]));
Q_ASSIGN U15539 ( .B(clk), .A(\g.we_clk [17235]));
Q_ASSIGN U15540 ( .B(clk), .A(\g.we_clk [17234]));
Q_ASSIGN U15541 ( .B(clk), .A(\g.we_clk [17233]));
Q_ASSIGN U15542 ( .B(clk), .A(\g.we_clk [17232]));
Q_ASSIGN U15543 ( .B(clk), .A(\g.we_clk [17231]));
Q_ASSIGN U15544 ( .B(clk), .A(\g.we_clk [17230]));
Q_ASSIGN U15545 ( .B(clk), .A(\g.we_clk [17229]));
Q_ASSIGN U15546 ( .B(clk), .A(\g.we_clk [17228]));
Q_ASSIGN U15547 ( .B(clk), .A(\g.we_clk [17227]));
Q_ASSIGN U15548 ( .B(clk), .A(\g.we_clk [17226]));
Q_ASSIGN U15549 ( .B(clk), .A(\g.we_clk [17225]));
Q_ASSIGN U15550 ( .B(clk), .A(\g.we_clk [17224]));
Q_ASSIGN U15551 ( .B(clk), .A(\g.we_clk [17223]));
Q_ASSIGN U15552 ( .B(clk), .A(\g.we_clk [17222]));
Q_ASSIGN U15553 ( .B(clk), .A(\g.we_clk [17221]));
Q_ASSIGN U15554 ( .B(clk), .A(\g.we_clk [17220]));
Q_ASSIGN U15555 ( .B(clk), .A(\g.we_clk [17219]));
Q_ASSIGN U15556 ( .B(clk), .A(\g.we_clk [17218]));
Q_ASSIGN U15557 ( .B(clk), .A(\g.we_clk [17217]));
Q_ASSIGN U15558 ( .B(clk), .A(\g.we_clk [17216]));
Q_ASSIGN U15559 ( .B(clk), .A(\g.we_clk [17215]));
Q_ASSIGN U15560 ( .B(clk), .A(\g.we_clk [17214]));
Q_ASSIGN U15561 ( .B(clk), .A(\g.we_clk [17213]));
Q_ASSIGN U15562 ( .B(clk), .A(\g.we_clk [17212]));
Q_ASSIGN U15563 ( .B(clk), .A(\g.we_clk [17211]));
Q_ASSIGN U15564 ( .B(clk), .A(\g.we_clk [17210]));
Q_ASSIGN U15565 ( .B(clk), .A(\g.we_clk [17209]));
Q_ASSIGN U15566 ( .B(clk), .A(\g.we_clk [17208]));
Q_ASSIGN U15567 ( .B(clk), .A(\g.we_clk [17207]));
Q_ASSIGN U15568 ( .B(clk), .A(\g.we_clk [17206]));
Q_ASSIGN U15569 ( .B(clk), .A(\g.we_clk [17205]));
Q_ASSIGN U15570 ( .B(clk), .A(\g.we_clk [17204]));
Q_ASSIGN U15571 ( .B(clk), .A(\g.we_clk [17203]));
Q_ASSIGN U15572 ( .B(clk), .A(\g.we_clk [17202]));
Q_ASSIGN U15573 ( .B(clk), .A(\g.we_clk [17201]));
Q_ASSIGN U15574 ( .B(clk), .A(\g.we_clk [17200]));
Q_ASSIGN U15575 ( .B(clk), .A(\g.we_clk [17199]));
Q_ASSIGN U15576 ( .B(clk), .A(\g.we_clk [17198]));
Q_ASSIGN U15577 ( .B(clk), .A(\g.we_clk [17197]));
Q_ASSIGN U15578 ( .B(clk), .A(\g.we_clk [17196]));
Q_ASSIGN U15579 ( .B(clk), .A(\g.we_clk [17195]));
Q_ASSIGN U15580 ( .B(clk), .A(\g.we_clk [17194]));
Q_ASSIGN U15581 ( .B(clk), .A(\g.we_clk [17193]));
Q_ASSIGN U15582 ( .B(clk), .A(\g.we_clk [17192]));
Q_ASSIGN U15583 ( .B(clk), .A(\g.we_clk [17191]));
Q_ASSIGN U15584 ( .B(clk), .A(\g.we_clk [17190]));
Q_ASSIGN U15585 ( .B(clk), .A(\g.we_clk [17189]));
Q_ASSIGN U15586 ( .B(clk), .A(\g.we_clk [17188]));
Q_ASSIGN U15587 ( .B(clk), .A(\g.we_clk [17187]));
Q_ASSIGN U15588 ( .B(clk), .A(\g.we_clk [17186]));
Q_ASSIGN U15589 ( .B(clk), .A(\g.we_clk [17185]));
Q_ASSIGN U15590 ( .B(clk), .A(\g.we_clk [17184]));
Q_ASSIGN U15591 ( .B(clk), .A(\g.we_clk [17183]));
Q_ASSIGN U15592 ( .B(clk), .A(\g.we_clk [17182]));
Q_ASSIGN U15593 ( .B(clk), .A(\g.we_clk [17181]));
Q_ASSIGN U15594 ( .B(clk), .A(\g.we_clk [17180]));
Q_ASSIGN U15595 ( .B(clk), .A(\g.we_clk [17179]));
Q_ASSIGN U15596 ( .B(clk), .A(\g.we_clk [17178]));
Q_ASSIGN U15597 ( .B(clk), .A(\g.we_clk [17177]));
Q_ASSIGN U15598 ( .B(clk), .A(\g.we_clk [17176]));
Q_ASSIGN U15599 ( .B(clk), .A(\g.we_clk [17175]));
Q_ASSIGN U15600 ( .B(clk), .A(\g.we_clk [17174]));
Q_ASSIGN U15601 ( .B(clk), .A(\g.we_clk [17173]));
Q_ASSIGN U15602 ( .B(clk), .A(\g.we_clk [17172]));
Q_ASSIGN U15603 ( .B(clk), .A(\g.we_clk [17171]));
Q_ASSIGN U15604 ( .B(clk), .A(\g.we_clk [17170]));
Q_ASSIGN U15605 ( .B(clk), .A(\g.we_clk [17169]));
Q_ASSIGN U15606 ( .B(clk), .A(\g.we_clk [17168]));
Q_ASSIGN U15607 ( .B(clk), .A(\g.we_clk [17167]));
Q_ASSIGN U15608 ( .B(clk), .A(\g.we_clk [17166]));
Q_ASSIGN U15609 ( .B(clk), .A(\g.we_clk [17165]));
Q_ASSIGN U15610 ( .B(clk), .A(\g.we_clk [17164]));
Q_ASSIGN U15611 ( .B(clk), .A(\g.we_clk [17163]));
Q_ASSIGN U15612 ( .B(clk), .A(\g.we_clk [17162]));
Q_ASSIGN U15613 ( .B(clk), .A(\g.we_clk [17161]));
Q_ASSIGN U15614 ( .B(clk), .A(\g.we_clk [17160]));
Q_ASSIGN U15615 ( .B(clk), .A(\g.we_clk [17159]));
Q_ASSIGN U15616 ( .B(clk), .A(\g.we_clk [17158]));
Q_ASSIGN U15617 ( .B(clk), .A(\g.we_clk [17157]));
Q_ASSIGN U15618 ( .B(clk), .A(\g.we_clk [17156]));
Q_ASSIGN U15619 ( .B(clk), .A(\g.we_clk [17155]));
Q_ASSIGN U15620 ( .B(clk), .A(\g.we_clk [17154]));
Q_ASSIGN U15621 ( .B(clk), .A(\g.we_clk [17153]));
Q_ASSIGN U15622 ( .B(clk), .A(\g.we_clk [17152]));
Q_ASSIGN U15623 ( .B(clk), .A(\g.we_clk [17151]));
Q_ASSIGN U15624 ( .B(clk), .A(\g.we_clk [17150]));
Q_ASSIGN U15625 ( .B(clk), .A(\g.we_clk [17149]));
Q_ASSIGN U15626 ( .B(clk), .A(\g.we_clk [17148]));
Q_ASSIGN U15627 ( .B(clk), .A(\g.we_clk [17147]));
Q_ASSIGN U15628 ( .B(clk), .A(\g.we_clk [17146]));
Q_ASSIGN U15629 ( .B(clk), .A(\g.we_clk [17145]));
Q_ASSIGN U15630 ( .B(clk), .A(\g.we_clk [17144]));
Q_ASSIGN U15631 ( .B(clk), .A(\g.we_clk [17143]));
Q_ASSIGN U15632 ( .B(clk), .A(\g.we_clk [17142]));
Q_ASSIGN U15633 ( .B(clk), .A(\g.we_clk [17141]));
Q_ASSIGN U15634 ( .B(clk), .A(\g.we_clk [17140]));
Q_ASSIGN U15635 ( .B(clk), .A(\g.we_clk [17139]));
Q_ASSIGN U15636 ( .B(clk), .A(\g.we_clk [17138]));
Q_ASSIGN U15637 ( .B(clk), .A(\g.we_clk [17137]));
Q_ASSIGN U15638 ( .B(clk), .A(\g.we_clk [17136]));
Q_ASSIGN U15639 ( .B(clk), .A(\g.we_clk [17135]));
Q_ASSIGN U15640 ( .B(clk), .A(\g.we_clk [17134]));
Q_ASSIGN U15641 ( .B(clk), .A(\g.we_clk [17133]));
Q_ASSIGN U15642 ( .B(clk), .A(\g.we_clk [17132]));
Q_ASSIGN U15643 ( .B(clk), .A(\g.we_clk [17131]));
Q_ASSIGN U15644 ( .B(clk), .A(\g.we_clk [17130]));
Q_ASSIGN U15645 ( .B(clk), .A(\g.we_clk [17129]));
Q_ASSIGN U15646 ( .B(clk), .A(\g.we_clk [17128]));
Q_ASSIGN U15647 ( .B(clk), .A(\g.we_clk [17127]));
Q_ASSIGN U15648 ( .B(clk), .A(\g.we_clk [17126]));
Q_ASSIGN U15649 ( .B(clk), .A(\g.we_clk [17125]));
Q_ASSIGN U15650 ( .B(clk), .A(\g.we_clk [17124]));
Q_ASSIGN U15651 ( .B(clk), .A(\g.we_clk [17123]));
Q_ASSIGN U15652 ( .B(clk), .A(\g.we_clk [17122]));
Q_ASSIGN U15653 ( .B(clk), .A(\g.we_clk [17121]));
Q_ASSIGN U15654 ( .B(clk), .A(\g.we_clk [17120]));
Q_ASSIGN U15655 ( .B(clk), .A(\g.we_clk [17119]));
Q_ASSIGN U15656 ( .B(clk), .A(\g.we_clk [17118]));
Q_ASSIGN U15657 ( .B(clk), .A(\g.we_clk [17117]));
Q_ASSIGN U15658 ( .B(clk), .A(\g.we_clk [17116]));
Q_ASSIGN U15659 ( .B(clk), .A(\g.we_clk [17115]));
Q_ASSIGN U15660 ( .B(clk), .A(\g.we_clk [17114]));
Q_ASSIGN U15661 ( .B(clk), .A(\g.we_clk [17113]));
Q_ASSIGN U15662 ( .B(clk), .A(\g.we_clk [17112]));
Q_ASSIGN U15663 ( .B(clk), .A(\g.we_clk [17111]));
Q_ASSIGN U15664 ( .B(clk), .A(\g.we_clk [17110]));
Q_ASSIGN U15665 ( .B(clk), .A(\g.we_clk [17109]));
Q_ASSIGN U15666 ( .B(clk), .A(\g.we_clk [17108]));
Q_ASSIGN U15667 ( .B(clk), .A(\g.we_clk [17107]));
Q_ASSIGN U15668 ( .B(clk), .A(\g.we_clk [17106]));
Q_ASSIGN U15669 ( .B(clk), .A(\g.we_clk [17105]));
Q_ASSIGN U15670 ( .B(clk), .A(\g.we_clk [17104]));
Q_ASSIGN U15671 ( .B(clk), .A(\g.we_clk [17103]));
Q_ASSIGN U15672 ( .B(clk), .A(\g.we_clk [17102]));
Q_ASSIGN U15673 ( .B(clk), .A(\g.we_clk [17101]));
Q_ASSIGN U15674 ( .B(clk), .A(\g.we_clk [17100]));
Q_ASSIGN U15675 ( .B(clk), .A(\g.we_clk [17099]));
Q_ASSIGN U15676 ( .B(clk), .A(\g.we_clk [17098]));
Q_ASSIGN U15677 ( .B(clk), .A(\g.we_clk [17097]));
Q_ASSIGN U15678 ( .B(clk), .A(\g.we_clk [17096]));
Q_ASSIGN U15679 ( .B(clk), .A(\g.we_clk [17095]));
Q_ASSIGN U15680 ( .B(clk), .A(\g.we_clk [17094]));
Q_ASSIGN U15681 ( .B(clk), .A(\g.we_clk [17093]));
Q_ASSIGN U15682 ( .B(clk), .A(\g.we_clk [17092]));
Q_ASSIGN U15683 ( .B(clk), .A(\g.we_clk [17091]));
Q_ASSIGN U15684 ( .B(clk), .A(\g.we_clk [17090]));
Q_ASSIGN U15685 ( .B(clk), .A(\g.we_clk [17089]));
Q_ASSIGN U15686 ( .B(clk), .A(\g.we_clk [17088]));
Q_ASSIGN U15687 ( .B(clk), .A(\g.we_clk [17087]));
Q_ASSIGN U15688 ( .B(clk), .A(\g.we_clk [17086]));
Q_ASSIGN U15689 ( .B(clk), .A(\g.we_clk [17085]));
Q_ASSIGN U15690 ( .B(clk), .A(\g.we_clk [17084]));
Q_ASSIGN U15691 ( .B(clk), .A(\g.we_clk [17083]));
Q_ASSIGN U15692 ( .B(clk), .A(\g.we_clk [17082]));
Q_ASSIGN U15693 ( .B(clk), .A(\g.we_clk [17081]));
Q_ASSIGN U15694 ( .B(clk), .A(\g.we_clk [17080]));
Q_ASSIGN U15695 ( .B(clk), .A(\g.we_clk [17079]));
Q_ASSIGN U15696 ( .B(clk), .A(\g.we_clk [17078]));
Q_ASSIGN U15697 ( .B(clk), .A(\g.we_clk [17077]));
Q_ASSIGN U15698 ( .B(clk), .A(\g.we_clk [17076]));
Q_ASSIGN U15699 ( .B(clk), .A(\g.we_clk [17075]));
Q_ASSIGN U15700 ( .B(clk), .A(\g.we_clk [17074]));
Q_ASSIGN U15701 ( .B(clk), .A(\g.we_clk [17073]));
Q_ASSIGN U15702 ( .B(clk), .A(\g.we_clk [17072]));
Q_ASSIGN U15703 ( .B(clk), .A(\g.we_clk [17071]));
Q_ASSIGN U15704 ( .B(clk), .A(\g.we_clk [17070]));
Q_ASSIGN U15705 ( .B(clk), .A(\g.we_clk [17069]));
Q_ASSIGN U15706 ( .B(clk), .A(\g.we_clk [17068]));
Q_ASSIGN U15707 ( .B(clk), .A(\g.we_clk [17067]));
Q_ASSIGN U15708 ( .B(clk), .A(\g.we_clk [17066]));
Q_ASSIGN U15709 ( .B(clk), .A(\g.we_clk [17065]));
Q_ASSIGN U15710 ( .B(clk), .A(\g.we_clk [17064]));
Q_ASSIGN U15711 ( .B(clk), .A(\g.we_clk [17063]));
Q_ASSIGN U15712 ( .B(clk), .A(\g.we_clk [17062]));
Q_ASSIGN U15713 ( .B(clk), .A(\g.we_clk [17061]));
Q_ASSIGN U15714 ( .B(clk), .A(\g.we_clk [17060]));
Q_ASSIGN U15715 ( .B(clk), .A(\g.we_clk [17059]));
Q_ASSIGN U15716 ( .B(clk), .A(\g.we_clk [17058]));
Q_ASSIGN U15717 ( .B(clk), .A(\g.we_clk [17057]));
Q_ASSIGN U15718 ( .B(clk), .A(\g.we_clk [17056]));
Q_ASSIGN U15719 ( .B(clk), .A(\g.we_clk [17055]));
Q_ASSIGN U15720 ( .B(clk), .A(\g.we_clk [17054]));
Q_ASSIGN U15721 ( .B(clk), .A(\g.we_clk [17053]));
Q_ASSIGN U15722 ( .B(clk), .A(\g.we_clk [17052]));
Q_ASSIGN U15723 ( .B(clk), .A(\g.we_clk [17051]));
Q_ASSIGN U15724 ( .B(clk), .A(\g.we_clk [17050]));
Q_ASSIGN U15725 ( .B(clk), .A(\g.we_clk [17049]));
Q_ASSIGN U15726 ( .B(clk), .A(\g.we_clk [17048]));
Q_ASSIGN U15727 ( .B(clk), .A(\g.we_clk [17047]));
Q_ASSIGN U15728 ( .B(clk), .A(\g.we_clk [17046]));
Q_ASSIGN U15729 ( .B(clk), .A(\g.we_clk [17045]));
Q_ASSIGN U15730 ( .B(clk), .A(\g.we_clk [17044]));
Q_ASSIGN U15731 ( .B(clk), .A(\g.we_clk [17043]));
Q_ASSIGN U15732 ( .B(clk), .A(\g.we_clk [17042]));
Q_ASSIGN U15733 ( .B(clk), .A(\g.we_clk [17041]));
Q_ASSIGN U15734 ( .B(clk), .A(\g.we_clk [17040]));
Q_ASSIGN U15735 ( .B(clk), .A(\g.we_clk [17039]));
Q_ASSIGN U15736 ( .B(clk), .A(\g.we_clk [17038]));
Q_ASSIGN U15737 ( .B(clk), .A(\g.we_clk [17037]));
Q_ASSIGN U15738 ( .B(clk), .A(\g.we_clk [17036]));
Q_ASSIGN U15739 ( .B(clk), .A(\g.we_clk [17035]));
Q_ASSIGN U15740 ( .B(clk), .A(\g.we_clk [17034]));
Q_ASSIGN U15741 ( .B(clk), .A(\g.we_clk [17033]));
Q_ASSIGN U15742 ( .B(clk), .A(\g.we_clk [17032]));
Q_ASSIGN U15743 ( .B(clk), .A(\g.we_clk [17031]));
Q_ASSIGN U15744 ( .B(clk), .A(\g.we_clk [17030]));
Q_ASSIGN U15745 ( .B(clk), .A(\g.we_clk [17029]));
Q_ASSIGN U15746 ( .B(clk), .A(\g.we_clk [17028]));
Q_ASSIGN U15747 ( .B(clk), .A(\g.we_clk [17027]));
Q_ASSIGN U15748 ( .B(clk), .A(\g.we_clk [17026]));
Q_ASSIGN U15749 ( .B(clk), .A(\g.we_clk [17025]));
Q_ASSIGN U15750 ( .B(clk), .A(\g.we_clk [17024]));
Q_ASSIGN U15751 ( .B(clk), .A(\g.we_clk [17023]));
Q_ASSIGN U15752 ( .B(clk), .A(\g.we_clk [17022]));
Q_ASSIGN U15753 ( .B(clk), .A(\g.we_clk [17021]));
Q_ASSIGN U15754 ( .B(clk), .A(\g.we_clk [17020]));
Q_ASSIGN U15755 ( .B(clk), .A(\g.we_clk [17019]));
Q_ASSIGN U15756 ( .B(clk), .A(\g.we_clk [17018]));
Q_ASSIGN U15757 ( .B(clk), .A(\g.we_clk [17017]));
Q_ASSIGN U15758 ( .B(clk), .A(\g.we_clk [17016]));
Q_ASSIGN U15759 ( .B(clk), .A(\g.we_clk [17015]));
Q_ASSIGN U15760 ( .B(clk), .A(\g.we_clk [17014]));
Q_ASSIGN U15761 ( .B(clk), .A(\g.we_clk [17013]));
Q_ASSIGN U15762 ( .B(clk), .A(\g.we_clk [17012]));
Q_ASSIGN U15763 ( .B(clk), .A(\g.we_clk [17011]));
Q_ASSIGN U15764 ( .B(clk), .A(\g.we_clk [17010]));
Q_ASSIGN U15765 ( .B(clk), .A(\g.we_clk [17009]));
Q_ASSIGN U15766 ( .B(clk), .A(\g.we_clk [17008]));
Q_ASSIGN U15767 ( .B(clk), .A(\g.we_clk [17007]));
Q_ASSIGN U15768 ( .B(clk), .A(\g.we_clk [17006]));
Q_ASSIGN U15769 ( .B(clk), .A(\g.we_clk [17005]));
Q_ASSIGN U15770 ( .B(clk), .A(\g.we_clk [17004]));
Q_ASSIGN U15771 ( .B(clk), .A(\g.we_clk [17003]));
Q_ASSIGN U15772 ( .B(clk), .A(\g.we_clk [17002]));
Q_ASSIGN U15773 ( .B(clk), .A(\g.we_clk [17001]));
Q_ASSIGN U15774 ( .B(clk), .A(\g.we_clk [17000]));
Q_ASSIGN U15775 ( .B(clk), .A(\g.we_clk [16999]));
Q_ASSIGN U15776 ( .B(clk), .A(\g.we_clk [16998]));
Q_ASSIGN U15777 ( .B(clk), .A(\g.we_clk [16997]));
Q_ASSIGN U15778 ( .B(clk), .A(\g.we_clk [16996]));
Q_ASSIGN U15779 ( .B(clk), .A(\g.we_clk [16995]));
Q_ASSIGN U15780 ( .B(clk), .A(\g.we_clk [16994]));
Q_ASSIGN U15781 ( .B(clk), .A(\g.we_clk [16993]));
Q_ASSIGN U15782 ( .B(clk), .A(\g.we_clk [16992]));
Q_ASSIGN U15783 ( .B(clk), .A(\g.we_clk [16991]));
Q_ASSIGN U15784 ( .B(clk), .A(\g.we_clk [16990]));
Q_ASSIGN U15785 ( .B(clk), .A(\g.we_clk [16989]));
Q_ASSIGN U15786 ( .B(clk), .A(\g.we_clk [16988]));
Q_ASSIGN U15787 ( .B(clk), .A(\g.we_clk [16987]));
Q_ASSIGN U15788 ( .B(clk), .A(\g.we_clk [16986]));
Q_ASSIGN U15789 ( .B(clk), .A(\g.we_clk [16985]));
Q_ASSIGN U15790 ( .B(clk), .A(\g.we_clk [16984]));
Q_ASSIGN U15791 ( .B(clk), .A(\g.we_clk [16983]));
Q_ASSIGN U15792 ( .B(clk), .A(\g.we_clk [16982]));
Q_ASSIGN U15793 ( .B(clk), .A(\g.we_clk [16981]));
Q_ASSIGN U15794 ( .B(clk), .A(\g.we_clk [16980]));
Q_ASSIGN U15795 ( .B(clk), .A(\g.we_clk [16979]));
Q_ASSIGN U15796 ( .B(clk), .A(\g.we_clk [16978]));
Q_ASSIGN U15797 ( .B(clk), .A(\g.we_clk [16977]));
Q_ASSIGN U15798 ( .B(clk), .A(\g.we_clk [16976]));
Q_ASSIGN U15799 ( .B(clk), .A(\g.we_clk [16975]));
Q_ASSIGN U15800 ( .B(clk), .A(\g.we_clk [16974]));
Q_ASSIGN U15801 ( .B(clk), .A(\g.we_clk [16973]));
Q_ASSIGN U15802 ( .B(clk), .A(\g.we_clk [16972]));
Q_ASSIGN U15803 ( .B(clk), .A(\g.we_clk [16971]));
Q_ASSIGN U15804 ( .B(clk), .A(\g.we_clk [16970]));
Q_ASSIGN U15805 ( .B(clk), .A(\g.we_clk [16969]));
Q_ASSIGN U15806 ( .B(clk), .A(\g.we_clk [16968]));
Q_ASSIGN U15807 ( .B(clk), .A(\g.we_clk [16967]));
Q_ASSIGN U15808 ( .B(clk), .A(\g.we_clk [16966]));
Q_ASSIGN U15809 ( .B(clk), .A(\g.we_clk [16965]));
Q_ASSIGN U15810 ( .B(clk), .A(\g.we_clk [16964]));
Q_ASSIGN U15811 ( .B(clk), .A(\g.we_clk [16963]));
Q_ASSIGN U15812 ( .B(clk), .A(\g.we_clk [16962]));
Q_ASSIGN U15813 ( .B(clk), .A(\g.we_clk [16961]));
Q_ASSIGN U15814 ( .B(clk), .A(\g.we_clk [16960]));
Q_ASSIGN U15815 ( .B(clk), .A(\g.we_clk [16959]));
Q_ASSIGN U15816 ( .B(clk), .A(\g.we_clk [16958]));
Q_ASSIGN U15817 ( .B(clk), .A(\g.we_clk [16957]));
Q_ASSIGN U15818 ( .B(clk), .A(\g.we_clk [16956]));
Q_ASSIGN U15819 ( .B(clk), .A(\g.we_clk [16955]));
Q_ASSIGN U15820 ( .B(clk), .A(\g.we_clk [16954]));
Q_ASSIGN U15821 ( .B(clk), .A(\g.we_clk [16953]));
Q_ASSIGN U15822 ( .B(clk), .A(\g.we_clk [16952]));
Q_ASSIGN U15823 ( .B(clk), .A(\g.we_clk [16951]));
Q_ASSIGN U15824 ( .B(clk), .A(\g.we_clk [16950]));
Q_ASSIGN U15825 ( .B(clk), .A(\g.we_clk [16949]));
Q_ASSIGN U15826 ( .B(clk), .A(\g.we_clk [16948]));
Q_ASSIGN U15827 ( .B(clk), .A(\g.we_clk [16947]));
Q_ASSIGN U15828 ( .B(clk), .A(\g.we_clk [16946]));
Q_ASSIGN U15829 ( .B(clk), .A(\g.we_clk [16945]));
Q_ASSIGN U15830 ( .B(clk), .A(\g.we_clk [16944]));
Q_ASSIGN U15831 ( .B(clk), .A(\g.we_clk [16943]));
Q_ASSIGN U15832 ( .B(clk), .A(\g.we_clk [16942]));
Q_ASSIGN U15833 ( .B(clk), .A(\g.we_clk [16941]));
Q_ASSIGN U15834 ( .B(clk), .A(\g.we_clk [16940]));
Q_ASSIGN U15835 ( .B(clk), .A(\g.we_clk [16939]));
Q_ASSIGN U15836 ( .B(clk), .A(\g.we_clk [16938]));
Q_ASSIGN U15837 ( .B(clk), .A(\g.we_clk [16937]));
Q_ASSIGN U15838 ( .B(clk), .A(\g.we_clk [16936]));
Q_ASSIGN U15839 ( .B(clk), .A(\g.we_clk [16935]));
Q_ASSIGN U15840 ( .B(clk), .A(\g.we_clk [16934]));
Q_ASSIGN U15841 ( .B(clk), .A(\g.we_clk [16933]));
Q_ASSIGN U15842 ( .B(clk), .A(\g.we_clk [16932]));
Q_ASSIGN U15843 ( .B(clk), .A(\g.we_clk [16931]));
Q_ASSIGN U15844 ( .B(clk), .A(\g.we_clk [16930]));
Q_ASSIGN U15845 ( .B(clk), .A(\g.we_clk [16929]));
Q_ASSIGN U15846 ( .B(clk), .A(\g.we_clk [16928]));
Q_ASSIGN U15847 ( .B(clk), .A(\g.we_clk [16927]));
Q_ASSIGN U15848 ( .B(clk), .A(\g.we_clk [16926]));
Q_ASSIGN U15849 ( .B(clk), .A(\g.we_clk [16925]));
Q_ASSIGN U15850 ( .B(clk), .A(\g.we_clk [16924]));
Q_ASSIGN U15851 ( .B(clk), .A(\g.we_clk [16923]));
Q_ASSIGN U15852 ( .B(clk), .A(\g.we_clk [16922]));
Q_ASSIGN U15853 ( .B(clk), .A(\g.we_clk [16921]));
Q_ASSIGN U15854 ( .B(clk), .A(\g.we_clk [16920]));
Q_ASSIGN U15855 ( .B(clk), .A(\g.we_clk [16919]));
Q_ASSIGN U15856 ( .B(clk), .A(\g.we_clk [16918]));
Q_ASSIGN U15857 ( .B(clk), .A(\g.we_clk [16917]));
Q_ASSIGN U15858 ( .B(clk), .A(\g.we_clk [16916]));
Q_ASSIGN U15859 ( .B(clk), .A(\g.we_clk [16915]));
Q_ASSIGN U15860 ( .B(clk), .A(\g.we_clk [16914]));
Q_ASSIGN U15861 ( .B(clk), .A(\g.we_clk [16913]));
Q_ASSIGN U15862 ( .B(clk), .A(\g.we_clk [16912]));
Q_ASSIGN U15863 ( .B(clk), .A(\g.we_clk [16911]));
Q_ASSIGN U15864 ( .B(clk), .A(\g.we_clk [16910]));
Q_ASSIGN U15865 ( .B(clk), .A(\g.we_clk [16909]));
Q_ASSIGN U15866 ( .B(clk), .A(\g.we_clk [16908]));
Q_ASSIGN U15867 ( .B(clk), .A(\g.we_clk [16907]));
Q_ASSIGN U15868 ( .B(clk), .A(\g.we_clk [16906]));
Q_ASSIGN U15869 ( .B(clk), .A(\g.we_clk [16905]));
Q_ASSIGN U15870 ( .B(clk), .A(\g.we_clk [16904]));
Q_ASSIGN U15871 ( .B(clk), .A(\g.we_clk [16903]));
Q_ASSIGN U15872 ( .B(clk), .A(\g.we_clk [16902]));
Q_ASSIGN U15873 ( .B(clk), .A(\g.we_clk [16901]));
Q_ASSIGN U15874 ( .B(clk), .A(\g.we_clk [16900]));
Q_ASSIGN U15875 ( .B(clk), .A(\g.we_clk [16899]));
Q_ASSIGN U15876 ( .B(clk), .A(\g.we_clk [16898]));
Q_ASSIGN U15877 ( .B(clk), .A(\g.we_clk [16897]));
Q_ASSIGN U15878 ( .B(clk), .A(\g.we_clk [16896]));
Q_ASSIGN U15879 ( .B(clk), .A(\g.we_clk [16895]));
Q_ASSIGN U15880 ( .B(clk), .A(\g.we_clk [16894]));
Q_ASSIGN U15881 ( .B(clk), .A(\g.we_clk [16893]));
Q_ASSIGN U15882 ( .B(clk), .A(\g.we_clk [16892]));
Q_ASSIGN U15883 ( .B(clk), .A(\g.we_clk [16891]));
Q_ASSIGN U15884 ( .B(clk), .A(\g.we_clk [16890]));
Q_ASSIGN U15885 ( .B(clk), .A(\g.we_clk [16889]));
Q_ASSIGN U15886 ( .B(clk), .A(\g.we_clk [16888]));
Q_ASSIGN U15887 ( .B(clk), .A(\g.we_clk [16887]));
Q_ASSIGN U15888 ( .B(clk), .A(\g.we_clk [16886]));
Q_ASSIGN U15889 ( .B(clk), .A(\g.we_clk [16885]));
Q_ASSIGN U15890 ( .B(clk), .A(\g.we_clk [16884]));
Q_ASSIGN U15891 ( .B(clk), .A(\g.we_clk [16883]));
Q_ASSIGN U15892 ( .B(clk), .A(\g.we_clk [16882]));
Q_ASSIGN U15893 ( .B(clk), .A(\g.we_clk [16881]));
Q_ASSIGN U15894 ( .B(clk), .A(\g.we_clk [16880]));
Q_ASSIGN U15895 ( .B(clk), .A(\g.we_clk [16879]));
Q_ASSIGN U15896 ( .B(clk), .A(\g.we_clk [16878]));
Q_ASSIGN U15897 ( .B(clk), .A(\g.we_clk [16877]));
Q_ASSIGN U15898 ( .B(clk), .A(\g.we_clk [16876]));
Q_ASSIGN U15899 ( .B(clk), .A(\g.we_clk [16875]));
Q_ASSIGN U15900 ( .B(clk), .A(\g.we_clk [16874]));
Q_ASSIGN U15901 ( .B(clk), .A(\g.we_clk [16873]));
Q_ASSIGN U15902 ( .B(clk), .A(\g.we_clk [16872]));
Q_ASSIGN U15903 ( .B(clk), .A(\g.we_clk [16871]));
Q_ASSIGN U15904 ( .B(clk), .A(\g.we_clk [16870]));
Q_ASSIGN U15905 ( .B(clk), .A(\g.we_clk [16869]));
Q_ASSIGN U15906 ( .B(clk), .A(\g.we_clk [16868]));
Q_ASSIGN U15907 ( .B(clk), .A(\g.we_clk [16867]));
Q_ASSIGN U15908 ( .B(clk), .A(\g.we_clk [16866]));
Q_ASSIGN U15909 ( .B(clk), .A(\g.we_clk [16865]));
Q_ASSIGN U15910 ( .B(clk), .A(\g.we_clk [16864]));
Q_ASSIGN U15911 ( .B(clk), .A(\g.we_clk [16863]));
Q_ASSIGN U15912 ( .B(clk), .A(\g.we_clk [16862]));
Q_ASSIGN U15913 ( .B(clk), .A(\g.we_clk [16861]));
Q_ASSIGN U15914 ( .B(clk), .A(\g.we_clk [16860]));
Q_ASSIGN U15915 ( .B(clk), .A(\g.we_clk [16859]));
Q_ASSIGN U15916 ( .B(clk), .A(\g.we_clk [16858]));
Q_ASSIGN U15917 ( .B(clk), .A(\g.we_clk [16857]));
Q_ASSIGN U15918 ( .B(clk), .A(\g.we_clk [16856]));
Q_ASSIGN U15919 ( .B(clk), .A(\g.we_clk [16855]));
Q_ASSIGN U15920 ( .B(clk), .A(\g.we_clk [16854]));
Q_ASSIGN U15921 ( .B(clk), .A(\g.we_clk [16853]));
Q_ASSIGN U15922 ( .B(clk), .A(\g.we_clk [16852]));
Q_ASSIGN U15923 ( .B(clk), .A(\g.we_clk [16851]));
Q_ASSIGN U15924 ( .B(clk), .A(\g.we_clk [16850]));
Q_ASSIGN U15925 ( .B(clk), .A(\g.we_clk [16849]));
Q_ASSIGN U15926 ( .B(clk), .A(\g.we_clk [16848]));
Q_ASSIGN U15927 ( .B(clk), .A(\g.we_clk [16847]));
Q_ASSIGN U15928 ( .B(clk), .A(\g.we_clk [16846]));
Q_ASSIGN U15929 ( .B(clk), .A(\g.we_clk [16845]));
Q_ASSIGN U15930 ( .B(clk), .A(\g.we_clk [16844]));
Q_ASSIGN U15931 ( .B(clk), .A(\g.we_clk [16843]));
Q_ASSIGN U15932 ( .B(clk), .A(\g.we_clk [16842]));
Q_ASSIGN U15933 ( .B(clk), .A(\g.we_clk [16841]));
Q_ASSIGN U15934 ( .B(clk), .A(\g.we_clk [16840]));
Q_ASSIGN U15935 ( .B(clk), .A(\g.we_clk [16839]));
Q_ASSIGN U15936 ( .B(clk), .A(\g.we_clk [16838]));
Q_ASSIGN U15937 ( .B(clk), .A(\g.we_clk [16837]));
Q_ASSIGN U15938 ( .B(clk), .A(\g.we_clk [16836]));
Q_ASSIGN U15939 ( .B(clk), .A(\g.we_clk [16835]));
Q_ASSIGN U15940 ( .B(clk), .A(\g.we_clk [16834]));
Q_ASSIGN U15941 ( .B(clk), .A(\g.we_clk [16833]));
Q_ASSIGN U15942 ( .B(clk), .A(\g.we_clk [16832]));
Q_ASSIGN U15943 ( .B(clk), .A(\g.we_clk [16831]));
Q_ASSIGN U15944 ( .B(clk), .A(\g.we_clk [16830]));
Q_ASSIGN U15945 ( .B(clk), .A(\g.we_clk [16829]));
Q_ASSIGN U15946 ( .B(clk), .A(\g.we_clk [16828]));
Q_ASSIGN U15947 ( .B(clk), .A(\g.we_clk [16827]));
Q_ASSIGN U15948 ( .B(clk), .A(\g.we_clk [16826]));
Q_ASSIGN U15949 ( .B(clk), .A(\g.we_clk [16825]));
Q_ASSIGN U15950 ( .B(clk), .A(\g.we_clk [16824]));
Q_ASSIGN U15951 ( .B(clk), .A(\g.we_clk [16823]));
Q_ASSIGN U15952 ( .B(clk), .A(\g.we_clk [16822]));
Q_ASSIGN U15953 ( .B(clk), .A(\g.we_clk [16821]));
Q_ASSIGN U15954 ( .B(clk), .A(\g.we_clk [16820]));
Q_ASSIGN U15955 ( .B(clk), .A(\g.we_clk [16819]));
Q_ASSIGN U15956 ( .B(clk), .A(\g.we_clk [16818]));
Q_ASSIGN U15957 ( .B(clk), .A(\g.we_clk [16817]));
Q_ASSIGN U15958 ( .B(clk), .A(\g.we_clk [16816]));
Q_ASSIGN U15959 ( .B(clk), .A(\g.we_clk [16815]));
Q_ASSIGN U15960 ( .B(clk), .A(\g.we_clk [16814]));
Q_ASSIGN U15961 ( .B(clk), .A(\g.we_clk [16813]));
Q_ASSIGN U15962 ( .B(clk), .A(\g.we_clk [16812]));
Q_ASSIGN U15963 ( .B(clk), .A(\g.we_clk [16811]));
Q_ASSIGN U15964 ( .B(clk), .A(\g.we_clk [16810]));
Q_ASSIGN U15965 ( .B(clk), .A(\g.we_clk [16809]));
Q_ASSIGN U15966 ( .B(clk), .A(\g.we_clk [16808]));
Q_ASSIGN U15967 ( .B(clk), .A(\g.we_clk [16807]));
Q_ASSIGN U15968 ( .B(clk), .A(\g.we_clk [16806]));
Q_ASSIGN U15969 ( .B(clk), .A(\g.we_clk [16805]));
Q_ASSIGN U15970 ( .B(clk), .A(\g.we_clk [16804]));
Q_ASSIGN U15971 ( .B(clk), .A(\g.we_clk [16803]));
Q_ASSIGN U15972 ( .B(clk), .A(\g.we_clk [16802]));
Q_ASSIGN U15973 ( .B(clk), .A(\g.we_clk [16801]));
Q_ASSIGN U15974 ( .B(clk), .A(\g.we_clk [16800]));
Q_ASSIGN U15975 ( .B(clk), .A(\g.we_clk [16799]));
Q_ASSIGN U15976 ( .B(clk), .A(\g.we_clk [16798]));
Q_ASSIGN U15977 ( .B(clk), .A(\g.we_clk [16797]));
Q_ASSIGN U15978 ( .B(clk), .A(\g.we_clk [16796]));
Q_ASSIGN U15979 ( .B(clk), .A(\g.we_clk [16795]));
Q_ASSIGN U15980 ( .B(clk), .A(\g.we_clk [16794]));
Q_ASSIGN U15981 ( .B(clk), .A(\g.we_clk [16793]));
Q_ASSIGN U15982 ( .B(clk), .A(\g.we_clk [16792]));
Q_ASSIGN U15983 ( .B(clk), .A(\g.we_clk [16791]));
Q_ASSIGN U15984 ( .B(clk), .A(\g.we_clk [16790]));
Q_ASSIGN U15985 ( .B(clk), .A(\g.we_clk [16789]));
Q_ASSIGN U15986 ( .B(clk), .A(\g.we_clk [16788]));
Q_ASSIGN U15987 ( .B(clk), .A(\g.we_clk [16787]));
Q_ASSIGN U15988 ( .B(clk), .A(\g.we_clk [16786]));
Q_ASSIGN U15989 ( .B(clk), .A(\g.we_clk [16785]));
Q_ASSIGN U15990 ( .B(clk), .A(\g.we_clk [16784]));
Q_ASSIGN U15991 ( .B(clk), .A(\g.we_clk [16783]));
Q_ASSIGN U15992 ( .B(clk), .A(\g.we_clk [16782]));
Q_ASSIGN U15993 ( .B(clk), .A(\g.we_clk [16781]));
Q_ASSIGN U15994 ( .B(clk), .A(\g.we_clk [16780]));
Q_ASSIGN U15995 ( .B(clk), .A(\g.we_clk [16779]));
Q_ASSIGN U15996 ( .B(clk), .A(\g.we_clk [16778]));
Q_ASSIGN U15997 ( .B(clk), .A(\g.we_clk [16777]));
Q_ASSIGN U15998 ( .B(clk), .A(\g.we_clk [16776]));
Q_ASSIGN U15999 ( .B(clk), .A(\g.we_clk [16775]));
Q_ASSIGN U16000 ( .B(clk), .A(\g.we_clk [16774]));
Q_ASSIGN U16001 ( .B(clk), .A(\g.we_clk [16773]));
Q_ASSIGN U16002 ( .B(clk), .A(\g.we_clk [16772]));
Q_ASSIGN U16003 ( .B(clk), .A(\g.we_clk [16771]));
Q_ASSIGN U16004 ( .B(clk), .A(\g.we_clk [16770]));
Q_ASSIGN U16005 ( .B(clk), .A(\g.we_clk [16769]));
Q_ASSIGN U16006 ( .B(clk), .A(\g.we_clk [16768]));
Q_ASSIGN U16007 ( .B(clk), .A(\g.we_clk [16767]));
Q_ASSIGN U16008 ( .B(clk), .A(\g.we_clk [16766]));
Q_ASSIGN U16009 ( .B(clk), .A(\g.we_clk [16765]));
Q_ASSIGN U16010 ( .B(clk), .A(\g.we_clk [16764]));
Q_ASSIGN U16011 ( .B(clk), .A(\g.we_clk [16763]));
Q_ASSIGN U16012 ( .B(clk), .A(\g.we_clk [16762]));
Q_ASSIGN U16013 ( .B(clk), .A(\g.we_clk [16761]));
Q_ASSIGN U16014 ( .B(clk), .A(\g.we_clk [16760]));
Q_ASSIGN U16015 ( .B(clk), .A(\g.we_clk [16759]));
Q_ASSIGN U16016 ( .B(clk), .A(\g.we_clk [16758]));
Q_ASSIGN U16017 ( .B(clk), .A(\g.we_clk [16757]));
Q_ASSIGN U16018 ( .B(clk), .A(\g.we_clk [16756]));
Q_ASSIGN U16019 ( .B(clk), .A(\g.we_clk [16755]));
Q_ASSIGN U16020 ( .B(clk), .A(\g.we_clk [16754]));
Q_ASSIGN U16021 ( .B(clk), .A(\g.we_clk [16753]));
Q_ASSIGN U16022 ( .B(clk), .A(\g.we_clk [16752]));
Q_ASSIGN U16023 ( .B(clk), .A(\g.we_clk [16751]));
Q_ASSIGN U16024 ( .B(clk), .A(\g.we_clk [16750]));
Q_ASSIGN U16025 ( .B(clk), .A(\g.we_clk [16749]));
Q_ASSIGN U16026 ( .B(clk), .A(\g.we_clk [16748]));
Q_ASSIGN U16027 ( .B(clk), .A(\g.we_clk [16747]));
Q_ASSIGN U16028 ( .B(clk), .A(\g.we_clk [16746]));
Q_ASSIGN U16029 ( .B(clk), .A(\g.we_clk [16745]));
Q_ASSIGN U16030 ( .B(clk), .A(\g.we_clk [16744]));
Q_ASSIGN U16031 ( .B(clk), .A(\g.we_clk [16743]));
Q_ASSIGN U16032 ( .B(clk), .A(\g.we_clk [16742]));
Q_ASSIGN U16033 ( .B(clk), .A(\g.we_clk [16741]));
Q_ASSIGN U16034 ( .B(clk), .A(\g.we_clk [16740]));
Q_ASSIGN U16035 ( .B(clk), .A(\g.we_clk [16739]));
Q_ASSIGN U16036 ( .B(clk), .A(\g.we_clk [16738]));
Q_ASSIGN U16037 ( .B(clk), .A(\g.we_clk [16737]));
Q_ASSIGN U16038 ( .B(clk), .A(\g.we_clk [16736]));
Q_ASSIGN U16039 ( .B(clk), .A(\g.we_clk [16735]));
Q_ASSIGN U16040 ( .B(clk), .A(\g.we_clk [16734]));
Q_ASSIGN U16041 ( .B(clk), .A(\g.we_clk [16733]));
Q_ASSIGN U16042 ( .B(clk), .A(\g.we_clk [16732]));
Q_ASSIGN U16043 ( .B(clk), .A(\g.we_clk [16731]));
Q_ASSIGN U16044 ( .B(clk), .A(\g.we_clk [16730]));
Q_ASSIGN U16045 ( .B(clk), .A(\g.we_clk [16729]));
Q_ASSIGN U16046 ( .B(clk), .A(\g.we_clk [16728]));
Q_ASSIGN U16047 ( .B(clk), .A(\g.we_clk [16727]));
Q_ASSIGN U16048 ( .B(clk), .A(\g.we_clk [16726]));
Q_ASSIGN U16049 ( .B(clk), .A(\g.we_clk [16725]));
Q_ASSIGN U16050 ( .B(clk), .A(\g.we_clk [16724]));
Q_ASSIGN U16051 ( .B(clk), .A(\g.we_clk [16723]));
Q_ASSIGN U16052 ( .B(clk), .A(\g.we_clk [16722]));
Q_ASSIGN U16053 ( .B(clk), .A(\g.we_clk [16721]));
Q_ASSIGN U16054 ( .B(clk), .A(\g.we_clk [16720]));
Q_ASSIGN U16055 ( .B(clk), .A(\g.we_clk [16719]));
Q_ASSIGN U16056 ( .B(clk), .A(\g.we_clk [16718]));
Q_ASSIGN U16057 ( .B(clk), .A(\g.we_clk [16717]));
Q_ASSIGN U16058 ( .B(clk), .A(\g.we_clk [16716]));
Q_ASSIGN U16059 ( .B(clk), .A(\g.we_clk [16715]));
Q_ASSIGN U16060 ( .B(clk), .A(\g.we_clk [16714]));
Q_ASSIGN U16061 ( .B(clk), .A(\g.we_clk [16713]));
Q_ASSIGN U16062 ( .B(clk), .A(\g.we_clk [16712]));
Q_ASSIGN U16063 ( .B(clk), .A(\g.we_clk [16711]));
Q_ASSIGN U16064 ( .B(clk), .A(\g.we_clk [16710]));
Q_ASSIGN U16065 ( .B(clk), .A(\g.we_clk [16709]));
Q_ASSIGN U16066 ( .B(clk), .A(\g.we_clk [16708]));
Q_ASSIGN U16067 ( .B(clk), .A(\g.we_clk [16707]));
Q_ASSIGN U16068 ( .B(clk), .A(\g.we_clk [16706]));
Q_ASSIGN U16069 ( .B(clk), .A(\g.we_clk [16705]));
Q_ASSIGN U16070 ( .B(clk), .A(\g.we_clk [16704]));
Q_ASSIGN U16071 ( .B(clk), .A(\g.we_clk [16703]));
Q_ASSIGN U16072 ( .B(clk), .A(\g.we_clk [16702]));
Q_ASSIGN U16073 ( .B(clk), .A(\g.we_clk [16701]));
Q_ASSIGN U16074 ( .B(clk), .A(\g.we_clk [16700]));
Q_ASSIGN U16075 ( .B(clk), .A(\g.we_clk [16699]));
Q_ASSIGN U16076 ( .B(clk), .A(\g.we_clk [16698]));
Q_ASSIGN U16077 ( .B(clk), .A(\g.we_clk [16697]));
Q_ASSIGN U16078 ( .B(clk), .A(\g.we_clk [16696]));
Q_ASSIGN U16079 ( .B(clk), .A(\g.we_clk [16695]));
Q_ASSIGN U16080 ( .B(clk), .A(\g.we_clk [16694]));
Q_ASSIGN U16081 ( .B(clk), .A(\g.we_clk [16693]));
Q_ASSIGN U16082 ( .B(clk), .A(\g.we_clk [16692]));
Q_ASSIGN U16083 ( .B(clk), .A(\g.we_clk [16691]));
Q_ASSIGN U16084 ( .B(clk), .A(\g.we_clk [16690]));
Q_ASSIGN U16085 ( .B(clk), .A(\g.we_clk [16689]));
Q_ASSIGN U16086 ( .B(clk), .A(\g.we_clk [16688]));
Q_ASSIGN U16087 ( .B(clk), .A(\g.we_clk [16687]));
Q_ASSIGN U16088 ( .B(clk), .A(\g.we_clk [16686]));
Q_ASSIGN U16089 ( .B(clk), .A(\g.we_clk [16685]));
Q_ASSIGN U16090 ( .B(clk), .A(\g.we_clk [16684]));
Q_ASSIGN U16091 ( .B(clk), .A(\g.we_clk [16683]));
Q_ASSIGN U16092 ( .B(clk), .A(\g.we_clk [16682]));
Q_ASSIGN U16093 ( .B(clk), .A(\g.we_clk [16681]));
Q_ASSIGN U16094 ( .B(clk), .A(\g.we_clk [16680]));
Q_ASSIGN U16095 ( .B(clk), .A(\g.we_clk [16679]));
Q_ASSIGN U16096 ( .B(clk), .A(\g.we_clk [16678]));
Q_ASSIGN U16097 ( .B(clk), .A(\g.we_clk [16677]));
Q_ASSIGN U16098 ( .B(clk), .A(\g.we_clk [16676]));
Q_ASSIGN U16099 ( .B(clk), .A(\g.we_clk [16675]));
Q_ASSIGN U16100 ( .B(clk), .A(\g.we_clk [16674]));
Q_ASSIGN U16101 ( .B(clk), .A(\g.we_clk [16673]));
Q_ASSIGN U16102 ( .B(clk), .A(\g.we_clk [16672]));
Q_ASSIGN U16103 ( .B(clk), .A(\g.we_clk [16671]));
Q_ASSIGN U16104 ( .B(clk), .A(\g.we_clk [16670]));
Q_ASSIGN U16105 ( .B(clk), .A(\g.we_clk [16669]));
Q_ASSIGN U16106 ( .B(clk), .A(\g.we_clk [16668]));
Q_ASSIGN U16107 ( .B(clk), .A(\g.we_clk [16667]));
Q_ASSIGN U16108 ( .B(clk), .A(\g.we_clk [16666]));
Q_ASSIGN U16109 ( .B(clk), .A(\g.we_clk [16665]));
Q_ASSIGN U16110 ( .B(clk), .A(\g.we_clk [16664]));
Q_ASSIGN U16111 ( .B(clk), .A(\g.we_clk [16663]));
Q_ASSIGN U16112 ( .B(clk), .A(\g.we_clk [16662]));
Q_ASSIGN U16113 ( .B(clk), .A(\g.we_clk [16661]));
Q_ASSIGN U16114 ( .B(clk), .A(\g.we_clk [16660]));
Q_ASSIGN U16115 ( .B(clk), .A(\g.we_clk [16659]));
Q_ASSIGN U16116 ( .B(clk), .A(\g.we_clk [16658]));
Q_ASSIGN U16117 ( .B(clk), .A(\g.we_clk [16657]));
Q_ASSIGN U16118 ( .B(clk), .A(\g.we_clk [16656]));
Q_ASSIGN U16119 ( .B(clk), .A(\g.we_clk [16655]));
Q_ASSIGN U16120 ( .B(clk), .A(\g.we_clk [16654]));
Q_ASSIGN U16121 ( .B(clk), .A(\g.we_clk [16653]));
Q_ASSIGN U16122 ( .B(clk), .A(\g.we_clk [16652]));
Q_ASSIGN U16123 ( .B(clk), .A(\g.we_clk [16651]));
Q_ASSIGN U16124 ( .B(clk), .A(\g.we_clk [16650]));
Q_ASSIGN U16125 ( .B(clk), .A(\g.we_clk [16649]));
Q_ASSIGN U16126 ( .B(clk), .A(\g.we_clk [16648]));
Q_ASSIGN U16127 ( .B(clk), .A(\g.we_clk [16647]));
Q_ASSIGN U16128 ( .B(clk), .A(\g.we_clk [16646]));
Q_ASSIGN U16129 ( .B(clk), .A(\g.we_clk [16645]));
Q_ASSIGN U16130 ( .B(clk), .A(\g.we_clk [16644]));
Q_ASSIGN U16131 ( .B(clk), .A(\g.we_clk [16643]));
Q_ASSIGN U16132 ( .B(clk), .A(\g.we_clk [16642]));
Q_ASSIGN U16133 ( .B(clk), .A(\g.we_clk [16641]));
Q_ASSIGN U16134 ( .B(clk), .A(\g.we_clk [16640]));
Q_ASSIGN U16135 ( .B(clk), .A(\g.we_clk [16639]));
Q_ASSIGN U16136 ( .B(clk), .A(\g.we_clk [16638]));
Q_ASSIGN U16137 ( .B(clk), .A(\g.we_clk [16637]));
Q_ASSIGN U16138 ( .B(clk), .A(\g.we_clk [16636]));
Q_ASSIGN U16139 ( .B(clk), .A(\g.we_clk [16635]));
Q_ASSIGN U16140 ( .B(clk), .A(\g.we_clk [16634]));
Q_ASSIGN U16141 ( .B(clk), .A(\g.we_clk [16633]));
Q_ASSIGN U16142 ( .B(clk), .A(\g.we_clk [16632]));
Q_ASSIGN U16143 ( .B(clk), .A(\g.we_clk [16631]));
Q_ASSIGN U16144 ( .B(clk), .A(\g.we_clk [16630]));
Q_ASSIGN U16145 ( .B(clk), .A(\g.we_clk [16629]));
Q_ASSIGN U16146 ( .B(clk), .A(\g.we_clk [16628]));
Q_ASSIGN U16147 ( .B(clk), .A(\g.we_clk [16627]));
Q_ASSIGN U16148 ( .B(clk), .A(\g.we_clk [16626]));
Q_ASSIGN U16149 ( .B(clk), .A(\g.we_clk [16625]));
Q_ASSIGN U16150 ( .B(clk), .A(\g.we_clk [16624]));
Q_ASSIGN U16151 ( .B(clk), .A(\g.we_clk [16623]));
Q_ASSIGN U16152 ( .B(clk), .A(\g.we_clk [16622]));
Q_ASSIGN U16153 ( .B(clk), .A(\g.we_clk [16621]));
Q_ASSIGN U16154 ( .B(clk), .A(\g.we_clk [16620]));
Q_ASSIGN U16155 ( .B(clk), .A(\g.we_clk [16619]));
Q_ASSIGN U16156 ( .B(clk), .A(\g.we_clk [16618]));
Q_ASSIGN U16157 ( .B(clk), .A(\g.we_clk [16617]));
Q_ASSIGN U16158 ( .B(clk), .A(\g.we_clk [16616]));
Q_ASSIGN U16159 ( .B(clk), .A(\g.we_clk [16615]));
Q_ASSIGN U16160 ( .B(clk), .A(\g.we_clk [16614]));
Q_ASSIGN U16161 ( .B(clk), .A(\g.we_clk [16613]));
Q_ASSIGN U16162 ( .B(clk), .A(\g.we_clk [16612]));
Q_ASSIGN U16163 ( .B(clk), .A(\g.we_clk [16611]));
Q_ASSIGN U16164 ( .B(clk), .A(\g.we_clk [16610]));
Q_ASSIGN U16165 ( .B(clk), .A(\g.we_clk [16609]));
Q_ASSIGN U16166 ( .B(clk), .A(\g.we_clk [16608]));
Q_ASSIGN U16167 ( .B(clk), .A(\g.we_clk [16607]));
Q_ASSIGN U16168 ( .B(clk), .A(\g.we_clk [16606]));
Q_ASSIGN U16169 ( .B(clk), .A(\g.we_clk [16605]));
Q_ASSIGN U16170 ( .B(clk), .A(\g.we_clk [16604]));
Q_ASSIGN U16171 ( .B(clk), .A(\g.we_clk [16603]));
Q_ASSIGN U16172 ( .B(clk), .A(\g.we_clk [16602]));
Q_ASSIGN U16173 ( .B(clk), .A(\g.we_clk [16601]));
Q_ASSIGN U16174 ( .B(clk), .A(\g.we_clk [16600]));
Q_ASSIGN U16175 ( .B(clk), .A(\g.we_clk [16599]));
Q_ASSIGN U16176 ( .B(clk), .A(\g.we_clk [16598]));
Q_ASSIGN U16177 ( .B(clk), .A(\g.we_clk [16597]));
Q_ASSIGN U16178 ( .B(clk), .A(\g.we_clk [16596]));
Q_ASSIGN U16179 ( .B(clk), .A(\g.we_clk [16595]));
Q_ASSIGN U16180 ( .B(clk), .A(\g.we_clk [16594]));
Q_ASSIGN U16181 ( .B(clk), .A(\g.we_clk [16593]));
Q_ASSIGN U16182 ( .B(clk), .A(\g.we_clk [16592]));
Q_ASSIGN U16183 ( .B(clk), .A(\g.we_clk [16591]));
Q_ASSIGN U16184 ( .B(clk), .A(\g.we_clk [16590]));
Q_ASSIGN U16185 ( .B(clk), .A(\g.we_clk [16589]));
Q_ASSIGN U16186 ( .B(clk), .A(\g.we_clk [16588]));
Q_ASSIGN U16187 ( .B(clk), .A(\g.we_clk [16587]));
Q_ASSIGN U16188 ( .B(clk), .A(\g.we_clk [16586]));
Q_ASSIGN U16189 ( .B(clk), .A(\g.we_clk [16585]));
Q_ASSIGN U16190 ( .B(clk), .A(\g.we_clk [16584]));
Q_ASSIGN U16191 ( .B(clk), .A(\g.we_clk [16583]));
Q_ASSIGN U16192 ( .B(clk), .A(\g.we_clk [16582]));
Q_ASSIGN U16193 ( .B(clk), .A(\g.we_clk [16581]));
Q_ASSIGN U16194 ( .B(clk), .A(\g.we_clk [16580]));
Q_ASSIGN U16195 ( .B(clk), .A(\g.we_clk [16579]));
Q_ASSIGN U16196 ( .B(clk), .A(\g.we_clk [16578]));
Q_ASSIGN U16197 ( .B(clk), .A(\g.we_clk [16577]));
Q_ASSIGN U16198 ( .B(clk), .A(\g.we_clk [16576]));
Q_ASSIGN U16199 ( .B(clk), .A(\g.we_clk [16575]));
Q_ASSIGN U16200 ( .B(clk), .A(\g.we_clk [16574]));
Q_ASSIGN U16201 ( .B(clk), .A(\g.we_clk [16573]));
Q_ASSIGN U16202 ( .B(clk), .A(\g.we_clk [16572]));
Q_ASSIGN U16203 ( .B(clk), .A(\g.we_clk [16571]));
Q_ASSIGN U16204 ( .B(clk), .A(\g.we_clk [16570]));
Q_ASSIGN U16205 ( .B(clk), .A(\g.we_clk [16569]));
Q_ASSIGN U16206 ( .B(clk), .A(\g.we_clk [16568]));
Q_ASSIGN U16207 ( .B(clk), .A(\g.we_clk [16567]));
Q_ASSIGN U16208 ( .B(clk), .A(\g.we_clk [16566]));
Q_ASSIGN U16209 ( .B(clk), .A(\g.we_clk [16565]));
Q_ASSIGN U16210 ( .B(clk), .A(\g.we_clk [16564]));
Q_ASSIGN U16211 ( .B(clk), .A(\g.we_clk [16563]));
Q_ASSIGN U16212 ( .B(clk), .A(\g.we_clk [16562]));
Q_ASSIGN U16213 ( .B(clk), .A(\g.we_clk [16561]));
Q_ASSIGN U16214 ( .B(clk), .A(\g.we_clk [16560]));
Q_ASSIGN U16215 ( .B(clk), .A(\g.we_clk [16559]));
Q_ASSIGN U16216 ( .B(clk), .A(\g.we_clk [16558]));
Q_ASSIGN U16217 ( .B(clk), .A(\g.we_clk [16557]));
Q_ASSIGN U16218 ( .B(clk), .A(\g.we_clk [16556]));
Q_ASSIGN U16219 ( .B(clk), .A(\g.we_clk [16555]));
Q_ASSIGN U16220 ( .B(clk), .A(\g.we_clk [16554]));
Q_ASSIGN U16221 ( .B(clk), .A(\g.we_clk [16553]));
Q_ASSIGN U16222 ( .B(clk), .A(\g.we_clk [16552]));
Q_ASSIGN U16223 ( .B(clk), .A(\g.we_clk [16551]));
Q_ASSIGN U16224 ( .B(clk), .A(\g.we_clk [16550]));
Q_ASSIGN U16225 ( .B(clk), .A(\g.we_clk [16549]));
Q_ASSIGN U16226 ( .B(clk), .A(\g.we_clk [16548]));
Q_ASSIGN U16227 ( .B(clk), .A(\g.we_clk [16547]));
Q_ASSIGN U16228 ( .B(clk), .A(\g.we_clk [16546]));
Q_ASSIGN U16229 ( .B(clk), .A(\g.we_clk [16545]));
Q_ASSIGN U16230 ( .B(clk), .A(\g.we_clk [16544]));
Q_ASSIGN U16231 ( .B(clk), .A(\g.we_clk [16543]));
Q_ASSIGN U16232 ( .B(clk), .A(\g.we_clk [16542]));
Q_ASSIGN U16233 ( .B(clk), .A(\g.we_clk [16541]));
Q_ASSIGN U16234 ( .B(clk), .A(\g.we_clk [16540]));
Q_ASSIGN U16235 ( .B(clk), .A(\g.we_clk [16539]));
Q_ASSIGN U16236 ( .B(clk), .A(\g.we_clk [16538]));
Q_ASSIGN U16237 ( .B(clk), .A(\g.we_clk [16537]));
Q_ASSIGN U16238 ( .B(clk), .A(\g.we_clk [16536]));
Q_ASSIGN U16239 ( .B(clk), .A(\g.we_clk [16535]));
Q_ASSIGN U16240 ( .B(clk), .A(\g.we_clk [16534]));
Q_ASSIGN U16241 ( .B(clk), .A(\g.we_clk [16533]));
Q_ASSIGN U16242 ( .B(clk), .A(\g.we_clk [16532]));
Q_ASSIGN U16243 ( .B(clk), .A(\g.we_clk [16531]));
Q_ASSIGN U16244 ( .B(clk), .A(\g.we_clk [16530]));
Q_ASSIGN U16245 ( .B(clk), .A(\g.we_clk [16529]));
Q_ASSIGN U16246 ( .B(clk), .A(\g.we_clk [16528]));
Q_ASSIGN U16247 ( .B(clk), .A(\g.we_clk [16527]));
Q_ASSIGN U16248 ( .B(clk), .A(\g.we_clk [16526]));
Q_ASSIGN U16249 ( .B(clk), .A(\g.we_clk [16525]));
Q_ASSIGN U16250 ( .B(clk), .A(\g.we_clk [16524]));
Q_ASSIGN U16251 ( .B(clk), .A(\g.we_clk [16523]));
Q_ASSIGN U16252 ( .B(clk), .A(\g.we_clk [16522]));
Q_ASSIGN U16253 ( .B(clk), .A(\g.we_clk [16521]));
Q_ASSIGN U16254 ( .B(clk), .A(\g.we_clk [16520]));
Q_ASSIGN U16255 ( .B(clk), .A(\g.we_clk [16519]));
Q_ASSIGN U16256 ( .B(clk), .A(\g.we_clk [16518]));
Q_ASSIGN U16257 ( .B(clk), .A(\g.we_clk [16517]));
Q_ASSIGN U16258 ( .B(clk), .A(\g.we_clk [16516]));
Q_ASSIGN U16259 ( .B(clk), .A(\g.we_clk [16515]));
Q_ASSIGN U16260 ( .B(clk), .A(\g.we_clk [16514]));
Q_ASSIGN U16261 ( .B(clk), .A(\g.we_clk [16513]));
Q_ASSIGN U16262 ( .B(clk), .A(\g.we_clk [16512]));
Q_ASSIGN U16263 ( .B(clk), .A(\g.we_clk [16511]));
Q_ASSIGN U16264 ( .B(clk), .A(\g.we_clk [16510]));
Q_ASSIGN U16265 ( .B(clk), .A(\g.we_clk [16509]));
Q_ASSIGN U16266 ( .B(clk), .A(\g.we_clk [16508]));
Q_ASSIGN U16267 ( .B(clk), .A(\g.we_clk [16507]));
Q_ASSIGN U16268 ( .B(clk), .A(\g.we_clk [16506]));
Q_ASSIGN U16269 ( .B(clk), .A(\g.we_clk [16505]));
Q_ASSIGN U16270 ( .B(clk), .A(\g.we_clk [16504]));
Q_ASSIGN U16271 ( .B(clk), .A(\g.we_clk [16503]));
Q_ASSIGN U16272 ( .B(clk), .A(\g.we_clk [16502]));
Q_ASSIGN U16273 ( .B(clk), .A(\g.we_clk [16501]));
Q_ASSIGN U16274 ( .B(clk), .A(\g.we_clk [16500]));
Q_ASSIGN U16275 ( .B(clk), .A(\g.we_clk [16499]));
Q_ASSIGN U16276 ( .B(clk), .A(\g.we_clk [16498]));
Q_ASSIGN U16277 ( .B(clk), .A(\g.we_clk [16497]));
Q_ASSIGN U16278 ( .B(clk), .A(\g.we_clk [16496]));
Q_ASSIGN U16279 ( .B(clk), .A(\g.we_clk [16495]));
Q_ASSIGN U16280 ( .B(clk), .A(\g.we_clk [16494]));
Q_ASSIGN U16281 ( .B(clk), .A(\g.we_clk [16493]));
Q_ASSIGN U16282 ( .B(clk), .A(\g.we_clk [16492]));
Q_ASSIGN U16283 ( .B(clk), .A(\g.we_clk [16491]));
Q_ASSIGN U16284 ( .B(clk), .A(\g.we_clk [16490]));
Q_ASSIGN U16285 ( .B(clk), .A(\g.we_clk [16489]));
Q_ASSIGN U16286 ( .B(clk), .A(\g.we_clk [16488]));
Q_ASSIGN U16287 ( .B(clk), .A(\g.we_clk [16487]));
Q_ASSIGN U16288 ( .B(clk), .A(\g.we_clk [16486]));
Q_ASSIGN U16289 ( .B(clk), .A(\g.we_clk [16485]));
Q_ASSIGN U16290 ( .B(clk), .A(\g.we_clk [16484]));
Q_ASSIGN U16291 ( .B(clk), .A(\g.we_clk [16483]));
Q_ASSIGN U16292 ( .B(clk), .A(\g.we_clk [16482]));
Q_ASSIGN U16293 ( .B(clk), .A(\g.we_clk [16481]));
Q_ASSIGN U16294 ( .B(clk), .A(\g.we_clk [16480]));
Q_ASSIGN U16295 ( .B(clk), .A(\g.we_clk [16479]));
Q_ASSIGN U16296 ( .B(clk), .A(\g.we_clk [16478]));
Q_ASSIGN U16297 ( .B(clk), .A(\g.we_clk [16477]));
Q_ASSIGN U16298 ( .B(clk), .A(\g.we_clk [16476]));
Q_ASSIGN U16299 ( .B(clk), .A(\g.we_clk [16475]));
Q_ASSIGN U16300 ( .B(clk), .A(\g.we_clk [16474]));
Q_ASSIGN U16301 ( .B(clk), .A(\g.we_clk [16473]));
Q_ASSIGN U16302 ( .B(clk), .A(\g.we_clk [16472]));
Q_ASSIGN U16303 ( .B(clk), .A(\g.we_clk [16471]));
Q_ASSIGN U16304 ( .B(clk), .A(\g.we_clk [16470]));
Q_ASSIGN U16305 ( .B(clk), .A(\g.we_clk [16469]));
Q_ASSIGN U16306 ( .B(clk), .A(\g.we_clk [16468]));
Q_ASSIGN U16307 ( .B(clk), .A(\g.we_clk [16467]));
Q_ASSIGN U16308 ( .B(clk), .A(\g.we_clk [16466]));
Q_ASSIGN U16309 ( .B(clk), .A(\g.we_clk [16465]));
Q_ASSIGN U16310 ( .B(clk), .A(\g.we_clk [16464]));
Q_ASSIGN U16311 ( .B(clk), .A(\g.we_clk [16463]));
Q_ASSIGN U16312 ( .B(clk), .A(\g.we_clk [16462]));
Q_ASSIGN U16313 ( .B(clk), .A(\g.we_clk [16461]));
Q_ASSIGN U16314 ( .B(clk), .A(\g.we_clk [16460]));
Q_ASSIGN U16315 ( .B(clk), .A(\g.we_clk [16459]));
Q_ASSIGN U16316 ( .B(clk), .A(\g.we_clk [16458]));
Q_ASSIGN U16317 ( .B(clk), .A(\g.we_clk [16457]));
Q_ASSIGN U16318 ( .B(clk), .A(\g.we_clk [16456]));
Q_ASSIGN U16319 ( .B(clk), .A(\g.we_clk [16455]));
Q_ASSIGN U16320 ( .B(clk), .A(\g.we_clk [16454]));
Q_ASSIGN U16321 ( .B(clk), .A(\g.we_clk [16453]));
Q_ASSIGN U16322 ( .B(clk), .A(\g.we_clk [16452]));
Q_ASSIGN U16323 ( .B(clk), .A(\g.we_clk [16451]));
Q_ASSIGN U16324 ( .B(clk), .A(\g.we_clk [16450]));
Q_ASSIGN U16325 ( .B(clk), .A(\g.we_clk [16449]));
Q_ASSIGN U16326 ( .B(clk), .A(\g.we_clk [16448]));
Q_ASSIGN U16327 ( .B(clk), .A(\g.we_clk [16447]));
Q_ASSIGN U16328 ( .B(clk), .A(\g.we_clk [16446]));
Q_ASSIGN U16329 ( .B(clk), .A(\g.we_clk [16445]));
Q_ASSIGN U16330 ( .B(clk), .A(\g.we_clk [16444]));
Q_ASSIGN U16331 ( .B(clk), .A(\g.we_clk [16443]));
Q_ASSIGN U16332 ( .B(clk), .A(\g.we_clk [16442]));
Q_ASSIGN U16333 ( .B(clk), .A(\g.we_clk [16441]));
Q_ASSIGN U16334 ( .B(clk), .A(\g.we_clk [16440]));
Q_ASSIGN U16335 ( .B(clk), .A(\g.we_clk [16439]));
Q_ASSIGN U16336 ( .B(clk), .A(\g.we_clk [16438]));
Q_ASSIGN U16337 ( .B(clk), .A(\g.we_clk [16437]));
Q_ASSIGN U16338 ( .B(clk), .A(\g.we_clk [16436]));
Q_ASSIGN U16339 ( .B(clk), .A(\g.we_clk [16435]));
Q_ASSIGN U16340 ( .B(clk), .A(\g.we_clk [16434]));
Q_ASSIGN U16341 ( .B(clk), .A(\g.we_clk [16433]));
Q_ASSIGN U16342 ( .B(clk), .A(\g.we_clk [16432]));
Q_ASSIGN U16343 ( .B(clk), .A(\g.we_clk [16431]));
Q_ASSIGN U16344 ( .B(clk), .A(\g.we_clk [16430]));
Q_ASSIGN U16345 ( .B(clk), .A(\g.we_clk [16429]));
Q_ASSIGN U16346 ( .B(clk), .A(\g.we_clk [16428]));
Q_ASSIGN U16347 ( .B(clk), .A(\g.we_clk [16427]));
Q_ASSIGN U16348 ( .B(clk), .A(\g.we_clk [16426]));
Q_ASSIGN U16349 ( .B(clk), .A(\g.we_clk [16425]));
Q_ASSIGN U16350 ( .B(clk), .A(\g.we_clk [16424]));
Q_ASSIGN U16351 ( .B(clk), .A(\g.we_clk [16423]));
Q_ASSIGN U16352 ( .B(clk), .A(\g.we_clk [16422]));
Q_ASSIGN U16353 ( .B(clk), .A(\g.we_clk [16421]));
Q_ASSIGN U16354 ( .B(clk), .A(\g.we_clk [16420]));
Q_ASSIGN U16355 ( .B(clk), .A(\g.we_clk [16419]));
Q_ASSIGN U16356 ( .B(clk), .A(\g.we_clk [16418]));
Q_ASSIGN U16357 ( .B(clk), .A(\g.we_clk [16417]));
Q_ASSIGN U16358 ( .B(clk), .A(\g.we_clk [16416]));
Q_ASSIGN U16359 ( .B(clk), .A(\g.we_clk [16415]));
Q_ASSIGN U16360 ( .B(clk), .A(\g.we_clk [16414]));
Q_ASSIGN U16361 ( .B(clk), .A(\g.we_clk [16413]));
Q_ASSIGN U16362 ( .B(clk), .A(\g.we_clk [16412]));
Q_ASSIGN U16363 ( .B(clk), .A(\g.we_clk [16411]));
Q_ASSIGN U16364 ( .B(clk), .A(\g.we_clk [16410]));
Q_ASSIGN U16365 ( .B(clk), .A(\g.we_clk [16409]));
Q_ASSIGN U16366 ( .B(clk), .A(\g.we_clk [16408]));
Q_ASSIGN U16367 ( .B(clk), .A(\g.we_clk [16407]));
Q_ASSIGN U16368 ( .B(clk), .A(\g.we_clk [16406]));
Q_ASSIGN U16369 ( .B(clk), .A(\g.we_clk [16405]));
Q_ASSIGN U16370 ( .B(clk), .A(\g.we_clk [16404]));
Q_ASSIGN U16371 ( .B(clk), .A(\g.we_clk [16403]));
Q_ASSIGN U16372 ( .B(clk), .A(\g.we_clk [16402]));
Q_ASSIGN U16373 ( .B(clk), .A(\g.we_clk [16401]));
Q_ASSIGN U16374 ( .B(clk), .A(\g.we_clk [16400]));
Q_ASSIGN U16375 ( .B(clk), .A(\g.we_clk [16399]));
Q_ASSIGN U16376 ( .B(clk), .A(\g.we_clk [16398]));
Q_ASSIGN U16377 ( .B(clk), .A(\g.we_clk [16397]));
Q_ASSIGN U16378 ( .B(clk), .A(\g.we_clk [16396]));
Q_ASSIGN U16379 ( .B(clk), .A(\g.we_clk [16395]));
Q_ASSIGN U16380 ( .B(clk), .A(\g.we_clk [16394]));
Q_ASSIGN U16381 ( .B(clk), .A(\g.we_clk [16393]));
Q_ASSIGN U16382 ( .B(clk), .A(\g.we_clk [16392]));
Q_ASSIGN U16383 ( .B(clk), .A(\g.we_clk [16391]));
Q_ASSIGN U16384 ( .B(clk), .A(\g.we_clk [16390]));
Q_ASSIGN U16385 ( .B(clk), .A(\g.we_clk [16389]));
Q_ASSIGN U16386 ( .B(clk), .A(\g.we_clk [16388]));
Q_ASSIGN U16387 ( .B(clk), .A(\g.we_clk [16387]));
Q_ASSIGN U16388 ( .B(clk), .A(\g.we_clk [16386]));
Q_ASSIGN U16389 ( .B(clk), .A(\g.we_clk [16385]));
Q_ASSIGN U16390 ( .B(clk), .A(\g.we_clk [16384]));
Q_ASSIGN U16391 ( .B(clk), .A(\g.we_clk [16383]));
Q_ASSIGN U16392 ( .B(clk), .A(\g.we_clk [16382]));
Q_ASSIGN U16393 ( .B(clk), .A(\g.we_clk [16381]));
Q_ASSIGN U16394 ( .B(clk), .A(\g.we_clk [16380]));
Q_ASSIGN U16395 ( .B(clk), .A(\g.we_clk [16379]));
Q_ASSIGN U16396 ( .B(clk), .A(\g.we_clk [16378]));
Q_ASSIGN U16397 ( .B(clk), .A(\g.we_clk [16377]));
Q_ASSIGN U16398 ( .B(clk), .A(\g.we_clk [16376]));
Q_ASSIGN U16399 ( .B(clk), .A(\g.we_clk [16375]));
Q_ASSIGN U16400 ( .B(clk), .A(\g.we_clk [16374]));
Q_ASSIGN U16401 ( .B(clk), .A(\g.we_clk [16373]));
Q_ASSIGN U16402 ( .B(clk), .A(\g.we_clk [16372]));
Q_ASSIGN U16403 ( .B(clk), .A(\g.we_clk [16371]));
Q_ASSIGN U16404 ( .B(clk), .A(\g.we_clk [16370]));
Q_ASSIGN U16405 ( .B(clk), .A(\g.we_clk [16369]));
Q_ASSIGN U16406 ( .B(clk), .A(\g.we_clk [16368]));
Q_ASSIGN U16407 ( .B(clk), .A(\g.we_clk [16367]));
Q_ASSIGN U16408 ( .B(clk), .A(\g.we_clk [16366]));
Q_ASSIGN U16409 ( .B(clk), .A(\g.we_clk [16365]));
Q_ASSIGN U16410 ( .B(clk), .A(\g.we_clk [16364]));
Q_ASSIGN U16411 ( .B(clk), .A(\g.we_clk [16363]));
Q_ASSIGN U16412 ( .B(clk), .A(\g.we_clk [16362]));
Q_ASSIGN U16413 ( .B(clk), .A(\g.we_clk [16361]));
Q_ASSIGN U16414 ( .B(clk), .A(\g.we_clk [16360]));
Q_ASSIGN U16415 ( .B(clk), .A(\g.we_clk [16359]));
Q_ASSIGN U16416 ( .B(clk), .A(\g.we_clk [16358]));
Q_ASSIGN U16417 ( .B(clk), .A(\g.we_clk [16357]));
Q_ASSIGN U16418 ( .B(clk), .A(\g.we_clk [16356]));
Q_ASSIGN U16419 ( .B(clk), .A(\g.we_clk [16355]));
Q_ASSIGN U16420 ( .B(clk), .A(\g.we_clk [16354]));
Q_ASSIGN U16421 ( .B(clk), .A(\g.we_clk [16353]));
Q_ASSIGN U16422 ( .B(clk), .A(\g.we_clk [16352]));
Q_ASSIGN U16423 ( .B(clk), .A(\g.we_clk [16351]));
Q_ASSIGN U16424 ( .B(clk), .A(\g.we_clk [16350]));
Q_ASSIGN U16425 ( .B(clk), .A(\g.we_clk [16349]));
Q_ASSIGN U16426 ( .B(clk), .A(\g.we_clk [16348]));
Q_ASSIGN U16427 ( .B(clk), .A(\g.we_clk [16347]));
Q_ASSIGN U16428 ( .B(clk), .A(\g.we_clk [16346]));
Q_ASSIGN U16429 ( .B(clk), .A(\g.we_clk [16345]));
Q_ASSIGN U16430 ( .B(clk), .A(\g.we_clk [16344]));
Q_ASSIGN U16431 ( .B(clk), .A(\g.we_clk [16343]));
Q_ASSIGN U16432 ( .B(clk), .A(\g.we_clk [16342]));
Q_ASSIGN U16433 ( .B(clk), .A(\g.we_clk [16341]));
Q_ASSIGN U16434 ( .B(clk), .A(\g.we_clk [16340]));
Q_ASSIGN U16435 ( .B(clk), .A(\g.we_clk [16339]));
Q_ASSIGN U16436 ( .B(clk), .A(\g.we_clk [16338]));
Q_ASSIGN U16437 ( .B(clk), .A(\g.we_clk [16337]));
Q_ASSIGN U16438 ( .B(clk), .A(\g.we_clk [16336]));
Q_ASSIGN U16439 ( .B(clk), .A(\g.we_clk [16335]));
Q_ASSIGN U16440 ( .B(clk), .A(\g.we_clk [16334]));
Q_ASSIGN U16441 ( .B(clk), .A(\g.we_clk [16333]));
Q_ASSIGN U16442 ( .B(clk), .A(\g.we_clk [16332]));
Q_ASSIGN U16443 ( .B(clk), .A(\g.we_clk [16331]));
Q_ASSIGN U16444 ( .B(clk), .A(\g.we_clk [16330]));
Q_ASSIGN U16445 ( .B(clk), .A(\g.we_clk [16329]));
Q_ASSIGN U16446 ( .B(clk), .A(\g.we_clk [16328]));
Q_ASSIGN U16447 ( .B(clk), .A(\g.we_clk [16327]));
Q_ASSIGN U16448 ( .B(clk), .A(\g.we_clk [16326]));
Q_ASSIGN U16449 ( .B(clk), .A(\g.we_clk [16325]));
Q_ASSIGN U16450 ( .B(clk), .A(\g.we_clk [16324]));
Q_ASSIGN U16451 ( .B(clk), .A(\g.we_clk [16323]));
Q_ASSIGN U16452 ( .B(clk), .A(\g.we_clk [16322]));
Q_ASSIGN U16453 ( .B(clk), .A(\g.we_clk [16321]));
Q_ASSIGN U16454 ( .B(clk), .A(\g.we_clk [16320]));
Q_ASSIGN U16455 ( .B(clk), .A(\g.we_clk [16319]));
Q_ASSIGN U16456 ( .B(clk), .A(\g.we_clk [16318]));
Q_ASSIGN U16457 ( .B(clk), .A(\g.we_clk [16317]));
Q_ASSIGN U16458 ( .B(clk), .A(\g.we_clk [16316]));
Q_ASSIGN U16459 ( .B(clk), .A(\g.we_clk [16315]));
Q_ASSIGN U16460 ( .B(clk), .A(\g.we_clk [16314]));
Q_ASSIGN U16461 ( .B(clk), .A(\g.we_clk [16313]));
Q_ASSIGN U16462 ( .B(clk), .A(\g.we_clk [16312]));
Q_ASSIGN U16463 ( .B(clk), .A(\g.we_clk [16311]));
Q_ASSIGN U16464 ( .B(clk), .A(\g.we_clk [16310]));
Q_ASSIGN U16465 ( .B(clk), .A(\g.we_clk [16309]));
Q_ASSIGN U16466 ( .B(clk), .A(\g.we_clk [16308]));
Q_ASSIGN U16467 ( .B(clk), .A(\g.we_clk [16307]));
Q_ASSIGN U16468 ( .B(clk), .A(\g.we_clk [16306]));
Q_ASSIGN U16469 ( .B(clk), .A(\g.we_clk [16305]));
Q_ASSIGN U16470 ( .B(clk), .A(\g.we_clk [16304]));
Q_ASSIGN U16471 ( .B(clk), .A(\g.we_clk [16303]));
Q_ASSIGN U16472 ( .B(clk), .A(\g.we_clk [16302]));
Q_ASSIGN U16473 ( .B(clk), .A(\g.we_clk [16301]));
Q_ASSIGN U16474 ( .B(clk), .A(\g.we_clk [16300]));
Q_ASSIGN U16475 ( .B(clk), .A(\g.we_clk [16299]));
Q_ASSIGN U16476 ( .B(clk), .A(\g.we_clk [16298]));
Q_ASSIGN U16477 ( .B(clk), .A(\g.we_clk [16297]));
Q_ASSIGN U16478 ( .B(clk), .A(\g.we_clk [16296]));
Q_ASSIGN U16479 ( .B(clk), .A(\g.we_clk [16295]));
Q_ASSIGN U16480 ( .B(clk), .A(\g.we_clk [16294]));
Q_ASSIGN U16481 ( .B(clk), .A(\g.we_clk [16293]));
Q_ASSIGN U16482 ( .B(clk), .A(\g.we_clk [16292]));
Q_ASSIGN U16483 ( .B(clk), .A(\g.we_clk [16291]));
Q_ASSIGN U16484 ( .B(clk), .A(\g.we_clk [16290]));
Q_ASSIGN U16485 ( .B(clk), .A(\g.we_clk [16289]));
Q_ASSIGN U16486 ( .B(clk), .A(\g.we_clk [16288]));
Q_ASSIGN U16487 ( .B(clk), .A(\g.we_clk [16287]));
Q_ASSIGN U16488 ( .B(clk), .A(\g.we_clk [16286]));
Q_ASSIGN U16489 ( .B(clk), .A(\g.we_clk [16285]));
Q_ASSIGN U16490 ( .B(clk), .A(\g.we_clk [16284]));
Q_ASSIGN U16491 ( .B(clk), .A(\g.we_clk [16283]));
Q_ASSIGN U16492 ( .B(clk), .A(\g.we_clk [16282]));
Q_ASSIGN U16493 ( .B(clk), .A(\g.we_clk [16281]));
Q_ASSIGN U16494 ( .B(clk), .A(\g.we_clk [16280]));
Q_ASSIGN U16495 ( .B(clk), .A(\g.we_clk [16279]));
Q_ASSIGN U16496 ( .B(clk), .A(\g.we_clk [16278]));
Q_ASSIGN U16497 ( .B(clk), .A(\g.we_clk [16277]));
Q_ASSIGN U16498 ( .B(clk), .A(\g.we_clk [16276]));
Q_ASSIGN U16499 ( .B(clk), .A(\g.we_clk [16275]));
Q_ASSIGN U16500 ( .B(clk), .A(\g.we_clk [16274]));
Q_ASSIGN U16501 ( .B(clk), .A(\g.we_clk [16273]));
Q_ASSIGN U16502 ( .B(clk), .A(\g.we_clk [16272]));
Q_ASSIGN U16503 ( .B(clk), .A(\g.we_clk [16271]));
Q_ASSIGN U16504 ( .B(clk), .A(\g.we_clk [16270]));
Q_ASSIGN U16505 ( .B(clk), .A(\g.we_clk [16269]));
Q_ASSIGN U16506 ( .B(clk), .A(\g.we_clk [16268]));
Q_ASSIGN U16507 ( .B(clk), .A(\g.we_clk [16267]));
Q_ASSIGN U16508 ( .B(clk), .A(\g.we_clk [16266]));
Q_ASSIGN U16509 ( .B(clk), .A(\g.we_clk [16265]));
Q_ASSIGN U16510 ( .B(clk), .A(\g.we_clk [16264]));
Q_ASSIGN U16511 ( .B(clk), .A(\g.we_clk [16263]));
Q_ASSIGN U16512 ( .B(clk), .A(\g.we_clk [16262]));
Q_ASSIGN U16513 ( .B(clk), .A(\g.we_clk [16261]));
Q_ASSIGN U16514 ( .B(clk), .A(\g.we_clk [16260]));
Q_ASSIGN U16515 ( .B(clk), .A(\g.we_clk [16259]));
Q_ASSIGN U16516 ( .B(clk), .A(\g.we_clk [16258]));
Q_ASSIGN U16517 ( .B(clk), .A(\g.we_clk [16257]));
Q_ASSIGN U16518 ( .B(clk), .A(\g.we_clk [16256]));
Q_ASSIGN U16519 ( .B(clk), .A(\g.we_clk [16255]));
Q_ASSIGN U16520 ( .B(clk), .A(\g.we_clk [16254]));
Q_ASSIGN U16521 ( .B(clk), .A(\g.we_clk [16253]));
Q_ASSIGN U16522 ( .B(clk), .A(\g.we_clk [16252]));
Q_ASSIGN U16523 ( .B(clk), .A(\g.we_clk [16251]));
Q_ASSIGN U16524 ( .B(clk), .A(\g.we_clk [16250]));
Q_ASSIGN U16525 ( .B(clk), .A(\g.we_clk [16249]));
Q_ASSIGN U16526 ( .B(clk), .A(\g.we_clk [16248]));
Q_ASSIGN U16527 ( .B(clk), .A(\g.we_clk [16247]));
Q_ASSIGN U16528 ( .B(clk), .A(\g.we_clk [16246]));
Q_ASSIGN U16529 ( .B(clk), .A(\g.we_clk [16245]));
Q_ASSIGN U16530 ( .B(clk), .A(\g.we_clk [16244]));
Q_ASSIGN U16531 ( .B(clk), .A(\g.we_clk [16243]));
Q_ASSIGN U16532 ( .B(clk), .A(\g.we_clk [16242]));
Q_ASSIGN U16533 ( .B(clk), .A(\g.we_clk [16241]));
Q_ASSIGN U16534 ( .B(clk), .A(\g.we_clk [16240]));
Q_ASSIGN U16535 ( .B(clk), .A(\g.we_clk [16239]));
Q_ASSIGN U16536 ( .B(clk), .A(\g.we_clk [16238]));
Q_ASSIGN U16537 ( .B(clk), .A(\g.we_clk [16237]));
Q_ASSIGN U16538 ( .B(clk), .A(\g.we_clk [16236]));
Q_ASSIGN U16539 ( .B(clk), .A(\g.we_clk [16235]));
Q_ASSIGN U16540 ( .B(clk), .A(\g.we_clk [16234]));
Q_ASSIGN U16541 ( .B(clk), .A(\g.we_clk [16233]));
Q_ASSIGN U16542 ( .B(clk), .A(\g.we_clk [16232]));
Q_ASSIGN U16543 ( .B(clk), .A(\g.we_clk [16231]));
Q_ASSIGN U16544 ( .B(clk), .A(\g.we_clk [16230]));
Q_ASSIGN U16545 ( .B(clk), .A(\g.we_clk [16229]));
Q_ASSIGN U16546 ( .B(clk), .A(\g.we_clk [16228]));
Q_ASSIGN U16547 ( .B(clk), .A(\g.we_clk [16227]));
Q_ASSIGN U16548 ( .B(clk), .A(\g.we_clk [16226]));
Q_ASSIGN U16549 ( .B(clk), .A(\g.we_clk [16225]));
Q_ASSIGN U16550 ( .B(clk), .A(\g.we_clk [16224]));
Q_ASSIGN U16551 ( .B(clk), .A(\g.we_clk [16223]));
Q_ASSIGN U16552 ( .B(clk), .A(\g.we_clk [16222]));
Q_ASSIGN U16553 ( .B(clk), .A(\g.we_clk [16221]));
Q_ASSIGN U16554 ( .B(clk), .A(\g.we_clk [16220]));
Q_ASSIGN U16555 ( .B(clk), .A(\g.we_clk [16219]));
Q_ASSIGN U16556 ( .B(clk), .A(\g.we_clk [16218]));
Q_ASSIGN U16557 ( .B(clk), .A(\g.we_clk [16217]));
Q_ASSIGN U16558 ( .B(clk), .A(\g.we_clk [16216]));
Q_ASSIGN U16559 ( .B(clk), .A(\g.we_clk [16215]));
Q_ASSIGN U16560 ( .B(clk), .A(\g.we_clk [16214]));
Q_ASSIGN U16561 ( .B(clk), .A(\g.we_clk [16213]));
Q_ASSIGN U16562 ( .B(clk), .A(\g.we_clk [16212]));
Q_ASSIGN U16563 ( .B(clk), .A(\g.we_clk [16211]));
Q_ASSIGN U16564 ( .B(clk), .A(\g.we_clk [16210]));
Q_ASSIGN U16565 ( .B(clk), .A(\g.we_clk [16209]));
Q_ASSIGN U16566 ( .B(clk), .A(\g.we_clk [16208]));
Q_ASSIGN U16567 ( .B(clk), .A(\g.we_clk [16207]));
Q_ASSIGN U16568 ( .B(clk), .A(\g.we_clk [16206]));
Q_ASSIGN U16569 ( .B(clk), .A(\g.we_clk [16205]));
Q_ASSIGN U16570 ( .B(clk), .A(\g.we_clk [16204]));
Q_ASSIGN U16571 ( .B(clk), .A(\g.we_clk [16203]));
Q_ASSIGN U16572 ( .B(clk), .A(\g.we_clk [16202]));
Q_ASSIGN U16573 ( .B(clk), .A(\g.we_clk [16201]));
Q_ASSIGN U16574 ( .B(clk), .A(\g.we_clk [16200]));
Q_ASSIGN U16575 ( .B(clk), .A(\g.we_clk [16199]));
Q_ASSIGN U16576 ( .B(clk), .A(\g.we_clk [16198]));
Q_ASSIGN U16577 ( .B(clk), .A(\g.we_clk [16197]));
Q_ASSIGN U16578 ( .B(clk), .A(\g.we_clk [16196]));
Q_ASSIGN U16579 ( .B(clk), .A(\g.we_clk [16195]));
Q_ASSIGN U16580 ( .B(clk), .A(\g.we_clk [16194]));
Q_ASSIGN U16581 ( .B(clk), .A(\g.we_clk [16193]));
Q_ASSIGN U16582 ( .B(clk), .A(\g.we_clk [16192]));
Q_ASSIGN U16583 ( .B(clk), .A(\g.we_clk [16191]));
Q_ASSIGN U16584 ( .B(clk), .A(\g.we_clk [16190]));
Q_ASSIGN U16585 ( .B(clk), .A(\g.we_clk [16189]));
Q_ASSIGN U16586 ( .B(clk), .A(\g.we_clk [16188]));
Q_ASSIGN U16587 ( .B(clk), .A(\g.we_clk [16187]));
Q_ASSIGN U16588 ( .B(clk), .A(\g.we_clk [16186]));
Q_ASSIGN U16589 ( .B(clk), .A(\g.we_clk [16185]));
Q_ASSIGN U16590 ( .B(clk), .A(\g.we_clk [16184]));
Q_ASSIGN U16591 ( .B(clk), .A(\g.we_clk [16183]));
Q_ASSIGN U16592 ( .B(clk), .A(\g.we_clk [16182]));
Q_ASSIGN U16593 ( .B(clk), .A(\g.we_clk [16181]));
Q_ASSIGN U16594 ( .B(clk), .A(\g.we_clk [16180]));
Q_ASSIGN U16595 ( .B(clk), .A(\g.we_clk [16179]));
Q_ASSIGN U16596 ( .B(clk), .A(\g.we_clk [16178]));
Q_ASSIGN U16597 ( .B(clk), .A(\g.we_clk [16177]));
Q_ASSIGN U16598 ( .B(clk), .A(\g.we_clk [16176]));
Q_ASSIGN U16599 ( .B(clk), .A(\g.we_clk [16175]));
Q_ASSIGN U16600 ( .B(clk), .A(\g.we_clk [16174]));
Q_ASSIGN U16601 ( .B(clk), .A(\g.we_clk [16173]));
Q_ASSIGN U16602 ( .B(clk), .A(\g.we_clk [16172]));
Q_ASSIGN U16603 ( .B(clk), .A(\g.we_clk [16171]));
Q_ASSIGN U16604 ( .B(clk), .A(\g.we_clk [16170]));
Q_ASSIGN U16605 ( .B(clk), .A(\g.we_clk [16169]));
Q_ASSIGN U16606 ( .B(clk), .A(\g.we_clk [16168]));
Q_ASSIGN U16607 ( .B(clk), .A(\g.we_clk [16167]));
Q_ASSIGN U16608 ( .B(clk), .A(\g.we_clk [16166]));
Q_ASSIGN U16609 ( .B(clk), .A(\g.we_clk [16165]));
Q_ASSIGN U16610 ( .B(clk), .A(\g.we_clk [16164]));
Q_ASSIGN U16611 ( .B(clk), .A(\g.we_clk [16163]));
Q_ASSIGN U16612 ( .B(clk), .A(\g.we_clk [16162]));
Q_ASSIGN U16613 ( .B(clk), .A(\g.we_clk [16161]));
Q_ASSIGN U16614 ( .B(clk), .A(\g.we_clk [16160]));
Q_ASSIGN U16615 ( .B(clk), .A(\g.we_clk [16159]));
Q_ASSIGN U16616 ( .B(clk), .A(\g.we_clk [16158]));
Q_ASSIGN U16617 ( .B(clk), .A(\g.we_clk [16157]));
Q_ASSIGN U16618 ( .B(clk), .A(\g.we_clk [16156]));
Q_ASSIGN U16619 ( .B(clk), .A(\g.we_clk [16155]));
Q_ASSIGN U16620 ( .B(clk), .A(\g.we_clk [16154]));
Q_ASSIGN U16621 ( .B(clk), .A(\g.we_clk [16153]));
Q_ASSIGN U16622 ( .B(clk), .A(\g.we_clk [16152]));
Q_ASSIGN U16623 ( .B(clk), .A(\g.we_clk [16151]));
Q_ASSIGN U16624 ( .B(clk), .A(\g.we_clk [16150]));
Q_ASSIGN U16625 ( .B(clk), .A(\g.we_clk [16149]));
Q_ASSIGN U16626 ( .B(clk), .A(\g.we_clk [16148]));
Q_ASSIGN U16627 ( .B(clk), .A(\g.we_clk [16147]));
Q_ASSIGN U16628 ( .B(clk), .A(\g.we_clk [16146]));
Q_ASSIGN U16629 ( .B(clk), .A(\g.we_clk [16145]));
Q_ASSIGN U16630 ( .B(clk), .A(\g.we_clk [16144]));
Q_ASSIGN U16631 ( .B(clk), .A(\g.we_clk [16143]));
Q_ASSIGN U16632 ( .B(clk), .A(\g.we_clk [16142]));
Q_ASSIGN U16633 ( .B(clk), .A(\g.we_clk [16141]));
Q_ASSIGN U16634 ( .B(clk), .A(\g.we_clk [16140]));
Q_ASSIGN U16635 ( .B(clk), .A(\g.we_clk [16139]));
Q_ASSIGN U16636 ( .B(clk), .A(\g.we_clk [16138]));
Q_ASSIGN U16637 ( .B(clk), .A(\g.we_clk [16137]));
Q_ASSIGN U16638 ( .B(clk), .A(\g.we_clk [16136]));
Q_ASSIGN U16639 ( .B(clk), .A(\g.we_clk [16135]));
Q_ASSIGN U16640 ( .B(clk), .A(\g.we_clk [16134]));
Q_ASSIGN U16641 ( .B(clk), .A(\g.we_clk [16133]));
Q_ASSIGN U16642 ( .B(clk), .A(\g.we_clk [16132]));
Q_ASSIGN U16643 ( .B(clk), .A(\g.we_clk [16131]));
Q_ASSIGN U16644 ( .B(clk), .A(\g.we_clk [16130]));
Q_ASSIGN U16645 ( .B(clk), .A(\g.we_clk [16129]));
Q_ASSIGN U16646 ( .B(clk), .A(\g.we_clk [16128]));
Q_ASSIGN U16647 ( .B(clk), .A(\g.we_clk [16127]));
Q_ASSIGN U16648 ( .B(clk), .A(\g.we_clk [16126]));
Q_ASSIGN U16649 ( .B(clk), .A(\g.we_clk [16125]));
Q_ASSIGN U16650 ( .B(clk), .A(\g.we_clk [16124]));
Q_ASSIGN U16651 ( .B(clk), .A(\g.we_clk [16123]));
Q_ASSIGN U16652 ( .B(clk), .A(\g.we_clk [16122]));
Q_ASSIGN U16653 ( .B(clk), .A(\g.we_clk [16121]));
Q_ASSIGN U16654 ( .B(clk), .A(\g.we_clk [16120]));
Q_ASSIGN U16655 ( .B(clk), .A(\g.we_clk [16119]));
Q_ASSIGN U16656 ( .B(clk), .A(\g.we_clk [16118]));
Q_ASSIGN U16657 ( .B(clk), .A(\g.we_clk [16117]));
Q_ASSIGN U16658 ( .B(clk), .A(\g.we_clk [16116]));
Q_ASSIGN U16659 ( .B(clk), .A(\g.we_clk [16115]));
Q_ASSIGN U16660 ( .B(clk), .A(\g.we_clk [16114]));
Q_ASSIGN U16661 ( .B(clk), .A(\g.we_clk [16113]));
Q_ASSIGN U16662 ( .B(clk), .A(\g.we_clk [16112]));
Q_ASSIGN U16663 ( .B(clk), .A(\g.we_clk [16111]));
Q_ASSIGN U16664 ( .B(clk), .A(\g.we_clk [16110]));
Q_ASSIGN U16665 ( .B(clk), .A(\g.we_clk [16109]));
Q_ASSIGN U16666 ( .B(clk), .A(\g.we_clk [16108]));
Q_ASSIGN U16667 ( .B(clk), .A(\g.we_clk [16107]));
Q_ASSIGN U16668 ( .B(clk), .A(\g.we_clk [16106]));
Q_ASSIGN U16669 ( .B(clk), .A(\g.we_clk [16105]));
Q_ASSIGN U16670 ( .B(clk), .A(\g.we_clk [16104]));
Q_ASSIGN U16671 ( .B(clk), .A(\g.we_clk [16103]));
Q_ASSIGN U16672 ( .B(clk), .A(\g.we_clk [16102]));
Q_ASSIGN U16673 ( .B(clk), .A(\g.we_clk [16101]));
Q_ASSIGN U16674 ( .B(clk), .A(\g.we_clk [16100]));
Q_ASSIGN U16675 ( .B(clk), .A(\g.we_clk [16099]));
Q_ASSIGN U16676 ( .B(clk), .A(\g.we_clk [16098]));
Q_ASSIGN U16677 ( .B(clk), .A(\g.we_clk [16097]));
Q_ASSIGN U16678 ( .B(clk), .A(\g.we_clk [16096]));
Q_ASSIGN U16679 ( .B(clk), .A(\g.we_clk [16095]));
Q_ASSIGN U16680 ( .B(clk), .A(\g.we_clk [16094]));
Q_ASSIGN U16681 ( .B(clk), .A(\g.we_clk [16093]));
Q_ASSIGN U16682 ( .B(clk), .A(\g.we_clk [16092]));
Q_ASSIGN U16683 ( .B(clk), .A(\g.we_clk [16091]));
Q_ASSIGN U16684 ( .B(clk), .A(\g.we_clk [16090]));
Q_ASSIGN U16685 ( .B(clk), .A(\g.we_clk [16089]));
Q_ASSIGN U16686 ( .B(clk), .A(\g.we_clk [16088]));
Q_ASSIGN U16687 ( .B(clk), .A(\g.we_clk [16087]));
Q_ASSIGN U16688 ( .B(clk), .A(\g.we_clk [16086]));
Q_ASSIGN U16689 ( .B(clk), .A(\g.we_clk [16085]));
Q_ASSIGN U16690 ( .B(clk), .A(\g.we_clk [16084]));
Q_ASSIGN U16691 ( .B(clk), .A(\g.we_clk [16083]));
Q_ASSIGN U16692 ( .B(clk), .A(\g.we_clk [16082]));
Q_ASSIGN U16693 ( .B(clk), .A(\g.we_clk [16081]));
Q_ASSIGN U16694 ( .B(clk), .A(\g.we_clk [16080]));
Q_ASSIGN U16695 ( .B(clk), .A(\g.we_clk [16079]));
Q_ASSIGN U16696 ( .B(clk), .A(\g.we_clk [16078]));
Q_ASSIGN U16697 ( .B(clk), .A(\g.we_clk [16077]));
Q_ASSIGN U16698 ( .B(clk), .A(\g.we_clk [16076]));
Q_ASSIGN U16699 ( .B(clk), .A(\g.we_clk [16075]));
Q_ASSIGN U16700 ( .B(clk), .A(\g.we_clk [16074]));
Q_ASSIGN U16701 ( .B(clk), .A(\g.we_clk [16073]));
Q_ASSIGN U16702 ( .B(clk), .A(\g.we_clk [16072]));
Q_ASSIGN U16703 ( .B(clk), .A(\g.we_clk [16071]));
Q_ASSIGN U16704 ( .B(clk), .A(\g.we_clk [16070]));
Q_ASSIGN U16705 ( .B(clk), .A(\g.we_clk [16069]));
Q_ASSIGN U16706 ( .B(clk), .A(\g.we_clk [16068]));
Q_ASSIGN U16707 ( .B(clk), .A(\g.we_clk [16067]));
Q_ASSIGN U16708 ( .B(clk), .A(\g.we_clk [16066]));
Q_ASSIGN U16709 ( .B(clk), .A(\g.we_clk [16065]));
Q_ASSIGN U16710 ( .B(clk), .A(\g.we_clk [16064]));
Q_ASSIGN U16711 ( .B(clk), .A(\g.we_clk [16063]));
Q_ASSIGN U16712 ( .B(clk), .A(\g.we_clk [16062]));
Q_ASSIGN U16713 ( .B(clk), .A(\g.we_clk [16061]));
Q_ASSIGN U16714 ( .B(clk), .A(\g.we_clk [16060]));
Q_ASSIGN U16715 ( .B(clk), .A(\g.we_clk [16059]));
Q_ASSIGN U16716 ( .B(clk), .A(\g.we_clk [16058]));
Q_ASSIGN U16717 ( .B(clk), .A(\g.we_clk [16057]));
Q_ASSIGN U16718 ( .B(clk), .A(\g.we_clk [16056]));
Q_ASSIGN U16719 ( .B(clk), .A(\g.we_clk [16055]));
Q_ASSIGN U16720 ( .B(clk), .A(\g.we_clk [16054]));
Q_ASSIGN U16721 ( .B(clk), .A(\g.we_clk [16053]));
Q_ASSIGN U16722 ( .B(clk), .A(\g.we_clk [16052]));
Q_ASSIGN U16723 ( .B(clk), .A(\g.we_clk [16051]));
Q_ASSIGN U16724 ( .B(clk), .A(\g.we_clk [16050]));
Q_ASSIGN U16725 ( .B(clk), .A(\g.we_clk [16049]));
Q_ASSIGN U16726 ( .B(clk), .A(\g.we_clk [16048]));
Q_ASSIGN U16727 ( .B(clk), .A(\g.we_clk [16047]));
Q_ASSIGN U16728 ( .B(clk), .A(\g.we_clk [16046]));
Q_ASSIGN U16729 ( .B(clk), .A(\g.we_clk [16045]));
Q_ASSIGN U16730 ( .B(clk), .A(\g.we_clk [16044]));
Q_ASSIGN U16731 ( .B(clk), .A(\g.we_clk [16043]));
Q_ASSIGN U16732 ( .B(clk), .A(\g.we_clk [16042]));
Q_ASSIGN U16733 ( .B(clk), .A(\g.we_clk [16041]));
Q_ASSIGN U16734 ( .B(clk), .A(\g.we_clk [16040]));
Q_ASSIGN U16735 ( .B(clk), .A(\g.we_clk [16039]));
Q_ASSIGN U16736 ( .B(clk), .A(\g.we_clk [16038]));
Q_ASSIGN U16737 ( .B(clk), .A(\g.we_clk [16037]));
Q_ASSIGN U16738 ( .B(clk), .A(\g.we_clk [16036]));
Q_ASSIGN U16739 ( .B(clk), .A(\g.we_clk [16035]));
Q_ASSIGN U16740 ( .B(clk), .A(\g.we_clk [16034]));
Q_ASSIGN U16741 ( .B(clk), .A(\g.we_clk [16033]));
Q_ASSIGN U16742 ( .B(clk), .A(\g.we_clk [16032]));
Q_ASSIGN U16743 ( .B(clk), .A(\g.we_clk [16031]));
Q_ASSIGN U16744 ( .B(clk), .A(\g.we_clk [16030]));
Q_ASSIGN U16745 ( .B(clk), .A(\g.we_clk [16029]));
Q_ASSIGN U16746 ( .B(clk), .A(\g.we_clk [16028]));
Q_ASSIGN U16747 ( .B(clk), .A(\g.we_clk [16027]));
Q_ASSIGN U16748 ( .B(clk), .A(\g.we_clk [16026]));
Q_ASSIGN U16749 ( .B(clk), .A(\g.we_clk [16025]));
Q_ASSIGN U16750 ( .B(clk), .A(\g.we_clk [16024]));
Q_ASSIGN U16751 ( .B(clk), .A(\g.we_clk [16023]));
Q_ASSIGN U16752 ( .B(clk), .A(\g.we_clk [16022]));
Q_ASSIGN U16753 ( .B(clk), .A(\g.we_clk [16021]));
Q_ASSIGN U16754 ( .B(clk), .A(\g.we_clk [16020]));
Q_ASSIGN U16755 ( .B(clk), .A(\g.we_clk [16019]));
Q_ASSIGN U16756 ( .B(clk), .A(\g.we_clk [16018]));
Q_ASSIGN U16757 ( .B(clk), .A(\g.we_clk [16017]));
Q_ASSIGN U16758 ( .B(clk), .A(\g.we_clk [16016]));
Q_ASSIGN U16759 ( .B(clk), .A(\g.we_clk [16015]));
Q_ASSIGN U16760 ( .B(clk), .A(\g.we_clk [16014]));
Q_ASSIGN U16761 ( .B(clk), .A(\g.we_clk [16013]));
Q_ASSIGN U16762 ( .B(clk), .A(\g.we_clk [16012]));
Q_ASSIGN U16763 ( .B(clk), .A(\g.we_clk [16011]));
Q_ASSIGN U16764 ( .B(clk), .A(\g.we_clk [16010]));
Q_ASSIGN U16765 ( .B(clk), .A(\g.we_clk [16009]));
Q_ASSIGN U16766 ( .B(clk), .A(\g.we_clk [16008]));
Q_ASSIGN U16767 ( .B(clk), .A(\g.we_clk [16007]));
Q_ASSIGN U16768 ( .B(clk), .A(\g.we_clk [16006]));
Q_ASSIGN U16769 ( .B(clk), .A(\g.we_clk [16005]));
Q_ASSIGN U16770 ( .B(clk), .A(\g.we_clk [16004]));
Q_ASSIGN U16771 ( .B(clk), .A(\g.we_clk [16003]));
Q_ASSIGN U16772 ( .B(clk), .A(\g.we_clk [16002]));
Q_ASSIGN U16773 ( .B(clk), .A(\g.we_clk [16001]));
Q_ASSIGN U16774 ( .B(clk), .A(\g.we_clk [16000]));
Q_ASSIGN U16775 ( .B(clk), .A(\g.we_clk [15999]));
Q_ASSIGN U16776 ( .B(clk), .A(\g.we_clk [15998]));
Q_ASSIGN U16777 ( .B(clk), .A(\g.we_clk [15997]));
Q_ASSIGN U16778 ( .B(clk), .A(\g.we_clk [15996]));
Q_ASSIGN U16779 ( .B(clk), .A(\g.we_clk [15995]));
Q_ASSIGN U16780 ( .B(clk), .A(\g.we_clk [15994]));
Q_ASSIGN U16781 ( .B(clk), .A(\g.we_clk [15993]));
Q_ASSIGN U16782 ( .B(clk), .A(\g.we_clk [15992]));
Q_ASSIGN U16783 ( .B(clk), .A(\g.we_clk [15991]));
Q_ASSIGN U16784 ( .B(clk), .A(\g.we_clk [15990]));
Q_ASSIGN U16785 ( .B(clk), .A(\g.we_clk [15989]));
Q_ASSIGN U16786 ( .B(clk), .A(\g.we_clk [15988]));
Q_ASSIGN U16787 ( .B(clk), .A(\g.we_clk [15987]));
Q_ASSIGN U16788 ( .B(clk), .A(\g.we_clk [15986]));
Q_ASSIGN U16789 ( .B(clk), .A(\g.we_clk [15985]));
Q_ASSIGN U16790 ( .B(clk), .A(\g.we_clk [15984]));
Q_ASSIGN U16791 ( .B(clk), .A(\g.we_clk [15983]));
Q_ASSIGN U16792 ( .B(clk), .A(\g.we_clk [15982]));
Q_ASSIGN U16793 ( .B(clk), .A(\g.we_clk [15981]));
Q_ASSIGN U16794 ( .B(clk), .A(\g.we_clk [15980]));
Q_ASSIGN U16795 ( .B(clk), .A(\g.we_clk [15979]));
Q_ASSIGN U16796 ( .B(clk), .A(\g.we_clk [15978]));
Q_ASSIGN U16797 ( .B(clk), .A(\g.we_clk [15977]));
Q_ASSIGN U16798 ( .B(clk), .A(\g.we_clk [15976]));
Q_ASSIGN U16799 ( .B(clk), .A(\g.we_clk [15975]));
Q_ASSIGN U16800 ( .B(clk), .A(\g.we_clk [15974]));
Q_ASSIGN U16801 ( .B(clk), .A(\g.we_clk [15973]));
Q_ASSIGN U16802 ( .B(clk), .A(\g.we_clk [15972]));
Q_ASSIGN U16803 ( .B(clk), .A(\g.we_clk [15971]));
Q_ASSIGN U16804 ( .B(clk), .A(\g.we_clk [15970]));
Q_ASSIGN U16805 ( .B(clk), .A(\g.we_clk [15969]));
Q_ASSIGN U16806 ( .B(clk), .A(\g.we_clk [15968]));
Q_ASSIGN U16807 ( .B(clk), .A(\g.we_clk [15967]));
Q_ASSIGN U16808 ( .B(clk), .A(\g.we_clk [15966]));
Q_ASSIGN U16809 ( .B(clk), .A(\g.we_clk [15965]));
Q_ASSIGN U16810 ( .B(clk), .A(\g.we_clk [15964]));
Q_ASSIGN U16811 ( .B(clk), .A(\g.we_clk [15963]));
Q_ASSIGN U16812 ( .B(clk), .A(\g.we_clk [15962]));
Q_ASSIGN U16813 ( .B(clk), .A(\g.we_clk [15961]));
Q_ASSIGN U16814 ( .B(clk), .A(\g.we_clk [15960]));
Q_ASSIGN U16815 ( .B(clk), .A(\g.we_clk [15959]));
Q_ASSIGN U16816 ( .B(clk), .A(\g.we_clk [15958]));
Q_ASSIGN U16817 ( .B(clk), .A(\g.we_clk [15957]));
Q_ASSIGN U16818 ( .B(clk), .A(\g.we_clk [15956]));
Q_ASSIGN U16819 ( .B(clk), .A(\g.we_clk [15955]));
Q_ASSIGN U16820 ( .B(clk), .A(\g.we_clk [15954]));
Q_ASSIGN U16821 ( .B(clk), .A(\g.we_clk [15953]));
Q_ASSIGN U16822 ( .B(clk), .A(\g.we_clk [15952]));
Q_ASSIGN U16823 ( .B(clk), .A(\g.we_clk [15951]));
Q_ASSIGN U16824 ( .B(clk), .A(\g.we_clk [15950]));
Q_ASSIGN U16825 ( .B(clk), .A(\g.we_clk [15949]));
Q_ASSIGN U16826 ( .B(clk), .A(\g.we_clk [15948]));
Q_ASSIGN U16827 ( .B(clk), .A(\g.we_clk [15947]));
Q_ASSIGN U16828 ( .B(clk), .A(\g.we_clk [15946]));
Q_ASSIGN U16829 ( .B(clk), .A(\g.we_clk [15945]));
Q_ASSIGN U16830 ( .B(clk), .A(\g.we_clk [15944]));
Q_ASSIGN U16831 ( .B(clk), .A(\g.we_clk [15943]));
Q_ASSIGN U16832 ( .B(clk), .A(\g.we_clk [15942]));
Q_ASSIGN U16833 ( .B(clk), .A(\g.we_clk [15941]));
Q_ASSIGN U16834 ( .B(clk), .A(\g.we_clk [15940]));
Q_ASSIGN U16835 ( .B(clk), .A(\g.we_clk [15939]));
Q_ASSIGN U16836 ( .B(clk), .A(\g.we_clk [15938]));
Q_ASSIGN U16837 ( .B(clk), .A(\g.we_clk [15937]));
Q_ASSIGN U16838 ( .B(clk), .A(\g.we_clk [15936]));
Q_ASSIGN U16839 ( .B(clk), .A(\g.we_clk [15935]));
Q_ASSIGN U16840 ( .B(clk), .A(\g.we_clk [15934]));
Q_ASSIGN U16841 ( .B(clk), .A(\g.we_clk [15933]));
Q_ASSIGN U16842 ( .B(clk), .A(\g.we_clk [15932]));
Q_ASSIGN U16843 ( .B(clk), .A(\g.we_clk [15931]));
Q_ASSIGN U16844 ( .B(clk), .A(\g.we_clk [15930]));
Q_ASSIGN U16845 ( .B(clk), .A(\g.we_clk [15929]));
Q_ASSIGN U16846 ( .B(clk), .A(\g.we_clk [15928]));
Q_ASSIGN U16847 ( .B(clk), .A(\g.we_clk [15927]));
Q_ASSIGN U16848 ( .B(clk), .A(\g.we_clk [15926]));
Q_ASSIGN U16849 ( .B(clk), .A(\g.we_clk [15925]));
Q_ASSIGN U16850 ( .B(clk), .A(\g.we_clk [15924]));
Q_ASSIGN U16851 ( .B(clk), .A(\g.we_clk [15923]));
Q_ASSIGN U16852 ( .B(clk), .A(\g.we_clk [15922]));
Q_ASSIGN U16853 ( .B(clk), .A(\g.we_clk [15921]));
Q_ASSIGN U16854 ( .B(clk), .A(\g.we_clk [15920]));
Q_ASSIGN U16855 ( .B(clk), .A(\g.we_clk [15919]));
Q_ASSIGN U16856 ( .B(clk), .A(\g.we_clk [15918]));
Q_ASSIGN U16857 ( .B(clk), .A(\g.we_clk [15917]));
Q_ASSIGN U16858 ( .B(clk), .A(\g.we_clk [15916]));
Q_ASSIGN U16859 ( .B(clk), .A(\g.we_clk [15915]));
Q_ASSIGN U16860 ( .B(clk), .A(\g.we_clk [15914]));
Q_ASSIGN U16861 ( .B(clk), .A(\g.we_clk [15913]));
Q_ASSIGN U16862 ( .B(clk), .A(\g.we_clk [15912]));
Q_ASSIGN U16863 ( .B(clk), .A(\g.we_clk [15911]));
Q_ASSIGN U16864 ( .B(clk), .A(\g.we_clk [15910]));
Q_ASSIGN U16865 ( .B(clk), .A(\g.we_clk [15909]));
Q_ASSIGN U16866 ( .B(clk), .A(\g.we_clk [15908]));
Q_ASSIGN U16867 ( .B(clk), .A(\g.we_clk [15907]));
Q_ASSIGN U16868 ( .B(clk), .A(\g.we_clk [15906]));
Q_ASSIGN U16869 ( .B(clk), .A(\g.we_clk [15905]));
Q_ASSIGN U16870 ( .B(clk), .A(\g.we_clk [15904]));
Q_ASSIGN U16871 ( .B(clk), .A(\g.we_clk [15903]));
Q_ASSIGN U16872 ( .B(clk), .A(\g.we_clk [15902]));
Q_ASSIGN U16873 ( .B(clk), .A(\g.we_clk [15901]));
Q_ASSIGN U16874 ( .B(clk), .A(\g.we_clk [15900]));
Q_ASSIGN U16875 ( .B(clk), .A(\g.we_clk [15899]));
Q_ASSIGN U16876 ( .B(clk), .A(\g.we_clk [15898]));
Q_ASSIGN U16877 ( .B(clk), .A(\g.we_clk [15897]));
Q_ASSIGN U16878 ( .B(clk), .A(\g.we_clk [15896]));
Q_ASSIGN U16879 ( .B(clk), .A(\g.we_clk [15895]));
Q_ASSIGN U16880 ( .B(clk), .A(\g.we_clk [15894]));
Q_ASSIGN U16881 ( .B(clk), .A(\g.we_clk [15893]));
Q_ASSIGN U16882 ( .B(clk), .A(\g.we_clk [15892]));
Q_ASSIGN U16883 ( .B(clk), .A(\g.we_clk [15891]));
Q_ASSIGN U16884 ( .B(clk), .A(\g.we_clk [15890]));
Q_ASSIGN U16885 ( .B(clk), .A(\g.we_clk [15889]));
Q_ASSIGN U16886 ( .B(clk), .A(\g.we_clk [15888]));
Q_ASSIGN U16887 ( .B(clk), .A(\g.we_clk [15887]));
Q_ASSIGN U16888 ( .B(clk), .A(\g.we_clk [15886]));
Q_ASSIGN U16889 ( .B(clk), .A(\g.we_clk [15885]));
Q_ASSIGN U16890 ( .B(clk), .A(\g.we_clk [15884]));
Q_ASSIGN U16891 ( .B(clk), .A(\g.we_clk [15883]));
Q_ASSIGN U16892 ( .B(clk), .A(\g.we_clk [15882]));
Q_ASSIGN U16893 ( .B(clk), .A(\g.we_clk [15881]));
Q_ASSIGN U16894 ( .B(clk), .A(\g.we_clk [15880]));
Q_ASSIGN U16895 ( .B(clk), .A(\g.we_clk [15879]));
Q_ASSIGN U16896 ( .B(clk), .A(\g.we_clk [15878]));
Q_ASSIGN U16897 ( .B(clk), .A(\g.we_clk [15877]));
Q_ASSIGN U16898 ( .B(clk), .A(\g.we_clk [15876]));
Q_ASSIGN U16899 ( .B(clk), .A(\g.we_clk [15875]));
Q_ASSIGN U16900 ( .B(clk), .A(\g.we_clk [15874]));
Q_ASSIGN U16901 ( .B(clk), .A(\g.we_clk [15873]));
Q_ASSIGN U16902 ( .B(clk), .A(\g.we_clk [15872]));
Q_ASSIGN U16903 ( .B(clk), .A(\g.we_clk [15871]));
Q_ASSIGN U16904 ( .B(clk), .A(\g.we_clk [15870]));
Q_ASSIGN U16905 ( .B(clk), .A(\g.we_clk [15869]));
Q_ASSIGN U16906 ( .B(clk), .A(\g.we_clk [15868]));
Q_ASSIGN U16907 ( .B(clk), .A(\g.we_clk [15867]));
Q_ASSIGN U16908 ( .B(clk), .A(\g.we_clk [15866]));
Q_ASSIGN U16909 ( .B(clk), .A(\g.we_clk [15865]));
Q_ASSIGN U16910 ( .B(clk), .A(\g.we_clk [15864]));
Q_ASSIGN U16911 ( .B(clk), .A(\g.we_clk [15863]));
Q_ASSIGN U16912 ( .B(clk), .A(\g.we_clk [15862]));
Q_ASSIGN U16913 ( .B(clk), .A(\g.we_clk [15861]));
Q_ASSIGN U16914 ( .B(clk), .A(\g.we_clk [15860]));
Q_ASSIGN U16915 ( .B(clk), .A(\g.we_clk [15859]));
Q_ASSIGN U16916 ( .B(clk), .A(\g.we_clk [15858]));
Q_ASSIGN U16917 ( .B(clk), .A(\g.we_clk [15857]));
Q_ASSIGN U16918 ( .B(clk), .A(\g.we_clk [15856]));
Q_ASSIGN U16919 ( .B(clk), .A(\g.we_clk [15855]));
Q_ASSIGN U16920 ( .B(clk), .A(\g.we_clk [15854]));
Q_ASSIGN U16921 ( .B(clk), .A(\g.we_clk [15853]));
Q_ASSIGN U16922 ( .B(clk), .A(\g.we_clk [15852]));
Q_ASSIGN U16923 ( .B(clk), .A(\g.we_clk [15851]));
Q_ASSIGN U16924 ( .B(clk), .A(\g.we_clk [15850]));
Q_ASSIGN U16925 ( .B(clk), .A(\g.we_clk [15849]));
Q_ASSIGN U16926 ( .B(clk), .A(\g.we_clk [15848]));
Q_ASSIGN U16927 ( .B(clk), .A(\g.we_clk [15847]));
Q_ASSIGN U16928 ( .B(clk), .A(\g.we_clk [15846]));
Q_ASSIGN U16929 ( .B(clk), .A(\g.we_clk [15845]));
Q_ASSIGN U16930 ( .B(clk), .A(\g.we_clk [15844]));
Q_ASSIGN U16931 ( .B(clk), .A(\g.we_clk [15843]));
Q_ASSIGN U16932 ( .B(clk), .A(\g.we_clk [15842]));
Q_ASSIGN U16933 ( .B(clk), .A(\g.we_clk [15841]));
Q_ASSIGN U16934 ( .B(clk), .A(\g.we_clk [15840]));
Q_ASSIGN U16935 ( .B(clk), .A(\g.we_clk [15839]));
Q_ASSIGN U16936 ( .B(clk), .A(\g.we_clk [15838]));
Q_ASSIGN U16937 ( .B(clk), .A(\g.we_clk [15837]));
Q_ASSIGN U16938 ( .B(clk), .A(\g.we_clk [15836]));
Q_ASSIGN U16939 ( .B(clk), .A(\g.we_clk [15835]));
Q_ASSIGN U16940 ( .B(clk), .A(\g.we_clk [15834]));
Q_ASSIGN U16941 ( .B(clk), .A(\g.we_clk [15833]));
Q_ASSIGN U16942 ( .B(clk), .A(\g.we_clk [15832]));
Q_ASSIGN U16943 ( .B(clk), .A(\g.we_clk [15831]));
Q_ASSIGN U16944 ( .B(clk), .A(\g.we_clk [15830]));
Q_ASSIGN U16945 ( .B(clk), .A(\g.we_clk [15829]));
Q_ASSIGN U16946 ( .B(clk), .A(\g.we_clk [15828]));
Q_ASSIGN U16947 ( .B(clk), .A(\g.we_clk [15827]));
Q_ASSIGN U16948 ( .B(clk), .A(\g.we_clk [15826]));
Q_ASSIGN U16949 ( .B(clk), .A(\g.we_clk [15825]));
Q_ASSIGN U16950 ( .B(clk), .A(\g.we_clk [15824]));
Q_ASSIGN U16951 ( .B(clk), .A(\g.we_clk [15823]));
Q_ASSIGN U16952 ( .B(clk), .A(\g.we_clk [15822]));
Q_ASSIGN U16953 ( .B(clk), .A(\g.we_clk [15821]));
Q_ASSIGN U16954 ( .B(clk), .A(\g.we_clk [15820]));
Q_ASSIGN U16955 ( .B(clk), .A(\g.we_clk [15819]));
Q_ASSIGN U16956 ( .B(clk), .A(\g.we_clk [15818]));
Q_ASSIGN U16957 ( .B(clk), .A(\g.we_clk [15817]));
Q_ASSIGN U16958 ( .B(clk), .A(\g.we_clk [15816]));
Q_ASSIGN U16959 ( .B(clk), .A(\g.we_clk [15815]));
Q_ASSIGN U16960 ( .B(clk), .A(\g.we_clk [15814]));
Q_ASSIGN U16961 ( .B(clk), .A(\g.we_clk [15813]));
Q_ASSIGN U16962 ( .B(clk), .A(\g.we_clk [15812]));
Q_ASSIGN U16963 ( .B(clk), .A(\g.we_clk [15811]));
Q_ASSIGN U16964 ( .B(clk), .A(\g.we_clk [15810]));
Q_ASSIGN U16965 ( .B(clk), .A(\g.we_clk [15809]));
Q_ASSIGN U16966 ( .B(clk), .A(\g.we_clk [15808]));
Q_ASSIGN U16967 ( .B(clk), .A(\g.we_clk [15807]));
Q_ASSIGN U16968 ( .B(clk), .A(\g.we_clk [15806]));
Q_ASSIGN U16969 ( .B(clk), .A(\g.we_clk [15805]));
Q_ASSIGN U16970 ( .B(clk), .A(\g.we_clk [15804]));
Q_ASSIGN U16971 ( .B(clk), .A(\g.we_clk [15803]));
Q_ASSIGN U16972 ( .B(clk), .A(\g.we_clk [15802]));
Q_ASSIGN U16973 ( .B(clk), .A(\g.we_clk [15801]));
Q_ASSIGN U16974 ( .B(clk), .A(\g.we_clk [15800]));
Q_ASSIGN U16975 ( .B(clk), .A(\g.we_clk [15799]));
Q_ASSIGN U16976 ( .B(clk), .A(\g.we_clk [15798]));
Q_ASSIGN U16977 ( .B(clk), .A(\g.we_clk [15797]));
Q_ASSIGN U16978 ( .B(clk), .A(\g.we_clk [15796]));
Q_ASSIGN U16979 ( .B(clk), .A(\g.we_clk [15795]));
Q_ASSIGN U16980 ( .B(clk), .A(\g.we_clk [15794]));
Q_ASSIGN U16981 ( .B(clk), .A(\g.we_clk [15793]));
Q_ASSIGN U16982 ( .B(clk), .A(\g.we_clk [15792]));
Q_ASSIGN U16983 ( .B(clk), .A(\g.we_clk [15791]));
Q_ASSIGN U16984 ( .B(clk), .A(\g.we_clk [15790]));
Q_ASSIGN U16985 ( .B(clk), .A(\g.we_clk [15789]));
Q_ASSIGN U16986 ( .B(clk), .A(\g.we_clk [15788]));
Q_ASSIGN U16987 ( .B(clk), .A(\g.we_clk [15787]));
Q_ASSIGN U16988 ( .B(clk), .A(\g.we_clk [15786]));
Q_ASSIGN U16989 ( .B(clk), .A(\g.we_clk [15785]));
Q_ASSIGN U16990 ( .B(clk), .A(\g.we_clk [15784]));
Q_ASSIGN U16991 ( .B(clk), .A(\g.we_clk [15783]));
Q_ASSIGN U16992 ( .B(clk), .A(\g.we_clk [15782]));
Q_ASSIGN U16993 ( .B(clk), .A(\g.we_clk [15781]));
Q_ASSIGN U16994 ( .B(clk), .A(\g.we_clk [15780]));
Q_ASSIGN U16995 ( .B(clk), .A(\g.we_clk [15779]));
Q_ASSIGN U16996 ( .B(clk), .A(\g.we_clk [15778]));
Q_ASSIGN U16997 ( .B(clk), .A(\g.we_clk [15777]));
Q_ASSIGN U16998 ( .B(clk), .A(\g.we_clk [15776]));
Q_ASSIGN U16999 ( .B(clk), .A(\g.we_clk [15775]));
Q_ASSIGN U17000 ( .B(clk), .A(\g.we_clk [15774]));
Q_ASSIGN U17001 ( .B(clk), .A(\g.we_clk [15773]));
Q_ASSIGN U17002 ( .B(clk), .A(\g.we_clk [15772]));
Q_ASSIGN U17003 ( .B(clk), .A(\g.we_clk [15771]));
Q_ASSIGN U17004 ( .B(clk), .A(\g.we_clk [15770]));
Q_ASSIGN U17005 ( .B(clk), .A(\g.we_clk [15769]));
Q_ASSIGN U17006 ( .B(clk), .A(\g.we_clk [15768]));
Q_ASSIGN U17007 ( .B(clk), .A(\g.we_clk [15767]));
Q_ASSIGN U17008 ( .B(clk), .A(\g.we_clk [15766]));
Q_ASSIGN U17009 ( .B(clk), .A(\g.we_clk [15765]));
Q_ASSIGN U17010 ( .B(clk), .A(\g.we_clk [15764]));
Q_ASSIGN U17011 ( .B(clk), .A(\g.we_clk [15763]));
Q_ASSIGN U17012 ( .B(clk), .A(\g.we_clk [15762]));
Q_ASSIGN U17013 ( .B(clk), .A(\g.we_clk [15761]));
Q_ASSIGN U17014 ( .B(clk), .A(\g.we_clk [15760]));
Q_ASSIGN U17015 ( .B(clk), .A(\g.we_clk [15759]));
Q_ASSIGN U17016 ( .B(clk), .A(\g.we_clk [15758]));
Q_ASSIGN U17017 ( .B(clk), .A(\g.we_clk [15757]));
Q_ASSIGN U17018 ( .B(clk), .A(\g.we_clk [15756]));
Q_ASSIGN U17019 ( .B(clk), .A(\g.we_clk [15755]));
Q_ASSIGN U17020 ( .B(clk), .A(\g.we_clk [15754]));
Q_ASSIGN U17021 ( .B(clk), .A(\g.we_clk [15753]));
Q_ASSIGN U17022 ( .B(clk), .A(\g.we_clk [15752]));
Q_ASSIGN U17023 ( .B(clk), .A(\g.we_clk [15751]));
Q_ASSIGN U17024 ( .B(clk), .A(\g.we_clk [15750]));
Q_ASSIGN U17025 ( .B(clk), .A(\g.we_clk [15749]));
Q_ASSIGN U17026 ( .B(clk), .A(\g.we_clk [15748]));
Q_ASSIGN U17027 ( .B(clk), .A(\g.we_clk [15747]));
Q_ASSIGN U17028 ( .B(clk), .A(\g.we_clk [15746]));
Q_ASSIGN U17029 ( .B(clk), .A(\g.we_clk [15745]));
Q_ASSIGN U17030 ( .B(clk), .A(\g.we_clk [15744]));
Q_ASSIGN U17031 ( .B(clk), .A(\g.we_clk [15743]));
Q_ASSIGN U17032 ( .B(clk), .A(\g.we_clk [15742]));
Q_ASSIGN U17033 ( .B(clk), .A(\g.we_clk [15741]));
Q_ASSIGN U17034 ( .B(clk), .A(\g.we_clk [15740]));
Q_ASSIGN U17035 ( .B(clk), .A(\g.we_clk [15739]));
Q_ASSIGN U17036 ( .B(clk), .A(\g.we_clk [15738]));
Q_ASSIGN U17037 ( .B(clk), .A(\g.we_clk [15737]));
Q_ASSIGN U17038 ( .B(clk), .A(\g.we_clk [15736]));
Q_ASSIGN U17039 ( .B(clk), .A(\g.we_clk [15735]));
Q_ASSIGN U17040 ( .B(clk), .A(\g.we_clk [15734]));
Q_ASSIGN U17041 ( .B(clk), .A(\g.we_clk [15733]));
Q_ASSIGN U17042 ( .B(clk), .A(\g.we_clk [15732]));
Q_ASSIGN U17043 ( .B(clk), .A(\g.we_clk [15731]));
Q_ASSIGN U17044 ( .B(clk), .A(\g.we_clk [15730]));
Q_ASSIGN U17045 ( .B(clk), .A(\g.we_clk [15729]));
Q_ASSIGN U17046 ( .B(clk), .A(\g.we_clk [15728]));
Q_ASSIGN U17047 ( .B(clk), .A(\g.we_clk [15727]));
Q_ASSIGN U17048 ( .B(clk), .A(\g.we_clk [15726]));
Q_ASSIGN U17049 ( .B(clk), .A(\g.we_clk [15725]));
Q_ASSIGN U17050 ( .B(clk), .A(\g.we_clk [15724]));
Q_ASSIGN U17051 ( .B(clk), .A(\g.we_clk [15723]));
Q_ASSIGN U17052 ( .B(clk), .A(\g.we_clk [15722]));
Q_ASSIGN U17053 ( .B(clk), .A(\g.we_clk [15721]));
Q_ASSIGN U17054 ( .B(clk), .A(\g.we_clk [15720]));
Q_ASSIGN U17055 ( .B(clk), .A(\g.we_clk [15719]));
Q_ASSIGN U17056 ( .B(clk), .A(\g.we_clk [15718]));
Q_ASSIGN U17057 ( .B(clk), .A(\g.we_clk [15717]));
Q_ASSIGN U17058 ( .B(clk), .A(\g.we_clk [15716]));
Q_ASSIGN U17059 ( .B(clk), .A(\g.we_clk [15715]));
Q_ASSIGN U17060 ( .B(clk), .A(\g.we_clk [15714]));
Q_ASSIGN U17061 ( .B(clk), .A(\g.we_clk [15713]));
Q_ASSIGN U17062 ( .B(clk), .A(\g.we_clk [15712]));
Q_ASSIGN U17063 ( .B(clk), .A(\g.we_clk [15711]));
Q_ASSIGN U17064 ( .B(clk), .A(\g.we_clk [15710]));
Q_ASSIGN U17065 ( .B(clk), .A(\g.we_clk [15709]));
Q_ASSIGN U17066 ( .B(clk), .A(\g.we_clk [15708]));
Q_ASSIGN U17067 ( .B(clk), .A(\g.we_clk [15707]));
Q_ASSIGN U17068 ( .B(clk), .A(\g.we_clk [15706]));
Q_ASSIGN U17069 ( .B(clk), .A(\g.we_clk [15705]));
Q_ASSIGN U17070 ( .B(clk), .A(\g.we_clk [15704]));
Q_ASSIGN U17071 ( .B(clk), .A(\g.we_clk [15703]));
Q_ASSIGN U17072 ( .B(clk), .A(\g.we_clk [15702]));
Q_ASSIGN U17073 ( .B(clk), .A(\g.we_clk [15701]));
Q_ASSIGN U17074 ( .B(clk), .A(\g.we_clk [15700]));
Q_ASSIGN U17075 ( .B(clk), .A(\g.we_clk [15699]));
Q_ASSIGN U17076 ( .B(clk), .A(\g.we_clk [15698]));
Q_ASSIGN U17077 ( .B(clk), .A(\g.we_clk [15697]));
Q_ASSIGN U17078 ( .B(clk), .A(\g.we_clk [15696]));
Q_ASSIGN U17079 ( .B(clk), .A(\g.we_clk [15695]));
Q_ASSIGN U17080 ( .B(clk), .A(\g.we_clk [15694]));
Q_ASSIGN U17081 ( .B(clk), .A(\g.we_clk [15693]));
Q_ASSIGN U17082 ( .B(clk), .A(\g.we_clk [15692]));
Q_ASSIGN U17083 ( .B(clk), .A(\g.we_clk [15691]));
Q_ASSIGN U17084 ( .B(clk), .A(\g.we_clk [15690]));
Q_ASSIGN U17085 ( .B(clk), .A(\g.we_clk [15689]));
Q_ASSIGN U17086 ( .B(clk), .A(\g.we_clk [15688]));
Q_ASSIGN U17087 ( .B(clk), .A(\g.we_clk [15687]));
Q_ASSIGN U17088 ( .B(clk), .A(\g.we_clk [15686]));
Q_ASSIGN U17089 ( .B(clk), .A(\g.we_clk [15685]));
Q_ASSIGN U17090 ( .B(clk), .A(\g.we_clk [15684]));
Q_ASSIGN U17091 ( .B(clk), .A(\g.we_clk [15683]));
Q_ASSIGN U17092 ( .B(clk), .A(\g.we_clk [15682]));
Q_ASSIGN U17093 ( .B(clk), .A(\g.we_clk [15681]));
Q_ASSIGN U17094 ( .B(clk), .A(\g.we_clk [15680]));
Q_ASSIGN U17095 ( .B(clk), .A(\g.we_clk [15679]));
Q_ASSIGN U17096 ( .B(clk), .A(\g.we_clk [15678]));
Q_ASSIGN U17097 ( .B(clk), .A(\g.we_clk [15677]));
Q_ASSIGN U17098 ( .B(clk), .A(\g.we_clk [15676]));
Q_ASSIGN U17099 ( .B(clk), .A(\g.we_clk [15675]));
Q_ASSIGN U17100 ( .B(clk), .A(\g.we_clk [15674]));
Q_ASSIGN U17101 ( .B(clk), .A(\g.we_clk [15673]));
Q_ASSIGN U17102 ( .B(clk), .A(\g.we_clk [15672]));
Q_ASSIGN U17103 ( .B(clk), .A(\g.we_clk [15671]));
Q_ASSIGN U17104 ( .B(clk), .A(\g.we_clk [15670]));
Q_ASSIGN U17105 ( .B(clk), .A(\g.we_clk [15669]));
Q_ASSIGN U17106 ( .B(clk), .A(\g.we_clk [15668]));
Q_ASSIGN U17107 ( .B(clk), .A(\g.we_clk [15667]));
Q_ASSIGN U17108 ( .B(clk), .A(\g.we_clk [15666]));
Q_ASSIGN U17109 ( .B(clk), .A(\g.we_clk [15665]));
Q_ASSIGN U17110 ( .B(clk), .A(\g.we_clk [15664]));
Q_ASSIGN U17111 ( .B(clk), .A(\g.we_clk [15663]));
Q_ASSIGN U17112 ( .B(clk), .A(\g.we_clk [15662]));
Q_ASSIGN U17113 ( .B(clk), .A(\g.we_clk [15661]));
Q_ASSIGN U17114 ( .B(clk), .A(\g.we_clk [15660]));
Q_ASSIGN U17115 ( .B(clk), .A(\g.we_clk [15659]));
Q_ASSIGN U17116 ( .B(clk), .A(\g.we_clk [15658]));
Q_ASSIGN U17117 ( .B(clk), .A(\g.we_clk [15657]));
Q_ASSIGN U17118 ( .B(clk), .A(\g.we_clk [15656]));
Q_ASSIGN U17119 ( .B(clk), .A(\g.we_clk [15655]));
Q_ASSIGN U17120 ( .B(clk), .A(\g.we_clk [15654]));
Q_ASSIGN U17121 ( .B(clk), .A(\g.we_clk [15653]));
Q_ASSIGN U17122 ( .B(clk), .A(\g.we_clk [15652]));
Q_ASSIGN U17123 ( .B(clk), .A(\g.we_clk [15651]));
Q_ASSIGN U17124 ( .B(clk), .A(\g.we_clk [15650]));
Q_ASSIGN U17125 ( .B(clk), .A(\g.we_clk [15649]));
Q_ASSIGN U17126 ( .B(clk), .A(\g.we_clk [15648]));
Q_ASSIGN U17127 ( .B(clk), .A(\g.we_clk [15647]));
Q_ASSIGN U17128 ( .B(clk), .A(\g.we_clk [15646]));
Q_ASSIGN U17129 ( .B(clk), .A(\g.we_clk [15645]));
Q_ASSIGN U17130 ( .B(clk), .A(\g.we_clk [15644]));
Q_ASSIGN U17131 ( .B(clk), .A(\g.we_clk [15643]));
Q_ASSIGN U17132 ( .B(clk), .A(\g.we_clk [15642]));
Q_ASSIGN U17133 ( .B(clk), .A(\g.we_clk [15641]));
Q_ASSIGN U17134 ( .B(clk), .A(\g.we_clk [15640]));
Q_ASSIGN U17135 ( .B(clk), .A(\g.we_clk [15639]));
Q_ASSIGN U17136 ( .B(clk), .A(\g.we_clk [15638]));
Q_ASSIGN U17137 ( .B(clk), .A(\g.we_clk [15637]));
Q_ASSIGN U17138 ( .B(clk), .A(\g.we_clk [15636]));
Q_ASSIGN U17139 ( .B(clk), .A(\g.we_clk [15635]));
Q_ASSIGN U17140 ( .B(clk), .A(\g.we_clk [15634]));
Q_ASSIGN U17141 ( .B(clk), .A(\g.we_clk [15633]));
Q_ASSIGN U17142 ( .B(clk), .A(\g.we_clk [15632]));
Q_ASSIGN U17143 ( .B(clk), .A(\g.we_clk [15631]));
Q_ASSIGN U17144 ( .B(clk), .A(\g.we_clk [15630]));
Q_ASSIGN U17145 ( .B(clk), .A(\g.we_clk [15629]));
Q_ASSIGN U17146 ( .B(clk), .A(\g.we_clk [15628]));
Q_ASSIGN U17147 ( .B(clk), .A(\g.we_clk [15627]));
Q_ASSIGN U17148 ( .B(clk), .A(\g.we_clk [15626]));
Q_ASSIGN U17149 ( .B(clk), .A(\g.we_clk [15625]));
Q_ASSIGN U17150 ( .B(clk), .A(\g.we_clk [15624]));
Q_ASSIGN U17151 ( .B(clk), .A(\g.we_clk [15623]));
Q_ASSIGN U17152 ( .B(clk), .A(\g.we_clk [15622]));
Q_ASSIGN U17153 ( .B(clk), .A(\g.we_clk [15621]));
Q_ASSIGN U17154 ( .B(clk), .A(\g.we_clk [15620]));
Q_ASSIGN U17155 ( .B(clk), .A(\g.we_clk [15619]));
Q_ASSIGN U17156 ( .B(clk), .A(\g.we_clk [15618]));
Q_ASSIGN U17157 ( .B(clk), .A(\g.we_clk [15617]));
Q_ASSIGN U17158 ( .B(clk), .A(\g.we_clk [15616]));
Q_ASSIGN U17159 ( .B(clk), .A(\g.we_clk [15615]));
Q_ASSIGN U17160 ( .B(clk), .A(\g.we_clk [15614]));
Q_ASSIGN U17161 ( .B(clk), .A(\g.we_clk [15613]));
Q_ASSIGN U17162 ( .B(clk), .A(\g.we_clk [15612]));
Q_ASSIGN U17163 ( .B(clk), .A(\g.we_clk [15611]));
Q_ASSIGN U17164 ( .B(clk), .A(\g.we_clk [15610]));
Q_ASSIGN U17165 ( .B(clk), .A(\g.we_clk [15609]));
Q_ASSIGN U17166 ( .B(clk), .A(\g.we_clk [15608]));
Q_ASSIGN U17167 ( .B(clk), .A(\g.we_clk [15607]));
Q_ASSIGN U17168 ( .B(clk), .A(\g.we_clk [15606]));
Q_ASSIGN U17169 ( .B(clk), .A(\g.we_clk [15605]));
Q_ASSIGN U17170 ( .B(clk), .A(\g.we_clk [15604]));
Q_ASSIGN U17171 ( .B(clk), .A(\g.we_clk [15603]));
Q_ASSIGN U17172 ( .B(clk), .A(\g.we_clk [15602]));
Q_ASSIGN U17173 ( .B(clk), .A(\g.we_clk [15601]));
Q_ASSIGN U17174 ( .B(clk), .A(\g.we_clk [15600]));
Q_ASSIGN U17175 ( .B(clk), .A(\g.we_clk [15599]));
Q_ASSIGN U17176 ( .B(clk), .A(\g.we_clk [15598]));
Q_ASSIGN U17177 ( .B(clk), .A(\g.we_clk [15597]));
Q_ASSIGN U17178 ( .B(clk), .A(\g.we_clk [15596]));
Q_ASSIGN U17179 ( .B(clk), .A(\g.we_clk [15595]));
Q_ASSIGN U17180 ( .B(clk), .A(\g.we_clk [15594]));
Q_ASSIGN U17181 ( .B(clk), .A(\g.we_clk [15593]));
Q_ASSIGN U17182 ( .B(clk), .A(\g.we_clk [15592]));
Q_ASSIGN U17183 ( .B(clk), .A(\g.we_clk [15591]));
Q_ASSIGN U17184 ( .B(clk), .A(\g.we_clk [15590]));
Q_ASSIGN U17185 ( .B(clk), .A(\g.we_clk [15589]));
Q_ASSIGN U17186 ( .B(clk), .A(\g.we_clk [15588]));
Q_ASSIGN U17187 ( .B(clk), .A(\g.we_clk [15587]));
Q_ASSIGN U17188 ( .B(clk), .A(\g.we_clk [15586]));
Q_ASSIGN U17189 ( .B(clk), .A(\g.we_clk [15585]));
Q_ASSIGN U17190 ( .B(clk), .A(\g.we_clk [15584]));
Q_ASSIGN U17191 ( .B(clk), .A(\g.we_clk [15583]));
Q_ASSIGN U17192 ( .B(clk), .A(\g.we_clk [15582]));
Q_ASSIGN U17193 ( .B(clk), .A(\g.we_clk [15581]));
Q_ASSIGN U17194 ( .B(clk), .A(\g.we_clk [15580]));
Q_ASSIGN U17195 ( .B(clk), .A(\g.we_clk [15579]));
Q_ASSIGN U17196 ( .B(clk), .A(\g.we_clk [15578]));
Q_ASSIGN U17197 ( .B(clk), .A(\g.we_clk [15577]));
Q_ASSIGN U17198 ( .B(clk), .A(\g.we_clk [15576]));
Q_ASSIGN U17199 ( .B(clk), .A(\g.we_clk [15575]));
Q_ASSIGN U17200 ( .B(clk), .A(\g.we_clk [15574]));
Q_ASSIGN U17201 ( .B(clk), .A(\g.we_clk [15573]));
Q_ASSIGN U17202 ( .B(clk), .A(\g.we_clk [15572]));
Q_ASSIGN U17203 ( .B(clk), .A(\g.we_clk [15571]));
Q_ASSIGN U17204 ( .B(clk), .A(\g.we_clk [15570]));
Q_ASSIGN U17205 ( .B(clk), .A(\g.we_clk [15569]));
Q_ASSIGN U17206 ( .B(clk), .A(\g.we_clk [15568]));
Q_ASSIGN U17207 ( .B(clk), .A(\g.we_clk [15567]));
Q_ASSIGN U17208 ( .B(clk), .A(\g.we_clk [15566]));
Q_ASSIGN U17209 ( .B(clk), .A(\g.we_clk [15565]));
Q_ASSIGN U17210 ( .B(clk), .A(\g.we_clk [15564]));
Q_ASSIGN U17211 ( .B(clk), .A(\g.we_clk [15563]));
Q_ASSIGN U17212 ( .B(clk), .A(\g.we_clk [15562]));
Q_ASSIGN U17213 ( .B(clk), .A(\g.we_clk [15561]));
Q_ASSIGN U17214 ( .B(clk), .A(\g.we_clk [15560]));
Q_ASSIGN U17215 ( .B(clk), .A(\g.we_clk [15559]));
Q_ASSIGN U17216 ( .B(clk), .A(\g.we_clk [15558]));
Q_ASSIGN U17217 ( .B(clk), .A(\g.we_clk [15557]));
Q_ASSIGN U17218 ( .B(clk), .A(\g.we_clk [15556]));
Q_ASSIGN U17219 ( .B(clk), .A(\g.we_clk [15555]));
Q_ASSIGN U17220 ( .B(clk), .A(\g.we_clk [15554]));
Q_ASSIGN U17221 ( .B(clk), .A(\g.we_clk [15553]));
Q_ASSIGN U17222 ( .B(clk), .A(\g.we_clk [15552]));
Q_ASSIGN U17223 ( .B(clk), .A(\g.we_clk [15551]));
Q_ASSIGN U17224 ( .B(clk), .A(\g.we_clk [15550]));
Q_ASSIGN U17225 ( .B(clk), .A(\g.we_clk [15549]));
Q_ASSIGN U17226 ( .B(clk), .A(\g.we_clk [15548]));
Q_ASSIGN U17227 ( .B(clk), .A(\g.we_clk [15547]));
Q_ASSIGN U17228 ( .B(clk), .A(\g.we_clk [15546]));
Q_ASSIGN U17229 ( .B(clk), .A(\g.we_clk [15545]));
Q_ASSIGN U17230 ( .B(clk), .A(\g.we_clk [15544]));
Q_ASSIGN U17231 ( .B(clk), .A(\g.we_clk [15543]));
Q_ASSIGN U17232 ( .B(clk), .A(\g.we_clk [15542]));
Q_ASSIGN U17233 ( .B(clk), .A(\g.we_clk [15541]));
Q_ASSIGN U17234 ( .B(clk), .A(\g.we_clk [15540]));
Q_ASSIGN U17235 ( .B(clk), .A(\g.we_clk [15539]));
Q_ASSIGN U17236 ( .B(clk), .A(\g.we_clk [15538]));
Q_ASSIGN U17237 ( .B(clk), .A(\g.we_clk [15537]));
Q_ASSIGN U17238 ( .B(clk), .A(\g.we_clk [15536]));
Q_ASSIGN U17239 ( .B(clk), .A(\g.we_clk [15535]));
Q_ASSIGN U17240 ( .B(clk), .A(\g.we_clk [15534]));
Q_ASSIGN U17241 ( .B(clk), .A(\g.we_clk [15533]));
Q_ASSIGN U17242 ( .B(clk), .A(\g.we_clk [15532]));
Q_ASSIGN U17243 ( .B(clk), .A(\g.we_clk [15531]));
Q_ASSIGN U17244 ( .B(clk), .A(\g.we_clk [15530]));
Q_ASSIGN U17245 ( .B(clk), .A(\g.we_clk [15529]));
Q_ASSIGN U17246 ( .B(clk), .A(\g.we_clk [15528]));
Q_ASSIGN U17247 ( .B(clk), .A(\g.we_clk [15527]));
Q_ASSIGN U17248 ( .B(clk), .A(\g.we_clk [15526]));
Q_ASSIGN U17249 ( .B(clk), .A(\g.we_clk [15525]));
Q_ASSIGN U17250 ( .B(clk), .A(\g.we_clk [15524]));
Q_ASSIGN U17251 ( .B(clk), .A(\g.we_clk [15523]));
Q_ASSIGN U17252 ( .B(clk), .A(\g.we_clk [15522]));
Q_ASSIGN U17253 ( .B(clk), .A(\g.we_clk [15521]));
Q_ASSIGN U17254 ( .B(clk), .A(\g.we_clk [15520]));
Q_ASSIGN U17255 ( .B(clk), .A(\g.we_clk [15519]));
Q_ASSIGN U17256 ( .B(clk), .A(\g.we_clk [15518]));
Q_ASSIGN U17257 ( .B(clk), .A(\g.we_clk [15517]));
Q_ASSIGN U17258 ( .B(clk), .A(\g.we_clk [15516]));
Q_ASSIGN U17259 ( .B(clk), .A(\g.we_clk [15515]));
Q_ASSIGN U17260 ( .B(clk), .A(\g.we_clk [15514]));
Q_ASSIGN U17261 ( .B(clk), .A(\g.we_clk [15513]));
Q_ASSIGN U17262 ( .B(clk), .A(\g.we_clk [15512]));
Q_ASSIGN U17263 ( .B(clk), .A(\g.we_clk [15511]));
Q_ASSIGN U17264 ( .B(clk), .A(\g.we_clk [15510]));
Q_ASSIGN U17265 ( .B(clk), .A(\g.we_clk [15509]));
Q_ASSIGN U17266 ( .B(clk), .A(\g.we_clk [15508]));
Q_ASSIGN U17267 ( .B(clk), .A(\g.we_clk [15507]));
Q_ASSIGN U17268 ( .B(clk), .A(\g.we_clk [15506]));
Q_ASSIGN U17269 ( .B(clk), .A(\g.we_clk [15505]));
Q_ASSIGN U17270 ( .B(clk), .A(\g.we_clk [15504]));
Q_ASSIGN U17271 ( .B(clk), .A(\g.we_clk [15503]));
Q_ASSIGN U17272 ( .B(clk), .A(\g.we_clk [15502]));
Q_ASSIGN U17273 ( .B(clk), .A(\g.we_clk [15501]));
Q_ASSIGN U17274 ( .B(clk), .A(\g.we_clk [15500]));
Q_ASSIGN U17275 ( .B(clk), .A(\g.we_clk [15499]));
Q_ASSIGN U17276 ( .B(clk), .A(\g.we_clk [15498]));
Q_ASSIGN U17277 ( .B(clk), .A(\g.we_clk [15497]));
Q_ASSIGN U17278 ( .B(clk), .A(\g.we_clk [15496]));
Q_ASSIGN U17279 ( .B(clk), .A(\g.we_clk [15495]));
Q_ASSIGN U17280 ( .B(clk), .A(\g.we_clk [15494]));
Q_ASSIGN U17281 ( .B(clk), .A(\g.we_clk [15493]));
Q_ASSIGN U17282 ( .B(clk), .A(\g.we_clk [15492]));
Q_ASSIGN U17283 ( .B(clk), .A(\g.we_clk [15491]));
Q_ASSIGN U17284 ( .B(clk), .A(\g.we_clk [15490]));
Q_ASSIGN U17285 ( .B(clk), .A(\g.we_clk [15489]));
Q_ASSIGN U17286 ( .B(clk), .A(\g.we_clk [15488]));
Q_ASSIGN U17287 ( .B(clk), .A(\g.we_clk [15487]));
Q_ASSIGN U17288 ( .B(clk), .A(\g.we_clk [15486]));
Q_ASSIGN U17289 ( .B(clk), .A(\g.we_clk [15485]));
Q_ASSIGN U17290 ( .B(clk), .A(\g.we_clk [15484]));
Q_ASSIGN U17291 ( .B(clk), .A(\g.we_clk [15483]));
Q_ASSIGN U17292 ( .B(clk), .A(\g.we_clk [15482]));
Q_ASSIGN U17293 ( .B(clk), .A(\g.we_clk [15481]));
Q_ASSIGN U17294 ( .B(clk), .A(\g.we_clk [15480]));
Q_ASSIGN U17295 ( .B(clk), .A(\g.we_clk [15479]));
Q_ASSIGN U17296 ( .B(clk), .A(\g.we_clk [15478]));
Q_ASSIGN U17297 ( .B(clk), .A(\g.we_clk [15477]));
Q_ASSIGN U17298 ( .B(clk), .A(\g.we_clk [15476]));
Q_ASSIGN U17299 ( .B(clk), .A(\g.we_clk [15475]));
Q_ASSIGN U17300 ( .B(clk), .A(\g.we_clk [15474]));
Q_ASSIGN U17301 ( .B(clk), .A(\g.we_clk [15473]));
Q_ASSIGN U17302 ( .B(clk), .A(\g.we_clk [15472]));
Q_ASSIGN U17303 ( .B(clk), .A(\g.we_clk [15471]));
Q_ASSIGN U17304 ( .B(clk), .A(\g.we_clk [15470]));
Q_ASSIGN U17305 ( .B(clk), .A(\g.we_clk [15469]));
Q_ASSIGN U17306 ( .B(clk), .A(\g.we_clk [15468]));
Q_ASSIGN U17307 ( .B(clk), .A(\g.we_clk [15467]));
Q_ASSIGN U17308 ( .B(clk), .A(\g.we_clk [15466]));
Q_ASSIGN U17309 ( .B(clk), .A(\g.we_clk [15465]));
Q_ASSIGN U17310 ( .B(clk), .A(\g.we_clk [15464]));
Q_ASSIGN U17311 ( .B(clk), .A(\g.we_clk [15463]));
Q_ASSIGN U17312 ( .B(clk), .A(\g.we_clk [15462]));
Q_ASSIGN U17313 ( .B(clk), .A(\g.we_clk [15461]));
Q_ASSIGN U17314 ( .B(clk), .A(\g.we_clk [15460]));
Q_ASSIGN U17315 ( .B(clk), .A(\g.we_clk [15459]));
Q_ASSIGN U17316 ( .B(clk), .A(\g.we_clk [15458]));
Q_ASSIGN U17317 ( .B(clk), .A(\g.we_clk [15457]));
Q_ASSIGN U17318 ( .B(clk), .A(\g.we_clk [15456]));
Q_ASSIGN U17319 ( .B(clk), .A(\g.we_clk [15455]));
Q_ASSIGN U17320 ( .B(clk), .A(\g.we_clk [15454]));
Q_ASSIGN U17321 ( .B(clk), .A(\g.we_clk [15453]));
Q_ASSIGN U17322 ( .B(clk), .A(\g.we_clk [15452]));
Q_ASSIGN U17323 ( .B(clk), .A(\g.we_clk [15451]));
Q_ASSIGN U17324 ( .B(clk), .A(\g.we_clk [15450]));
Q_ASSIGN U17325 ( .B(clk), .A(\g.we_clk [15449]));
Q_ASSIGN U17326 ( .B(clk), .A(\g.we_clk [15448]));
Q_ASSIGN U17327 ( .B(clk), .A(\g.we_clk [15447]));
Q_ASSIGN U17328 ( .B(clk), .A(\g.we_clk [15446]));
Q_ASSIGN U17329 ( .B(clk), .A(\g.we_clk [15445]));
Q_ASSIGN U17330 ( .B(clk), .A(\g.we_clk [15444]));
Q_ASSIGN U17331 ( .B(clk), .A(\g.we_clk [15443]));
Q_ASSIGN U17332 ( .B(clk), .A(\g.we_clk [15442]));
Q_ASSIGN U17333 ( .B(clk), .A(\g.we_clk [15441]));
Q_ASSIGN U17334 ( .B(clk), .A(\g.we_clk [15440]));
Q_ASSIGN U17335 ( .B(clk), .A(\g.we_clk [15439]));
Q_ASSIGN U17336 ( .B(clk), .A(\g.we_clk [15438]));
Q_ASSIGN U17337 ( .B(clk), .A(\g.we_clk [15437]));
Q_ASSIGN U17338 ( .B(clk), .A(\g.we_clk [15436]));
Q_ASSIGN U17339 ( .B(clk), .A(\g.we_clk [15435]));
Q_ASSIGN U17340 ( .B(clk), .A(\g.we_clk [15434]));
Q_ASSIGN U17341 ( .B(clk), .A(\g.we_clk [15433]));
Q_ASSIGN U17342 ( .B(clk), .A(\g.we_clk [15432]));
Q_ASSIGN U17343 ( .B(clk), .A(\g.we_clk [15431]));
Q_ASSIGN U17344 ( .B(clk), .A(\g.we_clk [15430]));
Q_ASSIGN U17345 ( .B(clk), .A(\g.we_clk [15429]));
Q_ASSIGN U17346 ( .B(clk), .A(\g.we_clk [15428]));
Q_ASSIGN U17347 ( .B(clk), .A(\g.we_clk [15427]));
Q_ASSIGN U17348 ( .B(clk), .A(\g.we_clk [15426]));
Q_ASSIGN U17349 ( .B(clk), .A(\g.we_clk [15425]));
Q_ASSIGN U17350 ( .B(clk), .A(\g.we_clk [15424]));
Q_ASSIGN U17351 ( .B(clk), .A(\g.we_clk [15423]));
Q_ASSIGN U17352 ( .B(clk), .A(\g.we_clk [15422]));
Q_ASSIGN U17353 ( .B(clk), .A(\g.we_clk [15421]));
Q_ASSIGN U17354 ( .B(clk), .A(\g.we_clk [15420]));
Q_ASSIGN U17355 ( .B(clk), .A(\g.we_clk [15419]));
Q_ASSIGN U17356 ( .B(clk), .A(\g.we_clk [15418]));
Q_ASSIGN U17357 ( .B(clk), .A(\g.we_clk [15417]));
Q_ASSIGN U17358 ( .B(clk), .A(\g.we_clk [15416]));
Q_ASSIGN U17359 ( .B(clk), .A(\g.we_clk [15415]));
Q_ASSIGN U17360 ( .B(clk), .A(\g.we_clk [15414]));
Q_ASSIGN U17361 ( .B(clk), .A(\g.we_clk [15413]));
Q_ASSIGN U17362 ( .B(clk), .A(\g.we_clk [15412]));
Q_ASSIGN U17363 ( .B(clk), .A(\g.we_clk [15411]));
Q_ASSIGN U17364 ( .B(clk), .A(\g.we_clk [15410]));
Q_ASSIGN U17365 ( .B(clk), .A(\g.we_clk [15409]));
Q_ASSIGN U17366 ( .B(clk), .A(\g.we_clk [15408]));
Q_ASSIGN U17367 ( .B(clk), .A(\g.we_clk [15407]));
Q_ASSIGN U17368 ( .B(clk), .A(\g.we_clk [15406]));
Q_ASSIGN U17369 ( .B(clk), .A(\g.we_clk [15405]));
Q_ASSIGN U17370 ( .B(clk), .A(\g.we_clk [15404]));
Q_ASSIGN U17371 ( .B(clk), .A(\g.we_clk [15403]));
Q_ASSIGN U17372 ( .B(clk), .A(\g.we_clk [15402]));
Q_ASSIGN U17373 ( .B(clk), .A(\g.we_clk [15401]));
Q_ASSIGN U17374 ( .B(clk), .A(\g.we_clk [15400]));
Q_ASSIGN U17375 ( .B(clk), .A(\g.we_clk [15399]));
Q_ASSIGN U17376 ( .B(clk), .A(\g.we_clk [15398]));
Q_ASSIGN U17377 ( .B(clk), .A(\g.we_clk [15397]));
Q_ASSIGN U17378 ( .B(clk), .A(\g.we_clk [15396]));
Q_ASSIGN U17379 ( .B(clk), .A(\g.we_clk [15395]));
Q_ASSIGN U17380 ( .B(clk), .A(\g.we_clk [15394]));
Q_ASSIGN U17381 ( .B(clk), .A(\g.we_clk [15393]));
Q_ASSIGN U17382 ( .B(clk), .A(\g.we_clk [15392]));
Q_ASSIGN U17383 ( .B(clk), .A(\g.we_clk [15391]));
Q_ASSIGN U17384 ( .B(clk), .A(\g.we_clk [15390]));
Q_ASSIGN U17385 ( .B(clk), .A(\g.we_clk [15389]));
Q_ASSIGN U17386 ( .B(clk), .A(\g.we_clk [15388]));
Q_ASSIGN U17387 ( .B(clk), .A(\g.we_clk [15387]));
Q_ASSIGN U17388 ( .B(clk), .A(\g.we_clk [15386]));
Q_ASSIGN U17389 ( .B(clk), .A(\g.we_clk [15385]));
Q_ASSIGN U17390 ( .B(clk), .A(\g.we_clk [15384]));
Q_ASSIGN U17391 ( .B(clk), .A(\g.we_clk [15383]));
Q_ASSIGN U17392 ( .B(clk), .A(\g.we_clk [15382]));
Q_ASSIGN U17393 ( .B(clk), .A(\g.we_clk [15381]));
Q_ASSIGN U17394 ( .B(clk), .A(\g.we_clk [15380]));
Q_ASSIGN U17395 ( .B(clk), .A(\g.we_clk [15379]));
Q_ASSIGN U17396 ( .B(clk), .A(\g.we_clk [15378]));
Q_ASSIGN U17397 ( .B(clk), .A(\g.we_clk [15377]));
Q_ASSIGN U17398 ( .B(clk), .A(\g.we_clk [15376]));
Q_ASSIGN U17399 ( .B(clk), .A(\g.we_clk [15375]));
Q_ASSIGN U17400 ( .B(clk), .A(\g.we_clk [15374]));
Q_ASSIGN U17401 ( .B(clk), .A(\g.we_clk [15373]));
Q_ASSIGN U17402 ( .B(clk), .A(\g.we_clk [15372]));
Q_ASSIGN U17403 ( .B(clk), .A(\g.we_clk [15371]));
Q_ASSIGN U17404 ( .B(clk), .A(\g.we_clk [15370]));
Q_ASSIGN U17405 ( .B(clk), .A(\g.we_clk [15369]));
Q_ASSIGN U17406 ( .B(clk), .A(\g.we_clk [15368]));
Q_ASSIGN U17407 ( .B(clk), .A(\g.we_clk [15367]));
Q_ASSIGN U17408 ( .B(clk), .A(\g.we_clk [15366]));
Q_ASSIGN U17409 ( .B(clk), .A(\g.we_clk [15365]));
Q_ASSIGN U17410 ( .B(clk), .A(\g.we_clk [15364]));
Q_ASSIGN U17411 ( .B(clk), .A(\g.we_clk [15363]));
Q_ASSIGN U17412 ( .B(clk), .A(\g.we_clk [15362]));
Q_ASSIGN U17413 ( .B(clk), .A(\g.we_clk [15361]));
Q_ASSIGN U17414 ( .B(clk), .A(\g.we_clk [15360]));
Q_ASSIGN U17415 ( .B(clk), .A(\g.we_clk [15359]));
Q_ASSIGN U17416 ( .B(clk), .A(\g.we_clk [15358]));
Q_ASSIGN U17417 ( .B(clk), .A(\g.we_clk [15357]));
Q_ASSIGN U17418 ( .B(clk), .A(\g.we_clk [15356]));
Q_ASSIGN U17419 ( .B(clk), .A(\g.we_clk [15355]));
Q_ASSIGN U17420 ( .B(clk), .A(\g.we_clk [15354]));
Q_ASSIGN U17421 ( .B(clk), .A(\g.we_clk [15353]));
Q_ASSIGN U17422 ( .B(clk), .A(\g.we_clk [15352]));
Q_ASSIGN U17423 ( .B(clk), .A(\g.we_clk [15351]));
Q_ASSIGN U17424 ( .B(clk), .A(\g.we_clk [15350]));
Q_ASSIGN U17425 ( .B(clk), .A(\g.we_clk [15349]));
Q_ASSIGN U17426 ( .B(clk), .A(\g.we_clk [15348]));
Q_ASSIGN U17427 ( .B(clk), .A(\g.we_clk [15347]));
Q_ASSIGN U17428 ( .B(clk), .A(\g.we_clk [15346]));
Q_ASSIGN U17429 ( .B(clk), .A(\g.we_clk [15345]));
Q_ASSIGN U17430 ( .B(clk), .A(\g.we_clk [15344]));
Q_ASSIGN U17431 ( .B(clk), .A(\g.we_clk [15343]));
Q_ASSIGN U17432 ( .B(clk), .A(\g.we_clk [15342]));
Q_ASSIGN U17433 ( .B(clk), .A(\g.we_clk [15341]));
Q_ASSIGN U17434 ( .B(clk), .A(\g.we_clk [15340]));
Q_ASSIGN U17435 ( .B(clk), .A(\g.we_clk [15339]));
Q_ASSIGN U17436 ( .B(clk), .A(\g.we_clk [15338]));
Q_ASSIGN U17437 ( .B(clk), .A(\g.we_clk [15337]));
Q_ASSIGN U17438 ( .B(clk), .A(\g.we_clk [15336]));
Q_ASSIGN U17439 ( .B(clk), .A(\g.we_clk [15335]));
Q_ASSIGN U17440 ( .B(clk), .A(\g.we_clk [15334]));
Q_ASSIGN U17441 ( .B(clk), .A(\g.we_clk [15333]));
Q_ASSIGN U17442 ( .B(clk), .A(\g.we_clk [15332]));
Q_ASSIGN U17443 ( .B(clk), .A(\g.we_clk [15331]));
Q_ASSIGN U17444 ( .B(clk), .A(\g.we_clk [15330]));
Q_ASSIGN U17445 ( .B(clk), .A(\g.we_clk [15329]));
Q_ASSIGN U17446 ( .B(clk), .A(\g.we_clk [15328]));
Q_ASSIGN U17447 ( .B(clk), .A(\g.we_clk [15327]));
Q_ASSIGN U17448 ( .B(clk), .A(\g.we_clk [15326]));
Q_ASSIGN U17449 ( .B(clk), .A(\g.we_clk [15325]));
Q_ASSIGN U17450 ( .B(clk), .A(\g.we_clk [15324]));
Q_ASSIGN U17451 ( .B(clk), .A(\g.we_clk [15323]));
Q_ASSIGN U17452 ( .B(clk), .A(\g.we_clk [15322]));
Q_ASSIGN U17453 ( .B(clk), .A(\g.we_clk [15321]));
Q_ASSIGN U17454 ( .B(clk), .A(\g.we_clk [15320]));
Q_ASSIGN U17455 ( .B(clk), .A(\g.we_clk [15319]));
Q_ASSIGN U17456 ( .B(clk), .A(\g.we_clk [15318]));
Q_ASSIGN U17457 ( .B(clk), .A(\g.we_clk [15317]));
Q_ASSIGN U17458 ( .B(clk), .A(\g.we_clk [15316]));
Q_ASSIGN U17459 ( .B(clk), .A(\g.we_clk [15315]));
Q_ASSIGN U17460 ( .B(clk), .A(\g.we_clk [15314]));
Q_ASSIGN U17461 ( .B(clk), .A(\g.we_clk [15313]));
Q_ASSIGN U17462 ( .B(clk), .A(\g.we_clk [15312]));
Q_ASSIGN U17463 ( .B(clk), .A(\g.we_clk [15311]));
Q_ASSIGN U17464 ( .B(clk), .A(\g.we_clk [15310]));
Q_ASSIGN U17465 ( .B(clk), .A(\g.we_clk [15309]));
Q_ASSIGN U17466 ( .B(clk), .A(\g.we_clk [15308]));
Q_ASSIGN U17467 ( .B(clk), .A(\g.we_clk [15307]));
Q_ASSIGN U17468 ( .B(clk), .A(\g.we_clk [15306]));
Q_ASSIGN U17469 ( .B(clk), .A(\g.we_clk [15305]));
Q_ASSIGN U17470 ( .B(clk), .A(\g.we_clk [15304]));
Q_ASSIGN U17471 ( .B(clk), .A(\g.we_clk [15303]));
Q_ASSIGN U17472 ( .B(clk), .A(\g.we_clk [15302]));
Q_ASSIGN U17473 ( .B(clk), .A(\g.we_clk [15301]));
Q_ASSIGN U17474 ( .B(clk), .A(\g.we_clk [15300]));
Q_ASSIGN U17475 ( .B(clk), .A(\g.we_clk [15299]));
Q_ASSIGN U17476 ( .B(clk), .A(\g.we_clk [15298]));
Q_ASSIGN U17477 ( .B(clk), .A(\g.we_clk [15297]));
Q_ASSIGN U17478 ( .B(clk), .A(\g.we_clk [15296]));
Q_ASSIGN U17479 ( .B(clk), .A(\g.we_clk [15295]));
Q_ASSIGN U17480 ( .B(clk), .A(\g.we_clk [15294]));
Q_ASSIGN U17481 ( .B(clk), .A(\g.we_clk [15293]));
Q_ASSIGN U17482 ( .B(clk), .A(\g.we_clk [15292]));
Q_ASSIGN U17483 ( .B(clk), .A(\g.we_clk [15291]));
Q_ASSIGN U17484 ( .B(clk), .A(\g.we_clk [15290]));
Q_ASSIGN U17485 ( .B(clk), .A(\g.we_clk [15289]));
Q_ASSIGN U17486 ( .B(clk), .A(\g.we_clk [15288]));
Q_ASSIGN U17487 ( .B(clk), .A(\g.we_clk [15287]));
Q_ASSIGN U17488 ( .B(clk), .A(\g.we_clk [15286]));
Q_ASSIGN U17489 ( .B(clk), .A(\g.we_clk [15285]));
Q_ASSIGN U17490 ( .B(clk), .A(\g.we_clk [15284]));
Q_ASSIGN U17491 ( .B(clk), .A(\g.we_clk [15283]));
Q_ASSIGN U17492 ( .B(clk), .A(\g.we_clk [15282]));
Q_ASSIGN U17493 ( .B(clk), .A(\g.we_clk [15281]));
Q_ASSIGN U17494 ( .B(clk), .A(\g.we_clk [15280]));
Q_ASSIGN U17495 ( .B(clk), .A(\g.we_clk [15279]));
Q_ASSIGN U17496 ( .B(clk), .A(\g.we_clk [15278]));
Q_ASSIGN U17497 ( .B(clk), .A(\g.we_clk [15277]));
Q_ASSIGN U17498 ( .B(clk), .A(\g.we_clk [15276]));
Q_ASSIGN U17499 ( .B(clk), .A(\g.we_clk [15275]));
Q_ASSIGN U17500 ( .B(clk), .A(\g.we_clk [15274]));
Q_ASSIGN U17501 ( .B(clk), .A(\g.we_clk [15273]));
Q_ASSIGN U17502 ( .B(clk), .A(\g.we_clk [15272]));
Q_ASSIGN U17503 ( .B(clk), .A(\g.we_clk [15271]));
Q_ASSIGN U17504 ( .B(clk), .A(\g.we_clk [15270]));
Q_ASSIGN U17505 ( .B(clk), .A(\g.we_clk [15269]));
Q_ASSIGN U17506 ( .B(clk), .A(\g.we_clk [15268]));
Q_ASSIGN U17507 ( .B(clk), .A(\g.we_clk [15267]));
Q_ASSIGN U17508 ( .B(clk), .A(\g.we_clk [15266]));
Q_ASSIGN U17509 ( .B(clk), .A(\g.we_clk [15265]));
Q_ASSIGN U17510 ( .B(clk), .A(\g.we_clk [15264]));
Q_ASSIGN U17511 ( .B(clk), .A(\g.we_clk [15263]));
Q_ASSIGN U17512 ( .B(clk), .A(\g.we_clk [15262]));
Q_ASSIGN U17513 ( .B(clk), .A(\g.we_clk [15261]));
Q_ASSIGN U17514 ( .B(clk), .A(\g.we_clk [15260]));
Q_ASSIGN U17515 ( .B(clk), .A(\g.we_clk [15259]));
Q_ASSIGN U17516 ( .B(clk), .A(\g.we_clk [15258]));
Q_ASSIGN U17517 ( .B(clk), .A(\g.we_clk [15257]));
Q_ASSIGN U17518 ( .B(clk), .A(\g.we_clk [15256]));
Q_ASSIGN U17519 ( .B(clk), .A(\g.we_clk [15255]));
Q_ASSIGN U17520 ( .B(clk), .A(\g.we_clk [15254]));
Q_ASSIGN U17521 ( .B(clk), .A(\g.we_clk [15253]));
Q_ASSIGN U17522 ( .B(clk), .A(\g.we_clk [15252]));
Q_ASSIGN U17523 ( .B(clk), .A(\g.we_clk [15251]));
Q_ASSIGN U17524 ( .B(clk), .A(\g.we_clk [15250]));
Q_ASSIGN U17525 ( .B(clk), .A(\g.we_clk [15249]));
Q_ASSIGN U17526 ( .B(clk), .A(\g.we_clk [15248]));
Q_ASSIGN U17527 ( .B(clk), .A(\g.we_clk [15247]));
Q_ASSIGN U17528 ( .B(clk), .A(\g.we_clk [15246]));
Q_ASSIGN U17529 ( .B(clk), .A(\g.we_clk [15245]));
Q_ASSIGN U17530 ( .B(clk), .A(\g.we_clk [15244]));
Q_ASSIGN U17531 ( .B(clk), .A(\g.we_clk [15243]));
Q_ASSIGN U17532 ( .B(clk), .A(\g.we_clk [15242]));
Q_ASSIGN U17533 ( .B(clk), .A(\g.we_clk [15241]));
Q_ASSIGN U17534 ( .B(clk), .A(\g.we_clk [15240]));
Q_ASSIGN U17535 ( .B(clk), .A(\g.we_clk [15239]));
Q_ASSIGN U17536 ( .B(clk), .A(\g.we_clk [15238]));
Q_ASSIGN U17537 ( .B(clk), .A(\g.we_clk [15237]));
Q_ASSIGN U17538 ( .B(clk), .A(\g.we_clk [15236]));
Q_ASSIGN U17539 ( .B(clk), .A(\g.we_clk [15235]));
Q_ASSIGN U17540 ( .B(clk), .A(\g.we_clk [15234]));
Q_ASSIGN U17541 ( .B(clk), .A(\g.we_clk [15233]));
Q_ASSIGN U17542 ( .B(clk), .A(\g.we_clk [15232]));
Q_ASSIGN U17543 ( .B(clk), .A(\g.we_clk [15231]));
Q_ASSIGN U17544 ( .B(clk), .A(\g.we_clk [15230]));
Q_ASSIGN U17545 ( .B(clk), .A(\g.we_clk [15229]));
Q_ASSIGN U17546 ( .B(clk), .A(\g.we_clk [15228]));
Q_ASSIGN U17547 ( .B(clk), .A(\g.we_clk [15227]));
Q_ASSIGN U17548 ( .B(clk), .A(\g.we_clk [15226]));
Q_ASSIGN U17549 ( .B(clk), .A(\g.we_clk [15225]));
Q_ASSIGN U17550 ( .B(clk), .A(\g.we_clk [15224]));
Q_ASSIGN U17551 ( .B(clk), .A(\g.we_clk [15223]));
Q_ASSIGN U17552 ( .B(clk), .A(\g.we_clk [15222]));
Q_ASSIGN U17553 ( .B(clk), .A(\g.we_clk [15221]));
Q_ASSIGN U17554 ( .B(clk), .A(\g.we_clk [15220]));
Q_ASSIGN U17555 ( .B(clk), .A(\g.we_clk [15219]));
Q_ASSIGN U17556 ( .B(clk), .A(\g.we_clk [15218]));
Q_ASSIGN U17557 ( .B(clk), .A(\g.we_clk [15217]));
Q_ASSIGN U17558 ( .B(clk), .A(\g.we_clk [15216]));
Q_ASSIGN U17559 ( .B(clk), .A(\g.we_clk [15215]));
Q_ASSIGN U17560 ( .B(clk), .A(\g.we_clk [15214]));
Q_ASSIGN U17561 ( .B(clk), .A(\g.we_clk [15213]));
Q_ASSIGN U17562 ( .B(clk), .A(\g.we_clk [15212]));
Q_ASSIGN U17563 ( .B(clk), .A(\g.we_clk [15211]));
Q_ASSIGN U17564 ( .B(clk), .A(\g.we_clk [15210]));
Q_ASSIGN U17565 ( .B(clk), .A(\g.we_clk [15209]));
Q_ASSIGN U17566 ( .B(clk), .A(\g.we_clk [15208]));
Q_ASSIGN U17567 ( .B(clk), .A(\g.we_clk [15207]));
Q_ASSIGN U17568 ( .B(clk), .A(\g.we_clk [15206]));
Q_ASSIGN U17569 ( .B(clk), .A(\g.we_clk [15205]));
Q_ASSIGN U17570 ( .B(clk), .A(\g.we_clk [15204]));
Q_ASSIGN U17571 ( .B(clk), .A(\g.we_clk [15203]));
Q_ASSIGN U17572 ( .B(clk), .A(\g.we_clk [15202]));
Q_ASSIGN U17573 ( .B(clk), .A(\g.we_clk [15201]));
Q_ASSIGN U17574 ( .B(clk), .A(\g.we_clk [15200]));
Q_ASSIGN U17575 ( .B(clk), .A(\g.we_clk [15199]));
Q_ASSIGN U17576 ( .B(clk), .A(\g.we_clk [15198]));
Q_ASSIGN U17577 ( .B(clk), .A(\g.we_clk [15197]));
Q_ASSIGN U17578 ( .B(clk), .A(\g.we_clk [15196]));
Q_ASSIGN U17579 ( .B(clk), .A(\g.we_clk [15195]));
Q_ASSIGN U17580 ( .B(clk), .A(\g.we_clk [15194]));
Q_ASSIGN U17581 ( .B(clk), .A(\g.we_clk [15193]));
Q_ASSIGN U17582 ( .B(clk), .A(\g.we_clk [15192]));
Q_ASSIGN U17583 ( .B(clk), .A(\g.we_clk [15191]));
Q_ASSIGN U17584 ( .B(clk), .A(\g.we_clk [15190]));
Q_ASSIGN U17585 ( .B(clk), .A(\g.we_clk [15189]));
Q_ASSIGN U17586 ( .B(clk), .A(\g.we_clk [15188]));
Q_ASSIGN U17587 ( .B(clk), .A(\g.we_clk [15187]));
Q_ASSIGN U17588 ( .B(clk), .A(\g.we_clk [15186]));
Q_ASSIGN U17589 ( .B(clk), .A(\g.we_clk [15185]));
Q_ASSIGN U17590 ( .B(clk), .A(\g.we_clk [15184]));
Q_ASSIGN U17591 ( .B(clk), .A(\g.we_clk [15183]));
Q_ASSIGN U17592 ( .B(clk), .A(\g.we_clk [15182]));
Q_ASSIGN U17593 ( .B(clk), .A(\g.we_clk [15181]));
Q_ASSIGN U17594 ( .B(clk), .A(\g.we_clk [15180]));
Q_ASSIGN U17595 ( .B(clk), .A(\g.we_clk [15179]));
Q_ASSIGN U17596 ( .B(clk), .A(\g.we_clk [15178]));
Q_ASSIGN U17597 ( .B(clk), .A(\g.we_clk [15177]));
Q_ASSIGN U17598 ( .B(clk), .A(\g.we_clk [15176]));
Q_ASSIGN U17599 ( .B(clk), .A(\g.we_clk [15175]));
Q_ASSIGN U17600 ( .B(clk), .A(\g.we_clk [15174]));
Q_ASSIGN U17601 ( .B(clk), .A(\g.we_clk [15173]));
Q_ASSIGN U17602 ( .B(clk), .A(\g.we_clk [15172]));
Q_ASSIGN U17603 ( .B(clk), .A(\g.we_clk [15171]));
Q_ASSIGN U17604 ( .B(clk), .A(\g.we_clk [15170]));
Q_ASSIGN U17605 ( .B(clk), .A(\g.we_clk [15169]));
Q_ASSIGN U17606 ( .B(clk), .A(\g.we_clk [15168]));
Q_ASSIGN U17607 ( .B(clk), .A(\g.we_clk [15167]));
Q_ASSIGN U17608 ( .B(clk), .A(\g.we_clk [15166]));
Q_ASSIGN U17609 ( .B(clk), .A(\g.we_clk [15165]));
Q_ASSIGN U17610 ( .B(clk), .A(\g.we_clk [15164]));
Q_ASSIGN U17611 ( .B(clk), .A(\g.we_clk [15163]));
Q_ASSIGN U17612 ( .B(clk), .A(\g.we_clk [15162]));
Q_ASSIGN U17613 ( .B(clk), .A(\g.we_clk [15161]));
Q_ASSIGN U17614 ( .B(clk), .A(\g.we_clk [15160]));
Q_ASSIGN U17615 ( .B(clk), .A(\g.we_clk [15159]));
Q_ASSIGN U17616 ( .B(clk), .A(\g.we_clk [15158]));
Q_ASSIGN U17617 ( .B(clk), .A(\g.we_clk [15157]));
Q_ASSIGN U17618 ( .B(clk), .A(\g.we_clk [15156]));
Q_ASSIGN U17619 ( .B(clk), .A(\g.we_clk [15155]));
Q_ASSIGN U17620 ( .B(clk), .A(\g.we_clk [15154]));
Q_ASSIGN U17621 ( .B(clk), .A(\g.we_clk [15153]));
Q_ASSIGN U17622 ( .B(clk), .A(\g.we_clk [15152]));
Q_ASSIGN U17623 ( .B(clk), .A(\g.we_clk [15151]));
Q_ASSIGN U17624 ( .B(clk), .A(\g.we_clk [15150]));
Q_ASSIGN U17625 ( .B(clk), .A(\g.we_clk [15149]));
Q_ASSIGN U17626 ( .B(clk), .A(\g.we_clk [15148]));
Q_ASSIGN U17627 ( .B(clk), .A(\g.we_clk [15147]));
Q_ASSIGN U17628 ( .B(clk), .A(\g.we_clk [15146]));
Q_ASSIGN U17629 ( .B(clk), .A(\g.we_clk [15145]));
Q_ASSIGN U17630 ( .B(clk), .A(\g.we_clk [15144]));
Q_ASSIGN U17631 ( .B(clk), .A(\g.we_clk [15143]));
Q_ASSIGN U17632 ( .B(clk), .A(\g.we_clk [15142]));
Q_ASSIGN U17633 ( .B(clk), .A(\g.we_clk [15141]));
Q_ASSIGN U17634 ( .B(clk), .A(\g.we_clk [15140]));
Q_ASSIGN U17635 ( .B(clk), .A(\g.we_clk [15139]));
Q_ASSIGN U17636 ( .B(clk), .A(\g.we_clk [15138]));
Q_ASSIGN U17637 ( .B(clk), .A(\g.we_clk [15137]));
Q_ASSIGN U17638 ( .B(clk), .A(\g.we_clk [15136]));
Q_ASSIGN U17639 ( .B(clk), .A(\g.we_clk [15135]));
Q_ASSIGN U17640 ( .B(clk), .A(\g.we_clk [15134]));
Q_ASSIGN U17641 ( .B(clk), .A(\g.we_clk [15133]));
Q_ASSIGN U17642 ( .B(clk), .A(\g.we_clk [15132]));
Q_ASSIGN U17643 ( .B(clk), .A(\g.we_clk [15131]));
Q_ASSIGN U17644 ( .B(clk), .A(\g.we_clk [15130]));
Q_ASSIGN U17645 ( .B(clk), .A(\g.we_clk [15129]));
Q_ASSIGN U17646 ( .B(clk), .A(\g.we_clk [15128]));
Q_ASSIGN U17647 ( .B(clk), .A(\g.we_clk [15127]));
Q_ASSIGN U17648 ( .B(clk), .A(\g.we_clk [15126]));
Q_ASSIGN U17649 ( .B(clk), .A(\g.we_clk [15125]));
Q_ASSIGN U17650 ( .B(clk), .A(\g.we_clk [15124]));
Q_ASSIGN U17651 ( .B(clk), .A(\g.we_clk [15123]));
Q_ASSIGN U17652 ( .B(clk), .A(\g.we_clk [15122]));
Q_ASSIGN U17653 ( .B(clk), .A(\g.we_clk [15121]));
Q_ASSIGN U17654 ( .B(clk), .A(\g.we_clk [15120]));
Q_ASSIGN U17655 ( .B(clk), .A(\g.we_clk [15119]));
Q_ASSIGN U17656 ( .B(clk), .A(\g.we_clk [15118]));
Q_ASSIGN U17657 ( .B(clk), .A(\g.we_clk [15117]));
Q_ASSIGN U17658 ( .B(clk), .A(\g.we_clk [15116]));
Q_ASSIGN U17659 ( .B(clk), .A(\g.we_clk [15115]));
Q_ASSIGN U17660 ( .B(clk), .A(\g.we_clk [15114]));
Q_ASSIGN U17661 ( .B(clk), .A(\g.we_clk [15113]));
Q_ASSIGN U17662 ( .B(clk), .A(\g.we_clk [15112]));
Q_ASSIGN U17663 ( .B(clk), .A(\g.we_clk [15111]));
Q_ASSIGN U17664 ( .B(clk), .A(\g.we_clk [15110]));
Q_ASSIGN U17665 ( .B(clk), .A(\g.we_clk [15109]));
Q_ASSIGN U17666 ( .B(clk), .A(\g.we_clk [15108]));
Q_ASSIGN U17667 ( .B(clk), .A(\g.we_clk [15107]));
Q_ASSIGN U17668 ( .B(clk), .A(\g.we_clk [15106]));
Q_ASSIGN U17669 ( .B(clk), .A(\g.we_clk [15105]));
Q_ASSIGN U17670 ( .B(clk), .A(\g.we_clk [15104]));
Q_ASSIGN U17671 ( .B(clk), .A(\g.we_clk [15103]));
Q_ASSIGN U17672 ( .B(clk), .A(\g.we_clk [15102]));
Q_ASSIGN U17673 ( .B(clk), .A(\g.we_clk [15101]));
Q_ASSIGN U17674 ( .B(clk), .A(\g.we_clk [15100]));
Q_ASSIGN U17675 ( .B(clk), .A(\g.we_clk [15099]));
Q_ASSIGN U17676 ( .B(clk), .A(\g.we_clk [15098]));
Q_ASSIGN U17677 ( .B(clk), .A(\g.we_clk [15097]));
Q_ASSIGN U17678 ( .B(clk), .A(\g.we_clk [15096]));
Q_ASSIGN U17679 ( .B(clk), .A(\g.we_clk [15095]));
Q_ASSIGN U17680 ( .B(clk), .A(\g.we_clk [15094]));
Q_ASSIGN U17681 ( .B(clk), .A(\g.we_clk [15093]));
Q_ASSIGN U17682 ( .B(clk), .A(\g.we_clk [15092]));
Q_ASSIGN U17683 ( .B(clk), .A(\g.we_clk [15091]));
Q_ASSIGN U17684 ( .B(clk), .A(\g.we_clk [15090]));
Q_ASSIGN U17685 ( .B(clk), .A(\g.we_clk [15089]));
Q_ASSIGN U17686 ( .B(clk), .A(\g.we_clk [15088]));
Q_ASSIGN U17687 ( .B(clk), .A(\g.we_clk [15087]));
Q_ASSIGN U17688 ( .B(clk), .A(\g.we_clk [15086]));
Q_ASSIGN U17689 ( .B(clk), .A(\g.we_clk [15085]));
Q_ASSIGN U17690 ( .B(clk), .A(\g.we_clk [15084]));
Q_ASSIGN U17691 ( .B(clk), .A(\g.we_clk [15083]));
Q_ASSIGN U17692 ( .B(clk), .A(\g.we_clk [15082]));
Q_ASSIGN U17693 ( .B(clk), .A(\g.we_clk [15081]));
Q_ASSIGN U17694 ( .B(clk), .A(\g.we_clk [15080]));
Q_ASSIGN U17695 ( .B(clk), .A(\g.we_clk [15079]));
Q_ASSIGN U17696 ( .B(clk), .A(\g.we_clk [15078]));
Q_ASSIGN U17697 ( .B(clk), .A(\g.we_clk [15077]));
Q_ASSIGN U17698 ( .B(clk), .A(\g.we_clk [15076]));
Q_ASSIGN U17699 ( .B(clk), .A(\g.we_clk [15075]));
Q_ASSIGN U17700 ( .B(clk), .A(\g.we_clk [15074]));
Q_ASSIGN U17701 ( .B(clk), .A(\g.we_clk [15073]));
Q_ASSIGN U17702 ( .B(clk), .A(\g.we_clk [15072]));
Q_ASSIGN U17703 ( .B(clk), .A(\g.we_clk [15071]));
Q_ASSIGN U17704 ( .B(clk), .A(\g.we_clk [15070]));
Q_ASSIGN U17705 ( .B(clk), .A(\g.we_clk [15069]));
Q_ASSIGN U17706 ( .B(clk), .A(\g.we_clk [15068]));
Q_ASSIGN U17707 ( .B(clk), .A(\g.we_clk [15067]));
Q_ASSIGN U17708 ( .B(clk), .A(\g.we_clk [15066]));
Q_ASSIGN U17709 ( .B(clk), .A(\g.we_clk [15065]));
Q_ASSIGN U17710 ( .B(clk), .A(\g.we_clk [15064]));
Q_ASSIGN U17711 ( .B(clk), .A(\g.we_clk [15063]));
Q_ASSIGN U17712 ( .B(clk), .A(\g.we_clk [15062]));
Q_ASSIGN U17713 ( .B(clk), .A(\g.we_clk [15061]));
Q_ASSIGN U17714 ( .B(clk), .A(\g.we_clk [15060]));
Q_ASSIGN U17715 ( .B(clk), .A(\g.we_clk [15059]));
Q_ASSIGN U17716 ( .B(clk), .A(\g.we_clk [15058]));
Q_ASSIGN U17717 ( .B(clk), .A(\g.we_clk [15057]));
Q_ASSIGN U17718 ( .B(clk), .A(\g.we_clk [15056]));
Q_ASSIGN U17719 ( .B(clk), .A(\g.we_clk [15055]));
Q_ASSIGN U17720 ( .B(clk), .A(\g.we_clk [15054]));
Q_ASSIGN U17721 ( .B(clk), .A(\g.we_clk [15053]));
Q_ASSIGN U17722 ( .B(clk), .A(\g.we_clk [15052]));
Q_ASSIGN U17723 ( .B(clk), .A(\g.we_clk [15051]));
Q_ASSIGN U17724 ( .B(clk), .A(\g.we_clk [15050]));
Q_ASSIGN U17725 ( .B(clk), .A(\g.we_clk [15049]));
Q_ASSIGN U17726 ( .B(clk), .A(\g.we_clk [15048]));
Q_ASSIGN U17727 ( .B(clk), .A(\g.we_clk [15047]));
Q_ASSIGN U17728 ( .B(clk), .A(\g.we_clk [15046]));
Q_ASSIGN U17729 ( .B(clk), .A(\g.we_clk [15045]));
Q_ASSIGN U17730 ( .B(clk), .A(\g.we_clk [15044]));
Q_ASSIGN U17731 ( .B(clk), .A(\g.we_clk [15043]));
Q_ASSIGN U17732 ( .B(clk), .A(\g.we_clk [15042]));
Q_ASSIGN U17733 ( .B(clk), .A(\g.we_clk [15041]));
Q_ASSIGN U17734 ( .B(clk), .A(\g.we_clk [15040]));
Q_ASSIGN U17735 ( .B(clk), .A(\g.we_clk [15039]));
Q_ASSIGN U17736 ( .B(clk), .A(\g.we_clk [15038]));
Q_ASSIGN U17737 ( .B(clk), .A(\g.we_clk [15037]));
Q_ASSIGN U17738 ( .B(clk), .A(\g.we_clk [15036]));
Q_ASSIGN U17739 ( .B(clk), .A(\g.we_clk [15035]));
Q_ASSIGN U17740 ( .B(clk), .A(\g.we_clk [15034]));
Q_ASSIGN U17741 ( .B(clk), .A(\g.we_clk [15033]));
Q_ASSIGN U17742 ( .B(clk), .A(\g.we_clk [15032]));
Q_ASSIGN U17743 ( .B(clk), .A(\g.we_clk [15031]));
Q_ASSIGN U17744 ( .B(clk), .A(\g.we_clk [15030]));
Q_ASSIGN U17745 ( .B(clk), .A(\g.we_clk [15029]));
Q_ASSIGN U17746 ( .B(clk), .A(\g.we_clk [15028]));
Q_ASSIGN U17747 ( .B(clk), .A(\g.we_clk [15027]));
Q_ASSIGN U17748 ( .B(clk), .A(\g.we_clk [15026]));
Q_ASSIGN U17749 ( .B(clk), .A(\g.we_clk [15025]));
Q_ASSIGN U17750 ( .B(clk), .A(\g.we_clk [15024]));
Q_ASSIGN U17751 ( .B(clk), .A(\g.we_clk [15023]));
Q_ASSIGN U17752 ( .B(clk), .A(\g.we_clk [15022]));
Q_ASSIGN U17753 ( .B(clk), .A(\g.we_clk [15021]));
Q_ASSIGN U17754 ( .B(clk), .A(\g.we_clk [15020]));
Q_ASSIGN U17755 ( .B(clk), .A(\g.we_clk [15019]));
Q_ASSIGN U17756 ( .B(clk), .A(\g.we_clk [15018]));
Q_ASSIGN U17757 ( .B(clk), .A(\g.we_clk [15017]));
Q_ASSIGN U17758 ( .B(clk), .A(\g.we_clk [15016]));
Q_ASSIGN U17759 ( .B(clk), .A(\g.we_clk [15015]));
Q_ASSIGN U17760 ( .B(clk), .A(\g.we_clk [15014]));
Q_ASSIGN U17761 ( .B(clk), .A(\g.we_clk [15013]));
Q_ASSIGN U17762 ( .B(clk), .A(\g.we_clk [15012]));
Q_ASSIGN U17763 ( .B(clk), .A(\g.we_clk [15011]));
Q_ASSIGN U17764 ( .B(clk), .A(\g.we_clk [15010]));
Q_ASSIGN U17765 ( .B(clk), .A(\g.we_clk [15009]));
Q_ASSIGN U17766 ( .B(clk), .A(\g.we_clk [15008]));
Q_ASSIGN U17767 ( .B(clk), .A(\g.we_clk [15007]));
Q_ASSIGN U17768 ( .B(clk), .A(\g.we_clk [15006]));
Q_ASSIGN U17769 ( .B(clk), .A(\g.we_clk [15005]));
Q_ASSIGN U17770 ( .B(clk), .A(\g.we_clk [15004]));
Q_ASSIGN U17771 ( .B(clk), .A(\g.we_clk [15003]));
Q_ASSIGN U17772 ( .B(clk), .A(\g.we_clk [15002]));
Q_ASSIGN U17773 ( .B(clk), .A(\g.we_clk [15001]));
Q_ASSIGN U17774 ( .B(clk), .A(\g.we_clk [15000]));
Q_ASSIGN U17775 ( .B(clk), .A(\g.we_clk [14999]));
Q_ASSIGN U17776 ( .B(clk), .A(\g.we_clk [14998]));
Q_ASSIGN U17777 ( .B(clk), .A(\g.we_clk [14997]));
Q_ASSIGN U17778 ( .B(clk), .A(\g.we_clk [14996]));
Q_ASSIGN U17779 ( .B(clk), .A(\g.we_clk [14995]));
Q_ASSIGN U17780 ( .B(clk), .A(\g.we_clk [14994]));
Q_ASSIGN U17781 ( .B(clk), .A(\g.we_clk [14993]));
Q_ASSIGN U17782 ( .B(clk), .A(\g.we_clk [14992]));
Q_ASSIGN U17783 ( .B(clk), .A(\g.we_clk [14991]));
Q_ASSIGN U17784 ( .B(clk), .A(\g.we_clk [14990]));
Q_ASSIGN U17785 ( .B(clk), .A(\g.we_clk [14989]));
Q_ASSIGN U17786 ( .B(clk), .A(\g.we_clk [14988]));
Q_ASSIGN U17787 ( .B(clk), .A(\g.we_clk [14987]));
Q_ASSIGN U17788 ( .B(clk), .A(\g.we_clk [14986]));
Q_ASSIGN U17789 ( .B(clk), .A(\g.we_clk [14985]));
Q_ASSIGN U17790 ( .B(clk), .A(\g.we_clk [14984]));
Q_ASSIGN U17791 ( .B(clk), .A(\g.we_clk [14983]));
Q_ASSIGN U17792 ( .B(clk), .A(\g.we_clk [14982]));
Q_ASSIGN U17793 ( .B(clk), .A(\g.we_clk [14981]));
Q_ASSIGN U17794 ( .B(clk), .A(\g.we_clk [14980]));
Q_ASSIGN U17795 ( .B(clk), .A(\g.we_clk [14979]));
Q_ASSIGN U17796 ( .B(clk), .A(\g.we_clk [14978]));
Q_ASSIGN U17797 ( .B(clk), .A(\g.we_clk [14977]));
Q_ASSIGN U17798 ( .B(clk), .A(\g.we_clk [14976]));
Q_ASSIGN U17799 ( .B(clk), .A(\g.we_clk [14975]));
Q_ASSIGN U17800 ( .B(clk), .A(\g.we_clk [14974]));
Q_ASSIGN U17801 ( .B(clk), .A(\g.we_clk [14973]));
Q_ASSIGN U17802 ( .B(clk), .A(\g.we_clk [14972]));
Q_ASSIGN U17803 ( .B(clk), .A(\g.we_clk [14971]));
Q_ASSIGN U17804 ( .B(clk), .A(\g.we_clk [14970]));
Q_ASSIGN U17805 ( .B(clk), .A(\g.we_clk [14969]));
Q_ASSIGN U17806 ( .B(clk), .A(\g.we_clk [14968]));
Q_ASSIGN U17807 ( .B(clk), .A(\g.we_clk [14967]));
Q_ASSIGN U17808 ( .B(clk), .A(\g.we_clk [14966]));
Q_ASSIGN U17809 ( .B(clk), .A(\g.we_clk [14965]));
Q_ASSIGN U17810 ( .B(clk), .A(\g.we_clk [14964]));
Q_ASSIGN U17811 ( .B(clk), .A(\g.we_clk [14963]));
Q_ASSIGN U17812 ( .B(clk), .A(\g.we_clk [14962]));
Q_ASSIGN U17813 ( .B(clk), .A(\g.we_clk [14961]));
Q_ASSIGN U17814 ( .B(clk), .A(\g.we_clk [14960]));
Q_ASSIGN U17815 ( .B(clk), .A(\g.we_clk [14959]));
Q_ASSIGN U17816 ( .B(clk), .A(\g.we_clk [14958]));
Q_ASSIGN U17817 ( .B(clk), .A(\g.we_clk [14957]));
Q_ASSIGN U17818 ( .B(clk), .A(\g.we_clk [14956]));
Q_ASSIGN U17819 ( .B(clk), .A(\g.we_clk [14955]));
Q_ASSIGN U17820 ( .B(clk), .A(\g.we_clk [14954]));
Q_ASSIGN U17821 ( .B(clk), .A(\g.we_clk [14953]));
Q_ASSIGN U17822 ( .B(clk), .A(\g.we_clk [14952]));
Q_ASSIGN U17823 ( .B(clk), .A(\g.we_clk [14951]));
Q_ASSIGN U17824 ( .B(clk), .A(\g.we_clk [14950]));
Q_ASSIGN U17825 ( .B(clk), .A(\g.we_clk [14949]));
Q_ASSIGN U17826 ( .B(clk), .A(\g.we_clk [14948]));
Q_ASSIGN U17827 ( .B(clk), .A(\g.we_clk [14947]));
Q_ASSIGN U17828 ( .B(clk), .A(\g.we_clk [14946]));
Q_ASSIGN U17829 ( .B(clk), .A(\g.we_clk [14945]));
Q_ASSIGN U17830 ( .B(clk), .A(\g.we_clk [14944]));
Q_ASSIGN U17831 ( .B(clk), .A(\g.we_clk [14943]));
Q_ASSIGN U17832 ( .B(clk), .A(\g.we_clk [14942]));
Q_ASSIGN U17833 ( .B(clk), .A(\g.we_clk [14941]));
Q_ASSIGN U17834 ( .B(clk), .A(\g.we_clk [14940]));
Q_ASSIGN U17835 ( .B(clk), .A(\g.we_clk [14939]));
Q_ASSIGN U17836 ( .B(clk), .A(\g.we_clk [14938]));
Q_ASSIGN U17837 ( .B(clk), .A(\g.we_clk [14937]));
Q_ASSIGN U17838 ( .B(clk), .A(\g.we_clk [14936]));
Q_ASSIGN U17839 ( .B(clk), .A(\g.we_clk [14935]));
Q_ASSIGN U17840 ( .B(clk), .A(\g.we_clk [14934]));
Q_ASSIGN U17841 ( .B(clk), .A(\g.we_clk [14933]));
Q_ASSIGN U17842 ( .B(clk), .A(\g.we_clk [14932]));
Q_ASSIGN U17843 ( .B(clk), .A(\g.we_clk [14931]));
Q_ASSIGN U17844 ( .B(clk), .A(\g.we_clk [14930]));
Q_ASSIGN U17845 ( .B(clk), .A(\g.we_clk [14929]));
Q_ASSIGN U17846 ( .B(clk), .A(\g.we_clk [14928]));
Q_ASSIGN U17847 ( .B(clk), .A(\g.we_clk [14927]));
Q_ASSIGN U17848 ( .B(clk), .A(\g.we_clk [14926]));
Q_ASSIGN U17849 ( .B(clk), .A(\g.we_clk [14925]));
Q_ASSIGN U17850 ( .B(clk), .A(\g.we_clk [14924]));
Q_ASSIGN U17851 ( .B(clk), .A(\g.we_clk [14923]));
Q_ASSIGN U17852 ( .B(clk), .A(\g.we_clk [14922]));
Q_ASSIGN U17853 ( .B(clk), .A(\g.we_clk [14921]));
Q_ASSIGN U17854 ( .B(clk), .A(\g.we_clk [14920]));
Q_ASSIGN U17855 ( .B(clk), .A(\g.we_clk [14919]));
Q_ASSIGN U17856 ( .B(clk), .A(\g.we_clk [14918]));
Q_ASSIGN U17857 ( .B(clk), .A(\g.we_clk [14917]));
Q_ASSIGN U17858 ( .B(clk), .A(\g.we_clk [14916]));
Q_ASSIGN U17859 ( .B(clk), .A(\g.we_clk [14915]));
Q_ASSIGN U17860 ( .B(clk), .A(\g.we_clk [14914]));
Q_ASSIGN U17861 ( .B(clk), .A(\g.we_clk [14913]));
Q_ASSIGN U17862 ( .B(clk), .A(\g.we_clk [14912]));
Q_ASSIGN U17863 ( .B(clk), .A(\g.we_clk [14911]));
Q_ASSIGN U17864 ( .B(clk), .A(\g.we_clk [14910]));
Q_ASSIGN U17865 ( .B(clk), .A(\g.we_clk [14909]));
Q_ASSIGN U17866 ( .B(clk), .A(\g.we_clk [14908]));
Q_ASSIGN U17867 ( .B(clk), .A(\g.we_clk [14907]));
Q_ASSIGN U17868 ( .B(clk), .A(\g.we_clk [14906]));
Q_ASSIGN U17869 ( .B(clk), .A(\g.we_clk [14905]));
Q_ASSIGN U17870 ( .B(clk), .A(\g.we_clk [14904]));
Q_ASSIGN U17871 ( .B(clk), .A(\g.we_clk [14903]));
Q_ASSIGN U17872 ( .B(clk), .A(\g.we_clk [14902]));
Q_ASSIGN U17873 ( .B(clk), .A(\g.we_clk [14901]));
Q_ASSIGN U17874 ( .B(clk), .A(\g.we_clk [14900]));
Q_ASSIGN U17875 ( .B(clk), .A(\g.we_clk [14899]));
Q_ASSIGN U17876 ( .B(clk), .A(\g.we_clk [14898]));
Q_ASSIGN U17877 ( .B(clk), .A(\g.we_clk [14897]));
Q_ASSIGN U17878 ( .B(clk), .A(\g.we_clk [14896]));
Q_ASSIGN U17879 ( .B(clk), .A(\g.we_clk [14895]));
Q_ASSIGN U17880 ( .B(clk), .A(\g.we_clk [14894]));
Q_ASSIGN U17881 ( .B(clk), .A(\g.we_clk [14893]));
Q_ASSIGN U17882 ( .B(clk), .A(\g.we_clk [14892]));
Q_ASSIGN U17883 ( .B(clk), .A(\g.we_clk [14891]));
Q_ASSIGN U17884 ( .B(clk), .A(\g.we_clk [14890]));
Q_ASSIGN U17885 ( .B(clk), .A(\g.we_clk [14889]));
Q_ASSIGN U17886 ( .B(clk), .A(\g.we_clk [14888]));
Q_ASSIGN U17887 ( .B(clk), .A(\g.we_clk [14887]));
Q_ASSIGN U17888 ( .B(clk), .A(\g.we_clk [14886]));
Q_ASSIGN U17889 ( .B(clk), .A(\g.we_clk [14885]));
Q_ASSIGN U17890 ( .B(clk), .A(\g.we_clk [14884]));
Q_ASSIGN U17891 ( .B(clk), .A(\g.we_clk [14883]));
Q_ASSIGN U17892 ( .B(clk), .A(\g.we_clk [14882]));
Q_ASSIGN U17893 ( .B(clk), .A(\g.we_clk [14881]));
Q_ASSIGN U17894 ( .B(clk), .A(\g.we_clk [14880]));
Q_ASSIGN U17895 ( .B(clk), .A(\g.we_clk [14879]));
Q_ASSIGN U17896 ( .B(clk), .A(\g.we_clk [14878]));
Q_ASSIGN U17897 ( .B(clk), .A(\g.we_clk [14877]));
Q_ASSIGN U17898 ( .B(clk), .A(\g.we_clk [14876]));
Q_ASSIGN U17899 ( .B(clk), .A(\g.we_clk [14875]));
Q_ASSIGN U17900 ( .B(clk), .A(\g.we_clk [14874]));
Q_ASSIGN U17901 ( .B(clk), .A(\g.we_clk [14873]));
Q_ASSIGN U17902 ( .B(clk), .A(\g.we_clk [14872]));
Q_ASSIGN U17903 ( .B(clk), .A(\g.we_clk [14871]));
Q_ASSIGN U17904 ( .B(clk), .A(\g.we_clk [14870]));
Q_ASSIGN U17905 ( .B(clk), .A(\g.we_clk [14869]));
Q_ASSIGN U17906 ( .B(clk), .A(\g.we_clk [14868]));
Q_ASSIGN U17907 ( .B(clk), .A(\g.we_clk [14867]));
Q_ASSIGN U17908 ( .B(clk), .A(\g.we_clk [14866]));
Q_ASSIGN U17909 ( .B(clk), .A(\g.we_clk [14865]));
Q_ASSIGN U17910 ( .B(clk), .A(\g.we_clk [14864]));
Q_ASSIGN U17911 ( .B(clk), .A(\g.we_clk [14863]));
Q_ASSIGN U17912 ( .B(clk), .A(\g.we_clk [14862]));
Q_ASSIGN U17913 ( .B(clk), .A(\g.we_clk [14861]));
Q_ASSIGN U17914 ( .B(clk), .A(\g.we_clk [14860]));
Q_ASSIGN U17915 ( .B(clk), .A(\g.we_clk [14859]));
Q_ASSIGN U17916 ( .B(clk), .A(\g.we_clk [14858]));
Q_ASSIGN U17917 ( .B(clk), .A(\g.we_clk [14857]));
Q_ASSIGN U17918 ( .B(clk), .A(\g.we_clk [14856]));
Q_ASSIGN U17919 ( .B(clk), .A(\g.we_clk [14855]));
Q_ASSIGN U17920 ( .B(clk), .A(\g.we_clk [14854]));
Q_ASSIGN U17921 ( .B(clk), .A(\g.we_clk [14853]));
Q_ASSIGN U17922 ( .B(clk), .A(\g.we_clk [14852]));
Q_ASSIGN U17923 ( .B(clk), .A(\g.we_clk [14851]));
Q_ASSIGN U17924 ( .B(clk), .A(\g.we_clk [14850]));
Q_ASSIGN U17925 ( .B(clk), .A(\g.we_clk [14849]));
Q_ASSIGN U17926 ( .B(clk), .A(\g.we_clk [14848]));
Q_ASSIGN U17927 ( .B(clk), .A(\g.we_clk [14847]));
Q_ASSIGN U17928 ( .B(clk), .A(\g.we_clk [14846]));
Q_ASSIGN U17929 ( .B(clk), .A(\g.we_clk [14845]));
Q_ASSIGN U17930 ( .B(clk), .A(\g.we_clk [14844]));
Q_ASSIGN U17931 ( .B(clk), .A(\g.we_clk [14843]));
Q_ASSIGN U17932 ( .B(clk), .A(\g.we_clk [14842]));
Q_ASSIGN U17933 ( .B(clk), .A(\g.we_clk [14841]));
Q_ASSIGN U17934 ( .B(clk), .A(\g.we_clk [14840]));
Q_ASSIGN U17935 ( .B(clk), .A(\g.we_clk [14839]));
Q_ASSIGN U17936 ( .B(clk), .A(\g.we_clk [14838]));
Q_ASSIGN U17937 ( .B(clk), .A(\g.we_clk [14837]));
Q_ASSIGN U17938 ( .B(clk), .A(\g.we_clk [14836]));
Q_ASSIGN U17939 ( .B(clk), .A(\g.we_clk [14835]));
Q_ASSIGN U17940 ( .B(clk), .A(\g.we_clk [14834]));
Q_ASSIGN U17941 ( .B(clk), .A(\g.we_clk [14833]));
Q_ASSIGN U17942 ( .B(clk), .A(\g.we_clk [14832]));
Q_ASSIGN U17943 ( .B(clk), .A(\g.we_clk [14831]));
Q_ASSIGN U17944 ( .B(clk), .A(\g.we_clk [14830]));
Q_ASSIGN U17945 ( .B(clk), .A(\g.we_clk [14829]));
Q_ASSIGN U17946 ( .B(clk), .A(\g.we_clk [14828]));
Q_ASSIGN U17947 ( .B(clk), .A(\g.we_clk [14827]));
Q_ASSIGN U17948 ( .B(clk), .A(\g.we_clk [14826]));
Q_ASSIGN U17949 ( .B(clk), .A(\g.we_clk [14825]));
Q_ASSIGN U17950 ( .B(clk), .A(\g.we_clk [14824]));
Q_ASSIGN U17951 ( .B(clk), .A(\g.we_clk [14823]));
Q_ASSIGN U17952 ( .B(clk), .A(\g.we_clk [14822]));
Q_ASSIGN U17953 ( .B(clk), .A(\g.we_clk [14821]));
Q_ASSIGN U17954 ( .B(clk), .A(\g.we_clk [14820]));
Q_ASSIGN U17955 ( .B(clk), .A(\g.we_clk [14819]));
Q_ASSIGN U17956 ( .B(clk), .A(\g.we_clk [14818]));
Q_ASSIGN U17957 ( .B(clk), .A(\g.we_clk [14817]));
Q_ASSIGN U17958 ( .B(clk), .A(\g.we_clk [14816]));
Q_ASSIGN U17959 ( .B(clk), .A(\g.we_clk [14815]));
Q_ASSIGN U17960 ( .B(clk), .A(\g.we_clk [14814]));
Q_ASSIGN U17961 ( .B(clk), .A(\g.we_clk [14813]));
Q_ASSIGN U17962 ( .B(clk), .A(\g.we_clk [14812]));
Q_ASSIGN U17963 ( .B(clk), .A(\g.we_clk [14811]));
Q_ASSIGN U17964 ( .B(clk), .A(\g.we_clk [14810]));
Q_ASSIGN U17965 ( .B(clk), .A(\g.we_clk [14809]));
Q_ASSIGN U17966 ( .B(clk), .A(\g.we_clk [14808]));
Q_ASSIGN U17967 ( .B(clk), .A(\g.we_clk [14807]));
Q_ASSIGN U17968 ( .B(clk), .A(\g.we_clk [14806]));
Q_ASSIGN U17969 ( .B(clk), .A(\g.we_clk [14805]));
Q_ASSIGN U17970 ( .B(clk), .A(\g.we_clk [14804]));
Q_ASSIGN U17971 ( .B(clk), .A(\g.we_clk [14803]));
Q_ASSIGN U17972 ( .B(clk), .A(\g.we_clk [14802]));
Q_ASSIGN U17973 ( .B(clk), .A(\g.we_clk [14801]));
Q_ASSIGN U17974 ( .B(clk), .A(\g.we_clk [14800]));
Q_ASSIGN U17975 ( .B(clk), .A(\g.we_clk [14799]));
Q_ASSIGN U17976 ( .B(clk), .A(\g.we_clk [14798]));
Q_ASSIGN U17977 ( .B(clk), .A(\g.we_clk [14797]));
Q_ASSIGN U17978 ( .B(clk), .A(\g.we_clk [14796]));
Q_ASSIGN U17979 ( .B(clk), .A(\g.we_clk [14795]));
Q_ASSIGN U17980 ( .B(clk), .A(\g.we_clk [14794]));
Q_ASSIGN U17981 ( .B(clk), .A(\g.we_clk [14793]));
Q_ASSIGN U17982 ( .B(clk), .A(\g.we_clk [14792]));
Q_ASSIGN U17983 ( .B(clk), .A(\g.we_clk [14791]));
Q_ASSIGN U17984 ( .B(clk), .A(\g.we_clk [14790]));
Q_ASSIGN U17985 ( .B(clk), .A(\g.we_clk [14789]));
Q_ASSIGN U17986 ( .B(clk), .A(\g.we_clk [14788]));
Q_ASSIGN U17987 ( .B(clk), .A(\g.we_clk [14787]));
Q_ASSIGN U17988 ( .B(clk), .A(\g.we_clk [14786]));
Q_ASSIGN U17989 ( .B(clk), .A(\g.we_clk [14785]));
Q_ASSIGN U17990 ( .B(clk), .A(\g.we_clk [14784]));
Q_ASSIGN U17991 ( .B(clk), .A(\g.we_clk [14783]));
Q_ASSIGN U17992 ( .B(clk), .A(\g.we_clk [14782]));
Q_ASSIGN U17993 ( .B(clk), .A(\g.we_clk [14781]));
Q_ASSIGN U17994 ( .B(clk), .A(\g.we_clk [14780]));
Q_ASSIGN U17995 ( .B(clk), .A(\g.we_clk [14779]));
Q_ASSIGN U17996 ( .B(clk), .A(\g.we_clk [14778]));
Q_ASSIGN U17997 ( .B(clk), .A(\g.we_clk [14777]));
Q_ASSIGN U17998 ( .B(clk), .A(\g.we_clk [14776]));
Q_ASSIGN U17999 ( .B(clk), .A(\g.we_clk [14775]));
Q_ASSIGN U18000 ( .B(clk), .A(\g.we_clk [14774]));
Q_ASSIGN U18001 ( .B(clk), .A(\g.we_clk [14773]));
Q_ASSIGN U18002 ( .B(clk), .A(\g.we_clk [14772]));
Q_ASSIGN U18003 ( .B(clk), .A(\g.we_clk [14771]));
Q_ASSIGN U18004 ( .B(clk), .A(\g.we_clk [14770]));
Q_ASSIGN U18005 ( .B(clk), .A(\g.we_clk [14769]));
Q_ASSIGN U18006 ( .B(clk), .A(\g.we_clk [14768]));
Q_ASSIGN U18007 ( .B(clk), .A(\g.we_clk [14767]));
Q_ASSIGN U18008 ( .B(clk), .A(\g.we_clk [14766]));
Q_ASSIGN U18009 ( .B(clk), .A(\g.we_clk [14765]));
Q_ASSIGN U18010 ( .B(clk), .A(\g.we_clk [14764]));
Q_ASSIGN U18011 ( .B(clk), .A(\g.we_clk [14763]));
Q_ASSIGN U18012 ( .B(clk), .A(\g.we_clk [14762]));
Q_ASSIGN U18013 ( .B(clk), .A(\g.we_clk [14761]));
Q_ASSIGN U18014 ( .B(clk), .A(\g.we_clk [14760]));
Q_ASSIGN U18015 ( .B(clk), .A(\g.we_clk [14759]));
Q_ASSIGN U18016 ( .B(clk), .A(\g.we_clk [14758]));
Q_ASSIGN U18017 ( .B(clk), .A(\g.we_clk [14757]));
Q_ASSIGN U18018 ( .B(clk), .A(\g.we_clk [14756]));
Q_ASSIGN U18019 ( .B(clk), .A(\g.we_clk [14755]));
Q_ASSIGN U18020 ( .B(clk), .A(\g.we_clk [14754]));
Q_ASSIGN U18021 ( .B(clk), .A(\g.we_clk [14753]));
Q_ASSIGN U18022 ( .B(clk), .A(\g.we_clk [14752]));
Q_ASSIGN U18023 ( .B(clk), .A(\g.we_clk [14751]));
Q_ASSIGN U18024 ( .B(clk), .A(\g.we_clk [14750]));
Q_ASSIGN U18025 ( .B(clk), .A(\g.we_clk [14749]));
Q_ASSIGN U18026 ( .B(clk), .A(\g.we_clk [14748]));
Q_ASSIGN U18027 ( .B(clk), .A(\g.we_clk [14747]));
Q_ASSIGN U18028 ( .B(clk), .A(\g.we_clk [14746]));
Q_ASSIGN U18029 ( .B(clk), .A(\g.we_clk [14745]));
Q_ASSIGN U18030 ( .B(clk), .A(\g.we_clk [14744]));
Q_ASSIGN U18031 ( .B(clk), .A(\g.we_clk [14743]));
Q_ASSIGN U18032 ( .B(clk), .A(\g.we_clk [14742]));
Q_ASSIGN U18033 ( .B(clk), .A(\g.we_clk [14741]));
Q_ASSIGN U18034 ( .B(clk), .A(\g.we_clk [14740]));
Q_ASSIGN U18035 ( .B(clk), .A(\g.we_clk [14739]));
Q_ASSIGN U18036 ( .B(clk), .A(\g.we_clk [14738]));
Q_ASSIGN U18037 ( .B(clk), .A(\g.we_clk [14737]));
Q_ASSIGN U18038 ( .B(clk), .A(\g.we_clk [14736]));
Q_ASSIGN U18039 ( .B(clk), .A(\g.we_clk [14735]));
Q_ASSIGN U18040 ( .B(clk), .A(\g.we_clk [14734]));
Q_ASSIGN U18041 ( .B(clk), .A(\g.we_clk [14733]));
Q_ASSIGN U18042 ( .B(clk), .A(\g.we_clk [14732]));
Q_ASSIGN U18043 ( .B(clk), .A(\g.we_clk [14731]));
Q_ASSIGN U18044 ( .B(clk), .A(\g.we_clk [14730]));
Q_ASSIGN U18045 ( .B(clk), .A(\g.we_clk [14729]));
Q_ASSIGN U18046 ( .B(clk), .A(\g.we_clk [14728]));
Q_ASSIGN U18047 ( .B(clk), .A(\g.we_clk [14727]));
Q_ASSIGN U18048 ( .B(clk), .A(\g.we_clk [14726]));
Q_ASSIGN U18049 ( .B(clk), .A(\g.we_clk [14725]));
Q_ASSIGN U18050 ( .B(clk), .A(\g.we_clk [14724]));
Q_ASSIGN U18051 ( .B(clk), .A(\g.we_clk [14723]));
Q_ASSIGN U18052 ( .B(clk), .A(\g.we_clk [14722]));
Q_ASSIGN U18053 ( .B(clk), .A(\g.we_clk [14721]));
Q_ASSIGN U18054 ( .B(clk), .A(\g.we_clk [14720]));
Q_ASSIGN U18055 ( .B(clk), .A(\g.we_clk [14719]));
Q_ASSIGN U18056 ( .B(clk), .A(\g.we_clk [14718]));
Q_ASSIGN U18057 ( .B(clk), .A(\g.we_clk [14717]));
Q_ASSIGN U18058 ( .B(clk), .A(\g.we_clk [14716]));
Q_ASSIGN U18059 ( .B(clk), .A(\g.we_clk [14715]));
Q_ASSIGN U18060 ( .B(clk), .A(\g.we_clk [14714]));
Q_ASSIGN U18061 ( .B(clk), .A(\g.we_clk [14713]));
Q_ASSIGN U18062 ( .B(clk), .A(\g.we_clk [14712]));
Q_ASSIGN U18063 ( .B(clk), .A(\g.we_clk [14711]));
Q_ASSIGN U18064 ( .B(clk), .A(\g.we_clk [14710]));
Q_ASSIGN U18065 ( .B(clk), .A(\g.we_clk [14709]));
Q_ASSIGN U18066 ( .B(clk), .A(\g.we_clk [14708]));
Q_ASSIGN U18067 ( .B(clk), .A(\g.we_clk [14707]));
Q_ASSIGN U18068 ( .B(clk), .A(\g.we_clk [14706]));
Q_ASSIGN U18069 ( .B(clk), .A(\g.we_clk [14705]));
Q_ASSIGN U18070 ( .B(clk), .A(\g.we_clk [14704]));
Q_ASSIGN U18071 ( .B(clk), .A(\g.we_clk [14703]));
Q_ASSIGN U18072 ( .B(clk), .A(\g.we_clk [14702]));
Q_ASSIGN U18073 ( .B(clk), .A(\g.we_clk [14701]));
Q_ASSIGN U18074 ( .B(clk), .A(\g.we_clk [14700]));
Q_ASSIGN U18075 ( .B(clk), .A(\g.we_clk [14699]));
Q_ASSIGN U18076 ( .B(clk), .A(\g.we_clk [14698]));
Q_ASSIGN U18077 ( .B(clk), .A(\g.we_clk [14697]));
Q_ASSIGN U18078 ( .B(clk), .A(\g.we_clk [14696]));
Q_ASSIGN U18079 ( .B(clk), .A(\g.we_clk [14695]));
Q_ASSIGN U18080 ( .B(clk), .A(\g.we_clk [14694]));
Q_ASSIGN U18081 ( .B(clk), .A(\g.we_clk [14693]));
Q_ASSIGN U18082 ( .B(clk), .A(\g.we_clk [14692]));
Q_ASSIGN U18083 ( .B(clk), .A(\g.we_clk [14691]));
Q_ASSIGN U18084 ( .B(clk), .A(\g.we_clk [14690]));
Q_ASSIGN U18085 ( .B(clk), .A(\g.we_clk [14689]));
Q_ASSIGN U18086 ( .B(clk), .A(\g.we_clk [14688]));
Q_ASSIGN U18087 ( .B(clk), .A(\g.we_clk [14687]));
Q_ASSIGN U18088 ( .B(clk), .A(\g.we_clk [14686]));
Q_ASSIGN U18089 ( .B(clk), .A(\g.we_clk [14685]));
Q_ASSIGN U18090 ( .B(clk), .A(\g.we_clk [14684]));
Q_ASSIGN U18091 ( .B(clk), .A(\g.we_clk [14683]));
Q_ASSIGN U18092 ( .B(clk), .A(\g.we_clk [14682]));
Q_ASSIGN U18093 ( .B(clk), .A(\g.we_clk [14681]));
Q_ASSIGN U18094 ( .B(clk), .A(\g.we_clk [14680]));
Q_ASSIGN U18095 ( .B(clk), .A(\g.we_clk [14679]));
Q_ASSIGN U18096 ( .B(clk), .A(\g.we_clk [14678]));
Q_ASSIGN U18097 ( .B(clk), .A(\g.we_clk [14677]));
Q_ASSIGN U18098 ( .B(clk), .A(\g.we_clk [14676]));
Q_ASSIGN U18099 ( .B(clk), .A(\g.we_clk [14675]));
Q_ASSIGN U18100 ( .B(clk), .A(\g.we_clk [14674]));
Q_ASSIGN U18101 ( .B(clk), .A(\g.we_clk [14673]));
Q_ASSIGN U18102 ( .B(clk), .A(\g.we_clk [14672]));
Q_ASSIGN U18103 ( .B(clk), .A(\g.we_clk [14671]));
Q_ASSIGN U18104 ( .B(clk), .A(\g.we_clk [14670]));
Q_ASSIGN U18105 ( .B(clk), .A(\g.we_clk [14669]));
Q_ASSIGN U18106 ( .B(clk), .A(\g.we_clk [14668]));
Q_ASSIGN U18107 ( .B(clk), .A(\g.we_clk [14667]));
Q_ASSIGN U18108 ( .B(clk), .A(\g.we_clk [14666]));
Q_ASSIGN U18109 ( .B(clk), .A(\g.we_clk [14665]));
Q_ASSIGN U18110 ( .B(clk), .A(\g.we_clk [14664]));
Q_ASSIGN U18111 ( .B(clk), .A(\g.we_clk [14663]));
Q_ASSIGN U18112 ( .B(clk), .A(\g.we_clk [14662]));
Q_ASSIGN U18113 ( .B(clk), .A(\g.we_clk [14661]));
Q_ASSIGN U18114 ( .B(clk), .A(\g.we_clk [14660]));
Q_ASSIGN U18115 ( .B(clk), .A(\g.we_clk [14659]));
Q_ASSIGN U18116 ( .B(clk), .A(\g.we_clk [14658]));
Q_ASSIGN U18117 ( .B(clk), .A(\g.we_clk [14657]));
Q_ASSIGN U18118 ( .B(clk), .A(\g.we_clk [14656]));
Q_ASSIGN U18119 ( .B(clk), .A(\g.we_clk [14655]));
Q_ASSIGN U18120 ( .B(clk), .A(\g.we_clk [14654]));
Q_ASSIGN U18121 ( .B(clk), .A(\g.we_clk [14653]));
Q_ASSIGN U18122 ( .B(clk), .A(\g.we_clk [14652]));
Q_ASSIGN U18123 ( .B(clk), .A(\g.we_clk [14651]));
Q_ASSIGN U18124 ( .B(clk), .A(\g.we_clk [14650]));
Q_ASSIGN U18125 ( .B(clk), .A(\g.we_clk [14649]));
Q_ASSIGN U18126 ( .B(clk), .A(\g.we_clk [14648]));
Q_ASSIGN U18127 ( .B(clk), .A(\g.we_clk [14647]));
Q_ASSIGN U18128 ( .B(clk), .A(\g.we_clk [14646]));
Q_ASSIGN U18129 ( .B(clk), .A(\g.we_clk [14645]));
Q_ASSIGN U18130 ( .B(clk), .A(\g.we_clk [14644]));
Q_ASSIGN U18131 ( .B(clk), .A(\g.we_clk [14643]));
Q_ASSIGN U18132 ( .B(clk), .A(\g.we_clk [14642]));
Q_ASSIGN U18133 ( .B(clk), .A(\g.we_clk [14641]));
Q_ASSIGN U18134 ( .B(clk), .A(\g.we_clk [14640]));
Q_ASSIGN U18135 ( .B(clk), .A(\g.we_clk [14639]));
Q_ASSIGN U18136 ( .B(clk), .A(\g.we_clk [14638]));
Q_ASSIGN U18137 ( .B(clk), .A(\g.we_clk [14637]));
Q_ASSIGN U18138 ( .B(clk), .A(\g.we_clk [14636]));
Q_ASSIGN U18139 ( .B(clk), .A(\g.we_clk [14635]));
Q_ASSIGN U18140 ( .B(clk), .A(\g.we_clk [14634]));
Q_ASSIGN U18141 ( .B(clk), .A(\g.we_clk [14633]));
Q_ASSIGN U18142 ( .B(clk), .A(\g.we_clk [14632]));
Q_ASSIGN U18143 ( .B(clk), .A(\g.we_clk [14631]));
Q_ASSIGN U18144 ( .B(clk), .A(\g.we_clk [14630]));
Q_ASSIGN U18145 ( .B(clk), .A(\g.we_clk [14629]));
Q_ASSIGN U18146 ( .B(clk), .A(\g.we_clk [14628]));
Q_ASSIGN U18147 ( .B(clk), .A(\g.we_clk [14627]));
Q_ASSIGN U18148 ( .B(clk), .A(\g.we_clk [14626]));
Q_ASSIGN U18149 ( .B(clk), .A(\g.we_clk [14625]));
Q_ASSIGN U18150 ( .B(clk), .A(\g.we_clk [14624]));
Q_ASSIGN U18151 ( .B(clk), .A(\g.we_clk [14623]));
Q_ASSIGN U18152 ( .B(clk), .A(\g.we_clk [14622]));
Q_ASSIGN U18153 ( .B(clk), .A(\g.we_clk [14621]));
Q_ASSIGN U18154 ( .B(clk), .A(\g.we_clk [14620]));
Q_ASSIGN U18155 ( .B(clk), .A(\g.we_clk [14619]));
Q_ASSIGN U18156 ( .B(clk), .A(\g.we_clk [14618]));
Q_ASSIGN U18157 ( .B(clk), .A(\g.we_clk [14617]));
Q_ASSIGN U18158 ( .B(clk), .A(\g.we_clk [14616]));
Q_ASSIGN U18159 ( .B(clk), .A(\g.we_clk [14615]));
Q_ASSIGN U18160 ( .B(clk), .A(\g.we_clk [14614]));
Q_ASSIGN U18161 ( .B(clk), .A(\g.we_clk [14613]));
Q_ASSIGN U18162 ( .B(clk), .A(\g.we_clk [14612]));
Q_ASSIGN U18163 ( .B(clk), .A(\g.we_clk [14611]));
Q_ASSIGN U18164 ( .B(clk), .A(\g.we_clk [14610]));
Q_ASSIGN U18165 ( .B(clk), .A(\g.we_clk [14609]));
Q_ASSIGN U18166 ( .B(clk), .A(\g.we_clk [14608]));
Q_ASSIGN U18167 ( .B(clk), .A(\g.we_clk [14607]));
Q_ASSIGN U18168 ( .B(clk), .A(\g.we_clk [14606]));
Q_ASSIGN U18169 ( .B(clk), .A(\g.we_clk [14605]));
Q_ASSIGN U18170 ( .B(clk), .A(\g.we_clk [14604]));
Q_ASSIGN U18171 ( .B(clk), .A(\g.we_clk [14603]));
Q_ASSIGN U18172 ( .B(clk), .A(\g.we_clk [14602]));
Q_ASSIGN U18173 ( .B(clk), .A(\g.we_clk [14601]));
Q_ASSIGN U18174 ( .B(clk), .A(\g.we_clk [14600]));
Q_ASSIGN U18175 ( .B(clk), .A(\g.we_clk [14599]));
Q_ASSIGN U18176 ( .B(clk), .A(\g.we_clk [14598]));
Q_ASSIGN U18177 ( .B(clk), .A(\g.we_clk [14597]));
Q_ASSIGN U18178 ( .B(clk), .A(\g.we_clk [14596]));
Q_ASSIGN U18179 ( .B(clk), .A(\g.we_clk [14595]));
Q_ASSIGN U18180 ( .B(clk), .A(\g.we_clk [14594]));
Q_ASSIGN U18181 ( .B(clk), .A(\g.we_clk [14593]));
Q_ASSIGN U18182 ( .B(clk), .A(\g.we_clk [14592]));
Q_ASSIGN U18183 ( .B(clk), .A(\g.we_clk [14591]));
Q_ASSIGN U18184 ( .B(clk), .A(\g.we_clk [14590]));
Q_ASSIGN U18185 ( .B(clk), .A(\g.we_clk [14589]));
Q_ASSIGN U18186 ( .B(clk), .A(\g.we_clk [14588]));
Q_ASSIGN U18187 ( .B(clk), .A(\g.we_clk [14587]));
Q_ASSIGN U18188 ( .B(clk), .A(\g.we_clk [14586]));
Q_ASSIGN U18189 ( .B(clk), .A(\g.we_clk [14585]));
Q_ASSIGN U18190 ( .B(clk), .A(\g.we_clk [14584]));
Q_ASSIGN U18191 ( .B(clk), .A(\g.we_clk [14583]));
Q_ASSIGN U18192 ( .B(clk), .A(\g.we_clk [14582]));
Q_ASSIGN U18193 ( .B(clk), .A(\g.we_clk [14581]));
Q_ASSIGN U18194 ( .B(clk), .A(\g.we_clk [14580]));
Q_ASSIGN U18195 ( .B(clk), .A(\g.we_clk [14579]));
Q_ASSIGN U18196 ( .B(clk), .A(\g.we_clk [14578]));
Q_ASSIGN U18197 ( .B(clk), .A(\g.we_clk [14577]));
Q_ASSIGN U18198 ( .B(clk), .A(\g.we_clk [14576]));
Q_ASSIGN U18199 ( .B(clk), .A(\g.we_clk [14575]));
Q_ASSIGN U18200 ( .B(clk), .A(\g.we_clk [14574]));
Q_ASSIGN U18201 ( .B(clk), .A(\g.we_clk [14573]));
Q_ASSIGN U18202 ( .B(clk), .A(\g.we_clk [14572]));
Q_ASSIGN U18203 ( .B(clk), .A(\g.we_clk [14571]));
Q_ASSIGN U18204 ( .B(clk), .A(\g.we_clk [14570]));
Q_ASSIGN U18205 ( .B(clk), .A(\g.we_clk [14569]));
Q_ASSIGN U18206 ( .B(clk), .A(\g.we_clk [14568]));
Q_ASSIGN U18207 ( .B(clk), .A(\g.we_clk [14567]));
Q_ASSIGN U18208 ( .B(clk), .A(\g.we_clk [14566]));
Q_ASSIGN U18209 ( .B(clk), .A(\g.we_clk [14565]));
Q_ASSIGN U18210 ( .B(clk), .A(\g.we_clk [14564]));
Q_ASSIGN U18211 ( .B(clk), .A(\g.we_clk [14563]));
Q_ASSIGN U18212 ( .B(clk), .A(\g.we_clk [14562]));
Q_ASSIGN U18213 ( .B(clk), .A(\g.we_clk [14561]));
Q_ASSIGN U18214 ( .B(clk), .A(\g.we_clk [14560]));
Q_ASSIGN U18215 ( .B(clk), .A(\g.we_clk [14559]));
Q_ASSIGN U18216 ( .B(clk), .A(\g.we_clk [14558]));
Q_ASSIGN U18217 ( .B(clk), .A(\g.we_clk [14557]));
Q_ASSIGN U18218 ( .B(clk), .A(\g.we_clk [14556]));
Q_ASSIGN U18219 ( .B(clk), .A(\g.we_clk [14555]));
Q_ASSIGN U18220 ( .B(clk), .A(\g.we_clk [14554]));
Q_ASSIGN U18221 ( .B(clk), .A(\g.we_clk [14553]));
Q_ASSIGN U18222 ( .B(clk), .A(\g.we_clk [14552]));
Q_ASSIGN U18223 ( .B(clk), .A(\g.we_clk [14551]));
Q_ASSIGN U18224 ( .B(clk), .A(\g.we_clk [14550]));
Q_ASSIGN U18225 ( .B(clk), .A(\g.we_clk [14549]));
Q_ASSIGN U18226 ( .B(clk), .A(\g.we_clk [14548]));
Q_ASSIGN U18227 ( .B(clk), .A(\g.we_clk [14547]));
Q_ASSIGN U18228 ( .B(clk), .A(\g.we_clk [14546]));
Q_ASSIGN U18229 ( .B(clk), .A(\g.we_clk [14545]));
Q_ASSIGN U18230 ( .B(clk), .A(\g.we_clk [14544]));
Q_ASSIGN U18231 ( .B(clk), .A(\g.we_clk [14543]));
Q_ASSIGN U18232 ( .B(clk), .A(\g.we_clk [14542]));
Q_ASSIGN U18233 ( .B(clk), .A(\g.we_clk [14541]));
Q_ASSIGN U18234 ( .B(clk), .A(\g.we_clk [14540]));
Q_ASSIGN U18235 ( .B(clk), .A(\g.we_clk [14539]));
Q_ASSIGN U18236 ( .B(clk), .A(\g.we_clk [14538]));
Q_ASSIGN U18237 ( .B(clk), .A(\g.we_clk [14537]));
Q_ASSIGN U18238 ( .B(clk), .A(\g.we_clk [14536]));
Q_ASSIGN U18239 ( .B(clk), .A(\g.we_clk [14535]));
Q_ASSIGN U18240 ( .B(clk), .A(\g.we_clk [14534]));
Q_ASSIGN U18241 ( .B(clk), .A(\g.we_clk [14533]));
Q_ASSIGN U18242 ( .B(clk), .A(\g.we_clk [14532]));
Q_ASSIGN U18243 ( .B(clk), .A(\g.we_clk [14531]));
Q_ASSIGN U18244 ( .B(clk), .A(\g.we_clk [14530]));
Q_ASSIGN U18245 ( .B(clk), .A(\g.we_clk [14529]));
Q_ASSIGN U18246 ( .B(clk), .A(\g.we_clk [14528]));
Q_ASSIGN U18247 ( .B(clk), .A(\g.we_clk [14527]));
Q_ASSIGN U18248 ( .B(clk), .A(\g.we_clk [14526]));
Q_ASSIGN U18249 ( .B(clk), .A(\g.we_clk [14525]));
Q_ASSIGN U18250 ( .B(clk), .A(\g.we_clk [14524]));
Q_ASSIGN U18251 ( .B(clk), .A(\g.we_clk [14523]));
Q_ASSIGN U18252 ( .B(clk), .A(\g.we_clk [14522]));
Q_ASSIGN U18253 ( .B(clk), .A(\g.we_clk [14521]));
Q_ASSIGN U18254 ( .B(clk), .A(\g.we_clk [14520]));
Q_ASSIGN U18255 ( .B(clk), .A(\g.we_clk [14519]));
Q_ASSIGN U18256 ( .B(clk), .A(\g.we_clk [14518]));
Q_ASSIGN U18257 ( .B(clk), .A(\g.we_clk [14517]));
Q_ASSIGN U18258 ( .B(clk), .A(\g.we_clk [14516]));
Q_ASSIGN U18259 ( .B(clk), .A(\g.we_clk [14515]));
Q_ASSIGN U18260 ( .B(clk), .A(\g.we_clk [14514]));
Q_ASSIGN U18261 ( .B(clk), .A(\g.we_clk [14513]));
Q_ASSIGN U18262 ( .B(clk), .A(\g.we_clk [14512]));
Q_ASSIGN U18263 ( .B(clk), .A(\g.we_clk [14511]));
Q_ASSIGN U18264 ( .B(clk), .A(\g.we_clk [14510]));
Q_ASSIGN U18265 ( .B(clk), .A(\g.we_clk [14509]));
Q_ASSIGN U18266 ( .B(clk), .A(\g.we_clk [14508]));
Q_ASSIGN U18267 ( .B(clk), .A(\g.we_clk [14507]));
Q_ASSIGN U18268 ( .B(clk), .A(\g.we_clk [14506]));
Q_ASSIGN U18269 ( .B(clk), .A(\g.we_clk [14505]));
Q_ASSIGN U18270 ( .B(clk), .A(\g.we_clk [14504]));
Q_ASSIGN U18271 ( .B(clk), .A(\g.we_clk [14503]));
Q_ASSIGN U18272 ( .B(clk), .A(\g.we_clk [14502]));
Q_ASSIGN U18273 ( .B(clk), .A(\g.we_clk [14501]));
Q_ASSIGN U18274 ( .B(clk), .A(\g.we_clk [14500]));
Q_ASSIGN U18275 ( .B(clk), .A(\g.we_clk [14499]));
Q_ASSIGN U18276 ( .B(clk), .A(\g.we_clk [14498]));
Q_ASSIGN U18277 ( .B(clk), .A(\g.we_clk [14497]));
Q_ASSIGN U18278 ( .B(clk), .A(\g.we_clk [14496]));
Q_ASSIGN U18279 ( .B(clk), .A(\g.we_clk [14495]));
Q_ASSIGN U18280 ( .B(clk), .A(\g.we_clk [14494]));
Q_ASSIGN U18281 ( .B(clk), .A(\g.we_clk [14493]));
Q_ASSIGN U18282 ( .B(clk), .A(\g.we_clk [14492]));
Q_ASSIGN U18283 ( .B(clk), .A(\g.we_clk [14491]));
Q_ASSIGN U18284 ( .B(clk), .A(\g.we_clk [14490]));
Q_ASSIGN U18285 ( .B(clk), .A(\g.we_clk [14489]));
Q_ASSIGN U18286 ( .B(clk), .A(\g.we_clk [14488]));
Q_ASSIGN U18287 ( .B(clk), .A(\g.we_clk [14487]));
Q_ASSIGN U18288 ( .B(clk), .A(\g.we_clk [14486]));
Q_ASSIGN U18289 ( .B(clk), .A(\g.we_clk [14485]));
Q_ASSIGN U18290 ( .B(clk), .A(\g.we_clk [14484]));
Q_ASSIGN U18291 ( .B(clk), .A(\g.we_clk [14483]));
Q_ASSIGN U18292 ( .B(clk), .A(\g.we_clk [14482]));
Q_ASSIGN U18293 ( .B(clk), .A(\g.we_clk [14481]));
Q_ASSIGN U18294 ( .B(clk), .A(\g.we_clk [14480]));
Q_ASSIGN U18295 ( .B(clk), .A(\g.we_clk [14479]));
Q_ASSIGN U18296 ( .B(clk), .A(\g.we_clk [14478]));
Q_ASSIGN U18297 ( .B(clk), .A(\g.we_clk [14477]));
Q_ASSIGN U18298 ( .B(clk), .A(\g.we_clk [14476]));
Q_ASSIGN U18299 ( .B(clk), .A(\g.we_clk [14475]));
Q_ASSIGN U18300 ( .B(clk), .A(\g.we_clk [14474]));
Q_ASSIGN U18301 ( .B(clk), .A(\g.we_clk [14473]));
Q_ASSIGN U18302 ( .B(clk), .A(\g.we_clk [14472]));
Q_ASSIGN U18303 ( .B(clk), .A(\g.we_clk [14471]));
Q_ASSIGN U18304 ( .B(clk), .A(\g.we_clk [14470]));
Q_ASSIGN U18305 ( .B(clk), .A(\g.we_clk [14469]));
Q_ASSIGN U18306 ( .B(clk), .A(\g.we_clk [14468]));
Q_ASSIGN U18307 ( .B(clk), .A(\g.we_clk [14467]));
Q_ASSIGN U18308 ( .B(clk), .A(\g.we_clk [14466]));
Q_ASSIGN U18309 ( .B(clk), .A(\g.we_clk [14465]));
Q_ASSIGN U18310 ( .B(clk), .A(\g.we_clk [14464]));
Q_ASSIGN U18311 ( .B(clk), .A(\g.we_clk [14463]));
Q_ASSIGN U18312 ( .B(clk), .A(\g.we_clk [14462]));
Q_ASSIGN U18313 ( .B(clk), .A(\g.we_clk [14461]));
Q_ASSIGN U18314 ( .B(clk), .A(\g.we_clk [14460]));
Q_ASSIGN U18315 ( .B(clk), .A(\g.we_clk [14459]));
Q_ASSIGN U18316 ( .B(clk), .A(\g.we_clk [14458]));
Q_ASSIGN U18317 ( .B(clk), .A(\g.we_clk [14457]));
Q_ASSIGN U18318 ( .B(clk), .A(\g.we_clk [14456]));
Q_ASSIGN U18319 ( .B(clk), .A(\g.we_clk [14455]));
Q_ASSIGN U18320 ( .B(clk), .A(\g.we_clk [14454]));
Q_ASSIGN U18321 ( .B(clk), .A(\g.we_clk [14453]));
Q_ASSIGN U18322 ( .B(clk), .A(\g.we_clk [14452]));
Q_ASSIGN U18323 ( .B(clk), .A(\g.we_clk [14451]));
Q_ASSIGN U18324 ( .B(clk), .A(\g.we_clk [14450]));
Q_ASSIGN U18325 ( .B(clk), .A(\g.we_clk [14449]));
Q_ASSIGN U18326 ( .B(clk), .A(\g.we_clk [14448]));
Q_ASSIGN U18327 ( .B(clk), .A(\g.we_clk [14447]));
Q_ASSIGN U18328 ( .B(clk), .A(\g.we_clk [14446]));
Q_ASSIGN U18329 ( .B(clk), .A(\g.we_clk [14445]));
Q_ASSIGN U18330 ( .B(clk), .A(\g.we_clk [14444]));
Q_ASSIGN U18331 ( .B(clk), .A(\g.we_clk [14443]));
Q_ASSIGN U18332 ( .B(clk), .A(\g.we_clk [14442]));
Q_ASSIGN U18333 ( .B(clk), .A(\g.we_clk [14441]));
Q_ASSIGN U18334 ( .B(clk), .A(\g.we_clk [14440]));
Q_ASSIGN U18335 ( .B(clk), .A(\g.we_clk [14439]));
Q_ASSIGN U18336 ( .B(clk), .A(\g.we_clk [14438]));
Q_ASSIGN U18337 ( .B(clk), .A(\g.we_clk [14437]));
Q_ASSIGN U18338 ( .B(clk), .A(\g.we_clk [14436]));
Q_ASSIGN U18339 ( .B(clk), .A(\g.we_clk [14435]));
Q_ASSIGN U18340 ( .B(clk), .A(\g.we_clk [14434]));
Q_ASSIGN U18341 ( .B(clk), .A(\g.we_clk [14433]));
Q_ASSIGN U18342 ( .B(clk), .A(\g.we_clk [14432]));
Q_ASSIGN U18343 ( .B(clk), .A(\g.we_clk [14431]));
Q_ASSIGN U18344 ( .B(clk), .A(\g.we_clk [14430]));
Q_ASSIGN U18345 ( .B(clk), .A(\g.we_clk [14429]));
Q_ASSIGN U18346 ( .B(clk), .A(\g.we_clk [14428]));
Q_ASSIGN U18347 ( .B(clk), .A(\g.we_clk [14427]));
Q_ASSIGN U18348 ( .B(clk), .A(\g.we_clk [14426]));
Q_ASSIGN U18349 ( .B(clk), .A(\g.we_clk [14425]));
Q_ASSIGN U18350 ( .B(clk), .A(\g.we_clk [14424]));
Q_ASSIGN U18351 ( .B(clk), .A(\g.we_clk [14423]));
Q_ASSIGN U18352 ( .B(clk), .A(\g.we_clk [14422]));
Q_ASSIGN U18353 ( .B(clk), .A(\g.we_clk [14421]));
Q_ASSIGN U18354 ( .B(clk), .A(\g.we_clk [14420]));
Q_ASSIGN U18355 ( .B(clk), .A(\g.we_clk [14419]));
Q_ASSIGN U18356 ( .B(clk), .A(\g.we_clk [14418]));
Q_ASSIGN U18357 ( .B(clk), .A(\g.we_clk [14417]));
Q_ASSIGN U18358 ( .B(clk), .A(\g.we_clk [14416]));
Q_ASSIGN U18359 ( .B(clk), .A(\g.we_clk [14415]));
Q_ASSIGN U18360 ( .B(clk), .A(\g.we_clk [14414]));
Q_ASSIGN U18361 ( .B(clk), .A(\g.we_clk [14413]));
Q_ASSIGN U18362 ( .B(clk), .A(\g.we_clk [14412]));
Q_ASSIGN U18363 ( .B(clk), .A(\g.we_clk [14411]));
Q_ASSIGN U18364 ( .B(clk), .A(\g.we_clk [14410]));
Q_ASSIGN U18365 ( .B(clk), .A(\g.we_clk [14409]));
Q_ASSIGN U18366 ( .B(clk), .A(\g.we_clk [14408]));
Q_ASSIGN U18367 ( .B(clk), .A(\g.we_clk [14407]));
Q_ASSIGN U18368 ( .B(clk), .A(\g.we_clk [14406]));
Q_ASSIGN U18369 ( .B(clk), .A(\g.we_clk [14405]));
Q_ASSIGN U18370 ( .B(clk), .A(\g.we_clk [14404]));
Q_ASSIGN U18371 ( .B(clk), .A(\g.we_clk [14403]));
Q_ASSIGN U18372 ( .B(clk), .A(\g.we_clk [14402]));
Q_ASSIGN U18373 ( .B(clk), .A(\g.we_clk [14401]));
Q_ASSIGN U18374 ( .B(clk), .A(\g.we_clk [14400]));
Q_ASSIGN U18375 ( .B(clk), .A(\g.we_clk [14399]));
Q_ASSIGN U18376 ( .B(clk), .A(\g.we_clk [14398]));
Q_ASSIGN U18377 ( .B(clk), .A(\g.we_clk [14397]));
Q_ASSIGN U18378 ( .B(clk), .A(\g.we_clk [14396]));
Q_ASSIGN U18379 ( .B(clk), .A(\g.we_clk [14395]));
Q_ASSIGN U18380 ( .B(clk), .A(\g.we_clk [14394]));
Q_ASSIGN U18381 ( .B(clk), .A(\g.we_clk [14393]));
Q_ASSIGN U18382 ( .B(clk), .A(\g.we_clk [14392]));
Q_ASSIGN U18383 ( .B(clk), .A(\g.we_clk [14391]));
Q_ASSIGN U18384 ( .B(clk), .A(\g.we_clk [14390]));
Q_ASSIGN U18385 ( .B(clk), .A(\g.we_clk [14389]));
Q_ASSIGN U18386 ( .B(clk), .A(\g.we_clk [14388]));
Q_ASSIGN U18387 ( .B(clk), .A(\g.we_clk [14387]));
Q_ASSIGN U18388 ( .B(clk), .A(\g.we_clk [14386]));
Q_ASSIGN U18389 ( .B(clk), .A(\g.we_clk [14385]));
Q_ASSIGN U18390 ( .B(clk), .A(\g.we_clk [14384]));
Q_ASSIGN U18391 ( .B(clk), .A(\g.we_clk [14383]));
Q_ASSIGN U18392 ( .B(clk), .A(\g.we_clk [14382]));
Q_ASSIGN U18393 ( .B(clk), .A(\g.we_clk [14381]));
Q_ASSIGN U18394 ( .B(clk), .A(\g.we_clk [14380]));
Q_ASSIGN U18395 ( .B(clk), .A(\g.we_clk [14379]));
Q_ASSIGN U18396 ( .B(clk), .A(\g.we_clk [14378]));
Q_ASSIGN U18397 ( .B(clk), .A(\g.we_clk [14377]));
Q_ASSIGN U18398 ( .B(clk), .A(\g.we_clk [14376]));
Q_ASSIGN U18399 ( .B(clk), .A(\g.we_clk [14375]));
Q_ASSIGN U18400 ( .B(clk), .A(\g.we_clk [14374]));
Q_ASSIGN U18401 ( .B(clk), .A(\g.we_clk [14373]));
Q_ASSIGN U18402 ( .B(clk), .A(\g.we_clk [14372]));
Q_ASSIGN U18403 ( .B(clk), .A(\g.we_clk [14371]));
Q_ASSIGN U18404 ( .B(clk), .A(\g.we_clk [14370]));
Q_ASSIGN U18405 ( .B(clk), .A(\g.we_clk [14369]));
Q_ASSIGN U18406 ( .B(clk), .A(\g.we_clk [14368]));
Q_ASSIGN U18407 ( .B(clk), .A(\g.we_clk [14367]));
Q_ASSIGN U18408 ( .B(clk), .A(\g.we_clk [14366]));
Q_ASSIGN U18409 ( .B(clk), .A(\g.we_clk [14365]));
Q_ASSIGN U18410 ( .B(clk), .A(\g.we_clk [14364]));
Q_ASSIGN U18411 ( .B(clk), .A(\g.we_clk [14363]));
Q_ASSIGN U18412 ( .B(clk), .A(\g.we_clk [14362]));
Q_ASSIGN U18413 ( .B(clk), .A(\g.we_clk [14361]));
Q_ASSIGN U18414 ( .B(clk), .A(\g.we_clk [14360]));
Q_ASSIGN U18415 ( .B(clk), .A(\g.we_clk [14359]));
Q_ASSIGN U18416 ( .B(clk), .A(\g.we_clk [14358]));
Q_ASSIGN U18417 ( .B(clk), .A(\g.we_clk [14357]));
Q_ASSIGN U18418 ( .B(clk), .A(\g.we_clk [14356]));
Q_ASSIGN U18419 ( .B(clk), .A(\g.we_clk [14355]));
Q_ASSIGN U18420 ( .B(clk), .A(\g.we_clk [14354]));
Q_ASSIGN U18421 ( .B(clk), .A(\g.we_clk [14353]));
Q_ASSIGN U18422 ( .B(clk), .A(\g.we_clk [14352]));
Q_ASSIGN U18423 ( .B(clk), .A(\g.we_clk [14351]));
Q_ASSIGN U18424 ( .B(clk), .A(\g.we_clk [14350]));
Q_ASSIGN U18425 ( .B(clk), .A(\g.we_clk [14349]));
Q_ASSIGN U18426 ( .B(clk), .A(\g.we_clk [14348]));
Q_ASSIGN U18427 ( .B(clk), .A(\g.we_clk [14347]));
Q_ASSIGN U18428 ( .B(clk), .A(\g.we_clk [14346]));
Q_ASSIGN U18429 ( .B(clk), .A(\g.we_clk [14345]));
Q_ASSIGN U18430 ( .B(clk), .A(\g.we_clk [14344]));
Q_ASSIGN U18431 ( .B(clk), .A(\g.we_clk [14343]));
Q_ASSIGN U18432 ( .B(clk), .A(\g.we_clk [14342]));
Q_ASSIGN U18433 ( .B(clk), .A(\g.we_clk [14341]));
Q_ASSIGN U18434 ( .B(clk), .A(\g.we_clk [14340]));
Q_ASSIGN U18435 ( .B(clk), .A(\g.we_clk [14339]));
Q_ASSIGN U18436 ( .B(clk), .A(\g.we_clk [14338]));
Q_ASSIGN U18437 ( .B(clk), .A(\g.we_clk [14337]));
Q_ASSIGN U18438 ( .B(clk), .A(\g.we_clk [14336]));
Q_ASSIGN U18439 ( .B(clk), .A(\g.we_clk [14335]));
Q_ASSIGN U18440 ( .B(clk), .A(\g.we_clk [14334]));
Q_ASSIGN U18441 ( .B(clk), .A(\g.we_clk [14333]));
Q_ASSIGN U18442 ( .B(clk), .A(\g.we_clk [14332]));
Q_ASSIGN U18443 ( .B(clk), .A(\g.we_clk [14331]));
Q_ASSIGN U18444 ( .B(clk), .A(\g.we_clk [14330]));
Q_ASSIGN U18445 ( .B(clk), .A(\g.we_clk [14329]));
Q_ASSIGN U18446 ( .B(clk), .A(\g.we_clk [14328]));
Q_ASSIGN U18447 ( .B(clk), .A(\g.we_clk [14327]));
Q_ASSIGN U18448 ( .B(clk), .A(\g.we_clk [14326]));
Q_ASSIGN U18449 ( .B(clk), .A(\g.we_clk [14325]));
Q_ASSIGN U18450 ( .B(clk), .A(\g.we_clk [14324]));
Q_ASSIGN U18451 ( .B(clk), .A(\g.we_clk [14323]));
Q_ASSIGN U18452 ( .B(clk), .A(\g.we_clk [14322]));
Q_ASSIGN U18453 ( .B(clk), .A(\g.we_clk [14321]));
Q_ASSIGN U18454 ( .B(clk), .A(\g.we_clk [14320]));
Q_ASSIGN U18455 ( .B(clk), .A(\g.we_clk [14319]));
Q_ASSIGN U18456 ( .B(clk), .A(\g.we_clk [14318]));
Q_ASSIGN U18457 ( .B(clk), .A(\g.we_clk [14317]));
Q_ASSIGN U18458 ( .B(clk), .A(\g.we_clk [14316]));
Q_ASSIGN U18459 ( .B(clk), .A(\g.we_clk [14315]));
Q_ASSIGN U18460 ( .B(clk), .A(\g.we_clk [14314]));
Q_ASSIGN U18461 ( .B(clk), .A(\g.we_clk [14313]));
Q_ASSIGN U18462 ( .B(clk), .A(\g.we_clk [14312]));
Q_ASSIGN U18463 ( .B(clk), .A(\g.we_clk [14311]));
Q_ASSIGN U18464 ( .B(clk), .A(\g.we_clk [14310]));
Q_ASSIGN U18465 ( .B(clk), .A(\g.we_clk [14309]));
Q_ASSIGN U18466 ( .B(clk), .A(\g.we_clk [14308]));
Q_ASSIGN U18467 ( .B(clk), .A(\g.we_clk [14307]));
Q_ASSIGN U18468 ( .B(clk), .A(\g.we_clk [14306]));
Q_ASSIGN U18469 ( .B(clk), .A(\g.we_clk [14305]));
Q_ASSIGN U18470 ( .B(clk), .A(\g.we_clk [14304]));
Q_ASSIGN U18471 ( .B(clk), .A(\g.we_clk [14303]));
Q_ASSIGN U18472 ( .B(clk), .A(\g.we_clk [14302]));
Q_ASSIGN U18473 ( .B(clk), .A(\g.we_clk [14301]));
Q_ASSIGN U18474 ( .B(clk), .A(\g.we_clk [14300]));
Q_ASSIGN U18475 ( .B(clk), .A(\g.we_clk [14299]));
Q_ASSIGN U18476 ( .B(clk), .A(\g.we_clk [14298]));
Q_ASSIGN U18477 ( .B(clk), .A(\g.we_clk [14297]));
Q_ASSIGN U18478 ( .B(clk), .A(\g.we_clk [14296]));
Q_ASSIGN U18479 ( .B(clk), .A(\g.we_clk [14295]));
Q_ASSIGN U18480 ( .B(clk), .A(\g.we_clk [14294]));
Q_ASSIGN U18481 ( .B(clk), .A(\g.we_clk [14293]));
Q_ASSIGN U18482 ( .B(clk), .A(\g.we_clk [14292]));
Q_ASSIGN U18483 ( .B(clk), .A(\g.we_clk [14291]));
Q_ASSIGN U18484 ( .B(clk), .A(\g.we_clk [14290]));
Q_ASSIGN U18485 ( .B(clk), .A(\g.we_clk [14289]));
Q_ASSIGN U18486 ( .B(clk), .A(\g.we_clk [14288]));
Q_ASSIGN U18487 ( .B(clk), .A(\g.we_clk [14287]));
Q_ASSIGN U18488 ( .B(clk), .A(\g.we_clk [14286]));
Q_ASSIGN U18489 ( .B(clk), .A(\g.we_clk [14285]));
Q_ASSIGN U18490 ( .B(clk), .A(\g.we_clk [14284]));
Q_ASSIGN U18491 ( .B(clk), .A(\g.we_clk [14283]));
Q_ASSIGN U18492 ( .B(clk), .A(\g.we_clk [14282]));
Q_ASSIGN U18493 ( .B(clk), .A(\g.we_clk [14281]));
Q_ASSIGN U18494 ( .B(clk), .A(\g.we_clk [14280]));
Q_ASSIGN U18495 ( .B(clk), .A(\g.we_clk [14279]));
Q_ASSIGN U18496 ( .B(clk), .A(\g.we_clk [14278]));
Q_ASSIGN U18497 ( .B(clk), .A(\g.we_clk [14277]));
Q_ASSIGN U18498 ( .B(clk), .A(\g.we_clk [14276]));
Q_ASSIGN U18499 ( .B(clk), .A(\g.we_clk [14275]));
Q_ASSIGN U18500 ( .B(clk), .A(\g.we_clk [14274]));
Q_ASSIGN U18501 ( .B(clk), .A(\g.we_clk [14273]));
Q_ASSIGN U18502 ( .B(clk), .A(\g.we_clk [14272]));
Q_ASSIGN U18503 ( .B(clk), .A(\g.we_clk [14271]));
Q_ASSIGN U18504 ( .B(clk), .A(\g.we_clk [14270]));
Q_ASSIGN U18505 ( .B(clk), .A(\g.we_clk [14269]));
Q_ASSIGN U18506 ( .B(clk), .A(\g.we_clk [14268]));
Q_ASSIGN U18507 ( .B(clk), .A(\g.we_clk [14267]));
Q_ASSIGN U18508 ( .B(clk), .A(\g.we_clk [14266]));
Q_ASSIGN U18509 ( .B(clk), .A(\g.we_clk [14265]));
Q_ASSIGN U18510 ( .B(clk), .A(\g.we_clk [14264]));
Q_ASSIGN U18511 ( .B(clk), .A(\g.we_clk [14263]));
Q_ASSIGN U18512 ( .B(clk), .A(\g.we_clk [14262]));
Q_ASSIGN U18513 ( .B(clk), .A(\g.we_clk [14261]));
Q_ASSIGN U18514 ( .B(clk), .A(\g.we_clk [14260]));
Q_ASSIGN U18515 ( .B(clk), .A(\g.we_clk [14259]));
Q_ASSIGN U18516 ( .B(clk), .A(\g.we_clk [14258]));
Q_ASSIGN U18517 ( .B(clk), .A(\g.we_clk [14257]));
Q_ASSIGN U18518 ( .B(clk), .A(\g.we_clk [14256]));
Q_ASSIGN U18519 ( .B(clk), .A(\g.we_clk [14255]));
Q_ASSIGN U18520 ( .B(clk), .A(\g.we_clk [14254]));
Q_ASSIGN U18521 ( .B(clk), .A(\g.we_clk [14253]));
Q_ASSIGN U18522 ( .B(clk), .A(\g.we_clk [14252]));
Q_ASSIGN U18523 ( .B(clk), .A(\g.we_clk [14251]));
Q_ASSIGN U18524 ( .B(clk), .A(\g.we_clk [14250]));
Q_ASSIGN U18525 ( .B(clk), .A(\g.we_clk [14249]));
Q_ASSIGN U18526 ( .B(clk), .A(\g.we_clk [14248]));
Q_ASSIGN U18527 ( .B(clk), .A(\g.we_clk [14247]));
Q_ASSIGN U18528 ( .B(clk), .A(\g.we_clk [14246]));
Q_ASSIGN U18529 ( .B(clk), .A(\g.we_clk [14245]));
Q_ASSIGN U18530 ( .B(clk), .A(\g.we_clk [14244]));
Q_ASSIGN U18531 ( .B(clk), .A(\g.we_clk [14243]));
Q_ASSIGN U18532 ( .B(clk), .A(\g.we_clk [14242]));
Q_ASSIGN U18533 ( .B(clk), .A(\g.we_clk [14241]));
Q_ASSIGN U18534 ( .B(clk), .A(\g.we_clk [14240]));
Q_ASSIGN U18535 ( .B(clk), .A(\g.we_clk [14239]));
Q_ASSIGN U18536 ( .B(clk), .A(\g.we_clk [14238]));
Q_ASSIGN U18537 ( .B(clk), .A(\g.we_clk [14237]));
Q_ASSIGN U18538 ( .B(clk), .A(\g.we_clk [14236]));
Q_ASSIGN U18539 ( .B(clk), .A(\g.we_clk [14235]));
Q_ASSIGN U18540 ( .B(clk), .A(\g.we_clk [14234]));
Q_ASSIGN U18541 ( .B(clk), .A(\g.we_clk [14233]));
Q_ASSIGN U18542 ( .B(clk), .A(\g.we_clk [14232]));
Q_ASSIGN U18543 ( .B(clk), .A(\g.we_clk [14231]));
Q_ASSIGN U18544 ( .B(clk), .A(\g.we_clk [14230]));
Q_ASSIGN U18545 ( .B(clk), .A(\g.we_clk [14229]));
Q_ASSIGN U18546 ( .B(clk), .A(\g.we_clk [14228]));
Q_ASSIGN U18547 ( .B(clk), .A(\g.we_clk [14227]));
Q_ASSIGN U18548 ( .B(clk), .A(\g.we_clk [14226]));
Q_ASSIGN U18549 ( .B(clk), .A(\g.we_clk [14225]));
Q_ASSIGN U18550 ( .B(clk), .A(\g.we_clk [14224]));
Q_ASSIGN U18551 ( .B(clk), .A(\g.we_clk [14223]));
Q_ASSIGN U18552 ( .B(clk), .A(\g.we_clk [14222]));
Q_ASSIGN U18553 ( .B(clk), .A(\g.we_clk [14221]));
Q_ASSIGN U18554 ( .B(clk), .A(\g.we_clk [14220]));
Q_ASSIGN U18555 ( .B(clk), .A(\g.we_clk [14219]));
Q_ASSIGN U18556 ( .B(clk), .A(\g.we_clk [14218]));
Q_ASSIGN U18557 ( .B(clk), .A(\g.we_clk [14217]));
Q_ASSIGN U18558 ( .B(clk), .A(\g.we_clk [14216]));
Q_ASSIGN U18559 ( .B(clk), .A(\g.we_clk [14215]));
Q_ASSIGN U18560 ( .B(clk), .A(\g.we_clk [14214]));
Q_ASSIGN U18561 ( .B(clk), .A(\g.we_clk [14213]));
Q_ASSIGN U18562 ( .B(clk), .A(\g.we_clk [14212]));
Q_ASSIGN U18563 ( .B(clk), .A(\g.we_clk [14211]));
Q_ASSIGN U18564 ( .B(clk), .A(\g.we_clk [14210]));
Q_ASSIGN U18565 ( .B(clk), .A(\g.we_clk [14209]));
Q_ASSIGN U18566 ( .B(clk), .A(\g.we_clk [14208]));
Q_ASSIGN U18567 ( .B(clk), .A(\g.we_clk [14207]));
Q_ASSIGN U18568 ( .B(clk), .A(\g.we_clk [14206]));
Q_ASSIGN U18569 ( .B(clk), .A(\g.we_clk [14205]));
Q_ASSIGN U18570 ( .B(clk), .A(\g.we_clk [14204]));
Q_ASSIGN U18571 ( .B(clk), .A(\g.we_clk [14203]));
Q_ASSIGN U18572 ( .B(clk), .A(\g.we_clk [14202]));
Q_ASSIGN U18573 ( .B(clk), .A(\g.we_clk [14201]));
Q_ASSIGN U18574 ( .B(clk), .A(\g.we_clk [14200]));
Q_ASSIGN U18575 ( .B(clk), .A(\g.we_clk [14199]));
Q_ASSIGN U18576 ( .B(clk), .A(\g.we_clk [14198]));
Q_ASSIGN U18577 ( .B(clk), .A(\g.we_clk [14197]));
Q_ASSIGN U18578 ( .B(clk), .A(\g.we_clk [14196]));
Q_ASSIGN U18579 ( .B(clk), .A(\g.we_clk [14195]));
Q_ASSIGN U18580 ( .B(clk), .A(\g.we_clk [14194]));
Q_ASSIGN U18581 ( .B(clk), .A(\g.we_clk [14193]));
Q_ASSIGN U18582 ( .B(clk), .A(\g.we_clk [14192]));
Q_ASSIGN U18583 ( .B(clk), .A(\g.we_clk [14191]));
Q_ASSIGN U18584 ( .B(clk), .A(\g.we_clk [14190]));
Q_ASSIGN U18585 ( .B(clk), .A(\g.we_clk [14189]));
Q_ASSIGN U18586 ( .B(clk), .A(\g.we_clk [14188]));
Q_ASSIGN U18587 ( .B(clk), .A(\g.we_clk [14187]));
Q_ASSIGN U18588 ( .B(clk), .A(\g.we_clk [14186]));
Q_ASSIGN U18589 ( .B(clk), .A(\g.we_clk [14185]));
Q_ASSIGN U18590 ( .B(clk), .A(\g.we_clk [14184]));
Q_ASSIGN U18591 ( .B(clk), .A(\g.we_clk [14183]));
Q_ASSIGN U18592 ( .B(clk), .A(\g.we_clk [14182]));
Q_ASSIGN U18593 ( .B(clk), .A(\g.we_clk [14181]));
Q_ASSIGN U18594 ( .B(clk), .A(\g.we_clk [14180]));
Q_ASSIGN U18595 ( .B(clk), .A(\g.we_clk [14179]));
Q_ASSIGN U18596 ( .B(clk), .A(\g.we_clk [14178]));
Q_ASSIGN U18597 ( .B(clk), .A(\g.we_clk [14177]));
Q_ASSIGN U18598 ( .B(clk), .A(\g.we_clk [14176]));
Q_ASSIGN U18599 ( .B(clk), .A(\g.we_clk [14175]));
Q_ASSIGN U18600 ( .B(clk), .A(\g.we_clk [14174]));
Q_ASSIGN U18601 ( .B(clk), .A(\g.we_clk [14173]));
Q_ASSIGN U18602 ( .B(clk), .A(\g.we_clk [14172]));
Q_ASSIGN U18603 ( .B(clk), .A(\g.we_clk [14171]));
Q_ASSIGN U18604 ( .B(clk), .A(\g.we_clk [14170]));
Q_ASSIGN U18605 ( .B(clk), .A(\g.we_clk [14169]));
Q_ASSIGN U18606 ( .B(clk), .A(\g.we_clk [14168]));
Q_ASSIGN U18607 ( .B(clk), .A(\g.we_clk [14167]));
Q_ASSIGN U18608 ( .B(clk), .A(\g.we_clk [14166]));
Q_ASSIGN U18609 ( .B(clk), .A(\g.we_clk [14165]));
Q_ASSIGN U18610 ( .B(clk), .A(\g.we_clk [14164]));
Q_ASSIGN U18611 ( .B(clk), .A(\g.we_clk [14163]));
Q_ASSIGN U18612 ( .B(clk), .A(\g.we_clk [14162]));
Q_ASSIGN U18613 ( .B(clk), .A(\g.we_clk [14161]));
Q_ASSIGN U18614 ( .B(clk), .A(\g.we_clk [14160]));
Q_ASSIGN U18615 ( .B(clk), .A(\g.we_clk [14159]));
Q_ASSIGN U18616 ( .B(clk), .A(\g.we_clk [14158]));
Q_ASSIGN U18617 ( .B(clk), .A(\g.we_clk [14157]));
Q_ASSIGN U18618 ( .B(clk), .A(\g.we_clk [14156]));
Q_ASSIGN U18619 ( .B(clk), .A(\g.we_clk [14155]));
Q_ASSIGN U18620 ( .B(clk), .A(\g.we_clk [14154]));
Q_ASSIGN U18621 ( .B(clk), .A(\g.we_clk [14153]));
Q_ASSIGN U18622 ( .B(clk), .A(\g.we_clk [14152]));
Q_ASSIGN U18623 ( .B(clk), .A(\g.we_clk [14151]));
Q_ASSIGN U18624 ( .B(clk), .A(\g.we_clk [14150]));
Q_ASSIGN U18625 ( .B(clk), .A(\g.we_clk [14149]));
Q_ASSIGN U18626 ( .B(clk), .A(\g.we_clk [14148]));
Q_ASSIGN U18627 ( .B(clk), .A(\g.we_clk [14147]));
Q_ASSIGN U18628 ( .B(clk), .A(\g.we_clk [14146]));
Q_ASSIGN U18629 ( .B(clk), .A(\g.we_clk [14145]));
Q_ASSIGN U18630 ( .B(clk), .A(\g.we_clk [14144]));
Q_ASSIGN U18631 ( .B(clk), .A(\g.we_clk [14143]));
Q_ASSIGN U18632 ( .B(clk), .A(\g.we_clk [14142]));
Q_ASSIGN U18633 ( .B(clk), .A(\g.we_clk [14141]));
Q_ASSIGN U18634 ( .B(clk), .A(\g.we_clk [14140]));
Q_ASSIGN U18635 ( .B(clk), .A(\g.we_clk [14139]));
Q_ASSIGN U18636 ( .B(clk), .A(\g.we_clk [14138]));
Q_ASSIGN U18637 ( .B(clk), .A(\g.we_clk [14137]));
Q_ASSIGN U18638 ( .B(clk), .A(\g.we_clk [14136]));
Q_ASSIGN U18639 ( .B(clk), .A(\g.we_clk [14135]));
Q_ASSIGN U18640 ( .B(clk), .A(\g.we_clk [14134]));
Q_ASSIGN U18641 ( .B(clk), .A(\g.we_clk [14133]));
Q_ASSIGN U18642 ( .B(clk), .A(\g.we_clk [14132]));
Q_ASSIGN U18643 ( .B(clk), .A(\g.we_clk [14131]));
Q_ASSIGN U18644 ( .B(clk), .A(\g.we_clk [14130]));
Q_ASSIGN U18645 ( .B(clk), .A(\g.we_clk [14129]));
Q_ASSIGN U18646 ( .B(clk), .A(\g.we_clk [14128]));
Q_ASSIGN U18647 ( .B(clk), .A(\g.we_clk [14127]));
Q_ASSIGN U18648 ( .B(clk), .A(\g.we_clk [14126]));
Q_ASSIGN U18649 ( .B(clk), .A(\g.we_clk [14125]));
Q_ASSIGN U18650 ( .B(clk), .A(\g.we_clk [14124]));
Q_ASSIGN U18651 ( .B(clk), .A(\g.we_clk [14123]));
Q_ASSIGN U18652 ( .B(clk), .A(\g.we_clk [14122]));
Q_ASSIGN U18653 ( .B(clk), .A(\g.we_clk [14121]));
Q_ASSIGN U18654 ( .B(clk), .A(\g.we_clk [14120]));
Q_ASSIGN U18655 ( .B(clk), .A(\g.we_clk [14119]));
Q_ASSIGN U18656 ( .B(clk), .A(\g.we_clk [14118]));
Q_ASSIGN U18657 ( .B(clk), .A(\g.we_clk [14117]));
Q_ASSIGN U18658 ( .B(clk), .A(\g.we_clk [14116]));
Q_ASSIGN U18659 ( .B(clk), .A(\g.we_clk [14115]));
Q_ASSIGN U18660 ( .B(clk), .A(\g.we_clk [14114]));
Q_ASSIGN U18661 ( .B(clk), .A(\g.we_clk [14113]));
Q_ASSIGN U18662 ( .B(clk), .A(\g.we_clk [14112]));
Q_ASSIGN U18663 ( .B(clk), .A(\g.we_clk [14111]));
Q_ASSIGN U18664 ( .B(clk), .A(\g.we_clk [14110]));
Q_ASSIGN U18665 ( .B(clk), .A(\g.we_clk [14109]));
Q_ASSIGN U18666 ( .B(clk), .A(\g.we_clk [14108]));
Q_ASSIGN U18667 ( .B(clk), .A(\g.we_clk [14107]));
Q_ASSIGN U18668 ( .B(clk), .A(\g.we_clk [14106]));
Q_ASSIGN U18669 ( .B(clk), .A(\g.we_clk [14105]));
Q_ASSIGN U18670 ( .B(clk), .A(\g.we_clk [14104]));
Q_ASSIGN U18671 ( .B(clk), .A(\g.we_clk [14103]));
Q_ASSIGN U18672 ( .B(clk), .A(\g.we_clk [14102]));
Q_ASSIGN U18673 ( .B(clk), .A(\g.we_clk [14101]));
Q_ASSIGN U18674 ( .B(clk), .A(\g.we_clk [14100]));
Q_ASSIGN U18675 ( .B(clk), .A(\g.we_clk [14099]));
Q_ASSIGN U18676 ( .B(clk), .A(\g.we_clk [14098]));
Q_ASSIGN U18677 ( .B(clk), .A(\g.we_clk [14097]));
Q_ASSIGN U18678 ( .B(clk), .A(\g.we_clk [14096]));
Q_ASSIGN U18679 ( .B(clk), .A(\g.we_clk [14095]));
Q_ASSIGN U18680 ( .B(clk), .A(\g.we_clk [14094]));
Q_ASSIGN U18681 ( .B(clk), .A(\g.we_clk [14093]));
Q_ASSIGN U18682 ( .B(clk), .A(\g.we_clk [14092]));
Q_ASSIGN U18683 ( .B(clk), .A(\g.we_clk [14091]));
Q_ASSIGN U18684 ( .B(clk), .A(\g.we_clk [14090]));
Q_ASSIGN U18685 ( .B(clk), .A(\g.we_clk [14089]));
Q_ASSIGN U18686 ( .B(clk), .A(\g.we_clk [14088]));
Q_ASSIGN U18687 ( .B(clk), .A(\g.we_clk [14087]));
Q_ASSIGN U18688 ( .B(clk), .A(\g.we_clk [14086]));
Q_ASSIGN U18689 ( .B(clk), .A(\g.we_clk [14085]));
Q_ASSIGN U18690 ( .B(clk), .A(\g.we_clk [14084]));
Q_ASSIGN U18691 ( .B(clk), .A(\g.we_clk [14083]));
Q_ASSIGN U18692 ( .B(clk), .A(\g.we_clk [14082]));
Q_ASSIGN U18693 ( .B(clk), .A(\g.we_clk [14081]));
Q_ASSIGN U18694 ( .B(clk), .A(\g.we_clk [14080]));
Q_ASSIGN U18695 ( .B(clk), .A(\g.we_clk [14079]));
Q_ASSIGN U18696 ( .B(clk), .A(\g.we_clk [14078]));
Q_ASSIGN U18697 ( .B(clk), .A(\g.we_clk [14077]));
Q_ASSIGN U18698 ( .B(clk), .A(\g.we_clk [14076]));
Q_ASSIGN U18699 ( .B(clk), .A(\g.we_clk [14075]));
Q_ASSIGN U18700 ( .B(clk), .A(\g.we_clk [14074]));
Q_ASSIGN U18701 ( .B(clk), .A(\g.we_clk [14073]));
Q_ASSIGN U18702 ( .B(clk), .A(\g.we_clk [14072]));
Q_ASSIGN U18703 ( .B(clk), .A(\g.we_clk [14071]));
Q_ASSIGN U18704 ( .B(clk), .A(\g.we_clk [14070]));
Q_ASSIGN U18705 ( .B(clk), .A(\g.we_clk [14069]));
Q_ASSIGN U18706 ( .B(clk), .A(\g.we_clk [14068]));
Q_ASSIGN U18707 ( .B(clk), .A(\g.we_clk [14067]));
Q_ASSIGN U18708 ( .B(clk), .A(\g.we_clk [14066]));
Q_ASSIGN U18709 ( .B(clk), .A(\g.we_clk [14065]));
Q_ASSIGN U18710 ( .B(clk), .A(\g.we_clk [14064]));
Q_ASSIGN U18711 ( .B(clk), .A(\g.we_clk [14063]));
Q_ASSIGN U18712 ( .B(clk), .A(\g.we_clk [14062]));
Q_ASSIGN U18713 ( .B(clk), .A(\g.we_clk [14061]));
Q_ASSIGN U18714 ( .B(clk), .A(\g.we_clk [14060]));
Q_ASSIGN U18715 ( .B(clk), .A(\g.we_clk [14059]));
Q_ASSIGN U18716 ( .B(clk), .A(\g.we_clk [14058]));
Q_ASSIGN U18717 ( .B(clk), .A(\g.we_clk [14057]));
Q_ASSIGN U18718 ( .B(clk), .A(\g.we_clk [14056]));
Q_ASSIGN U18719 ( .B(clk), .A(\g.we_clk [14055]));
Q_ASSIGN U18720 ( .B(clk), .A(\g.we_clk [14054]));
Q_ASSIGN U18721 ( .B(clk), .A(\g.we_clk [14053]));
Q_ASSIGN U18722 ( .B(clk), .A(\g.we_clk [14052]));
Q_ASSIGN U18723 ( .B(clk), .A(\g.we_clk [14051]));
Q_ASSIGN U18724 ( .B(clk), .A(\g.we_clk [14050]));
Q_ASSIGN U18725 ( .B(clk), .A(\g.we_clk [14049]));
Q_ASSIGN U18726 ( .B(clk), .A(\g.we_clk [14048]));
Q_ASSIGN U18727 ( .B(clk), .A(\g.we_clk [14047]));
Q_ASSIGN U18728 ( .B(clk), .A(\g.we_clk [14046]));
Q_ASSIGN U18729 ( .B(clk), .A(\g.we_clk [14045]));
Q_ASSIGN U18730 ( .B(clk), .A(\g.we_clk [14044]));
Q_ASSIGN U18731 ( .B(clk), .A(\g.we_clk [14043]));
Q_ASSIGN U18732 ( .B(clk), .A(\g.we_clk [14042]));
Q_ASSIGN U18733 ( .B(clk), .A(\g.we_clk [14041]));
Q_ASSIGN U18734 ( .B(clk), .A(\g.we_clk [14040]));
Q_ASSIGN U18735 ( .B(clk), .A(\g.we_clk [14039]));
Q_ASSIGN U18736 ( .B(clk), .A(\g.we_clk [14038]));
Q_ASSIGN U18737 ( .B(clk), .A(\g.we_clk [14037]));
Q_ASSIGN U18738 ( .B(clk), .A(\g.we_clk [14036]));
Q_ASSIGN U18739 ( .B(clk), .A(\g.we_clk [14035]));
Q_ASSIGN U18740 ( .B(clk), .A(\g.we_clk [14034]));
Q_ASSIGN U18741 ( .B(clk), .A(\g.we_clk [14033]));
Q_ASSIGN U18742 ( .B(clk), .A(\g.we_clk [14032]));
Q_ASSIGN U18743 ( .B(clk), .A(\g.we_clk [14031]));
Q_ASSIGN U18744 ( .B(clk), .A(\g.we_clk [14030]));
Q_ASSIGN U18745 ( .B(clk), .A(\g.we_clk [14029]));
Q_ASSIGN U18746 ( .B(clk), .A(\g.we_clk [14028]));
Q_ASSIGN U18747 ( .B(clk), .A(\g.we_clk [14027]));
Q_ASSIGN U18748 ( .B(clk), .A(\g.we_clk [14026]));
Q_ASSIGN U18749 ( .B(clk), .A(\g.we_clk [14025]));
Q_ASSIGN U18750 ( .B(clk), .A(\g.we_clk [14024]));
Q_ASSIGN U18751 ( .B(clk), .A(\g.we_clk [14023]));
Q_ASSIGN U18752 ( .B(clk), .A(\g.we_clk [14022]));
Q_ASSIGN U18753 ( .B(clk), .A(\g.we_clk [14021]));
Q_ASSIGN U18754 ( .B(clk), .A(\g.we_clk [14020]));
Q_ASSIGN U18755 ( .B(clk), .A(\g.we_clk [14019]));
Q_ASSIGN U18756 ( .B(clk), .A(\g.we_clk [14018]));
Q_ASSIGN U18757 ( .B(clk), .A(\g.we_clk [14017]));
Q_ASSIGN U18758 ( .B(clk), .A(\g.we_clk [14016]));
Q_ASSIGN U18759 ( .B(clk), .A(\g.we_clk [14015]));
Q_ASSIGN U18760 ( .B(clk), .A(\g.we_clk [14014]));
Q_ASSIGN U18761 ( .B(clk), .A(\g.we_clk [14013]));
Q_ASSIGN U18762 ( .B(clk), .A(\g.we_clk [14012]));
Q_ASSIGN U18763 ( .B(clk), .A(\g.we_clk [14011]));
Q_ASSIGN U18764 ( .B(clk), .A(\g.we_clk [14010]));
Q_ASSIGN U18765 ( .B(clk), .A(\g.we_clk [14009]));
Q_ASSIGN U18766 ( .B(clk), .A(\g.we_clk [14008]));
Q_ASSIGN U18767 ( .B(clk), .A(\g.we_clk [14007]));
Q_ASSIGN U18768 ( .B(clk), .A(\g.we_clk [14006]));
Q_ASSIGN U18769 ( .B(clk), .A(\g.we_clk [14005]));
Q_ASSIGN U18770 ( .B(clk), .A(\g.we_clk [14004]));
Q_ASSIGN U18771 ( .B(clk), .A(\g.we_clk [14003]));
Q_ASSIGN U18772 ( .B(clk), .A(\g.we_clk [14002]));
Q_ASSIGN U18773 ( .B(clk), .A(\g.we_clk [14001]));
Q_ASSIGN U18774 ( .B(clk), .A(\g.we_clk [14000]));
Q_ASSIGN U18775 ( .B(clk), .A(\g.we_clk [13999]));
Q_ASSIGN U18776 ( .B(clk), .A(\g.we_clk [13998]));
Q_ASSIGN U18777 ( .B(clk), .A(\g.we_clk [13997]));
Q_ASSIGN U18778 ( .B(clk), .A(\g.we_clk [13996]));
Q_ASSIGN U18779 ( .B(clk), .A(\g.we_clk [13995]));
Q_ASSIGN U18780 ( .B(clk), .A(\g.we_clk [13994]));
Q_ASSIGN U18781 ( .B(clk), .A(\g.we_clk [13993]));
Q_ASSIGN U18782 ( .B(clk), .A(\g.we_clk [13992]));
Q_ASSIGN U18783 ( .B(clk), .A(\g.we_clk [13991]));
Q_ASSIGN U18784 ( .B(clk), .A(\g.we_clk [13990]));
Q_ASSIGN U18785 ( .B(clk), .A(\g.we_clk [13989]));
Q_ASSIGN U18786 ( .B(clk), .A(\g.we_clk [13988]));
Q_ASSIGN U18787 ( .B(clk), .A(\g.we_clk [13987]));
Q_ASSIGN U18788 ( .B(clk), .A(\g.we_clk [13986]));
Q_ASSIGN U18789 ( .B(clk), .A(\g.we_clk [13985]));
Q_ASSIGN U18790 ( .B(clk), .A(\g.we_clk [13984]));
Q_ASSIGN U18791 ( .B(clk), .A(\g.we_clk [13983]));
Q_ASSIGN U18792 ( .B(clk), .A(\g.we_clk [13982]));
Q_ASSIGN U18793 ( .B(clk), .A(\g.we_clk [13981]));
Q_ASSIGN U18794 ( .B(clk), .A(\g.we_clk [13980]));
Q_ASSIGN U18795 ( .B(clk), .A(\g.we_clk [13979]));
Q_ASSIGN U18796 ( .B(clk), .A(\g.we_clk [13978]));
Q_ASSIGN U18797 ( .B(clk), .A(\g.we_clk [13977]));
Q_ASSIGN U18798 ( .B(clk), .A(\g.we_clk [13976]));
Q_ASSIGN U18799 ( .B(clk), .A(\g.we_clk [13975]));
Q_ASSIGN U18800 ( .B(clk), .A(\g.we_clk [13974]));
Q_ASSIGN U18801 ( .B(clk), .A(\g.we_clk [13973]));
Q_ASSIGN U18802 ( .B(clk), .A(\g.we_clk [13972]));
Q_ASSIGN U18803 ( .B(clk), .A(\g.we_clk [13971]));
Q_ASSIGN U18804 ( .B(clk), .A(\g.we_clk [13970]));
Q_ASSIGN U18805 ( .B(clk), .A(\g.we_clk [13969]));
Q_ASSIGN U18806 ( .B(clk), .A(\g.we_clk [13968]));
Q_ASSIGN U18807 ( .B(clk), .A(\g.we_clk [13967]));
Q_ASSIGN U18808 ( .B(clk), .A(\g.we_clk [13966]));
Q_ASSIGN U18809 ( .B(clk), .A(\g.we_clk [13965]));
Q_ASSIGN U18810 ( .B(clk), .A(\g.we_clk [13964]));
Q_ASSIGN U18811 ( .B(clk), .A(\g.we_clk [13963]));
Q_ASSIGN U18812 ( .B(clk), .A(\g.we_clk [13962]));
Q_ASSIGN U18813 ( .B(clk), .A(\g.we_clk [13961]));
Q_ASSIGN U18814 ( .B(clk), .A(\g.we_clk [13960]));
Q_ASSIGN U18815 ( .B(clk), .A(\g.we_clk [13959]));
Q_ASSIGN U18816 ( .B(clk), .A(\g.we_clk [13958]));
Q_ASSIGN U18817 ( .B(clk), .A(\g.we_clk [13957]));
Q_ASSIGN U18818 ( .B(clk), .A(\g.we_clk [13956]));
Q_ASSIGN U18819 ( .B(clk), .A(\g.we_clk [13955]));
Q_ASSIGN U18820 ( .B(clk), .A(\g.we_clk [13954]));
Q_ASSIGN U18821 ( .B(clk), .A(\g.we_clk [13953]));
Q_ASSIGN U18822 ( .B(clk), .A(\g.we_clk [13952]));
Q_ASSIGN U18823 ( .B(clk), .A(\g.we_clk [13951]));
Q_ASSIGN U18824 ( .B(clk), .A(\g.we_clk [13950]));
Q_ASSIGN U18825 ( .B(clk), .A(\g.we_clk [13949]));
Q_ASSIGN U18826 ( .B(clk), .A(\g.we_clk [13948]));
Q_ASSIGN U18827 ( .B(clk), .A(\g.we_clk [13947]));
Q_ASSIGN U18828 ( .B(clk), .A(\g.we_clk [13946]));
Q_ASSIGN U18829 ( .B(clk), .A(\g.we_clk [13945]));
Q_ASSIGN U18830 ( .B(clk), .A(\g.we_clk [13944]));
Q_ASSIGN U18831 ( .B(clk), .A(\g.we_clk [13943]));
Q_ASSIGN U18832 ( .B(clk), .A(\g.we_clk [13942]));
Q_ASSIGN U18833 ( .B(clk), .A(\g.we_clk [13941]));
Q_ASSIGN U18834 ( .B(clk), .A(\g.we_clk [13940]));
Q_ASSIGN U18835 ( .B(clk), .A(\g.we_clk [13939]));
Q_ASSIGN U18836 ( .B(clk), .A(\g.we_clk [13938]));
Q_ASSIGN U18837 ( .B(clk), .A(\g.we_clk [13937]));
Q_ASSIGN U18838 ( .B(clk), .A(\g.we_clk [13936]));
Q_ASSIGN U18839 ( .B(clk), .A(\g.we_clk [13935]));
Q_ASSIGN U18840 ( .B(clk), .A(\g.we_clk [13934]));
Q_ASSIGN U18841 ( .B(clk), .A(\g.we_clk [13933]));
Q_ASSIGN U18842 ( .B(clk), .A(\g.we_clk [13932]));
Q_ASSIGN U18843 ( .B(clk), .A(\g.we_clk [13931]));
Q_ASSIGN U18844 ( .B(clk), .A(\g.we_clk [13930]));
Q_ASSIGN U18845 ( .B(clk), .A(\g.we_clk [13929]));
Q_ASSIGN U18846 ( .B(clk), .A(\g.we_clk [13928]));
Q_ASSIGN U18847 ( .B(clk), .A(\g.we_clk [13927]));
Q_ASSIGN U18848 ( .B(clk), .A(\g.we_clk [13926]));
Q_ASSIGN U18849 ( .B(clk), .A(\g.we_clk [13925]));
Q_ASSIGN U18850 ( .B(clk), .A(\g.we_clk [13924]));
Q_ASSIGN U18851 ( .B(clk), .A(\g.we_clk [13923]));
Q_ASSIGN U18852 ( .B(clk), .A(\g.we_clk [13922]));
Q_ASSIGN U18853 ( .B(clk), .A(\g.we_clk [13921]));
Q_ASSIGN U18854 ( .B(clk), .A(\g.we_clk [13920]));
Q_ASSIGN U18855 ( .B(clk), .A(\g.we_clk [13919]));
Q_ASSIGN U18856 ( .B(clk), .A(\g.we_clk [13918]));
Q_ASSIGN U18857 ( .B(clk), .A(\g.we_clk [13917]));
Q_ASSIGN U18858 ( .B(clk), .A(\g.we_clk [13916]));
Q_ASSIGN U18859 ( .B(clk), .A(\g.we_clk [13915]));
Q_ASSIGN U18860 ( .B(clk), .A(\g.we_clk [13914]));
Q_ASSIGN U18861 ( .B(clk), .A(\g.we_clk [13913]));
Q_ASSIGN U18862 ( .B(clk), .A(\g.we_clk [13912]));
Q_ASSIGN U18863 ( .B(clk), .A(\g.we_clk [13911]));
Q_ASSIGN U18864 ( .B(clk), .A(\g.we_clk [13910]));
Q_ASSIGN U18865 ( .B(clk), .A(\g.we_clk [13909]));
Q_ASSIGN U18866 ( .B(clk), .A(\g.we_clk [13908]));
Q_ASSIGN U18867 ( .B(clk), .A(\g.we_clk [13907]));
Q_ASSIGN U18868 ( .B(clk), .A(\g.we_clk [13906]));
Q_ASSIGN U18869 ( .B(clk), .A(\g.we_clk [13905]));
Q_ASSIGN U18870 ( .B(clk), .A(\g.we_clk [13904]));
Q_ASSIGN U18871 ( .B(clk), .A(\g.we_clk [13903]));
Q_ASSIGN U18872 ( .B(clk), .A(\g.we_clk [13902]));
Q_ASSIGN U18873 ( .B(clk), .A(\g.we_clk [13901]));
Q_ASSIGN U18874 ( .B(clk), .A(\g.we_clk [13900]));
Q_ASSIGN U18875 ( .B(clk), .A(\g.we_clk [13899]));
Q_ASSIGN U18876 ( .B(clk), .A(\g.we_clk [13898]));
Q_ASSIGN U18877 ( .B(clk), .A(\g.we_clk [13897]));
Q_ASSIGN U18878 ( .B(clk), .A(\g.we_clk [13896]));
Q_ASSIGN U18879 ( .B(clk), .A(\g.we_clk [13895]));
Q_ASSIGN U18880 ( .B(clk), .A(\g.we_clk [13894]));
Q_ASSIGN U18881 ( .B(clk), .A(\g.we_clk [13893]));
Q_ASSIGN U18882 ( .B(clk), .A(\g.we_clk [13892]));
Q_ASSIGN U18883 ( .B(clk), .A(\g.we_clk [13891]));
Q_ASSIGN U18884 ( .B(clk), .A(\g.we_clk [13890]));
Q_ASSIGN U18885 ( .B(clk), .A(\g.we_clk [13889]));
Q_ASSIGN U18886 ( .B(clk), .A(\g.we_clk [13888]));
Q_ASSIGN U18887 ( .B(clk), .A(\g.we_clk [13887]));
Q_ASSIGN U18888 ( .B(clk), .A(\g.we_clk [13886]));
Q_ASSIGN U18889 ( .B(clk), .A(\g.we_clk [13885]));
Q_ASSIGN U18890 ( .B(clk), .A(\g.we_clk [13884]));
Q_ASSIGN U18891 ( .B(clk), .A(\g.we_clk [13883]));
Q_ASSIGN U18892 ( .B(clk), .A(\g.we_clk [13882]));
Q_ASSIGN U18893 ( .B(clk), .A(\g.we_clk [13881]));
Q_ASSIGN U18894 ( .B(clk), .A(\g.we_clk [13880]));
Q_ASSIGN U18895 ( .B(clk), .A(\g.we_clk [13879]));
Q_ASSIGN U18896 ( .B(clk), .A(\g.we_clk [13878]));
Q_ASSIGN U18897 ( .B(clk), .A(\g.we_clk [13877]));
Q_ASSIGN U18898 ( .B(clk), .A(\g.we_clk [13876]));
Q_ASSIGN U18899 ( .B(clk), .A(\g.we_clk [13875]));
Q_ASSIGN U18900 ( .B(clk), .A(\g.we_clk [13874]));
Q_ASSIGN U18901 ( .B(clk), .A(\g.we_clk [13873]));
Q_ASSIGN U18902 ( .B(clk), .A(\g.we_clk [13872]));
Q_ASSIGN U18903 ( .B(clk), .A(\g.we_clk [13871]));
Q_ASSIGN U18904 ( .B(clk), .A(\g.we_clk [13870]));
Q_ASSIGN U18905 ( .B(clk), .A(\g.we_clk [13869]));
Q_ASSIGN U18906 ( .B(clk), .A(\g.we_clk [13868]));
Q_ASSIGN U18907 ( .B(clk), .A(\g.we_clk [13867]));
Q_ASSIGN U18908 ( .B(clk), .A(\g.we_clk [13866]));
Q_ASSIGN U18909 ( .B(clk), .A(\g.we_clk [13865]));
Q_ASSIGN U18910 ( .B(clk), .A(\g.we_clk [13864]));
Q_ASSIGN U18911 ( .B(clk), .A(\g.we_clk [13863]));
Q_ASSIGN U18912 ( .B(clk), .A(\g.we_clk [13862]));
Q_ASSIGN U18913 ( .B(clk), .A(\g.we_clk [13861]));
Q_ASSIGN U18914 ( .B(clk), .A(\g.we_clk [13860]));
Q_ASSIGN U18915 ( .B(clk), .A(\g.we_clk [13859]));
Q_ASSIGN U18916 ( .B(clk), .A(\g.we_clk [13858]));
Q_ASSIGN U18917 ( .B(clk), .A(\g.we_clk [13857]));
Q_ASSIGN U18918 ( .B(clk), .A(\g.we_clk [13856]));
Q_ASSIGN U18919 ( .B(clk), .A(\g.we_clk [13855]));
Q_ASSIGN U18920 ( .B(clk), .A(\g.we_clk [13854]));
Q_ASSIGN U18921 ( .B(clk), .A(\g.we_clk [13853]));
Q_ASSIGN U18922 ( .B(clk), .A(\g.we_clk [13852]));
Q_ASSIGN U18923 ( .B(clk), .A(\g.we_clk [13851]));
Q_ASSIGN U18924 ( .B(clk), .A(\g.we_clk [13850]));
Q_ASSIGN U18925 ( .B(clk), .A(\g.we_clk [13849]));
Q_ASSIGN U18926 ( .B(clk), .A(\g.we_clk [13848]));
Q_ASSIGN U18927 ( .B(clk), .A(\g.we_clk [13847]));
Q_ASSIGN U18928 ( .B(clk), .A(\g.we_clk [13846]));
Q_ASSIGN U18929 ( .B(clk), .A(\g.we_clk [13845]));
Q_ASSIGN U18930 ( .B(clk), .A(\g.we_clk [13844]));
Q_ASSIGN U18931 ( .B(clk), .A(\g.we_clk [13843]));
Q_ASSIGN U18932 ( .B(clk), .A(\g.we_clk [13842]));
Q_ASSIGN U18933 ( .B(clk), .A(\g.we_clk [13841]));
Q_ASSIGN U18934 ( .B(clk), .A(\g.we_clk [13840]));
Q_ASSIGN U18935 ( .B(clk), .A(\g.we_clk [13839]));
Q_ASSIGN U18936 ( .B(clk), .A(\g.we_clk [13838]));
Q_ASSIGN U18937 ( .B(clk), .A(\g.we_clk [13837]));
Q_ASSIGN U18938 ( .B(clk), .A(\g.we_clk [13836]));
Q_ASSIGN U18939 ( .B(clk), .A(\g.we_clk [13835]));
Q_ASSIGN U18940 ( .B(clk), .A(\g.we_clk [13834]));
Q_ASSIGN U18941 ( .B(clk), .A(\g.we_clk [13833]));
Q_ASSIGN U18942 ( .B(clk), .A(\g.we_clk [13832]));
Q_ASSIGN U18943 ( .B(clk), .A(\g.we_clk [13831]));
Q_ASSIGN U18944 ( .B(clk), .A(\g.we_clk [13830]));
Q_ASSIGN U18945 ( .B(clk), .A(\g.we_clk [13829]));
Q_ASSIGN U18946 ( .B(clk), .A(\g.we_clk [13828]));
Q_ASSIGN U18947 ( .B(clk), .A(\g.we_clk [13827]));
Q_ASSIGN U18948 ( .B(clk), .A(\g.we_clk [13826]));
Q_ASSIGN U18949 ( .B(clk), .A(\g.we_clk [13825]));
Q_ASSIGN U18950 ( .B(clk), .A(\g.we_clk [13824]));
Q_ASSIGN U18951 ( .B(clk), .A(\g.we_clk [13823]));
Q_ASSIGN U18952 ( .B(clk), .A(\g.we_clk [13822]));
Q_ASSIGN U18953 ( .B(clk), .A(\g.we_clk [13821]));
Q_ASSIGN U18954 ( .B(clk), .A(\g.we_clk [13820]));
Q_ASSIGN U18955 ( .B(clk), .A(\g.we_clk [13819]));
Q_ASSIGN U18956 ( .B(clk), .A(\g.we_clk [13818]));
Q_ASSIGN U18957 ( .B(clk), .A(\g.we_clk [13817]));
Q_ASSIGN U18958 ( .B(clk), .A(\g.we_clk [13816]));
Q_ASSIGN U18959 ( .B(clk), .A(\g.we_clk [13815]));
Q_ASSIGN U18960 ( .B(clk), .A(\g.we_clk [13814]));
Q_ASSIGN U18961 ( .B(clk), .A(\g.we_clk [13813]));
Q_ASSIGN U18962 ( .B(clk), .A(\g.we_clk [13812]));
Q_ASSIGN U18963 ( .B(clk), .A(\g.we_clk [13811]));
Q_ASSIGN U18964 ( .B(clk), .A(\g.we_clk [13810]));
Q_ASSIGN U18965 ( .B(clk), .A(\g.we_clk [13809]));
Q_ASSIGN U18966 ( .B(clk), .A(\g.we_clk [13808]));
Q_ASSIGN U18967 ( .B(clk), .A(\g.we_clk [13807]));
Q_ASSIGN U18968 ( .B(clk), .A(\g.we_clk [13806]));
Q_ASSIGN U18969 ( .B(clk), .A(\g.we_clk [13805]));
Q_ASSIGN U18970 ( .B(clk), .A(\g.we_clk [13804]));
Q_ASSIGN U18971 ( .B(clk), .A(\g.we_clk [13803]));
Q_ASSIGN U18972 ( .B(clk), .A(\g.we_clk [13802]));
Q_ASSIGN U18973 ( .B(clk), .A(\g.we_clk [13801]));
Q_ASSIGN U18974 ( .B(clk), .A(\g.we_clk [13800]));
Q_ASSIGN U18975 ( .B(clk), .A(\g.we_clk [13799]));
Q_ASSIGN U18976 ( .B(clk), .A(\g.we_clk [13798]));
Q_ASSIGN U18977 ( .B(clk), .A(\g.we_clk [13797]));
Q_ASSIGN U18978 ( .B(clk), .A(\g.we_clk [13796]));
Q_ASSIGN U18979 ( .B(clk), .A(\g.we_clk [13795]));
Q_ASSIGN U18980 ( .B(clk), .A(\g.we_clk [13794]));
Q_ASSIGN U18981 ( .B(clk), .A(\g.we_clk [13793]));
Q_ASSIGN U18982 ( .B(clk), .A(\g.we_clk [13792]));
Q_ASSIGN U18983 ( .B(clk), .A(\g.we_clk [13791]));
Q_ASSIGN U18984 ( .B(clk), .A(\g.we_clk [13790]));
Q_ASSIGN U18985 ( .B(clk), .A(\g.we_clk [13789]));
Q_ASSIGN U18986 ( .B(clk), .A(\g.we_clk [13788]));
Q_ASSIGN U18987 ( .B(clk), .A(\g.we_clk [13787]));
Q_ASSIGN U18988 ( .B(clk), .A(\g.we_clk [13786]));
Q_ASSIGN U18989 ( .B(clk), .A(\g.we_clk [13785]));
Q_ASSIGN U18990 ( .B(clk), .A(\g.we_clk [13784]));
Q_ASSIGN U18991 ( .B(clk), .A(\g.we_clk [13783]));
Q_ASSIGN U18992 ( .B(clk), .A(\g.we_clk [13782]));
Q_ASSIGN U18993 ( .B(clk), .A(\g.we_clk [13781]));
Q_ASSIGN U18994 ( .B(clk), .A(\g.we_clk [13780]));
Q_ASSIGN U18995 ( .B(clk), .A(\g.we_clk [13779]));
Q_ASSIGN U18996 ( .B(clk), .A(\g.we_clk [13778]));
Q_ASSIGN U18997 ( .B(clk), .A(\g.we_clk [13777]));
Q_ASSIGN U18998 ( .B(clk), .A(\g.we_clk [13776]));
Q_ASSIGN U18999 ( .B(clk), .A(\g.we_clk [13775]));
Q_ASSIGN U19000 ( .B(clk), .A(\g.we_clk [13774]));
Q_ASSIGN U19001 ( .B(clk), .A(\g.we_clk [13773]));
Q_ASSIGN U19002 ( .B(clk), .A(\g.we_clk [13772]));
Q_ASSIGN U19003 ( .B(clk), .A(\g.we_clk [13771]));
Q_ASSIGN U19004 ( .B(clk), .A(\g.we_clk [13770]));
Q_ASSIGN U19005 ( .B(clk), .A(\g.we_clk [13769]));
Q_ASSIGN U19006 ( .B(clk), .A(\g.we_clk [13768]));
Q_ASSIGN U19007 ( .B(clk), .A(\g.we_clk [13767]));
Q_ASSIGN U19008 ( .B(clk), .A(\g.we_clk [13766]));
Q_ASSIGN U19009 ( .B(clk), .A(\g.we_clk [13765]));
Q_ASSIGN U19010 ( .B(clk), .A(\g.we_clk [13764]));
Q_ASSIGN U19011 ( .B(clk), .A(\g.we_clk [13763]));
Q_ASSIGN U19012 ( .B(clk), .A(\g.we_clk [13762]));
Q_ASSIGN U19013 ( .B(clk), .A(\g.we_clk [13761]));
Q_ASSIGN U19014 ( .B(clk), .A(\g.we_clk [13760]));
Q_ASSIGN U19015 ( .B(clk), .A(\g.we_clk [13759]));
Q_ASSIGN U19016 ( .B(clk), .A(\g.we_clk [13758]));
Q_ASSIGN U19017 ( .B(clk), .A(\g.we_clk [13757]));
Q_ASSIGN U19018 ( .B(clk), .A(\g.we_clk [13756]));
Q_ASSIGN U19019 ( .B(clk), .A(\g.we_clk [13755]));
Q_ASSIGN U19020 ( .B(clk), .A(\g.we_clk [13754]));
Q_ASSIGN U19021 ( .B(clk), .A(\g.we_clk [13753]));
Q_ASSIGN U19022 ( .B(clk), .A(\g.we_clk [13752]));
Q_ASSIGN U19023 ( .B(clk), .A(\g.we_clk [13751]));
Q_ASSIGN U19024 ( .B(clk), .A(\g.we_clk [13750]));
Q_ASSIGN U19025 ( .B(clk), .A(\g.we_clk [13749]));
Q_ASSIGN U19026 ( .B(clk), .A(\g.we_clk [13748]));
Q_ASSIGN U19027 ( .B(clk), .A(\g.we_clk [13747]));
Q_ASSIGN U19028 ( .B(clk), .A(\g.we_clk [13746]));
Q_ASSIGN U19029 ( .B(clk), .A(\g.we_clk [13745]));
Q_ASSIGN U19030 ( .B(clk), .A(\g.we_clk [13744]));
Q_ASSIGN U19031 ( .B(clk), .A(\g.we_clk [13743]));
Q_ASSIGN U19032 ( .B(clk), .A(\g.we_clk [13742]));
Q_ASSIGN U19033 ( .B(clk), .A(\g.we_clk [13741]));
Q_ASSIGN U19034 ( .B(clk), .A(\g.we_clk [13740]));
Q_ASSIGN U19035 ( .B(clk), .A(\g.we_clk [13739]));
Q_ASSIGN U19036 ( .B(clk), .A(\g.we_clk [13738]));
Q_ASSIGN U19037 ( .B(clk), .A(\g.we_clk [13737]));
Q_ASSIGN U19038 ( .B(clk), .A(\g.we_clk [13736]));
Q_ASSIGN U19039 ( .B(clk), .A(\g.we_clk [13735]));
Q_ASSIGN U19040 ( .B(clk), .A(\g.we_clk [13734]));
Q_ASSIGN U19041 ( .B(clk), .A(\g.we_clk [13733]));
Q_ASSIGN U19042 ( .B(clk), .A(\g.we_clk [13732]));
Q_ASSIGN U19043 ( .B(clk), .A(\g.we_clk [13731]));
Q_ASSIGN U19044 ( .B(clk), .A(\g.we_clk [13730]));
Q_ASSIGN U19045 ( .B(clk), .A(\g.we_clk [13729]));
Q_ASSIGN U19046 ( .B(clk), .A(\g.we_clk [13728]));
Q_ASSIGN U19047 ( .B(clk), .A(\g.we_clk [13727]));
Q_ASSIGN U19048 ( .B(clk), .A(\g.we_clk [13726]));
Q_ASSIGN U19049 ( .B(clk), .A(\g.we_clk [13725]));
Q_ASSIGN U19050 ( .B(clk), .A(\g.we_clk [13724]));
Q_ASSIGN U19051 ( .B(clk), .A(\g.we_clk [13723]));
Q_ASSIGN U19052 ( .B(clk), .A(\g.we_clk [13722]));
Q_ASSIGN U19053 ( .B(clk), .A(\g.we_clk [13721]));
Q_ASSIGN U19054 ( .B(clk), .A(\g.we_clk [13720]));
Q_ASSIGN U19055 ( .B(clk), .A(\g.we_clk [13719]));
Q_ASSIGN U19056 ( .B(clk), .A(\g.we_clk [13718]));
Q_ASSIGN U19057 ( .B(clk), .A(\g.we_clk [13717]));
Q_ASSIGN U19058 ( .B(clk), .A(\g.we_clk [13716]));
Q_ASSIGN U19059 ( .B(clk), .A(\g.we_clk [13715]));
Q_ASSIGN U19060 ( .B(clk), .A(\g.we_clk [13714]));
Q_ASSIGN U19061 ( .B(clk), .A(\g.we_clk [13713]));
Q_ASSIGN U19062 ( .B(clk), .A(\g.we_clk [13712]));
Q_ASSIGN U19063 ( .B(clk), .A(\g.we_clk [13711]));
Q_ASSIGN U19064 ( .B(clk), .A(\g.we_clk [13710]));
Q_ASSIGN U19065 ( .B(clk), .A(\g.we_clk [13709]));
Q_ASSIGN U19066 ( .B(clk), .A(\g.we_clk [13708]));
Q_ASSIGN U19067 ( .B(clk), .A(\g.we_clk [13707]));
Q_ASSIGN U19068 ( .B(clk), .A(\g.we_clk [13706]));
Q_ASSIGN U19069 ( .B(clk), .A(\g.we_clk [13705]));
Q_ASSIGN U19070 ( .B(clk), .A(\g.we_clk [13704]));
Q_ASSIGN U19071 ( .B(clk), .A(\g.we_clk [13703]));
Q_ASSIGN U19072 ( .B(clk), .A(\g.we_clk [13702]));
Q_ASSIGN U19073 ( .B(clk), .A(\g.we_clk [13701]));
Q_ASSIGN U19074 ( .B(clk), .A(\g.we_clk [13700]));
Q_ASSIGN U19075 ( .B(clk), .A(\g.we_clk [13699]));
Q_ASSIGN U19076 ( .B(clk), .A(\g.we_clk [13698]));
Q_ASSIGN U19077 ( .B(clk), .A(\g.we_clk [13697]));
Q_ASSIGN U19078 ( .B(clk), .A(\g.we_clk [13696]));
Q_ASSIGN U19079 ( .B(clk), .A(\g.we_clk [13695]));
Q_ASSIGN U19080 ( .B(clk), .A(\g.we_clk [13694]));
Q_ASSIGN U19081 ( .B(clk), .A(\g.we_clk [13693]));
Q_ASSIGN U19082 ( .B(clk), .A(\g.we_clk [13692]));
Q_ASSIGN U19083 ( .B(clk), .A(\g.we_clk [13691]));
Q_ASSIGN U19084 ( .B(clk), .A(\g.we_clk [13690]));
Q_ASSIGN U19085 ( .B(clk), .A(\g.we_clk [13689]));
Q_ASSIGN U19086 ( .B(clk), .A(\g.we_clk [13688]));
Q_ASSIGN U19087 ( .B(clk), .A(\g.we_clk [13687]));
Q_ASSIGN U19088 ( .B(clk), .A(\g.we_clk [13686]));
Q_ASSIGN U19089 ( .B(clk), .A(\g.we_clk [13685]));
Q_ASSIGN U19090 ( .B(clk), .A(\g.we_clk [13684]));
Q_ASSIGN U19091 ( .B(clk), .A(\g.we_clk [13683]));
Q_ASSIGN U19092 ( .B(clk), .A(\g.we_clk [13682]));
Q_ASSIGN U19093 ( .B(clk), .A(\g.we_clk [13681]));
Q_ASSIGN U19094 ( .B(clk), .A(\g.we_clk [13680]));
Q_ASSIGN U19095 ( .B(clk), .A(\g.we_clk [13679]));
Q_ASSIGN U19096 ( .B(clk), .A(\g.we_clk [13678]));
Q_ASSIGN U19097 ( .B(clk), .A(\g.we_clk [13677]));
Q_ASSIGN U19098 ( .B(clk), .A(\g.we_clk [13676]));
Q_ASSIGN U19099 ( .B(clk), .A(\g.we_clk [13675]));
Q_ASSIGN U19100 ( .B(clk), .A(\g.we_clk [13674]));
Q_ASSIGN U19101 ( .B(clk), .A(\g.we_clk [13673]));
Q_ASSIGN U19102 ( .B(clk), .A(\g.we_clk [13672]));
Q_ASSIGN U19103 ( .B(clk), .A(\g.we_clk [13671]));
Q_ASSIGN U19104 ( .B(clk), .A(\g.we_clk [13670]));
Q_ASSIGN U19105 ( .B(clk), .A(\g.we_clk [13669]));
Q_ASSIGN U19106 ( .B(clk), .A(\g.we_clk [13668]));
Q_ASSIGN U19107 ( .B(clk), .A(\g.we_clk [13667]));
Q_ASSIGN U19108 ( .B(clk), .A(\g.we_clk [13666]));
Q_ASSIGN U19109 ( .B(clk), .A(\g.we_clk [13665]));
Q_ASSIGN U19110 ( .B(clk), .A(\g.we_clk [13664]));
Q_ASSIGN U19111 ( .B(clk), .A(\g.we_clk [13663]));
Q_ASSIGN U19112 ( .B(clk), .A(\g.we_clk [13662]));
Q_ASSIGN U19113 ( .B(clk), .A(\g.we_clk [13661]));
Q_ASSIGN U19114 ( .B(clk), .A(\g.we_clk [13660]));
Q_ASSIGN U19115 ( .B(clk), .A(\g.we_clk [13659]));
Q_ASSIGN U19116 ( .B(clk), .A(\g.we_clk [13658]));
Q_ASSIGN U19117 ( .B(clk), .A(\g.we_clk [13657]));
Q_ASSIGN U19118 ( .B(clk), .A(\g.we_clk [13656]));
Q_ASSIGN U19119 ( .B(clk), .A(\g.we_clk [13655]));
Q_ASSIGN U19120 ( .B(clk), .A(\g.we_clk [13654]));
Q_ASSIGN U19121 ( .B(clk), .A(\g.we_clk [13653]));
Q_ASSIGN U19122 ( .B(clk), .A(\g.we_clk [13652]));
Q_ASSIGN U19123 ( .B(clk), .A(\g.we_clk [13651]));
Q_ASSIGN U19124 ( .B(clk), .A(\g.we_clk [13650]));
Q_ASSIGN U19125 ( .B(clk), .A(\g.we_clk [13649]));
Q_ASSIGN U19126 ( .B(clk), .A(\g.we_clk [13648]));
Q_ASSIGN U19127 ( .B(clk), .A(\g.we_clk [13647]));
Q_ASSIGN U19128 ( .B(clk), .A(\g.we_clk [13646]));
Q_ASSIGN U19129 ( .B(clk), .A(\g.we_clk [13645]));
Q_ASSIGN U19130 ( .B(clk), .A(\g.we_clk [13644]));
Q_ASSIGN U19131 ( .B(clk), .A(\g.we_clk [13643]));
Q_ASSIGN U19132 ( .B(clk), .A(\g.we_clk [13642]));
Q_ASSIGN U19133 ( .B(clk), .A(\g.we_clk [13641]));
Q_ASSIGN U19134 ( .B(clk), .A(\g.we_clk [13640]));
Q_ASSIGN U19135 ( .B(clk), .A(\g.we_clk [13639]));
Q_ASSIGN U19136 ( .B(clk), .A(\g.we_clk [13638]));
Q_ASSIGN U19137 ( .B(clk), .A(\g.we_clk [13637]));
Q_ASSIGN U19138 ( .B(clk), .A(\g.we_clk [13636]));
Q_ASSIGN U19139 ( .B(clk), .A(\g.we_clk [13635]));
Q_ASSIGN U19140 ( .B(clk), .A(\g.we_clk [13634]));
Q_ASSIGN U19141 ( .B(clk), .A(\g.we_clk [13633]));
Q_ASSIGN U19142 ( .B(clk), .A(\g.we_clk [13632]));
Q_ASSIGN U19143 ( .B(clk), .A(\g.we_clk [13631]));
Q_ASSIGN U19144 ( .B(clk), .A(\g.we_clk [13630]));
Q_ASSIGN U19145 ( .B(clk), .A(\g.we_clk [13629]));
Q_ASSIGN U19146 ( .B(clk), .A(\g.we_clk [13628]));
Q_ASSIGN U19147 ( .B(clk), .A(\g.we_clk [13627]));
Q_ASSIGN U19148 ( .B(clk), .A(\g.we_clk [13626]));
Q_ASSIGN U19149 ( .B(clk), .A(\g.we_clk [13625]));
Q_ASSIGN U19150 ( .B(clk), .A(\g.we_clk [13624]));
Q_ASSIGN U19151 ( .B(clk), .A(\g.we_clk [13623]));
Q_ASSIGN U19152 ( .B(clk), .A(\g.we_clk [13622]));
Q_ASSIGN U19153 ( .B(clk), .A(\g.we_clk [13621]));
Q_ASSIGN U19154 ( .B(clk), .A(\g.we_clk [13620]));
Q_ASSIGN U19155 ( .B(clk), .A(\g.we_clk [13619]));
Q_ASSIGN U19156 ( .B(clk), .A(\g.we_clk [13618]));
Q_ASSIGN U19157 ( .B(clk), .A(\g.we_clk [13617]));
Q_ASSIGN U19158 ( .B(clk), .A(\g.we_clk [13616]));
Q_ASSIGN U19159 ( .B(clk), .A(\g.we_clk [13615]));
Q_ASSIGN U19160 ( .B(clk), .A(\g.we_clk [13614]));
Q_ASSIGN U19161 ( .B(clk), .A(\g.we_clk [13613]));
Q_ASSIGN U19162 ( .B(clk), .A(\g.we_clk [13612]));
Q_ASSIGN U19163 ( .B(clk), .A(\g.we_clk [13611]));
Q_ASSIGN U19164 ( .B(clk), .A(\g.we_clk [13610]));
Q_ASSIGN U19165 ( .B(clk), .A(\g.we_clk [13609]));
Q_ASSIGN U19166 ( .B(clk), .A(\g.we_clk [13608]));
Q_ASSIGN U19167 ( .B(clk), .A(\g.we_clk [13607]));
Q_ASSIGN U19168 ( .B(clk), .A(\g.we_clk [13606]));
Q_ASSIGN U19169 ( .B(clk), .A(\g.we_clk [13605]));
Q_ASSIGN U19170 ( .B(clk), .A(\g.we_clk [13604]));
Q_ASSIGN U19171 ( .B(clk), .A(\g.we_clk [13603]));
Q_ASSIGN U19172 ( .B(clk), .A(\g.we_clk [13602]));
Q_ASSIGN U19173 ( .B(clk), .A(\g.we_clk [13601]));
Q_ASSIGN U19174 ( .B(clk), .A(\g.we_clk [13600]));
Q_ASSIGN U19175 ( .B(clk), .A(\g.we_clk [13599]));
Q_ASSIGN U19176 ( .B(clk), .A(\g.we_clk [13598]));
Q_ASSIGN U19177 ( .B(clk), .A(\g.we_clk [13597]));
Q_ASSIGN U19178 ( .B(clk), .A(\g.we_clk [13596]));
Q_ASSIGN U19179 ( .B(clk), .A(\g.we_clk [13595]));
Q_ASSIGN U19180 ( .B(clk), .A(\g.we_clk [13594]));
Q_ASSIGN U19181 ( .B(clk), .A(\g.we_clk [13593]));
Q_ASSIGN U19182 ( .B(clk), .A(\g.we_clk [13592]));
Q_ASSIGN U19183 ( .B(clk), .A(\g.we_clk [13591]));
Q_ASSIGN U19184 ( .B(clk), .A(\g.we_clk [13590]));
Q_ASSIGN U19185 ( .B(clk), .A(\g.we_clk [13589]));
Q_ASSIGN U19186 ( .B(clk), .A(\g.we_clk [13588]));
Q_ASSIGN U19187 ( .B(clk), .A(\g.we_clk [13587]));
Q_ASSIGN U19188 ( .B(clk), .A(\g.we_clk [13586]));
Q_ASSIGN U19189 ( .B(clk), .A(\g.we_clk [13585]));
Q_ASSIGN U19190 ( .B(clk), .A(\g.we_clk [13584]));
Q_ASSIGN U19191 ( .B(clk), .A(\g.we_clk [13583]));
Q_ASSIGN U19192 ( .B(clk), .A(\g.we_clk [13582]));
Q_ASSIGN U19193 ( .B(clk), .A(\g.we_clk [13581]));
Q_ASSIGN U19194 ( .B(clk), .A(\g.we_clk [13580]));
Q_ASSIGN U19195 ( .B(clk), .A(\g.we_clk [13579]));
Q_ASSIGN U19196 ( .B(clk), .A(\g.we_clk [13578]));
Q_ASSIGN U19197 ( .B(clk), .A(\g.we_clk [13577]));
Q_ASSIGN U19198 ( .B(clk), .A(\g.we_clk [13576]));
Q_ASSIGN U19199 ( .B(clk), .A(\g.we_clk [13575]));
Q_ASSIGN U19200 ( .B(clk), .A(\g.we_clk [13574]));
Q_ASSIGN U19201 ( .B(clk), .A(\g.we_clk [13573]));
Q_ASSIGN U19202 ( .B(clk), .A(\g.we_clk [13572]));
Q_ASSIGN U19203 ( .B(clk), .A(\g.we_clk [13571]));
Q_ASSIGN U19204 ( .B(clk), .A(\g.we_clk [13570]));
Q_ASSIGN U19205 ( .B(clk), .A(\g.we_clk [13569]));
Q_ASSIGN U19206 ( .B(clk), .A(\g.we_clk [13568]));
Q_ASSIGN U19207 ( .B(clk), .A(\g.we_clk [13567]));
Q_ASSIGN U19208 ( .B(clk), .A(\g.we_clk [13566]));
Q_ASSIGN U19209 ( .B(clk), .A(\g.we_clk [13565]));
Q_ASSIGN U19210 ( .B(clk), .A(\g.we_clk [13564]));
Q_ASSIGN U19211 ( .B(clk), .A(\g.we_clk [13563]));
Q_ASSIGN U19212 ( .B(clk), .A(\g.we_clk [13562]));
Q_ASSIGN U19213 ( .B(clk), .A(\g.we_clk [13561]));
Q_ASSIGN U19214 ( .B(clk), .A(\g.we_clk [13560]));
Q_ASSIGN U19215 ( .B(clk), .A(\g.we_clk [13559]));
Q_ASSIGN U19216 ( .B(clk), .A(\g.we_clk [13558]));
Q_ASSIGN U19217 ( .B(clk), .A(\g.we_clk [13557]));
Q_ASSIGN U19218 ( .B(clk), .A(\g.we_clk [13556]));
Q_ASSIGN U19219 ( .B(clk), .A(\g.we_clk [13555]));
Q_ASSIGN U19220 ( .B(clk), .A(\g.we_clk [13554]));
Q_ASSIGN U19221 ( .B(clk), .A(\g.we_clk [13553]));
Q_ASSIGN U19222 ( .B(clk), .A(\g.we_clk [13552]));
Q_ASSIGN U19223 ( .B(clk), .A(\g.we_clk [13551]));
Q_ASSIGN U19224 ( .B(clk), .A(\g.we_clk [13550]));
Q_ASSIGN U19225 ( .B(clk), .A(\g.we_clk [13549]));
Q_ASSIGN U19226 ( .B(clk), .A(\g.we_clk [13548]));
Q_ASSIGN U19227 ( .B(clk), .A(\g.we_clk [13547]));
Q_ASSIGN U19228 ( .B(clk), .A(\g.we_clk [13546]));
Q_ASSIGN U19229 ( .B(clk), .A(\g.we_clk [13545]));
Q_ASSIGN U19230 ( .B(clk), .A(\g.we_clk [13544]));
Q_ASSIGN U19231 ( .B(clk), .A(\g.we_clk [13543]));
Q_ASSIGN U19232 ( .B(clk), .A(\g.we_clk [13542]));
Q_ASSIGN U19233 ( .B(clk), .A(\g.we_clk [13541]));
Q_ASSIGN U19234 ( .B(clk), .A(\g.we_clk [13540]));
Q_ASSIGN U19235 ( .B(clk), .A(\g.we_clk [13539]));
Q_ASSIGN U19236 ( .B(clk), .A(\g.we_clk [13538]));
Q_ASSIGN U19237 ( .B(clk), .A(\g.we_clk [13537]));
Q_ASSIGN U19238 ( .B(clk), .A(\g.we_clk [13536]));
Q_ASSIGN U19239 ( .B(clk), .A(\g.we_clk [13535]));
Q_ASSIGN U19240 ( .B(clk), .A(\g.we_clk [13534]));
Q_ASSIGN U19241 ( .B(clk), .A(\g.we_clk [13533]));
Q_ASSIGN U19242 ( .B(clk), .A(\g.we_clk [13532]));
Q_ASSIGN U19243 ( .B(clk), .A(\g.we_clk [13531]));
Q_ASSIGN U19244 ( .B(clk), .A(\g.we_clk [13530]));
Q_ASSIGN U19245 ( .B(clk), .A(\g.we_clk [13529]));
Q_ASSIGN U19246 ( .B(clk), .A(\g.we_clk [13528]));
Q_ASSIGN U19247 ( .B(clk), .A(\g.we_clk [13527]));
Q_ASSIGN U19248 ( .B(clk), .A(\g.we_clk [13526]));
Q_ASSIGN U19249 ( .B(clk), .A(\g.we_clk [13525]));
Q_ASSIGN U19250 ( .B(clk), .A(\g.we_clk [13524]));
Q_ASSIGN U19251 ( .B(clk), .A(\g.we_clk [13523]));
Q_ASSIGN U19252 ( .B(clk), .A(\g.we_clk [13522]));
Q_ASSIGN U19253 ( .B(clk), .A(\g.we_clk [13521]));
Q_ASSIGN U19254 ( .B(clk), .A(\g.we_clk [13520]));
Q_ASSIGN U19255 ( .B(clk), .A(\g.we_clk [13519]));
Q_ASSIGN U19256 ( .B(clk), .A(\g.we_clk [13518]));
Q_ASSIGN U19257 ( .B(clk), .A(\g.we_clk [13517]));
Q_ASSIGN U19258 ( .B(clk), .A(\g.we_clk [13516]));
Q_ASSIGN U19259 ( .B(clk), .A(\g.we_clk [13515]));
Q_ASSIGN U19260 ( .B(clk), .A(\g.we_clk [13514]));
Q_ASSIGN U19261 ( .B(clk), .A(\g.we_clk [13513]));
Q_ASSIGN U19262 ( .B(clk), .A(\g.we_clk [13512]));
Q_ASSIGN U19263 ( .B(clk), .A(\g.we_clk [13511]));
Q_ASSIGN U19264 ( .B(clk), .A(\g.we_clk [13510]));
Q_ASSIGN U19265 ( .B(clk), .A(\g.we_clk [13509]));
Q_ASSIGN U19266 ( .B(clk), .A(\g.we_clk [13508]));
Q_ASSIGN U19267 ( .B(clk), .A(\g.we_clk [13507]));
Q_ASSIGN U19268 ( .B(clk), .A(\g.we_clk [13506]));
Q_ASSIGN U19269 ( .B(clk), .A(\g.we_clk [13505]));
Q_ASSIGN U19270 ( .B(clk), .A(\g.we_clk [13504]));
Q_ASSIGN U19271 ( .B(clk), .A(\g.we_clk [13503]));
Q_ASSIGN U19272 ( .B(clk), .A(\g.we_clk [13502]));
Q_ASSIGN U19273 ( .B(clk), .A(\g.we_clk [13501]));
Q_ASSIGN U19274 ( .B(clk), .A(\g.we_clk [13500]));
Q_ASSIGN U19275 ( .B(clk), .A(\g.we_clk [13499]));
Q_ASSIGN U19276 ( .B(clk), .A(\g.we_clk [13498]));
Q_ASSIGN U19277 ( .B(clk), .A(\g.we_clk [13497]));
Q_ASSIGN U19278 ( .B(clk), .A(\g.we_clk [13496]));
Q_ASSIGN U19279 ( .B(clk), .A(\g.we_clk [13495]));
Q_ASSIGN U19280 ( .B(clk), .A(\g.we_clk [13494]));
Q_ASSIGN U19281 ( .B(clk), .A(\g.we_clk [13493]));
Q_ASSIGN U19282 ( .B(clk), .A(\g.we_clk [13492]));
Q_ASSIGN U19283 ( .B(clk), .A(\g.we_clk [13491]));
Q_ASSIGN U19284 ( .B(clk), .A(\g.we_clk [13490]));
Q_ASSIGN U19285 ( .B(clk), .A(\g.we_clk [13489]));
Q_ASSIGN U19286 ( .B(clk), .A(\g.we_clk [13488]));
Q_ASSIGN U19287 ( .B(clk), .A(\g.we_clk [13487]));
Q_ASSIGN U19288 ( .B(clk), .A(\g.we_clk [13486]));
Q_ASSIGN U19289 ( .B(clk), .A(\g.we_clk [13485]));
Q_ASSIGN U19290 ( .B(clk), .A(\g.we_clk [13484]));
Q_ASSIGN U19291 ( .B(clk), .A(\g.we_clk [13483]));
Q_ASSIGN U19292 ( .B(clk), .A(\g.we_clk [13482]));
Q_ASSIGN U19293 ( .B(clk), .A(\g.we_clk [13481]));
Q_ASSIGN U19294 ( .B(clk), .A(\g.we_clk [13480]));
Q_ASSIGN U19295 ( .B(clk), .A(\g.we_clk [13479]));
Q_ASSIGN U19296 ( .B(clk), .A(\g.we_clk [13478]));
Q_ASSIGN U19297 ( .B(clk), .A(\g.we_clk [13477]));
Q_ASSIGN U19298 ( .B(clk), .A(\g.we_clk [13476]));
Q_ASSIGN U19299 ( .B(clk), .A(\g.we_clk [13475]));
Q_ASSIGN U19300 ( .B(clk), .A(\g.we_clk [13474]));
Q_ASSIGN U19301 ( .B(clk), .A(\g.we_clk [13473]));
Q_ASSIGN U19302 ( .B(clk), .A(\g.we_clk [13472]));
Q_ASSIGN U19303 ( .B(clk), .A(\g.we_clk [13471]));
Q_ASSIGN U19304 ( .B(clk), .A(\g.we_clk [13470]));
Q_ASSIGN U19305 ( .B(clk), .A(\g.we_clk [13469]));
Q_ASSIGN U19306 ( .B(clk), .A(\g.we_clk [13468]));
Q_ASSIGN U19307 ( .B(clk), .A(\g.we_clk [13467]));
Q_ASSIGN U19308 ( .B(clk), .A(\g.we_clk [13466]));
Q_ASSIGN U19309 ( .B(clk), .A(\g.we_clk [13465]));
Q_ASSIGN U19310 ( .B(clk), .A(\g.we_clk [13464]));
Q_ASSIGN U19311 ( .B(clk), .A(\g.we_clk [13463]));
Q_ASSIGN U19312 ( .B(clk), .A(\g.we_clk [13462]));
Q_ASSIGN U19313 ( .B(clk), .A(\g.we_clk [13461]));
Q_ASSIGN U19314 ( .B(clk), .A(\g.we_clk [13460]));
Q_ASSIGN U19315 ( .B(clk), .A(\g.we_clk [13459]));
Q_ASSIGN U19316 ( .B(clk), .A(\g.we_clk [13458]));
Q_ASSIGN U19317 ( .B(clk), .A(\g.we_clk [13457]));
Q_ASSIGN U19318 ( .B(clk), .A(\g.we_clk [13456]));
Q_ASSIGN U19319 ( .B(clk), .A(\g.we_clk [13455]));
Q_ASSIGN U19320 ( .B(clk), .A(\g.we_clk [13454]));
Q_ASSIGN U19321 ( .B(clk), .A(\g.we_clk [13453]));
Q_ASSIGN U19322 ( .B(clk), .A(\g.we_clk [13452]));
Q_ASSIGN U19323 ( .B(clk), .A(\g.we_clk [13451]));
Q_ASSIGN U19324 ( .B(clk), .A(\g.we_clk [13450]));
Q_ASSIGN U19325 ( .B(clk), .A(\g.we_clk [13449]));
Q_ASSIGN U19326 ( .B(clk), .A(\g.we_clk [13448]));
Q_ASSIGN U19327 ( .B(clk), .A(\g.we_clk [13447]));
Q_ASSIGN U19328 ( .B(clk), .A(\g.we_clk [13446]));
Q_ASSIGN U19329 ( .B(clk), .A(\g.we_clk [13445]));
Q_ASSIGN U19330 ( .B(clk), .A(\g.we_clk [13444]));
Q_ASSIGN U19331 ( .B(clk), .A(\g.we_clk [13443]));
Q_ASSIGN U19332 ( .B(clk), .A(\g.we_clk [13442]));
Q_ASSIGN U19333 ( .B(clk), .A(\g.we_clk [13441]));
Q_ASSIGN U19334 ( .B(clk), .A(\g.we_clk [13440]));
Q_ASSIGN U19335 ( .B(clk), .A(\g.we_clk [13439]));
Q_ASSIGN U19336 ( .B(clk), .A(\g.we_clk [13438]));
Q_ASSIGN U19337 ( .B(clk), .A(\g.we_clk [13437]));
Q_ASSIGN U19338 ( .B(clk), .A(\g.we_clk [13436]));
Q_ASSIGN U19339 ( .B(clk), .A(\g.we_clk [13435]));
Q_ASSIGN U19340 ( .B(clk), .A(\g.we_clk [13434]));
Q_ASSIGN U19341 ( .B(clk), .A(\g.we_clk [13433]));
Q_ASSIGN U19342 ( .B(clk), .A(\g.we_clk [13432]));
Q_ASSIGN U19343 ( .B(clk), .A(\g.we_clk [13431]));
Q_ASSIGN U19344 ( .B(clk), .A(\g.we_clk [13430]));
Q_ASSIGN U19345 ( .B(clk), .A(\g.we_clk [13429]));
Q_ASSIGN U19346 ( .B(clk), .A(\g.we_clk [13428]));
Q_ASSIGN U19347 ( .B(clk), .A(\g.we_clk [13427]));
Q_ASSIGN U19348 ( .B(clk), .A(\g.we_clk [13426]));
Q_ASSIGN U19349 ( .B(clk), .A(\g.we_clk [13425]));
Q_ASSIGN U19350 ( .B(clk), .A(\g.we_clk [13424]));
Q_ASSIGN U19351 ( .B(clk), .A(\g.we_clk [13423]));
Q_ASSIGN U19352 ( .B(clk), .A(\g.we_clk [13422]));
Q_ASSIGN U19353 ( .B(clk), .A(\g.we_clk [13421]));
Q_ASSIGN U19354 ( .B(clk), .A(\g.we_clk [13420]));
Q_ASSIGN U19355 ( .B(clk), .A(\g.we_clk [13419]));
Q_ASSIGN U19356 ( .B(clk), .A(\g.we_clk [13418]));
Q_ASSIGN U19357 ( .B(clk), .A(\g.we_clk [13417]));
Q_ASSIGN U19358 ( .B(clk), .A(\g.we_clk [13416]));
Q_ASSIGN U19359 ( .B(clk), .A(\g.we_clk [13415]));
Q_ASSIGN U19360 ( .B(clk), .A(\g.we_clk [13414]));
Q_ASSIGN U19361 ( .B(clk), .A(\g.we_clk [13413]));
Q_ASSIGN U19362 ( .B(clk), .A(\g.we_clk [13412]));
Q_ASSIGN U19363 ( .B(clk), .A(\g.we_clk [13411]));
Q_ASSIGN U19364 ( .B(clk), .A(\g.we_clk [13410]));
Q_ASSIGN U19365 ( .B(clk), .A(\g.we_clk [13409]));
Q_ASSIGN U19366 ( .B(clk), .A(\g.we_clk [13408]));
Q_ASSIGN U19367 ( .B(clk), .A(\g.we_clk [13407]));
Q_ASSIGN U19368 ( .B(clk), .A(\g.we_clk [13406]));
Q_ASSIGN U19369 ( .B(clk), .A(\g.we_clk [13405]));
Q_ASSIGN U19370 ( .B(clk), .A(\g.we_clk [13404]));
Q_ASSIGN U19371 ( .B(clk), .A(\g.we_clk [13403]));
Q_ASSIGN U19372 ( .B(clk), .A(\g.we_clk [13402]));
Q_ASSIGN U19373 ( .B(clk), .A(\g.we_clk [13401]));
Q_ASSIGN U19374 ( .B(clk), .A(\g.we_clk [13400]));
Q_ASSIGN U19375 ( .B(clk), .A(\g.we_clk [13399]));
Q_ASSIGN U19376 ( .B(clk), .A(\g.we_clk [13398]));
Q_ASSIGN U19377 ( .B(clk), .A(\g.we_clk [13397]));
Q_ASSIGN U19378 ( .B(clk), .A(\g.we_clk [13396]));
Q_ASSIGN U19379 ( .B(clk), .A(\g.we_clk [13395]));
Q_ASSIGN U19380 ( .B(clk), .A(\g.we_clk [13394]));
Q_ASSIGN U19381 ( .B(clk), .A(\g.we_clk [13393]));
Q_ASSIGN U19382 ( .B(clk), .A(\g.we_clk [13392]));
Q_ASSIGN U19383 ( .B(clk), .A(\g.we_clk [13391]));
Q_ASSIGN U19384 ( .B(clk), .A(\g.we_clk [13390]));
Q_ASSIGN U19385 ( .B(clk), .A(\g.we_clk [13389]));
Q_ASSIGN U19386 ( .B(clk), .A(\g.we_clk [13388]));
Q_ASSIGN U19387 ( .B(clk), .A(\g.we_clk [13387]));
Q_ASSIGN U19388 ( .B(clk), .A(\g.we_clk [13386]));
Q_ASSIGN U19389 ( .B(clk), .A(\g.we_clk [13385]));
Q_ASSIGN U19390 ( .B(clk), .A(\g.we_clk [13384]));
Q_ASSIGN U19391 ( .B(clk), .A(\g.we_clk [13383]));
Q_ASSIGN U19392 ( .B(clk), .A(\g.we_clk [13382]));
Q_ASSIGN U19393 ( .B(clk), .A(\g.we_clk [13381]));
Q_ASSIGN U19394 ( .B(clk), .A(\g.we_clk [13380]));
Q_ASSIGN U19395 ( .B(clk), .A(\g.we_clk [13379]));
Q_ASSIGN U19396 ( .B(clk), .A(\g.we_clk [13378]));
Q_ASSIGN U19397 ( .B(clk), .A(\g.we_clk [13377]));
Q_ASSIGN U19398 ( .B(clk), .A(\g.we_clk [13376]));
Q_ASSIGN U19399 ( .B(clk), .A(\g.we_clk [13375]));
Q_ASSIGN U19400 ( .B(clk), .A(\g.we_clk [13374]));
Q_ASSIGN U19401 ( .B(clk), .A(\g.we_clk [13373]));
Q_ASSIGN U19402 ( .B(clk), .A(\g.we_clk [13372]));
Q_ASSIGN U19403 ( .B(clk), .A(\g.we_clk [13371]));
Q_ASSIGN U19404 ( .B(clk), .A(\g.we_clk [13370]));
Q_ASSIGN U19405 ( .B(clk), .A(\g.we_clk [13369]));
Q_ASSIGN U19406 ( .B(clk), .A(\g.we_clk [13368]));
Q_ASSIGN U19407 ( .B(clk), .A(\g.we_clk [13367]));
Q_ASSIGN U19408 ( .B(clk), .A(\g.we_clk [13366]));
Q_ASSIGN U19409 ( .B(clk), .A(\g.we_clk [13365]));
Q_ASSIGN U19410 ( .B(clk), .A(\g.we_clk [13364]));
Q_ASSIGN U19411 ( .B(clk), .A(\g.we_clk [13363]));
Q_ASSIGN U19412 ( .B(clk), .A(\g.we_clk [13362]));
Q_ASSIGN U19413 ( .B(clk), .A(\g.we_clk [13361]));
Q_ASSIGN U19414 ( .B(clk), .A(\g.we_clk [13360]));
Q_ASSIGN U19415 ( .B(clk), .A(\g.we_clk [13359]));
Q_ASSIGN U19416 ( .B(clk), .A(\g.we_clk [13358]));
Q_ASSIGN U19417 ( .B(clk), .A(\g.we_clk [13357]));
Q_ASSIGN U19418 ( .B(clk), .A(\g.we_clk [13356]));
Q_ASSIGN U19419 ( .B(clk), .A(\g.we_clk [13355]));
Q_ASSIGN U19420 ( .B(clk), .A(\g.we_clk [13354]));
Q_ASSIGN U19421 ( .B(clk), .A(\g.we_clk [13353]));
Q_ASSIGN U19422 ( .B(clk), .A(\g.we_clk [13352]));
Q_ASSIGN U19423 ( .B(clk), .A(\g.we_clk [13351]));
Q_ASSIGN U19424 ( .B(clk), .A(\g.we_clk [13350]));
Q_ASSIGN U19425 ( .B(clk), .A(\g.we_clk [13349]));
Q_ASSIGN U19426 ( .B(clk), .A(\g.we_clk [13348]));
Q_ASSIGN U19427 ( .B(clk), .A(\g.we_clk [13347]));
Q_ASSIGN U19428 ( .B(clk), .A(\g.we_clk [13346]));
Q_ASSIGN U19429 ( .B(clk), .A(\g.we_clk [13345]));
Q_ASSIGN U19430 ( .B(clk), .A(\g.we_clk [13344]));
Q_ASSIGN U19431 ( .B(clk), .A(\g.we_clk [13343]));
Q_ASSIGN U19432 ( .B(clk), .A(\g.we_clk [13342]));
Q_ASSIGN U19433 ( .B(clk), .A(\g.we_clk [13341]));
Q_ASSIGN U19434 ( .B(clk), .A(\g.we_clk [13340]));
Q_ASSIGN U19435 ( .B(clk), .A(\g.we_clk [13339]));
Q_ASSIGN U19436 ( .B(clk), .A(\g.we_clk [13338]));
Q_ASSIGN U19437 ( .B(clk), .A(\g.we_clk [13337]));
Q_ASSIGN U19438 ( .B(clk), .A(\g.we_clk [13336]));
Q_ASSIGN U19439 ( .B(clk), .A(\g.we_clk [13335]));
Q_ASSIGN U19440 ( .B(clk), .A(\g.we_clk [13334]));
Q_ASSIGN U19441 ( .B(clk), .A(\g.we_clk [13333]));
Q_ASSIGN U19442 ( .B(clk), .A(\g.we_clk [13332]));
Q_ASSIGN U19443 ( .B(clk), .A(\g.we_clk [13331]));
Q_ASSIGN U19444 ( .B(clk), .A(\g.we_clk [13330]));
Q_ASSIGN U19445 ( .B(clk), .A(\g.we_clk [13329]));
Q_ASSIGN U19446 ( .B(clk), .A(\g.we_clk [13328]));
Q_ASSIGN U19447 ( .B(clk), .A(\g.we_clk [13327]));
Q_ASSIGN U19448 ( .B(clk), .A(\g.we_clk [13326]));
Q_ASSIGN U19449 ( .B(clk), .A(\g.we_clk [13325]));
Q_ASSIGN U19450 ( .B(clk), .A(\g.we_clk [13324]));
Q_ASSIGN U19451 ( .B(clk), .A(\g.we_clk [13323]));
Q_ASSIGN U19452 ( .B(clk), .A(\g.we_clk [13322]));
Q_ASSIGN U19453 ( .B(clk), .A(\g.we_clk [13321]));
Q_ASSIGN U19454 ( .B(clk), .A(\g.we_clk [13320]));
Q_ASSIGN U19455 ( .B(clk), .A(\g.we_clk [13319]));
Q_ASSIGN U19456 ( .B(clk), .A(\g.we_clk [13318]));
Q_ASSIGN U19457 ( .B(clk), .A(\g.we_clk [13317]));
Q_ASSIGN U19458 ( .B(clk), .A(\g.we_clk [13316]));
Q_ASSIGN U19459 ( .B(clk), .A(\g.we_clk [13315]));
Q_ASSIGN U19460 ( .B(clk), .A(\g.we_clk [13314]));
Q_ASSIGN U19461 ( .B(clk), .A(\g.we_clk [13313]));
Q_ASSIGN U19462 ( .B(clk), .A(\g.we_clk [13312]));
Q_ASSIGN U19463 ( .B(clk), .A(\g.we_clk [13311]));
Q_ASSIGN U19464 ( .B(clk), .A(\g.we_clk [13310]));
Q_ASSIGN U19465 ( .B(clk), .A(\g.we_clk [13309]));
Q_ASSIGN U19466 ( .B(clk), .A(\g.we_clk [13308]));
Q_ASSIGN U19467 ( .B(clk), .A(\g.we_clk [13307]));
Q_ASSIGN U19468 ( .B(clk), .A(\g.we_clk [13306]));
Q_ASSIGN U19469 ( .B(clk), .A(\g.we_clk [13305]));
Q_ASSIGN U19470 ( .B(clk), .A(\g.we_clk [13304]));
Q_ASSIGN U19471 ( .B(clk), .A(\g.we_clk [13303]));
Q_ASSIGN U19472 ( .B(clk), .A(\g.we_clk [13302]));
Q_ASSIGN U19473 ( .B(clk), .A(\g.we_clk [13301]));
Q_ASSIGN U19474 ( .B(clk), .A(\g.we_clk [13300]));
Q_ASSIGN U19475 ( .B(clk), .A(\g.we_clk [13299]));
Q_ASSIGN U19476 ( .B(clk), .A(\g.we_clk [13298]));
Q_ASSIGN U19477 ( .B(clk), .A(\g.we_clk [13297]));
Q_ASSIGN U19478 ( .B(clk), .A(\g.we_clk [13296]));
Q_ASSIGN U19479 ( .B(clk), .A(\g.we_clk [13295]));
Q_ASSIGN U19480 ( .B(clk), .A(\g.we_clk [13294]));
Q_ASSIGN U19481 ( .B(clk), .A(\g.we_clk [13293]));
Q_ASSIGN U19482 ( .B(clk), .A(\g.we_clk [13292]));
Q_ASSIGN U19483 ( .B(clk), .A(\g.we_clk [13291]));
Q_ASSIGN U19484 ( .B(clk), .A(\g.we_clk [13290]));
Q_ASSIGN U19485 ( .B(clk), .A(\g.we_clk [13289]));
Q_ASSIGN U19486 ( .B(clk), .A(\g.we_clk [13288]));
Q_ASSIGN U19487 ( .B(clk), .A(\g.we_clk [13287]));
Q_ASSIGN U19488 ( .B(clk), .A(\g.we_clk [13286]));
Q_ASSIGN U19489 ( .B(clk), .A(\g.we_clk [13285]));
Q_ASSIGN U19490 ( .B(clk), .A(\g.we_clk [13284]));
Q_ASSIGN U19491 ( .B(clk), .A(\g.we_clk [13283]));
Q_ASSIGN U19492 ( .B(clk), .A(\g.we_clk [13282]));
Q_ASSIGN U19493 ( .B(clk), .A(\g.we_clk [13281]));
Q_ASSIGN U19494 ( .B(clk), .A(\g.we_clk [13280]));
Q_ASSIGN U19495 ( .B(clk), .A(\g.we_clk [13279]));
Q_ASSIGN U19496 ( .B(clk), .A(\g.we_clk [13278]));
Q_ASSIGN U19497 ( .B(clk), .A(\g.we_clk [13277]));
Q_ASSIGN U19498 ( .B(clk), .A(\g.we_clk [13276]));
Q_ASSIGN U19499 ( .B(clk), .A(\g.we_clk [13275]));
Q_ASSIGN U19500 ( .B(clk), .A(\g.we_clk [13274]));
Q_ASSIGN U19501 ( .B(clk), .A(\g.we_clk [13273]));
Q_ASSIGN U19502 ( .B(clk), .A(\g.we_clk [13272]));
Q_ASSIGN U19503 ( .B(clk), .A(\g.we_clk [13271]));
Q_ASSIGN U19504 ( .B(clk), .A(\g.we_clk [13270]));
Q_ASSIGN U19505 ( .B(clk), .A(\g.we_clk [13269]));
Q_ASSIGN U19506 ( .B(clk), .A(\g.we_clk [13268]));
Q_ASSIGN U19507 ( .B(clk), .A(\g.we_clk [13267]));
Q_ASSIGN U19508 ( .B(clk), .A(\g.we_clk [13266]));
Q_ASSIGN U19509 ( .B(clk), .A(\g.we_clk [13265]));
Q_ASSIGN U19510 ( .B(clk), .A(\g.we_clk [13264]));
Q_ASSIGN U19511 ( .B(clk), .A(\g.we_clk [13263]));
Q_ASSIGN U19512 ( .B(clk), .A(\g.we_clk [13262]));
Q_ASSIGN U19513 ( .B(clk), .A(\g.we_clk [13261]));
Q_ASSIGN U19514 ( .B(clk), .A(\g.we_clk [13260]));
Q_ASSIGN U19515 ( .B(clk), .A(\g.we_clk [13259]));
Q_ASSIGN U19516 ( .B(clk), .A(\g.we_clk [13258]));
Q_ASSIGN U19517 ( .B(clk), .A(\g.we_clk [13257]));
Q_ASSIGN U19518 ( .B(clk), .A(\g.we_clk [13256]));
Q_ASSIGN U19519 ( .B(clk), .A(\g.we_clk [13255]));
Q_ASSIGN U19520 ( .B(clk), .A(\g.we_clk [13254]));
Q_ASSIGN U19521 ( .B(clk), .A(\g.we_clk [13253]));
Q_ASSIGN U19522 ( .B(clk), .A(\g.we_clk [13252]));
Q_ASSIGN U19523 ( .B(clk), .A(\g.we_clk [13251]));
Q_ASSIGN U19524 ( .B(clk), .A(\g.we_clk [13250]));
Q_ASSIGN U19525 ( .B(clk), .A(\g.we_clk [13249]));
Q_ASSIGN U19526 ( .B(clk), .A(\g.we_clk [13248]));
Q_ASSIGN U19527 ( .B(clk), .A(\g.we_clk [13247]));
Q_ASSIGN U19528 ( .B(clk), .A(\g.we_clk [13246]));
Q_ASSIGN U19529 ( .B(clk), .A(\g.we_clk [13245]));
Q_ASSIGN U19530 ( .B(clk), .A(\g.we_clk [13244]));
Q_ASSIGN U19531 ( .B(clk), .A(\g.we_clk [13243]));
Q_ASSIGN U19532 ( .B(clk), .A(\g.we_clk [13242]));
Q_ASSIGN U19533 ( .B(clk), .A(\g.we_clk [13241]));
Q_ASSIGN U19534 ( .B(clk), .A(\g.we_clk [13240]));
Q_ASSIGN U19535 ( .B(clk), .A(\g.we_clk [13239]));
Q_ASSIGN U19536 ( .B(clk), .A(\g.we_clk [13238]));
Q_ASSIGN U19537 ( .B(clk), .A(\g.we_clk [13237]));
Q_ASSIGN U19538 ( .B(clk), .A(\g.we_clk [13236]));
Q_ASSIGN U19539 ( .B(clk), .A(\g.we_clk [13235]));
Q_ASSIGN U19540 ( .B(clk), .A(\g.we_clk [13234]));
Q_ASSIGN U19541 ( .B(clk), .A(\g.we_clk [13233]));
Q_ASSIGN U19542 ( .B(clk), .A(\g.we_clk [13232]));
Q_ASSIGN U19543 ( .B(clk), .A(\g.we_clk [13231]));
Q_ASSIGN U19544 ( .B(clk), .A(\g.we_clk [13230]));
Q_ASSIGN U19545 ( .B(clk), .A(\g.we_clk [13229]));
Q_ASSIGN U19546 ( .B(clk), .A(\g.we_clk [13228]));
Q_ASSIGN U19547 ( .B(clk), .A(\g.we_clk [13227]));
Q_ASSIGN U19548 ( .B(clk), .A(\g.we_clk [13226]));
Q_ASSIGN U19549 ( .B(clk), .A(\g.we_clk [13225]));
Q_ASSIGN U19550 ( .B(clk), .A(\g.we_clk [13224]));
Q_ASSIGN U19551 ( .B(clk), .A(\g.we_clk [13223]));
Q_ASSIGN U19552 ( .B(clk), .A(\g.we_clk [13222]));
Q_ASSIGN U19553 ( .B(clk), .A(\g.we_clk [13221]));
Q_ASSIGN U19554 ( .B(clk), .A(\g.we_clk [13220]));
Q_ASSIGN U19555 ( .B(clk), .A(\g.we_clk [13219]));
Q_ASSIGN U19556 ( .B(clk), .A(\g.we_clk [13218]));
Q_ASSIGN U19557 ( .B(clk), .A(\g.we_clk [13217]));
Q_ASSIGN U19558 ( .B(clk), .A(\g.we_clk [13216]));
Q_ASSIGN U19559 ( .B(clk), .A(\g.we_clk [13215]));
Q_ASSIGN U19560 ( .B(clk), .A(\g.we_clk [13214]));
Q_ASSIGN U19561 ( .B(clk), .A(\g.we_clk [13213]));
Q_ASSIGN U19562 ( .B(clk), .A(\g.we_clk [13212]));
Q_ASSIGN U19563 ( .B(clk), .A(\g.we_clk [13211]));
Q_ASSIGN U19564 ( .B(clk), .A(\g.we_clk [13210]));
Q_ASSIGN U19565 ( .B(clk), .A(\g.we_clk [13209]));
Q_ASSIGN U19566 ( .B(clk), .A(\g.we_clk [13208]));
Q_ASSIGN U19567 ( .B(clk), .A(\g.we_clk [13207]));
Q_ASSIGN U19568 ( .B(clk), .A(\g.we_clk [13206]));
Q_ASSIGN U19569 ( .B(clk), .A(\g.we_clk [13205]));
Q_ASSIGN U19570 ( .B(clk), .A(\g.we_clk [13204]));
Q_ASSIGN U19571 ( .B(clk), .A(\g.we_clk [13203]));
Q_ASSIGN U19572 ( .B(clk), .A(\g.we_clk [13202]));
Q_ASSIGN U19573 ( .B(clk), .A(\g.we_clk [13201]));
Q_ASSIGN U19574 ( .B(clk), .A(\g.we_clk [13200]));
Q_ASSIGN U19575 ( .B(clk), .A(\g.we_clk [13199]));
Q_ASSIGN U19576 ( .B(clk), .A(\g.we_clk [13198]));
Q_ASSIGN U19577 ( .B(clk), .A(\g.we_clk [13197]));
Q_ASSIGN U19578 ( .B(clk), .A(\g.we_clk [13196]));
Q_ASSIGN U19579 ( .B(clk), .A(\g.we_clk [13195]));
Q_ASSIGN U19580 ( .B(clk), .A(\g.we_clk [13194]));
Q_ASSIGN U19581 ( .B(clk), .A(\g.we_clk [13193]));
Q_ASSIGN U19582 ( .B(clk), .A(\g.we_clk [13192]));
Q_ASSIGN U19583 ( .B(clk), .A(\g.we_clk [13191]));
Q_ASSIGN U19584 ( .B(clk), .A(\g.we_clk [13190]));
Q_ASSIGN U19585 ( .B(clk), .A(\g.we_clk [13189]));
Q_ASSIGN U19586 ( .B(clk), .A(\g.we_clk [13188]));
Q_ASSIGN U19587 ( .B(clk), .A(\g.we_clk [13187]));
Q_ASSIGN U19588 ( .B(clk), .A(\g.we_clk [13186]));
Q_ASSIGN U19589 ( .B(clk), .A(\g.we_clk [13185]));
Q_ASSIGN U19590 ( .B(clk), .A(\g.we_clk [13184]));
Q_ASSIGN U19591 ( .B(clk), .A(\g.we_clk [13183]));
Q_ASSIGN U19592 ( .B(clk), .A(\g.we_clk [13182]));
Q_ASSIGN U19593 ( .B(clk), .A(\g.we_clk [13181]));
Q_ASSIGN U19594 ( .B(clk), .A(\g.we_clk [13180]));
Q_ASSIGN U19595 ( .B(clk), .A(\g.we_clk [13179]));
Q_ASSIGN U19596 ( .B(clk), .A(\g.we_clk [13178]));
Q_ASSIGN U19597 ( .B(clk), .A(\g.we_clk [13177]));
Q_ASSIGN U19598 ( .B(clk), .A(\g.we_clk [13176]));
Q_ASSIGN U19599 ( .B(clk), .A(\g.we_clk [13175]));
Q_ASSIGN U19600 ( .B(clk), .A(\g.we_clk [13174]));
Q_ASSIGN U19601 ( .B(clk), .A(\g.we_clk [13173]));
Q_ASSIGN U19602 ( .B(clk), .A(\g.we_clk [13172]));
Q_ASSIGN U19603 ( .B(clk), .A(\g.we_clk [13171]));
Q_ASSIGN U19604 ( .B(clk), .A(\g.we_clk [13170]));
Q_ASSIGN U19605 ( .B(clk), .A(\g.we_clk [13169]));
Q_ASSIGN U19606 ( .B(clk), .A(\g.we_clk [13168]));
Q_ASSIGN U19607 ( .B(clk), .A(\g.we_clk [13167]));
Q_ASSIGN U19608 ( .B(clk), .A(\g.we_clk [13166]));
Q_ASSIGN U19609 ( .B(clk), .A(\g.we_clk [13165]));
Q_ASSIGN U19610 ( .B(clk), .A(\g.we_clk [13164]));
Q_ASSIGN U19611 ( .B(clk), .A(\g.we_clk [13163]));
Q_ASSIGN U19612 ( .B(clk), .A(\g.we_clk [13162]));
Q_ASSIGN U19613 ( .B(clk), .A(\g.we_clk [13161]));
Q_ASSIGN U19614 ( .B(clk), .A(\g.we_clk [13160]));
Q_ASSIGN U19615 ( .B(clk), .A(\g.we_clk [13159]));
Q_ASSIGN U19616 ( .B(clk), .A(\g.we_clk [13158]));
Q_ASSIGN U19617 ( .B(clk), .A(\g.we_clk [13157]));
Q_ASSIGN U19618 ( .B(clk), .A(\g.we_clk [13156]));
Q_ASSIGN U19619 ( .B(clk), .A(\g.we_clk [13155]));
Q_ASSIGN U19620 ( .B(clk), .A(\g.we_clk [13154]));
Q_ASSIGN U19621 ( .B(clk), .A(\g.we_clk [13153]));
Q_ASSIGN U19622 ( .B(clk), .A(\g.we_clk [13152]));
Q_ASSIGN U19623 ( .B(clk), .A(\g.we_clk [13151]));
Q_ASSIGN U19624 ( .B(clk), .A(\g.we_clk [13150]));
Q_ASSIGN U19625 ( .B(clk), .A(\g.we_clk [13149]));
Q_ASSIGN U19626 ( .B(clk), .A(\g.we_clk [13148]));
Q_ASSIGN U19627 ( .B(clk), .A(\g.we_clk [13147]));
Q_ASSIGN U19628 ( .B(clk), .A(\g.we_clk [13146]));
Q_ASSIGN U19629 ( .B(clk), .A(\g.we_clk [13145]));
Q_ASSIGN U19630 ( .B(clk), .A(\g.we_clk [13144]));
Q_ASSIGN U19631 ( .B(clk), .A(\g.we_clk [13143]));
Q_ASSIGN U19632 ( .B(clk), .A(\g.we_clk [13142]));
Q_ASSIGN U19633 ( .B(clk), .A(\g.we_clk [13141]));
Q_ASSIGN U19634 ( .B(clk), .A(\g.we_clk [13140]));
Q_ASSIGN U19635 ( .B(clk), .A(\g.we_clk [13139]));
Q_ASSIGN U19636 ( .B(clk), .A(\g.we_clk [13138]));
Q_ASSIGN U19637 ( .B(clk), .A(\g.we_clk [13137]));
Q_ASSIGN U19638 ( .B(clk), .A(\g.we_clk [13136]));
Q_ASSIGN U19639 ( .B(clk), .A(\g.we_clk [13135]));
Q_ASSIGN U19640 ( .B(clk), .A(\g.we_clk [13134]));
Q_ASSIGN U19641 ( .B(clk), .A(\g.we_clk [13133]));
Q_ASSIGN U19642 ( .B(clk), .A(\g.we_clk [13132]));
Q_ASSIGN U19643 ( .B(clk), .A(\g.we_clk [13131]));
Q_ASSIGN U19644 ( .B(clk), .A(\g.we_clk [13130]));
Q_ASSIGN U19645 ( .B(clk), .A(\g.we_clk [13129]));
Q_ASSIGN U19646 ( .B(clk), .A(\g.we_clk [13128]));
Q_ASSIGN U19647 ( .B(clk), .A(\g.we_clk [13127]));
Q_ASSIGN U19648 ( .B(clk), .A(\g.we_clk [13126]));
Q_ASSIGN U19649 ( .B(clk), .A(\g.we_clk [13125]));
Q_ASSIGN U19650 ( .B(clk), .A(\g.we_clk [13124]));
Q_ASSIGN U19651 ( .B(clk), .A(\g.we_clk [13123]));
Q_ASSIGN U19652 ( .B(clk), .A(\g.we_clk [13122]));
Q_ASSIGN U19653 ( .B(clk), .A(\g.we_clk [13121]));
Q_ASSIGN U19654 ( .B(clk), .A(\g.we_clk [13120]));
Q_ASSIGN U19655 ( .B(clk), .A(\g.we_clk [13119]));
Q_ASSIGN U19656 ( .B(clk), .A(\g.we_clk [13118]));
Q_ASSIGN U19657 ( .B(clk), .A(\g.we_clk [13117]));
Q_ASSIGN U19658 ( .B(clk), .A(\g.we_clk [13116]));
Q_ASSIGN U19659 ( .B(clk), .A(\g.we_clk [13115]));
Q_ASSIGN U19660 ( .B(clk), .A(\g.we_clk [13114]));
Q_ASSIGN U19661 ( .B(clk), .A(\g.we_clk [13113]));
Q_ASSIGN U19662 ( .B(clk), .A(\g.we_clk [13112]));
Q_ASSIGN U19663 ( .B(clk), .A(\g.we_clk [13111]));
Q_ASSIGN U19664 ( .B(clk), .A(\g.we_clk [13110]));
Q_ASSIGN U19665 ( .B(clk), .A(\g.we_clk [13109]));
Q_ASSIGN U19666 ( .B(clk), .A(\g.we_clk [13108]));
Q_ASSIGN U19667 ( .B(clk), .A(\g.we_clk [13107]));
Q_ASSIGN U19668 ( .B(clk), .A(\g.we_clk [13106]));
Q_ASSIGN U19669 ( .B(clk), .A(\g.we_clk [13105]));
Q_ASSIGN U19670 ( .B(clk), .A(\g.we_clk [13104]));
Q_ASSIGN U19671 ( .B(clk), .A(\g.we_clk [13103]));
Q_ASSIGN U19672 ( .B(clk), .A(\g.we_clk [13102]));
Q_ASSIGN U19673 ( .B(clk), .A(\g.we_clk [13101]));
Q_ASSIGN U19674 ( .B(clk), .A(\g.we_clk [13100]));
Q_ASSIGN U19675 ( .B(clk), .A(\g.we_clk [13099]));
Q_ASSIGN U19676 ( .B(clk), .A(\g.we_clk [13098]));
Q_ASSIGN U19677 ( .B(clk), .A(\g.we_clk [13097]));
Q_ASSIGN U19678 ( .B(clk), .A(\g.we_clk [13096]));
Q_ASSIGN U19679 ( .B(clk), .A(\g.we_clk [13095]));
Q_ASSIGN U19680 ( .B(clk), .A(\g.we_clk [13094]));
Q_ASSIGN U19681 ( .B(clk), .A(\g.we_clk [13093]));
Q_ASSIGN U19682 ( .B(clk), .A(\g.we_clk [13092]));
Q_ASSIGN U19683 ( .B(clk), .A(\g.we_clk [13091]));
Q_ASSIGN U19684 ( .B(clk), .A(\g.we_clk [13090]));
Q_ASSIGN U19685 ( .B(clk), .A(\g.we_clk [13089]));
Q_ASSIGN U19686 ( .B(clk), .A(\g.we_clk [13088]));
Q_ASSIGN U19687 ( .B(clk), .A(\g.we_clk [13087]));
Q_ASSIGN U19688 ( .B(clk), .A(\g.we_clk [13086]));
Q_ASSIGN U19689 ( .B(clk), .A(\g.we_clk [13085]));
Q_ASSIGN U19690 ( .B(clk), .A(\g.we_clk [13084]));
Q_ASSIGN U19691 ( .B(clk), .A(\g.we_clk [13083]));
Q_ASSIGN U19692 ( .B(clk), .A(\g.we_clk [13082]));
Q_ASSIGN U19693 ( .B(clk), .A(\g.we_clk [13081]));
Q_ASSIGN U19694 ( .B(clk), .A(\g.we_clk [13080]));
Q_ASSIGN U19695 ( .B(clk), .A(\g.we_clk [13079]));
Q_ASSIGN U19696 ( .B(clk), .A(\g.we_clk [13078]));
Q_ASSIGN U19697 ( .B(clk), .A(\g.we_clk [13077]));
Q_ASSIGN U19698 ( .B(clk), .A(\g.we_clk [13076]));
Q_ASSIGN U19699 ( .B(clk), .A(\g.we_clk [13075]));
Q_ASSIGN U19700 ( .B(clk), .A(\g.we_clk [13074]));
Q_ASSIGN U19701 ( .B(clk), .A(\g.we_clk [13073]));
Q_ASSIGN U19702 ( .B(clk), .A(\g.we_clk [13072]));
Q_ASSIGN U19703 ( .B(clk), .A(\g.we_clk [13071]));
Q_ASSIGN U19704 ( .B(clk), .A(\g.we_clk [13070]));
Q_ASSIGN U19705 ( .B(clk), .A(\g.we_clk [13069]));
Q_ASSIGN U19706 ( .B(clk), .A(\g.we_clk [13068]));
Q_ASSIGN U19707 ( .B(clk), .A(\g.we_clk [13067]));
Q_ASSIGN U19708 ( .B(clk), .A(\g.we_clk [13066]));
Q_ASSIGN U19709 ( .B(clk), .A(\g.we_clk [13065]));
Q_ASSIGN U19710 ( .B(clk), .A(\g.we_clk [13064]));
Q_ASSIGN U19711 ( .B(clk), .A(\g.we_clk [13063]));
Q_ASSIGN U19712 ( .B(clk), .A(\g.we_clk [13062]));
Q_ASSIGN U19713 ( .B(clk), .A(\g.we_clk [13061]));
Q_ASSIGN U19714 ( .B(clk), .A(\g.we_clk [13060]));
Q_ASSIGN U19715 ( .B(clk), .A(\g.we_clk [13059]));
Q_ASSIGN U19716 ( .B(clk), .A(\g.we_clk [13058]));
Q_ASSIGN U19717 ( .B(clk), .A(\g.we_clk [13057]));
Q_ASSIGN U19718 ( .B(clk), .A(\g.we_clk [13056]));
Q_ASSIGN U19719 ( .B(clk), .A(\g.we_clk [13055]));
Q_ASSIGN U19720 ( .B(clk), .A(\g.we_clk [13054]));
Q_ASSIGN U19721 ( .B(clk), .A(\g.we_clk [13053]));
Q_ASSIGN U19722 ( .B(clk), .A(\g.we_clk [13052]));
Q_ASSIGN U19723 ( .B(clk), .A(\g.we_clk [13051]));
Q_ASSIGN U19724 ( .B(clk), .A(\g.we_clk [13050]));
Q_ASSIGN U19725 ( .B(clk), .A(\g.we_clk [13049]));
Q_ASSIGN U19726 ( .B(clk), .A(\g.we_clk [13048]));
Q_ASSIGN U19727 ( .B(clk), .A(\g.we_clk [13047]));
Q_ASSIGN U19728 ( .B(clk), .A(\g.we_clk [13046]));
Q_ASSIGN U19729 ( .B(clk), .A(\g.we_clk [13045]));
Q_ASSIGN U19730 ( .B(clk), .A(\g.we_clk [13044]));
Q_ASSIGN U19731 ( .B(clk), .A(\g.we_clk [13043]));
Q_ASSIGN U19732 ( .B(clk), .A(\g.we_clk [13042]));
Q_ASSIGN U19733 ( .B(clk), .A(\g.we_clk [13041]));
Q_ASSIGN U19734 ( .B(clk), .A(\g.we_clk [13040]));
Q_ASSIGN U19735 ( .B(clk), .A(\g.we_clk [13039]));
Q_ASSIGN U19736 ( .B(clk), .A(\g.we_clk [13038]));
Q_ASSIGN U19737 ( .B(clk), .A(\g.we_clk [13037]));
Q_ASSIGN U19738 ( .B(clk), .A(\g.we_clk [13036]));
Q_ASSIGN U19739 ( .B(clk), .A(\g.we_clk [13035]));
Q_ASSIGN U19740 ( .B(clk), .A(\g.we_clk [13034]));
Q_ASSIGN U19741 ( .B(clk), .A(\g.we_clk [13033]));
Q_ASSIGN U19742 ( .B(clk), .A(\g.we_clk [13032]));
Q_ASSIGN U19743 ( .B(clk), .A(\g.we_clk [13031]));
Q_ASSIGN U19744 ( .B(clk), .A(\g.we_clk [13030]));
Q_ASSIGN U19745 ( .B(clk), .A(\g.we_clk [13029]));
Q_ASSIGN U19746 ( .B(clk), .A(\g.we_clk [13028]));
Q_ASSIGN U19747 ( .B(clk), .A(\g.we_clk [13027]));
Q_ASSIGN U19748 ( .B(clk), .A(\g.we_clk [13026]));
Q_ASSIGN U19749 ( .B(clk), .A(\g.we_clk [13025]));
Q_ASSIGN U19750 ( .B(clk), .A(\g.we_clk [13024]));
Q_ASSIGN U19751 ( .B(clk), .A(\g.we_clk [13023]));
Q_ASSIGN U19752 ( .B(clk), .A(\g.we_clk [13022]));
Q_ASSIGN U19753 ( .B(clk), .A(\g.we_clk [13021]));
Q_ASSIGN U19754 ( .B(clk), .A(\g.we_clk [13020]));
Q_ASSIGN U19755 ( .B(clk), .A(\g.we_clk [13019]));
Q_ASSIGN U19756 ( .B(clk), .A(\g.we_clk [13018]));
Q_ASSIGN U19757 ( .B(clk), .A(\g.we_clk [13017]));
Q_ASSIGN U19758 ( .B(clk), .A(\g.we_clk [13016]));
Q_ASSIGN U19759 ( .B(clk), .A(\g.we_clk [13015]));
Q_ASSIGN U19760 ( .B(clk), .A(\g.we_clk [13014]));
Q_ASSIGN U19761 ( .B(clk), .A(\g.we_clk [13013]));
Q_ASSIGN U19762 ( .B(clk), .A(\g.we_clk [13012]));
Q_ASSIGN U19763 ( .B(clk), .A(\g.we_clk [13011]));
Q_ASSIGN U19764 ( .B(clk), .A(\g.we_clk [13010]));
Q_ASSIGN U19765 ( .B(clk), .A(\g.we_clk [13009]));
Q_ASSIGN U19766 ( .B(clk), .A(\g.we_clk [13008]));
Q_ASSIGN U19767 ( .B(clk), .A(\g.we_clk [13007]));
Q_ASSIGN U19768 ( .B(clk), .A(\g.we_clk [13006]));
Q_ASSIGN U19769 ( .B(clk), .A(\g.we_clk [13005]));
Q_ASSIGN U19770 ( .B(clk), .A(\g.we_clk [13004]));
Q_ASSIGN U19771 ( .B(clk), .A(\g.we_clk [13003]));
Q_ASSIGN U19772 ( .B(clk), .A(\g.we_clk [13002]));
Q_ASSIGN U19773 ( .B(clk), .A(\g.we_clk [13001]));
Q_ASSIGN U19774 ( .B(clk), .A(\g.we_clk [13000]));
Q_ASSIGN U19775 ( .B(clk), .A(\g.we_clk [12999]));
Q_ASSIGN U19776 ( .B(clk), .A(\g.we_clk [12998]));
Q_ASSIGN U19777 ( .B(clk), .A(\g.we_clk [12997]));
Q_ASSIGN U19778 ( .B(clk), .A(\g.we_clk [12996]));
Q_ASSIGN U19779 ( .B(clk), .A(\g.we_clk [12995]));
Q_ASSIGN U19780 ( .B(clk), .A(\g.we_clk [12994]));
Q_ASSIGN U19781 ( .B(clk), .A(\g.we_clk [12993]));
Q_ASSIGN U19782 ( .B(clk), .A(\g.we_clk [12992]));
Q_ASSIGN U19783 ( .B(clk), .A(\g.we_clk [12991]));
Q_ASSIGN U19784 ( .B(clk), .A(\g.we_clk [12990]));
Q_ASSIGN U19785 ( .B(clk), .A(\g.we_clk [12989]));
Q_ASSIGN U19786 ( .B(clk), .A(\g.we_clk [12988]));
Q_ASSIGN U19787 ( .B(clk), .A(\g.we_clk [12987]));
Q_ASSIGN U19788 ( .B(clk), .A(\g.we_clk [12986]));
Q_ASSIGN U19789 ( .B(clk), .A(\g.we_clk [12985]));
Q_ASSIGN U19790 ( .B(clk), .A(\g.we_clk [12984]));
Q_ASSIGN U19791 ( .B(clk), .A(\g.we_clk [12983]));
Q_ASSIGN U19792 ( .B(clk), .A(\g.we_clk [12982]));
Q_ASSIGN U19793 ( .B(clk), .A(\g.we_clk [12981]));
Q_ASSIGN U19794 ( .B(clk), .A(\g.we_clk [12980]));
Q_ASSIGN U19795 ( .B(clk), .A(\g.we_clk [12979]));
Q_ASSIGN U19796 ( .B(clk), .A(\g.we_clk [12978]));
Q_ASSIGN U19797 ( .B(clk), .A(\g.we_clk [12977]));
Q_ASSIGN U19798 ( .B(clk), .A(\g.we_clk [12976]));
Q_ASSIGN U19799 ( .B(clk), .A(\g.we_clk [12975]));
Q_ASSIGN U19800 ( .B(clk), .A(\g.we_clk [12974]));
Q_ASSIGN U19801 ( .B(clk), .A(\g.we_clk [12973]));
Q_ASSIGN U19802 ( .B(clk), .A(\g.we_clk [12972]));
Q_ASSIGN U19803 ( .B(clk), .A(\g.we_clk [12971]));
Q_ASSIGN U19804 ( .B(clk), .A(\g.we_clk [12970]));
Q_ASSIGN U19805 ( .B(clk), .A(\g.we_clk [12969]));
Q_ASSIGN U19806 ( .B(clk), .A(\g.we_clk [12968]));
Q_ASSIGN U19807 ( .B(clk), .A(\g.we_clk [12967]));
Q_ASSIGN U19808 ( .B(clk), .A(\g.we_clk [12966]));
Q_ASSIGN U19809 ( .B(clk), .A(\g.we_clk [12965]));
Q_ASSIGN U19810 ( .B(clk), .A(\g.we_clk [12964]));
Q_ASSIGN U19811 ( .B(clk), .A(\g.we_clk [12963]));
Q_ASSIGN U19812 ( .B(clk), .A(\g.we_clk [12962]));
Q_ASSIGN U19813 ( .B(clk), .A(\g.we_clk [12961]));
Q_ASSIGN U19814 ( .B(clk), .A(\g.we_clk [12960]));
Q_ASSIGN U19815 ( .B(clk), .A(\g.we_clk [12959]));
Q_ASSIGN U19816 ( .B(clk), .A(\g.we_clk [12958]));
Q_ASSIGN U19817 ( .B(clk), .A(\g.we_clk [12957]));
Q_ASSIGN U19818 ( .B(clk), .A(\g.we_clk [12956]));
Q_ASSIGN U19819 ( .B(clk), .A(\g.we_clk [12955]));
Q_ASSIGN U19820 ( .B(clk), .A(\g.we_clk [12954]));
Q_ASSIGN U19821 ( .B(clk), .A(\g.we_clk [12953]));
Q_ASSIGN U19822 ( .B(clk), .A(\g.we_clk [12952]));
Q_ASSIGN U19823 ( .B(clk), .A(\g.we_clk [12951]));
Q_ASSIGN U19824 ( .B(clk), .A(\g.we_clk [12950]));
Q_ASSIGN U19825 ( .B(clk), .A(\g.we_clk [12949]));
Q_ASSIGN U19826 ( .B(clk), .A(\g.we_clk [12948]));
Q_ASSIGN U19827 ( .B(clk), .A(\g.we_clk [12947]));
Q_ASSIGN U19828 ( .B(clk), .A(\g.we_clk [12946]));
Q_ASSIGN U19829 ( .B(clk), .A(\g.we_clk [12945]));
Q_ASSIGN U19830 ( .B(clk), .A(\g.we_clk [12944]));
Q_ASSIGN U19831 ( .B(clk), .A(\g.we_clk [12943]));
Q_ASSIGN U19832 ( .B(clk), .A(\g.we_clk [12942]));
Q_ASSIGN U19833 ( .B(clk), .A(\g.we_clk [12941]));
Q_ASSIGN U19834 ( .B(clk), .A(\g.we_clk [12940]));
Q_ASSIGN U19835 ( .B(clk), .A(\g.we_clk [12939]));
Q_ASSIGN U19836 ( .B(clk), .A(\g.we_clk [12938]));
Q_ASSIGN U19837 ( .B(clk), .A(\g.we_clk [12937]));
Q_ASSIGN U19838 ( .B(clk), .A(\g.we_clk [12936]));
Q_ASSIGN U19839 ( .B(clk), .A(\g.we_clk [12935]));
Q_ASSIGN U19840 ( .B(clk), .A(\g.we_clk [12934]));
Q_ASSIGN U19841 ( .B(clk), .A(\g.we_clk [12933]));
Q_ASSIGN U19842 ( .B(clk), .A(\g.we_clk [12932]));
Q_ASSIGN U19843 ( .B(clk), .A(\g.we_clk [12931]));
Q_ASSIGN U19844 ( .B(clk), .A(\g.we_clk [12930]));
Q_ASSIGN U19845 ( .B(clk), .A(\g.we_clk [12929]));
Q_ASSIGN U19846 ( .B(clk), .A(\g.we_clk [12928]));
Q_ASSIGN U19847 ( .B(clk), .A(\g.we_clk [12927]));
Q_ASSIGN U19848 ( .B(clk), .A(\g.we_clk [12926]));
Q_ASSIGN U19849 ( .B(clk), .A(\g.we_clk [12925]));
Q_ASSIGN U19850 ( .B(clk), .A(\g.we_clk [12924]));
Q_ASSIGN U19851 ( .B(clk), .A(\g.we_clk [12923]));
Q_ASSIGN U19852 ( .B(clk), .A(\g.we_clk [12922]));
Q_ASSIGN U19853 ( .B(clk), .A(\g.we_clk [12921]));
Q_ASSIGN U19854 ( .B(clk), .A(\g.we_clk [12920]));
Q_ASSIGN U19855 ( .B(clk), .A(\g.we_clk [12919]));
Q_ASSIGN U19856 ( .B(clk), .A(\g.we_clk [12918]));
Q_ASSIGN U19857 ( .B(clk), .A(\g.we_clk [12917]));
Q_ASSIGN U19858 ( .B(clk), .A(\g.we_clk [12916]));
Q_ASSIGN U19859 ( .B(clk), .A(\g.we_clk [12915]));
Q_ASSIGN U19860 ( .B(clk), .A(\g.we_clk [12914]));
Q_ASSIGN U19861 ( .B(clk), .A(\g.we_clk [12913]));
Q_ASSIGN U19862 ( .B(clk), .A(\g.we_clk [12912]));
Q_ASSIGN U19863 ( .B(clk), .A(\g.we_clk [12911]));
Q_ASSIGN U19864 ( .B(clk), .A(\g.we_clk [12910]));
Q_ASSIGN U19865 ( .B(clk), .A(\g.we_clk [12909]));
Q_ASSIGN U19866 ( .B(clk), .A(\g.we_clk [12908]));
Q_ASSIGN U19867 ( .B(clk), .A(\g.we_clk [12907]));
Q_ASSIGN U19868 ( .B(clk), .A(\g.we_clk [12906]));
Q_ASSIGN U19869 ( .B(clk), .A(\g.we_clk [12905]));
Q_ASSIGN U19870 ( .B(clk), .A(\g.we_clk [12904]));
Q_ASSIGN U19871 ( .B(clk), .A(\g.we_clk [12903]));
Q_ASSIGN U19872 ( .B(clk), .A(\g.we_clk [12902]));
Q_ASSIGN U19873 ( .B(clk), .A(\g.we_clk [12901]));
Q_ASSIGN U19874 ( .B(clk), .A(\g.we_clk [12900]));
Q_ASSIGN U19875 ( .B(clk), .A(\g.we_clk [12899]));
Q_ASSIGN U19876 ( .B(clk), .A(\g.we_clk [12898]));
Q_ASSIGN U19877 ( .B(clk), .A(\g.we_clk [12897]));
Q_ASSIGN U19878 ( .B(clk), .A(\g.we_clk [12896]));
Q_ASSIGN U19879 ( .B(clk), .A(\g.we_clk [12895]));
Q_ASSIGN U19880 ( .B(clk), .A(\g.we_clk [12894]));
Q_ASSIGN U19881 ( .B(clk), .A(\g.we_clk [12893]));
Q_ASSIGN U19882 ( .B(clk), .A(\g.we_clk [12892]));
Q_ASSIGN U19883 ( .B(clk), .A(\g.we_clk [12891]));
Q_ASSIGN U19884 ( .B(clk), .A(\g.we_clk [12890]));
Q_ASSIGN U19885 ( .B(clk), .A(\g.we_clk [12889]));
Q_ASSIGN U19886 ( .B(clk), .A(\g.we_clk [12888]));
Q_ASSIGN U19887 ( .B(clk), .A(\g.we_clk [12887]));
Q_ASSIGN U19888 ( .B(clk), .A(\g.we_clk [12886]));
Q_ASSIGN U19889 ( .B(clk), .A(\g.we_clk [12885]));
Q_ASSIGN U19890 ( .B(clk), .A(\g.we_clk [12884]));
Q_ASSIGN U19891 ( .B(clk), .A(\g.we_clk [12883]));
Q_ASSIGN U19892 ( .B(clk), .A(\g.we_clk [12882]));
Q_ASSIGN U19893 ( .B(clk), .A(\g.we_clk [12881]));
Q_ASSIGN U19894 ( .B(clk), .A(\g.we_clk [12880]));
Q_ASSIGN U19895 ( .B(clk), .A(\g.we_clk [12879]));
Q_ASSIGN U19896 ( .B(clk), .A(\g.we_clk [12878]));
Q_ASSIGN U19897 ( .B(clk), .A(\g.we_clk [12877]));
Q_ASSIGN U19898 ( .B(clk), .A(\g.we_clk [12876]));
Q_ASSIGN U19899 ( .B(clk), .A(\g.we_clk [12875]));
Q_ASSIGN U19900 ( .B(clk), .A(\g.we_clk [12874]));
Q_ASSIGN U19901 ( .B(clk), .A(\g.we_clk [12873]));
Q_ASSIGN U19902 ( .B(clk), .A(\g.we_clk [12872]));
Q_ASSIGN U19903 ( .B(clk), .A(\g.we_clk [12871]));
Q_ASSIGN U19904 ( .B(clk), .A(\g.we_clk [12870]));
Q_ASSIGN U19905 ( .B(clk), .A(\g.we_clk [12869]));
Q_ASSIGN U19906 ( .B(clk), .A(\g.we_clk [12868]));
Q_ASSIGN U19907 ( .B(clk), .A(\g.we_clk [12867]));
Q_ASSIGN U19908 ( .B(clk), .A(\g.we_clk [12866]));
Q_ASSIGN U19909 ( .B(clk), .A(\g.we_clk [12865]));
Q_ASSIGN U19910 ( .B(clk), .A(\g.we_clk [12864]));
Q_ASSIGN U19911 ( .B(clk), .A(\g.we_clk [12863]));
Q_ASSIGN U19912 ( .B(clk), .A(\g.we_clk [12862]));
Q_ASSIGN U19913 ( .B(clk), .A(\g.we_clk [12861]));
Q_ASSIGN U19914 ( .B(clk), .A(\g.we_clk [12860]));
Q_ASSIGN U19915 ( .B(clk), .A(\g.we_clk [12859]));
Q_ASSIGN U19916 ( .B(clk), .A(\g.we_clk [12858]));
Q_ASSIGN U19917 ( .B(clk), .A(\g.we_clk [12857]));
Q_ASSIGN U19918 ( .B(clk), .A(\g.we_clk [12856]));
Q_ASSIGN U19919 ( .B(clk), .A(\g.we_clk [12855]));
Q_ASSIGN U19920 ( .B(clk), .A(\g.we_clk [12854]));
Q_ASSIGN U19921 ( .B(clk), .A(\g.we_clk [12853]));
Q_ASSIGN U19922 ( .B(clk), .A(\g.we_clk [12852]));
Q_ASSIGN U19923 ( .B(clk), .A(\g.we_clk [12851]));
Q_ASSIGN U19924 ( .B(clk), .A(\g.we_clk [12850]));
Q_ASSIGN U19925 ( .B(clk), .A(\g.we_clk [12849]));
Q_ASSIGN U19926 ( .B(clk), .A(\g.we_clk [12848]));
Q_ASSIGN U19927 ( .B(clk), .A(\g.we_clk [12847]));
Q_ASSIGN U19928 ( .B(clk), .A(\g.we_clk [12846]));
Q_ASSIGN U19929 ( .B(clk), .A(\g.we_clk [12845]));
Q_ASSIGN U19930 ( .B(clk), .A(\g.we_clk [12844]));
Q_ASSIGN U19931 ( .B(clk), .A(\g.we_clk [12843]));
Q_ASSIGN U19932 ( .B(clk), .A(\g.we_clk [12842]));
Q_ASSIGN U19933 ( .B(clk), .A(\g.we_clk [12841]));
Q_ASSIGN U19934 ( .B(clk), .A(\g.we_clk [12840]));
Q_ASSIGN U19935 ( .B(clk), .A(\g.we_clk [12839]));
Q_ASSIGN U19936 ( .B(clk), .A(\g.we_clk [12838]));
Q_ASSIGN U19937 ( .B(clk), .A(\g.we_clk [12837]));
Q_ASSIGN U19938 ( .B(clk), .A(\g.we_clk [12836]));
Q_ASSIGN U19939 ( .B(clk), .A(\g.we_clk [12835]));
Q_ASSIGN U19940 ( .B(clk), .A(\g.we_clk [12834]));
Q_ASSIGN U19941 ( .B(clk), .A(\g.we_clk [12833]));
Q_ASSIGN U19942 ( .B(clk), .A(\g.we_clk [12832]));
Q_ASSIGN U19943 ( .B(clk), .A(\g.we_clk [12831]));
Q_ASSIGN U19944 ( .B(clk), .A(\g.we_clk [12830]));
Q_ASSIGN U19945 ( .B(clk), .A(\g.we_clk [12829]));
Q_ASSIGN U19946 ( .B(clk), .A(\g.we_clk [12828]));
Q_ASSIGN U19947 ( .B(clk), .A(\g.we_clk [12827]));
Q_ASSIGN U19948 ( .B(clk), .A(\g.we_clk [12826]));
Q_ASSIGN U19949 ( .B(clk), .A(\g.we_clk [12825]));
Q_ASSIGN U19950 ( .B(clk), .A(\g.we_clk [12824]));
Q_ASSIGN U19951 ( .B(clk), .A(\g.we_clk [12823]));
Q_ASSIGN U19952 ( .B(clk), .A(\g.we_clk [12822]));
Q_ASSIGN U19953 ( .B(clk), .A(\g.we_clk [12821]));
Q_ASSIGN U19954 ( .B(clk), .A(\g.we_clk [12820]));
Q_ASSIGN U19955 ( .B(clk), .A(\g.we_clk [12819]));
Q_ASSIGN U19956 ( .B(clk), .A(\g.we_clk [12818]));
Q_ASSIGN U19957 ( .B(clk), .A(\g.we_clk [12817]));
Q_ASSIGN U19958 ( .B(clk), .A(\g.we_clk [12816]));
Q_ASSIGN U19959 ( .B(clk), .A(\g.we_clk [12815]));
Q_ASSIGN U19960 ( .B(clk), .A(\g.we_clk [12814]));
Q_ASSIGN U19961 ( .B(clk), .A(\g.we_clk [12813]));
Q_ASSIGN U19962 ( .B(clk), .A(\g.we_clk [12812]));
Q_ASSIGN U19963 ( .B(clk), .A(\g.we_clk [12811]));
Q_ASSIGN U19964 ( .B(clk), .A(\g.we_clk [12810]));
Q_ASSIGN U19965 ( .B(clk), .A(\g.we_clk [12809]));
Q_ASSIGN U19966 ( .B(clk), .A(\g.we_clk [12808]));
Q_ASSIGN U19967 ( .B(clk), .A(\g.we_clk [12807]));
Q_ASSIGN U19968 ( .B(clk), .A(\g.we_clk [12806]));
Q_ASSIGN U19969 ( .B(clk), .A(\g.we_clk [12805]));
Q_ASSIGN U19970 ( .B(clk), .A(\g.we_clk [12804]));
Q_ASSIGN U19971 ( .B(clk), .A(\g.we_clk [12803]));
Q_ASSIGN U19972 ( .B(clk), .A(\g.we_clk [12802]));
Q_ASSIGN U19973 ( .B(clk), .A(\g.we_clk [12801]));
Q_ASSIGN U19974 ( .B(clk), .A(\g.we_clk [12800]));
Q_ASSIGN U19975 ( .B(clk), .A(\g.we_clk [12799]));
Q_ASSIGN U19976 ( .B(clk), .A(\g.we_clk [12798]));
Q_ASSIGN U19977 ( .B(clk), .A(\g.we_clk [12797]));
Q_ASSIGN U19978 ( .B(clk), .A(\g.we_clk [12796]));
Q_ASSIGN U19979 ( .B(clk), .A(\g.we_clk [12795]));
Q_ASSIGN U19980 ( .B(clk), .A(\g.we_clk [12794]));
Q_ASSIGN U19981 ( .B(clk), .A(\g.we_clk [12793]));
Q_ASSIGN U19982 ( .B(clk), .A(\g.we_clk [12792]));
Q_ASSIGN U19983 ( .B(clk), .A(\g.we_clk [12791]));
Q_ASSIGN U19984 ( .B(clk), .A(\g.we_clk [12790]));
Q_ASSIGN U19985 ( .B(clk), .A(\g.we_clk [12789]));
Q_ASSIGN U19986 ( .B(clk), .A(\g.we_clk [12788]));
Q_ASSIGN U19987 ( .B(clk), .A(\g.we_clk [12787]));
Q_ASSIGN U19988 ( .B(clk), .A(\g.we_clk [12786]));
Q_ASSIGN U19989 ( .B(clk), .A(\g.we_clk [12785]));
Q_ASSIGN U19990 ( .B(clk), .A(\g.we_clk [12784]));
Q_ASSIGN U19991 ( .B(clk), .A(\g.we_clk [12783]));
Q_ASSIGN U19992 ( .B(clk), .A(\g.we_clk [12782]));
Q_ASSIGN U19993 ( .B(clk), .A(\g.we_clk [12781]));
Q_ASSIGN U19994 ( .B(clk), .A(\g.we_clk [12780]));
Q_ASSIGN U19995 ( .B(clk), .A(\g.we_clk [12779]));
Q_ASSIGN U19996 ( .B(clk), .A(\g.we_clk [12778]));
Q_ASSIGN U19997 ( .B(clk), .A(\g.we_clk [12777]));
Q_ASSIGN U19998 ( .B(clk), .A(\g.we_clk [12776]));
Q_ASSIGN U19999 ( .B(clk), .A(\g.we_clk [12775]));
Q_ASSIGN U20000 ( .B(clk), .A(\g.we_clk [12774]));
Q_ASSIGN U20001 ( .B(clk), .A(\g.we_clk [12773]));
Q_ASSIGN U20002 ( .B(clk), .A(\g.we_clk [12772]));
Q_ASSIGN U20003 ( .B(clk), .A(\g.we_clk [12771]));
Q_ASSIGN U20004 ( .B(clk), .A(\g.we_clk [12770]));
Q_ASSIGN U20005 ( .B(clk), .A(\g.we_clk [12769]));
Q_ASSIGN U20006 ( .B(clk), .A(\g.we_clk [12768]));
Q_ASSIGN U20007 ( .B(clk), .A(\g.we_clk [12767]));
Q_ASSIGN U20008 ( .B(clk), .A(\g.we_clk [12766]));
Q_ASSIGN U20009 ( .B(clk), .A(\g.we_clk [12765]));
Q_ASSIGN U20010 ( .B(clk), .A(\g.we_clk [12764]));
Q_ASSIGN U20011 ( .B(clk), .A(\g.we_clk [12763]));
Q_ASSIGN U20012 ( .B(clk), .A(\g.we_clk [12762]));
Q_ASSIGN U20013 ( .B(clk), .A(\g.we_clk [12761]));
Q_ASSIGN U20014 ( .B(clk), .A(\g.we_clk [12760]));
Q_ASSIGN U20015 ( .B(clk), .A(\g.we_clk [12759]));
Q_ASSIGN U20016 ( .B(clk), .A(\g.we_clk [12758]));
Q_ASSIGN U20017 ( .B(clk), .A(\g.we_clk [12757]));
Q_ASSIGN U20018 ( .B(clk), .A(\g.we_clk [12756]));
Q_ASSIGN U20019 ( .B(clk), .A(\g.we_clk [12755]));
Q_ASSIGN U20020 ( .B(clk), .A(\g.we_clk [12754]));
Q_ASSIGN U20021 ( .B(clk), .A(\g.we_clk [12753]));
Q_ASSIGN U20022 ( .B(clk), .A(\g.we_clk [12752]));
Q_ASSIGN U20023 ( .B(clk), .A(\g.we_clk [12751]));
Q_ASSIGN U20024 ( .B(clk), .A(\g.we_clk [12750]));
Q_ASSIGN U20025 ( .B(clk), .A(\g.we_clk [12749]));
Q_ASSIGN U20026 ( .B(clk), .A(\g.we_clk [12748]));
Q_ASSIGN U20027 ( .B(clk), .A(\g.we_clk [12747]));
Q_ASSIGN U20028 ( .B(clk), .A(\g.we_clk [12746]));
Q_ASSIGN U20029 ( .B(clk), .A(\g.we_clk [12745]));
Q_ASSIGN U20030 ( .B(clk), .A(\g.we_clk [12744]));
Q_ASSIGN U20031 ( .B(clk), .A(\g.we_clk [12743]));
Q_ASSIGN U20032 ( .B(clk), .A(\g.we_clk [12742]));
Q_ASSIGN U20033 ( .B(clk), .A(\g.we_clk [12741]));
Q_ASSIGN U20034 ( .B(clk), .A(\g.we_clk [12740]));
Q_ASSIGN U20035 ( .B(clk), .A(\g.we_clk [12739]));
Q_ASSIGN U20036 ( .B(clk), .A(\g.we_clk [12738]));
Q_ASSIGN U20037 ( .B(clk), .A(\g.we_clk [12737]));
Q_ASSIGN U20038 ( .B(clk), .A(\g.we_clk [12736]));
Q_ASSIGN U20039 ( .B(clk), .A(\g.we_clk [12735]));
Q_ASSIGN U20040 ( .B(clk), .A(\g.we_clk [12734]));
Q_ASSIGN U20041 ( .B(clk), .A(\g.we_clk [12733]));
Q_ASSIGN U20042 ( .B(clk), .A(\g.we_clk [12732]));
Q_ASSIGN U20043 ( .B(clk), .A(\g.we_clk [12731]));
Q_ASSIGN U20044 ( .B(clk), .A(\g.we_clk [12730]));
Q_ASSIGN U20045 ( .B(clk), .A(\g.we_clk [12729]));
Q_ASSIGN U20046 ( .B(clk), .A(\g.we_clk [12728]));
Q_ASSIGN U20047 ( .B(clk), .A(\g.we_clk [12727]));
Q_ASSIGN U20048 ( .B(clk), .A(\g.we_clk [12726]));
Q_ASSIGN U20049 ( .B(clk), .A(\g.we_clk [12725]));
Q_ASSIGN U20050 ( .B(clk), .A(\g.we_clk [12724]));
Q_ASSIGN U20051 ( .B(clk), .A(\g.we_clk [12723]));
Q_ASSIGN U20052 ( .B(clk), .A(\g.we_clk [12722]));
Q_ASSIGN U20053 ( .B(clk), .A(\g.we_clk [12721]));
Q_ASSIGN U20054 ( .B(clk), .A(\g.we_clk [12720]));
Q_ASSIGN U20055 ( .B(clk), .A(\g.we_clk [12719]));
Q_ASSIGN U20056 ( .B(clk), .A(\g.we_clk [12718]));
Q_ASSIGN U20057 ( .B(clk), .A(\g.we_clk [12717]));
Q_ASSIGN U20058 ( .B(clk), .A(\g.we_clk [12716]));
Q_ASSIGN U20059 ( .B(clk), .A(\g.we_clk [12715]));
Q_ASSIGN U20060 ( .B(clk), .A(\g.we_clk [12714]));
Q_ASSIGN U20061 ( .B(clk), .A(\g.we_clk [12713]));
Q_ASSIGN U20062 ( .B(clk), .A(\g.we_clk [12712]));
Q_ASSIGN U20063 ( .B(clk), .A(\g.we_clk [12711]));
Q_ASSIGN U20064 ( .B(clk), .A(\g.we_clk [12710]));
Q_ASSIGN U20065 ( .B(clk), .A(\g.we_clk [12709]));
Q_ASSIGN U20066 ( .B(clk), .A(\g.we_clk [12708]));
Q_ASSIGN U20067 ( .B(clk), .A(\g.we_clk [12707]));
Q_ASSIGN U20068 ( .B(clk), .A(\g.we_clk [12706]));
Q_ASSIGN U20069 ( .B(clk), .A(\g.we_clk [12705]));
Q_ASSIGN U20070 ( .B(clk), .A(\g.we_clk [12704]));
Q_ASSIGN U20071 ( .B(clk), .A(\g.we_clk [12703]));
Q_ASSIGN U20072 ( .B(clk), .A(\g.we_clk [12702]));
Q_ASSIGN U20073 ( .B(clk), .A(\g.we_clk [12701]));
Q_ASSIGN U20074 ( .B(clk), .A(\g.we_clk [12700]));
Q_ASSIGN U20075 ( .B(clk), .A(\g.we_clk [12699]));
Q_ASSIGN U20076 ( .B(clk), .A(\g.we_clk [12698]));
Q_ASSIGN U20077 ( .B(clk), .A(\g.we_clk [12697]));
Q_ASSIGN U20078 ( .B(clk), .A(\g.we_clk [12696]));
Q_ASSIGN U20079 ( .B(clk), .A(\g.we_clk [12695]));
Q_ASSIGN U20080 ( .B(clk), .A(\g.we_clk [12694]));
Q_ASSIGN U20081 ( .B(clk), .A(\g.we_clk [12693]));
Q_ASSIGN U20082 ( .B(clk), .A(\g.we_clk [12692]));
Q_ASSIGN U20083 ( .B(clk), .A(\g.we_clk [12691]));
Q_ASSIGN U20084 ( .B(clk), .A(\g.we_clk [12690]));
Q_ASSIGN U20085 ( .B(clk), .A(\g.we_clk [12689]));
Q_ASSIGN U20086 ( .B(clk), .A(\g.we_clk [12688]));
Q_ASSIGN U20087 ( .B(clk), .A(\g.we_clk [12687]));
Q_ASSIGN U20088 ( .B(clk), .A(\g.we_clk [12686]));
Q_ASSIGN U20089 ( .B(clk), .A(\g.we_clk [12685]));
Q_ASSIGN U20090 ( .B(clk), .A(\g.we_clk [12684]));
Q_ASSIGN U20091 ( .B(clk), .A(\g.we_clk [12683]));
Q_ASSIGN U20092 ( .B(clk), .A(\g.we_clk [12682]));
Q_ASSIGN U20093 ( .B(clk), .A(\g.we_clk [12681]));
Q_ASSIGN U20094 ( .B(clk), .A(\g.we_clk [12680]));
Q_ASSIGN U20095 ( .B(clk), .A(\g.we_clk [12679]));
Q_ASSIGN U20096 ( .B(clk), .A(\g.we_clk [12678]));
Q_ASSIGN U20097 ( .B(clk), .A(\g.we_clk [12677]));
Q_ASSIGN U20098 ( .B(clk), .A(\g.we_clk [12676]));
Q_ASSIGN U20099 ( .B(clk), .A(\g.we_clk [12675]));
Q_ASSIGN U20100 ( .B(clk), .A(\g.we_clk [12674]));
Q_ASSIGN U20101 ( .B(clk), .A(\g.we_clk [12673]));
Q_ASSIGN U20102 ( .B(clk), .A(\g.we_clk [12672]));
Q_ASSIGN U20103 ( .B(clk), .A(\g.we_clk [12671]));
Q_ASSIGN U20104 ( .B(clk), .A(\g.we_clk [12670]));
Q_ASSIGN U20105 ( .B(clk), .A(\g.we_clk [12669]));
Q_ASSIGN U20106 ( .B(clk), .A(\g.we_clk [12668]));
Q_ASSIGN U20107 ( .B(clk), .A(\g.we_clk [12667]));
Q_ASSIGN U20108 ( .B(clk), .A(\g.we_clk [12666]));
Q_ASSIGN U20109 ( .B(clk), .A(\g.we_clk [12665]));
Q_ASSIGN U20110 ( .B(clk), .A(\g.we_clk [12664]));
Q_ASSIGN U20111 ( .B(clk), .A(\g.we_clk [12663]));
Q_ASSIGN U20112 ( .B(clk), .A(\g.we_clk [12662]));
Q_ASSIGN U20113 ( .B(clk), .A(\g.we_clk [12661]));
Q_ASSIGN U20114 ( .B(clk), .A(\g.we_clk [12660]));
Q_ASSIGN U20115 ( .B(clk), .A(\g.we_clk [12659]));
Q_ASSIGN U20116 ( .B(clk), .A(\g.we_clk [12658]));
Q_ASSIGN U20117 ( .B(clk), .A(\g.we_clk [12657]));
Q_ASSIGN U20118 ( .B(clk), .A(\g.we_clk [12656]));
Q_ASSIGN U20119 ( .B(clk), .A(\g.we_clk [12655]));
Q_ASSIGN U20120 ( .B(clk), .A(\g.we_clk [12654]));
Q_ASSIGN U20121 ( .B(clk), .A(\g.we_clk [12653]));
Q_ASSIGN U20122 ( .B(clk), .A(\g.we_clk [12652]));
Q_ASSIGN U20123 ( .B(clk), .A(\g.we_clk [12651]));
Q_ASSIGN U20124 ( .B(clk), .A(\g.we_clk [12650]));
Q_ASSIGN U20125 ( .B(clk), .A(\g.we_clk [12649]));
Q_ASSIGN U20126 ( .B(clk), .A(\g.we_clk [12648]));
Q_ASSIGN U20127 ( .B(clk), .A(\g.we_clk [12647]));
Q_ASSIGN U20128 ( .B(clk), .A(\g.we_clk [12646]));
Q_ASSIGN U20129 ( .B(clk), .A(\g.we_clk [12645]));
Q_ASSIGN U20130 ( .B(clk), .A(\g.we_clk [12644]));
Q_ASSIGN U20131 ( .B(clk), .A(\g.we_clk [12643]));
Q_ASSIGN U20132 ( .B(clk), .A(\g.we_clk [12642]));
Q_ASSIGN U20133 ( .B(clk), .A(\g.we_clk [12641]));
Q_ASSIGN U20134 ( .B(clk), .A(\g.we_clk [12640]));
Q_ASSIGN U20135 ( .B(clk), .A(\g.we_clk [12639]));
Q_ASSIGN U20136 ( .B(clk), .A(\g.we_clk [12638]));
Q_ASSIGN U20137 ( .B(clk), .A(\g.we_clk [12637]));
Q_ASSIGN U20138 ( .B(clk), .A(\g.we_clk [12636]));
Q_ASSIGN U20139 ( .B(clk), .A(\g.we_clk [12635]));
Q_ASSIGN U20140 ( .B(clk), .A(\g.we_clk [12634]));
Q_ASSIGN U20141 ( .B(clk), .A(\g.we_clk [12633]));
Q_ASSIGN U20142 ( .B(clk), .A(\g.we_clk [12632]));
Q_ASSIGN U20143 ( .B(clk), .A(\g.we_clk [12631]));
Q_ASSIGN U20144 ( .B(clk), .A(\g.we_clk [12630]));
Q_ASSIGN U20145 ( .B(clk), .A(\g.we_clk [12629]));
Q_ASSIGN U20146 ( .B(clk), .A(\g.we_clk [12628]));
Q_ASSIGN U20147 ( .B(clk), .A(\g.we_clk [12627]));
Q_ASSIGN U20148 ( .B(clk), .A(\g.we_clk [12626]));
Q_ASSIGN U20149 ( .B(clk), .A(\g.we_clk [12625]));
Q_ASSIGN U20150 ( .B(clk), .A(\g.we_clk [12624]));
Q_ASSIGN U20151 ( .B(clk), .A(\g.we_clk [12623]));
Q_ASSIGN U20152 ( .B(clk), .A(\g.we_clk [12622]));
Q_ASSIGN U20153 ( .B(clk), .A(\g.we_clk [12621]));
Q_ASSIGN U20154 ( .B(clk), .A(\g.we_clk [12620]));
Q_ASSIGN U20155 ( .B(clk), .A(\g.we_clk [12619]));
Q_ASSIGN U20156 ( .B(clk), .A(\g.we_clk [12618]));
Q_ASSIGN U20157 ( .B(clk), .A(\g.we_clk [12617]));
Q_ASSIGN U20158 ( .B(clk), .A(\g.we_clk [12616]));
Q_ASSIGN U20159 ( .B(clk), .A(\g.we_clk [12615]));
Q_ASSIGN U20160 ( .B(clk), .A(\g.we_clk [12614]));
Q_ASSIGN U20161 ( .B(clk), .A(\g.we_clk [12613]));
Q_ASSIGN U20162 ( .B(clk), .A(\g.we_clk [12612]));
Q_ASSIGN U20163 ( .B(clk), .A(\g.we_clk [12611]));
Q_ASSIGN U20164 ( .B(clk), .A(\g.we_clk [12610]));
Q_ASSIGN U20165 ( .B(clk), .A(\g.we_clk [12609]));
Q_ASSIGN U20166 ( .B(clk), .A(\g.we_clk [12608]));
Q_ASSIGN U20167 ( .B(clk), .A(\g.we_clk [12607]));
Q_ASSIGN U20168 ( .B(clk), .A(\g.we_clk [12606]));
Q_ASSIGN U20169 ( .B(clk), .A(\g.we_clk [12605]));
Q_ASSIGN U20170 ( .B(clk), .A(\g.we_clk [12604]));
Q_ASSIGN U20171 ( .B(clk), .A(\g.we_clk [12603]));
Q_ASSIGN U20172 ( .B(clk), .A(\g.we_clk [12602]));
Q_ASSIGN U20173 ( .B(clk), .A(\g.we_clk [12601]));
Q_ASSIGN U20174 ( .B(clk), .A(\g.we_clk [12600]));
Q_ASSIGN U20175 ( .B(clk), .A(\g.we_clk [12599]));
Q_ASSIGN U20176 ( .B(clk), .A(\g.we_clk [12598]));
Q_ASSIGN U20177 ( .B(clk), .A(\g.we_clk [12597]));
Q_ASSIGN U20178 ( .B(clk), .A(\g.we_clk [12596]));
Q_ASSIGN U20179 ( .B(clk), .A(\g.we_clk [12595]));
Q_ASSIGN U20180 ( .B(clk), .A(\g.we_clk [12594]));
Q_ASSIGN U20181 ( .B(clk), .A(\g.we_clk [12593]));
Q_ASSIGN U20182 ( .B(clk), .A(\g.we_clk [12592]));
Q_ASSIGN U20183 ( .B(clk), .A(\g.we_clk [12591]));
Q_ASSIGN U20184 ( .B(clk), .A(\g.we_clk [12590]));
Q_ASSIGN U20185 ( .B(clk), .A(\g.we_clk [12589]));
Q_ASSIGN U20186 ( .B(clk), .A(\g.we_clk [12588]));
Q_ASSIGN U20187 ( .B(clk), .A(\g.we_clk [12587]));
Q_ASSIGN U20188 ( .B(clk), .A(\g.we_clk [12586]));
Q_ASSIGN U20189 ( .B(clk), .A(\g.we_clk [12585]));
Q_ASSIGN U20190 ( .B(clk), .A(\g.we_clk [12584]));
Q_ASSIGN U20191 ( .B(clk), .A(\g.we_clk [12583]));
Q_ASSIGN U20192 ( .B(clk), .A(\g.we_clk [12582]));
Q_ASSIGN U20193 ( .B(clk), .A(\g.we_clk [12581]));
Q_ASSIGN U20194 ( .B(clk), .A(\g.we_clk [12580]));
Q_ASSIGN U20195 ( .B(clk), .A(\g.we_clk [12579]));
Q_ASSIGN U20196 ( .B(clk), .A(\g.we_clk [12578]));
Q_ASSIGN U20197 ( .B(clk), .A(\g.we_clk [12577]));
Q_ASSIGN U20198 ( .B(clk), .A(\g.we_clk [12576]));
Q_ASSIGN U20199 ( .B(clk), .A(\g.we_clk [12575]));
Q_ASSIGN U20200 ( .B(clk), .A(\g.we_clk [12574]));
Q_ASSIGN U20201 ( .B(clk), .A(\g.we_clk [12573]));
Q_ASSIGN U20202 ( .B(clk), .A(\g.we_clk [12572]));
Q_ASSIGN U20203 ( .B(clk), .A(\g.we_clk [12571]));
Q_ASSIGN U20204 ( .B(clk), .A(\g.we_clk [12570]));
Q_ASSIGN U20205 ( .B(clk), .A(\g.we_clk [12569]));
Q_ASSIGN U20206 ( .B(clk), .A(\g.we_clk [12568]));
Q_ASSIGN U20207 ( .B(clk), .A(\g.we_clk [12567]));
Q_ASSIGN U20208 ( .B(clk), .A(\g.we_clk [12566]));
Q_ASSIGN U20209 ( .B(clk), .A(\g.we_clk [12565]));
Q_ASSIGN U20210 ( .B(clk), .A(\g.we_clk [12564]));
Q_ASSIGN U20211 ( .B(clk), .A(\g.we_clk [12563]));
Q_ASSIGN U20212 ( .B(clk), .A(\g.we_clk [12562]));
Q_ASSIGN U20213 ( .B(clk), .A(\g.we_clk [12561]));
Q_ASSIGN U20214 ( .B(clk), .A(\g.we_clk [12560]));
Q_ASSIGN U20215 ( .B(clk), .A(\g.we_clk [12559]));
Q_ASSIGN U20216 ( .B(clk), .A(\g.we_clk [12558]));
Q_ASSIGN U20217 ( .B(clk), .A(\g.we_clk [12557]));
Q_ASSIGN U20218 ( .B(clk), .A(\g.we_clk [12556]));
Q_ASSIGN U20219 ( .B(clk), .A(\g.we_clk [12555]));
Q_ASSIGN U20220 ( .B(clk), .A(\g.we_clk [12554]));
Q_ASSIGN U20221 ( .B(clk), .A(\g.we_clk [12553]));
Q_ASSIGN U20222 ( .B(clk), .A(\g.we_clk [12552]));
Q_ASSIGN U20223 ( .B(clk), .A(\g.we_clk [12551]));
Q_ASSIGN U20224 ( .B(clk), .A(\g.we_clk [12550]));
Q_ASSIGN U20225 ( .B(clk), .A(\g.we_clk [12549]));
Q_ASSIGN U20226 ( .B(clk), .A(\g.we_clk [12548]));
Q_ASSIGN U20227 ( .B(clk), .A(\g.we_clk [12547]));
Q_ASSIGN U20228 ( .B(clk), .A(\g.we_clk [12546]));
Q_ASSIGN U20229 ( .B(clk), .A(\g.we_clk [12545]));
Q_ASSIGN U20230 ( .B(clk), .A(\g.we_clk [12544]));
Q_ASSIGN U20231 ( .B(clk), .A(\g.we_clk [12543]));
Q_ASSIGN U20232 ( .B(clk), .A(\g.we_clk [12542]));
Q_ASSIGN U20233 ( .B(clk), .A(\g.we_clk [12541]));
Q_ASSIGN U20234 ( .B(clk), .A(\g.we_clk [12540]));
Q_ASSIGN U20235 ( .B(clk), .A(\g.we_clk [12539]));
Q_ASSIGN U20236 ( .B(clk), .A(\g.we_clk [12538]));
Q_ASSIGN U20237 ( .B(clk), .A(\g.we_clk [12537]));
Q_ASSIGN U20238 ( .B(clk), .A(\g.we_clk [12536]));
Q_ASSIGN U20239 ( .B(clk), .A(\g.we_clk [12535]));
Q_ASSIGN U20240 ( .B(clk), .A(\g.we_clk [12534]));
Q_ASSIGN U20241 ( .B(clk), .A(\g.we_clk [12533]));
Q_ASSIGN U20242 ( .B(clk), .A(\g.we_clk [12532]));
Q_ASSIGN U20243 ( .B(clk), .A(\g.we_clk [12531]));
Q_ASSIGN U20244 ( .B(clk), .A(\g.we_clk [12530]));
Q_ASSIGN U20245 ( .B(clk), .A(\g.we_clk [12529]));
Q_ASSIGN U20246 ( .B(clk), .A(\g.we_clk [12528]));
Q_ASSIGN U20247 ( .B(clk), .A(\g.we_clk [12527]));
Q_ASSIGN U20248 ( .B(clk), .A(\g.we_clk [12526]));
Q_ASSIGN U20249 ( .B(clk), .A(\g.we_clk [12525]));
Q_ASSIGN U20250 ( .B(clk), .A(\g.we_clk [12524]));
Q_ASSIGN U20251 ( .B(clk), .A(\g.we_clk [12523]));
Q_ASSIGN U20252 ( .B(clk), .A(\g.we_clk [12522]));
Q_ASSIGN U20253 ( .B(clk), .A(\g.we_clk [12521]));
Q_ASSIGN U20254 ( .B(clk), .A(\g.we_clk [12520]));
Q_ASSIGN U20255 ( .B(clk), .A(\g.we_clk [12519]));
Q_ASSIGN U20256 ( .B(clk), .A(\g.we_clk [12518]));
Q_ASSIGN U20257 ( .B(clk), .A(\g.we_clk [12517]));
Q_ASSIGN U20258 ( .B(clk), .A(\g.we_clk [12516]));
Q_ASSIGN U20259 ( .B(clk), .A(\g.we_clk [12515]));
Q_ASSIGN U20260 ( .B(clk), .A(\g.we_clk [12514]));
Q_ASSIGN U20261 ( .B(clk), .A(\g.we_clk [12513]));
Q_ASSIGN U20262 ( .B(clk), .A(\g.we_clk [12512]));
Q_ASSIGN U20263 ( .B(clk), .A(\g.we_clk [12511]));
Q_ASSIGN U20264 ( .B(clk), .A(\g.we_clk [12510]));
Q_ASSIGN U20265 ( .B(clk), .A(\g.we_clk [12509]));
Q_ASSIGN U20266 ( .B(clk), .A(\g.we_clk [12508]));
Q_ASSIGN U20267 ( .B(clk), .A(\g.we_clk [12507]));
Q_ASSIGN U20268 ( .B(clk), .A(\g.we_clk [12506]));
Q_ASSIGN U20269 ( .B(clk), .A(\g.we_clk [12505]));
Q_ASSIGN U20270 ( .B(clk), .A(\g.we_clk [12504]));
Q_ASSIGN U20271 ( .B(clk), .A(\g.we_clk [12503]));
Q_ASSIGN U20272 ( .B(clk), .A(\g.we_clk [12502]));
Q_ASSIGN U20273 ( .B(clk), .A(\g.we_clk [12501]));
Q_ASSIGN U20274 ( .B(clk), .A(\g.we_clk [12500]));
Q_ASSIGN U20275 ( .B(clk), .A(\g.we_clk [12499]));
Q_ASSIGN U20276 ( .B(clk), .A(\g.we_clk [12498]));
Q_ASSIGN U20277 ( .B(clk), .A(\g.we_clk [12497]));
Q_ASSIGN U20278 ( .B(clk), .A(\g.we_clk [12496]));
Q_ASSIGN U20279 ( .B(clk), .A(\g.we_clk [12495]));
Q_ASSIGN U20280 ( .B(clk), .A(\g.we_clk [12494]));
Q_ASSIGN U20281 ( .B(clk), .A(\g.we_clk [12493]));
Q_ASSIGN U20282 ( .B(clk), .A(\g.we_clk [12492]));
Q_ASSIGN U20283 ( .B(clk), .A(\g.we_clk [12491]));
Q_ASSIGN U20284 ( .B(clk), .A(\g.we_clk [12490]));
Q_ASSIGN U20285 ( .B(clk), .A(\g.we_clk [12489]));
Q_ASSIGN U20286 ( .B(clk), .A(\g.we_clk [12488]));
Q_ASSIGN U20287 ( .B(clk), .A(\g.we_clk [12487]));
Q_ASSIGN U20288 ( .B(clk), .A(\g.we_clk [12486]));
Q_ASSIGN U20289 ( .B(clk), .A(\g.we_clk [12485]));
Q_ASSIGN U20290 ( .B(clk), .A(\g.we_clk [12484]));
Q_ASSIGN U20291 ( .B(clk), .A(\g.we_clk [12483]));
Q_ASSIGN U20292 ( .B(clk), .A(\g.we_clk [12482]));
Q_ASSIGN U20293 ( .B(clk), .A(\g.we_clk [12481]));
Q_ASSIGN U20294 ( .B(clk), .A(\g.we_clk [12480]));
Q_ASSIGN U20295 ( .B(clk), .A(\g.we_clk [12479]));
Q_ASSIGN U20296 ( .B(clk), .A(\g.we_clk [12478]));
Q_ASSIGN U20297 ( .B(clk), .A(\g.we_clk [12477]));
Q_ASSIGN U20298 ( .B(clk), .A(\g.we_clk [12476]));
Q_ASSIGN U20299 ( .B(clk), .A(\g.we_clk [12475]));
Q_ASSIGN U20300 ( .B(clk), .A(\g.we_clk [12474]));
Q_ASSIGN U20301 ( .B(clk), .A(\g.we_clk [12473]));
Q_ASSIGN U20302 ( .B(clk), .A(\g.we_clk [12472]));
Q_ASSIGN U20303 ( .B(clk), .A(\g.we_clk [12471]));
Q_ASSIGN U20304 ( .B(clk), .A(\g.we_clk [12470]));
Q_ASSIGN U20305 ( .B(clk), .A(\g.we_clk [12469]));
Q_ASSIGN U20306 ( .B(clk), .A(\g.we_clk [12468]));
Q_ASSIGN U20307 ( .B(clk), .A(\g.we_clk [12467]));
Q_ASSIGN U20308 ( .B(clk), .A(\g.we_clk [12466]));
Q_ASSIGN U20309 ( .B(clk), .A(\g.we_clk [12465]));
Q_ASSIGN U20310 ( .B(clk), .A(\g.we_clk [12464]));
Q_ASSIGN U20311 ( .B(clk), .A(\g.we_clk [12463]));
Q_ASSIGN U20312 ( .B(clk), .A(\g.we_clk [12462]));
Q_ASSIGN U20313 ( .B(clk), .A(\g.we_clk [12461]));
Q_ASSIGN U20314 ( .B(clk), .A(\g.we_clk [12460]));
Q_ASSIGN U20315 ( .B(clk), .A(\g.we_clk [12459]));
Q_ASSIGN U20316 ( .B(clk), .A(\g.we_clk [12458]));
Q_ASSIGN U20317 ( .B(clk), .A(\g.we_clk [12457]));
Q_ASSIGN U20318 ( .B(clk), .A(\g.we_clk [12456]));
Q_ASSIGN U20319 ( .B(clk), .A(\g.we_clk [12455]));
Q_ASSIGN U20320 ( .B(clk), .A(\g.we_clk [12454]));
Q_ASSIGN U20321 ( .B(clk), .A(\g.we_clk [12453]));
Q_ASSIGN U20322 ( .B(clk), .A(\g.we_clk [12452]));
Q_ASSIGN U20323 ( .B(clk), .A(\g.we_clk [12451]));
Q_ASSIGN U20324 ( .B(clk), .A(\g.we_clk [12450]));
Q_ASSIGN U20325 ( .B(clk), .A(\g.we_clk [12449]));
Q_ASSIGN U20326 ( .B(clk), .A(\g.we_clk [12448]));
Q_ASSIGN U20327 ( .B(clk), .A(\g.we_clk [12447]));
Q_ASSIGN U20328 ( .B(clk), .A(\g.we_clk [12446]));
Q_ASSIGN U20329 ( .B(clk), .A(\g.we_clk [12445]));
Q_ASSIGN U20330 ( .B(clk), .A(\g.we_clk [12444]));
Q_ASSIGN U20331 ( .B(clk), .A(\g.we_clk [12443]));
Q_ASSIGN U20332 ( .B(clk), .A(\g.we_clk [12442]));
Q_ASSIGN U20333 ( .B(clk), .A(\g.we_clk [12441]));
Q_ASSIGN U20334 ( .B(clk), .A(\g.we_clk [12440]));
Q_ASSIGN U20335 ( .B(clk), .A(\g.we_clk [12439]));
Q_ASSIGN U20336 ( .B(clk), .A(\g.we_clk [12438]));
Q_ASSIGN U20337 ( .B(clk), .A(\g.we_clk [12437]));
Q_ASSIGN U20338 ( .B(clk), .A(\g.we_clk [12436]));
Q_ASSIGN U20339 ( .B(clk), .A(\g.we_clk [12435]));
Q_ASSIGN U20340 ( .B(clk), .A(\g.we_clk [12434]));
Q_ASSIGN U20341 ( .B(clk), .A(\g.we_clk [12433]));
Q_ASSIGN U20342 ( .B(clk), .A(\g.we_clk [12432]));
Q_ASSIGN U20343 ( .B(clk), .A(\g.we_clk [12431]));
Q_ASSIGN U20344 ( .B(clk), .A(\g.we_clk [12430]));
Q_ASSIGN U20345 ( .B(clk), .A(\g.we_clk [12429]));
Q_ASSIGN U20346 ( .B(clk), .A(\g.we_clk [12428]));
Q_ASSIGN U20347 ( .B(clk), .A(\g.we_clk [12427]));
Q_ASSIGN U20348 ( .B(clk), .A(\g.we_clk [12426]));
Q_ASSIGN U20349 ( .B(clk), .A(\g.we_clk [12425]));
Q_ASSIGN U20350 ( .B(clk), .A(\g.we_clk [12424]));
Q_ASSIGN U20351 ( .B(clk), .A(\g.we_clk [12423]));
Q_ASSIGN U20352 ( .B(clk), .A(\g.we_clk [12422]));
Q_ASSIGN U20353 ( .B(clk), .A(\g.we_clk [12421]));
Q_ASSIGN U20354 ( .B(clk), .A(\g.we_clk [12420]));
Q_ASSIGN U20355 ( .B(clk), .A(\g.we_clk [12419]));
Q_ASSIGN U20356 ( .B(clk), .A(\g.we_clk [12418]));
Q_ASSIGN U20357 ( .B(clk), .A(\g.we_clk [12417]));
Q_ASSIGN U20358 ( .B(clk), .A(\g.we_clk [12416]));
Q_ASSIGN U20359 ( .B(clk), .A(\g.we_clk [12415]));
Q_ASSIGN U20360 ( .B(clk), .A(\g.we_clk [12414]));
Q_ASSIGN U20361 ( .B(clk), .A(\g.we_clk [12413]));
Q_ASSIGN U20362 ( .B(clk), .A(\g.we_clk [12412]));
Q_ASSIGN U20363 ( .B(clk), .A(\g.we_clk [12411]));
Q_ASSIGN U20364 ( .B(clk), .A(\g.we_clk [12410]));
Q_ASSIGN U20365 ( .B(clk), .A(\g.we_clk [12409]));
Q_ASSIGN U20366 ( .B(clk), .A(\g.we_clk [12408]));
Q_ASSIGN U20367 ( .B(clk), .A(\g.we_clk [12407]));
Q_ASSIGN U20368 ( .B(clk), .A(\g.we_clk [12406]));
Q_ASSIGN U20369 ( .B(clk), .A(\g.we_clk [12405]));
Q_ASSIGN U20370 ( .B(clk), .A(\g.we_clk [12404]));
Q_ASSIGN U20371 ( .B(clk), .A(\g.we_clk [12403]));
Q_ASSIGN U20372 ( .B(clk), .A(\g.we_clk [12402]));
Q_ASSIGN U20373 ( .B(clk), .A(\g.we_clk [12401]));
Q_ASSIGN U20374 ( .B(clk), .A(\g.we_clk [12400]));
Q_ASSIGN U20375 ( .B(clk), .A(\g.we_clk [12399]));
Q_ASSIGN U20376 ( .B(clk), .A(\g.we_clk [12398]));
Q_ASSIGN U20377 ( .B(clk), .A(\g.we_clk [12397]));
Q_ASSIGN U20378 ( .B(clk), .A(\g.we_clk [12396]));
Q_ASSIGN U20379 ( .B(clk), .A(\g.we_clk [12395]));
Q_ASSIGN U20380 ( .B(clk), .A(\g.we_clk [12394]));
Q_ASSIGN U20381 ( .B(clk), .A(\g.we_clk [12393]));
Q_ASSIGN U20382 ( .B(clk), .A(\g.we_clk [12392]));
Q_ASSIGN U20383 ( .B(clk), .A(\g.we_clk [12391]));
Q_ASSIGN U20384 ( .B(clk), .A(\g.we_clk [12390]));
Q_ASSIGN U20385 ( .B(clk), .A(\g.we_clk [12389]));
Q_ASSIGN U20386 ( .B(clk), .A(\g.we_clk [12388]));
Q_ASSIGN U20387 ( .B(clk), .A(\g.we_clk [12387]));
Q_ASSIGN U20388 ( .B(clk), .A(\g.we_clk [12386]));
Q_ASSIGN U20389 ( .B(clk), .A(\g.we_clk [12385]));
Q_ASSIGN U20390 ( .B(clk), .A(\g.we_clk [12384]));
Q_ASSIGN U20391 ( .B(clk), .A(\g.we_clk [12383]));
Q_ASSIGN U20392 ( .B(clk), .A(\g.we_clk [12382]));
Q_ASSIGN U20393 ( .B(clk), .A(\g.we_clk [12381]));
Q_ASSIGN U20394 ( .B(clk), .A(\g.we_clk [12380]));
Q_ASSIGN U20395 ( .B(clk), .A(\g.we_clk [12379]));
Q_ASSIGN U20396 ( .B(clk), .A(\g.we_clk [12378]));
Q_ASSIGN U20397 ( .B(clk), .A(\g.we_clk [12377]));
Q_ASSIGN U20398 ( .B(clk), .A(\g.we_clk [12376]));
Q_ASSIGN U20399 ( .B(clk), .A(\g.we_clk [12375]));
Q_ASSIGN U20400 ( .B(clk), .A(\g.we_clk [12374]));
Q_ASSIGN U20401 ( .B(clk), .A(\g.we_clk [12373]));
Q_ASSIGN U20402 ( .B(clk), .A(\g.we_clk [12372]));
Q_ASSIGN U20403 ( .B(clk), .A(\g.we_clk [12371]));
Q_ASSIGN U20404 ( .B(clk), .A(\g.we_clk [12370]));
Q_ASSIGN U20405 ( .B(clk), .A(\g.we_clk [12369]));
Q_ASSIGN U20406 ( .B(clk), .A(\g.we_clk [12368]));
Q_ASSIGN U20407 ( .B(clk), .A(\g.we_clk [12367]));
Q_ASSIGN U20408 ( .B(clk), .A(\g.we_clk [12366]));
Q_ASSIGN U20409 ( .B(clk), .A(\g.we_clk [12365]));
Q_ASSIGN U20410 ( .B(clk), .A(\g.we_clk [12364]));
Q_ASSIGN U20411 ( .B(clk), .A(\g.we_clk [12363]));
Q_ASSIGN U20412 ( .B(clk), .A(\g.we_clk [12362]));
Q_ASSIGN U20413 ( .B(clk), .A(\g.we_clk [12361]));
Q_ASSIGN U20414 ( .B(clk), .A(\g.we_clk [12360]));
Q_ASSIGN U20415 ( .B(clk), .A(\g.we_clk [12359]));
Q_ASSIGN U20416 ( .B(clk), .A(\g.we_clk [12358]));
Q_ASSIGN U20417 ( .B(clk), .A(\g.we_clk [12357]));
Q_ASSIGN U20418 ( .B(clk), .A(\g.we_clk [12356]));
Q_ASSIGN U20419 ( .B(clk), .A(\g.we_clk [12355]));
Q_ASSIGN U20420 ( .B(clk), .A(\g.we_clk [12354]));
Q_ASSIGN U20421 ( .B(clk), .A(\g.we_clk [12353]));
Q_ASSIGN U20422 ( .B(clk), .A(\g.we_clk [12352]));
Q_ASSIGN U20423 ( .B(clk), .A(\g.we_clk [12351]));
Q_ASSIGN U20424 ( .B(clk), .A(\g.we_clk [12350]));
Q_ASSIGN U20425 ( .B(clk), .A(\g.we_clk [12349]));
Q_ASSIGN U20426 ( .B(clk), .A(\g.we_clk [12348]));
Q_ASSIGN U20427 ( .B(clk), .A(\g.we_clk [12347]));
Q_ASSIGN U20428 ( .B(clk), .A(\g.we_clk [12346]));
Q_ASSIGN U20429 ( .B(clk), .A(\g.we_clk [12345]));
Q_ASSIGN U20430 ( .B(clk), .A(\g.we_clk [12344]));
Q_ASSIGN U20431 ( .B(clk), .A(\g.we_clk [12343]));
Q_ASSIGN U20432 ( .B(clk), .A(\g.we_clk [12342]));
Q_ASSIGN U20433 ( .B(clk), .A(\g.we_clk [12341]));
Q_ASSIGN U20434 ( .B(clk), .A(\g.we_clk [12340]));
Q_ASSIGN U20435 ( .B(clk), .A(\g.we_clk [12339]));
Q_ASSIGN U20436 ( .B(clk), .A(\g.we_clk [12338]));
Q_ASSIGN U20437 ( .B(clk), .A(\g.we_clk [12337]));
Q_ASSIGN U20438 ( .B(clk), .A(\g.we_clk [12336]));
Q_ASSIGN U20439 ( .B(clk), .A(\g.we_clk [12335]));
Q_ASSIGN U20440 ( .B(clk), .A(\g.we_clk [12334]));
Q_ASSIGN U20441 ( .B(clk), .A(\g.we_clk [12333]));
Q_ASSIGN U20442 ( .B(clk), .A(\g.we_clk [12332]));
Q_ASSIGN U20443 ( .B(clk), .A(\g.we_clk [12331]));
Q_ASSIGN U20444 ( .B(clk), .A(\g.we_clk [12330]));
Q_ASSIGN U20445 ( .B(clk), .A(\g.we_clk [12329]));
Q_ASSIGN U20446 ( .B(clk), .A(\g.we_clk [12328]));
Q_ASSIGN U20447 ( .B(clk), .A(\g.we_clk [12327]));
Q_ASSIGN U20448 ( .B(clk), .A(\g.we_clk [12326]));
Q_ASSIGN U20449 ( .B(clk), .A(\g.we_clk [12325]));
Q_ASSIGN U20450 ( .B(clk), .A(\g.we_clk [12324]));
Q_ASSIGN U20451 ( .B(clk), .A(\g.we_clk [12323]));
Q_ASSIGN U20452 ( .B(clk), .A(\g.we_clk [12322]));
Q_ASSIGN U20453 ( .B(clk), .A(\g.we_clk [12321]));
Q_ASSIGN U20454 ( .B(clk), .A(\g.we_clk [12320]));
Q_ASSIGN U20455 ( .B(clk), .A(\g.we_clk [12319]));
Q_ASSIGN U20456 ( .B(clk), .A(\g.we_clk [12318]));
Q_ASSIGN U20457 ( .B(clk), .A(\g.we_clk [12317]));
Q_ASSIGN U20458 ( .B(clk), .A(\g.we_clk [12316]));
Q_ASSIGN U20459 ( .B(clk), .A(\g.we_clk [12315]));
Q_ASSIGN U20460 ( .B(clk), .A(\g.we_clk [12314]));
Q_ASSIGN U20461 ( .B(clk), .A(\g.we_clk [12313]));
Q_ASSIGN U20462 ( .B(clk), .A(\g.we_clk [12312]));
Q_ASSIGN U20463 ( .B(clk), .A(\g.we_clk [12311]));
Q_ASSIGN U20464 ( .B(clk), .A(\g.we_clk [12310]));
Q_ASSIGN U20465 ( .B(clk), .A(\g.we_clk [12309]));
Q_ASSIGN U20466 ( .B(clk), .A(\g.we_clk [12308]));
Q_ASSIGN U20467 ( .B(clk), .A(\g.we_clk [12307]));
Q_ASSIGN U20468 ( .B(clk), .A(\g.we_clk [12306]));
Q_ASSIGN U20469 ( .B(clk), .A(\g.we_clk [12305]));
Q_ASSIGN U20470 ( .B(clk), .A(\g.we_clk [12304]));
Q_ASSIGN U20471 ( .B(clk), .A(\g.we_clk [12303]));
Q_ASSIGN U20472 ( .B(clk), .A(\g.we_clk [12302]));
Q_ASSIGN U20473 ( .B(clk), .A(\g.we_clk [12301]));
Q_ASSIGN U20474 ( .B(clk), .A(\g.we_clk [12300]));
Q_ASSIGN U20475 ( .B(clk), .A(\g.we_clk [12299]));
Q_ASSIGN U20476 ( .B(clk), .A(\g.we_clk [12298]));
Q_ASSIGN U20477 ( .B(clk), .A(\g.we_clk [12297]));
Q_ASSIGN U20478 ( .B(clk), .A(\g.we_clk [12296]));
Q_ASSIGN U20479 ( .B(clk), .A(\g.we_clk [12295]));
Q_ASSIGN U20480 ( .B(clk), .A(\g.we_clk [12294]));
Q_ASSIGN U20481 ( .B(clk), .A(\g.we_clk [12293]));
Q_ASSIGN U20482 ( .B(clk), .A(\g.we_clk [12292]));
Q_ASSIGN U20483 ( .B(clk), .A(\g.we_clk [12291]));
Q_ASSIGN U20484 ( .B(clk), .A(\g.we_clk [12290]));
Q_ASSIGN U20485 ( .B(clk), .A(\g.we_clk [12289]));
Q_ASSIGN U20486 ( .B(clk), .A(\g.we_clk [12288]));
Q_ASSIGN U20487 ( .B(clk), .A(\g.we_clk [12287]));
Q_ASSIGN U20488 ( .B(clk), .A(\g.we_clk [12286]));
Q_ASSIGN U20489 ( .B(clk), .A(\g.we_clk [12285]));
Q_ASSIGN U20490 ( .B(clk), .A(\g.we_clk [12284]));
Q_ASSIGN U20491 ( .B(clk), .A(\g.we_clk [12283]));
Q_ASSIGN U20492 ( .B(clk), .A(\g.we_clk [12282]));
Q_ASSIGN U20493 ( .B(clk), .A(\g.we_clk [12281]));
Q_ASSIGN U20494 ( .B(clk), .A(\g.we_clk [12280]));
Q_ASSIGN U20495 ( .B(clk), .A(\g.we_clk [12279]));
Q_ASSIGN U20496 ( .B(clk), .A(\g.we_clk [12278]));
Q_ASSIGN U20497 ( .B(clk), .A(\g.we_clk [12277]));
Q_ASSIGN U20498 ( .B(clk), .A(\g.we_clk [12276]));
Q_ASSIGN U20499 ( .B(clk), .A(\g.we_clk [12275]));
Q_ASSIGN U20500 ( .B(clk), .A(\g.we_clk [12274]));
Q_ASSIGN U20501 ( .B(clk), .A(\g.we_clk [12273]));
Q_ASSIGN U20502 ( .B(clk), .A(\g.we_clk [12272]));
Q_ASSIGN U20503 ( .B(clk), .A(\g.we_clk [12271]));
Q_ASSIGN U20504 ( .B(clk), .A(\g.we_clk [12270]));
Q_ASSIGN U20505 ( .B(clk), .A(\g.we_clk [12269]));
Q_ASSIGN U20506 ( .B(clk), .A(\g.we_clk [12268]));
Q_ASSIGN U20507 ( .B(clk), .A(\g.we_clk [12267]));
Q_ASSIGN U20508 ( .B(clk), .A(\g.we_clk [12266]));
Q_ASSIGN U20509 ( .B(clk), .A(\g.we_clk [12265]));
Q_ASSIGN U20510 ( .B(clk), .A(\g.we_clk [12264]));
Q_ASSIGN U20511 ( .B(clk), .A(\g.we_clk [12263]));
Q_ASSIGN U20512 ( .B(clk), .A(\g.we_clk [12262]));
Q_ASSIGN U20513 ( .B(clk), .A(\g.we_clk [12261]));
Q_ASSIGN U20514 ( .B(clk), .A(\g.we_clk [12260]));
Q_ASSIGN U20515 ( .B(clk), .A(\g.we_clk [12259]));
Q_ASSIGN U20516 ( .B(clk), .A(\g.we_clk [12258]));
Q_ASSIGN U20517 ( .B(clk), .A(\g.we_clk [12257]));
Q_ASSIGN U20518 ( .B(clk), .A(\g.we_clk [12256]));
Q_ASSIGN U20519 ( .B(clk), .A(\g.we_clk [12255]));
Q_ASSIGN U20520 ( .B(clk), .A(\g.we_clk [12254]));
Q_ASSIGN U20521 ( .B(clk), .A(\g.we_clk [12253]));
Q_ASSIGN U20522 ( .B(clk), .A(\g.we_clk [12252]));
Q_ASSIGN U20523 ( .B(clk), .A(\g.we_clk [12251]));
Q_ASSIGN U20524 ( .B(clk), .A(\g.we_clk [12250]));
Q_ASSIGN U20525 ( .B(clk), .A(\g.we_clk [12249]));
Q_ASSIGN U20526 ( .B(clk), .A(\g.we_clk [12248]));
Q_ASSIGN U20527 ( .B(clk), .A(\g.we_clk [12247]));
Q_ASSIGN U20528 ( .B(clk), .A(\g.we_clk [12246]));
Q_ASSIGN U20529 ( .B(clk), .A(\g.we_clk [12245]));
Q_ASSIGN U20530 ( .B(clk), .A(\g.we_clk [12244]));
Q_ASSIGN U20531 ( .B(clk), .A(\g.we_clk [12243]));
Q_ASSIGN U20532 ( .B(clk), .A(\g.we_clk [12242]));
Q_ASSIGN U20533 ( .B(clk), .A(\g.we_clk [12241]));
Q_ASSIGN U20534 ( .B(clk), .A(\g.we_clk [12240]));
Q_ASSIGN U20535 ( .B(clk), .A(\g.we_clk [12239]));
Q_ASSIGN U20536 ( .B(clk), .A(\g.we_clk [12238]));
Q_ASSIGN U20537 ( .B(clk), .A(\g.we_clk [12237]));
Q_ASSIGN U20538 ( .B(clk), .A(\g.we_clk [12236]));
Q_ASSIGN U20539 ( .B(clk), .A(\g.we_clk [12235]));
Q_ASSIGN U20540 ( .B(clk), .A(\g.we_clk [12234]));
Q_ASSIGN U20541 ( .B(clk), .A(\g.we_clk [12233]));
Q_ASSIGN U20542 ( .B(clk), .A(\g.we_clk [12232]));
Q_ASSIGN U20543 ( .B(clk), .A(\g.we_clk [12231]));
Q_ASSIGN U20544 ( .B(clk), .A(\g.we_clk [12230]));
Q_ASSIGN U20545 ( .B(clk), .A(\g.we_clk [12229]));
Q_ASSIGN U20546 ( .B(clk), .A(\g.we_clk [12228]));
Q_ASSIGN U20547 ( .B(clk), .A(\g.we_clk [12227]));
Q_ASSIGN U20548 ( .B(clk), .A(\g.we_clk [12226]));
Q_ASSIGN U20549 ( .B(clk), .A(\g.we_clk [12225]));
Q_ASSIGN U20550 ( .B(clk), .A(\g.we_clk [12224]));
Q_ASSIGN U20551 ( .B(clk), .A(\g.we_clk [12223]));
Q_ASSIGN U20552 ( .B(clk), .A(\g.we_clk [12222]));
Q_ASSIGN U20553 ( .B(clk), .A(\g.we_clk [12221]));
Q_ASSIGN U20554 ( .B(clk), .A(\g.we_clk [12220]));
Q_ASSIGN U20555 ( .B(clk), .A(\g.we_clk [12219]));
Q_ASSIGN U20556 ( .B(clk), .A(\g.we_clk [12218]));
Q_ASSIGN U20557 ( .B(clk), .A(\g.we_clk [12217]));
Q_ASSIGN U20558 ( .B(clk), .A(\g.we_clk [12216]));
Q_ASSIGN U20559 ( .B(clk), .A(\g.we_clk [12215]));
Q_ASSIGN U20560 ( .B(clk), .A(\g.we_clk [12214]));
Q_ASSIGN U20561 ( .B(clk), .A(\g.we_clk [12213]));
Q_ASSIGN U20562 ( .B(clk), .A(\g.we_clk [12212]));
Q_ASSIGN U20563 ( .B(clk), .A(\g.we_clk [12211]));
Q_ASSIGN U20564 ( .B(clk), .A(\g.we_clk [12210]));
Q_ASSIGN U20565 ( .B(clk), .A(\g.we_clk [12209]));
Q_ASSIGN U20566 ( .B(clk), .A(\g.we_clk [12208]));
Q_ASSIGN U20567 ( .B(clk), .A(\g.we_clk [12207]));
Q_ASSIGN U20568 ( .B(clk), .A(\g.we_clk [12206]));
Q_ASSIGN U20569 ( .B(clk), .A(\g.we_clk [12205]));
Q_ASSIGN U20570 ( .B(clk), .A(\g.we_clk [12204]));
Q_ASSIGN U20571 ( .B(clk), .A(\g.we_clk [12203]));
Q_ASSIGN U20572 ( .B(clk), .A(\g.we_clk [12202]));
Q_ASSIGN U20573 ( .B(clk), .A(\g.we_clk [12201]));
Q_ASSIGN U20574 ( .B(clk), .A(\g.we_clk [12200]));
Q_ASSIGN U20575 ( .B(clk), .A(\g.we_clk [12199]));
Q_ASSIGN U20576 ( .B(clk), .A(\g.we_clk [12198]));
Q_ASSIGN U20577 ( .B(clk), .A(\g.we_clk [12197]));
Q_ASSIGN U20578 ( .B(clk), .A(\g.we_clk [12196]));
Q_ASSIGN U20579 ( .B(clk), .A(\g.we_clk [12195]));
Q_ASSIGN U20580 ( .B(clk), .A(\g.we_clk [12194]));
Q_ASSIGN U20581 ( .B(clk), .A(\g.we_clk [12193]));
Q_ASSIGN U20582 ( .B(clk), .A(\g.we_clk [12192]));
Q_ASSIGN U20583 ( .B(clk), .A(\g.we_clk [12191]));
Q_ASSIGN U20584 ( .B(clk), .A(\g.we_clk [12190]));
Q_ASSIGN U20585 ( .B(clk), .A(\g.we_clk [12189]));
Q_ASSIGN U20586 ( .B(clk), .A(\g.we_clk [12188]));
Q_ASSIGN U20587 ( .B(clk), .A(\g.we_clk [12187]));
Q_ASSIGN U20588 ( .B(clk), .A(\g.we_clk [12186]));
Q_ASSIGN U20589 ( .B(clk), .A(\g.we_clk [12185]));
Q_ASSIGN U20590 ( .B(clk), .A(\g.we_clk [12184]));
Q_ASSIGN U20591 ( .B(clk), .A(\g.we_clk [12183]));
Q_ASSIGN U20592 ( .B(clk), .A(\g.we_clk [12182]));
Q_ASSIGN U20593 ( .B(clk), .A(\g.we_clk [12181]));
Q_ASSIGN U20594 ( .B(clk), .A(\g.we_clk [12180]));
Q_ASSIGN U20595 ( .B(clk), .A(\g.we_clk [12179]));
Q_ASSIGN U20596 ( .B(clk), .A(\g.we_clk [12178]));
Q_ASSIGN U20597 ( .B(clk), .A(\g.we_clk [12177]));
Q_ASSIGN U20598 ( .B(clk), .A(\g.we_clk [12176]));
Q_ASSIGN U20599 ( .B(clk), .A(\g.we_clk [12175]));
Q_ASSIGN U20600 ( .B(clk), .A(\g.we_clk [12174]));
Q_ASSIGN U20601 ( .B(clk), .A(\g.we_clk [12173]));
Q_ASSIGN U20602 ( .B(clk), .A(\g.we_clk [12172]));
Q_ASSIGN U20603 ( .B(clk), .A(\g.we_clk [12171]));
Q_ASSIGN U20604 ( .B(clk), .A(\g.we_clk [12170]));
Q_ASSIGN U20605 ( .B(clk), .A(\g.we_clk [12169]));
Q_ASSIGN U20606 ( .B(clk), .A(\g.we_clk [12168]));
Q_ASSIGN U20607 ( .B(clk), .A(\g.we_clk [12167]));
Q_ASSIGN U20608 ( .B(clk), .A(\g.we_clk [12166]));
Q_ASSIGN U20609 ( .B(clk), .A(\g.we_clk [12165]));
Q_ASSIGN U20610 ( .B(clk), .A(\g.we_clk [12164]));
Q_ASSIGN U20611 ( .B(clk), .A(\g.we_clk [12163]));
Q_ASSIGN U20612 ( .B(clk), .A(\g.we_clk [12162]));
Q_ASSIGN U20613 ( .B(clk), .A(\g.we_clk [12161]));
Q_ASSIGN U20614 ( .B(clk), .A(\g.we_clk [12160]));
Q_ASSIGN U20615 ( .B(clk), .A(\g.we_clk [12159]));
Q_ASSIGN U20616 ( .B(clk), .A(\g.we_clk [12158]));
Q_ASSIGN U20617 ( .B(clk), .A(\g.we_clk [12157]));
Q_ASSIGN U20618 ( .B(clk), .A(\g.we_clk [12156]));
Q_ASSIGN U20619 ( .B(clk), .A(\g.we_clk [12155]));
Q_ASSIGN U20620 ( .B(clk), .A(\g.we_clk [12154]));
Q_ASSIGN U20621 ( .B(clk), .A(\g.we_clk [12153]));
Q_ASSIGN U20622 ( .B(clk), .A(\g.we_clk [12152]));
Q_ASSIGN U20623 ( .B(clk), .A(\g.we_clk [12151]));
Q_ASSIGN U20624 ( .B(clk), .A(\g.we_clk [12150]));
Q_ASSIGN U20625 ( .B(clk), .A(\g.we_clk [12149]));
Q_ASSIGN U20626 ( .B(clk), .A(\g.we_clk [12148]));
Q_ASSIGN U20627 ( .B(clk), .A(\g.we_clk [12147]));
Q_ASSIGN U20628 ( .B(clk), .A(\g.we_clk [12146]));
Q_ASSIGN U20629 ( .B(clk), .A(\g.we_clk [12145]));
Q_ASSIGN U20630 ( .B(clk), .A(\g.we_clk [12144]));
Q_ASSIGN U20631 ( .B(clk), .A(\g.we_clk [12143]));
Q_ASSIGN U20632 ( .B(clk), .A(\g.we_clk [12142]));
Q_ASSIGN U20633 ( .B(clk), .A(\g.we_clk [12141]));
Q_ASSIGN U20634 ( .B(clk), .A(\g.we_clk [12140]));
Q_ASSIGN U20635 ( .B(clk), .A(\g.we_clk [12139]));
Q_ASSIGN U20636 ( .B(clk), .A(\g.we_clk [12138]));
Q_ASSIGN U20637 ( .B(clk), .A(\g.we_clk [12137]));
Q_ASSIGN U20638 ( .B(clk), .A(\g.we_clk [12136]));
Q_ASSIGN U20639 ( .B(clk), .A(\g.we_clk [12135]));
Q_ASSIGN U20640 ( .B(clk), .A(\g.we_clk [12134]));
Q_ASSIGN U20641 ( .B(clk), .A(\g.we_clk [12133]));
Q_ASSIGN U20642 ( .B(clk), .A(\g.we_clk [12132]));
Q_ASSIGN U20643 ( .B(clk), .A(\g.we_clk [12131]));
Q_ASSIGN U20644 ( .B(clk), .A(\g.we_clk [12130]));
Q_ASSIGN U20645 ( .B(clk), .A(\g.we_clk [12129]));
Q_ASSIGN U20646 ( .B(clk), .A(\g.we_clk [12128]));
Q_ASSIGN U20647 ( .B(clk), .A(\g.we_clk [12127]));
Q_ASSIGN U20648 ( .B(clk), .A(\g.we_clk [12126]));
Q_ASSIGN U20649 ( .B(clk), .A(\g.we_clk [12125]));
Q_ASSIGN U20650 ( .B(clk), .A(\g.we_clk [12124]));
Q_ASSIGN U20651 ( .B(clk), .A(\g.we_clk [12123]));
Q_ASSIGN U20652 ( .B(clk), .A(\g.we_clk [12122]));
Q_ASSIGN U20653 ( .B(clk), .A(\g.we_clk [12121]));
Q_ASSIGN U20654 ( .B(clk), .A(\g.we_clk [12120]));
Q_ASSIGN U20655 ( .B(clk), .A(\g.we_clk [12119]));
Q_ASSIGN U20656 ( .B(clk), .A(\g.we_clk [12118]));
Q_ASSIGN U20657 ( .B(clk), .A(\g.we_clk [12117]));
Q_ASSIGN U20658 ( .B(clk), .A(\g.we_clk [12116]));
Q_ASSIGN U20659 ( .B(clk), .A(\g.we_clk [12115]));
Q_ASSIGN U20660 ( .B(clk), .A(\g.we_clk [12114]));
Q_ASSIGN U20661 ( .B(clk), .A(\g.we_clk [12113]));
Q_ASSIGN U20662 ( .B(clk), .A(\g.we_clk [12112]));
Q_ASSIGN U20663 ( .B(clk), .A(\g.we_clk [12111]));
Q_ASSIGN U20664 ( .B(clk), .A(\g.we_clk [12110]));
Q_ASSIGN U20665 ( .B(clk), .A(\g.we_clk [12109]));
Q_ASSIGN U20666 ( .B(clk), .A(\g.we_clk [12108]));
Q_ASSIGN U20667 ( .B(clk), .A(\g.we_clk [12107]));
Q_ASSIGN U20668 ( .B(clk), .A(\g.we_clk [12106]));
Q_ASSIGN U20669 ( .B(clk), .A(\g.we_clk [12105]));
Q_ASSIGN U20670 ( .B(clk), .A(\g.we_clk [12104]));
Q_ASSIGN U20671 ( .B(clk), .A(\g.we_clk [12103]));
Q_ASSIGN U20672 ( .B(clk), .A(\g.we_clk [12102]));
Q_ASSIGN U20673 ( .B(clk), .A(\g.we_clk [12101]));
Q_ASSIGN U20674 ( .B(clk), .A(\g.we_clk [12100]));
Q_ASSIGN U20675 ( .B(clk), .A(\g.we_clk [12099]));
Q_ASSIGN U20676 ( .B(clk), .A(\g.we_clk [12098]));
Q_ASSIGN U20677 ( .B(clk), .A(\g.we_clk [12097]));
Q_ASSIGN U20678 ( .B(clk), .A(\g.we_clk [12096]));
Q_ASSIGN U20679 ( .B(clk), .A(\g.we_clk [12095]));
Q_ASSIGN U20680 ( .B(clk), .A(\g.we_clk [12094]));
Q_ASSIGN U20681 ( .B(clk), .A(\g.we_clk [12093]));
Q_ASSIGN U20682 ( .B(clk), .A(\g.we_clk [12092]));
Q_ASSIGN U20683 ( .B(clk), .A(\g.we_clk [12091]));
Q_ASSIGN U20684 ( .B(clk), .A(\g.we_clk [12090]));
Q_ASSIGN U20685 ( .B(clk), .A(\g.we_clk [12089]));
Q_ASSIGN U20686 ( .B(clk), .A(\g.we_clk [12088]));
Q_ASSIGN U20687 ( .B(clk), .A(\g.we_clk [12087]));
Q_ASSIGN U20688 ( .B(clk), .A(\g.we_clk [12086]));
Q_ASSIGN U20689 ( .B(clk), .A(\g.we_clk [12085]));
Q_ASSIGN U20690 ( .B(clk), .A(\g.we_clk [12084]));
Q_ASSIGN U20691 ( .B(clk), .A(\g.we_clk [12083]));
Q_ASSIGN U20692 ( .B(clk), .A(\g.we_clk [12082]));
Q_ASSIGN U20693 ( .B(clk), .A(\g.we_clk [12081]));
Q_ASSIGN U20694 ( .B(clk), .A(\g.we_clk [12080]));
Q_ASSIGN U20695 ( .B(clk), .A(\g.we_clk [12079]));
Q_ASSIGN U20696 ( .B(clk), .A(\g.we_clk [12078]));
Q_ASSIGN U20697 ( .B(clk), .A(\g.we_clk [12077]));
Q_ASSIGN U20698 ( .B(clk), .A(\g.we_clk [12076]));
Q_ASSIGN U20699 ( .B(clk), .A(\g.we_clk [12075]));
Q_ASSIGN U20700 ( .B(clk), .A(\g.we_clk [12074]));
Q_ASSIGN U20701 ( .B(clk), .A(\g.we_clk [12073]));
Q_ASSIGN U20702 ( .B(clk), .A(\g.we_clk [12072]));
Q_ASSIGN U20703 ( .B(clk), .A(\g.we_clk [12071]));
Q_ASSIGN U20704 ( .B(clk), .A(\g.we_clk [12070]));
Q_ASSIGN U20705 ( .B(clk), .A(\g.we_clk [12069]));
Q_ASSIGN U20706 ( .B(clk), .A(\g.we_clk [12068]));
Q_ASSIGN U20707 ( .B(clk), .A(\g.we_clk [12067]));
Q_ASSIGN U20708 ( .B(clk), .A(\g.we_clk [12066]));
Q_ASSIGN U20709 ( .B(clk), .A(\g.we_clk [12065]));
Q_ASSIGN U20710 ( .B(clk), .A(\g.we_clk [12064]));
Q_ASSIGN U20711 ( .B(clk), .A(\g.we_clk [12063]));
Q_ASSIGN U20712 ( .B(clk), .A(\g.we_clk [12062]));
Q_ASSIGN U20713 ( .B(clk), .A(\g.we_clk [12061]));
Q_ASSIGN U20714 ( .B(clk), .A(\g.we_clk [12060]));
Q_ASSIGN U20715 ( .B(clk), .A(\g.we_clk [12059]));
Q_ASSIGN U20716 ( .B(clk), .A(\g.we_clk [12058]));
Q_ASSIGN U20717 ( .B(clk), .A(\g.we_clk [12057]));
Q_ASSIGN U20718 ( .B(clk), .A(\g.we_clk [12056]));
Q_ASSIGN U20719 ( .B(clk), .A(\g.we_clk [12055]));
Q_ASSIGN U20720 ( .B(clk), .A(\g.we_clk [12054]));
Q_ASSIGN U20721 ( .B(clk), .A(\g.we_clk [12053]));
Q_ASSIGN U20722 ( .B(clk), .A(\g.we_clk [12052]));
Q_ASSIGN U20723 ( .B(clk), .A(\g.we_clk [12051]));
Q_ASSIGN U20724 ( .B(clk), .A(\g.we_clk [12050]));
Q_ASSIGN U20725 ( .B(clk), .A(\g.we_clk [12049]));
Q_ASSIGN U20726 ( .B(clk), .A(\g.we_clk [12048]));
Q_ASSIGN U20727 ( .B(clk), .A(\g.we_clk [12047]));
Q_ASSIGN U20728 ( .B(clk), .A(\g.we_clk [12046]));
Q_ASSIGN U20729 ( .B(clk), .A(\g.we_clk [12045]));
Q_ASSIGN U20730 ( .B(clk), .A(\g.we_clk [12044]));
Q_ASSIGN U20731 ( .B(clk), .A(\g.we_clk [12043]));
Q_ASSIGN U20732 ( .B(clk), .A(\g.we_clk [12042]));
Q_ASSIGN U20733 ( .B(clk), .A(\g.we_clk [12041]));
Q_ASSIGN U20734 ( .B(clk), .A(\g.we_clk [12040]));
Q_ASSIGN U20735 ( .B(clk), .A(\g.we_clk [12039]));
Q_ASSIGN U20736 ( .B(clk), .A(\g.we_clk [12038]));
Q_ASSIGN U20737 ( .B(clk), .A(\g.we_clk [12037]));
Q_ASSIGN U20738 ( .B(clk), .A(\g.we_clk [12036]));
Q_ASSIGN U20739 ( .B(clk), .A(\g.we_clk [12035]));
Q_ASSIGN U20740 ( .B(clk), .A(\g.we_clk [12034]));
Q_ASSIGN U20741 ( .B(clk), .A(\g.we_clk [12033]));
Q_ASSIGN U20742 ( .B(clk), .A(\g.we_clk [12032]));
Q_ASSIGN U20743 ( .B(clk), .A(\g.we_clk [12031]));
Q_ASSIGN U20744 ( .B(clk), .A(\g.we_clk [12030]));
Q_ASSIGN U20745 ( .B(clk), .A(\g.we_clk [12029]));
Q_ASSIGN U20746 ( .B(clk), .A(\g.we_clk [12028]));
Q_ASSIGN U20747 ( .B(clk), .A(\g.we_clk [12027]));
Q_ASSIGN U20748 ( .B(clk), .A(\g.we_clk [12026]));
Q_ASSIGN U20749 ( .B(clk), .A(\g.we_clk [12025]));
Q_ASSIGN U20750 ( .B(clk), .A(\g.we_clk [12024]));
Q_ASSIGN U20751 ( .B(clk), .A(\g.we_clk [12023]));
Q_ASSIGN U20752 ( .B(clk), .A(\g.we_clk [12022]));
Q_ASSIGN U20753 ( .B(clk), .A(\g.we_clk [12021]));
Q_ASSIGN U20754 ( .B(clk), .A(\g.we_clk [12020]));
Q_ASSIGN U20755 ( .B(clk), .A(\g.we_clk [12019]));
Q_ASSIGN U20756 ( .B(clk), .A(\g.we_clk [12018]));
Q_ASSIGN U20757 ( .B(clk), .A(\g.we_clk [12017]));
Q_ASSIGN U20758 ( .B(clk), .A(\g.we_clk [12016]));
Q_ASSIGN U20759 ( .B(clk), .A(\g.we_clk [12015]));
Q_ASSIGN U20760 ( .B(clk), .A(\g.we_clk [12014]));
Q_ASSIGN U20761 ( .B(clk), .A(\g.we_clk [12013]));
Q_ASSIGN U20762 ( .B(clk), .A(\g.we_clk [12012]));
Q_ASSIGN U20763 ( .B(clk), .A(\g.we_clk [12011]));
Q_ASSIGN U20764 ( .B(clk), .A(\g.we_clk [12010]));
Q_ASSIGN U20765 ( .B(clk), .A(\g.we_clk [12009]));
Q_ASSIGN U20766 ( .B(clk), .A(\g.we_clk [12008]));
Q_ASSIGN U20767 ( .B(clk), .A(\g.we_clk [12007]));
Q_ASSIGN U20768 ( .B(clk), .A(\g.we_clk [12006]));
Q_ASSIGN U20769 ( .B(clk), .A(\g.we_clk [12005]));
Q_ASSIGN U20770 ( .B(clk), .A(\g.we_clk [12004]));
Q_ASSIGN U20771 ( .B(clk), .A(\g.we_clk [12003]));
Q_ASSIGN U20772 ( .B(clk), .A(\g.we_clk [12002]));
Q_ASSIGN U20773 ( .B(clk), .A(\g.we_clk [12001]));
Q_ASSIGN U20774 ( .B(clk), .A(\g.we_clk [12000]));
Q_ASSIGN U20775 ( .B(clk), .A(\g.we_clk [11999]));
Q_ASSIGN U20776 ( .B(clk), .A(\g.we_clk [11998]));
Q_ASSIGN U20777 ( .B(clk), .A(\g.we_clk [11997]));
Q_ASSIGN U20778 ( .B(clk), .A(\g.we_clk [11996]));
Q_ASSIGN U20779 ( .B(clk), .A(\g.we_clk [11995]));
Q_ASSIGN U20780 ( .B(clk), .A(\g.we_clk [11994]));
Q_ASSIGN U20781 ( .B(clk), .A(\g.we_clk [11993]));
Q_ASSIGN U20782 ( .B(clk), .A(\g.we_clk [11992]));
Q_ASSIGN U20783 ( .B(clk), .A(\g.we_clk [11991]));
Q_ASSIGN U20784 ( .B(clk), .A(\g.we_clk [11990]));
Q_ASSIGN U20785 ( .B(clk), .A(\g.we_clk [11989]));
Q_ASSIGN U20786 ( .B(clk), .A(\g.we_clk [11988]));
Q_ASSIGN U20787 ( .B(clk), .A(\g.we_clk [11987]));
Q_ASSIGN U20788 ( .B(clk), .A(\g.we_clk [11986]));
Q_ASSIGN U20789 ( .B(clk), .A(\g.we_clk [11985]));
Q_ASSIGN U20790 ( .B(clk), .A(\g.we_clk [11984]));
Q_ASSIGN U20791 ( .B(clk), .A(\g.we_clk [11983]));
Q_ASSIGN U20792 ( .B(clk), .A(\g.we_clk [11982]));
Q_ASSIGN U20793 ( .B(clk), .A(\g.we_clk [11981]));
Q_ASSIGN U20794 ( .B(clk), .A(\g.we_clk [11980]));
Q_ASSIGN U20795 ( .B(clk), .A(\g.we_clk [11979]));
Q_ASSIGN U20796 ( .B(clk), .A(\g.we_clk [11978]));
Q_ASSIGN U20797 ( .B(clk), .A(\g.we_clk [11977]));
Q_ASSIGN U20798 ( .B(clk), .A(\g.we_clk [11976]));
Q_ASSIGN U20799 ( .B(clk), .A(\g.we_clk [11975]));
Q_ASSIGN U20800 ( .B(clk), .A(\g.we_clk [11974]));
Q_ASSIGN U20801 ( .B(clk), .A(\g.we_clk [11973]));
Q_ASSIGN U20802 ( .B(clk), .A(\g.we_clk [11972]));
Q_ASSIGN U20803 ( .B(clk), .A(\g.we_clk [11971]));
Q_ASSIGN U20804 ( .B(clk), .A(\g.we_clk [11970]));
Q_ASSIGN U20805 ( .B(clk), .A(\g.we_clk [11969]));
Q_ASSIGN U20806 ( .B(clk), .A(\g.we_clk [11968]));
Q_ASSIGN U20807 ( .B(clk), .A(\g.we_clk [11967]));
Q_ASSIGN U20808 ( .B(clk), .A(\g.we_clk [11966]));
Q_ASSIGN U20809 ( .B(clk), .A(\g.we_clk [11965]));
Q_ASSIGN U20810 ( .B(clk), .A(\g.we_clk [11964]));
Q_ASSIGN U20811 ( .B(clk), .A(\g.we_clk [11963]));
Q_ASSIGN U20812 ( .B(clk), .A(\g.we_clk [11962]));
Q_ASSIGN U20813 ( .B(clk), .A(\g.we_clk [11961]));
Q_ASSIGN U20814 ( .B(clk), .A(\g.we_clk [11960]));
Q_ASSIGN U20815 ( .B(clk), .A(\g.we_clk [11959]));
Q_ASSIGN U20816 ( .B(clk), .A(\g.we_clk [11958]));
Q_ASSIGN U20817 ( .B(clk), .A(\g.we_clk [11957]));
Q_ASSIGN U20818 ( .B(clk), .A(\g.we_clk [11956]));
Q_ASSIGN U20819 ( .B(clk), .A(\g.we_clk [11955]));
Q_ASSIGN U20820 ( .B(clk), .A(\g.we_clk [11954]));
Q_ASSIGN U20821 ( .B(clk), .A(\g.we_clk [11953]));
Q_ASSIGN U20822 ( .B(clk), .A(\g.we_clk [11952]));
Q_ASSIGN U20823 ( .B(clk), .A(\g.we_clk [11951]));
Q_ASSIGN U20824 ( .B(clk), .A(\g.we_clk [11950]));
Q_ASSIGN U20825 ( .B(clk), .A(\g.we_clk [11949]));
Q_ASSIGN U20826 ( .B(clk), .A(\g.we_clk [11948]));
Q_ASSIGN U20827 ( .B(clk), .A(\g.we_clk [11947]));
Q_ASSIGN U20828 ( .B(clk), .A(\g.we_clk [11946]));
Q_ASSIGN U20829 ( .B(clk), .A(\g.we_clk [11945]));
Q_ASSIGN U20830 ( .B(clk), .A(\g.we_clk [11944]));
Q_ASSIGN U20831 ( .B(clk), .A(\g.we_clk [11943]));
Q_ASSIGN U20832 ( .B(clk), .A(\g.we_clk [11942]));
Q_ASSIGN U20833 ( .B(clk), .A(\g.we_clk [11941]));
Q_ASSIGN U20834 ( .B(clk), .A(\g.we_clk [11940]));
Q_ASSIGN U20835 ( .B(clk), .A(\g.we_clk [11939]));
Q_ASSIGN U20836 ( .B(clk), .A(\g.we_clk [11938]));
Q_ASSIGN U20837 ( .B(clk), .A(\g.we_clk [11937]));
Q_ASSIGN U20838 ( .B(clk), .A(\g.we_clk [11936]));
Q_ASSIGN U20839 ( .B(clk), .A(\g.we_clk [11935]));
Q_ASSIGN U20840 ( .B(clk), .A(\g.we_clk [11934]));
Q_ASSIGN U20841 ( .B(clk), .A(\g.we_clk [11933]));
Q_ASSIGN U20842 ( .B(clk), .A(\g.we_clk [11932]));
Q_ASSIGN U20843 ( .B(clk), .A(\g.we_clk [11931]));
Q_ASSIGN U20844 ( .B(clk), .A(\g.we_clk [11930]));
Q_ASSIGN U20845 ( .B(clk), .A(\g.we_clk [11929]));
Q_ASSIGN U20846 ( .B(clk), .A(\g.we_clk [11928]));
Q_ASSIGN U20847 ( .B(clk), .A(\g.we_clk [11927]));
Q_ASSIGN U20848 ( .B(clk), .A(\g.we_clk [11926]));
Q_ASSIGN U20849 ( .B(clk), .A(\g.we_clk [11925]));
Q_ASSIGN U20850 ( .B(clk), .A(\g.we_clk [11924]));
Q_ASSIGN U20851 ( .B(clk), .A(\g.we_clk [11923]));
Q_ASSIGN U20852 ( .B(clk), .A(\g.we_clk [11922]));
Q_ASSIGN U20853 ( .B(clk), .A(\g.we_clk [11921]));
Q_ASSIGN U20854 ( .B(clk), .A(\g.we_clk [11920]));
Q_ASSIGN U20855 ( .B(clk), .A(\g.we_clk [11919]));
Q_ASSIGN U20856 ( .B(clk), .A(\g.we_clk [11918]));
Q_ASSIGN U20857 ( .B(clk), .A(\g.we_clk [11917]));
Q_ASSIGN U20858 ( .B(clk), .A(\g.we_clk [11916]));
Q_ASSIGN U20859 ( .B(clk), .A(\g.we_clk [11915]));
Q_ASSIGN U20860 ( .B(clk), .A(\g.we_clk [11914]));
Q_ASSIGN U20861 ( .B(clk), .A(\g.we_clk [11913]));
Q_ASSIGN U20862 ( .B(clk), .A(\g.we_clk [11912]));
Q_ASSIGN U20863 ( .B(clk), .A(\g.we_clk [11911]));
Q_ASSIGN U20864 ( .B(clk), .A(\g.we_clk [11910]));
Q_ASSIGN U20865 ( .B(clk), .A(\g.we_clk [11909]));
Q_ASSIGN U20866 ( .B(clk), .A(\g.we_clk [11908]));
Q_ASSIGN U20867 ( .B(clk), .A(\g.we_clk [11907]));
Q_ASSIGN U20868 ( .B(clk), .A(\g.we_clk [11906]));
Q_ASSIGN U20869 ( .B(clk), .A(\g.we_clk [11905]));
Q_ASSIGN U20870 ( .B(clk), .A(\g.we_clk [11904]));
Q_ASSIGN U20871 ( .B(clk), .A(\g.we_clk [11903]));
Q_ASSIGN U20872 ( .B(clk), .A(\g.we_clk [11902]));
Q_ASSIGN U20873 ( .B(clk), .A(\g.we_clk [11901]));
Q_ASSIGN U20874 ( .B(clk), .A(\g.we_clk [11900]));
Q_ASSIGN U20875 ( .B(clk), .A(\g.we_clk [11899]));
Q_ASSIGN U20876 ( .B(clk), .A(\g.we_clk [11898]));
Q_ASSIGN U20877 ( .B(clk), .A(\g.we_clk [11897]));
Q_ASSIGN U20878 ( .B(clk), .A(\g.we_clk [11896]));
Q_ASSIGN U20879 ( .B(clk), .A(\g.we_clk [11895]));
Q_ASSIGN U20880 ( .B(clk), .A(\g.we_clk [11894]));
Q_ASSIGN U20881 ( .B(clk), .A(\g.we_clk [11893]));
Q_ASSIGN U20882 ( .B(clk), .A(\g.we_clk [11892]));
Q_ASSIGN U20883 ( .B(clk), .A(\g.we_clk [11891]));
Q_ASSIGN U20884 ( .B(clk), .A(\g.we_clk [11890]));
Q_ASSIGN U20885 ( .B(clk), .A(\g.we_clk [11889]));
Q_ASSIGN U20886 ( .B(clk), .A(\g.we_clk [11888]));
Q_ASSIGN U20887 ( .B(clk), .A(\g.we_clk [11887]));
Q_ASSIGN U20888 ( .B(clk), .A(\g.we_clk [11886]));
Q_ASSIGN U20889 ( .B(clk), .A(\g.we_clk [11885]));
Q_ASSIGN U20890 ( .B(clk), .A(\g.we_clk [11884]));
Q_ASSIGN U20891 ( .B(clk), .A(\g.we_clk [11883]));
Q_ASSIGN U20892 ( .B(clk), .A(\g.we_clk [11882]));
Q_ASSIGN U20893 ( .B(clk), .A(\g.we_clk [11881]));
Q_ASSIGN U20894 ( .B(clk), .A(\g.we_clk [11880]));
Q_ASSIGN U20895 ( .B(clk), .A(\g.we_clk [11879]));
Q_ASSIGN U20896 ( .B(clk), .A(\g.we_clk [11878]));
Q_ASSIGN U20897 ( .B(clk), .A(\g.we_clk [11877]));
Q_ASSIGN U20898 ( .B(clk), .A(\g.we_clk [11876]));
Q_ASSIGN U20899 ( .B(clk), .A(\g.we_clk [11875]));
Q_ASSIGN U20900 ( .B(clk), .A(\g.we_clk [11874]));
Q_ASSIGN U20901 ( .B(clk), .A(\g.we_clk [11873]));
Q_ASSIGN U20902 ( .B(clk), .A(\g.we_clk [11872]));
Q_ASSIGN U20903 ( .B(clk), .A(\g.we_clk [11871]));
Q_ASSIGN U20904 ( .B(clk), .A(\g.we_clk [11870]));
Q_ASSIGN U20905 ( .B(clk), .A(\g.we_clk [11869]));
Q_ASSIGN U20906 ( .B(clk), .A(\g.we_clk [11868]));
Q_ASSIGN U20907 ( .B(clk), .A(\g.we_clk [11867]));
Q_ASSIGN U20908 ( .B(clk), .A(\g.we_clk [11866]));
Q_ASSIGN U20909 ( .B(clk), .A(\g.we_clk [11865]));
Q_ASSIGN U20910 ( .B(clk), .A(\g.we_clk [11864]));
Q_ASSIGN U20911 ( .B(clk), .A(\g.we_clk [11863]));
Q_ASSIGN U20912 ( .B(clk), .A(\g.we_clk [11862]));
Q_ASSIGN U20913 ( .B(clk), .A(\g.we_clk [11861]));
Q_ASSIGN U20914 ( .B(clk), .A(\g.we_clk [11860]));
Q_ASSIGN U20915 ( .B(clk), .A(\g.we_clk [11859]));
Q_ASSIGN U20916 ( .B(clk), .A(\g.we_clk [11858]));
Q_ASSIGN U20917 ( .B(clk), .A(\g.we_clk [11857]));
Q_ASSIGN U20918 ( .B(clk), .A(\g.we_clk [11856]));
Q_ASSIGN U20919 ( .B(clk), .A(\g.we_clk [11855]));
Q_ASSIGN U20920 ( .B(clk), .A(\g.we_clk [11854]));
Q_ASSIGN U20921 ( .B(clk), .A(\g.we_clk [11853]));
Q_ASSIGN U20922 ( .B(clk), .A(\g.we_clk [11852]));
Q_ASSIGN U20923 ( .B(clk), .A(\g.we_clk [11851]));
Q_ASSIGN U20924 ( .B(clk), .A(\g.we_clk [11850]));
Q_ASSIGN U20925 ( .B(clk), .A(\g.we_clk [11849]));
Q_ASSIGN U20926 ( .B(clk), .A(\g.we_clk [11848]));
Q_ASSIGN U20927 ( .B(clk), .A(\g.we_clk [11847]));
Q_ASSIGN U20928 ( .B(clk), .A(\g.we_clk [11846]));
Q_ASSIGN U20929 ( .B(clk), .A(\g.we_clk [11845]));
Q_ASSIGN U20930 ( .B(clk), .A(\g.we_clk [11844]));
Q_ASSIGN U20931 ( .B(clk), .A(\g.we_clk [11843]));
Q_ASSIGN U20932 ( .B(clk), .A(\g.we_clk [11842]));
Q_ASSIGN U20933 ( .B(clk), .A(\g.we_clk [11841]));
Q_ASSIGN U20934 ( .B(clk), .A(\g.we_clk [11840]));
Q_ASSIGN U20935 ( .B(clk), .A(\g.we_clk [11839]));
Q_ASSIGN U20936 ( .B(clk), .A(\g.we_clk [11838]));
Q_ASSIGN U20937 ( .B(clk), .A(\g.we_clk [11837]));
Q_ASSIGN U20938 ( .B(clk), .A(\g.we_clk [11836]));
Q_ASSIGN U20939 ( .B(clk), .A(\g.we_clk [11835]));
Q_ASSIGN U20940 ( .B(clk), .A(\g.we_clk [11834]));
Q_ASSIGN U20941 ( .B(clk), .A(\g.we_clk [11833]));
Q_ASSIGN U20942 ( .B(clk), .A(\g.we_clk [11832]));
Q_ASSIGN U20943 ( .B(clk), .A(\g.we_clk [11831]));
Q_ASSIGN U20944 ( .B(clk), .A(\g.we_clk [11830]));
Q_ASSIGN U20945 ( .B(clk), .A(\g.we_clk [11829]));
Q_ASSIGN U20946 ( .B(clk), .A(\g.we_clk [11828]));
Q_ASSIGN U20947 ( .B(clk), .A(\g.we_clk [11827]));
Q_ASSIGN U20948 ( .B(clk), .A(\g.we_clk [11826]));
Q_ASSIGN U20949 ( .B(clk), .A(\g.we_clk [11825]));
Q_ASSIGN U20950 ( .B(clk), .A(\g.we_clk [11824]));
Q_ASSIGN U20951 ( .B(clk), .A(\g.we_clk [11823]));
Q_ASSIGN U20952 ( .B(clk), .A(\g.we_clk [11822]));
Q_ASSIGN U20953 ( .B(clk), .A(\g.we_clk [11821]));
Q_ASSIGN U20954 ( .B(clk), .A(\g.we_clk [11820]));
Q_ASSIGN U20955 ( .B(clk), .A(\g.we_clk [11819]));
Q_ASSIGN U20956 ( .B(clk), .A(\g.we_clk [11818]));
Q_ASSIGN U20957 ( .B(clk), .A(\g.we_clk [11817]));
Q_ASSIGN U20958 ( .B(clk), .A(\g.we_clk [11816]));
Q_ASSIGN U20959 ( .B(clk), .A(\g.we_clk [11815]));
Q_ASSIGN U20960 ( .B(clk), .A(\g.we_clk [11814]));
Q_ASSIGN U20961 ( .B(clk), .A(\g.we_clk [11813]));
Q_ASSIGN U20962 ( .B(clk), .A(\g.we_clk [11812]));
Q_ASSIGN U20963 ( .B(clk), .A(\g.we_clk [11811]));
Q_ASSIGN U20964 ( .B(clk), .A(\g.we_clk [11810]));
Q_ASSIGN U20965 ( .B(clk), .A(\g.we_clk [11809]));
Q_ASSIGN U20966 ( .B(clk), .A(\g.we_clk [11808]));
Q_ASSIGN U20967 ( .B(clk), .A(\g.we_clk [11807]));
Q_ASSIGN U20968 ( .B(clk), .A(\g.we_clk [11806]));
Q_ASSIGN U20969 ( .B(clk), .A(\g.we_clk [11805]));
Q_ASSIGN U20970 ( .B(clk), .A(\g.we_clk [11804]));
Q_ASSIGN U20971 ( .B(clk), .A(\g.we_clk [11803]));
Q_ASSIGN U20972 ( .B(clk), .A(\g.we_clk [11802]));
Q_ASSIGN U20973 ( .B(clk), .A(\g.we_clk [11801]));
Q_ASSIGN U20974 ( .B(clk), .A(\g.we_clk [11800]));
Q_ASSIGN U20975 ( .B(clk), .A(\g.we_clk [11799]));
Q_ASSIGN U20976 ( .B(clk), .A(\g.we_clk [11798]));
Q_ASSIGN U20977 ( .B(clk), .A(\g.we_clk [11797]));
Q_ASSIGN U20978 ( .B(clk), .A(\g.we_clk [11796]));
Q_ASSIGN U20979 ( .B(clk), .A(\g.we_clk [11795]));
Q_ASSIGN U20980 ( .B(clk), .A(\g.we_clk [11794]));
Q_ASSIGN U20981 ( .B(clk), .A(\g.we_clk [11793]));
Q_ASSIGN U20982 ( .B(clk), .A(\g.we_clk [11792]));
Q_ASSIGN U20983 ( .B(clk), .A(\g.we_clk [11791]));
Q_ASSIGN U20984 ( .B(clk), .A(\g.we_clk [11790]));
Q_ASSIGN U20985 ( .B(clk), .A(\g.we_clk [11789]));
Q_ASSIGN U20986 ( .B(clk), .A(\g.we_clk [11788]));
Q_ASSIGN U20987 ( .B(clk), .A(\g.we_clk [11787]));
Q_ASSIGN U20988 ( .B(clk), .A(\g.we_clk [11786]));
Q_ASSIGN U20989 ( .B(clk), .A(\g.we_clk [11785]));
Q_ASSIGN U20990 ( .B(clk), .A(\g.we_clk [11784]));
Q_ASSIGN U20991 ( .B(clk), .A(\g.we_clk [11783]));
Q_ASSIGN U20992 ( .B(clk), .A(\g.we_clk [11782]));
Q_ASSIGN U20993 ( .B(clk), .A(\g.we_clk [11781]));
Q_ASSIGN U20994 ( .B(clk), .A(\g.we_clk [11780]));
Q_ASSIGN U20995 ( .B(clk), .A(\g.we_clk [11779]));
Q_ASSIGN U20996 ( .B(clk), .A(\g.we_clk [11778]));
Q_ASSIGN U20997 ( .B(clk), .A(\g.we_clk [11777]));
Q_ASSIGN U20998 ( .B(clk), .A(\g.we_clk [11776]));
Q_ASSIGN U20999 ( .B(clk), .A(\g.we_clk [11775]));
Q_ASSIGN U21000 ( .B(clk), .A(\g.we_clk [11774]));
Q_ASSIGN U21001 ( .B(clk), .A(\g.we_clk [11773]));
Q_ASSIGN U21002 ( .B(clk), .A(\g.we_clk [11772]));
Q_ASSIGN U21003 ( .B(clk), .A(\g.we_clk [11771]));
Q_ASSIGN U21004 ( .B(clk), .A(\g.we_clk [11770]));
Q_ASSIGN U21005 ( .B(clk), .A(\g.we_clk [11769]));
Q_ASSIGN U21006 ( .B(clk), .A(\g.we_clk [11768]));
Q_ASSIGN U21007 ( .B(clk), .A(\g.we_clk [11767]));
Q_ASSIGN U21008 ( .B(clk), .A(\g.we_clk [11766]));
Q_ASSIGN U21009 ( .B(clk), .A(\g.we_clk [11765]));
Q_ASSIGN U21010 ( .B(clk), .A(\g.we_clk [11764]));
Q_ASSIGN U21011 ( .B(clk), .A(\g.we_clk [11763]));
Q_ASSIGN U21012 ( .B(clk), .A(\g.we_clk [11762]));
Q_ASSIGN U21013 ( .B(clk), .A(\g.we_clk [11761]));
Q_ASSIGN U21014 ( .B(clk), .A(\g.we_clk [11760]));
Q_ASSIGN U21015 ( .B(clk), .A(\g.we_clk [11759]));
Q_ASSIGN U21016 ( .B(clk), .A(\g.we_clk [11758]));
Q_ASSIGN U21017 ( .B(clk), .A(\g.we_clk [11757]));
Q_ASSIGN U21018 ( .B(clk), .A(\g.we_clk [11756]));
Q_ASSIGN U21019 ( .B(clk), .A(\g.we_clk [11755]));
Q_ASSIGN U21020 ( .B(clk), .A(\g.we_clk [11754]));
Q_ASSIGN U21021 ( .B(clk), .A(\g.we_clk [11753]));
Q_ASSIGN U21022 ( .B(clk), .A(\g.we_clk [11752]));
Q_ASSIGN U21023 ( .B(clk), .A(\g.we_clk [11751]));
Q_ASSIGN U21024 ( .B(clk), .A(\g.we_clk [11750]));
Q_ASSIGN U21025 ( .B(clk), .A(\g.we_clk [11749]));
Q_ASSIGN U21026 ( .B(clk), .A(\g.we_clk [11748]));
Q_ASSIGN U21027 ( .B(clk), .A(\g.we_clk [11747]));
Q_ASSIGN U21028 ( .B(clk), .A(\g.we_clk [11746]));
Q_ASSIGN U21029 ( .B(clk), .A(\g.we_clk [11745]));
Q_ASSIGN U21030 ( .B(clk), .A(\g.we_clk [11744]));
Q_ASSIGN U21031 ( .B(clk), .A(\g.we_clk [11743]));
Q_ASSIGN U21032 ( .B(clk), .A(\g.we_clk [11742]));
Q_ASSIGN U21033 ( .B(clk), .A(\g.we_clk [11741]));
Q_ASSIGN U21034 ( .B(clk), .A(\g.we_clk [11740]));
Q_ASSIGN U21035 ( .B(clk), .A(\g.we_clk [11739]));
Q_ASSIGN U21036 ( .B(clk), .A(\g.we_clk [11738]));
Q_ASSIGN U21037 ( .B(clk), .A(\g.we_clk [11737]));
Q_ASSIGN U21038 ( .B(clk), .A(\g.we_clk [11736]));
Q_ASSIGN U21039 ( .B(clk), .A(\g.we_clk [11735]));
Q_ASSIGN U21040 ( .B(clk), .A(\g.we_clk [11734]));
Q_ASSIGN U21041 ( .B(clk), .A(\g.we_clk [11733]));
Q_ASSIGN U21042 ( .B(clk), .A(\g.we_clk [11732]));
Q_ASSIGN U21043 ( .B(clk), .A(\g.we_clk [11731]));
Q_ASSIGN U21044 ( .B(clk), .A(\g.we_clk [11730]));
Q_ASSIGN U21045 ( .B(clk), .A(\g.we_clk [11729]));
Q_ASSIGN U21046 ( .B(clk), .A(\g.we_clk [11728]));
Q_ASSIGN U21047 ( .B(clk), .A(\g.we_clk [11727]));
Q_ASSIGN U21048 ( .B(clk), .A(\g.we_clk [11726]));
Q_ASSIGN U21049 ( .B(clk), .A(\g.we_clk [11725]));
Q_ASSIGN U21050 ( .B(clk), .A(\g.we_clk [11724]));
Q_ASSIGN U21051 ( .B(clk), .A(\g.we_clk [11723]));
Q_ASSIGN U21052 ( .B(clk), .A(\g.we_clk [11722]));
Q_ASSIGN U21053 ( .B(clk), .A(\g.we_clk [11721]));
Q_ASSIGN U21054 ( .B(clk), .A(\g.we_clk [11720]));
Q_ASSIGN U21055 ( .B(clk), .A(\g.we_clk [11719]));
Q_ASSIGN U21056 ( .B(clk), .A(\g.we_clk [11718]));
Q_ASSIGN U21057 ( .B(clk), .A(\g.we_clk [11717]));
Q_ASSIGN U21058 ( .B(clk), .A(\g.we_clk [11716]));
Q_ASSIGN U21059 ( .B(clk), .A(\g.we_clk [11715]));
Q_ASSIGN U21060 ( .B(clk), .A(\g.we_clk [11714]));
Q_ASSIGN U21061 ( .B(clk), .A(\g.we_clk [11713]));
Q_ASSIGN U21062 ( .B(clk), .A(\g.we_clk [11712]));
Q_ASSIGN U21063 ( .B(clk), .A(\g.we_clk [11711]));
Q_ASSIGN U21064 ( .B(clk), .A(\g.we_clk [11710]));
Q_ASSIGN U21065 ( .B(clk), .A(\g.we_clk [11709]));
Q_ASSIGN U21066 ( .B(clk), .A(\g.we_clk [11708]));
Q_ASSIGN U21067 ( .B(clk), .A(\g.we_clk [11707]));
Q_ASSIGN U21068 ( .B(clk), .A(\g.we_clk [11706]));
Q_ASSIGN U21069 ( .B(clk), .A(\g.we_clk [11705]));
Q_ASSIGN U21070 ( .B(clk), .A(\g.we_clk [11704]));
Q_ASSIGN U21071 ( .B(clk), .A(\g.we_clk [11703]));
Q_ASSIGN U21072 ( .B(clk), .A(\g.we_clk [11702]));
Q_ASSIGN U21073 ( .B(clk), .A(\g.we_clk [11701]));
Q_ASSIGN U21074 ( .B(clk), .A(\g.we_clk [11700]));
Q_ASSIGN U21075 ( .B(clk), .A(\g.we_clk [11699]));
Q_ASSIGN U21076 ( .B(clk), .A(\g.we_clk [11698]));
Q_ASSIGN U21077 ( .B(clk), .A(\g.we_clk [11697]));
Q_ASSIGN U21078 ( .B(clk), .A(\g.we_clk [11696]));
Q_ASSIGN U21079 ( .B(clk), .A(\g.we_clk [11695]));
Q_ASSIGN U21080 ( .B(clk), .A(\g.we_clk [11694]));
Q_ASSIGN U21081 ( .B(clk), .A(\g.we_clk [11693]));
Q_ASSIGN U21082 ( .B(clk), .A(\g.we_clk [11692]));
Q_ASSIGN U21083 ( .B(clk), .A(\g.we_clk [11691]));
Q_ASSIGN U21084 ( .B(clk), .A(\g.we_clk [11690]));
Q_ASSIGN U21085 ( .B(clk), .A(\g.we_clk [11689]));
Q_ASSIGN U21086 ( .B(clk), .A(\g.we_clk [11688]));
Q_ASSIGN U21087 ( .B(clk), .A(\g.we_clk [11687]));
Q_ASSIGN U21088 ( .B(clk), .A(\g.we_clk [11686]));
Q_ASSIGN U21089 ( .B(clk), .A(\g.we_clk [11685]));
Q_ASSIGN U21090 ( .B(clk), .A(\g.we_clk [11684]));
Q_ASSIGN U21091 ( .B(clk), .A(\g.we_clk [11683]));
Q_ASSIGN U21092 ( .B(clk), .A(\g.we_clk [11682]));
Q_ASSIGN U21093 ( .B(clk), .A(\g.we_clk [11681]));
Q_ASSIGN U21094 ( .B(clk), .A(\g.we_clk [11680]));
Q_ASSIGN U21095 ( .B(clk), .A(\g.we_clk [11679]));
Q_ASSIGN U21096 ( .B(clk), .A(\g.we_clk [11678]));
Q_ASSIGN U21097 ( .B(clk), .A(\g.we_clk [11677]));
Q_ASSIGN U21098 ( .B(clk), .A(\g.we_clk [11676]));
Q_ASSIGN U21099 ( .B(clk), .A(\g.we_clk [11675]));
Q_ASSIGN U21100 ( .B(clk), .A(\g.we_clk [11674]));
Q_ASSIGN U21101 ( .B(clk), .A(\g.we_clk [11673]));
Q_ASSIGN U21102 ( .B(clk), .A(\g.we_clk [11672]));
Q_ASSIGN U21103 ( .B(clk), .A(\g.we_clk [11671]));
Q_ASSIGN U21104 ( .B(clk), .A(\g.we_clk [11670]));
Q_ASSIGN U21105 ( .B(clk), .A(\g.we_clk [11669]));
Q_ASSIGN U21106 ( .B(clk), .A(\g.we_clk [11668]));
Q_ASSIGN U21107 ( .B(clk), .A(\g.we_clk [11667]));
Q_ASSIGN U21108 ( .B(clk), .A(\g.we_clk [11666]));
Q_ASSIGN U21109 ( .B(clk), .A(\g.we_clk [11665]));
Q_ASSIGN U21110 ( .B(clk), .A(\g.we_clk [11664]));
Q_ASSIGN U21111 ( .B(clk), .A(\g.we_clk [11663]));
Q_ASSIGN U21112 ( .B(clk), .A(\g.we_clk [11662]));
Q_ASSIGN U21113 ( .B(clk), .A(\g.we_clk [11661]));
Q_ASSIGN U21114 ( .B(clk), .A(\g.we_clk [11660]));
Q_ASSIGN U21115 ( .B(clk), .A(\g.we_clk [11659]));
Q_ASSIGN U21116 ( .B(clk), .A(\g.we_clk [11658]));
Q_ASSIGN U21117 ( .B(clk), .A(\g.we_clk [11657]));
Q_ASSIGN U21118 ( .B(clk), .A(\g.we_clk [11656]));
Q_ASSIGN U21119 ( .B(clk), .A(\g.we_clk [11655]));
Q_ASSIGN U21120 ( .B(clk), .A(\g.we_clk [11654]));
Q_ASSIGN U21121 ( .B(clk), .A(\g.we_clk [11653]));
Q_ASSIGN U21122 ( .B(clk), .A(\g.we_clk [11652]));
Q_ASSIGN U21123 ( .B(clk), .A(\g.we_clk [11651]));
Q_ASSIGN U21124 ( .B(clk), .A(\g.we_clk [11650]));
Q_ASSIGN U21125 ( .B(clk), .A(\g.we_clk [11649]));
Q_ASSIGN U21126 ( .B(clk), .A(\g.we_clk [11648]));
Q_ASSIGN U21127 ( .B(clk), .A(\g.we_clk [11647]));
Q_ASSIGN U21128 ( .B(clk), .A(\g.we_clk [11646]));
Q_ASSIGN U21129 ( .B(clk), .A(\g.we_clk [11645]));
Q_ASSIGN U21130 ( .B(clk), .A(\g.we_clk [11644]));
Q_ASSIGN U21131 ( .B(clk), .A(\g.we_clk [11643]));
Q_ASSIGN U21132 ( .B(clk), .A(\g.we_clk [11642]));
Q_ASSIGN U21133 ( .B(clk), .A(\g.we_clk [11641]));
Q_ASSIGN U21134 ( .B(clk), .A(\g.we_clk [11640]));
Q_ASSIGN U21135 ( .B(clk), .A(\g.we_clk [11639]));
Q_ASSIGN U21136 ( .B(clk), .A(\g.we_clk [11638]));
Q_ASSIGN U21137 ( .B(clk), .A(\g.we_clk [11637]));
Q_ASSIGN U21138 ( .B(clk), .A(\g.we_clk [11636]));
Q_ASSIGN U21139 ( .B(clk), .A(\g.we_clk [11635]));
Q_ASSIGN U21140 ( .B(clk), .A(\g.we_clk [11634]));
Q_ASSIGN U21141 ( .B(clk), .A(\g.we_clk [11633]));
Q_ASSIGN U21142 ( .B(clk), .A(\g.we_clk [11632]));
Q_ASSIGN U21143 ( .B(clk), .A(\g.we_clk [11631]));
Q_ASSIGN U21144 ( .B(clk), .A(\g.we_clk [11630]));
Q_ASSIGN U21145 ( .B(clk), .A(\g.we_clk [11629]));
Q_ASSIGN U21146 ( .B(clk), .A(\g.we_clk [11628]));
Q_ASSIGN U21147 ( .B(clk), .A(\g.we_clk [11627]));
Q_ASSIGN U21148 ( .B(clk), .A(\g.we_clk [11626]));
Q_ASSIGN U21149 ( .B(clk), .A(\g.we_clk [11625]));
Q_ASSIGN U21150 ( .B(clk), .A(\g.we_clk [11624]));
Q_ASSIGN U21151 ( .B(clk), .A(\g.we_clk [11623]));
Q_ASSIGN U21152 ( .B(clk), .A(\g.we_clk [11622]));
Q_ASSIGN U21153 ( .B(clk), .A(\g.we_clk [11621]));
Q_ASSIGN U21154 ( .B(clk), .A(\g.we_clk [11620]));
Q_ASSIGN U21155 ( .B(clk), .A(\g.we_clk [11619]));
Q_ASSIGN U21156 ( .B(clk), .A(\g.we_clk [11618]));
Q_ASSIGN U21157 ( .B(clk), .A(\g.we_clk [11617]));
Q_ASSIGN U21158 ( .B(clk), .A(\g.we_clk [11616]));
Q_ASSIGN U21159 ( .B(clk), .A(\g.we_clk [11615]));
Q_ASSIGN U21160 ( .B(clk), .A(\g.we_clk [11614]));
Q_ASSIGN U21161 ( .B(clk), .A(\g.we_clk [11613]));
Q_ASSIGN U21162 ( .B(clk), .A(\g.we_clk [11612]));
Q_ASSIGN U21163 ( .B(clk), .A(\g.we_clk [11611]));
Q_ASSIGN U21164 ( .B(clk), .A(\g.we_clk [11610]));
Q_ASSIGN U21165 ( .B(clk), .A(\g.we_clk [11609]));
Q_ASSIGN U21166 ( .B(clk), .A(\g.we_clk [11608]));
Q_ASSIGN U21167 ( .B(clk), .A(\g.we_clk [11607]));
Q_ASSIGN U21168 ( .B(clk), .A(\g.we_clk [11606]));
Q_ASSIGN U21169 ( .B(clk), .A(\g.we_clk [11605]));
Q_ASSIGN U21170 ( .B(clk), .A(\g.we_clk [11604]));
Q_ASSIGN U21171 ( .B(clk), .A(\g.we_clk [11603]));
Q_ASSIGN U21172 ( .B(clk), .A(\g.we_clk [11602]));
Q_ASSIGN U21173 ( .B(clk), .A(\g.we_clk [11601]));
Q_ASSIGN U21174 ( .B(clk), .A(\g.we_clk [11600]));
Q_ASSIGN U21175 ( .B(clk), .A(\g.we_clk [11599]));
Q_ASSIGN U21176 ( .B(clk), .A(\g.we_clk [11598]));
Q_ASSIGN U21177 ( .B(clk), .A(\g.we_clk [11597]));
Q_ASSIGN U21178 ( .B(clk), .A(\g.we_clk [11596]));
Q_ASSIGN U21179 ( .B(clk), .A(\g.we_clk [11595]));
Q_ASSIGN U21180 ( .B(clk), .A(\g.we_clk [11594]));
Q_ASSIGN U21181 ( .B(clk), .A(\g.we_clk [11593]));
Q_ASSIGN U21182 ( .B(clk), .A(\g.we_clk [11592]));
Q_ASSIGN U21183 ( .B(clk), .A(\g.we_clk [11591]));
Q_ASSIGN U21184 ( .B(clk), .A(\g.we_clk [11590]));
Q_ASSIGN U21185 ( .B(clk), .A(\g.we_clk [11589]));
Q_ASSIGN U21186 ( .B(clk), .A(\g.we_clk [11588]));
Q_ASSIGN U21187 ( .B(clk), .A(\g.we_clk [11587]));
Q_ASSIGN U21188 ( .B(clk), .A(\g.we_clk [11586]));
Q_ASSIGN U21189 ( .B(clk), .A(\g.we_clk [11585]));
Q_ASSIGN U21190 ( .B(clk), .A(\g.we_clk [11584]));
Q_ASSIGN U21191 ( .B(clk), .A(\g.we_clk [11583]));
Q_ASSIGN U21192 ( .B(clk), .A(\g.we_clk [11582]));
Q_ASSIGN U21193 ( .B(clk), .A(\g.we_clk [11581]));
Q_ASSIGN U21194 ( .B(clk), .A(\g.we_clk [11580]));
Q_ASSIGN U21195 ( .B(clk), .A(\g.we_clk [11579]));
Q_ASSIGN U21196 ( .B(clk), .A(\g.we_clk [11578]));
Q_ASSIGN U21197 ( .B(clk), .A(\g.we_clk [11577]));
Q_ASSIGN U21198 ( .B(clk), .A(\g.we_clk [11576]));
Q_ASSIGN U21199 ( .B(clk), .A(\g.we_clk [11575]));
Q_ASSIGN U21200 ( .B(clk), .A(\g.we_clk [11574]));
Q_ASSIGN U21201 ( .B(clk), .A(\g.we_clk [11573]));
Q_ASSIGN U21202 ( .B(clk), .A(\g.we_clk [11572]));
Q_ASSIGN U21203 ( .B(clk), .A(\g.we_clk [11571]));
Q_ASSIGN U21204 ( .B(clk), .A(\g.we_clk [11570]));
Q_ASSIGN U21205 ( .B(clk), .A(\g.we_clk [11569]));
Q_ASSIGN U21206 ( .B(clk), .A(\g.we_clk [11568]));
Q_ASSIGN U21207 ( .B(clk), .A(\g.we_clk [11567]));
Q_ASSIGN U21208 ( .B(clk), .A(\g.we_clk [11566]));
Q_ASSIGN U21209 ( .B(clk), .A(\g.we_clk [11565]));
Q_ASSIGN U21210 ( .B(clk), .A(\g.we_clk [11564]));
Q_ASSIGN U21211 ( .B(clk), .A(\g.we_clk [11563]));
Q_ASSIGN U21212 ( .B(clk), .A(\g.we_clk [11562]));
Q_ASSIGN U21213 ( .B(clk), .A(\g.we_clk [11561]));
Q_ASSIGN U21214 ( .B(clk), .A(\g.we_clk [11560]));
Q_ASSIGN U21215 ( .B(clk), .A(\g.we_clk [11559]));
Q_ASSIGN U21216 ( .B(clk), .A(\g.we_clk [11558]));
Q_ASSIGN U21217 ( .B(clk), .A(\g.we_clk [11557]));
Q_ASSIGN U21218 ( .B(clk), .A(\g.we_clk [11556]));
Q_ASSIGN U21219 ( .B(clk), .A(\g.we_clk [11555]));
Q_ASSIGN U21220 ( .B(clk), .A(\g.we_clk [11554]));
Q_ASSIGN U21221 ( .B(clk), .A(\g.we_clk [11553]));
Q_ASSIGN U21222 ( .B(clk), .A(\g.we_clk [11552]));
Q_ASSIGN U21223 ( .B(clk), .A(\g.we_clk [11551]));
Q_ASSIGN U21224 ( .B(clk), .A(\g.we_clk [11550]));
Q_ASSIGN U21225 ( .B(clk), .A(\g.we_clk [11549]));
Q_ASSIGN U21226 ( .B(clk), .A(\g.we_clk [11548]));
Q_ASSIGN U21227 ( .B(clk), .A(\g.we_clk [11547]));
Q_ASSIGN U21228 ( .B(clk), .A(\g.we_clk [11546]));
Q_ASSIGN U21229 ( .B(clk), .A(\g.we_clk [11545]));
Q_ASSIGN U21230 ( .B(clk), .A(\g.we_clk [11544]));
Q_ASSIGN U21231 ( .B(clk), .A(\g.we_clk [11543]));
Q_ASSIGN U21232 ( .B(clk), .A(\g.we_clk [11542]));
Q_ASSIGN U21233 ( .B(clk), .A(\g.we_clk [11541]));
Q_ASSIGN U21234 ( .B(clk), .A(\g.we_clk [11540]));
Q_ASSIGN U21235 ( .B(clk), .A(\g.we_clk [11539]));
Q_ASSIGN U21236 ( .B(clk), .A(\g.we_clk [11538]));
Q_ASSIGN U21237 ( .B(clk), .A(\g.we_clk [11537]));
Q_ASSIGN U21238 ( .B(clk), .A(\g.we_clk [11536]));
Q_ASSIGN U21239 ( .B(clk), .A(\g.we_clk [11535]));
Q_ASSIGN U21240 ( .B(clk), .A(\g.we_clk [11534]));
Q_ASSIGN U21241 ( .B(clk), .A(\g.we_clk [11533]));
Q_ASSIGN U21242 ( .B(clk), .A(\g.we_clk [11532]));
Q_ASSIGN U21243 ( .B(clk), .A(\g.we_clk [11531]));
Q_ASSIGN U21244 ( .B(clk), .A(\g.we_clk [11530]));
Q_ASSIGN U21245 ( .B(clk), .A(\g.we_clk [11529]));
Q_ASSIGN U21246 ( .B(clk), .A(\g.we_clk [11528]));
Q_ASSIGN U21247 ( .B(clk), .A(\g.we_clk [11527]));
Q_ASSIGN U21248 ( .B(clk), .A(\g.we_clk [11526]));
Q_ASSIGN U21249 ( .B(clk), .A(\g.we_clk [11525]));
Q_ASSIGN U21250 ( .B(clk), .A(\g.we_clk [11524]));
Q_ASSIGN U21251 ( .B(clk), .A(\g.we_clk [11523]));
Q_ASSIGN U21252 ( .B(clk), .A(\g.we_clk [11522]));
Q_ASSIGN U21253 ( .B(clk), .A(\g.we_clk [11521]));
Q_ASSIGN U21254 ( .B(clk), .A(\g.we_clk [11520]));
Q_ASSIGN U21255 ( .B(clk), .A(\g.we_clk [11519]));
Q_ASSIGN U21256 ( .B(clk), .A(\g.we_clk [11518]));
Q_ASSIGN U21257 ( .B(clk), .A(\g.we_clk [11517]));
Q_ASSIGN U21258 ( .B(clk), .A(\g.we_clk [11516]));
Q_ASSIGN U21259 ( .B(clk), .A(\g.we_clk [11515]));
Q_ASSIGN U21260 ( .B(clk), .A(\g.we_clk [11514]));
Q_ASSIGN U21261 ( .B(clk), .A(\g.we_clk [11513]));
Q_ASSIGN U21262 ( .B(clk), .A(\g.we_clk [11512]));
Q_ASSIGN U21263 ( .B(clk), .A(\g.we_clk [11511]));
Q_ASSIGN U21264 ( .B(clk), .A(\g.we_clk [11510]));
Q_ASSIGN U21265 ( .B(clk), .A(\g.we_clk [11509]));
Q_ASSIGN U21266 ( .B(clk), .A(\g.we_clk [11508]));
Q_ASSIGN U21267 ( .B(clk), .A(\g.we_clk [11507]));
Q_ASSIGN U21268 ( .B(clk), .A(\g.we_clk [11506]));
Q_ASSIGN U21269 ( .B(clk), .A(\g.we_clk [11505]));
Q_ASSIGN U21270 ( .B(clk), .A(\g.we_clk [11504]));
Q_ASSIGN U21271 ( .B(clk), .A(\g.we_clk [11503]));
Q_ASSIGN U21272 ( .B(clk), .A(\g.we_clk [11502]));
Q_ASSIGN U21273 ( .B(clk), .A(\g.we_clk [11501]));
Q_ASSIGN U21274 ( .B(clk), .A(\g.we_clk [11500]));
Q_ASSIGN U21275 ( .B(clk), .A(\g.we_clk [11499]));
Q_ASSIGN U21276 ( .B(clk), .A(\g.we_clk [11498]));
Q_ASSIGN U21277 ( .B(clk), .A(\g.we_clk [11497]));
Q_ASSIGN U21278 ( .B(clk), .A(\g.we_clk [11496]));
Q_ASSIGN U21279 ( .B(clk), .A(\g.we_clk [11495]));
Q_ASSIGN U21280 ( .B(clk), .A(\g.we_clk [11494]));
Q_ASSIGN U21281 ( .B(clk), .A(\g.we_clk [11493]));
Q_ASSIGN U21282 ( .B(clk), .A(\g.we_clk [11492]));
Q_ASSIGN U21283 ( .B(clk), .A(\g.we_clk [11491]));
Q_ASSIGN U21284 ( .B(clk), .A(\g.we_clk [11490]));
Q_ASSIGN U21285 ( .B(clk), .A(\g.we_clk [11489]));
Q_ASSIGN U21286 ( .B(clk), .A(\g.we_clk [11488]));
Q_ASSIGN U21287 ( .B(clk), .A(\g.we_clk [11487]));
Q_ASSIGN U21288 ( .B(clk), .A(\g.we_clk [11486]));
Q_ASSIGN U21289 ( .B(clk), .A(\g.we_clk [11485]));
Q_ASSIGN U21290 ( .B(clk), .A(\g.we_clk [11484]));
Q_ASSIGN U21291 ( .B(clk), .A(\g.we_clk [11483]));
Q_ASSIGN U21292 ( .B(clk), .A(\g.we_clk [11482]));
Q_ASSIGN U21293 ( .B(clk), .A(\g.we_clk [11481]));
Q_ASSIGN U21294 ( .B(clk), .A(\g.we_clk [11480]));
Q_ASSIGN U21295 ( .B(clk), .A(\g.we_clk [11479]));
Q_ASSIGN U21296 ( .B(clk), .A(\g.we_clk [11478]));
Q_ASSIGN U21297 ( .B(clk), .A(\g.we_clk [11477]));
Q_ASSIGN U21298 ( .B(clk), .A(\g.we_clk [11476]));
Q_ASSIGN U21299 ( .B(clk), .A(\g.we_clk [11475]));
Q_ASSIGN U21300 ( .B(clk), .A(\g.we_clk [11474]));
Q_ASSIGN U21301 ( .B(clk), .A(\g.we_clk [11473]));
Q_ASSIGN U21302 ( .B(clk), .A(\g.we_clk [11472]));
Q_ASSIGN U21303 ( .B(clk), .A(\g.we_clk [11471]));
Q_ASSIGN U21304 ( .B(clk), .A(\g.we_clk [11470]));
Q_ASSIGN U21305 ( .B(clk), .A(\g.we_clk [11469]));
Q_ASSIGN U21306 ( .B(clk), .A(\g.we_clk [11468]));
Q_ASSIGN U21307 ( .B(clk), .A(\g.we_clk [11467]));
Q_ASSIGN U21308 ( .B(clk), .A(\g.we_clk [11466]));
Q_ASSIGN U21309 ( .B(clk), .A(\g.we_clk [11465]));
Q_ASSIGN U21310 ( .B(clk), .A(\g.we_clk [11464]));
Q_ASSIGN U21311 ( .B(clk), .A(\g.we_clk [11463]));
Q_ASSIGN U21312 ( .B(clk), .A(\g.we_clk [11462]));
Q_ASSIGN U21313 ( .B(clk), .A(\g.we_clk [11461]));
Q_ASSIGN U21314 ( .B(clk), .A(\g.we_clk [11460]));
Q_ASSIGN U21315 ( .B(clk), .A(\g.we_clk [11459]));
Q_ASSIGN U21316 ( .B(clk), .A(\g.we_clk [11458]));
Q_ASSIGN U21317 ( .B(clk), .A(\g.we_clk [11457]));
Q_ASSIGN U21318 ( .B(clk), .A(\g.we_clk [11456]));
Q_ASSIGN U21319 ( .B(clk), .A(\g.we_clk [11455]));
Q_ASSIGN U21320 ( .B(clk), .A(\g.we_clk [11454]));
Q_ASSIGN U21321 ( .B(clk), .A(\g.we_clk [11453]));
Q_ASSIGN U21322 ( .B(clk), .A(\g.we_clk [11452]));
Q_ASSIGN U21323 ( .B(clk), .A(\g.we_clk [11451]));
Q_ASSIGN U21324 ( .B(clk), .A(\g.we_clk [11450]));
Q_ASSIGN U21325 ( .B(clk), .A(\g.we_clk [11449]));
Q_ASSIGN U21326 ( .B(clk), .A(\g.we_clk [11448]));
Q_ASSIGN U21327 ( .B(clk), .A(\g.we_clk [11447]));
Q_ASSIGN U21328 ( .B(clk), .A(\g.we_clk [11446]));
Q_ASSIGN U21329 ( .B(clk), .A(\g.we_clk [11445]));
Q_ASSIGN U21330 ( .B(clk), .A(\g.we_clk [11444]));
Q_ASSIGN U21331 ( .B(clk), .A(\g.we_clk [11443]));
Q_ASSIGN U21332 ( .B(clk), .A(\g.we_clk [11442]));
Q_ASSIGN U21333 ( .B(clk), .A(\g.we_clk [11441]));
Q_ASSIGN U21334 ( .B(clk), .A(\g.we_clk [11440]));
Q_ASSIGN U21335 ( .B(clk), .A(\g.we_clk [11439]));
Q_ASSIGN U21336 ( .B(clk), .A(\g.we_clk [11438]));
Q_ASSIGN U21337 ( .B(clk), .A(\g.we_clk [11437]));
Q_ASSIGN U21338 ( .B(clk), .A(\g.we_clk [11436]));
Q_ASSIGN U21339 ( .B(clk), .A(\g.we_clk [11435]));
Q_ASSIGN U21340 ( .B(clk), .A(\g.we_clk [11434]));
Q_ASSIGN U21341 ( .B(clk), .A(\g.we_clk [11433]));
Q_ASSIGN U21342 ( .B(clk), .A(\g.we_clk [11432]));
Q_ASSIGN U21343 ( .B(clk), .A(\g.we_clk [11431]));
Q_ASSIGN U21344 ( .B(clk), .A(\g.we_clk [11430]));
Q_ASSIGN U21345 ( .B(clk), .A(\g.we_clk [11429]));
Q_ASSIGN U21346 ( .B(clk), .A(\g.we_clk [11428]));
Q_ASSIGN U21347 ( .B(clk), .A(\g.we_clk [11427]));
Q_ASSIGN U21348 ( .B(clk), .A(\g.we_clk [11426]));
Q_ASSIGN U21349 ( .B(clk), .A(\g.we_clk [11425]));
Q_ASSIGN U21350 ( .B(clk), .A(\g.we_clk [11424]));
Q_ASSIGN U21351 ( .B(clk), .A(\g.we_clk [11423]));
Q_ASSIGN U21352 ( .B(clk), .A(\g.we_clk [11422]));
Q_ASSIGN U21353 ( .B(clk), .A(\g.we_clk [11421]));
Q_ASSIGN U21354 ( .B(clk), .A(\g.we_clk [11420]));
Q_ASSIGN U21355 ( .B(clk), .A(\g.we_clk [11419]));
Q_ASSIGN U21356 ( .B(clk), .A(\g.we_clk [11418]));
Q_ASSIGN U21357 ( .B(clk), .A(\g.we_clk [11417]));
Q_ASSIGN U21358 ( .B(clk), .A(\g.we_clk [11416]));
Q_ASSIGN U21359 ( .B(clk), .A(\g.we_clk [11415]));
Q_ASSIGN U21360 ( .B(clk), .A(\g.we_clk [11414]));
Q_ASSIGN U21361 ( .B(clk), .A(\g.we_clk [11413]));
Q_ASSIGN U21362 ( .B(clk), .A(\g.we_clk [11412]));
Q_ASSIGN U21363 ( .B(clk), .A(\g.we_clk [11411]));
Q_ASSIGN U21364 ( .B(clk), .A(\g.we_clk [11410]));
Q_ASSIGN U21365 ( .B(clk), .A(\g.we_clk [11409]));
Q_ASSIGN U21366 ( .B(clk), .A(\g.we_clk [11408]));
Q_ASSIGN U21367 ( .B(clk), .A(\g.we_clk [11407]));
Q_ASSIGN U21368 ( .B(clk), .A(\g.we_clk [11406]));
Q_ASSIGN U21369 ( .B(clk), .A(\g.we_clk [11405]));
Q_ASSIGN U21370 ( .B(clk), .A(\g.we_clk [11404]));
Q_ASSIGN U21371 ( .B(clk), .A(\g.we_clk [11403]));
Q_ASSIGN U21372 ( .B(clk), .A(\g.we_clk [11402]));
Q_ASSIGN U21373 ( .B(clk), .A(\g.we_clk [11401]));
Q_ASSIGN U21374 ( .B(clk), .A(\g.we_clk [11400]));
Q_ASSIGN U21375 ( .B(clk), .A(\g.we_clk [11399]));
Q_ASSIGN U21376 ( .B(clk), .A(\g.we_clk [11398]));
Q_ASSIGN U21377 ( .B(clk), .A(\g.we_clk [11397]));
Q_ASSIGN U21378 ( .B(clk), .A(\g.we_clk [11396]));
Q_ASSIGN U21379 ( .B(clk), .A(\g.we_clk [11395]));
Q_ASSIGN U21380 ( .B(clk), .A(\g.we_clk [11394]));
Q_ASSIGN U21381 ( .B(clk), .A(\g.we_clk [11393]));
Q_ASSIGN U21382 ( .B(clk), .A(\g.we_clk [11392]));
Q_ASSIGN U21383 ( .B(clk), .A(\g.we_clk [11391]));
Q_ASSIGN U21384 ( .B(clk), .A(\g.we_clk [11390]));
Q_ASSIGN U21385 ( .B(clk), .A(\g.we_clk [11389]));
Q_ASSIGN U21386 ( .B(clk), .A(\g.we_clk [11388]));
Q_ASSIGN U21387 ( .B(clk), .A(\g.we_clk [11387]));
Q_ASSIGN U21388 ( .B(clk), .A(\g.we_clk [11386]));
Q_ASSIGN U21389 ( .B(clk), .A(\g.we_clk [11385]));
Q_ASSIGN U21390 ( .B(clk), .A(\g.we_clk [11384]));
Q_ASSIGN U21391 ( .B(clk), .A(\g.we_clk [11383]));
Q_ASSIGN U21392 ( .B(clk), .A(\g.we_clk [11382]));
Q_ASSIGN U21393 ( .B(clk), .A(\g.we_clk [11381]));
Q_ASSIGN U21394 ( .B(clk), .A(\g.we_clk [11380]));
Q_ASSIGN U21395 ( .B(clk), .A(\g.we_clk [11379]));
Q_ASSIGN U21396 ( .B(clk), .A(\g.we_clk [11378]));
Q_ASSIGN U21397 ( .B(clk), .A(\g.we_clk [11377]));
Q_ASSIGN U21398 ( .B(clk), .A(\g.we_clk [11376]));
Q_ASSIGN U21399 ( .B(clk), .A(\g.we_clk [11375]));
Q_ASSIGN U21400 ( .B(clk), .A(\g.we_clk [11374]));
Q_ASSIGN U21401 ( .B(clk), .A(\g.we_clk [11373]));
Q_ASSIGN U21402 ( .B(clk), .A(\g.we_clk [11372]));
Q_ASSIGN U21403 ( .B(clk), .A(\g.we_clk [11371]));
Q_ASSIGN U21404 ( .B(clk), .A(\g.we_clk [11370]));
Q_ASSIGN U21405 ( .B(clk), .A(\g.we_clk [11369]));
Q_ASSIGN U21406 ( .B(clk), .A(\g.we_clk [11368]));
Q_ASSIGN U21407 ( .B(clk), .A(\g.we_clk [11367]));
Q_ASSIGN U21408 ( .B(clk), .A(\g.we_clk [11366]));
Q_ASSIGN U21409 ( .B(clk), .A(\g.we_clk [11365]));
Q_ASSIGN U21410 ( .B(clk), .A(\g.we_clk [11364]));
Q_ASSIGN U21411 ( .B(clk), .A(\g.we_clk [11363]));
Q_ASSIGN U21412 ( .B(clk), .A(\g.we_clk [11362]));
Q_ASSIGN U21413 ( .B(clk), .A(\g.we_clk [11361]));
Q_ASSIGN U21414 ( .B(clk), .A(\g.we_clk [11360]));
Q_ASSIGN U21415 ( .B(clk), .A(\g.we_clk [11359]));
Q_ASSIGN U21416 ( .B(clk), .A(\g.we_clk [11358]));
Q_ASSIGN U21417 ( .B(clk), .A(\g.we_clk [11357]));
Q_ASSIGN U21418 ( .B(clk), .A(\g.we_clk [11356]));
Q_ASSIGN U21419 ( .B(clk), .A(\g.we_clk [11355]));
Q_ASSIGN U21420 ( .B(clk), .A(\g.we_clk [11354]));
Q_ASSIGN U21421 ( .B(clk), .A(\g.we_clk [11353]));
Q_ASSIGN U21422 ( .B(clk), .A(\g.we_clk [11352]));
Q_ASSIGN U21423 ( .B(clk), .A(\g.we_clk [11351]));
Q_ASSIGN U21424 ( .B(clk), .A(\g.we_clk [11350]));
Q_ASSIGN U21425 ( .B(clk), .A(\g.we_clk [11349]));
Q_ASSIGN U21426 ( .B(clk), .A(\g.we_clk [11348]));
Q_ASSIGN U21427 ( .B(clk), .A(\g.we_clk [11347]));
Q_ASSIGN U21428 ( .B(clk), .A(\g.we_clk [11346]));
Q_ASSIGN U21429 ( .B(clk), .A(\g.we_clk [11345]));
Q_ASSIGN U21430 ( .B(clk), .A(\g.we_clk [11344]));
Q_ASSIGN U21431 ( .B(clk), .A(\g.we_clk [11343]));
Q_ASSIGN U21432 ( .B(clk), .A(\g.we_clk [11342]));
Q_ASSIGN U21433 ( .B(clk), .A(\g.we_clk [11341]));
Q_ASSIGN U21434 ( .B(clk), .A(\g.we_clk [11340]));
Q_ASSIGN U21435 ( .B(clk), .A(\g.we_clk [11339]));
Q_ASSIGN U21436 ( .B(clk), .A(\g.we_clk [11338]));
Q_ASSIGN U21437 ( .B(clk), .A(\g.we_clk [11337]));
Q_ASSIGN U21438 ( .B(clk), .A(\g.we_clk [11336]));
Q_ASSIGN U21439 ( .B(clk), .A(\g.we_clk [11335]));
Q_ASSIGN U21440 ( .B(clk), .A(\g.we_clk [11334]));
Q_ASSIGN U21441 ( .B(clk), .A(\g.we_clk [11333]));
Q_ASSIGN U21442 ( .B(clk), .A(\g.we_clk [11332]));
Q_ASSIGN U21443 ( .B(clk), .A(\g.we_clk [11331]));
Q_ASSIGN U21444 ( .B(clk), .A(\g.we_clk [11330]));
Q_ASSIGN U21445 ( .B(clk), .A(\g.we_clk [11329]));
Q_ASSIGN U21446 ( .B(clk), .A(\g.we_clk [11328]));
Q_ASSIGN U21447 ( .B(clk), .A(\g.we_clk [11327]));
Q_ASSIGN U21448 ( .B(clk), .A(\g.we_clk [11326]));
Q_ASSIGN U21449 ( .B(clk), .A(\g.we_clk [11325]));
Q_ASSIGN U21450 ( .B(clk), .A(\g.we_clk [11324]));
Q_ASSIGN U21451 ( .B(clk), .A(\g.we_clk [11323]));
Q_ASSIGN U21452 ( .B(clk), .A(\g.we_clk [11322]));
Q_ASSIGN U21453 ( .B(clk), .A(\g.we_clk [11321]));
Q_ASSIGN U21454 ( .B(clk), .A(\g.we_clk [11320]));
Q_ASSIGN U21455 ( .B(clk), .A(\g.we_clk [11319]));
Q_ASSIGN U21456 ( .B(clk), .A(\g.we_clk [11318]));
Q_ASSIGN U21457 ( .B(clk), .A(\g.we_clk [11317]));
Q_ASSIGN U21458 ( .B(clk), .A(\g.we_clk [11316]));
Q_ASSIGN U21459 ( .B(clk), .A(\g.we_clk [11315]));
Q_ASSIGN U21460 ( .B(clk), .A(\g.we_clk [11314]));
Q_ASSIGN U21461 ( .B(clk), .A(\g.we_clk [11313]));
Q_ASSIGN U21462 ( .B(clk), .A(\g.we_clk [11312]));
Q_ASSIGN U21463 ( .B(clk), .A(\g.we_clk [11311]));
Q_ASSIGN U21464 ( .B(clk), .A(\g.we_clk [11310]));
Q_ASSIGN U21465 ( .B(clk), .A(\g.we_clk [11309]));
Q_ASSIGN U21466 ( .B(clk), .A(\g.we_clk [11308]));
Q_ASSIGN U21467 ( .B(clk), .A(\g.we_clk [11307]));
Q_ASSIGN U21468 ( .B(clk), .A(\g.we_clk [11306]));
Q_ASSIGN U21469 ( .B(clk), .A(\g.we_clk [11305]));
Q_ASSIGN U21470 ( .B(clk), .A(\g.we_clk [11304]));
Q_ASSIGN U21471 ( .B(clk), .A(\g.we_clk [11303]));
Q_ASSIGN U21472 ( .B(clk), .A(\g.we_clk [11302]));
Q_ASSIGN U21473 ( .B(clk), .A(\g.we_clk [11301]));
Q_ASSIGN U21474 ( .B(clk), .A(\g.we_clk [11300]));
Q_ASSIGN U21475 ( .B(clk), .A(\g.we_clk [11299]));
Q_ASSIGN U21476 ( .B(clk), .A(\g.we_clk [11298]));
Q_ASSIGN U21477 ( .B(clk), .A(\g.we_clk [11297]));
Q_ASSIGN U21478 ( .B(clk), .A(\g.we_clk [11296]));
Q_ASSIGN U21479 ( .B(clk), .A(\g.we_clk [11295]));
Q_ASSIGN U21480 ( .B(clk), .A(\g.we_clk [11294]));
Q_ASSIGN U21481 ( .B(clk), .A(\g.we_clk [11293]));
Q_ASSIGN U21482 ( .B(clk), .A(\g.we_clk [11292]));
Q_ASSIGN U21483 ( .B(clk), .A(\g.we_clk [11291]));
Q_ASSIGN U21484 ( .B(clk), .A(\g.we_clk [11290]));
Q_ASSIGN U21485 ( .B(clk), .A(\g.we_clk [11289]));
Q_ASSIGN U21486 ( .B(clk), .A(\g.we_clk [11288]));
Q_ASSIGN U21487 ( .B(clk), .A(\g.we_clk [11287]));
Q_ASSIGN U21488 ( .B(clk), .A(\g.we_clk [11286]));
Q_ASSIGN U21489 ( .B(clk), .A(\g.we_clk [11285]));
Q_ASSIGN U21490 ( .B(clk), .A(\g.we_clk [11284]));
Q_ASSIGN U21491 ( .B(clk), .A(\g.we_clk [11283]));
Q_ASSIGN U21492 ( .B(clk), .A(\g.we_clk [11282]));
Q_ASSIGN U21493 ( .B(clk), .A(\g.we_clk [11281]));
Q_ASSIGN U21494 ( .B(clk), .A(\g.we_clk [11280]));
Q_ASSIGN U21495 ( .B(clk), .A(\g.we_clk [11279]));
Q_ASSIGN U21496 ( .B(clk), .A(\g.we_clk [11278]));
Q_ASSIGN U21497 ( .B(clk), .A(\g.we_clk [11277]));
Q_ASSIGN U21498 ( .B(clk), .A(\g.we_clk [11276]));
Q_ASSIGN U21499 ( .B(clk), .A(\g.we_clk [11275]));
Q_ASSIGN U21500 ( .B(clk), .A(\g.we_clk [11274]));
Q_ASSIGN U21501 ( .B(clk), .A(\g.we_clk [11273]));
Q_ASSIGN U21502 ( .B(clk), .A(\g.we_clk [11272]));
Q_ASSIGN U21503 ( .B(clk), .A(\g.we_clk [11271]));
Q_ASSIGN U21504 ( .B(clk), .A(\g.we_clk [11270]));
Q_ASSIGN U21505 ( .B(clk), .A(\g.we_clk [11269]));
Q_ASSIGN U21506 ( .B(clk), .A(\g.we_clk [11268]));
Q_ASSIGN U21507 ( .B(clk), .A(\g.we_clk [11267]));
Q_ASSIGN U21508 ( .B(clk), .A(\g.we_clk [11266]));
Q_ASSIGN U21509 ( .B(clk), .A(\g.we_clk [11265]));
Q_ASSIGN U21510 ( .B(clk), .A(\g.we_clk [11264]));
Q_ASSIGN U21511 ( .B(clk), .A(\g.we_clk [11263]));
Q_ASSIGN U21512 ( .B(clk), .A(\g.we_clk [11262]));
Q_ASSIGN U21513 ( .B(clk), .A(\g.we_clk [11261]));
Q_ASSIGN U21514 ( .B(clk), .A(\g.we_clk [11260]));
Q_ASSIGN U21515 ( .B(clk), .A(\g.we_clk [11259]));
Q_ASSIGN U21516 ( .B(clk), .A(\g.we_clk [11258]));
Q_ASSIGN U21517 ( .B(clk), .A(\g.we_clk [11257]));
Q_ASSIGN U21518 ( .B(clk), .A(\g.we_clk [11256]));
Q_ASSIGN U21519 ( .B(clk), .A(\g.we_clk [11255]));
Q_ASSIGN U21520 ( .B(clk), .A(\g.we_clk [11254]));
Q_ASSIGN U21521 ( .B(clk), .A(\g.we_clk [11253]));
Q_ASSIGN U21522 ( .B(clk), .A(\g.we_clk [11252]));
Q_ASSIGN U21523 ( .B(clk), .A(\g.we_clk [11251]));
Q_ASSIGN U21524 ( .B(clk), .A(\g.we_clk [11250]));
Q_ASSIGN U21525 ( .B(clk), .A(\g.we_clk [11249]));
Q_ASSIGN U21526 ( .B(clk), .A(\g.we_clk [11248]));
Q_ASSIGN U21527 ( .B(clk), .A(\g.we_clk [11247]));
Q_ASSIGN U21528 ( .B(clk), .A(\g.we_clk [11246]));
Q_ASSIGN U21529 ( .B(clk), .A(\g.we_clk [11245]));
Q_ASSIGN U21530 ( .B(clk), .A(\g.we_clk [11244]));
Q_ASSIGN U21531 ( .B(clk), .A(\g.we_clk [11243]));
Q_ASSIGN U21532 ( .B(clk), .A(\g.we_clk [11242]));
Q_ASSIGN U21533 ( .B(clk), .A(\g.we_clk [11241]));
Q_ASSIGN U21534 ( .B(clk), .A(\g.we_clk [11240]));
Q_ASSIGN U21535 ( .B(clk), .A(\g.we_clk [11239]));
Q_ASSIGN U21536 ( .B(clk), .A(\g.we_clk [11238]));
Q_ASSIGN U21537 ( .B(clk), .A(\g.we_clk [11237]));
Q_ASSIGN U21538 ( .B(clk), .A(\g.we_clk [11236]));
Q_ASSIGN U21539 ( .B(clk), .A(\g.we_clk [11235]));
Q_ASSIGN U21540 ( .B(clk), .A(\g.we_clk [11234]));
Q_ASSIGN U21541 ( .B(clk), .A(\g.we_clk [11233]));
Q_ASSIGN U21542 ( .B(clk), .A(\g.we_clk [11232]));
Q_ASSIGN U21543 ( .B(clk), .A(\g.we_clk [11231]));
Q_ASSIGN U21544 ( .B(clk), .A(\g.we_clk [11230]));
Q_ASSIGN U21545 ( .B(clk), .A(\g.we_clk [11229]));
Q_ASSIGN U21546 ( .B(clk), .A(\g.we_clk [11228]));
Q_ASSIGN U21547 ( .B(clk), .A(\g.we_clk [11227]));
Q_ASSIGN U21548 ( .B(clk), .A(\g.we_clk [11226]));
Q_ASSIGN U21549 ( .B(clk), .A(\g.we_clk [11225]));
Q_ASSIGN U21550 ( .B(clk), .A(\g.we_clk [11224]));
Q_ASSIGN U21551 ( .B(clk), .A(\g.we_clk [11223]));
Q_ASSIGN U21552 ( .B(clk), .A(\g.we_clk [11222]));
Q_ASSIGN U21553 ( .B(clk), .A(\g.we_clk [11221]));
Q_ASSIGN U21554 ( .B(clk), .A(\g.we_clk [11220]));
Q_ASSIGN U21555 ( .B(clk), .A(\g.we_clk [11219]));
Q_ASSIGN U21556 ( .B(clk), .A(\g.we_clk [11218]));
Q_ASSIGN U21557 ( .B(clk), .A(\g.we_clk [11217]));
Q_ASSIGN U21558 ( .B(clk), .A(\g.we_clk [11216]));
Q_ASSIGN U21559 ( .B(clk), .A(\g.we_clk [11215]));
Q_ASSIGN U21560 ( .B(clk), .A(\g.we_clk [11214]));
Q_ASSIGN U21561 ( .B(clk), .A(\g.we_clk [11213]));
Q_ASSIGN U21562 ( .B(clk), .A(\g.we_clk [11212]));
Q_ASSIGN U21563 ( .B(clk), .A(\g.we_clk [11211]));
Q_ASSIGN U21564 ( .B(clk), .A(\g.we_clk [11210]));
Q_ASSIGN U21565 ( .B(clk), .A(\g.we_clk [11209]));
Q_ASSIGN U21566 ( .B(clk), .A(\g.we_clk [11208]));
Q_ASSIGN U21567 ( .B(clk), .A(\g.we_clk [11207]));
Q_ASSIGN U21568 ( .B(clk), .A(\g.we_clk [11206]));
Q_ASSIGN U21569 ( .B(clk), .A(\g.we_clk [11205]));
Q_ASSIGN U21570 ( .B(clk), .A(\g.we_clk [11204]));
Q_ASSIGN U21571 ( .B(clk), .A(\g.we_clk [11203]));
Q_ASSIGN U21572 ( .B(clk), .A(\g.we_clk [11202]));
Q_ASSIGN U21573 ( .B(clk), .A(\g.we_clk [11201]));
Q_ASSIGN U21574 ( .B(clk), .A(\g.we_clk [11200]));
Q_ASSIGN U21575 ( .B(clk), .A(\g.we_clk [11199]));
Q_ASSIGN U21576 ( .B(clk), .A(\g.we_clk [11198]));
Q_ASSIGN U21577 ( .B(clk), .A(\g.we_clk [11197]));
Q_ASSIGN U21578 ( .B(clk), .A(\g.we_clk [11196]));
Q_ASSIGN U21579 ( .B(clk), .A(\g.we_clk [11195]));
Q_ASSIGN U21580 ( .B(clk), .A(\g.we_clk [11194]));
Q_ASSIGN U21581 ( .B(clk), .A(\g.we_clk [11193]));
Q_ASSIGN U21582 ( .B(clk), .A(\g.we_clk [11192]));
Q_ASSIGN U21583 ( .B(clk), .A(\g.we_clk [11191]));
Q_ASSIGN U21584 ( .B(clk), .A(\g.we_clk [11190]));
Q_ASSIGN U21585 ( .B(clk), .A(\g.we_clk [11189]));
Q_ASSIGN U21586 ( .B(clk), .A(\g.we_clk [11188]));
Q_ASSIGN U21587 ( .B(clk), .A(\g.we_clk [11187]));
Q_ASSIGN U21588 ( .B(clk), .A(\g.we_clk [11186]));
Q_ASSIGN U21589 ( .B(clk), .A(\g.we_clk [11185]));
Q_ASSIGN U21590 ( .B(clk), .A(\g.we_clk [11184]));
Q_ASSIGN U21591 ( .B(clk), .A(\g.we_clk [11183]));
Q_ASSIGN U21592 ( .B(clk), .A(\g.we_clk [11182]));
Q_ASSIGN U21593 ( .B(clk), .A(\g.we_clk [11181]));
Q_ASSIGN U21594 ( .B(clk), .A(\g.we_clk [11180]));
Q_ASSIGN U21595 ( .B(clk), .A(\g.we_clk [11179]));
Q_ASSIGN U21596 ( .B(clk), .A(\g.we_clk [11178]));
Q_ASSIGN U21597 ( .B(clk), .A(\g.we_clk [11177]));
Q_ASSIGN U21598 ( .B(clk), .A(\g.we_clk [11176]));
Q_ASSIGN U21599 ( .B(clk), .A(\g.we_clk [11175]));
Q_ASSIGN U21600 ( .B(clk), .A(\g.we_clk [11174]));
Q_ASSIGN U21601 ( .B(clk), .A(\g.we_clk [11173]));
Q_ASSIGN U21602 ( .B(clk), .A(\g.we_clk [11172]));
Q_ASSIGN U21603 ( .B(clk), .A(\g.we_clk [11171]));
Q_ASSIGN U21604 ( .B(clk), .A(\g.we_clk [11170]));
Q_ASSIGN U21605 ( .B(clk), .A(\g.we_clk [11169]));
Q_ASSIGN U21606 ( .B(clk), .A(\g.we_clk [11168]));
Q_ASSIGN U21607 ( .B(clk), .A(\g.we_clk [11167]));
Q_ASSIGN U21608 ( .B(clk), .A(\g.we_clk [11166]));
Q_ASSIGN U21609 ( .B(clk), .A(\g.we_clk [11165]));
Q_ASSIGN U21610 ( .B(clk), .A(\g.we_clk [11164]));
Q_ASSIGN U21611 ( .B(clk), .A(\g.we_clk [11163]));
Q_ASSIGN U21612 ( .B(clk), .A(\g.we_clk [11162]));
Q_ASSIGN U21613 ( .B(clk), .A(\g.we_clk [11161]));
Q_ASSIGN U21614 ( .B(clk), .A(\g.we_clk [11160]));
Q_ASSIGN U21615 ( .B(clk), .A(\g.we_clk [11159]));
Q_ASSIGN U21616 ( .B(clk), .A(\g.we_clk [11158]));
Q_ASSIGN U21617 ( .B(clk), .A(\g.we_clk [11157]));
Q_ASSIGN U21618 ( .B(clk), .A(\g.we_clk [11156]));
Q_ASSIGN U21619 ( .B(clk), .A(\g.we_clk [11155]));
Q_ASSIGN U21620 ( .B(clk), .A(\g.we_clk [11154]));
Q_ASSIGN U21621 ( .B(clk), .A(\g.we_clk [11153]));
Q_ASSIGN U21622 ( .B(clk), .A(\g.we_clk [11152]));
Q_ASSIGN U21623 ( .B(clk), .A(\g.we_clk [11151]));
Q_ASSIGN U21624 ( .B(clk), .A(\g.we_clk [11150]));
Q_ASSIGN U21625 ( .B(clk), .A(\g.we_clk [11149]));
Q_ASSIGN U21626 ( .B(clk), .A(\g.we_clk [11148]));
Q_ASSIGN U21627 ( .B(clk), .A(\g.we_clk [11147]));
Q_ASSIGN U21628 ( .B(clk), .A(\g.we_clk [11146]));
Q_ASSIGN U21629 ( .B(clk), .A(\g.we_clk [11145]));
Q_ASSIGN U21630 ( .B(clk), .A(\g.we_clk [11144]));
Q_ASSIGN U21631 ( .B(clk), .A(\g.we_clk [11143]));
Q_ASSIGN U21632 ( .B(clk), .A(\g.we_clk [11142]));
Q_ASSIGN U21633 ( .B(clk), .A(\g.we_clk [11141]));
Q_ASSIGN U21634 ( .B(clk), .A(\g.we_clk [11140]));
Q_ASSIGN U21635 ( .B(clk), .A(\g.we_clk [11139]));
Q_ASSIGN U21636 ( .B(clk), .A(\g.we_clk [11138]));
Q_ASSIGN U21637 ( .B(clk), .A(\g.we_clk [11137]));
Q_ASSIGN U21638 ( .B(clk), .A(\g.we_clk [11136]));
Q_ASSIGN U21639 ( .B(clk), .A(\g.we_clk [11135]));
Q_ASSIGN U21640 ( .B(clk), .A(\g.we_clk [11134]));
Q_ASSIGN U21641 ( .B(clk), .A(\g.we_clk [11133]));
Q_ASSIGN U21642 ( .B(clk), .A(\g.we_clk [11132]));
Q_ASSIGN U21643 ( .B(clk), .A(\g.we_clk [11131]));
Q_ASSIGN U21644 ( .B(clk), .A(\g.we_clk [11130]));
Q_ASSIGN U21645 ( .B(clk), .A(\g.we_clk [11129]));
Q_ASSIGN U21646 ( .B(clk), .A(\g.we_clk [11128]));
Q_ASSIGN U21647 ( .B(clk), .A(\g.we_clk [11127]));
Q_ASSIGN U21648 ( .B(clk), .A(\g.we_clk [11126]));
Q_ASSIGN U21649 ( .B(clk), .A(\g.we_clk [11125]));
Q_ASSIGN U21650 ( .B(clk), .A(\g.we_clk [11124]));
Q_ASSIGN U21651 ( .B(clk), .A(\g.we_clk [11123]));
Q_ASSIGN U21652 ( .B(clk), .A(\g.we_clk [11122]));
Q_ASSIGN U21653 ( .B(clk), .A(\g.we_clk [11121]));
Q_ASSIGN U21654 ( .B(clk), .A(\g.we_clk [11120]));
Q_ASSIGN U21655 ( .B(clk), .A(\g.we_clk [11119]));
Q_ASSIGN U21656 ( .B(clk), .A(\g.we_clk [11118]));
Q_ASSIGN U21657 ( .B(clk), .A(\g.we_clk [11117]));
Q_ASSIGN U21658 ( .B(clk), .A(\g.we_clk [11116]));
Q_ASSIGN U21659 ( .B(clk), .A(\g.we_clk [11115]));
Q_ASSIGN U21660 ( .B(clk), .A(\g.we_clk [11114]));
Q_ASSIGN U21661 ( .B(clk), .A(\g.we_clk [11113]));
Q_ASSIGN U21662 ( .B(clk), .A(\g.we_clk [11112]));
Q_ASSIGN U21663 ( .B(clk), .A(\g.we_clk [11111]));
Q_ASSIGN U21664 ( .B(clk), .A(\g.we_clk [11110]));
Q_ASSIGN U21665 ( .B(clk), .A(\g.we_clk [11109]));
Q_ASSIGN U21666 ( .B(clk), .A(\g.we_clk [11108]));
Q_ASSIGN U21667 ( .B(clk), .A(\g.we_clk [11107]));
Q_ASSIGN U21668 ( .B(clk), .A(\g.we_clk [11106]));
Q_ASSIGN U21669 ( .B(clk), .A(\g.we_clk [11105]));
Q_ASSIGN U21670 ( .B(clk), .A(\g.we_clk [11104]));
Q_ASSIGN U21671 ( .B(clk), .A(\g.we_clk [11103]));
Q_ASSIGN U21672 ( .B(clk), .A(\g.we_clk [11102]));
Q_ASSIGN U21673 ( .B(clk), .A(\g.we_clk [11101]));
Q_ASSIGN U21674 ( .B(clk), .A(\g.we_clk [11100]));
Q_ASSIGN U21675 ( .B(clk), .A(\g.we_clk [11099]));
Q_ASSIGN U21676 ( .B(clk), .A(\g.we_clk [11098]));
Q_ASSIGN U21677 ( .B(clk), .A(\g.we_clk [11097]));
Q_ASSIGN U21678 ( .B(clk), .A(\g.we_clk [11096]));
Q_ASSIGN U21679 ( .B(clk), .A(\g.we_clk [11095]));
Q_ASSIGN U21680 ( .B(clk), .A(\g.we_clk [11094]));
Q_ASSIGN U21681 ( .B(clk), .A(\g.we_clk [11093]));
Q_ASSIGN U21682 ( .B(clk), .A(\g.we_clk [11092]));
Q_ASSIGN U21683 ( .B(clk), .A(\g.we_clk [11091]));
Q_ASSIGN U21684 ( .B(clk), .A(\g.we_clk [11090]));
Q_ASSIGN U21685 ( .B(clk), .A(\g.we_clk [11089]));
Q_ASSIGN U21686 ( .B(clk), .A(\g.we_clk [11088]));
Q_ASSIGN U21687 ( .B(clk), .A(\g.we_clk [11087]));
Q_ASSIGN U21688 ( .B(clk), .A(\g.we_clk [11086]));
Q_ASSIGN U21689 ( .B(clk), .A(\g.we_clk [11085]));
Q_ASSIGN U21690 ( .B(clk), .A(\g.we_clk [11084]));
Q_ASSIGN U21691 ( .B(clk), .A(\g.we_clk [11083]));
Q_ASSIGN U21692 ( .B(clk), .A(\g.we_clk [11082]));
Q_ASSIGN U21693 ( .B(clk), .A(\g.we_clk [11081]));
Q_ASSIGN U21694 ( .B(clk), .A(\g.we_clk [11080]));
Q_ASSIGN U21695 ( .B(clk), .A(\g.we_clk [11079]));
Q_ASSIGN U21696 ( .B(clk), .A(\g.we_clk [11078]));
Q_ASSIGN U21697 ( .B(clk), .A(\g.we_clk [11077]));
Q_ASSIGN U21698 ( .B(clk), .A(\g.we_clk [11076]));
Q_ASSIGN U21699 ( .B(clk), .A(\g.we_clk [11075]));
Q_ASSIGN U21700 ( .B(clk), .A(\g.we_clk [11074]));
Q_ASSIGN U21701 ( .B(clk), .A(\g.we_clk [11073]));
Q_ASSIGN U21702 ( .B(clk), .A(\g.we_clk [11072]));
Q_ASSIGN U21703 ( .B(clk), .A(\g.we_clk [11071]));
Q_ASSIGN U21704 ( .B(clk), .A(\g.we_clk [11070]));
Q_ASSIGN U21705 ( .B(clk), .A(\g.we_clk [11069]));
Q_ASSIGN U21706 ( .B(clk), .A(\g.we_clk [11068]));
Q_ASSIGN U21707 ( .B(clk), .A(\g.we_clk [11067]));
Q_ASSIGN U21708 ( .B(clk), .A(\g.we_clk [11066]));
Q_ASSIGN U21709 ( .B(clk), .A(\g.we_clk [11065]));
Q_ASSIGN U21710 ( .B(clk), .A(\g.we_clk [11064]));
Q_ASSIGN U21711 ( .B(clk), .A(\g.we_clk [11063]));
Q_ASSIGN U21712 ( .B(clk), .A(\g.we_clk [11062]));
Q_ASSIGN U21713 ( .B(clk), .A(\g.we_clk [11061]));
Q_ASSIGN U21714 ( .B(clk), .A(\g.we_clk [11060]));
Q_ASSIGN U21715 ( .B(clk), .A(\g.we_clk [11059]));
Q_ASSIGN U21716 ( .B(clk), .A(\g.we_clk [11058]));
Q_ASSIGN U21717 ( .B(clk), .A(\g.we_clk [11057]));
Q_ASSIGN U21718 ( .B(clk), .A(\g.we_clk [11056]));
Q_ASSIGN U21719 ( .B(clk), .A(\g.we_clk [11055]));
Q_ASSIGN U21720 ( .B(clk), .A(\g.we_clk [11054]));
Q_ASSIGN U21721 ( .B(clk), .A(\g.we_clk [11053]));
Q_ASSIGN U21722 ( .B(clk), .A(\g.we_clk [11052]));
Q_ASSIGN U21723 ( .B(clk), .A(\g.we_clk [11051]));
Q_ASSIGN U21724 ( .B(clk), .A(\g.we_clk [11050]));
Q_ASSIGN U21725 ( .B(clk), .A(\g.we_clk [11049]));
Q_ASSIGN U21726 ( .B(clk), .A(\g.we_clk [11048]));
Q_ASSIGN U21727 ( .B(clk), .A(\g.we_clk [11047]));
Q_ASSIGN U21728 ( .B(clk), .A(\g.we_clk [11046]));
Q_ASSIGN U21729 ( .B(clk), .A(\g.we_clk [11045]));
Q_ASSIGN U21730 ( .B(clk), .A(\g.we_clk [11044]));
Q_ASSIGN U21731 ( .B(clk), .A(\g.we_clk [11043]));
Q_ASSIGN U21732 ( .B(clk), .A(\g.we_clk [11042]));
Q_ASSIGN U21733 ( .B(clk), .A(\g.we_clk [11041]));
Q_ASSIGN U21734 ( .B(clk), .A(\g.we_clk [11040]));
Q_ASSIGN U21735 ( .B(clk), .A(\g.we_clk [11039]));
Q_ASSIGN U21736 ( .B(clk), .A(\g.we_clk [11038]));
Q_ASSIGN U21737 ( .B(clk), .A(\g.we_clk [11037]));
Q_ASSIGN U21738 ( .B(clk), .A(\g.we_clk [11036]));
Q_ASSIGN U21739 ( .B(clk), .A(\g.we_clk [11035]));
Q_ASSIGN U21740 ( .B(clk), .A(\g.we_clk [11034]));
Q_ASSIGN U21741 ( .B(clk), .A(\g.we_clk [11033]));
Q_ASSIGN U21742 ( .B(clk), .A(\g.we_clk [11032]));
Q_ASSIGN U21743 ( .B(clk), .A(\g.we_clk [11031]));
Q_ASSIGN U21744 ( .B(clk), .A(\g.we_clk [11030]));
Q_ASSIGN U21745 ( .B(clk), .A(\g.we_clk [11029]));
Q_ASSIGN U21746 ( .B(clk), .A(\g.we_clk [11028]));
Q_ASSIGN U21747 ( .B(clk), .A(\g.we_clk [11027]));
Q_ASSIGN U21748 ( .B(clk), .A(\g.we_clk [11026]));
Q_ASSIGN U21749 ( .B(clk), .A(\g.we_clk [11025]));
Q_ASSIGN U21750 ( .B(clk), .A(\g.we_clk [11024]));
Q_ASSIGN U21751 ( .B(clk), .A(\g.we_clk [11023]));
Q_ASSIGN U21752 ( .B(clk), .A(\g.we_clk [11022]));
Q_ASSIGN U21753 ( .B(clk), .A(\g.we_clk [11021]));
Q_ASSIGN U21754 ( .B(clk), .A(\g.we_clk [11020]));
Q_ASSIGN U21755 ( .B(clk), .A(\g.we_clk [11019]));
Q_ASSIGN U21756 ( .B(clk), .A(\g.we_clk [11018]));
Q_ASSIGN U21757 ( .B(clk), .A(\g.we_clk [11017]));
Q_ASSIGN U21758 ( .B(clk), .A(\g.we_clk [11016]));
Q_ASSIGN U21759 ( .B(clk), .A(\g.we_clk [11015]));
Q_ASSIGN U21760 ( .B(clk), .A(\g.we_clk [11014]));
Q_ASSIGN U21761 ( .B(clk), .A(\g.we_clk [11013]));
Q_ASSIGN U21762 ( .B(clk), .A(\g.we_clk [11012]));
Q_ASSIGN U21763 ( .B(clk), .A(\g.we_clk [11011]));
Q_ASSIGN U21764 ( .B(clk), .A(\g.we_clk [11010]));
Q_ASSIGN U21765 ( .B(clk), .A(\g.we_clk [11009]));
Q_ASSIGN U21766 ( .B(clk), .A(\g.we_clk [11008]));
Q_ASSIGN U21767 ( .B(clk), .A(\g.we_clk [11007]));
Q_ASSIGN U21768 ( .B(clk), .A(\g.we_clk [11006]));
Q_ASSIGN U21769 ( .B(clk), .A(\g.we_clk [11005]));
Q_ASSIGN U21770 ( .B(clk), .A(\g.we_clk [11004]));
Q_ASSIGN U21771 ( .B(clk), .A(\g.we_clk [11003]));
Q_ASSIGN U21772 ( .B(clk), .A(\g.we_clk [11002]));
Q_ASSIGN U21773 ( .B(clk), .A(\g.we_clk [11001]));
Q_ASSIGN U21774 ( .B(clk), .A(\g.we_clk [11000]));
Q_ASSIGN U21775 ( .B(clk), .A(\g.we_clk [10999]));
Q_ASSIGN U21776 ( .B(clk), .A(\g.we_clk [10998]));
Q_ASSIGN U21777 ( .B(clk), .A(\g.we_clk [10997]));
Q_ASSIGN U21778 ( .B(clk), .A(\g.we_clk [10996]));
Q_ASSIGN U21779 ( .B(clk), .A(\g.we_clk [10995]));
Q_ASSIGN U21780 ( .B(clk), .A(\g.we_clk [10994]));
Q_ASSIGN U21781 ( .B(clk), .A(\g.we_clk [10993]));
Q_ASSIGN U21782 ( .B(clk), .A(\g.we_clk [10992]));
Q_ASSIGN U21783 ( .B(clk), .A(\g.we_clk [10991]));
Q_ASSIGN U21784 ( .B(clk), .A(\g.we_clk [10990]));
Q_ASSIGN U21785 ( .B(clk), .A(\g.we_clk [10989]));
Q_ASSIGN U21786 ( .B(clk), .A(\g.we_clk [10988]));
Q_ASSIGN U21787 ( .B(clk), .A(\g.we_clk [10987]));
Q_ASSIGN U21788 ( .B(clk), .A(\g.we_clk [10986]));
Q_ASSIGN U21789 ( .B(clk), .A(\g.we_clk [10985]));
Q_ASSIGN U21790 ( .B(clk), .A(\g.we_clk [10984]));
Q_ASSIGN U21791 ( .B(clk), .A(\g.we_clk [10983]));
Q_ASSIGN U21792 ( .B(clk), .A(\g.we_clk [10982]));
Q_ASSIGN U21793 ( .B(clk), .A(\g.we_clk [10981]));
Q_ASSIGN U21794 ( .B(clk), .A(\g.we_clk [10980]));
Q_ASSIGN U21795 ( .B(clk), .A(\g.we_clk [10979]));
Q_ASSIGN U21796 ( .B(clk), .A(\g.we_clk [10978]));
Q_ASSIGN U21797 ( .B(clk), .A(\g.we_clk [10977]));
Q_ASSIGN U21798 ( .B(clk), .A(\g.we_clk [10976]));
Q_ASSIGN U21799 ( .B(clk), .A(\g.we_clk [10975]));
Q_ASSIGN U21800 ( .B(clk), .A(\g.we_clk [10974]));
Q_ASSIGN U21801 ( .B(clk), .A(\g.we_clk [10973]));
Q_ASSIGN U21802 ( .B(clk), .A(\g.we_clk [10972]));
Q_ASSIGN U21803 ( .B(clk), .A(\g.we_clk [10971]));
Q_ASSIGN U21804 ( .B(clk), .A(\g.we_clk [10970]));
Q_ASSIGN U21805 ( .B(clk), .A(\g.we_clk [10969]));
Q_ASSIGN U21806 ( .B(clk), .A(\g.we_clk [10968]));
Q_ASSIGN U21807 ( .B(clk), .A(\g.we_clk [10967]));
Q_ASSIGN U21808 ( .B(clk), .A(\g.we_clk [10966]));
Q_ASSIGN U21809 ( .B(clk), .A(\g.we_clk [10965]));
Q_ASSIGN U21810 ( .B(clk), .A(\g.we_clk [10964]));
Q_ASSIGN U21811 ( .B(clk), .A(\g.we_clk [10963]));
Q_ASSIGN U21812 ( .B(clk), .A(\g.we_clk [10962]));
Q_ASSIGN U21813 ( .B(clk), .A(\g.we_clk [10961]));
Q_ASSIGN U21814 ( .B(clk), .A(\g.we_clk [10960]));
Q_ASSIGN U21815 ( .B(clk), .A(\g.we_clk [10959]));
Q_ASSIGN U21816 ( .B(clk), .A(\g.we_clk [10958]));
Q_ASSIGN U21817 ( .B(clk), .A(\g.we_clk [10957]));
Q_ASSIGN U21818 ( .B(clk), .A(\g.we_clk [10956]));
Q_ASSIGN U21819 ( .B(clk), .A(\g.we_clk [10955]));
Q_ASSIGN U21820 ( .B(clk), .A(\g.we_clk [10954]));
Q_ASSIGN U21821 ( .B(clk), .A(\g.we_clk [10953]));
Q_ASSIGN U21822 ( .B(clk), .A(\g.we_clk [10952]));
Q_ASSIGN U21823 ( .B(clk), .A(\g.we_clk [10951]));
Q_ASSIGN U21824 ( .B(clk), .A(\g.we_clk [10950]));
Q_ASSIGN U21825 ( .B(clk), .A(\g.we_clk [10949]));
Q_ASSIGN U21826 ( .B(clk), .A(\g.we_clk [10948]));
Q_ASSIGN U21827 ( .B(clk), .A(\g.we_clk [10947]));
Q_ASSIGN U21828 ( .B(clk), .A(\g.we_clk [10946]));
Q_ASSIGN U21829 ( .B(clk), .A(\g.we_clk [10945]));
Q_ASSIGN U21830 ( .B(clk), .A(\g.we_clk [10944]));
Q_ASSIGN U21831 ( .B(clk), .A(\g.we_clk [10943]));
Q_ASSIGN U21832 ( .B(clk), .A(\g.we_clk [10942]));
Q_ASSIGN U21833 ( .B(clk), .A(\g.we_clk [10941]));
Q_ASSIGN U21834 ( .B(clk), .A(\g.we_clk [10940]));
Q_ASSIGN U21835 ( .B(clk), .A(\g.we_clk [10939]));
Q_ASSIGN U21836 ( .B(clk), .A(\g.we_clk [10938]));
Q_ASSIGN U21837 ( .B(clk), .A(\g.we_clk [10937]));
Q_ASSIGN U21838 ( .B(clk), .A(\g.we_clk [10936]));
Q_ASSIGN U21839 ( .B(clk), .A(\g.we_clk [10935]));
Q_ASSIGN U21840 ( .B(clk), .A(\g.we_clk [10934]));
Q_ASSIGN U21841 ( .B(clk), .A(\g.we_clk [10933]));
Q_ASSIGN U21842 ( .B(clk), .A(\g.we_clk [10932]));
Q_ASSIGN U21843 ( .B(clk), .A(\g.we_clk [10931]));
Q_ASSIGN U21844 ( .B(clk), .A(\g.we_clk [10930]));
Q_ASSIGN U21845 ( .B(clk), .A(\g.we_clk [10929]));
Q_ASSIGN U21846 ( .B(clk), .A(\g.we_clk [10928]));
Q_ASSIGN U21847 ( .B(clk), .A(\g.we_clk [10927]));
Q_ASSIGN U21848 ( .B(clk), .A(\g.we_clk [10926]));
Q_ASSIGN U21849 ( .B(clk), .A(\g.we_clk [10925]));
Q_ASSIGN U21850 ( .B(clk), .A(\g.we_clk [10924]));
Q_ASSIGN U21851 ( .B(clk), .A(\g.we_clk [10923]));
Q_ASSIGN U21852 ( .B(clk), .A(\g.we_clk [10922]));
Q_ASSIGN U21853 ( .B(clk), .A(\g.we_clk [10921]));
Q_ASSIGN U21854 ( .B(clk), .A(\g.we_clk [10920]));
Q_ASSIGN U21855 ( .B(clk), .A(\g.we_clk [10919]));
Q_ASSIGN U21856 ( .B(clk), .A(\g.we_clk [10918]));
Q_ASSIGN U21857 ( .B(clk), .A(\g.we_clk [10917]));
Q_ASSIGN U21858 ( .B(clk), .A(\g.we_clk [10916]));
Q_ASSIGN U21859 ( .B(clk), .A(\g.we_clk [10915]));
Q_ASSIGN U21860 ( .B(clk), .A(\g.we_clk [10914]));
Q_ASSIGN U21861 ( .B(clk), .A(\g.we_clk [10913]));
Q_ASSIGN U21862 ( .B(clk), .A(\g.we_clk [10912]));
Q_ASSIGN U21863 ( .B(clk), .A(\g.we_clk [10911]));
Q_ASSIGN U21864 ( .B(clk), .A(\g.we_clk [10910]));
Q_ASSIGN U21865 ( .B(clk), .A(\g.we_clk [10909]));
Q_ASSIGN U21866 ( .B(clk), .A(\g.we_clk [10908]));
Q_ASSIGN U21867 ( .B(clk), .A(\g.we_clk [10907]));
Q_ASSIGN U21868 ( .B(clk), .A(\g.we_clk [10906]));
Q_ASSIGN U21869 ( .B(clk), .A(\g.we_clk [10905]));
Q_ASSIGN U21870 ( .B(clk), .A(\g.we_clk [10904]));
Q_ASSIGN U21871 ( .B(clk), .A(\g.we_clk [10903]));
Q_ASSIGN U21872 ( .B(clk), .A(\g.we_clk [10902]));
Q_ASSIGN U21873 ( .B(clk), .A(\g.we_clk [10901]));
Q_ASSIGN U21874 ( .B(clk), .A(\g.we_clk [10900]));
Q_ASSIGN U21875 ( .B(clk), .A(\g.we_clk [10899]));
Q_ASSIGN U21876 ( .B(clk), .A(\g.we_clk [10898]));
Q_ASSIGN U21877 ( .B(clk), .A(\g.we_clk [10897]));
Q_ASSIGN U21878 ( .B(clk), .A(\g.we_clk [10896]));
Q_ASSIGN U21879 ( .B(clk), .A(\g.we_clk [10895]));
Q_ASSIGN U21880 ( .B(clk), .A(\g.we_clk [10894]));
Q_ASSIGN U21881 ( .B(clk), .A(\g.we_clk [10893]));
Q_ASSIGN U21882 ( .B(clk), .A(\g.we_clk [10892]));
Q_ASSIGN U21883 ( .B(clk), .A(\g.we_clk [10891]));
Q_ASSIGN U21884 ( .B(clk), .A(\g.we_clk [10890]));
Q_ASSIGN U21885 ( .B(clk), .A(\g.we_clk [10889]));
Q_ASSIGN U21886 ( .B(clk), .A(\g.we_clk [10888]));
Q_ASSIGN U21887 ( .B(clk), .A(\g.we_clk [10887]));
Q_ASSIGN U21888 ( .B(clk), .A(\g.we_clk [10886]));
Q_ASSIGN U21889 ( .B(clk), .A(\g.we_clk [10885]));
Q_ASSIGN U21890 ( .B(clk), .A(\g.we_clk [10884]));
Q_ASSIGN U21891 ( .B(clk), .A(\g.we_clk [10883]));
Q_ASSIGN U21892 ( .B(clk), .A(\g.we_clk [10882]));
Q_ASSIGN U21893 ( .B(clk), .A(\g.we_clk [10881]));
Q_ASSIGN U21894 ( .B(clk), .A(\g.we_clk [10880]));
Q_ASSIGN U21895 ( .B(clk), .A(\g.we_clk [10879]));
Q_ASSIGN U21896 ( .B(clk), .A(\g.we_clk [10878]));
Q_ASSIGN U21897 ( .B(clk), .A(\g.we_clk [10877]));
Q_ASSIGN U21898 ( .B(clk), .A(\g.we_clk [10876]));
Q_ASSIGN U21899 ( .B(clk), .A(\g.we_clk [10875]));
Q_ASSIGN U21900 ( .B(clk), .A(\g.we_clk [10874]));
Q_ASSIGN U21901 ( .B(clk), .A(\g.we_clk [10873]));
Q_ASSIGN U21902 ( .B(clk), .A(\g.we_clk [10872]));
Q_ASSIGN U21903 ( .B(clk), .A(\g.we_clk [10871]));
Q_ASSIGN U21904 ( .B(clk), .A(\g.we_clk [10870]));
Q_ASSIGN U21905 ( .B(clk), .A(\g.we_clk [10869]));
Q_ASSIGN U21906 ( .B(clk), .A(\g.we_clk [10868]));
Q_ASSIGN U21907 ( .B(clk), .A(\g.we_clk [10867]));
Q_ASSIGN U21908 ( .B(clk), .A(\g.we_clk [10866]));
Q_ASSIGN U21909 ( .B(clk), .A(\g.we_clk [10865]));
Q_ASSIGN U21910 ( .B(clk), .A(\g.we_clk [10864]));
Q_ASSIGN U21911 ( .B(clk), .A(\g.we_clk [10863]));
Q_ASSIGN U21912 ( .B(clk), .A(\g.we_clk [10862]));
Q_ASSIGN U21913 ( .B(clk), .A(\g.we_clk [10861]));
Q_ASSIGN U21914 ( .B(clk), .A(\g.we_clk [10860]));
Q_ASSIGN U21915 ( .B(clk), .A(\g.we_clk [10859]));
Q_ASSIGN U21916 ( .B(clk), .A(\g.we_clk [10858]));
Q_ASSIGN U21917 ( .B(clk), .A(\g.we_clk [10857]));
Q_ASSIGN U21918 ( .B(clk), .A(\g.we_clk [10856]));
Q_ASSIGN U21919 ( .B(clk), .A(\g.we_clk [10855]));
Q_ASSIGN U21920 ( .B(clk), .A(\g.we_clk [10854]));
Q_ASSIGN U21921 ( .B(clk), .A(\g.we_clk [10853]));
Q_ASSIGN U21922 ( .B(clk), .A(\g.we_clk [10852]));
Q_ASSIGN U21923 ( .B(clk), .A(\g.we_clk [10851]));
Q_ASSIGN U21924 ( .B(clk), .A(\g.we_clk [10850]));
Q_ASSIGN U21925 ( .B(clk), .A(\g.we_clk [10849]));
Q_ASSIGN U21926 ( .B(clk), .A(\g.we_clk [10848]));
Q_ASSIGN U21927 ( .B(clk), .A(\g.we_clk [10847]));
Q_ASSIGN U21928 ( .B(clk), .A(\g.we_clk [10846]));
Q_ASSIGN U21929 ( .B(clk), .A(\g.we_clk [10845]));
Q_ASSIGN U21930 ( .B(clk), .A(\g.we_clk [10844]));
Q_ASSIGN U21931 ( .B(clk), .A(\g.we_clk [10843]));
Q_ASSIGN U21932 ( .B(clk), .A(\g.we_clk [10842]));
Q_ASSIGN U21933 ( .B(clk), .A(\g.we_clk [10841]));
Q_ASSIGN U21934 ( .B(clk), .A(\g.we_clk [10840]));
Q_ASSIGN U21935 ( .B(clk), .A(\g.we_clk [10839]));
Q_ASSIGN U21936 ( .B(clk), .A(\g.we_clk [10838]));
Q_ASSIGN U21937 ( .B(clk), .A(\g.we_clk [10837]));
Q_ASSIGN U21938 ( .B(clk), .A(\g.we_clk [10836]));
Q_ASSIGN U21939 ( .B(clk), .A(\g.we_clk [10835]));
Q_ASSIGN U21940 ( .B(clk), .A(\g.we_clk [10834]));
Q_ASSIGN U21941 ( .B(clk), .A(\g.we_clk [10833]));
Q_ASSIGN U21942 ( .B(clk), .A(\g.we_clk [10832]));
Q_ASSIGN U21943 ( .B(clk), .A(\g.we_clk [10831]));
Q_ASSIGN U21944 ( .B(clk), .A(\g.we_clk [10830]));
Q_ASSIGN U21945 ( .B(clk), .A(\g.we_clk [10829]));
Q_ASSIGN U21946 ( .B(clk), .A(\g.we_clk [10828]));
Q_ASSIGN U21947 ( .B(clk), .A(\g.we_clk [10827]));
Q_ASSIGN U21948 ( .B(clk), .A(\g.we_clk [10826]));
Q_ASSIGN U21949 ( .B(clk), .A(\g.we_clk [10825]));
Q_ASSIGN U21950 ( .B(clk), .A(\g.we_clk [10824]));
Q_ASSIGN U21951 ( .B(clk), .A(\g.we_clk [10823]));
Q_ASSIGN U21952 ( .B(clk), .A(\g.we_clk [10822]));
Q_ASSIGN U21953 ( .B(clk), .A(\g.we_clk [10821]));
Q_ASSIGN U21954 ( .B(clk), .A(\g.we_clk [10820]));
Q_ASSIGN U21955 ( .B(clk), .A(\g.we_clk [10819]));
Q_ASSIGN U21956 ( .B(clk), .A(\g.we_clk [10818]));
Q_ASSIGN U21957 ( .B(clk), .A(\g.we_clk [10817]));
Q_ASSIGN U21958 ( .B(clk), .A(\g.we_clk [10816]));
Q_ASSIGN U21959 ( .B(clk), .A(\g.we_clk [10815]));
Q_ASSIGN U21960 ( .B(clk), .A(\g.we_clk [10814]));
Q_ASSIGN U21961 ( .B(clk), .A(\g.we_clk [10813]));
Q_ASSIGN U21962 ( .B(clk), .A(\g.we_clk [10812]));
Q_ASSIGN U21963 ( .B(clk), .A(\g.we_clk [10811]));
Q_ASSIGN U21964 ( .B(clk), .A(\g.we_clk [10810]));
Q_ASSIGN U21965 ( .B(clk), .A(\g.we_clk [10809]));
Q_ASSIGN U21966 ( .B(clk), .A(\g.we_clk [10808]));
Q_ASSIGN U21967 ( .B(clk), .A(\g.we_clk [10807]));
Q_ASSIGN U21968 ( .B(clk), .A(\g.we_clk [10806]));
Q_ASSIGN U21969 ( .B(clk), .A(\g.we_clk [10805]));
Q_ASSIGN U21970 ( .B(clk), .A(\g.we_clk [10804]));
Q_ASSIGN U21971 ( .B(clk), .A(\g.we_clk [10803]));
Q_ASSIGN U21972 ( .B(clk), .A(\g.we_clk [10802]));
Q_ASSIGN U21973 ( .B(clk), .A(\g.we_clk [10801]));
Q_ASSIGN U21974 ( .B(clk), .A(\g.we_clk [10800]));
Q_ASSIGN U21975 ( .B(clk), .A(\g.we_clk [10799]));
Q_ASSIGN U21976 ( .B(clk), .A(\g.we_clk [10798]));
Q_ASSIGN U21977 ( .B(clk), .A(\g.we_clk [10797]));
Q_ASSIGN U21978 ( .B(clk), .A(\g.we_clk [10796]));
Q_ASSIGN U21979 ( .B(clk), .A(\g.we_clk [10795]));
Q_ASSIGN U21980 ( .B(clk), .A(\g.we_clk [10794]));
Q_ASSIGN U21981 ( .B(clk), .A(\g.we_clk [10793]));
Q_ASSIGN U21982 ( .B(clk), .A(\g.we_clk [10792]));
Q_ASSIGN U21983 ( .B(clk), .A(\g.we_clk [10791]));
Q_ASSIGN U21984 ( .B(clk), .A(\g.we_clk [10790]));
Q_ASSIGN U21985 ( .B(clk), .A(\g.we_clk [10789]));
Q_ASSIGN U21986 ( .B(clk), .A(\g.we_clk [10788]));
Q_ASSIGN U21987 ( .B(clk), .A(\g.we_clk [10787]));
Q_ASSIGN U21988 ( .B(clk), .A(\g.we_clk [10786]));
Q_ASSIGN U21989 ( .B(clk), .A(\g.we_clk [10785]));
Q_ASSIGN U21990 ( .B(clk), .A(\g.we_clk [10784]));
Q_ASSIGN U21991 ( .B(clk), .A(\g.we_clk [10783]));
Q_ASSIGN U21992 ( .B(clk), .A(\g.we_clk [10782]));
Q_ASSIGN U21993 ( .B(clk), .A(\g.we_clk [10781]));
Q_ASSIGN U21994 ( .B(clk), .A(\g.we_clk [10780]));
Q_ASSIGN U21995 ( .B(clk), .A(\g.we_clk [10779]));
Q_ASSIGN U21996 ( .B(clk), .A(\g.we_clk [10778]));
Q_ASSIGN U21997 ( .B(clk), .A(\g.we_clk [10777]));
Q_ASSIGN U21998 ( .B(clk), .A(\g.we_clk [10776]));
Q_ASSIGN U21999 ( .B(clk), .A(\g.we_clk [10775]));
Q_ASSIGN U22000 ( .B(clk), .A(\g.we_clk [10774]));
Q_ASSIGN U22001 ( .B(clk), .A(\g.we_clk [10773]));
Q_ASSIGN U22002 ( .B(clk), .A(\g.we_clk [10772]));
Q_ASSIGN U22003 ( .B(clk), .A(\g.we_clk [10771]));
Q_ASSIGN U22004 ( .B(clk), .A(\g.we_clk [10770]));
Q_ASSIGN U22005 ( .B(clk), .A(\g.we_clk [10769]));
Q_ASSIGN U22006 ( .B(clk), .A(\g.we_clk [10768]));
Q_ASSIGN U22007 ( .B(clk), .A(\g.we_clk [10767]));
Q_ASSIGN U22008 ( .B(clk), .A(\g.we_clk [10766]));
Q_ASSIGN U22009 ( .B(clk), .A(\g.we_clk [10765]));
Q_ASSIGN U22010 ( .B(clk), .A(\g.we_clk [10764]));
Q_ASSIGN U22011 ( .B(clk), .A(\g.we_clk [10763]));
Q_ASSIGN U22012 ( .B(clk), .A(\g.we_clk [10762]));
Q_ASSIGN U22013 ( .B(clk), .A(\g.we_clk [10761]));
Q_ASSIGN U22014 ( .B(clk), .A(\g.we_clk [10760]));
Q_ASSIGN U22015 ( .B(clk), .A(\g.we_clk [10759]));
Q_ASSIGN U22016 ( .B(clk), .A(\g.we_clk [10758]));
Q_ASSIGN U22017 ( .B(clk), .A(\g.we_clk [10757]));
Q_ASSIGN U22018 ( .B(clk), .A(\g.we_clk [10756]));
Q_ASSIGN U22019 ( .B(clk), .A(\g.we_clk [10755]));
Q_ASSIGN U22020 ( .B(clk), .A(\g.we_clk [10754]));
Q_ASSIGN U22021 ( .B(clk), .A(\g.we_clk [10753]));
Q_ASSIGN U22022 ( .B(clk), .A(\g.we_clk [10752]));
Q_ASSIGN U22023 ( .B(clk), .A(\g.we_clk [10751]));
Q_ASSIGN U22024 ( .B(clk), .A(\g.we_clk [10750]));
Q_ASSIGN U22025 ( .B(clk), .A(\g.we_clk [10749]));
Q_ASSIGN U22026 ( .B(clk), .A(\g.we_clk [10748]));
Q_ASSIGN U22027 ( .B(clk), .A(\g.we_clk [10747]));
Q_ASSIGN U22028 ( .B(clk), .A(\g.we_clk [10746]));
Q_ASSIGN U22029 ( .B(clk), .A(\g.we_clk [10745]));
Q_ASSIGN U22030 ( .B(clk), .A(\g.we_clk [10744]));
Q_ASSIGN U22031 ( .B(clk), .A(\g.we_clk [10743]));
Q_ASSIGN U22032 ( .B(clk), .A(\g.we_clk [10742]));
Q_ASSIGN U22033 ( .B(clk), .A(\g.we_clk [10741]));
Q_ASSIGN U22034 ( .B(clk), .A(\g.we_clk [10740]));
Q_ASSIGN U22035 ( .B(clk), .A(\g.we_clk [10739]));
Q_ASSIGN U22036 ( .B(clk), .A(\g.we_clk [10738]));
Q_ASSIGN U22037 ( .B(clk), .A(\g.we_clk [10737]));
Q_ASSIGN U22038 ( .B(clk), .A(\g.we_clk [10736]));
Q_ASSIGN U22039 ( .B(clk), .A(\g.we_clk [10735]));
Q_ASSIGN U22040 ( .B(clk), .A(\g.we_clk [10734]));
Q_ASSIGN U22041 ( .B(clk), .A(\g.we_clk [10733]));
Q_ASSIGN U22042 ( .B(clk), .A(\g.we_clk [10732]));
Q_ASSIGN U22043 ( .B(clk), .A(\g.we_clk [10731]));
Q_ASSIGN U22044 ( .B(clk), .A(\g.we_clk [10730]));
Q_ASSIGN U22045 ( .B(clk), .A(\g.we_clk [10729]));
Q_ASSIGN U22046 ( .B(clk), .A(\g.we_clk [10728]));
Q_ASSIGN U22047 ( .B(clk), .A(\g.we_clk [10727]));
Q_ASSIGN U22048 ( .B(clk), .A(\g.we_clk [10726]));
Q_ASSIGN U22049 ( .B(clk), .A(\g.we_clk [10725]));
Q_ASSIGN U22050 ( .B(clk), .A(\g.we_clk [10724]));
Q_ASSIGN U22051 ( .B(clk), .A(\g.we_clk [10723]));
Q_ASSIGN U22052 ( .B(clk), .A(\g.we_clk [10722]));
Q_ASSIGN U22053 ( .B(clk), .A(\g.we_clk [10721]));
Q_ASSIGN U22054 ( .B(clk), .A(\g.we_clk [10720]));
Q_ASSIGN U22055 ( .B(clk), .A(\g.we_clk [10719]));
Q_ASSIGN U22056 ( .B(clk), .A(\g.we_clk [10718]));
Q_ASSIGN U22057 ( .B(clk), .A(\g.we_clk [10717]));
Q_ASSIGN U22058 ( .B(clk), .A(\g.we_clk [10716]));
Q_ASSIGN U22059 ( .B(clk), .A(\g.we_clk [10715]));
Q_ASSIGN U22060 ( .B(clk), .A(\g.we_clk [10714]));
Q_ASSIGN U22061 ( .B(clk), .A(\g.we_clk [10713]));
Q_ASSIGN U22062 ( .B(clk), .A(\g.we_clk [10712]));
Q_ASSIGN U22063 ( .B(clk), .A(\g.we_clk [10711]));
Q_ASSIGN U22064 ( .B(clk), .A(\g.we_clk [10710]));
Q_ASSIGN U22065 ( .B(clk), .A(\g.we_clk [10709]));
Q_ASSIGN U22066 ( .B(clk), .A(\g.we_clk [10708]));
Q_ASSIGN U22067 ( .B(clk), .A(\g.we_clk [10707]));
Q_ASSIGN U22068 ( .B(clk), .A(\g.we_clk [10706]));
Q_ASSIGN U22069 ( .B(clk), .A(\g.we_clk [10705]));
Q_ASSIGN U22070 ( .B(clk), .A(\g.we_clk [10704]));
Q_ASSIGN U22071 ( .B(clk), .A(\g.we_clk [10703]));
Q_ASSIGN U22072 ( .B(clk), .A(\g.we_clk [10702]));
Q_ASSIGN U22073 ( .B(clk), .A(\g.we_clk [10701]));
Q_ASSIGN U22074 ( .B(clk), .A(\g.we_clk [10700]));
Q_ASSIGN U22075 ( .B(clk), .A(\g.we_clk [10699]));
Q_ASSIGN U22076 ( .B(clk), .A(\g.we_clk [10698]));
Q_ASSIGN U22077 ( .B(clk), .A(\g.we_clk [10697]));
Q_ASSIGN U22078 ( .B(clk), .A(\g.we_clk [10696]));
Q_ASSIGN U22079 ( .B(clk), .A(\g.we_clk [10695]));
Q_ASSIGN U22080 ( .B(clk), .A(\g.we_clk [10694]));
Q_ASSIGN U22081 ( .B(clk), .A(\g.we_clk [10693]));
Q_ASSIGN U22082 ( .B(clk), .A(\g.we_clk [10692]));
Q_ASSIGN U22083 ( .B(clk), .A(\g.we_clk [10691]));
Q_ASSIGN U22084 ( .B(clk), .A(\g.we_clk [10690]));
Q_ASSIGN U22085 ( .B(clk), .A(\g.we_clk [10689]));
Q_ASSIGN U22086 ( .B(clk), .A(\g.we_clk [10688]));
Q_ASSIGN U22087 ( .B(clk), .A(\g.we_clk [10687]));
Q_ASSIGN U22088 ( .B(clk), .A(\g.we_clk [10686]));
Q_ASSIGN U22089 ( .B(clk), .A(\g.we_clk [10685]));
Q_ASSIGN U22090 ( .B(clk), .A(\g.we_clk [10684]));
Q_ASSIGN U22091 ( .B(clk), .A(\g.we_clk [10683]));
Q_ASSIGN U22092 ( .B(clk), .A(\g.we_clk [10682]));
Q_ASSIGN U22093 ( .B(clk), .A(\g.we_clk [10681]));
Q_ASSIGN U22094 ( .B(clk), .A(\g.we_clk [10680]));
Q_ASSIGN U22095 ( .B(clk), .A(\g.we_clk [10679]));
Q_ASSIGN U22096 ( .B(clk), .A(\g.we_clk [10678]));
Q_ASSIGN U22097 ( .B(clk), .A(\g.we_clk [10677]));
Q_ASSIGN U22098 ( .B(clk), .A(\g.we_clk [10676]));
Q_ASSIGN U22099 ( .B(clk), .A(\g.we_clk [10675]));
Q_ASSIGN U22100 ( .B(clk), .A(\g.we_clk [10674]));
Q_ASSIGN U22101 ( .B(clk), .A(\g.we_clk [10673]));
Q_ASSIGN U22102 ( .B(clk), .A(\g.we_clk [10672]));
Q_ASSIGN U22103 ( .B(clk), .A(\g.we_clk [10671]));
Q_ASSIGN U22104 ( .B(clk), .A(\g.we_clk [10670]));
Q_ASSIGN U22105 ( .B(clk), .A(\g.we_clk [10669]));
Q_ASSIGN U22106 ( .B(clk), .A(\g.we_clk [10668]));
Q_ASSIGN U22107 ( .B(clk), .A(\g.we_clk [10667]));
Q_ASSIGN U22108 ( .B(clk), .A(\g.we_clk [10666]));
Q_ASSIGN U22109 ( .B(clk), .A(\g.we_clk [10665]));
Q_ASSIGN U22110 ( .B(clk), .A(\g.we_clk [10664]));
Q_ASSIGN U22111 ( .B(clk), .A(\g.we_clk [10663]));
Q_ASSIGN U22112 ( .B(clk), .A(\g.we_clk [10662]));
Q_ASSIGN U22113 ( .B(clk), .A(\g.we_clk [10661]));
Q_ASSIGN U22114 ( .B(clk), .A(\g.we_clk [10660]));
Q_ASSIGN U22115 ( .B(clk), .A(\g.we_clk [10659]));
Q_ASSIGN U22116 ( .B(clk), .A(\g.we_clk [10658]));
Q_ASSIGN U22117 ( .B(clk), .A(\g.we_clk [10657]));
Q_ASSIGN U22118 ( .B(clk), .A(\g.we_clk [10656]));
Q_ASSIGN U22119 ( .B(clk), .A(\g.we_clk [10655]));
Q_ASSIGN U22120 ( .B(clk), .A(\g.we_clk [10654]));
Q_ASSIGN U22121 ( .B(clk), .A(\g.we_clk [10653]));
Q_ASSIGN U22122 ( .B(clk), .A(\g.we_clk [10652]));
Q_ASSIGN U22123 ( .B(clk), .A(\g.we_clk [10651]));
Q_ASSIGN U22124 ( .B(clk), .A(\g.we_clk [10650]));
Q_ASSIGN U22125 ( .B(clk), .A(\g.we_clk [10649]));
Q_ASSIGN U22126 ( .B(clk), .A(\g.we_clk [10648]));
Q_ASSIGN U22127 ( .B(clk), .A(\g.we_clk [10647]));
Q_ASSIGN U22128 ( .B(clk), .A(\g.we_clk [10646]));
Q_ASSIGN U22129 ( .B(clk), .A(\g.we_clk [10645]));
Q_ASSIGN U22130 ( .B(clk), .A(\g.we_clk [10644]));
Q_ASSIGN U22131 ( .B(clk), .A(\g.we_clk [10643]));
Q_ASSIGN U22132 ( .B(clk), .A(\g.we_clk [10642]));
Q_ASSIGN U22133 ( .B(clk), .A(\g.we_clk [10641]));
Q_ASSIGN U22134 ( .B(clk), .A(\g.we_clk [10640]));
Q_ASSIGN U22135 ( .B(clk), .A(\g.we_clk [10639]));
Q_ASSIGN U22136 ( .B(clk), .A(\g.we_clk [10638]));
Q_ASSIGN U22137 ( .B(clk), .A(\g.we_clk [10637]));
Q_ASSIGN U22138 ( .B(clk), .A(\g.we_clk [10636]));
Q_ASSIGN U22139 ( .B(clk), .A(\g.we_clk [10635]));
Q_ASSIGN U22140 ( .B(clk), .A(\g.we_clk [10634]));
Q_ASSIGN U22141 ( .B(clk), .A(\g.we_clk [10633]));
Q_ASSIGN U22142 ( .B(clk), .A(\g.we_clk [10632]));
Q_ASSIGN U22143 ( .B(clk), .A(\g.we_clk [10631]));
Q_ASSIGN U22144 ( .B(clk), .A(\g.we_clk [10630]));
Q_ASSIGN U22145 ( .B(clk), .A(\g.we_clk [10629]));
Q_ASSIGN U22146 ( .B(clk), .A(\g.we_clk [10628]));
Q_ASSIGN U22147 ( .B(clk), .A(\g.we_clk [10627]));
Q_ASSIGN U22148 ( .B(clk), .A(\g.we_clk [10626]));
Q_ASSIGN U22149 ( .B(clk), .A(\g.we_clk [10625]));
Q_ASSIGN U22150 ( .B(clk), .A(\g.we_clk [10624]));
Q_ASSIGN U22151 ( .B(clk), .A(\g.we_clk [10623]));
Q_ASSIGN U22152 ( .B(clk), .A(\g.we_clk [10622]));
Q_ASSIGN U22153 ( .B(clk), .A(\g.we_clk [10621]));
Q_ASSIGN U22154 ( .B(clk), .A(\g.we_clk [10620]));
Q_ASSIGN U22155 ( .B(clk), .A(\g.we_clk [10619]));
Q_ASSIGN U22156 ( .B(clk), .A(\g.we_clk [10618]));
Q_ASSIGN U22157 ( .B(clk), .A(\g.we_clk [10617]));
Q_ASSIGN U22158 ( .B(clk), .A(\g.we_clk [10616]));
Q_ASSIGN U22159 ( .B(clk), .A(\g.we_clk [10615]));
Q_ASSIGN U22160 ( .B(clk), .A(\g.we_clk [10614]));
Q_ASSIGN U22161 ( .B(clk), .A(\g.we_clk [10613]));
Q_ASSIGN U22162 ( .B(clk), .A(\g.we_clk [10612]));
Q_ASSIGN U22163 ( .B(clk), .A(\g.we_clk [10611]));
Q_ASSIGN U22164 ( .B(clk), .A(\g.we_clk [10610]));
Q_ASSIGN U22165 ( .B(clk), .A(\g.we_clk [10609]));
Q_ASSIGN U22166 ( .B(clk), .A(\g.we_clk [10608]));
Q_ASSIGN U22167 ( .B(clk), .A(\g.we_clk [10607]));
Q_ASSIGN U22168 ( .B(clk), .A(\g.we_clk [10606]));
Q_ASSIGN U22169 ( .B(clk), .A(\g.we_clk [10605]));
Q_ASSIGN U22170 ( .B(clk), .A(\g.we_clk [10604]));
Q_ASSIGN U22171 ( .B(clk), .A(\g.we_clk [10603]));
Q_ASSIGN U22172 ( .B(clk), .A(\g.we_clk [10602]));
Q_ASSIGN U22173 ( .B(clk), .A(\g.we_clk [10601]));
Q_ASSIGN U22174 ( .B(clk), .A(\g.we_clk [10600]));
Q_ASSIGN U22175 ( .B(clk), .A(\g.we_clk [10599]));
Q_ASSIGN U22176 ( .B(clk), .A(\g.we_clk [10598]));
Q_ASSIGN U22177 ( .B(clk), .A(\g.we_clk [10597]));
Q_ASSIGN U22178 ( .B(clk), .A(\g.we_clk [10596]));
Q_ASSIGN U22179 ( .B(clk), .A(\g.we_clk [10595]));
Q_ASSIGN U22180 ( .B(clk), .A(\g.we_clk [10594]));
Q_ASSIGN U22181 ( .B(clk), .A(\g.we_clk [10593]));
Q_ASSIGN U22182 ( .B(clk), .A(\g.we_clk [10592]));
Q_ASSIGN U22183 ( .B(clk), .A(\g.we_clk [10591]));
Q_ASSIGN U22184 ( .B(clk), .A(\g.we_clk [10590]));
Q_ASSIGN U22185 ( .B(clk), .A(\g.we_clk [10589]));
Q_ASSIGN U22186 ( .B(clk), .A(\g.we_clk [10588]));
Q_ASSIGN U22187 ( .B(clk), .A(\g.we_clk [10587]));
Q_ASSIGN U22188 ( .B(clk), .A(\g.we_clk [10586]));
Q_ASSIGN U22189 ( .B(clk), .A(\g.we_clk [10585]));
Q_ASSIGN U22190 ( .B(clk), .A(\g.we_clk [10584]));
Q_ASSIGN U22191 ( .B(clk), .A(\g.we_clk [10583]));
Q_ASSIGN U22192 ( .B(clk), .A(\g.we_clk [10582]));
Q_ASSIGN U22193 ( .B(clk), .A(\g.we_clk [10581]));
Q_ASSIGN U22194 ( .B(clk), .A(\g.we_clk [10580]));
Q_ASSIGN U22195 ( .B(clk), .A(\g.we_clk [10579]));
Q_ASSIGN U22196 ( .B(clk), .A(\g.we_clk [10578]));
Q_ASSIGN U22197 ( .B(clk), .A(\g.we_clk [10577]));
Q_ASSIGN U22198 ( .B(clk), .A(\g.we_clk [10576]));
Q_ASSIGN U22199 ( .B(clk), .A(\g.we_clk [10575]));
Q_ASSIGN U22200 ( .B(clk), .A(\g.we_clk [10574]));
Q_ASSIGN U22201 ( .B(clk), .A(\g.we_clk [10573]));
Q_ASSIGN U22202 ( .B(clk), .A(\g.we_clk [10572]));
Q_ASSIGN U22203 ( .B(clk), .A(\g.we_clk [10571]));
Q_ASSIGN U22204 ( .B(clk), .A(\g.we_clk [10570]));
Q_ASSIGN U22205 ( .B(clk), .A(\g.we_clk [10569]));
Q_ASSIGN U22206 ( .B(clk), .A(\g.we_clk [10568]));
Q_ASSIGN U22207 ( .B(clk), .A(\g.we_clk [10567]));
Q_ASSIGN U22208 ( .B(clk), .A(\g.we_clk [10566]));
Q_ASSIGN U22209 ( .B(clk), .A(\g.we_clk [10565]));
Q_ASSIGN U22210 ( .B(clk), .A(\g.we_clk [10564]));
Q_ASSIGN U22211 ( .B(clk), .A(\g.we_clk [10563]));
Q_ASSIGN U22212 ( .B(clk), .A(\g.we_clk [10562]));
Q_ASSIGN U22213 ( .B(clk), .A(\g.we_clk [10561]));
Q_ASSIGN U22214 ( .B(clk), .A(\g.we_clk [10560]));
Q_ASSIGN U22215 ( .B(clk), .A(\g.we_clk [10559]));
Q_ASSIGN U22216 ( .B(clk), .A(\g.we_clk [10558]));
Q_ASSIGN U22217 ( .B(clk), .A(\g.we_clk [10557]));
Q_ASSIGN U22218 ( .B(clk), .A(\g.we_clk [10556]));
Q_ASSIGN U22219 ( .B(clk), .A(\g.we_clk [10555]));
Q_ASSIGN U22220 ( .B(clk), .A(\g.we_clk [10554]));
Q_ASSIGN U22221 ( .B(clk), .A(\g.we_clk [10553]));
Q_ASSIGN U22222 ( .B(clk), .A(\g.we_clk [10552]));
Q_ASSIGN U22223 ( .B(clk), .A(\g.we_clk [10551]));
Q_ASSIGN U22224 ( .B(clk), .A(\g.we_clk [10550]));
Q_ASSIGN U22225 ( .B(clk), .A(\g.we_clk [10549]));
Q_ASSIGN U22226 ( .B(clk), .A(\g.we_clk [10548]));
Q_ASSIGN U22227 ( .B(clk), .A(\g.we_clk [10547]));
Q_ASSIGN U22228 ( .B(clk), .A(\g.we_clk [10546]));
Q_ASSIGN U22229 ( .B(clk), .A(\g.we_clk [10545]));
Q_ASSIGN U22230 ( .B(clk), .A(\g.we_clk [10544]));
Q_ASSIGN U22231 ( .B(clk), .A(\g.we_clk [10543]));
Q_ASSIGN U22232 ( .B(clk), .A(\g.we_clk [10542]));
Q_ASSIGN U22233 ( .B(clk), .A(\g.we_clk [10541]));
Q_ASSIGN U22234 ( .B(clk), .A(\g.we_clk [10540]));
Q_ASSIGN U22235 ( .B(clk), .A(\g.we_clk [10539]));
Q_ASSIGN U22236 ( .B(clk), .A(\g.we_clk [10538]));
Q_ASSIGN U22237 ( .B(clk), .A(\g.we_clk [10537]));
Q_ASSIGN U22238 ( .B(clk), .A(\g.we_clk [10536]));
Q_ASSIGN U22239 ( .B(clk), .A(\g.we_clk [10535]));
Q_ASSIGN U22240 ( .B(clk), .A(\g.we_clk [10534]));
Q_ASSIGN U22241 ( .B(clk), .A(\g.we_clk [10533]));
Q_ASSIGN U22242 ( .B(clk), .A(\g.we_clk [10532]));
Q_ASSIGN U22243 ( .B(clk), .A(\g.we_clk [10531]));
Q_ASSIGN U22244 ( .B(clk), .A(\g.we_clk [10530]));
Q_ASSIGN U22245 ( .B(clk), .A(\g.we_clk [10529]));
Q_ASSIGN U22246 ( .B(clk), .A(\g.we_clk [10528]));
Q_ASSIGN U22247 ( .B(clk), .A(\g.we_clk [10527]));
Q_ASSIGN U22248 ( .B(clk), .A(\g.we_clk [10526]));
Q_ASSIGN U22249 ( .B(clk), .A(\g.we_clk [10525]));
Q_ASSIGN U22250 ( .B(clk), .A(\g.we_clk [10524]));
Q_ASSIGN U22251 ( .B(clk), .A(\g.we_clk [10523]));
Q_ASSIGN U22252 ( .B(clk), .A(\g.we_clk [10522]));
Q_ASSIGN U22253 ( .B(clk), .A(\g.we_clk [10521]));
Q_ASSIGN U22254 ( .B(clk), .A(\g.we_clk [10520]));
Q_ASSIGN U22255 ( .B(clk), .A(\g.we_clk [10519]));
Q_ASSIGN U22256 ( .B(clk), .A(\g.we_clk [10518]));
Q_ASSIGN U22257 ( .B(clk), .A(\g.we_clk [10517]));
Q_ASSIGN U22258 ( .B(clk), .A(\g.we_clk [10516]));
Q_ASSIGN U22259 ( .B(clk), .A(\g.we_clk [10515]));
Q_ASSIGN U22260 ( .B(clk), .A(\g.we_clk [10514]));
Q_ASSIGN U22261 ( .B(clk), .A(\g.we_clk [10513]));
Q_ASSIGN U22262 ( .B(clk), .A(\g.we_clk [10512]));
Q_ASSIGN U22263 ( .B(clk), .A(\g.we_clk [10511]));
Q_ASSIGN U22264 ( .B(clk), .A(\g.we_clk [10510]));
Q_ASSIGN U22265 ( .B(clk), .A(\g.we_clk [10509]));
Q_ASSIGN U22266 ( .B(clk), .A(\g.we_clk [10508]));
Q_ASSIGN U22267 ( .B(clk), .A(\g.we_clk [10507]));
Q_ASSIGN U22268 ( .B(clk), .A(\g.we_clk [10506]));
Q_ASSIGN U22269 ( .B(clk), .A(\g.we_clk [10505]));
Q_ASSIGN U22270 ( .B(clk), .A(\g.we_clk [10504]));
Q_ASSIGN U22271 ( .B(clk), .A(\g.we_clk [10503]));
Q_ASSIGN U22272 ( .B(clk), .A(\g.we_clk [10502]));
Q_ASSIGN U22273 ( .B(clk), .A(\g.we_clk [10501]));
Q_ASSIGN U22274 ( .B(clk), .A(\g.we_clk [10500]));
Q_ASSIGN U22275 ( .B(clk), .A(\g.we_clk [10499]));
Q_ASSIGN U22276 ( .B(clk), .A(\g.we_clk [10498]));
Q_ASSIGN U22277 ( .B(clk), .A(\g.we_clk [10497]));
Q_ASSIGN U22278 ( .B(clk), .A(\g.we_clk [10496]));
Q_ASSIGN U22279 ( .B(clk), .A(\g.we_clk [10495]));
Q_ASSIGN U22280 ( .B(clk), .A(\g.we_clk [10494]));
Q_ASSIGN U22281 ( .B(clk), .A(\g.we_clk [10493]));
Q_ASSIGN U22282 ( .B(clk), .A(\g.we_clk [10492]));
Q_ASSIGN U22283 ( .B(clk), .A(\g.we_clk [10491]));
Q_ASSIGN U22284 ( .B(clk), .A(\g.we_clk [10490]));
Q_ASSIGN U22285 ( .B(clk), .A(\g.we_clk [10489]));
Q_ASSIGN U22286 ( .B(clk), .A(\g.we_clk [10488]));
Q_ASSIGN U22287 ( .B(clk), .A(\g.we_clk [10487]));
Q_ASSIGN U22288 ( .B(clk), .A(\g.we_clk [10486]));
Q_ASSIGN U22289 ( .B(clk), .A(\g.we_clk [10485]));
Q_ASSIGN U22290 ( .B(clk), .A(\g.we_clk [10484]));
Q_ASSIGN U22291 ( .B(clk), .A(\g.we_clk [10483]));
Q_ASSIGN U22292 ( .B(clk), .A(\g.we_clk [10482]));
Q_ASSIGN U22293 ( .B(clk), .A(\g.we_clk [10481]));
Q_ASSIGN U22294 ( .B(clk), .A(\g.we_clk [10480]));
Q_ASSIGN U22295 ( .B(clk), .A(\g.we_clk [10479]));
Q_ASSIGN U22296 ( .B(clk), .A(\g.we_clk [10478]));
Q_ASSIGN U22297 ( .B(clk), .A(\g.we_clk [10477]));
Q_ASSIGN U22298 ( .B(clk), .A(\g.we_clk [10476]));
Q_ASSIGN U22299 ( .B(clk), .A(\g.we_clk [10475]));
Q_ASSIGN U22300 ( .B(clk), .A(\g.we_clk [10474]));
Q_ASSIGN U22301 ( .B(clk), .A(\g.we_clk [10473]));
Q_ASSIGN U22302 ( .B(clk), .A(\g.we_clk [10472]));
Q_ASSIGN U22303 ( .B(clk), .A(\g.we_clk [10471]));
Q_ASSIGN U22304 ( .B(clk), .A(\g.we_clk [10470]));
Q_ASSIGN U22305 ( .B(clk), .A(\g.we_clk [10469]));
Q_ASSIGN U22306 ( .B(clk), .A(\g.we_clk [10468]));
Q_ASSIGN U22307 ( .B(clk), .A(\g.we_clk [10467]));
Q_ASSIGN U22308 ( .B(clk), .A(\g.we_clk [10466]));
Q_ASSIGN U22309 ( .B(clk), .A(\g.we_clk [10465]));
Q_ASSIGN U22310 ( .B(clk), .A(\g.we_clk [10464]));
Q_ASSIGN U22311 ( .B(clk), .A(\g.we_clk [10463]));
Q_ASSIGN U22312 ( .B(clk), .A(\g.we_clk [10462]));
Q_ASSIGN U22313 ( .B(clk), .A(\g.we_clk [10461]));
Q_ASSIGN U22314 ( .B(clk), .A(\g.we_clk [10460]));
Q_ASSIGN U22315 ( .B(clk), .A(\g.we_clk [10459]));
Q_ASSIGN U22316 ( .B(clk), .A(\g.we_clk [10458]));
Q_ASSIGN U22317 ( .B(clk), .A(\g.we_clk [10457]));
Q_ASSIGN U22318 ( .B(clk), .A(\g.we_clk [10456]));
Q_ASSIGN U22319 ( .B(clk), .A(\g.we_clk [10455]));
Q_ASSIGN U22320 ( .B(clk), .A(\g.we_clk [10454]));
Q_ASSIGN U22321 ( .B(clk), .A(\g.we_clk [10453]));
Q_ASSIGN U22322 ( .B(clk), .A(\g.we_clk [10452]));
Q_ASSIGN U22323 ( .B(clk), .A(\g.we_clk [10451]));
Q_ASSIGN U22324 ( .B(clk), .A(\g.we_clk [10450]));
Q_ASSIGN U22325 ( .B(clk), .A(\g.we_clk [10449]));
Q_ASSIGN U22326 ( .B(clk), .A(\g.we_clk [10448]));
Q_ASSIGN U22327 ( .B(clk), .A(\g.we_clk [10447]));
Q_ASSIGN U22328 ( .B(clk), .A(\g.we_clk [10446]));
Q_ASSIGN U22329 ( .B(clk), .A(\g.we_clk [10445]));
Q_ASSIGN U22330 ( .B(clk), .A(\g.we_clk [10444]));
Q_ASSIGN U22331 ( .B(clk), .A(\g.we_clk [10443]));
Q_ASSIGN U22332 ( .B(clk), .A(\g.we_clk [10442]));
Q_ASSIGN U22333 ( .B(clk), .A(\g.we_clk [10441]));
Q_ASSIGN U22334 ( .B(clk), .A(\g.we_clk [10440]));
Q_ASSIGN U22335 ( .B(clk), .A(\g.we_clk [10439]));
Q_ASSIGN U22336 ( .B(clk), .A(\g.we_clk [10438]));
Q_ASSIGN U22337 ( .B(clk), .A(\g.we_clk [10437]));
Q_ASSIGN U22338 ( .B(clk), .A(\g.we_clk [10436]));
Q_ASSIGN U22339 ( .B(clk), .A(\g.we_clk [10435]));
Q_ASSIGN U22340 ( .B(clk), .A(\g.we_clk [10434]));
Q_ASSIGN U22341 ( .B(clk), .A(\g.we_clk [10433]));
Q_ASSIGN U22342 ( .B(clk), .A(\g.we_clk [10432]));
Q_ASSIGN U22343 ( .B(clk), .A(\g.we_clk [10431]));
Q_ASSIGN U22344 ( .B(clk), .A(\g.we_clk [10430]));
Q_ASSIGN U22345 ( .B(clk), .A(\g.we_clk [10429]));
Q_ASSIGN U22346 ( .B(clk), .A(\g.we_clk [10428]));
Q_ASSIGN U22347 ( .B(clk), .A(\g.we_clk [10427]));
Q_ASSIGN U22348 ( .B(clk), .A(\g.we_clk [10426]));
Q_ASSIGN U22349 ( .B(clk), .A(\g.we_clk [10425]));
Q_ASSIGN U22350 ( .B(clk), .A(\g.we_clk [10424]));
Q_ASSIGN U22351 ( .B(clk), .A(\g.we_clk [10423]));
Q_ASSIGN U22352 ( .B(clk), .A(\g.we_clk [10422]));
Q_ASSIGN U22353 ( .B(clk), .A(\g.we_clk [10421]));
Q_ASSIGN U22354 ( .B(clk), .A(\g.we_clk [10420]));
Q_ASSIGN U22355 ( .B(clk), .A(\g.we_clk [10419]));
Q_ASSIGN U22356 ( .B(clk), .A(\g.we_clk [10418]));
Q_ASSIGN U22357 ( .B(clk), .A(\g.we_clk [10417]));
Q_ASSIGN U22358 ( .B(clk), .A(\g.we_clk [10416]));
Q_ASSIGN U22359 ( .B(clk), .A(\g.we_clk [10415]));
Q_ASSIGN U22360 ( .B(clk), .A(\g.we_clk [10414]));
Q_ASSIGN U22361 ( .B(clk), .A(\g.we_clk [10413]));
Q_ASSIGN U22362 ( .B(clk), .A(\g.we_clk [10412]));
Q_ASSIGN U22363 ( .B(clk), .A(\g.we_clk [10411]));
Q_ASSIGN U22364 ( .B(clk), .A(\g.we_clk [10410]));
Q_ASSIGN U22365 ( .B(clk), .A(\g.we_clk [10409]));
Q_ASSIGN U22366 ( .B(clk), .A(\g.we_clk [10408]));
Q_ASSIGN U22367 ( .B(clk), .A(\g.we_clk [10407]));
Q_ASSIGN U22368 ( .B(clk), .A(\g.we_clk [10406]));
Q_ASSIGN U22369 ( .B(clk), .A(\g.we_clk [10405]));
Q_ASSIGN U22370 ( .B(clk), .A(\g.we_clk [10404]));
Q_ASSIGN U22371 ( .B(clk), .A(\g.we_clk [10403]));
Q_ASSIGN U22372 ( .B(clk), .A(\g.we_clk [10402]));
Q_ASSIGN U22373 ( .B(clk), .A(\g.we_clk [10401]));
Q_ASSIGN U22374 ( .B(clk), .A(\g.we_clk [10400]));
Q_ASSIGN U22375 ( .B(clk), .A(\g.we_clk [10399]));
Q_ASSIGN U22376 ( .B(clk), .A(\g.we_clk [10398]));
Q_ASSIGN U22377 ( .B(clk), .A(\g.we_clk [10397]));
Q_ASSIGN U22378 ( .B(clk), .A(\g.we_clk [10396]));
Q_ASSIGN U22379 ( .B(clk), .A(\g.we_clk [10395]));
Q_ASSIGN U22380 ( .B(clk), .A(\g.we_clk [10394]));
Q_ASSIGN U22381 ( .B(clk), .A(\g.we_clk [10393]));
Q_ASSIGN U22382 ( .B(clk), .A(\g.we_clk [10392]));
Q_ASSIGN U22383 ( .B(clk), .A(\g.we_clk [10391]));
Q_ASSIGN U22384 ( .B(clk), .A(\g.we_clk [10390]));
Q_ASSIGN U22385 ( .B(clk), .A(\g.we_clk [10389]));
Q_ASSIGN U22386 ( .B(clk), .A(\g.we_clk [10388]));
Q_ASSIGN U22387 ( .B(clk), .A(\g.we_clk [10387]));
Q_ASSIGN U22388 ( .B(clk), .A(\g.we_clk [10386]));
Q_ASSIGN U22389 ( .B(clk), .A(\g.we_clk [10385]));
Q_ASSIGN U22390 ( .B(clk), .A(\g.we_clk [10384]));
Q_ASSIGN U22391 ( .B(clk), .A(\g.we_clk [10383]));
Q_ASSIGN U22392 ( .B(clk), .A(\g.we_clk [10382]));
Q_ASSIGN U22393 ( .B(clk), .A(\g.we_clk [10381]));
Q_ASSIGN U22394 ( .B(clk), .A(\g.we_clk [10380]));
Q_ASSIGN U22395 ( .B(clk), .A(\g.we_clk [10379]));
Q_ASSIGN U22396 ( .B(clk), .A(\g.we_clk [10378]));
Q_ASSIGN U22397 ( .B(clk), .A(\g.we_clk [10377]));
Q_ASSIGN U22398 ( .B(clk), .A(\g.we_clk [10376]));
Q_ASSIGN U22399 ( .B(clk), .A(\g.we_clk [10375]));
Q_ASSIGN U22400 ( .B(clk), .A(\g.we_clk [10374]));
Q_ASSIGN U22401 ( .B(clk), .A(\g.we_clk [10373]));
Q_ASSIGN U22402 ( .B(clk), .A(\g.we_clk [10372]));
Q_ASSIGN U22403 ( .B(clk), .A(\g.we_clk [10371]));
Q_ASSIGN U22404 ( .B(clk), .A(\g.we_clk [10370]));
Q_ASSIGN U22405 ( .B(clk), .A(\g.we_clk [10369]));
Q_ASSIGN U22406 ( .B(clk), .A(\g.we_clk [10368]));
Q_ASSIGN U22407 ( .B(clk), .A(\g.we_clk [10367]));
Q_ASSIGN U22408 ( .B(clk), .A(\g.we_clk [10366]));
Q_ASSIGN U22409 ( .B(clk), .A(\g.we_clk [10365]));
Q_ASSIGN U22410 ( .B(clk), .A(\g.we_clk [10364]));
Q_ASSIGN U22411 ( .B(clk), .A(\g.we_clk [10363]));
Q_ASSIGN U22412 ( .B(clk), .A(\g.we_clk [10362]));
Q_ASSIGN U22413 ( .B(clk), .A(\g.we_clk [10361]));
Q_ASSIGN U22414 ( .B(clk), .A(\g.we_clk [10360]));
Q_ASSIGN U22415 ( .B(clk), .A(\g.we_clk [10359]));
Q_ASSIGN U22416 ( .B(clk), .A(\g.we_clk [10358]));
Q_ASSIGN U22417 ( .B(clk), .A(\g.we_clk [10357]));
Q_ASSIGN U22418 ( .B(clk), .A(\g.we_clk [10356]));
Q_ASSIGN U22419 ( .B(clk), .A(\g.we_clk [10355]));
Q_ASSIGN U22420 ( .B(clk), .A(\g.we_clk [10354]));
Q_ASSIGN U22421 ( .B(clk), .A(\g.we_clk [10353]));
Q_ASSIGN U22422 ( .B(clk), .A(\g.we_clk [10352]));
Q_ASSIGN U22423 ( .B(clk), .A(\g.we_clk [10351]));
Q_ASSIGN U22424 ( .B(clk), .A(\g.we_clk [10350]));
Q_ASSIGN U22425 ( .B(clk), .A(\g.we_clk [10349]));
Q_ASSIGN U22426 ( .B(clk), .A(\g.we_clk [10348]));
Q_ASSIGN U22427 ( .B(clk), .A(\g.we_clk [10347]));
Q_ASSIGN U22428 ( .B(clk), .A(\g.we_clk [10346]));
Q_ASSIGN U22429 ( .B(clk), .A(\g.we_clk [10345]));
Q_ASSIGN U22430 ( .B(clk), .A(\g.we_clk [10344]));
Q_ASSIGN U22431 ( .B(clk), .A(\g.we_clk [10343]));
Q_ASSIGN U22432 ( .B(clk), .A(\g.we_clk [10342]));
Q_ASSIGN U22433 ( .B(clk), .A(\g.we_clk [10341]));
Q_ASSIGN U22434 ( .B(clk), .A(\g.we_clk [10340]));
Q_ASSIGN U22435 ( .B(clk), .A(\g.we_clk [10339]));
Q_ASSIGN U22436 ( .B(clk), .A(\g.we_clk [10338]));
Q_ASSIGN U22437 ( .B(clk), .A(\g.we_clk [10337]));
Q_ASSIGN U22438 ( .B(clk), .A(\g.we_clk [10336]));
Q_ASSIGN U22439 ( .B(clk), .A(\g.we_clk [10335]));
Q_ASSIGN U22440 ( .B(clk), .A(\g.we_clk [10334]));
Q_ASSIGN U22441 ( .B(clk), .A(\g.we_clk [10333]));
Q_ASSIGN U22442 ( .B(clk), .A(\g.we_clk [10332]));
Q_ASSIGN U22443 ( .B(clk), .A(\g.we_clk [10331]));
Q_ASSIGN U22444 ( .B(clk), .A(\g.we_clk [10330]));
Q_ASSIGN U22445 ( .B(clk), .A(\g.we_clk [10329]));
Q_ASSIGN U22446 ( .B(clk), .A(\g.we_clk [10328]));
Q_ASSIGN U22447 ( .B(clk), .A(\g.we_clk [10327]));
Q_ASSIGN U22448 ( .B(clk), .A(\g.we_clk [10326]));
Q_ASSIGN U22449 ( .B(clk), .A(\g.we_clk [10325]));
Q_ASSIGN U22450 ( .B(clk), .A(\g.we_clk [10324]));
Q_ASSIGN U22451 ( .B(clk), .A(\g.we_clk [10323]));
Q_ASSIGN U22452 ( .B(clk), .A(\g.we_clk [10322]));
Q_ASSIGN U22453 ( .B(clk), .A(\g.we_clk [10321]));
Q_ASSIGN U22454 ( .B(clk), .A(\g.we_clk [10320]));
Q_ASSIGN U22455 ( .B(clk), .A(\g.we_clk [10319]));
Q_ASSIGN U22456 ( .B(clk), .A(\g.we_clk [10318]));
Q_ASSIGN U22457 ( .B(clk), .A(\g.we_clk [10317]));
Q_ASSIGN U22458 ( .B(clk), .A(\g.we_clk [10316]));
Q_ASSIGN U22459 ( .B(clk), .A(\g.we_clk [10315]));
Q_ASSIGN U22460 ( .B(clk), .A(\g.we_clk [10314]));
Q_ASSIGN U22461 ( .B(clk), .A(\g.we_clk [10313]));
Q_ASSIGN U22462 ( .B(clk), .A(\g.we_clk [10312]));
Q_ASSIGN U22463 ( .B(clk), .A(\g.we_clk [10311]));
Q_ASSIGN U22464 ( .B(clk), .A(\g.we_clk [10310]));
Q_ASSIGN U22465 ( .B(clk), .A(\g.we_clk [10309]));
Q_ASSIGN U22466 ( .B(clk), .A(\g.we_clk [10308]));
Q_ASSIGN U22467 ( .B(clk), .A(\g.we_clk [10307]));
Q_ASSIGN U22468 ( .B(clk), .A(\g.we_clk [10306]));
Q_ASSIGN U22469 ( .B(clk), .A(\g.we_clk [10305]));
Q_ASSIGN U22470 ( .B(clk), .A(\g.we_clk [10304]));
Q_ASSIGN U22471 ( .B(clk), .A(\g.we_clk [10303]));
Q_ASSIGN U22472 ( .B(clk), .A(\g.we_clk [10302]));
Q_ASSIGN U22473 ( .B(clk), .A(\g.we_clk [10301]));
Q_ASSIGN U22474 ( .B(clk), .A(\g.we_clk [10300]));
Q_ASSIGN U22475 ( .B(clk), .A(\g.we_clk [10299]));
Q_ASSIGN U22476 ( .B(clk), .A(\g.we_clk [10298]));
Q_ASSIGN U22477 ( .B(clk), .A(\g.we_clk [10297]));
Q_ASSIGN U22478 ( .B(clk), .A(\g.we_clk [10296]));
Q_ASSIGN U22479 ( .B(clk), .A(\g.we_clk [10295]));
Q_ASSIGN U22480 ( .B(clk), .A(\g.we_clk [10294]));
Q_ASSIGN U22481 ( .B(clk), .A(\g.we_clk [10293]));
Q_ASSIGN U22482 ( .B(clk), .A(\g.we_clk [10292]));
Q_ASSIGN U22483 ( .B(clk), .A(\g.we_clk [10291]));
Q_ASSIGN U22484 ( .B(clk), .A(\g.we_clk [10290]));
Q_ASSIGN U22485 ( .B(clk), .A(\g.we_clk [10289]));
Q_ASSIGN U22486 ( .B(clk), .A(\g.we_clk [10288]));
Q_ASSIGN U22487 ( .B(clk), .A(\g.we_clk [10287]));
Q_ASSIGN U22488 ( .B(clk), .A(\g.we_clk [10286]));
Q_ASSIGN U22489 ( .B(clk), .A(\g.we_clk [10285]));
Q_ASSIGN U22490 ( .B(clk), .A(\g.we_clk [10284]));
Q_ASSIGN U22491 ( .B(clk), .A(\g.we_clk [10283]));
Q_ASSIGN U22492 ( .B(clk), .A(\g.we_clk [10282]));
Q_ASSIGN U22493 ( .B(clk), .A(\g.we_clk [10281]));
Q_ASSIGN U22494 ( .B(clk), .A(\g.we_clk [10280]));
Q_ASSIGN U22495 ( .B(clk), .A(\g.we_clk [10279]));
Q_ASSIGN U22496 ( .B(clk), .A(\g.we_clk [10278]));
Q_ASSIGN U22497 ( .B(clk), .A(\g.we_clk [10277]));
Q_ASSIGN U22498 ( .B(clk), .A(\g.we_clk [10276]));
Q_ASSIGN U22499 ( .B(clk), .A(\g.we_clk [10275]));
Q_ASSIGN U22500 ( .B(clk), .A(\g.we_clk [10274]));
Q_ASSIGN U22501 ( .B(clk), .A(\g.we_clk [10273]));
Q_ASSIGN U22502 ( .B(clk), .A(\g.we_clk [10272]));
Q_ASSIGN U22503 ( .B(clk), .A(\g.we_clk [10271]));
Q_ASSIGN U22504 ( .B(clk), .A(\g.we_clk [10270]));
Q_ASSIGN U22505 ( .B(clk), .A(\g.we_clk [10269]));
Q_ASSIGN U22506 ( .B(clk), .A(\g.we_clk [10268]));
Q_ASSIGN U22507 ( .B(clk), .A(\g.we_clk [10267]));
Q_ASSIGN U22508 ( .B(clk), .A(\g.we_clk [10266]));
Q_ASSIGN U22509 ( .B(clk), .A(\g.we_clk [10265]));
Q_ASSIGN U22510 ( .B(clk), .A(\g.we_clk [10264]));
Q_ASSIGN U22511 ( .B(clk), .A(\g.we_clk [10263]));
Q_ASSIGN U22512 ( .B(clk), .A(\g.we_clk [10262]));
Q_ASSIGN U22513 ( .B(clk), .A(\g.we_clk [10261]));
Q_ASSIGN U22514 ( .B(clk), .A(\g.we_clk [10260]));
Q_ASSIGN U22515 ( .B(clk), .A(\g.we_clk [10259]));
Q_ASSIGN U22516 ( .B(clk), .A(\g.we_clk [10258]));
Q_ASSIGN U22517 ( .B(clk), .A(\g.we_clk [10257]));
Q_ASSIGN U22518 ( .B(clk), .A(\g.we_clk [10256]));
Q_ASSIGN U22519 ( .B(clk), .A(\g.we_clk [10255]));
Q_ASSIGN U22520 ( .B(clk), .A(\g.we_clk [10254]));
Q_ASSIGN U22521 ( .B(clk), .A(\g.we_clk [10253]));
Q_ASSIGN U22522 ( .B(clk), .A(\g.we_clk [10252]));
Q_ASSIGN U22523 ( .B(clk), .A(\g.we_clk [10251]));
Q_ASSIGN U22524 ( .B(clk), .A(\g.we_clk [10250]));
Q_ASSIGN U22525 ( .B(clk), .A(\g.we_clk [10249]));
Q_ASSIGN U22526 ( .B(clk), .A(\g.we_clk [10248]));
Q_ASSIGN U22527 ( .B(clk), .A(\g.we_clk [10247]));
Q_ASSIGN U22528 ( .B(clk), .A(\g.we_clk [10246]));
Q_ASSIGN U22529 ( .B(clk), .A(\g.we_clk [10245]));
Q_ASSIGN U22530 ( .B(clk), .A(\g.we_clk [10244]));
Q_ASSIGN U22531 ( .B(clk), .A(\g.we_clk [10243]));
Q_ASSIGN U22532 ( .B(clk), .A(\g.we_clk [10242]));
Q_ASSIGN U22533 ( .B(clk), .A(\g.we_clk [10241]));
Q_ASSIGN U22534 ( .B(clk), .A(\g.we_clk [10240]));
Q_ASSIGN U22535 ( .B(clk), .A(\g.we_clk [10239]));
Q_ASSIGN U22536 ( .B(clk), .A(\g.we_clk [10238]));
Q_ASSIGN U22537 ( .B(clk), .A(\g.we_clk [10237]));
Q_ASSIGN U22538 ( .B(clk), .A(\g.we_clk [10236]));
Q_ASSIGN U22539 ( .B(clk), .A(\g.we_clk [10235]));
Q_ASSIGN U22540 ( .B(clk), .A(\g.we_clk [10234]));
Q_ASSIGN U22541 ( .B(clk), .A(\g.we_clk [10233]));
Q_ASSIGN U22542 ( .B(clk), .A(\g.we_clk [10232]));
Q_ASSIGN U22543 ( .B(clk), .A(\g.we_clk [10231]));
Q_ASSIGN U22544 ( .B(clk), .A(\g.we_clk [10230]));
Q_ASSIGN U22545 ( .B(clk), .A(\g.we_clk [10229]));
Q_ASSIGN U22546 ( .B(clk), .A(\g.we_clk [10228]));
Q_ASSIGN U22547 ( .B(clk), .A(\g.we_clk [10227]));
Q_ASSIGN U22548 ( .B(clk), .A(\g.we_clk [10226]));
Q_ASSIGN U22549 ( .B(clk), .A(\g.we_clk [10225]));
Q_ASSIGN U22550 ( .B(clk), .A(\g.we_clk [10224]));
Q_ASSIGN U22551 ( .B(clk), .A(\g.we_clk [10223]));
Q_ASSIGN U22552 ( .B(clk), .A(\g.we_clk [10222]));
Q_ASSIGN U22553 ( .B(clk), .A(\g.we_clk [10221]));
Q_ASSIGN U22554 ( .B(clk), .A(\g.we_clk [10220]));
Q_ASSIGN U22555 ( .B(clk), .A(\g.we_clk [10219]));
Q_ASSIGN U22556 ( .B(clk), .A(\g.we_clk [10218]));
Q_ASSIGN U22557 ( .B(clk), .A(\g.we_clk [10217]));
Q_ASSIGN U22558 ( .B(clk), .A(\g.we_clk [10216]));
Q_ASSIGN U22559 ( .B(clk), .A(\g.we_clk [10215]));
Q_ASSIGN U22560 ( .B(clk), .A(\g.we_clk [10214]));
Q_ASSIGN U22561 ( .B(clk), .A(\g.we_clk [10213]));
Q_ASSIGN U22562 ( .B(clk), .A(\g.we_clk [10212]));
Q_ASSIGN U22563 ( .B(clk), .A(\g.we_clk [10211]));
Q_ASSIGN U22564 ( .B(clk), .A(\g.we_clk [10210]));
Q_ASSIGN U22565 ( .B(clk), .A(\g.we_clk [10209]));
Q_ASSIGN U22566 ( .B(clk), .A(\g.we_clk [10208]));
Q_ASSIGN U22567 ( .B(clk), .A(\g.we_clk [10207]));
Q_ASSIGN U22568 ( .B(clk), .A(\g.we_clk [10206]));
Q_ASSIGN U22569 ( .B(clk), .A(\g.we_clk [10205]));
Q_ASSIGN U22570 ( .B(clk), .A(\g.we_clk [10204]));
Q_ASSIGN U22571 ( .B(clk), .A(\g.we_clk [10203]));
Q_ASSIGN U22572 ( .B(clk), .A(\g.we_clk [10202]));
Q_ASSIGN U22573 ( .B(clk), .A(\g.we_clk [10201]));
Q_ASSIGN U22574 ( .B(clk), .A(\g.we_clk [10200]));
Q_ASSIGN U22575 ( .B(clk), .A(\g.we_clk [10199]));
Q_ASSIGN U22576 ( .B(clk), .A(\g.we_clk [10198]));
Q_ASSIGN U22577 ( .B(clk), .A(\g.we_clk [10197]));
Q_ASSIGN U22578 ( .B(clk), .A(\g.we_clk [10196]));
Q_ASSIGN U22579 ( .B(clk), .A(\g.we_clk [10195]));
Q_ASSIGN U22580 ( .B(clk), .A(\g.we_clk [10194]));
Q_ASSIGN U22581 ( .B(clk), .A(\g.we_clk [10193]));
Q_ASSIGN U22582 ( .B(clk), .A(\g.we_clk [10192]));
Q_ASSIGN U22583 ( .B(clk), .A(\g.we_clk [10191]));
Q_ASSIGN U22584 ( .B(clk), .A(\g.we_clk [10190]));
Q_ASSIGN U22585 ( .B(clk), .A(\g.we_clk [10189]));
Q_ASSIGN U22586 ( .B(clk), .A(\g.we_clk [10188]));
Q_ASSIGN U22587 ( .B(clk), .A(\g.we_clk [10187]));
Q_ASSIGN U22588 ( .B(clk), .A(\g.we_clk [10186]));
Q_ASSIGN U22589 ( .B(clk), .A(\g.we_clk [10185]));
Q_ASSIGN U22590 ( .B(clk), .A(\g.we_clk [10184]));
Q_ASSIGN U22591 ( .B(clk), .A(\g.we_clk [10183]));
Q_ASSIGN U22592 ( .B(clk), .A(\g.we_clk [10182]));
Q_ASSIGN U22593 ( .B(clk), .A(\g.we_clk [10181]));
Q_ASSIGN U22594 ( .B(clk), .A(\g.we_clk [10180]));
Q_ASSIGN U22595 ( .B(clk), .A(\g.we_clk [10179]));
Q_ASSIGN U22596 ( .B(clk), .A(\g.we_clk [10178]));
Q_ASSIGN U22597 ( .B(clk), .A(\g.we_clk [10177]));
Q_ASSIGN U22598 ( .B(clk), .A(\g.we_clk [10176]));
Q_ASSIGN U22599 ( .B(clk), .A(\g.we_clk [10175]));
Q_ASSIGN U22600 ( .B(clk), .A(\g.we_clk [10174]));
Q_ASSIGN U22601 ( .B(clk), .A(\g.we_clk [10173]));
Q_ASSIGN U22602 ( .B(clk), .A(\g.we_clk [10172]));
Q_ASSIGN U22603 ( .B(clk), .A(\g.we_clk [10171]));
Q_ASSIGN U22604 ( .B(clk), .A(\g.we_clk [10170]));
Q_ASSIGN U22605 ( .B(clk), .A(\g.we_clk [10169]));
Q_ASSIGN U22606 ( .B(clk), .A(\g.we_clk [10168]));
Q_ASSIGN U22607 ( .B(clk), .A(\g.we_clk [10167]));
Q_ASSIGN U22608 ( .B(clk), .A(\g.we_clk [10166]));
Q_ASSIGN U22609 ( .B(clk), .A(\g.we_clk [10165]));
Q_ASSIGN U22610 ( .B(clk), .A(\g.we_clk [10164]));
Q_ASSIGN U22611 ( .B(clk), .A(\g.we_clk [10163]));
Q_ASSIGN U22612 ( .B(clk), .A(\g.we_clk [10162]));
Q_ASSIGN U22613 ( .B(clk), .A(\g.we_clk [10161]));
Q_ASSIGN U22614 ( .B(clk), .A(\g.we_clk [10160]));
Q_ASSIGN U22615 ( .B(clk), .A(\g.we_clk [10159]));
Q_ASSIGN U22616 ( .B(clk), .A(\g.we_clk [10158]));
Q_ASSIGN U22617 ( .B(clk), .A(\g.we_clk [10157]));
Q_ASSIGN U22618 ( .B(clk), .A(\g.we_clk [10156]));
Q_ASSIGN U22619 ( .B(clk), .A(\g.we_clk [10155]));
Q_ASSIGN U22620 ( .B(clk), .A(\g.we_clk [10154]));
Q_ASSIGN U22621 ( .B(clk), .A(\g.we_clk [10153]));
Q_ASSIGN U22622 ( .B(clk), .A(\g.we_clk [10152]));
Q_ASSIGN U22623 ( .B(clk), .A(\g.we_clk [10151]));
Q_ASSIGN U22624 ( .B(clk), .A(\g.we_clk [10150]));
Q_ASSIGN U22625 ( .B(clk), .A(\g.we_clk [10149]));
Q_ASSIGN U22626 ( .B(clk), .A(\g.we_clk [10148]));
Q_ASSIGN U22627 ( .B(clk), .A(\g.we_clk [10147]));
Q_ASSIGN U22628 ( .B(clk), .A(\g.we_clk [10146]));
Q_ASSIGN U22629 ( .B(clk), .A(\g.we_clk [10145]));
Q_ASSIGN U22630 ( .B(clk), .A(\g.we_clk [10144]));
Q_ASSIGN U22631 ( .B(clk), .A(\g.we_clk [10143]));
Q_ASSIGN U22632 ( .B(clk), .A(\g.we_clk [10142]));
Q_ASSIGN U22633 ( .B(clk), .A(\g.we_clk [10141]));
Q_ASSIGN U22634 ( .B(clk), .A(\g.we_clk [10140]));
Q_ASSIGN U22635 ( .B(clk), .A(\g.we_clk [10139]));
Q_ASSIGN U22636 ( .B(clk), .A(\g.we_clk [10138]));
Q_ASSIGN U22637 ( .B(clk), .A(\g.we_clk [10137]));
Q_ASSIGN U22638 ( .B(clk), .A(\g.we_clk [10136]));
Q_ASSIGN U22639 ( .B(clk), .A(\g.we_clk [10135]));
Q_ASSIGN U22640 ( .B(clk), .A(\g.we_clk [10134]));
Q_ASSIGN U22641 ( .B(clk), .A(\g.we_clk [10133]));
Q_ASSIGN U22642 ( .B(clk), .A(\g.we_clk [10132]));
Q_ASSIGN U22643 ( .B(clk), .A(\g.we_clk [10131]));
Q_ASSIGN U22644 ( .B(clk), .A(\g.we_clk [10130]));
Q_ASSIGN U22645 ( .B(clk), .A(\g.we_clk [10129]));
Q_ASSIGN U22646 ( .B(clk), .A(\g.we_clk [10128]));
Q_ASSIGN U22647 ( .B(clk), .A(\g.we_clk [10127]));
Q_ASSIGN U22648 ( .B(clk), .A(\g.we_clk [10126]));
Q_ASSIGN U22649 ( .B(clk), .A(\g.we_clk [10125]));
Q_ASSIGN U22650 ( .B(clk), .A(\g.we_clk [10124]));
Q_ASSIGN U22651 ( .B(clk), .A(\g.we_clk [10123]));
Q_ASSIGN U22652 ( .B(clk), .A(\g.we_clk [10122]));
Q_ASSIGN U22653 ( .B(clk), .A(\g.we_clk [10121]));
Q_ASSIGN U22654 ( .B(clk), .A(\g.we_clk [10120]));
Q_ASSIGN U22655 ( .B(clk), .A(\g.we_clk [10119]));
Q_ASSIGN U22656 ( .B(clk), .A(\g.we_clk [10118]));
Q_ASSIGN U22657 ( .B(clk), .A(\g.we_clk [10117]));
Q_ASSIGN U22658 ( .B(clk), .A(\g.we_clk [10116]));
Q_ASSIGN U22659 ( .B(clk), .A(\g.we_clk [10115]));
Q_ASSIGN U22660 ( .B(clk), .A(\g.we_clk [10114]));
Q_ASSIGN U22661 ( .B(clk), .A(\g.we_clk [10113]));
Q_ASSIGN U22662 ( .B(clk), .A(\g.we_clk [10112]));
Q_ASSIGN U22663 ( .B(clk), .A(\g.we_clk [10111]));
Q_ASSIGN U22664 ( .B(clk), .A(\g.we_clk [10110]));
Q_ASSIGN U22665 ( .B(clk), .A(\g.we_clk [10109]));
Q_ASSIGN U22666 ( .B(clk), .A(\g.we_clk [10108]));
Q_ASSIGN U22667 ( .B(clk), .A(\g.we_clk [10107]));
Q_ASSIGN U22668 ( .B(clk), .A(\g.we_clk [10106]));
Q_ASSIGN U22669 ( .B(clk), .A(\g.we_clk [10105]));
Q_ASSIGN U22670 ( .B(clk), .A(\g.we_clk [10104]));
Q_ASSIGN U22671 ( .B(clk), .A(\g.we_clk [10103]));
Q_ASSIGN U22672 ( .B(clk), .A(\g.we_clk [10102]));
Q_ASSIGN U22673 ( .B(clk), .A(\g.we_clk [10101]));
Q_ASSIGN U22674 ( .B(clk), .A(\g.we_clk [10100]));
Q_ASSIGN U22675 ( .B(clk), .A(\g.we_clk [10099]));
Q_ASSIGN U22676 ( .B(clk), .A(\g.we_clk [10098]));
Q_ASSIGN U22677 ( .B(clk), .A(\g.we_clk [10097]));
Q_ASSIGN U22678 ( .B(clk), .A(\g.we_clk [10096]));
Q_ASSIGN U22679 ( .B(clk), .A(\g.we_clk [10095]));
Q_ASSIGN U22680 ( .B(clk), .A(\g.we_clk [10094]));
Q_ASSIGN U22681 ( .B(clk), .A(\g.we_clk [10093]));
Q_ASSIGN U22682 ( .B(clk), .A(\g.we_clk [10092]));
Q_ASSIGN U22683 ( .B(clk), .A(\g.we_clk [10091]));
Q_ASSIGN U22684 ( .B(clk), .A(\g.we_clk [10090]));
Q_ASSIGN U22685 ( .B(clk), .A(\g.we_clk [10089]));
Q_ASSIGN U22686 ( .B(clk), .A(\g.we_clk [10088]));
Q_ASSIGN U22687 ( .B(clk), .A(\g.we_clk [10087]));
Q_ASSIGN U22688 ( .B(clk), .A(\g.we_clk [10086]));
Q_ASSIGN U22689 ( .B(clk), .A(\g.we_clk [10085]));
Q_ASSIGN U22690 ( .B(clk), .A(\g.we_clk [10084]));
Q_ASSIGN U22691 ( .B(clk), .A(\g.we_clk [10083]));
Q_ASSIGN U22692 ( .B(clk), .A(\g.we_clk [10082]));
Q_ASSIGN U22693 ( .B(clk), .A(\g.we_clk [10081]));
Q_ASSIGN U22694 ( .B(clk), .A(\g.we_clk [10080]));
Q_ASSIGN U22695 ( .B(clk), .A(\g.we_clk [10079]));
Q_ASSIGN U22696 ( .B(clk), .A(\g.we_clk [10078]));
Q_ASSIGN U22697 ( .B(clk), .A(\g.we_clk [10077]));
Q_ASSIGN U22698 ( .B(clk), .A(\g.we_clk [10076]));
Q_ASSIGN U22699 ( .B(clk), .A(\g.we_clk [10075]));
Q_ASSIGN U22700 ( .B(clk), .A(\g.we_clk [10074]));
Q_ASSIGN U22701 ( .B(clk), .A(\g.we_clk [10073]));
Q_ASSIGN U22702 ( .B(clk), .A(\g.we_clk [10072]));
Q_ASSIGN U22703 ( .B(clk), .A(\g.we_clk [10071]));
Q_ASSIGN U22704 ( .B(clk), .A(\g.we_clk [10070]));
Q_ASSIGN U22705 ( .B(clk), .A(\g.we_clk [10069]));
Q_ASSIGN U22706 ( .B(clk), .A(\g.we_clk [10068]));
Q_ASSIGN U22707 ( .B(clk), .A(\g.we_clk [10067]));
Q_ASSIGN U22708 ( .B(clk), .A(\g.we_clk [10066]));
Q_ASSIGN U22709 ( .B(clk), .A(\g.we_clk [10065]));
Q_ASSIGN U22710 ( .B(clk), .A(\g.we_clk [10064]));
Q_ASSIGN U22711 ( .B(clk), .A(\g.we_clk [10063]));
Q_ASSIGN U22712 ( .B(clk), .A(\g.we_clk [10062]));
Q_ASSIGN U22713 ( .B(clk), .A(\g.we_clk [10061]));
Q_ASSIGN U22714 ( .B(clk), .A(\g.we_clk [10060]));
Q_ASSIGN U22715 ( .B(clk), .A(\g.we_clk [10059]));
Q_ASSIGN U22716 ( .B(clk), .A(\g.we_clk [10058]));
Q_ASSIGN U22717 ( .B(clk), .A(\g.we_clk [10057]));
Q_ASSIGN U22718 ( .B(clk), .A(\g.we_clk [10056]));
Q_ASSIGN U22719 ( .B(clk), .A(\g.we_clk [10055]));
Q_ASSIGN U22720 ( .B(clk), .A(\g.we_clk [10054]));
Q_ASSIGN U22721 ( .B(clk), .A(\g.we_clk [10053]));
Q_ASSIGN U22722 ( .B(clk), .A(\g.we_clk [10052]));
Q_ASSIGN U22723 ( .B(clk), .A(\g.we_clk [10051]));
Q_ASSIGN U22724 ( .B(clk), .A(\g.we_clk [10050]));
Q_ASSIGN U22725 ( .B(clk), .A(\g.we_clk [10049]));
Q_ASSIGN U22726 ( .B(clk), .A(\g.we_clk [10048]));
Q_ASSIGN U22727 ( .B(clk), .A(\g.we_clk [10047]));
Q_ASSIGN U22728 ( .B(clk), .A(\g.we_clk [10046]));
Q_ASSIGN U22729 ( .B(clk), .A(\g.we_clk [10045]));
Q_ASSIGN U22730 ( .B(clk), .A(\g.we_clk [10044]));
Q_ASSIGN U22731 ( .B(clk), .A(\g.we_clk [10043]));
Q_ASSIGN U22732 ( .B(clk), .A(\g.we_clk [10042]));
Q_ASSIGN U22733 ( .B(clk), .A(\g.we_clk [10041]));
Q_ASSIGN U22734 ( .B(clk), .A(\g.we_clk [10040]));
Q_ASSIGN U22735 ( .B(clk), .A(\g.we_clk [10039]));
Q_ASSIGN U22736 ( .B(clk), .A(\g.we_clk [10038]));
Q_ASSIGN U22737 ( .B(clk), .A(\g.we_clk [10037]));
Q_ASSIGN U22738 ( .B(clk), .A(\g.we_clk [10036]));
Q_ASSIGN U22739 ( .B(clk), .A(\g.we_clk [10035]));
Q_ASSIGN U22740 ( .B(clk), .A(\g.we_clk [10034]));
Q_ASSIGN U22741 ( .B(clk), .A(\g.we_clk [10033]));
Q_ASSIGN U22742 ( .B(clk), .A(\g.we_clk [10032]));
Q_ASSIGN U22743 ( .B(clk), .A(\g.we_clk [10031]));
Q_ASSIGN U22744 ( .B(clk), .A(\g.we_clk [10030]));
Q_ASSIGN U22745 ( .B(clk), .A(\g.we_clk [10029]));
Q_ASSIGN U22746 ( .B(clk), .A(\g.we_clk [10028]));
Q_ASSIGN U22747 ( .B(clk), .A(\g.we_clk [10027]));
Q_ASSIGN U22748 ( .B(clk), .A(\g.we_clk [10026]));
Q_ASSIGN U22749 ( .B(clk), .A(\g.we_clk [10025]));
Q_ASSIGN U22750 ( .B(clk), .A(\g.we_clk [10024]));
Q_ASSIGN U22751 ( .B(clk), .A(\g.we_clk [10023]));
Q_ASSIGN U22752 ( .B(clk), .A(\g.we_clk [10022]));
Q_ASSIGN U22753 ( .B(clk), .A(\g.we_clk [10021]));
Q_ASSIGN U22754 ( .B(clk), .A(\g.we_clk [10020]));
Q_ASSIGN U22755 ( .B(clk), .A(\g.we_clk [10019]));
Q_ASSIGN U22756 ( .B(clk), .A(\g.we_clk [10018]));
Q_ASSIGN U22757 ( .B(clk), .A(\g.we_clk [10017]));
Q_ASSIGN U22758 ( .B(clk), .A(\g.we_clk [10016]));
Q_ASSIGN U22759 ( .B(clk), .A(\g.we_clk [10015]));
Q_ASSIGN U22760 ( .B(clk), .A(\g.we_clk [10014]));
Q_ASSIGN U22761 ( .B(clk), .A(\g.we_clk [10013]));
Q_ASSIGN U22762 ( .B(clk), .A(\g.we_clk [10012]));
Q_ASSIGN U22763 ( .B(clk), .A(\g.we_clk [10011]));
Q_ASSIGN U22764 ( .B(clk), .A(\g.we_clk [10010]));
Q_ASSIGN U22765 ( .B(clk), .A(\g.we_clk [10009]));
Q_ASSIGN U22766 ( .B(clk), .A(\g.we_clk [10008]));
Q_ASSIGN U22767 ( .B(clk), .A(\g.we_clk [10007]));
Q_ASSIGN U22768 ( .B(clk), .A(\g.we_clk [10006]));
Q_ASSIGN U22769 ( .B(clk), .A(\g.we_clk [10005]));
Q_ASSIGN U22770 ( .B(clk), .A(\g.we_clk [10004]));
Q_ASSIGN U22771 ( .B(clk), .A(\g.we_clk [10003]));
Q_ASSIGN U22772 ( .B(clk), .A(\g.we_clk [10002]));
Q_ASSIGN U22773 ( .B(clk), .A(\g.we_clk [10001]));
Q_ASSIGN U22774 ( .B(clk), .A(\g.we_clk [10000]));
Q_ASSIGN U22775 ( .B(clk), .A(\g.we_clk [9999]));
Q_ASSIGN U22776 ( .B(clk), .A(\g.we_clk [9998]));
Q_ASSIGN U22777 ( .B(clk), .A(\g.we_clk [9997]));
Q_ASSIGN U22778 ( .B(clk), .A(\g.we_clk [9996]));
Q_ASSIGN U22779 ( .B(clk), .A(\g.we_clk [9995]));
Q_ASSIGN U22780 ( .B(clk), .A(\g.we_clk [9994]));
Q_ASSIGN U22781 ( .B(clk), .A(\g.we_clk [9993]));
Q_ASSIGN U22782 ( .B(clk), .A(\g.we_clk [9992]));
Q_ASSIGN U22783 ( .B(clk), .A(\g.we_clk [9991]));
Q_ASSIGN U22784 ( .B(clk), .A(\g.we_clk [9990]));
Q_ASSIGN U22785 ( .B(clk), .A(\g.we_clk [9989]));
Q_ASSIGN U22786 ( .B(clk), .A(\g.we_clk [9988]));
Q_ASSIGN U22787 ( .B(clk), .A(\g.we_clk [9987]));
Q_ASSIGN U22788 ( .B(clk), .A(\g.we_clk [9986]));
Q_ASSIGN U22789 ( .B(clk), .A(\g.we_clk [9985]));
Q_ASSIGN U22790 ( .B(clk), .A(\g.we_clk [9984]));
Q_ASSIGN U22791 ( .B(clk), .A(\g.we_clk [9983]));
Q_ASSIGN U22792 ( .B(clk), .A(\g.we_clk [9982]));
Q_ASSIGN U22793 ( .B(clk), .A(\g.we_clk [9981]));
Q_ASSIGN U22794 ( .B(clk), .A(\g.we_clk [9980]));
Q_ASSIGN U22795 ( .B(clk), .A(\g.we_clk [9979]));
Q_ASSIGN U22796 ( .B(clk), .A(\g.we_clk [9978]));
Q_ASSIGN U22797 ( .B(clk), .A(\g.we_clk [9977]));
Q_ASSIGN U22798 ( .B(clk), .A(\g.we_clk [9976]));
Q_ASSIGN U22799 ( .B(clk), .A(\g.we_clk [9975]));
Q_ASSIGN U22800 ( .B(clk), .A(\g.we_clk [9974]));
Q_ASSIGN U22801 ( .B(clk), .A(\g.we_clk [9973]));
Q_ASSIGN U22802 ( .B(clk), .A(\g.we_clk [9972]));
Q_ASSIGN U22803 ( .B(clk), .A(\g.we_clk [9971]));
Q_ASSIGN U22804 ( .B(clk), .A(\g.we_clk [9970]));
Q_ASSIGN U22805 ( .B(clk), .A(\g.we_clk [9969]));
Q_ASSIGN U22806 ( .B(clk), .A(\g.we_clk [9968]));
Q_ASSIGN U22807 ( .B(clk), .A(\g.we_clk [9967]));
Q_ASSIGN U22808 ( .B(clk), .A(\g.we_clk [9966]));
Q_ASSIGN U22809 ( .B(clk), .A(\g.we_clk [9965]));
Q_ASSIGN U22810 ( .B(clk), .A(\g.we_clk [9964]));
Q_ASSIGN U22811 ( .B(clk), .A(\g.we_clk [9963]));
Q_ASSIGN U22812 ( .B(clk), .A(\g.we_clk [9962]));
Q_ASSIGN U22813 ( .B(clk), .A(\g.we_clk [9961]));
Q_ASSIGN U22814 ( .B(clk), .A(\g.we_clk [9960]));
Q_ASSIGN U22815 ( .B(clk), .A(\g.we_clk [9959]));
Q_ASSIGN U22816 ( .B(clk), .A(\g.we_clk [9958]));
Q_ASSIGN U22817 ( .B(clk), .A(\g.we_clk [9957]));
Q_ASSIGN U22818 ( .B(clk), .A(\g.we_clk [9956]));
Q_ASSIGN U22819 ( .B(clk), .A(\g.we_clk [9955]));
Q_ASSIGN U22820 ( .B(clk), .A(\g.we_clk [9954]));
Q_ASSIGN U22821 ( .B(clk), .A(\g.we_clk [9953]));
Q_ASSIGN U22822 ( .B(clk), .A(\g.we_clk [9952]));
Q_ASSIGN U22823 ( .B(clk), .A(\g.we_clk [9951]));
Q_ASSIGN U22824 ( .B(clk), .A(\g.we_clk [9950]));
Q_ASSIGN U22825 ( .B(clk), .A(\g.we_clk [9949]));
Q_ASSIGN U22826 ( .B(clk), .A(\g.we_clk [9948]));
Q_ASSIGN U22827 ( .B(clk), .A(\g.we_clk [9947]));
Q_ASSIGN U22828 ( .B(clk), .A(\g.we_clk [9946]));
Q_ASSIGN U22829 ( .B(clk), .A(\g.we_clk [9945]));
Q_ASSIGN U22830 ( .B(clk), .A(\g.we_clk [9944]));
Q_ASSIGN U22831 ( .B(clk), .A(\g.we_clk [9943]));
Q_ASSIGN U22832 ( .B(clk), .A(\g.we_clk [9942]));
Q_ASSIGN U22833 ( .B(clk), .A(\g.we_clk [9941]));
Q_ASSIGN U22834 ( .B(clk), .A(\g.we_clk [9940]));
Q_ASSIGN U22835 ( .B(clk), .A(\g.we_clk [9939]));
Q_ASSIGN U22836 ( .B(clk), .A(\g.we_clk [9938]));
Q_ASSIGN U22837 ( .B(clk), .A(\g.we_clk [9937]));
Q_ASSIGN U22838 ( .B(clk), .A(\g.we_clk [9936]));
Q_ASSIGN U22839 ( .B(clk), .A(\g.we_clk [9935]));
Q_ASSIGN U22840 ( .B(clk), .A(\g.we_clk [9934]));
Q_ASSIGN U22841 ( .B(clk), .A(\g.we_clk [9933]));
Q_ASSIGN U22842 ( .B(clk), .A(\g.we_clk [9932]));
Q_ASSIGN U22843 ( .B(clk), .A(\g.we_clk [9931]));
Q_ASSIGN U22844 ( .B(clk), .A(\g.we_clk [9930]));
Q_ASSIGN U22845 ( .B(clk), .A(\g.we_clk [9929]));
Q_ASSIGN U22846 ( .B(clk), .A(\g.we_clk [9928]));
Q_ASSIGN U22847 ( .B(clk), .A(\g.we_clk [9927]));
Q_ASSIGN U22848 ( .B(clk), .A(\g.we_clk [9926]));
Q_ASSIGN U22849 ( .B(clk), .A(\g.we_clk [9925]));
Q_ASSIGN U22850 ( .B(clk), .A(\g.we_clk [9924]));
Q_ASSIGN U22851 ( .B(clk), .A(\g.we_clk [9923]));
Q_ASSIGN U22852 ( .B(clk), .A(\g.we_clk [9922]));
Q_ASSIGN U22853 ( .B(clk), .A(\g.we_clk [9921]));
Q_ASSIGN U22854 ( .B(clk), .A(\g.we_clk [9920]));
Q_ASSIGN U22855 ( .B(clk), .A(\g.we_clk [9919]));
Q_ASSIGN U22856 ( .B(clk), .A(\g.we_clk [9918]));
Q_ASSIGN U22857 ( .B(clk), .A(\g.we_clk [9917]));
Q_ASSIGN U22858 ( .B(clk), .A(\g.we_clk [9916]));
Q_ASSIGN U22859 ( .B(clk), .A(\g.we_clk [9915]));
Q_ASSIGN U22860 ( .B(clk), .A(\g.we_clk [9914]));
Q_ASSIGN U22861 ( .B(clk), .A(\g.we_clk [9913]));
Q_ASSIGN U22862 ( .B(clk), .A(\g.we_clk [9912]));
Q_ASSIGN U22863 ( .B(clk), .A(\g.we_clk [9911]));
Q_ASSIGN U22864 ( .B(clk), .A(\g.we_clk [9910]));
Q_ASSIGN U22865 ( .B(clk), .A(\g.we_clk [9909]));
Q_ASSIGN U22866 ( .B(clk), .A(\g.we_clk [9908]));
Q_ASSIGN U22867 ( .B(clk), .A(\g.we_clk [9907]));
Q_ASSIGN U22868 ( .B(clk), .A(\g.we_clk [9906]));
Q_ASSIGN U22869 ( .B(clk), .A(\g.we_clk [9905]));
Q_ASSIGN U22870 ( .B(clk), .A(\g.we_clk [9904]));
Q_ASSIGN U22871 ( .B(clk), .A(\g.we_clk [9903]));
Q_ASSIGN U22872 ( .B(clk), .A(\g.we_clk [9902]));
Q_ASSIGN U22873 ( .B(clk), .A(\g.we_clk [9901]));
Q_ASSIGN U22874 ( .B(clk), .A(\g.we_clk [9900]));
Q_ASSIGN U22875 ( .B(clk), .A(\g.we_clk [9899]));
Q_ASSIGN U22876 ( .B(clk), .A(\g.we_clk [9898]));
Q_ASSIGN U22877 ( .B(clk), .A(\g.we_clk [9897]));
Q_ASSIGN U22878 ( .B(clk), .A(\g.we_clk [9896]));
Q_ASSIGN U22879 ( .B(clk), .A(\g.we_clk [9895]));
Q_ASSIGN U22880 ( .B(clk), .A(\g.we_clk [9894]));
Q_ASSIGN U22881 ( .B(clk), .A(\g.we_clk [9893]));
Q_ASSIGN U22882 ( .B(clk), .A(\g.we_clk [9892]));
Q_ASSIGN U22883 ( .B(clk), .A(\g.we_clk [9891]));
Q_ASSIGN U22884 ( .B(clk), .A(\g.we_clk [9890]));
Q_ASSIGN U22885 ( .B(clk), .A(\g.we_clk [9889]));
Q_ASSIGN U22886 ( .B(clk), .A(\g.we_clk [9888]));
Q_ASSIGN U22887 ( .B(clk), .A(\g.we_clk [9887]));
Q_ASSIGN U22888 ( .B(clk), .A(\g.we_clk [9886]));
Q_ASSIGN U22889 ( .B(clk), .A(\g.we_clk [9885]));
Q_ASSIGN U22890 ( .B(clk), .A(\g.we_clk [9884]));
Q_ASSIGN U22891 ( .B(clk), .A(\g.we_clk [9883]));
Q_ASSIGN U22892 ( .B(clk), .A(\g.we_clk [9882]));
Q_ASSIGN U22893 ( .B(clk), .A(\g.we_clk [9881]));
Q_ASSIGN U22894 ( .B(clk), .A(\g.we_clk [9880]));
Q_ASSIGN U22895 ( .B(clk), .A(\g.we_clk [9879]));
Q_ASSIGN U22896 ( .B(clk), .A(\g.we_clk [9878]));
Q_ASSIGN U22897 ( .B(clk), .A(\g.we_clk [9877]));
Q_ASSIGN U22898 ( .B(clk), .A(\g.we_clk [9876]));
Q_ASSIGN U22899 ( .B(clk), .A(\g.we_clk [9875]));
Q_ASSIGN U22900 ( .B(clk), .A(\g.we_clk [9874]));
Q_ASSIGN U22901 ( .B(clk), .A(\g.we_clk [9873]));
Q_ASSIGN U22902 ( .B(clk), .A(\g.we_clk [9872]));
Q_ASSIGN U22903 ( .B(clk), .A(\g.we_clk [9871]));
Q_ASSIGN U22904 ( .B(clk), .A(\g.we_clk [9870]));
Q_ASSIGN U22905 ( .B(clk), .A(\g.we_clk [9869]));
Q_ASSIGN U22906 ( .B(clk), .A(\g.we_clk [9868]));
Q_ASSIGN U22907 ( .B(clk), .A(\g.we_clk [9867]));
Q_ASSIGN U22908 ( .B(clk), .A(\g.we_clk [9866]));
Q_ASSIGN U22909 ( .B(clk), .A(\g.we_clk [9865]));
Q_ASSIGN U22910 ( .B(clk), .A(\g.we_clk [9864]));
Q_ASSIGN U22911 ( .B(clk), .A(\g.we_clk [9863]));
Q_ASSIGN U22912 ( .B(clk), .A(\g.we_clk [9862]));
Q_ASSIGN U22913 ( .B(clk), .A(\g.we_clk [9861]));
Q_ASSIGN U22914 ( .B(clk), .A(\g.we_clk [9860]));
Q_ASSIGN U22915 ( .B(clk), .A(\g.we_clk [9859]));
Q_ASSIGN U22916 ( .B(clk), .A(\g.we_clk [9858]));
Q_ASSIGN U22917 ( .B(clk), .A(\g.we_clk [9857]));
Q_ASSIGN U22918 ( .B(clk), .A(\g.we_clk [9856]));
Q_ASSIGN U22919 ( .B(clk), .A(\g.we_clk [9855]));
Q_ASSIGN U22920 ( .B(clk), .A(\g.we_clk [9854]));
Q_ASSIGN U22921 ( .B(clk), .A(\g.we_clk [9853]));
Q_ASSIGN U22922 ( .B(clk), .A(\g.we_clk [9852]));
Q_ASSIGN U22923 ( .B(clk), .A(\g.we_clk [9851]));
Q_ASSIGN U22924 ( .B(clk), .A(\g.we_clk [9850]));
Q_ASSIGN U22925 ( .B(clk), .A(\g.we_clk [9849]));
Q_ASSIGN U22926 ( .B(clk), .A(\g.we_clk [9848]));
Q_ASSIGN U22927 ( .B(clk), .A(\g.we_clk [9847]));
Q_ASSIGN U22928 ( .B(clk), .A(\g.we_clk [9846]));
Q_ASSIGN U22929 ( .B(clk), .A(\g.we_clk [9845]));
Q_ASSIGN U22930 ( .B(clk), .A(\g.we_clk [9844]));
Q_ASSIGN U22931 ( .B(clk), .A(\g.we_clk [9843]));
Q_ASSIGN U22932 ( .B(clk), .A(\g.we_clk [9842]));
Q_ASSIGN U22933 ( .B(clk), .A(\g.we_clk [9841]));
Q_ASSIGN U22934 ( .B(clk), .A(\g.we_clk [9840]));
Q_ASSIGN U22935 ( .B(clk), .A(\g.we_clk [9839]));
Q_ASSIGN U22936 ( .B(clk), .A(\g.we_clk [9838]));
Q_ASSIGN U22937 ( .B(clk), .A(\g.we_clk [9837]));
Q_ASSIGN U22938 ( .B(clk), .A(\g.we_clk [9836]));
Q_ASSIGN U22939 ( .B(clk), .A(\g.we_clk [9835]));
Q_ASSIGN U22940 ( .B(clk), .A(\g.we_clk [9834]));
Q_ASSIGN U22941 ( .B(clk), .A(\g.we_clk [9833]));
Q_ASSIGN U22942 ( .B(clk), .A(\g.we_clk [9832]));
Q_ASSIGN U22943 ( .B(clk), .A(\g.we_clk [9831]));
Q_ASSIGN U22944 ( .B(clk), .A(\g.we_clk [9830]));
Q_ASSIGN U22945 ( .B(clk), .A(\g.we_clk [9829]));
Q_ASSIGN U22946 ( .B(clk), .A(\g.we_clk [9828]));
Q_ASSIGN U22947 ( .B(clk), .A(\g.we_clk [9827]));
Q_ASSIGN U22948 ( .B(clk), .A(\g.we_clk [9826]));
Q_ASSIGN U22949 ( .B(clk), .A(\g.we_clk [9825]));
Q_ASSIGN U22950 ( .B(clk), .A(\g.we_clk [9824]));
Q_ASSIGN U22951 ( .B(clk), .A(\g.we_clk [9823]));
Q_ASSIGN U22952 ( .B(clk), .A(\g.we_clk [9822]));
Q_ASSIGN U22953 ( .B(clk), .A(\g.we_clk [9821]));
Q_ASSIGN U22954 ( .B(clk), .A(\g.we_clk [9820]));
Q_ASSIGN U22955 ( .B(clk), .A(\g.we_clk [9819]));
Q_ASSIGN U22956 ( .B(clk), .A(\g.we_clk [9818]));
Q_ASSIGN U22957 ( .B(clk), .A(\g.we_clk [9817]));
Q_ASSIGN U22958 ( .B(clk), .A(\g.we_clk [9816]));
Q_ASSIGN U22959 ( .B(clk), .A(\g.we_clk [9815]));
Q_ASSIGN U22960 ( .B(clk), .A(\g.we_clk [9814]));
Q_ASSIGN U22961 ( .B(clk), .A(\g.we_clk [9813]));
Q_ASSIGN U22962 ( .B(clk), .A(\g.we_clk [9812]));
Q_ASSIGN U22963 ( .B(clk), .A(\g.we_clk [9811]));
Q_ASSIGN U22964 ( .B(clk), .A(\g.we_clk [9810]));
Q_ASSIGN U22965 ( .B(clk), .A(\g.we_clk [9809]));
Q_ASSIGN U22966 ( .B(clk), .A(\g.we_clk [9808]));
Q_ASSIGN U22967 ( .B(clk), .A(\g.we_clk [9807]));
Q_ASSIGN U22968 ( .B(clk), .A(\g.we_clk [9806]));
Q_ASSIGN U22969 ( .B(clk), .A(\g.we_clk [9805]));
Q_ASSIGN U22970 ( .B(clk), .A(\g.we_clk [9804]));
Q_ASSIGN U22971 ( .B(clk), .A(\g.we_clk [9803]));
Q_ASSIGN U22972 ( .B(clk), .A(\g.we_clk [9802]));
Q_ASSIGN U22973 ( .B(clk), .A(\g.we_clk [9801]));
Q_ASSIGN U22974 ( .B(clk), .A(\g.we_clk [9800]));
Q_ASSIGN U22975 ( .B(clk), .A(\g.we_clk [9799]));
Q_ASSIGN U22976 ( .B(clk), .A(\g.we_clk [9798]));
Q_ASSIGN U22977 ( .B(clk), .A(\g.we_clk [9797]));
Q_ASSIGN U22978 ( .B(clk), .A(\g.we_clk [9796]));
Q_ASSIGN U22979 ( .B(clk), .A(\g.we_clk [9795]));
Q_ASSIGN U22980 ( .B(clk), .A(\g.we_clk [9794]));
Q_ASSIGN U22981 ( .B(clk), .A(\g.we_clk [9793]));
Q_ASSIGN U22982 ( .B(clk), .A(\g.we_clk [9792]));
Q_ASSIGN U22983 ( .B(clk), .A(\g.we_clk [9791]));
Q_ASSIGN U22984 ( .B(clk), .A(\g.we_clk [9790]));
Q_ASSIGN U22985 ( .B(clk), .A(\g.we_clk [9789]));
Q_ASSIGN U22986 ( .B(clk), .A(\g.we_clk [9788]));
Q_ASSIGN U22987 ( .B(clk), .A(\g.we_clk [9787]));
Q_ASSIGN U22988 ( .B(clk), .A(\g.we_clk [9786]));
Q_ASSIGN U22989 ( .B(clk), .A(\g.we_clk [9785]));
Q_ASSIGN U22990 ( .B(clk), .A(\g.we_clk [9784]));
Q_ASSIGN U22991 ( .B(clk), .A(\g.we_clk [9783]));
Q_ASSIGN U22992 ( .B(clk), .A(\g.we_clk [9782]));
Q_ASSIGN U22993 ( .B(clk), .A(\g.we_clk [9781]));
Q_ASSIGN U22994 ( .B(clk), .A(\g.we_clk [9780]));
Q_ASSIGN U22995 ( .B(clk), .A(\g.we_clk [9779]));
Q_ASSIGN U22996 ( .B(clk), .A(\g.we_clk [9778]));
Q_ASSIGN U22997 ( .B(clk), .A(\g.we_clk [9777]));
Q_ASSIGN U22998 ( .B(clk), .A(\g.we_clk [9776]));
Q_ASSIGN U22999 ( .B(clk), .A(\g.we_clk [9775]));
Q_ASSIGN U23000 ( .B(clk), .A(\g.we_clk [9774]));
Q_ASSIGN U23001 ( .B(clk), .A(\g.we_clk [9773]));
Q_ASSIGN U23002 ( .B(clk), .A(\g.we_clk [9772]));
Q_ASSIGN U23003 ( .B(clk), .A(\g.we_clk [9771]));
Q_ASSIGN U23004 ( .B(clk), .A(\g.we_clk [9770]));
Q_ASSIGN U23005 ( .B(clk), .A(\g.we_clk [9769]));
Q_ASSIGN U23006 ( .B(clk), .A(\g.we_clk [9768]));
Q_ASSIGN U23007 ( .B(clk), .A(\g.we_clk [9767]));
Q_ASSIGN U23008 ( .B(clk), .A(\g.we_clk [9766]));
Q_ASSIGN U23009 ( .B(clk), .A(\g.we_clk [9765]));
Q_ASSIGN U23010 ( .B(clk), .A(\g.we_clk [9764]));
Q_ASSIGN U23011 ( .B(clk), .A(\g.we_clk [9763]));
Q_ASSIGN U23012 ( .B(clk), .A(\g.we_clk [9762]));
Q_ASSIGN U23013 ( .B(clk), .A(\g.we_clk [9761]));
Q_ASSIGN U23014 ( .B(clk), .A(\g.we_clk [9760]));
Q_ASSIGN U23015 ( .B(clk), .A(\g.we_clk [9759]));
Q_ASSIGN U23016 ( .B(clk), .A(\g.we_clk [9758]));
Q_ASSIGN U23017 ( .B(clk), .A(\g.we_clk [9757]));
Q_ASSIGN U23018 ( .B(clk), .A(\g.we_clk [9756]));
Q_ASSIGN U23019 ( .B(clk), .A(\g.we_clk [9755]));
Q_ASSIGN U23020 ( .B(clk), .A(\g.we_clk [9754]));
Q_ASSIGN U23021 ( .B(clk), .A(\g.we_clk [9753]));
Q_ASSIGN U23022 ( .B(clk), .A(\g.we_clk [9752]));
Q_ASSIGN U23023 ( .B(clk), .A(\g.we_clk [9751]));
Q_ASSIGN U23024 ( .B(clk), .A(\g.we_clk [9750]));
Q_ASSIGN U23025 ( .B(clk), .A(\g.we_clk [9749]));
Q_ASSIGN U23026 ( .B(clk), .A(\g.we_clk [9748]));
Q_ASSIGN U23027 ( .B(clk), .A(\g.we_clk [9747]));
Q_ASSIGN U23028 ( .B(clk), .A(\g.we_clk [9746]));
Q_ASSIGN U23029 ( .B(clk), .A(\g.we_clk [9745]));
Q_ASSIGN U23030 ( .B(clk), .A(\g.we_clk [9744]));
Q_ASSIGN U23031 ( .B(clk), .A(\g.we_clk [9743]));
Q_ASSIGN U23032 ( .B(clk), .A(\g.we_clk [9742]));
Q_ASSIGN U23033 ( .B(clk), .A(\g.we_clk [9741]));
Q_ASSIGN U23034 ( .B(clk), .A(\g.we_clk [9740]));
Q_ASSIGN U23035 ( .B(clk), .A(\g.we_clk [9739]));
Q_ASSIGN U23036 ( .B(clk), .A(\g.we_clk [9738]));
Q_ASSIGN U23037 ( .B(clk), .A(\g.we_clk [9737]));
Q_ASSIGN U23038 ( .B(clk), .A(\g.we_clk [9736]));
Q_ASSIGN U23039 ( .B(clk), .A(\g.we_clk [9735]));
Q_ASSIGN U23040 ( .B(clk), .A(\g.we_clk [9734]));
Q_ASSIGN U23041 ( .B(clk), .A(\g.we_clk [9733]));
Q_ASSIGN U23042 ( .B(clk), .A(\g.we_clk [9732]));
Q_ASSIGN U23043 ( .B(clk), .A(\g.we_clk [9731]));
Q_ASSIGN U23044 ( .B(clk), .A(\g.we_clk [9730]));
Q_ASSIGN U23045 ( .B(clk), .A(\g.we_clk [9729]));
Q_ASSIGN U23046 ( .B(clk), .A(\g.we_clk [9728]));
Q_ASSIGN U23047 ( .B(clk), .A(\g.we_clk [9727]));
Q_ASSIGN U23048 ( .B(clk), .A(\g.we_clk [9726]));
Q_ASSIGN U23049 ( .B(clk), .A(\g.we_clk [9725]));
Q_ASSIGN U23050 ( .B(clk), .A(\g.we_clk [9724]));
Q_ASSIGN U23051 ( .B(clk), .A(\g.we_clk [9723]));
Q_ASSIGN U23052 ( .B(clk), .A(\g.we_clk [9722]));
Q_ASSIGN U23053 ( .B(clk), .A(\g.we_clk [9721]));
Q_ASSIGN U23054 ( .B(clk), .A(\g.we_clk [9720]));
Q_ASSIGN U23055 ( .B(clk), .A(\g.we_clk [9719]));
Q_ASSIGN U23056 ( .B(clk), .A(\g.we_clk [9718]));
Q_ASSIGN U23057 ( .B(clk), .A(\g.we_clk [9717]));
Q_ASSIGN U23058 ( .B(clk), .A(\g.we_clk [9716]));
Q_ASSIGN U23059 ( .B(clk), .A(\g.we_clk [9715]));
Q_ASSIGN U23060 ( .B(clk), .A(\g.we_clk [9714]));
Q_ASSIGN U23061 ( .B(clk), .A(\g.we_clk [9713]));
Q_ASSIGN U23062 ( .B(clk), .A(\g.we_clk [9712]));
Q_ASSIGN U23063 ( .B(clk), .A(\g.we_clk [9711]));
Q_ASSIGN U23064 ( .B(clk), .A(\g.we_clk [9710]));
Q_ASSIGN U23065 ( .B(clk), .A(\g.we_clk [9709]));
Q_ASSIGN U23066 ( .B(clk), .A(\g.we_clk [9708]));
Q_ASSIGN U23067 ( .B(clk), .A(\g.we_clk [9707]));
Q_ASSIGN U23068 ( .B(clk), .A(\g.we_clk [9706]));
Q_ASSIGN U23069 ( .B(clk), .A(\g.we_clk [9705]));
Q_ASSIGN U23070 ( .B(clk), .A(\g.we_clk [9704]));
Q_ASSIGN U23071 ( .B(clk), .A(\g.we_clk [9703]));
Q_ASSIGN U23072 ( .B(clk), .A(\g.we_clk [9702]));
Q_ASSIGN U23073 ( .B(clk), .A(\g.we_clk [9701]));
Q_ASSIGN U23074 ( .B(clk), .A(\g.we_clk [9700]));
Q_ASSIGN U23075 ( .B(clk), .A(\g.we_clk [9699]));
Q_ASSIGN U23076 ( .B(clk), .A(\g.we_clk [9698]));
Q_ASSIGN U23077 ( .B(clk), .A(\g.we_clk [9697]));
Q_ASSIGN U23078 ( .B(clk), .A(\g.we_clk [9696]));
Q_ASSIGN U23079 ( .B(clk), .A(\g.we_clk [9695]));
Q_ASSIGN U23080 ( .B(clk), .A(\g.we_clk [9694]));
Q_ASSIGN U23081 ( .B(clk), .A(\g.we_clk [9693]));
Q_ASSIGN U23082 ( .B(clk), .A(\g.we_clk [9692]));
Q_ASSIGN U23083 ( .B(clk), .A(\g.we_clk [9691]));
Q_ASSIGN U23084 ( .B(clk), .A(\g.we_clk [9690]));
Q_ASSIGN U23085 ( .B(clk), .A(\g.we_clk [9689]));
Q_ASSIGN U23086 ( .B(clk), .A(\g.we_clk [9688]));
Q_ASSIGN U23087 ( .B(clk), .A(\g.we_clk [9687]));
Q_ASSIGN U23088 ( .B(clk), .A(\g.we_clk [9686]));
Q_ASSIGN U23089 ( .B(clk), .A(\g.we_clk [9685]));
Q_ASSIGN U23090 ( .B(clk), .A(\g.we_clk [9684]));
Q_ASSIGN U23091 ( .B(clk), .A(\g.we_clk [9683]));
Q_ASSIGN U23092 ( .B(clk), .A(\g.we_clk [9682]));
Q_ASSIGN U23093 ( .B(clk), .A(\g.we_clk [9681]));
Q_ASSIGN U23094 ( .B(clk), .A(\g.we_clk [9680]));
Q_ASSIGN U23095 ( .B(clk), .A(\g.we_clk [9679]));
Q_ASSIGN U23096 ( .B(clk), .A(\g.we_clk [9678]));
Q_ASSIGN U23097 ( .B(clk), .A(\g.we_clk [9677]));
Q_ASSIGN U23098 ( .B(clk), .A(\g.we_clk [9676]));
Q_ASSIGN U23099 ( .B(clk), .A(\g.we_clk [9675]));
Q_ASSIGN U23100 ( .B(clk), .A(\g.we_clk [9674]));
Q_ASSIGN U23101 ( .B(clk), .A(\g.we_clk [9673]));
Q_ASSIGN U23102 ( .B(clk), .A(\g.we_clk [9672]));
Q_ASSIGN U23103 ( .B(clk), .A(\g.we_clk [9671]));
Q_ASSIGN U23104 ( .B(clk), .A(\g.we_clk [9670]));
Q_ASSIGN U23105 ( .B(clk), .A(\g.we_clk [9669]));
Q_ASSIGN U23106 ( .B(clk), .A(\g.we_clk [9668]));
Q_ASSIGN U23107 ( .B(clk), .A(\g.we_clk [9667]));
Q_ASSIGN U23108 ( .B(clk), .A(\g.we_clk [9666]));
Q_ASSIGN U23109 ( .B(clk), .A(\g.we_clk [9665]));
Q_ASSIGN U23110 ( .B(clk), .A(\g.we_clk [9664]));
Q_ASSIGN U23111 ( .B(clk), .A(\g.we_clk [9663]));
Q_ASSIGN U23112 ( .B(clk), .A(\g.we_clk [9662]));
Q_ASSIGN U23113 ( .B(clk), .A(\g.we_clk [9661]));
Q_ASSIGN U23114 ( .B(clk), .A(\g.we_clk [9660]));
Q_ASSIGN U23115 ( .B(clk), .A(\g.we_clk [9659]));
Q_ASSIGN U23116 ( .B(clk), .A(\g.we_clk [9658]));
Q_ASSIGN U23117 ( .B(clk), .A(\g.we_clk [9657]));
Q_ASSIGN U23118 ( .B(clk), .A(\g.we_clk [9656]));
Q_ASSIGN U23119 ( .B(clk), .A(\g.we_clk [9655]));
Q_ASSIGN U23120 ( .B(clk), .A(\g.we_clk [9654]));
Q_ASSIGN U23121 ( .B(clk), .A(\g.we_clk [9653]));
Q_ASSIGN U23122 ( .B(clk), .A(\g.we_clk [9652]));
Q_ASSIGN U23123 ( .B(clk), .A(\g.we_clk [9651]));
Q_ASSIGN U23124 ( .B(clk), .A(\g.we_clk [9650]));
Q_ASSIGN U23125 ( .B(clk), .A(\g.we_clk [9649]));
Q_ASSIGN U23126 ( .B(clk), .A(\g.we_clk [9648]));
Q_ASSIGN U23127 ( .B(clk), .A(\g.we_clk [9647]));
Q_ASSIGN U23128 ( .B(clk), .A(\g.we_clk [9646]));
Q_ASSIGN U23129 ( .B(clk), .A(\g.we_clk [9645]));
Q_ASSIGN U23130 ( .B(clk), .A(\g.we_clk [9644]));
Q_ASSIGN U23131 ( .B(clk), .A(\g.we_clk [9643]));
Q_ASSIGN U23132 ( .B(clk), .A(\g.we_clk [9642]));
Q_ASSIGN U23133 ( .B(clk), .A(\g.we_clk [9641]));
Q_ASSIGN U23134 ( .B(clk), .A(\g.we_clk [9640]));
Q_ASSIGN U23135 ( .B(clk), .A(\g.we_clk [9639]));
Q_ASSIGN U23136 ( .B(clk), .A(\g.we_clk [9638]));
Q_ASSIGN U23137 ( .B(clk), .A(\g.we_clk [9637]));
Q_ASSIGN U23138 ( .B(clk), .A(\g.we_clk [9636]));
Q_ASSIGN U23139 ( .B(clk), .A(\g.we_clk [9635]));
Q_ASSIGN U23140 ( .B(clk), .A(\g.we_clk [9634]));
Q_ASSIGN U23141 ( .B(clk), .A(\g.we_clk [9633]));
Q_ASSIGN U23142 ( .B(clk), .A(\g.we_clk [9632]));
Q_ASSIGN U23143 ( .B(clk), .A(\g.we_clk [9631]));
Q_ASSIGN U23144 ( .B(clk), .A(\g.we_clk [9630]));
Q_ASSIGN U23145 ( .B(clk), .A(\g.we_clk [9629]));
Q_ASSIGN U23146 ( .B(clk), .A(\g.we_clk [9628]));
Q_ASSIGN U23147 ( .B(clk), .A(\g.we_clk [9627]));
Q_ASSIGN U23148 ( .B(clk), .A(\g.we_clk [9626]));
Q_ASSIGN U23149 ( .B(clk), .A(\g.we_clk [9625]));
Q_ASSIGN U23150 ( .B(clk), .A(\g.we_clk [9624]));
Q_ASSIGN U23151 ( .B(clk), .A(\g.we_clk [9623]));
Q_ASSIGN U23152 ( .B(clk), .A(\g.we_clk [9622]));
Q_ASSIGN U23153 ( .B(clk), .A(\g.we_clk [9621]));
Q_ASSIGN U23154 ( .B(clk), .A(\g.we_clk [9620]));
Q_ASSIGN U23155 ( .B(clk), .A(\g.we_clk [9619]));
Q_ASSIGN U23156 ( .B(clk), .A(\g.we_clk [9618]));
Q_ASSIGN U23157 ( .B(clk), .A(\g.we_clk [9617]));
Q_ASSIGN U23158 ( .B(clk), .A(\g.we_clk [9616]));
Q_ASSIGN U23159 ( .B(clk), .A(\g.we_clk [9615]));
Q_ASSIGN U23160 ( .B(clk), .A(\g.we_clk [9614]));
Q_ASSIGN U23161 ( .B(clk), .A(\g.we_clk [9613]));
Q_ASSIGN U23162 ( .B(clk), .A(\g.we_clk [9612]));
Q_ASSIGN U23163 ( .B(clk), .A(\g.we_clk [9611]));
Q_ASSIGN U23164 ( .B(clk), .A(\g.we_clk [9610]));
Q_ASSIGN U23165 ( .B(clk), .A(\g.we_clk [9609]));
Q_ASSIGN U23166 ( .B(clk), .A(\g.we_clk [9608]));
Q_ASSIGN U23167 ( .B(clk), .A(\g.we_clk [9607]));
Q_ASSIGN U23168 ( .B(clk), .A(\g.we_clk [9606]));
Q_ASSIGN U23169 ( .B(clk), .A(\g.we_clk [9605]));
Q_ASSIGN U23170 ( .B(clk), .A(\g.we_clk [9604]));
Q_ASSIGN U23171 ( .B(clk), .A(\g.we_clk [9603]));
Q_ASSIGN U23172 ( .B(clk), .A(\g.we_clk [9602]));
Q_ASSIGN U23173 ( .B(clk), .A(\g.we_clk [9601]));
Q_ASSIGN U23174 ( .B(clk), .A(\g.we_clk [9600]));
Q_ASSIGN U23175 ( .B(clk), .A(\g.we_clk [9599]));
Q_ASSIGN U23176 ( .B(clk), .A(\g.we_clk [9598]));
Q_ASSIGN U23177 ( .B(clk), .A(\g.we_clk [9597]));
Q_ASSIGN U23178 ( .B(clk), .A(\g.we_clk [9596]));
Q_ASSIGN U23179 ( .B(clk), .A(\g.we_clk [9595]));
Q_ASSIGN U23180 ( .B(clk), .A(\g.we_clk [9594]));
Q_ASSIGN U23181 ( .B(clk), .A(\g.we_clk [9593]));
Q_ASSIGN U23182 ( .B(clk), .A(\g.we_clk [9592]));
Q_ASSIGN U23183 ( .B(clk), .A(\g.we_clk [9591]));
Q_ASSIGN U23184 ( .B(clk), .A(\g.we_clk [9590]));
Q_ASSIGN U23185 ( .B(clk), .A(\g.we_clk [9589]));
Q_ASSIGN U23186 ( .B(clk), .A(\g.we_clk [9588]));
Q_ASSIGN U23187 ( .B(clk), .A(\g.we_clk [9587]));
Q_ASSIGN U23188 ( .B(clk), .A(\g.we_clk [9586]));
Q_ASSIGN U23189 ( .B(clk), .A(\g.we_clk [9585]));
Q_ASSIGN U23190 ( .B(clk), .A(\g.we_clk [9584]));
Q_ASSIGN U23191 ( .B(clk), .A(\g.we_clk [9583]));
Q_ASSIGN U23192 ( .B(clk), .A(\g.we_clk [9582]));
Q_ASSIGN U23193 ( .B(clk), .A(\g.we_clk [9581]));
Q_ASSIGN U23194 ( .B(clk), .A(\g.we_clk [9580]));
Q_ASSIGN U23195 ( .B(clk), .A(\g.we_clk [9579]));
Q_ASSIGN U23196 ( .B(clk), .A(\g.we_clk [9578]));
Q_ASSIGN U23197 ( .B(clk), .A(\g.we_clk [9577]));
Q_ASSIGN U23198 ( .B(clk), .A(\g.we_clk [9576]));
Q_ASSIGN U23199 ( .B(clk), .A(\g.we_clk [9575]));
Q_ASSIGN U23200 ( .B(clk), .A(\g.we_clk [9574]));
Q_ASSIGN U23201 ( .B(clk), .A(\g.we_clk [9573]));
Q_ASSIGN U23202 ( .B(clk), .A(\g.we_clk [9572]));
Q_ASSIGN U23203 ( .B(clk), .A(\g.we_clk [9571]));
Q_ASSIGN U23204 ( .B(clk), .A(\g.we_clk [9570]));
Q_ASSIGN U23205 ( .B(clk), .A(\g.we_clk [9569]));
Q_ASSIGN U23206 ( .B(clk), .A(\g.we_clk [9568]));
Q_ASSIGN U23207 ( .B(clk), .A(\g.we_clk [9567]));
Q_ASSIGN U23208 ( .B(clk), .A(\g.we_clk [9566]));
Q_ASSIGN U23209 ( .B(clk), .A(\g.we_clk [9565]));
Q_ASSIGN U23210 ( .B(clk), .A(\g.we_clk [9564]));
Q_ASSIGN U23211 ( .B(clk), .A(\g.we_clk [9563]));
Q_ASSIGN U23212 ( .B(clk), .A(\g.we_clk [9562]));
Q_ASSIGN U23213 ( .B(clk), .A(\g.we_clk [9561]));
Q_ASSIGN U23214 ( .B(clk), .A(\g.we_clk [9560]));
Q_ASSIGN U23215 ( .B(clk), .A(\g.we_clk [9559]));
Q_ASSIGN U23216 ( .B(clk), .A(\g.we_clk [9558]));
Q_ASSIGN U23217 ( .B(clk), .A(\g.we_clk [9557]));
Q_ASSIGN U23218 ( .B(clk), .A(\g.we_clk [9556]));
Q_ASSIGN U23219 ( .B(clk), .A(\g.we_clk [9555]));
Q_ASSIGN U23220 ( .B(clk), .A(\g.we_clk [9554]));
Q_ASSIGN U23221 ( .B(clk), .A(\g.we_clk [9553]));
Q_ASSIGN U23222 ( .B(clk), .A(\g.we_clk [9552]));
Q_ASSIGN U23223 ( .B(clk), .A(\g.we_clk [9551]));
Q_ASSIGN U23224 ( .B(clk), .A(\g.we_clk [9550]));
Q_ASSIGN U23225 ( .B(clk), .A(\g.we_clk [9549]));
Q_ASSIGN U23226 ( .B(clk), .A(\g.we_clk [9548]));
Q_ASSIGN U23227 ( .B(clk), .A(\g.we_clk [9547]));
Q_ASSIGN U23228 ( .B(clk), .A(\g.we_clk [9546]));
Q_ASSIGN U23229 ( .B(clk), .A(\g.we_clk [9545]));
Q_ASSIGN U23230 ( .B(clk), .A(\g.we_clk [9544]));
Q_ASSIGN U23231 ( .B(clk), .A(\g.we_clk [9543]));
Q_ASSIGN U23232 ( .B(clk), .A(\g.we_clk [9542]));
Q_ASSIGN U23233 ( .B(clk), .A(\g.we_clk [9541]));
Q_ASSIGN U23234 ( .B(clk), .A(\g.we_clk [9540]));
Q_ASSIGN U23235 ( .B(clk), .A(\g.we_clk [9539]));
Q_ASSIGN U23236 ( .B(clk), .A(\g.we_clk [9538]));
Q_ASSIGN U23237 ( .B(clk), .A(\g.we_clk [9537]));
Q_ASSIGN U23238 ( .B(clk), .A(\g.we_clk [9536]));
Q_ASSIGN U23239 ( .B(clk), .A(\g.we_clk [9535]));
Q_ASSIGN U23240 ( .B(clk), .A(\g.we_clk [9534]));
Q_ASSIGN U23241 ( .B(clk), .A(\g.we_clk [9533]));
Q_ASSIGN U23242 ( .B(clk), .A(\g.we_clk [9532]));
Q_ASSIGN U23243 ( .B(clk), .A(\g.we_clk [9531]));
Q_ASSIGN U23244 ( .B(clk), .A(\g.we_clk [9530]));
Q_ASSIGN U23245 ( .B(clk), .A(\g.we_clk [9529]));
Q_ASSIGN U23246 ( .B(clk), .A(\g.we_clk [9528]));
Q_ASSIGN U23247 ( .B(clk), .A(\g.we_clk [9527]));
Q_ASSIGN U23248 ( .B(clk), .A(\g.we_clk [9526]));
Q_ASSIGN U23249 ( .B(clk), .A(\g.we_clk [9525]));
Q_ASSIGN U23250 ( .B(clk), .A(\g.we_clk [9524]));
Q_ASSIGN U23251 ( .B(clk), .A(\g.we_clk [9523]));
Q_ASSIGN U23252 ( .B(clk), .A(\g.we_clk [9522]));
Q_ASSIGN U23253 ( .B(clk), .A(\g.we_clk [9521]));
Q_ASSIGN U23254 ( .B(clk), .A(\g.we_clk [9520]));
Q_ASSIGN U23255 ( .B(clk), .A(\g.we_clk [9519]));
Q_ASSIGN U23256 ( .B(clk), .A(\g.we_clk [9518]));
Q_ASSIGN U23257 ( .B(clk), .A(\g.we_clk [9517]));
Q_ASSIGN U23258 ( .B(clk), .A(\g.we_clk [9516]));
Q_ASSIGN U23259 ( .B(clk), .A(\g.we_clk [9515]));
Q_ASSIGN U23260 ( .B(clk), .A(\g.we_clk [9514]));
Q_ASSIGN U23261 ( .B(clk), .A(\g.we_clk [9513]));
Q_ASSIGN U23262 ( .B(clk), .A(\g.we_clk [9512]));
Q_ASSIGN U23263 ( .B(clk), .A(\g.we_clk [9511]));
Q_ASSIGN U23264 ( .B(clk), .A(\g.we_clk [9510]));
Q_ASSIGN U23265 ( .B(clk), .A(\g.we_clk [9509]));
Q_ASSIGN U23266 ( .B(clk), .A(\g.we_clk [9508]));
Q_ASSIGN U23267 ( .B(clk), .A(\g.we_clk [9507]));
Q_ASSIGN U23268 ( .B(clk), .A(\g.we_clk [9506]));
Q_ASSIGN U23269 ( .B(clk), .A(\g.we_clk [9505]));
Q_ASSIGN U23270 ( .B(clk), .A(\g.we_clk [9504]));
Q_ASSIGN U23271 ( .B(clk), .A(\g.we_clk [9503]));
Q_ASSIGN U23272 ( .B(clk), .A(\g.we_clk [9502]));
Q_ASSIGN U23273 ( .B(clk), .A(\g.we_clk [9501]));
Q_ASSIGN U23274 ( .B(clk), .A(\g.we_clk [9500]));
Q_ASSIGN U23275 ( .B(clk), .A(\g.we_clk [9499]));
Q_ASSIGN U23276 ( .B(clk), .A(\g.we_clk [9498]));
Q_ASSIGN U23277 ( .B(clk), .A(\g.we_clk [9497]));
Q_ASSIGN U23278 ( .B(clk), .A(\g.we_clk [9496]));
Q_ASSIGN U23279 ( .B(clk), .A(\g.we_clk [9495]));
Q_ASSIGN U23280 ( .B(clk), .A(\g.we_clk [9494]));
Q_ASSIGN U23281 ( .B(clk), .A(\g.we_clk [9493]));
Q_ASSIGN U23282 ( .B(clk), .A(\g.we_clk [9492]));
Q_ASSIGN U23283 ( .B(clk), .A(\g.we_clk [9491]));
Q_ASSIGN U23284 ( .B(clk), .A(\g.we_clk [9490]));
Q_ASSIGN U23285 ( .B(clk), .A(\g.we_clk [9489]));
Q_ASSIGN U23286 ( .B(clk), .A(\g.we_clk [9488]));
Q_ASSIGN U23287 ( .B(clk), .A(\g.we_clk [9487]));
Q_ASSIGN U23288 ( .B(clk), .A(\g.we_clk [9486]));
Q_ASSIGN U23289 ( .B(clk), .A(\g.we_clk [9485]));
Q_ASSIGN U23290 ( .B(clk), .A(\g.we_clk [9484]));
Q_ASSIGN U23291 ( .B(clk), .A(\g.we_clk [9483]));
Q_ASSIGN U23292 ( .B(clk), .A(\g.we_clk [9482]));
Q_ASSIGN U23293 ( .B(clk), .A(\g.we_clk [9481]));
Q_ASSIGN U23294 ( .B(clk), .A(\g.we_clk [9480]));
Q_ASSIGN U23295 ( .B(clk), .A(\g.we_clk [9479]));
Q_ASSIGN U23296 ( .B(clk), .A(\g.we_clk [9478]));
Q_ASSIGN U23297 ( .B(clk), .A(\g.we_clk [9477]));
Q_ASSIGN U23298 ( .B(clk), .A(\g.we_clk [9476]));
Q_ASSIGN U23299 ( .B(clk), .A(\g.we_clk [9475]));
Q_ASSIGN U23300 ( .B(clk), .A(\g.we_clk [9474]));
Q_ASSIGN U23301 ( .B(clk), .A(\g.we_clk [9473]));
Q_ASSIGN U23302 ( .B(clk), .A(\g.we_clk [9472]));
Q_ASSIGN U23303 ( .B(clk), .A(\g.we_clk [9471]));
Q_ASSIGN U23304 ( .B(clk), .A(\g.we_clk [9470]));
Q_ASSIGN U23305 ( .B(clk), .A(\g.we_clk [9469]));
Q_ASSIGN U23306 ( .B(clk), .A(\g.we_clk [9468]));
Q_ASSIGN U23307 ( .B(clk), .A(\g.we_clk [9467]));
Q_ASSIGN U23308 ( .B(clk), .A(\g.we_clk [9466]));
Q_ASSIGN U23309 ( .B(clk), .A(\g.we_clk [9465]));
Q_ASSIGN U23310 ( .B(clk), .A(\g.we_clk [9464]));
Q_ASSIGN U23311 ( .B(clk), .A(\g.we_clk [9463]));
Q_ASSIGN U23312 ( .B(clk), .A(\g.we_clk [9462]));
Q_ASSIGN U23313 ( .B(clk), .A(\g.we_clk [9461]));
Q_ASSIGN U23314 ( .B(clk), .A(\g.we_clk [9460]));
Q_ASSIGN U23315 ( .B(clk), .A(\g.we_clk [9459]));
Q_ASSIGN U23316 ( .B(clk), .A(\g.we_clk [9458]));
Q_ASSIGN U23317 ( .B(clk), .A(\g.we_clk [9457]));
Q_ASSIGN U23318 ( .B(clk), .A(\g.we_clk [9456]));
Q_ASSIGN U23319 ( .B(clk), .A(\g.we_clk [9455]));
Q_ASSIGN U23320 ( .B(clk), .A(\g.we_clk [9454]));
Q_ASSIGN U23321 ( .B(clk), .A(\g.we_clk [9453]));
Q_ASSIGN U23322 ( .B(clk), .A(\g.we_clk [9452]));
Q_ASSIGN U23323 ( .B(clk), .A(\g.we_clk [9451]));
Q_ASSIGN U23324 ( .B(clk), .A(\g.we_clk [9450]));
Q_ASSIGN U23325 ( .B(clk), .A(\g.we_clk [9449]));
Q_ASSIGN U23326 ( .B(clk), .A(\g.we_clk [9448]));
Q_ASSIGN U23327 ( .B(clk), .A(\g.we_clk [9447]));
Q_ASSIGN U23328 ( .B(clk), .A(\g.we_clk [9446]));
Q_ASSIGN U23329 ( .B(clk), .A(\g.we_clk [9445]));
Q_ASSIGN U23330 ( .B(clk), .A(\g.we_clk [9444]));
Q_ASSIGN U23331 ( .B(clk), .A(\g.we_clk [9443]));
Q_ASSIGN U23332 ( .B(clk), .A(\g.we_clk [9442]));
Q_ASSIGN U23333 ( .B(clk), .A(\g.we_clk [9441]));
Q_ASSIGN U23334 ( .B(clk), .A(\g.we_clk [9440]));
Q_ASSIGN U23335 ( .B(clk), .A(\g.we_clk [9439]));
Q_ASSIGN U23336 ( .B(clk), .A(\g.we_clk [9438]));
Q_ASSIGN U23337 ( .B(clk), .A(\g.we_clk [9437]));
Q_ASSIGN U23338 ( .B(clk), .A(\g.we_clk [9436]));
Q_ASSIGN U23339 ( .B(clk), .A(\g.we_clk [9435]));
Q_ASSIGN U23340 ( .B(clk), .A(\g.we_clk [9434]));
Q_ASSIGN U23341 ( .B(clk), .A(\g.we_clk [9433]));
Q_ASSIGN U23342 ( .B(clk), .A(\g.we_clk [9432]));
Q_ASSIGN U23343 ( .B(clk), .A(\g.we_clk [9431]));
Q_ASSIGN U23344 ( .B(clk), .A(\g.we_clk [9430]));
Q_ASSIGN U23345 ( .B(clk), .A(\g.we_clk [9429]));
Q_ASSIGN U23346 ( .B(clk), .A(\g.we_clk [9428]));
Q_ASSIGN U23347 ( .B(clk), .A(\g.we_clk [9427]));
Q_ASSIGN U23348 ( .B(clk), .A(\g.we_clk [9426]));
Q_ASSIGN U23349 ( .B(clk), .A(\g.we_clk [9425]));
Q_ASSIGN U23350 ( .B(clk), .A(\g.we_clk [9424]));
Q_ASSIGN U23351 ( .B(clk), .A(\g.we_clk [9423]));
Q_ASSIGN U23352 ( .B(clk), .A(\g.we_clk [9422]));
Q_ASSIGN U23353 ( .B(clk), .A(\g.we_clk [9421]));
Q_ASSIGN U23354 ( .B(clk), .A(\g.we_clk [9420]));
Q_ASSIGN U23355 ( .B(clk), .A(\g.we_clk [9419]));
Q_ASSIGN U23356 ( .B(clk), .A(\g.we_clk [9418]));
Q_ASSIGN U23357 ( .B(clk), .A(\g.we_clk [9417]));
Q_ASSIGN U23358 ( .B(clk), .A(\g.we_clk [9416]));
Q_ASSIGN U23359 ( .B(clk), .A(\g.we_clk [9415]));
Q_ASSIGN U23360 ( .B(clk), .A(\g.we_clk [9414]));
Q_ASSIGN U23361 ( .B(clk), .A(\g.we_clk [9413]));
Q_ASSIGN U23362 ( .B(clk), .A(\g.we_clk [9412]));
Q_ASSIGN U23363 ( .B(clk), .A(\g.we_clk [9411]));
Q_ASSIGN U23364 ( .B(clk), .A(\g.we_clk [9410]));
Q_ASSIGN U23365 ( .B(clk), .A(\g.we_clk [9409]));
Q_ASSIGN U23366 ( .B(clk), .A(\g.we_clk [9408]));
Q_ASSIGN U23367 ( .B(clk), .A(\g.we_clk [9407]));
Q_ASSIGN U23368 ( .B(clk), .A(\g.we_clk [9406]));
Q_ASSIGN U23369 ( .B(clk), .A(\g.we_clk [9405]));
Q_ASSIGN U23370 ( .B(clk), .A(\g.we_clk [9404]));
Q_ASSIGN U23371 ( .B(clk), .A(\g.we_clk [9403]));
Q_ASSIGN U23372 ( .B(clk), .A(\g.we_clk [9402]));
Q_ASSIGN U23373 ( .B(clk), .A(\g.we_clk [9401]));
Q_ASSIGN U23374 ( .B(clk), .A(\g.we_clk [9400]));
Q_ASSIGN U23375 ( .B(clk), .A(\g.we_clk [9399]));
Q_ASSIGN U23376 ( .B(clk), .A(\g.we_clk [9398]));
Q_ASSIGN U23377 ( .B(clk), .A(\g.we_clk [9397]));
Q_ASSIGN U23378 ( .B(clk), .A(\g.we_clk [9396]));
Q_ASSIGN U23379 ( .B(clk), .A(\g.we_clk [9395]));
Q_ASSIGN U23380 ( .B(clk), .A(\g.we_clk [9394]));
Q_ASSIGN U23381 ( .B(clk), .A(\g.we_clk [9393]));
Q_ASSIGN U23382 ( .B(clk), .A(\g.we_clk [9392]));
Q_ASSIGN U23383 ( .B(clk), .A(\g.we_clk [9391]));
Q_ASSIGN U23384 ( .B(clk), .A(\g.we_clk [9390]));
Q_ASSIGN U23385 ( .B(clk), .A(\g.we_clk [9389]));
Q_ASSIGN U23386 ( .B(clk), .A(\g.we_clk [9388]));
Q_ASSIGN U23387 ( .B(clk), .A(\g.we_clk [9387]));
Q_ASSIGN U23388 ( .B(clk), .A(\g.we_clk [9386]));
Q_ASSIGN U23389 ( .B(clk), .A(\g.we_clk [9385]));
Q_ASSIGN U23390 ( .B(clk), .A(\g.we_clk [9384]));
Q_ASSIGN U23391 ( .B(clk), .A(\g.we_clk [9383]));
Q_ASSIGN U23392 ( .B(clk), .A(\g.we_clk [9382]));
Q_ASSIGN U23393 ( .B(clk), .A(\g.we_clk [9381]));
Q_ASSIGN U23394 ( .B(clk), .A(\g.we_clk [9380]));
Q_ASSIGN U23395 ( .B(clk), .A(\g.we_clk [9379]));
Q_ASSIGN U23396 ( .B(clk), .A(\g.we_clk [9378]));
Q_ASSIGN U23397 ( .B(clk), .A(\g.we_clk [9377]));
Q_ASSIGN U23398 ( .B(clk), .A(\g.we_clk [9376]));
Q_ASSIGN U23399 ( .B(clk), .A(\g.we_clk [9375]));
Q_ASSIGN U23400 ( .B(clk), .A(\g.we_clk [9374]));
Q_ASSIGN U23401 ( .B(clk), .A(\g.we_clk [9373]));
Q_ASSIGN U23402 ( .B(clk), .A(\g.we_clk [9372]));
Q_ASSIGN U23403 ( .B(clk), .A(\g.we_clk [9371]));
Q_ASSIGN U23404 ( .B(clk), .A(\g.we_clk [9370]));
Q_ASSIGN U23405 ( .B(clk), .A(\g.we_clk [9369]));
Q_ASSIGN U23406 ( .B(clk), .A(\g.we_clk [9368]));
Q_ASSIGN U23407 ( .B(clk), .A(\g.we_clk [9367]));
Q_ASSIGN U23408 ( .B(clk), .A(\g.we_clk [9366]));
Q_ASSIGN U23409 ( .B(clk), .A(\g.we_clk [9365]));
Q_ASSIGN U23410 ( .B(clk), .A(\g.we_clk [9364]));
Q_ASSIGN U23411 ( .B(clk), .A(\g.we_clk [9363]));
Q_ASSIGN U23412 ( .B(clk), .A(\g.we_clk [9362]));
Q_ASSIGN U23413 ( .B(clk), .A(\g.we_clk [9361]));
Q_ASSIGN U23414 ( .B(clk), .A(\g.we_clk [9360]));
Q_ASSIGN U23415 ( .B(clk), .A(\g.we_clk [9359]));
Q_ASSIGN U23416 ( .B(clk), .A(\g.we_clk [9358]));
Q_ASSIGN U23417 ( .B(clk), .A(\g.we_clk [9357]));
Q_ASSIGN U23418 ( .B(clk), .A(\g.we_clk [9356]));
Q_ASSIGN U23419 ( .B(clk), .A(\g.we_clk [9355]));
Q_ASSIGN U23420 ( .B(clk), .A(\g.we_clk [9354]));
Q_ASSIGN U23421 ( .B(clk), .A(\g.we_clk [9353]));
Q_ASSIGN U23422 ( .B(clk), .A(\g.we_clk [9352]));
Q_ASSIGN U23423 ( .B(clk), .A(\g.we_clk [9351]));
Q_ASSIGN U23424 ( .B(clk), .A(\g.we_clk [9350]));
Q_ASSIGN U23425 ( .B(clk), .A(\g.we_clk [9349]));
Q_ASSIGN U23426 ( .B(clk), .A(\g.we_clk [9348]));
Q_ASSIGN U23427 ( .B(clk), .A(\g.we_clk [9347]));
Q_ASSIGN U23428 ( .B(clk), .A(\g.we_clk [9346]));
Q_ASSIGN U23429 ( .B(clk), .A(\g.we_clk [9345]));
Q_ASSIGN U23430 ( .B(clk), .A(\g.we_clk [9344]));
Q_ASSIGN U23431 ( .B(clk), .A(\g.we_clk [9343]));
Q_ASSIGN U23432 ( .B(clk), .A(\g.we_clk [9342]));
Q_ASSIGN U23433 ( .B(clk), .A(\g.we_clk [9341]));
Q_ASSIGN U23434 ( .B(clk), .A(\g.we_clk [9340]));
Q_ASSIGN U23435 ( .B(clk), .A(\g.we_clk [9339]));
Q_ASSIGN U23436 ( .B(clk), .A(\g.we_clk [9338]));
Q_ASSIGN U23437 ( .B(clk), .A(\g.we_clk [9337]));
Q_ASSIGN U23438 ( .B(clk), .A(\g.we_clk [9336]));
Q_ASSIGN U23439 ( .B(clk), .A(\g.we_clk [9335]));
Q_ASSIGN U23440 ( .B(clk), .A(\g.we_clk [9334]));
Q_ASSIGN U23441 ( .B(clk), .A(\g.we_clk [9333]));
Q_ASSIGN U23442 ( .B(clk), .A(\g.we_clk [9332]));
Q_ASSIGN U23443 ( .B(clk), .A(\g.we_clk [9331]));
Q_ASSIGN U23444 ( .B(clk), .A(\g.we_clk [9330]));
Q_ASSIGN U23445 ( .B(clk), .A(\g.we_clk [9329]));
Q_ASSIGN U23446 ( .B(clk), .A(\g.we_clk [9328]));
Q_ASSIGN U23447 ( .B(clk), .A(\g.we_clk [9327]));
Q_ASSIGN U23448 ( .B(clk), .A(\g.we_clk [9326]));
Q_ASSIGN U23449 ( .B(clk), .A(\g.we_clk [9325]));
Q_ASSIGN U23450 ( .B(clk), .A(\g.we_clk [9324]));
Q_ASSIGN U23451 ( .B(clk), .A(\g.we_clk [9323]));
Q_ASSIGN U23452 ( .B(clk), .A(\g.we_clk [9322]));
Q_ASSIGN U23453 ( .B(clk), .A(\g.we_clk [9321]));
Q_ASSIGN U23454 ( .B(clk), .A(\g.we_clk [9320]));
Q_ASSIGN U23455 ( .B(clk), .A(\g.we_clk [9319]));
Q_ASSIGN U23456 ( .B(clk), .A(\g.we_clk [9318]));
Q_ASSIGN U23457 ( .B(clk), .A(\g.we_clk [9317]));
Q_ASSIGN U23458 ( .B(clk), .A(\g.we_clk [9316]));
Q_ASSIGN U23459 ( .B(clk), .A(\g.we_clk [9315]));
Q_ASSIGN U23460 ( .B(clk), .A(\g.we_clk [9314]));
Q_ASSIGN U23461 ( .B(clk), .A(\g.we_clk [9313]));
Q_ASSIGN U23462 ( .B(clk), .A(\g.we_clk [9312]));
Q_ASSIGN U23463 ( .B(clk), .A(\g.we_clk [9311]));
Q_ASSIGN U23464 ( .B(clk), .A(\g.we_clk [9310]));
Q_ASSIGN U23465 ( .B(clk), .A(\g.we_clk [9309]));
Q_ASSIGN U23466 ( .B(clk), .A(\g.we_clk [9308]));
Q_ASSIGN U23467 ( .B(clk), .A(\g.we_clk [9307]));
Q_ASSIGN U23468 ( .B(clk), .A(\g.we_clk [9306]));
Q_ASSIGN U23469 ( .B(clk), .A(\g.we_clk [9305]));
Q_ASSIGN U23470 ( .B(clk), .A(\g.we_clk [9304]));
Q_ASSIGN U23471 ( .B(clk), .A(\g.we_clk [9303]));
Q_ASSIGN U23472 ( .B(clk), .A(\g.we_clk [9302]));
Q_ASSIGN U23473 ( .B(clk), .A(\g.we_clk [9301]));
Q_ASSIGN U23474 ( .B(clk), .A(\g.we_clk [9300]));
Q_ASSIGN U23475 ( .B(clk), .A(\g.we_clk [9299]));
Q_ASSIGN U23476 ( .B(clk), .A(\g.we_clk [9298]));
Q_ASSIGN U23477 ( .B(clk), .A(\g.we_clk [9297]));
Q_ASSIGN U23478 ( .B(clk), .A(\g.we_clk [9296]));
Q_ASSIGN U23479 ( .B(clk), .A(\g.we_clk [9295]));
Q_ASSIGN U23480 ( .B(clk), .A(\g.we_clk [9294]));
Q_ASSIGN U23481 ( .B(clk), .A(\g.we_clk [9293]));
Q_ASSIGN U23482 ( .B(clk), .A(\g.we_clk [9292]));
Q_ASSIGN U23483 ( .B(clk), .A(\g.we_clk [9291]));
Q_ASSIGN U23484 ( .B(clk), .A(\g.we_clk [9290]));
Q_ASSIGN U23485 ( .B(clk), .A(\g.we_clk [9289]));
Q_ASSIGN U23486 ( .B(clk), .A(\g.we_clk [9288]));
Q_ASSIGN U23487 ( .B(clk), .A(\g.we_clk [9287]));
Q_ASSIGN U23488 ( .B(clk), .A(\g.we_clk [9286]));
Q_ASSIGN U23489 ( .B(clk), .A(\g.we_clk [9285]));
Q_ASSIGN U23490 ( .B(clk), .A(\g.we_clk [9284]));
Q_ASSIGN U23491 ( .B(clk), .A(\g.we_clk [9283]));
Q_ASSIGN U23492 ( .B(clk), .A(\g.we_clk [9282]));
Q_ASSIGN U23493 ( .B(clk), .A(\g.we_clk [9281]));
Q_ASSIGN U23494 ( .B(clk), .A(\g.we_clk [9280]));
Q_ASSIGN U23495 ( .B(clk), .A(\g.we_clk [9279]));
Q_ASSIGN U23496 ( .B(clk), .A(\g.we_clk [9278]));
Q_ASSIGN U23497 ( .B(clk), .A(\g.we_clk [9277]));
Q_ASSIGN U23498 ( .B(clk), .A(\g.we_clk [9276]));
Q_ASSIGN U23499 ( .B(clk), .A(\g.we_clk [9275]));
Q_ASSIGN U23500 ( .B(clk), .A(\g.we_clk [9274]));
Q_ASSIGN U23501 ( .B(clk), .A(\g.we_clk [9273]));
Q_ASSIGN U23502 ( .B(clk), .A(\g.we_clk [9272]));
Q_ASSIGN U23503 ( .B(clk), .A(\g.we_clk [9271]));
Q_ASSIGN U23504 ( .B(clk), .A(\g.we_clk [9270]));
Q_ASSIGN U23505 ( .B(clk), .A(\g.we_clk [9269]));
Q_ASSIGN U23506 ( .B(clk), .A(\g.we_clk [9268]));
Q_ASSIGN U23507 ( .B(clk), .A(\g.we_clk [9267]));
Q_ASSIGN U23508 ( .B(clk), .A(\g.we_clk [9266]));
Q_ASSIGN U23509 ( .B(clk), .A(\g.we_clk [9265]));
Q_ASSIGN U23510 ( .B(clk), .A(\g.we_clk [9264]));
Q_ASSIGN U23511 ( .B(clk), .A(\g.we_clk [9263]));
Q_ASSIGN U23512 ( .B(clk), .A(\g.we_clk [9262]));
Q_ASSIGN U23513 ( .B(clk), .A(\g.we_clk [9261]));
Q_ASSIGN U23514 ( .B(clk), .A(\g.we_clk [9260]));
Q_ASSIGN U23515 ( .B(clk), .A(\g.we_clk [9259]));
Q_ASSIGN U23516 ( .B(clk), .A(\g.we_clk [9258]));
Q_ASSIGN U23517 ( .B(clk), .A(\g.we_clk [9257]));
Q_ASSIGN U23518 ( .B(clk), .A(\g.we_clk [9256]));
Q_ASSIGN U23519 ( .B(clk), .A(\g.we_clk [9255]));
Q_ASSIGN U23520 ( .B(clk), .A(\g.we_clk [9254]));
Q_ASSIGN U23521 ( .B(clk), .A(\g.we_clk [9253]));
Q_ASSIGN U23522 ( .B(clk), .A(\g.we_clk [9252]));
Q_ASSIGN U23523 ( .B(clk), .A(\g.we_clk [9251]));
Q_ASSIGN U23524 ( .B(clk), .A(\g.we_clk [9250]));
Q_ASSIGN U23525 ( .B(clk), .A(\g.we_clk [9249]));
Q_ASSIGN U23526 ( .B(clk), .A(\g.we_clk [9248]));
Q_ASSIGN U23527 ( .B(clk), .A(\g.we_clk [9247]));
Q_ASSIGN U23528 ( .B(clk), .A(\g.we_clk [9246]));
Q_ASSIGN U23529 ( .B(clk), .A(\g.we_clk [9245]));
Q_ASSIGN U23530 ( .B(clk), .A(\g.we_clk [9244]));
Q_ASSIGN U23531 ( .B(clk), .A(\g.we_clk [9243]));
Q_ASSIGN U23532 ( .B(clk), .A(\g.we_clk [9242]));
Q_ASSIGN U23533 ( .B(clk), .A(\g.we_clk [9241]));
Q_ASSIGN U23534 ( .B(clk), .A(\g.we_clk [9240]));
Q_ASSIGN U23535 ( .B(clk), .A(\g.we_clk [9239]));
Q_ASSIGN U23536 ( .B(clk), .A(\g.we_clk [9238]));
Q_ASSIGN U23537 ( .B(clk), .A(\g.we_clk [9237]));
Q_ASSIGN U23538 ( .B(clk), .A(\g.we_clk [9236]));
Q_ASSIGN U23539 ( .B(clk), .A(\g.we_clk [9235]));
Q_ASSIGN U23540 ( .B(clk), .A(\g.we_clk [9234]));
Q_ASSIGN U23541 ( .B(clk), .A(\g.we_clk [9233]));
Q_ASSIGN U23542 ( .B(clk), .A(\g.we_clk [9232]));
Q_ASSIGN U23543 ( .B(clk), .A(\g.we_clk [9231]));
Q_ASSIGN U23544 ( .B(clk), .A(\g.we_clk [9230]));
Q_ASSIGN U23545 ( .B(clk), .A(\g.we_clk [9229]));
Q_ASSIGN U23546 ( .B(clk), .A(\g.we_clk [9228]));
Q_ASSIGN U23547 ( .B(clk), .A(\g.we_clk [9227]));
Q_ASSIGN U23548 ( .B(clk), .A(\g.we_clk [9226]));
Q_ASSIGN U23549 ( .B(clk), .A(\g.we_clk [9225]));
Q_ASSIGN U23550 ( .B(clk), .A(\g.we_clk [9224]));
Q_ASSIGN U23551 ( .B(clk), .A(\g.we_clk [9223]));
Q_ASSIGN U23552 ( .B(clk), .A(\g.we_clk [9222]));
Q_ASSIGN U23553 ( .B(clk), .A(\g.we_clk [9221]));
Q_ASSIGN U23554 ( .B(clk), .A(\g.we_clk [9220]));
Q_ASSIGN U23555 ( .B(clk), .A(\g.we_clk [9219]));
Q_ASSIGN U23556 ( .B(clk), .A(\g.we_clk [9218]));
Q_ASSIGN U23557 ( .B(clk), .A(\g.we_clk [9217]));
Q_ASSIGN U23558 ( .B(clk), .A(\g.we_clk [9216]));
Q_ASSIGN U23559 ( .B(clk), .A(\g.we_clk [9215]));
Q_ASSIGN U23560 ( .B(clk), .A(\g.we_clk [9214]));
Q_ASSIGN U23561 ( .B(clk), .A(\g.we_clk [9213]));
Q_ASSIGN U23562 ( .B(clk), .A(\g.we_clk [9212]));
Q_ASSIGN U23563 ( .B(clk), .A(\g.we_clk [9211]));
Q_ASSIGN U23564 ( .B(clk), .A(\g.we_clk [9210]));
Q_ASSIGN U23565 ( .B(clk), .A(\g.we_clk [9209]));
Q_ASSIGN U23566 ( .B(clk), .A(\g.we_clk [9208]));
Q_ASSIGN U23567 ( .B(clk), .A(\g.we_clk [9207]));
Q_ASSIGN U23568 ( .B(clk), .A(\g.we_clk [9206]));
Q_ASSIGN U23569 ( .B(clk), .A(\g.we_clk [9205]));
Q_ASSIGN U23570 ( .B(clk), .A(\g.we_clk [9204]));
Q_ASSIGN U23571 ( .B(clk), .A(\g.we_clk [9203]));
Q_ASSIGN U23572 ( .B(clk), .A(\g.we_clk [9202]));
Q_ASSIGN U23573 ( .B(clk), .A(\g.we_clk [9201]));
Q_ASSIGN U23574 ( .B(clk), .A(\g.we_clk [9200]));
Q_ASSIGN U23575 ( .B(clk), .A(\g.we_clk [9199]));
Q_ASSIGN U23576 ( .B(clk), .A(\g.we_clk [9198]));
Q_ASSIGN U23577 ( .B(clk), .A(\g.we_clk [9197]));
Q_ASSIGN U23578 ( .B(clk), .A(\g.we_clk [9196]));
Q_ASSIGN U23579 ( .B(clk), .A(\g.we_clk [9195]));
Q_ASSIGN U23580 ( .B(clk), .A(\g.we_clk [9194]));
Q_ASSIGN U23581 ( .B(clk), .A(\g.we_clk [9193]));
Q_ASSIGN U23582 ( .B(clk), .A(\g.we_clk [9192]));
Q_ASSIGN U23583 ( .B(clk), .A(\g.we_clk [9191]));
Q_ASSIGN U23584 ( .B(clk), .A(\g.we_clk [9190]));
Q_ASSIGN U23585 ( .B(clk), .A(\g.we_clk [9189]));
Q_ASSIGN U23586 ( .B(clk), .A(\g.we_clk [9188]));
Q_ASSIGN U23587 ( .B(clk), .A(\g.we_clk [9187]));
Q_ASSIGN U23588 ( .B(clk), .A(\g.we_clk [9186]));
Q_ASSIGN U23589 ( .B(clk), .A(\g.we_clk [9185]));
Q_ASSIGN U23590 ( .B(clk), .A(\g.we_clk [9184]));
Q_ASSIGN U23591 ( .B(clk), .A(\g.we_clk [9183]));
Q_ASSIGN U23592 ( .B(clk), .A(\g.we_clk [9182]));
Q_ASSIGN U23593 ( .B(clk), .A(\g.we_clk [9181]));
Q_ASSIGN U23594 ( .B(clk), .A(\g.we_clk [9180]));
Q_ASSIGN U23595 ( .B(clk), .A(\g.we_clk [9179]));
Q_ASSIGN U23596 ( .B(clk), .A(\g.we_clk [9178]));
Q_ASSIGN U23597 ( .B(clk), .A(\g.we_clk [9177]));
Q_ASSIGN U23598 ( .B(clk), .A(\g.we_clk [9176]));
Q_ASSIGN U23599 ( .B(clk), .A(\g.we_clk [9175]));
Q_ASSIGN U23600 ( .B(clk), .A(\g.we_clk [9174]));
Q_ASSIGN U23601 ( .B(clk), .A(\g.we_clk [9173]));
Q_ASSIGN U23602 ( .B(clk), .A(\g.we_clk [9172]));
Q_ASSIGN U23603 ( .B(clk), .A(\g.we_clk [9171]));
Q_ASSIGN U23604 ( .B(clk), .A(\g.we_clk [9170]));
Q_ASSIGN U23605 ( .B(clk), .A(\g.we_clk [9169]));
Q_ASSIGN U23606 ( .B(clk), .A(\g.we_clk [9168]));
Q_ASSIGN U23607 ( .B(clk), .A(\g.we_clk [9167]));
Q_ASSIGN U23608 ( .B(clk), .A(\g.we_clk [9166]));
Q_ASSIGN U23609 ( .B(clk), .A(\g.we_clk [9165]));
Q_ASSIGN U23610 ( .B(clk), .A(\g.we_clk [9164]));
Q_ASSIGN U23611 ( .B(clk), .A(\g.we_clk [9163]));
Q_ASSIGN U23612 ( .B(clk), .A(\g.we_clk [9162]));
Q_ASSIGN U23613 ( .B(clk), .A(\g.we_clk [9161]));
Q_ASSIGN U23614 ( .B(clk), .A(\g.we_clk [9160]));
Q_ASSIGN U23615 ( .B(clk), .A(\g.we_clk [9159]));
Q_ASSIGN U23616 ( .B(clk), .A(\g.we_clk [9158]));
Q_ASSIGN U23617 ( .B(clk), .A(\g.we_clk [9157]));
Q_ASSIGN U23618 ( .B(clk), .A(\g.we_clk [9156]));
Q_ASSIGN U23619 ( .B(clk), .A(\g.we_clk [9155]));
Q_ASSIGN U23620 ( .B(clk), .A(\g.we_clk [9154]));
Q_ASSIGN U23621 ( .B(clk), .A(\g.we_clk [9153]));
Q_ASSIGN U23622 ( .B(clk), .A(\g.we_clk [9152]));
Q_ASSIGN U23623 ( .B(clk), .A(\g.we_clk [9151]));
Q_ASSIGN U23624 ( .B(clk), .A(\g.we_clk [9150]));
Q_ASSIGN U23625 ( .B(clk), .A(\g.we_clk [9149]));
Q_ASSIGN U23626 ( .B(clk), .A(\g.we_clk [9148]));
Q_ASSIGN U23627 ( .B(clk), .A(\g.we_clk [9147]));
Q_ASSIGN U23628 ( .B(clk), .A(\g.we_clk [9146]));
Q_ASSIGN U23629 ( .B(clk), .A(\g.we_clk [9145]));
Q_ASSIGN U23630 ( .B(clk), .A(\g.we_clk [9144]));
Q_ASSIGN U23631 ( .B(clk), .A(\g.we_clk [9143]));
Q_ASSIGN U23632 ( .B(clk), .A(\g.we_clk [9142]));
Q_ASSIGN U23633 ( .B(clk), .A(\g.we_clk [9141]));
Q_ASSIGN U23634 ( .B(clk), .A(\g.we_clk [9140]));
Q_ASSIGN U23635 ( .B(clk), .A(\g.we_clk [9139]));
Q_ASSIGN U23636 ( .B(clk), .A(\g.we_clk [9138]));
Q_ASSIGN U23637 ( .B(clk), .A(\g.we_clk [9137]));
Q_ASSIGN U23638 ( .B(clk), .A(\g.we_clk [9136]));
Q_ASSIGN U23639 ( .B(clk), .A(\g.we_clk [9135]));
Q_ASSIGN U23640 ( .B(clk), .A(\g.we_clk [9134]));
Q_ASSIGN U23641 ( .B(clk), .A(\g.we_clk [9133]));
Q_ASSIGN U23642 ( .B(clk), .A(\g.we_clk [9132]));
Q_ASSIGN U23643 ( .B(clk), .A(\g.we_clk [9131]));
Q_ASSIGN U23644 ( .B(clk), .A(\g.we_clk [9130]));
Q_ASSIGN U23645 ( .B(clk), .A(\g.we_clk [9129]));
Q_ASSIGN U23646 ( .B(clk), .A(\g.we_clk [9128]));
Q_ASSIGN U23647 ( .B(clk), .A(\g.we_clk [9127]));
Q_ASSIGN U23648 ( .B(clk), .A(\g.we_clk [9126]));
Q_ASSIGN U23649 ( .B(clk), .A(\g.we_clk [9125]));
Q_ASSIGN U23650 ( .B(clk), .A(\g.we_clk [9124]));
Q_ASSIGN U23651 ( .B(clk), .A(\g.we_clk [9123]));
Q_ASSIGN U23652 ( .B(clk), .A(\g.we_clk [9122]));
Q_ASSIGN U23653 ( .B(clk), .A(\g.we_clk [9121]));
Q_ASSIGN U23654 ( .B(clk), .A(\g.we_clk [9120]));
Q_ASSIGN U23655 ( .B(clk), .A(\g.we_clk [9119]));
Q_ASSIGN U23656 ( .B(clk), .A(\g.we_clk [9118]));
Q_ASSIGN U23657 ( .B(clk), .A(\g.we_clk [9117]));
Q_ASSIGN U23658 ( .B(clk), .A(\g.we_clk [9116]));
Q_ASSIGN U23659 ( .B(clk), .A(\g.we_clk [9115]));
Q_ASSIGN U23660 ( .B(clk), .A(\g.we_clk [9114]));
Q_ASSIGN U23661 ( .B(clk), .A(\g.we_clk [9113]));
Q_ASSIGN U23662 ( .B(clk), .A(\g.we_clk [9112]));
Q_ASSIGN U23663 ( .B(clk), .A(\g.we_clk [9111]));
Q_ASSIGN U23664 ( .B(clk), .A(\g.we_clk [9110]));
Q_ASSIGN U23665 ( .B(clk), .A(\g.we_clk [9109]));
Q_ASSIGN U23666 ( .B(clk), .A(\g.we_clk [9108]));
Q_ASSIGN U23667 ( .B(clk), .A(\g.we_clk [9107]));
Q_ASSIGN U23668 ( .B(clk), .A(\g.we_clk [9106]));
Q_ASSIGN U23669 ( .B(clk), .A(\g.we_clk [9105]));
Q_ASSIGN U23670 ( .B(clk), .A(\g.we_clk [9104]));
Q_ASSIGN U23671 ( .B(clk), .A(\g.we_clk [9103]));
Q_ASSIGN U23672 ( .B(clk), .A(\g.we_clk [9102]));
Q_ASSIGN U23673 ( .B(clk), .A(\g.we_clk [9101]));
Q_ASSIGN U23674 ( .B(clk), .A(\g.we_clk [9100]));
Q_ASSIGN U23675 ( .B(clk), .A(\g.we_clk [9099]));
Q_ASSIGN U23676 ( .B(clk), .A(\g.we_clk [9098]));
Q_ASSIGN U23677 ( .B(clk), .A(\g.we_clk [9097]));
Q_ASSIGN U23678 ( .B(clk), .A(\g.we_clk [9096]));
Q_ASSIGN U23679 ( .B(clk), .A(\g.we_clk [9095]));
Q_ASSIGN U23680 ( .B(clk), .A(\g.we_clk [9094]));
Q_ASSIGN U23681 ( .B(clk), .A(\g.we_clk [9093]));
Q_ASSIGN U23682 ( .B(clk), .A(\g.we_clk [9092]));
Q_ASSIGN U23683 ( .B(clk), .A(\g.we_clk [9091]));
Q_ASSIGN U23684 ( .B(clk), .A(\g.we_clk [9090]));
Q_ASSIGN U23685 ( .B(clk), .A(\g.we_clk [9089]));
Q_ASSIGN U23686 ( .B(clk), .A(\g.we_clk [9088]));
Q_ASSIGN U23687 ( .B(clk), .A(\g.we_clk [9087]));
Q_ASSIGN U23688 ( .B(clk), .A(\g.we_clk [9086]));
Q_ASSIGN U23689 ( .B(clk), .A(\g.we_clk [9085]));
Q_ASSIGN U23690 ( .B(clk), .A(\g.we_clk [9084]));
Q_ASSIGN U23691 ( .B(clk), .A(\g.we_clk [9083]));
Q_ASSIGN U23692 ( .B(clk), .A(\g.we_clk [9082]));
Q_ASSIGN U23693 ( .B(clk), .A(\g.we_clk [9081]));
Q_ASSIGN U23694 ( .B(clk), .A(\g.we_clk [9080]));
Q_ASSIGN U23695 ( .B(clk), .A(\g.we_clk [9079]));
Q_ASSIGN U23696 ( .B(clk), .A(\g.we_clk [9078]));
Q_ASSIGN U23697 ( .B(clk), .A(\g.we_clk [9077]));
Q_ASSIGN U23698 ( .B(clk), .A(\g.we_clk [9076]));
Q_ASSIGN U23699 ( .B(clk), .A(\g.we_clk [9075]));
Q_ASSIGN U23700 ( .B(clk), .A(\g.we_clk [9074]));
Q_ASSIGN U23701 ( .B(clk), .A(\g.we_clk [9073]));
Q_ASSIGN U23702 ( .B(clk), .A(\g.we_clk [9072]));
Q_ASSIGN U23703 ( .B(clk), .A(\g.we_clk [9071]));
Q_ASSIGN U23704 ( .B(clk), .A(\g.we_clk [9070]));
Q_ASSIGN U23705 ( .B(clk), .A(\g.we_clk [9069]));
Q_ASSIGN U23706 ( .B(clk), .A(\g.we_clk [9068]));
Q_ASSIGN U23707 ( .B(clk), .A(\g.we_clk [9067]));
Q_ASSIGN U23708 ( .B(clk), .A(\g.we_clk [9066]));
Q_ASSIGN U23709 ( .B(clk), .A(\g.we_clk [9065]));
Q_ASSIGN U23710 ( .B(clk), .A(\g.we_clk [9064]));
Q_ASSIGN U23711 ( .B(clk), .A(\g.we_clk [9063]));
Q_ASSIGN U23712 ( .B(clk), .A(\g.we_clk [9062]));
Q_ASSIGN U23713 ( .B(clk), .A(\g.we_clk [9061]));
Q_ASSIGN U23714 ( .B(clk), .A(\g.we_clk [9060]));
Q_ASSIGN U23715 ( .B(clk), .A(\g.we_clk [9059]));
Q_ASSIGN U23716 ( .B(clk), .A(\g.we_clk [9058]));
Q_ASSIGN U23717 ( .B(clk), .A(\g.we_clk [9057]));
Q_ASSIGN U23718 ( .B(clk), .A(\g.we_clk [9056]));
Q_ASSIGN U23719 ( .B(clk), .A(\g.we_clk [9055]));
Q_ASSIGN U23720 ( .B(clk), .A(\g.we_clk [9054]));
Q_ASSIGN U23721 ( .B(clk), .A(\g.we_clk [9053]));
Q_ASSIGN U23722 ( .B(clk), .A(\g.we_clk [9052]));
Q_ASSIGN U23723 ( .B(clk), .A(\g.we_clk [9051]));
Q_ASSIGN U23724 ( .B(clk), .A(\g.we_clk [9050]));
Q_ASSIGN U23725 ( .B(clk), .A(\g.we_clk [9049]));
Q_ASSIGN U23726 ( .B(clk), .A(\g.we_clk [9048]));
Q_ASSIGN U23727 ( .B(clk), .A(\g.we_clk [9047]));
Q_ASSIGN U23728 ( .B(clk), .A(\g.we_clk [9046]));
Q_ASSIGN U23729 ( .B(clk), .A(\g.we_clk [9045]));
Q_ASSIGN U23730 ( .B(clk), .A(\g.we_clk [9044]));
Q_ASSIGN U23731 ( .B(clk), .A(\g.we_clk [9043]));
Q_ASSIGN U23732 ( .B(clk), .A(\g.we_clk [9042]));
Q_ASSIGN U23733 ( .B(clk), .A(\g.we_clk [9041]));
Q_ASSIGN U23734 ( .B(clk), .A(\g.we_clk [9040]));
Q_ASSIGN U23735 ( .B(clk), .A(\g.we_clk [9039]));
Q_ASSIGN U23736 ( .B(clk), .A(\g.we_clk [9038]));
Q_ASSIGN U23737 ( .B(clk), .A(\g.we_clk [9037]));
Q_ASSIGN U23738 ( .B(clk), .A(\g.we_clk [9036]));
Q_ASSIGN U23739 ( .B(clk), .A(\g.we_clk [9035]));
Q_ASSIGN U23740 ( .B(clk), .A(\g.we_clk [9034]));
Q_ASSIGN U23741 ( .B(clk), .A(\g.we_clk [9033]));
Q_ASSIGN U23742 ( .B(clk), .A(\g.we_clk [9032]));
Q_ASSIGN U23743 ( .B(clk), .A(\g.we_clk [9031]));
Q_ASSIGN U23744 ( .B(clk), .A(\g.we_clk [9030]));
Q_ASSIGN U23745 ( .B(clk), .A(\g.we_clk [9029]));
Q_ASSIGN U23746 ( .B(clk), .A(\g.we_clk [9028]));
Q_ASSIGN U23747 ( .B(clk), .A(\g.we_clk [9027]));
Q_ASSIGN U23748 ( .B(clk), .A(\g.we_clk [9026]));
Q_ASSIGN U23749 ( .B(clk), .A(\g.we_clk [9025]));
Q_ASSIGN U23750 ( .B(clk), .A(\g.we_clk [9024]));
Q_ASSIGN U23751 ( .B(clk), .A(\g.we_clk [9023]));
Q_ASSIGN U23752 ( .B(clk), .A(\g.we_clk [9022]));
Q_ASSIGN U23753 ( .B(clk), .A(\g.we_clk [9021]));
Q_ASSIGN U23754 ( .B(clk), .A(\g.we_clk [9020]));
Q_ASSIGN U23755 ( .B(clk), .A(\g.we_clk [9019]));
Q_ASSIGN U23756 ( .B(clk), .A(\g.we_clk [9018]));
Q_ASSIGN U23757 ( .B(clk), .A(\g.we_clk [9017]));
Q_ASSIGN U23758 ( .B(clk), .A(\g.we_clk [9016]));
Q_ASSIGN U23759 ( .B(clk), .A(\g.we_clk [9015]));
Q_ASSIGN U23760 ( .B(clk), .A(\g.we_clk [9014]));
Q_ASSIGN U23761 ( .B(clk), .A(\g.we_clk [9013]));
Q_ASSIGN U23762 ( .B(clk), .A(\g.we_clk [9012]));
Q_ASSIGN U23763 ( .B(clk), .A(\g.we_clk [9011]));
Q_ASSIGN U23764 ( .B(clk), .A(\g.we_clk [9010]));
Q_ASSIGN U23765 ( .B(clk), .A(\g.we_clk [9009]));
Q_ASSIGN U23766 ( .B(clk), .A(\g.we_clk [9008]));
Q_ASSIGN U23767 ( .B(clk), .A(\g.we_clk [9007]));
Q_ASSIGN U23768 ( .B(clk), .A(\g.we_clk [9006]));
Q_ASSIGN U23769 ( .B(clk), .A(\g.we_clk [9005]));
Q_ASSIGN U23770 ( .B(clk), .A(\g.we_clk [9004]));
Q_ASSIGN U23771 ( .B(clk), .A(\g.we_clk [9003]));
Q_ASSIGN U23772 ( .B(clk), .A(\g.we_clk [9002]));
Q_ASSIGN U23773 ( .B(clk), .A(\g.we_clk [9001]));
Q_ASSIGN U23774 ( .B(clk), .A(\g.we_clk [9000]));
Q_ASSIGN U23775 ( .B(clk), .A(\g.we_clk [8999]));
Q_ASSIGN U23776 ( .B(clk), .A(\g.we_clk [8998]));
Q_ASSIGN U23777 ( .B(clk), .A(\g.we_clk [8997]));
Q_ASSIGN U23778 ( .B(clk), .A(\g.we_clk [8996]));
Q_ASSIGN U23779 ( .B(clk), .A(\g.we_clk [8995]));
Q_ASSIGN U23780 ( .B(clk), .A(\g.we_clk [8994]));
Q_ASSIGN U23781 ( .B(clk), .A(\g.we_clk [8993]));
Q_ASSIGN U23782 ( .B(clk), .A(\g.we_clk [8992]));
Q_ASSIGN U23783 ( .B(clk), .A(\g.we_clk [8991]));
Q_ASSIGN U23784 ( .B(clk), .A(\g.we_clk [8990]));
Q_ASSIGN U23785 ( .B(clk), .A(\g.we_clk [8989]));
Q_ASSIGN U23786 ( .B(clk), .A(\g.we_clk [8988]));
Q_ASSIGN U23787 ( .B(clk), .A(\g.we_clk [8987]));
Q_ASSIGN U23788 ( .B(clk), .A(\g.we_clk [8986]));
Q_ASSIGN U23789 ( .B(clk), .A(\g.we_clk [8985]));
Q_ASSIGN U23790 ( .B(clk), .A(\g.we_clk [8984]));
Q_ASSIGN U23791 ( .B(clk), .A(\g.we_clk [8983]));
Q_ASSIGN U23792 ( .B(clk), .A(\g.we_clk [8982]));
Q_ASSIGN U23793 ( .B(clk), .A(\g.we_clk [8981]));
Q_ASSIGN U23794 ( .B(clk), .A(\g.we_clk [8980]));
Q_ASSIGN U23795 ( .B(clk), .A(\g.we_clk [8979]));
Q_ASSIGN U23796 ( .B(clk), .A(\g.we_clk [8978]));
Q_ASSIGN U23797 ( .B(clk), .A(\g.we_clk [8977]));
Q_ASSIGN U23798 ( .B(clk), .A(\g.we_clk [8976]));
Q_ASSIGN U23799 ( .B(clk), .A(\g.we_clk [8975]));
Q_ASSIGN U23800 ( .B(clk), .A(\g.we_clk [8974]));
Q_ASSIGN U23801 ( .B(clk), .A(\g.we_clk [8973]));
Q_ASSIGN U23802 ( .B(clk), .A(\g.we_clk [8972]));
Q_ASSIGN U23803 ( .B(clk), .A(\g.we_clk [8971]));
Q_ASSIGN U23804 ( .B(clk), .A(\g.we_clk [8970]));
Q_ASSIGN U23805 ( .B(clk), .A(\g.we_clk [8969]));
Q_ASSIGN U23806 ( .B(clk), .A(\g.we_clk [8968]));
Q_ASSIGN U23807 ( .B(clk), .A(\g.we_clk [8967]));
Q_ASSIGN U23808 ( .B(clk), .A(\g.we_clk [8966]));
Q_ASSIGN U23809 ( .B(clk), .A(\g.we_clk [8965]));
Q_ASSIGN U23810 ( .B(clk), .A(\g.we_clk [8964]));
Q_ASSIGN U23811 ( .B(clk), .A(\g.we_clk [8963]));
Q_ASSIGN U23812 ( .B(clk), .A(\g.we_clk [8962]));
Q_ASSIGN U23813 ( .B(clk), .A(\g.we_clk [8961]));
Q_ASSIGN U23814 ( .B(clk), .A(\g.we_clk [8960]));
Q_ASSIGN U23815 ( .B(clk), .A(\g.we_clk [8959]));
Q_ASSIGN U23816 ( .B(clk), .A(\g.we_clk [8958]));
Q_ASSIGN U23817 ( .B(clk), .A(\g.we_clk [8957]));
Q_ASSIGN U23818 ( .B(clk), .A(\g.we_clk [8956]));
Q_ASSIGN U23819 ( .B(clk), .A(\g.we_clk [8955]));
Q_ASSIGN U23820 ( .B(clk), .A(\g.we_clk [8954]));
Q_ASSIGN U23821 ( .B(clk), .A(\g.we_clk [8953]));
Q_ASSIGN U23822 ( .B(clk), .A(\g.we_clk [8952]));
Q_ASSIGN U23823 ( .B(clk), .A(\g.we_clk [8951]));
Q_ASSIGN U23824 ( .B(clk), .A(\g.we_clk [8950]));
Q_ASSIGN U23825 ( .B(clk), .A(\g.we_clk [8949]));
Q_ASSIGN U23826 ( .B(clk), .A(\g.we_clk [8948]));
Q_ASSIGN U23827 ( .B(clk), .A(\g.we_clk [8947]));
Q_ASSIGN U23828 ( .B(clk), .A(\g.we_clk [8946]));
Q_ASSIGN U23829 ( .B(clk), .A(\g.we_clk [8945]));
Q_ASSIGN U23830 ( .B(clk), .A(\g.we_clk [8944]));
Q_ASSIGN U23831 ( .B(clk), .A(\g.we_clk [8943]));
Q_ASSIGN U23832 ( .B(clk), .A(\g.we_clk [8942]));
Q_ASSIGN U23833 ( .B(clk), .A(\g.we_clk [8941]));
Q_ASSIGN U23834 ( .B(clk), .A(\g.we_clk [8940]));
Q_ASSIGN U23835 ( .B(clk), .A(\g.we_clk [8939]));
Q_ASSIGN U23836 ( .B(clk), .A(\g.we_clk [8938]));
Q_ASSIGN U23837 ( .B(clk), .A(\g.we_clk [8937]));
Q_ASSIGN U23838 ( .B(clk), .A(\g.we_clk [8936]));
Q_ASSIGN U23839 ( .B(clk), .A(\g.we_clk [8935]));
Q_ASSIGN U23840 ( .B(clk), .A(\g.we_clk [8934]));
Q_ASSIGN U23841 ( .B(clk), .A(\g.we_clk [8933]));
Q_ASSIGN U23842 ( .B(clk), .A(\g.we_clk [8932]));
Q_ASSIGN U23843 ( .B(clk), .A(\g.we_clk [8931]));
Q_ASSIGN U23844 ( .B(clk), .A(\g.we_clk [8930]));
Q_ASSIGN U23845 ( .B(clk), .A(\g.we_clk [8929]));
Q_ASSIGN U23846 ( .B(clk), .A(\g.we_clk [8928]));
Q_ASSIGN U23847 ( .B(clk), .A(\g.we_clk [8927]));
Q_ASSIGN U23848 ( .B(clk), .A(\g.we_clk [8926]));
Q_ASSIGN U23849 ( .B(clk), .A(\g.we_clk [8925]));
Q_ASSIGN U23850 ( .B(clk), .A(\g.we_clk [8924]));
Q_ASSIGN U23851 ( .B(clk), .A(\g.we_clk [8923]));
Q_ASSIGN U23852 ( .B(clk), .A(\g.we_clk [8922]));
Q_ASSIGN U23853 ( .B(clk), .A(\g.we_clk [8921]));
Q_ASSIGN U23854 ( .B(clk), .A(\g.we_clk [8920]));
Q_ASSIGN U23855 ( .B(clk), .A(\g.we_clk [8919]));
Q_ASSIGN U23856 ( .B(clk), .A(\g.we_clk [8918]));
Q_ASSIGN U23857 ( .B(clk), .A(\g.we_clk [8917]));
Q_ASSIGN U23858 ( .B(clk), .A(\g.we_clk [8916]));
Q_ASSIGN U23859 ( .B(clk), .A(\g.we_clk [8915]));
Q_ASSIGN U23860 ( .B(clk), .A(\g.we_clk [8914]));
Q_ASSIGN U23861 ( .B(clk), .A(\g.we_clk [8913]));
Q_ASSIGN U23862 ( .B(clk), .A(\g.we_clk [8912]));
Q_ASSIGN U23863 ( .B(clk), .A(\g.we_clk [8911]));
Q_ASSIGN U23864 ( .B(clk), .A(\g.we_clk [8910]));
Q_ASSIGN U23865 ( .B(clk), .A(\g.we_clk [8909]));
Q_ASSIGN U23866 ( .B(clk), .A(\g.we_clk [8908]));
Q_ASSIGN U23867 ( .B(clk), .A(\g.we_clk [8907]));
Q_ASSIGN U23868 ( .B(clk), .A(\g.we_clk [8906]));
Q_ASSIGN U23869 ( .B(clk), .A(\g.we_clk [8905]));
Q_ASSIGN U23870 ( .B(clk), .A(\g.we_clk [8904]));
Q_ASSIGN U23871 ( .B(clk), .A(\g.we_clk [8903]));
Q_ASSIGN U23872 ( .B(clk), .A(\g.we_clk [8902]));
Q_ASSIGN U23873 ( .B(clk), .A(\g.we_clk [8901]));
Q_ASSIGN U23874 ( .B(clk), .A(\g.we_clk [8900]));
Q_ASSIGN U23875 ( .B(clk), .A(\g.we_clk [8899]));
Q_ASSIGN U23876 ( .B(clk), .A(\g.we_clk [8898]));
Q_ASSIGN U23877 ( .B(clk), .A(\g.we_clk [8897]));
Q_ASSIGN U23878 ( .B(clk), .A(\g.we_clk [8896]));
Q_ASSIGN U23879 ( .B(clk), .A(\g.we_clk [8895]));
Q_ASSIGN U23880 ( .B(clk), .A(\g.we_clk [8894]));
Q_ASSIGN U23881 ( .B(clk), .A(\g.we_clk [8893]));
Q_ASSIGN U23882 ( .B(clk), .A(\g.we_clk [8892]));
Q_ASSIGN U23883 ( .B(clk), .A(\g.we_clk [8891]));
Q_ASSIGN U23884 ( .B(clk), .A(\g.we_clk [8890]));
Q_ASSIGN U23885 ( .B(clk), .A(\g.we_clk [8889]));
Q_ASSIGN U23886 ( .B(clk), .A(\g.we_clk [8888]));
Q_ASSIGN U23887 ( .B(clk), .A(\g.we_clk [8887]));
Q_ASSIGN U23888 ( .B(clk), .A(\g.we_clk [8886]));
Q_ASSIGN U23889 ( .B(clk), .A(\g.we_clk [8885]));
Q_ASSIGN U23890 ( .B(clk), .A(\g.we_clk [8884]));
Q_ASSIGN U23891 ( .B(clk), .A(\g.we_clk [8883]));
Q_ASSIGN U23892 ( .B(clk), .A(\g.we_clk [8882]));
Q_ASSIGN U23893 ( .B(clk), .A(\g.we_clk [8881]));
Q_ASSIGN U23894 ( .B(clk), .A(\g.we_clk [8880]));
Q_ASSIGN U23895 ( .B(clk), .A(\g.we_clk [8879]));
Q_ASSIGN U23896 ( .B(clk), .A(\g.we_clk [8878]));
Q_ASSIGN U23897 ( .B(clk), .A(\g.we_clk [8877]));
Q_ASSIGN U23898 ( .B(clk), .A(\g.we_clk [8876]));
Q_ASSIGN U23899 ( .B(clk), .A(\g.we_clk [8875]));
Q_ASSIGN U23900 ( .B(clk), .A(\g.we_clk [8874]));
Q_ASSIGN U23901 ( .B(clk), .A(\g.we_clk [8873]));
Q_ASSIGN U23902 ( .B(clk), .A(\g.we_clk [8872]));
Q_ASSIGN U23903 ( .B(clk), .A(\g.we_clk [8871]));
Q_ASSIGN U23904 ( .B(clk), .A(\g.we_clk [8870]));
Q_ASSIGN U23905 ( .B(clk), .A(\g.we_clk [8869]));
Q_ASSIGN U23906 ( .B(clk), .A(\g.we_clk [8868]));
Q_ASSIGN U23907 ( .B(clk), .A(\g.we_clk [8867]));
Q_ASSIGN U23908 ( .B(clk), .A(\g.we_clk [8866]));
Q_ASSIGN U23909 ( .B(clk), .A(\g.we_clk [8865]));
Q_ASSIGN U23910 ( .B(clk), .A(\g.we_clk [8864]));
Q_ASSIGN U23911 ( .B(clk), .A(\g.we_clk [8863]));
Q_ASSIGN U23912 ( .B(clk), .A(\g.we_clk [8862]));
Q_ASSIGN U23913 ( .B(clk), .A(\g.we_clk [8861]));
Q_ASSIGN U23914 ( .B(clk), .A(\g.we_clk [8860]));
Q_ASSIGN U23915 ( .B(clk), .A(\g.we_clk [8859]));
Q_ASSIGN U23916 ( .B(clk), .A(\g.we_clk [8858]));
Q_ASSIGN U23917 ( .B(clk), .A(\g.we_clk [8857]));
Q_ASSIGN U23918 ( .B(clk), .A(\g.we_clk [8856]));
Q_ASSIGN U23919 ( .B(clk), .A(\g.we_clk [8855]));
Q_ASSIGN U23920 ( .B(clk), .A(\g.we_clk [8854]));
Q_ASSIGN U23921 ( .B(clk), .A(\g.we_clk [8853]));
Q_ASSIGN U23922 ( .B(clk), .A(\g.we_clk [8852]));
Q_ASSIGN U23923 ( .B(clk), .A(\g.we_clk [8851]));
Q_ASSIGN U23924 ( .B(clk), .A(\g.we_clk [8850]));
Q_ASSIGN U23925 ( .B(clk), .A(\g.we_clk [8849]));
Q_ASSIGN U23926 ( .B(clk), .A(\g.we_clk [8848]));
Q_ASSIGN U23927 ( .B(clk), .A(\g.we_clk [8847]));
Q_ASSIGN U23928 ( .B(clk), .A(\g.we_clk [8846]));
Q_ASSIGN U23929 ( .B(clk), .A(\g.we_clk [8845]));
Q_ASSIGN U23930 ( .B(clk), .A(\g.we_clk [8844]));
Q_ASSIGN U23931 ( .B(clk), .A(\g.we_clk [8843]));
Q_ASSIGN U23932 ( .B(clk), .A(\g.we_clk [8842]));
Q_ASSIGN U23933 ( .B(clk), .A(\g.we_clk [8841]));
Q_ASSIGN U23934 ( .B(clk), .A(\g.we_clk [8840]));
Q_ASSIGN U23935 ( .B(clk), .A(\g.we_clk [8839]));
Q_ASSIGN U23936 ( .B(clk), .A(\g.we_clk [8838]));
Q_ASSIGN U23937 ( .B(clk), .A(\g.we_clk [8837]));
Q_ASSIGN U23938 ( .B(clk), .A(\g.we_clk [8836]));
Q_ASSIGN U23939 ( .B(clk), .A(\g.we_clk [8835]));
Q_ASSIGN U23940 ( .B(clk), .A(\g.we_clk [8834]));
Q_ASSIGN U23941 ( .B(clk), .A(\g.we_clk [8833]));
Q_ASSIGN U23942 ( .B(clk), .A(\g.we_clk [8832]));
Q_ASSIGN U23943 ( .B(clk), .A(\g.we_clk [8831]));
Q_ASSIGN U23944 ( .B(clk), .A(\g.we_clk [8830]));
Q_ASSIGN U23945 ( .B(clk), .A(\g.we_clk [8829]));
Q_ASSIGN U23946 ( .B(clk), .A(\g.we_clk [8828]));
Q_ASSIGN U23947 ( .B(clk), .A(\g.we_clk [8827]));
Q_ASSIGN U23948 ( .B(clk), .A(\g.we_clk [8826]));
Q_ASSIGN U23949 ( .B(clk), .A(\g.we_clk [8825]));
Q_ASSIGN U23950 ( .B(clk), .A(\g.we_clk [8824]));
Q_ASSIGN U23951 ( .B(clk), .A(\g.we_clk [8823]));
Q_ASSIGN U23952 ( .B(clk), .A(\g.we_clk [8822]));
Q_ASSIGN U23953 ( .B(clk), .A(\g.we_clk [8821]));
Q_ASSIGN U23954 ( .B(clk), .A(\g.we_clk [8820]));
Q_ASSIGN U23955 ( .B(clk), .A(\g.we_clk [8819]));
Q_ASSIGN U23956 ( .B(clk), .A(\g.we_clk [8818]));
Q_ASSIGN U23957 ( .B(clk), .A(\g.we_clk [8817]));
Q_ASSIGN U23958 ( .B(clk), .A(\g.we_clk [8816]));
Q_ASSIGN U23959 ( .B(clk), .A(\g.we_clk [8815]));
Q_ASSIGN U23960 ( .B(clk), .A(\g.we_clk [8814]));
Q_ASSIGN U23961 ( .B(clk), .A(\g.we_clk [8813]));
Q_ASSIGN U23962 ( .B(clk), .A(\g.we_clk [8812]));
Q_ASSIGN U23963 ( .B(clk), .A(\g.we_clk [8811]));
Q_ASSIGN U23964 ( .B(clk), .A(\g.we_clk [8810]));
Q_ASSIGN U23965 ( .B(clk), .A(\g.we_clk [8809]));
Q_ASSIGN U23966 ( .B(clk), .A(\g.we_clk [8808]));
Q_ASSIGN U23967 ( .B(clk), .A(\g.we_clk [8807]));
Q_ASSIGN U23968 ( .B(clk), .A(\g.we_clk [8806]));
Q_ASSIGN U23969 ( .B(clk), .A(\g.we_clk [8805]));
Q_ASSIGN U23970 ( .B(clk), .A(\g.we_clk [8804]));
Q_ASSIGN U23971 ( .B(clk), .A(\g.we_clk [8803]));
Q_ASSIGN U23972 ( .B(clk), .A(\g.we_clk [8802]));
Q_ASSIGN U23973 ( .B(clk), .A(\g.we_clk [8801]));
Q_ASSIGN U23974 ( .B(clk), .A(\g.we_clk [8800]));
Q_ASSIGN U23975 ( .B(clk), .A(\g.we_clk [8799]));
Q_ASSIGN U23976 ( .B(clk), .A(\g.we_clk [8798]));
Q_ASSIGN U23977 ( .B(clk), .A(\g.we_clk [8797]));
Q_ASSIGN U23978 ( .B(clk), .A(\g.we_clk [8796]));
Q_ASSIGN U23979 ( .B(clk), .A(\g.we_clk [8795]));
Q_ASSIGN U23980 ( .B(clk), .A(\g.we_clk [8794]));
Q_ASSIGN U23981 ( .B(clk), .A(\g.we_clk [8793]));
Q_ASSIGN U23982 ( .B(clk), .A(\g.we_clk [8792]));
Q_ASSIGN U23983 ( .B(clk), .A(\g.we_clk [8791]));
Q_ASSIGN U23984 ( .B(clk), .A(\g.we_clk [8790]));
Q_ASSIGN U23985 ( .B(clk), .A(\g.we_clk [8789]));
Q_ASSIGN U23986 ( .B(clk), .A(\g.we_clk [8788]));
Q_ASSIGN U23987 ( .B(clk), .A(\g.we_clk [8787]));
Q_ASSIGN U23988 ( .B(clk), .A(\g.we_clk [8786]));
Q_ASSIGN U23989 ( .B(clk), .A(\g.we_clk [8785]));
Q_ASSIGN U23990 ( .B(clk), .A(\g.we_clk [8784]));
Q_ASSIGN U23991 ( .B(clk), .A(\g.we_clk [8783]));
Q_ASSIGN U23992 ( .B(clk), .A(\g.we_clk [8782]));
Q_ASSIGN U23993 ( .B(clk), .A(\g.we_clk [8781]));
Q_ASSIGN U23994 ( .B(clk), .A(\g.we_clk [8780]));
Q_ASSIGN U23995 ( .B(clk), .A(\g.we_clk [8779]));
Q_ASSIGN U23996 ( .B(clk), .A(\g.we_clk [8778]));
Q_ASSIGN U23997 ( .B(clk), .A(\g.we_clk [8777]));
Q_ASSIGN U23998 ( .B(clk), .A(\g.we_clk [8776]));
Q_ASSIGN U23999 ( .B(clk), .A(\g.we_clk [8775]));
Q_ASSIGN U24000 ( .B(clk), .A(\g.we_clk [8774]));
Q_ASSIGN U24001 ( .B(clk), .A(\g.we_clk [8773]));
Q_ASSIGN U24002 ( .B(clk), .A(\g.we_clk [8772]));
Q_ASSIGN U24003 ( .B(clk), .A(\g.we_clk [8771]));
Q_ASSIGN U24004 ( .B(clk), .A(\g.we_clk [8770]));
Q_ASSIGN U24005 ( .B(clk), .A(\g.we_clk [8769]));
Q_ASSIGN U24006 ( .B(clk), .A(\g.we_clk [8768]));
Q_ASSIGN U24007 ( .B(clk), .A(\g.we_clk [8767]));
Q_ASSIGN U24008 ( .B(clk), .A(\g.we_clk [8766]));
Q_ASSIGN U24009 ( .B(clk), .A(\g.we_clk [8765]));
Q_ASSIGN U24010 ( .B(clk), .A(\g.we_clk [8764]));
Q_ASSIGN U24011 ( .B(clk), .A(\g.we_clk [8763]));
Q_ASSIGN U24012 ( .B(clk), .A(\g.we_clk [8762]));
Q_ASSIGN U24013 ( .B(clk), .A(\g.we_clk [8761]));
Q_ASSIGN U24014 ( .B(clk), .A(\g.we_clk [8760]));
Q_ASSIGN U24015 ( .B(clk), .A(\g.we_clk [8759]));
Q_ASSIGN U24016 ( .B(clk), .A(\g.we_clk [8758]));
Q_ASSIGN U24017 ( .B(clk), .A(\g.we_clk [8757]));
Q_ASSIGN U24018 ( .B(clk), .A(\g.we_clk [8756]));
Q_ASSIGN U24019 ( .B(clk), .A(\g.we_clk [8755]));
Q_ASSIGN U24020 ( .B(clk), .A(\g.we_clk [8754]));
Q_ASSIGN U24021 ( .B(clk), .A(\g.we_clk [8753]));
Q_ASSIGN U24022 ( .B(clk), .A(\g.we_clk [8752]));
Q_ASSIGN U24023 ( .B(clk), .A(\g.we_clk [8751]));
Q_ASSIGN U24024 ( .B(clk), .A(\g.we_clk [8750]));
Q_ASSIGN U24025 ( .B(clk), .A(\g.we_clk [8749]));
Q_ASSIGN U24026 ( .B(clk), .A(\g.we_clk [8748]));
Q_ASSIGN U24027 ( .B(clk), .A(\g.we_clk [8747]));
Q_ASSIGN U24028 ( .B(clk), .A(\g.we_clk [8746]));
Q_ASSIGN U24029 ( .B(clk), .A(\g.we_clk [8745]));
Q_ASSIGN U24030 ( .B(clk), .A(\g.we_clk [8744]));
Q_ASSIGN U24031 ( .B(clk), .A(\g.we_clk [8743]));
Q_ASSIGN U24032 ( .B(clk), .A(\g.we_clk [8742]));
Q_ASSIGN U24033 ( .B(clk), .A(\g.we_clk [8741]));
Q_ASSIGN U24034 ( .B(clk), .A(\g.we_clk [8740]));
Q_ASSIGN U24035 ( .B(clk), .A(\g.we_clk [8739]));
Q_ASSIGN U24036 ( .B(clk), .A(\g.we_clk [8738]));
Q_ASSIGN U24037 ( .B(clk), .A(\g.we_clk [8737]));
Q_ASSIGN U24038 ( .B(clk), .A(\g.we_clk [8736]));
Q_ASSIGN U24039 ( .B(clk), .A(\g.we_clk [8735]));
Q_ASSIGN U24040 ( .B(clk), .A(\g.we_clk [8734]));
Q_ASSIGN U24041 ( .B(clk), .A(\g.we_clk [8733]));
Q_ASSIGN U24042 ( .B(clk), .A(\g.we_clk [8732]));
Q_ASSIGN U24043 ( .B(clk), .A(\g.we_clk [8731]));
Q_ASSIGN U24044 ( .B(clk), .A(\g.we_clk [8730]));
Q_ASSIGN U24045 ( .B(clk), .A(\g.we_clk [8729]));
Q_ASSIGN U24046 ( .B(clk), .A(\g.we_clk [8728]));
Q_ASSIGN U24047 ( .B(clk), .A(\g.we_clk [8727]));
Q_ASSIGN U24048 ( .B(clk), .A(\g.we_clk [8726]));
Q_ASSIGN U24049 ( .B(clk), .A(\g.we_clk [8725]));
Q_ASSIGN U24050 ( .B(clk), .A(\g.we_clk [8724]));
Q_ASSIGN U24051 ( .B(clk), .A(\g.we_clk [8723]));
Q_ASSIGN U24052 ( .B(clk), .A(\g.we_clk [8722]));
Q_ASSIGN U24053 ( .B(clk), .A(\g.we_clk [8721]));
Q_ASSIGN U24054 ( .B(clk), .A(\g.we_clk [8720]));
Q_ASSIGN U24055 ( .B(clk), .A(\g.we_clk [8719]));
Q_ASSIGN U24056 ( .B(clk), .A(\g.we_clk [8718]));
Q_ASSIGN U24057 ( .B(clk), .A(\g.we_clk [8717]));
Q_ASSIGN U24058 ( .B(clk), .A(\g.we_clk [8716]));
Q_ASSIGN U24059 ( .B(clk), .A(\g.we_clk [8715]));
Q_ASSIGN U24060 ( .B(clk), .A(\g.we_clk [8714]));
Q_ASSIGN U24061 ( .B(clk), .A(\g.we_clk [8713]));
Q_ASSIGN U24062 ( .B(clk), .A(\g.we_clk [8712]));
Q_ASSIGN U24063 ( .B(clk), .A(\g.we_clk [8711]));
Q_ASSIGN U24064 ( .B(clk), .A(\g.we_clk [8710]));
Q_ASSIGN U24065 ( .B(clk), .A(\g.we_clk [8709]));
Q_ASSIGN U24066 ( .B(clk), .A(\g.we_clk [8708]));
Q_ASSIGN U24067 ( .B(clk), .A(\g.we_clk [8707]));
Q_ASSIGN U24068 ( .B(clk), .A(\g.we_clk [8706]));
Q_ASSIGN U24069 ( .B(clk), .A(\g.we_clk [8705]));
Q_ASSIGN U24070 ( .B(clk), .A(\g.we_clk [8704]));
Q_ASSIGN U24071 ( .B(clk), .A(\g.we_clk [8703]));
Q_ASSIGN U24072 ( .B(clk), .A(\g.we_clk [8702]));
Q_ASSIGN U24073 ( .B(clk), .A(\g.we_clk [8701]));
Q_ASSIGN U24074 ( .B(clk), .A(\g.we_clk [8700]));
Q_ASSIGN U24075 ( .B(clk), .A(\g.we_clk [8699]));
Q_ASSIGN U24076 ( .B(clk), .A(\g.we_clk [8698]));
Q_ASSIGN U24077 ( .B(clk), .A(\g.we_clk [8697]));
Q_ASSIGN U24078 ( .B(clk), .A(\g.we_clk [8696]));
Q_ASSIGN U24079 ( .B(clk), .A(\g.we_clk [8695]));
Q_ASSIGN U24080 ( .B(clk), .A(\g.we_clk [8694]));
Q_ASSIGN U24081 ( .B(clk), .A(\g.we_clk [8693]));
Q_ASSIGN U24082 ( .B(clk), .A(\g.we_clk [8692]));
Q_ASSIGN U24083 ( .B(clk), .A(\g.we_clk [8691]));
Q_ASSIGN U24084 ( .B(clk), .A(\g.we_clk [8690]));
Q_ASSIGN U24085 ( .B(clk), .A(\g.we_clk [8689]));
Q_ASSIGN U24086 ( .B(clk), .A(\g.we_clk [8688]));
Q_ASSIGN U24087 ( .B(clk), .A(\g.we_clk [8687]));
Q_ASSIGN U24088 ( .B(clk), .A(\g.we_clk [8686]));
Q_ASSIGN U24089 ( .B(clk), .A(\g.we_clk [8685]));
Q_ASSIGN U24090 ( .B(clk), .A(\g.we_clk [8684]));
Q_ASSIGN U24091 ( .B(clk), .A(\g.we_clk [8683]));
Q_ASSIGN U24092 ( .B(clk), .A(\g.we_clk [8682]));
Q_ASSIGN U24093 ( .B(clk), .A(\g.we_clk [8681]));
Q_ASSIGN U24094 ( .B(clk), .A(\g.we_clk [8680]));
Q_ASSIGN U24095 ( .B(clk), .A(\g.we_clk [8679]));
Q_ASSIGN U24096 ( .B(clk), .A(\g.we_clk [8678]));
Q_ASSIGN U24097 ( .B(clk), .A(\g.we_clk [8677]));
Q_ASSIGN U24098 ( .B(clk), .A(\g.we_clk [8676]));
Q_ASSIGN U24099 ( .B(clk), .A(\g.we_clk [8675]));
Q_ASSIGN U24100 ( .B(clk), .A(\g.we_clk [8674]));
Q_ASSIGN U24101 ( .B(clk), .A(\g.we_clk [8673]));
Q_ASSIGN U24102 ( .B(clk), .A(\g.we_clk [8672]));
Q_ASSIGN U24103 ( .B(clk), .A(\g.we_clk [8671]));
Q_ASSIGN U24104 ( .B(clk), .A(\g.we_clk [8670]));
Q_ASSIGN U24105 ( .B(clk), .A(\g.we_clk [8669]));
Q_ASSIGN U24106 ( .B(clk), .A(\g.we_clk [8668]));
Q_ASSIGN U24107 ( .B(clk), .A(\g.we_clk [8667]));
Q_ASSIGN U24108 ( .B(clk), .A(\g.we_clk [8666]));
Q_ASSIGN U24109 ( .B(clk), .A(\g.we_clk [8665]));
Q_ASSIGN U24110 ( .B(clk), .A(\g.we_clk [8664]));
Q_ASSIGN U24111 ( .B(clk), .A(\g.we_clk [8663]));
Q_ASSIGN U24112 ( .B(clk), .A(\g.we_clk [8662]));
Q_ASSIGN U24113 ( .B(clk), .A(\g.we_clk [8661]));
Q_ASSIGN U24114 ( .B(clk), .A(\g.we_clk [8660]));
Q_ASSIGN U24115 ( .B(clk), .A(\g.we_clk [8659]));
Q_ASSIGN U24116 ( .B(clk), .A(\g.we_clk [8658]));
Q_ASSIGN U24117 ( .B(clk), .A(\g.we_clk [8657]));
Q_ASSIGN U24118 ( .B(clk), .A(\g.we_clk [8656]));
Q_ASSIGN U24119 ( .B(clk), .A(\g.we_clk [8655]));
Q_ASSIGN U24120 ( .B(clk), .A(\g.we_clk [8654]));
Q_ASSIGN U24121 ( .B(clk), .A(\g.we_clk [8653]));
Q_ASSIGN U24122 ( .B(clk), .A(\g.we_clk [8652]));
Q_ASSIGN U24123 ( .B(clk), .A(\g.we_clk [8651]));
Q_ASSIGN U24124 ( .B(clk), .A(\g.we_clk [8650]));
Q_ASSIGN U24125 ( .B(clk), .A(\g.we_clk [8649]));
Q_ASSIGN U24126 ( .B(clk), .A(\g.we_clk [8648]));
Q_ASSIGN U24127 ( .B(clk), .A(\g.we_clk [8647]));
Q_ASSIGN U24128 ( .B(clk), .A(\g.we_clk [8646]));
Q_ASSIGN U24129 ( .B(clk), .A(\g.we_clk [8645]));
Q_ASSIGN U24130 ( .B(clk), .A(\g.we_clk [8644]));
Q_ASSIGN U24131 ( .B(clk), .A(\g.we_clk [8643]));
Q_ASSIGN U24132 ( .B(clk), .A(\g.we_clk [8642]));
Q_ASSIGN U24133 ( .B(clk), .A(\g.we_clk [8641]));
Q_ASSIGN U24134 ( .B(clk), .A(\g.we_clk [8640]));
Q_ASSIGN U24135 ( .B(clk), .A(\g.we_clk [8639]));
Q_ASSIGN U24136 ( .B(clk), .A(\g.we_clk [8638]));
Q_ASSIGN U24137 ( .B(clk), .A(\g.we_clk [8637]));
Q_ASSIGN U24138 ( .B(clk), .A(\g.we_clk [8636]));
Q_ASSIGN U24139 ( .B(clk), .A(\g.we_clk [8635]));
Q_ASSIGN U24140 ( .B(clk), .A(\g.we_clk [8634]));
Q_ASSIGN U24141 ( .B(clk), .A(\g.we_clk [8633]));
Q_ASSIGN U24142 ( .B(clk), .A(\g.we_clk [8632]));
Q_ASSIGN U24143 ( .B(clk), .A(\g.we_clk [8631]));
Q_ASSIGN U24144 ( .B(clk), .A(\g.we_clk [8630]));
Q_ASSIGN U24145 ( .B(clk), .A(\g.we_clk [8629]));
Q_ASSIGN U24146 ( .B(clk), .A(\g.we_clk [8628]));
Q_ASSIGN U24147 ( .B(clk), .A(\g.we_clk [8627]));
Q_ASSIGN U24148 ( .B(clk), .A(\g.we_clk [8626]));
Q_ASSIGN U24149 ( .B(clk), .A(\g.we_clk [8625]));
Q_ASSIGN U24150 ( .B(clk), .A(\g.we_clk [8624]));
Q_ASSIGN U24151 ( .B(clk), .A(\g.we_clk [8623]));
Q_ASSIGN U24152 ( .B(clk), .A(\g.we_clk [8622]));
Q_ASSIGN U24153 ( .B(clk), .A(\g.we_clk [8621]));
Q_ASSIGN U24154 ( .B(clk), .A(\g.we_clk [8620]));
Q_ASSIGN U24155 ( .B(clk), .A(\g.we_clk [8619]));
Q_ASSIGN U24156 ( .B(clk), .A(\g.we_clk [8618]));
Q_ASSIGN U24157 ( .B(clk), .A(\g.we_clk [8617]));
Q_ASSIGN U24158 ( .B(clk), .A(\g.we_clk [8616]));
Q_ASSIGN U24159 ( .B(clk), .A(\g.we_clk [8615]));
Q_ASSIGN U24160 ( .B(clk), .A(\g.we_clk [8614]));
Q_ASSIGN U24161 ( .B(clk), .A(\g.we_clk [8613]));
Q_ASSIGN U24162 ( .B(clk), .A(\g.we_clk [8612]));
Q_ASSIGN U24163 ( .B(clk), .A(\g.we_clk [8611]));
Q_ASSIGN U24164 ( .B(clk), .A(\g.we_clk [8610]));
Q_ASSIGN U24165 ( .B(clk), .A(\g.we_clk [8609]));
Q_ASSIGN U24166 ( .B(clk), .A(\g.we_clk [8608]));
Q_ASSIGN U24167 ( .B(clk), .A(\g.we_clk [8607]));
Q_ASSIGN U24168 ( .B(clk), .A(\g.we_clk [8606]));
Q_ASSIGN U24169 ( .B(clk), .A(\g.we_clk [8605]));
Q_ASSIGN U24170 ( .B(clk), .A(\g.we_clk [8604]));
Q_ASSIGN U24171 ( .B(clk), .A(\g.we_clk [8603]));
Q_ASSIGN U24172 ( .B(clk), .A(\g.we_clk [8602]));
Q_ASSIGN U24173 ( .B(clk), .A(\g.we_clk [8601]));
Q_ASSIGN U24174 ( .B(clk), .A(\g.we_clk [8600]));
Q_ASSIGN U24175 ( .B(clk), .A(\g.we_clk [8599]));
Q_ASSIGN U24176 ( .B(clk), .A(\g.we_clk [8598]));
Q_ASSIGN U24177 ( .B(clk), .A(\g.we_clk [8597]));
Q_ASSIGN U24178 ( .B(clk), .A(\g.we_clk [8596]));
Q_ASSIGN U24179 ( .B(clk), .A(\g.we_clk [8595]));
Q_ASSIGN U24180 ( .B(clk), .A(\g.we_clk [8594]));
Q_ASSIGN U24181 ( .B(clk), .A(\g.we_clk [8593]));
Q_ASSIGN U24182 ( .B(clk), .A(\g.we_clk [8592]));
Q_ASSIGN U24183 ( .B(clk), .A(\g.we_clk [8591]));
Q_ASSIGN U24184 ( .B(clk), .A(\g.we_clk [8590]));
Q_ASSIGN U24185 ( .B(clk), .A(\g.we_clk [8589]));
Q_ASSIGN U24186 ( .B(clk), .A(\g.we_clk [8588]));
Q_ASSIGN U24187 ( .B(clk), .A(\g.we_clk [8587]));
Q_ASSIGN U24188 ( .B(clk), .A(\g.we_clk [8586]));
Q_ASSIGN U24189 ( .B(clk), .A(\g.we_clk [8585]));
Q_ASSIGN U24190 ( .B(clk), .A(\g.we_clk [8584]));
Q_ASSIGN U24191 ( .B(clk), .A(\g.we_clk [8583]));
Q_ASSIGN U24192 ( .B(clk), .A(\g.we_clk [8582]));
Q_ASSIGN U24193 ( .B(clk), .A(\g.we_clk [8581]));
Q_ASSIGN U24194 ( .B(clk), .A(\g.we_clk [8580]));
Q_ASSIGN U24195 ( .B(clk), .A(\g.we_clk [8579]));
Q_ASSIGN U24196 ( .B(clk), .A(\g.we_clk [8578]));
Q_ASSIGN U24197 ( .B(clk), .A(\g.we_clk [8577]));
Q_ASSIGN U24198 ( .B(clk), .A(\g.we_clk [8576]));
Q_ASSIGN U24199 ( .B(clk), .A(\g.we_clk [8575]));
Q_ASSIGN U24200 ( .B(clk), .A(\g.we_clk [8574]));
Q_ASSIGN U24201 ( .B(clk), .A(\g.we_clk [8573]));
Q_ASSIGN U24202 ( .B(clk), .A(\g.we_clk [8572]));
Q_ASSIGN U24203 ( .B(clk), .A(\g.we_clk [8571]));
Q_ASSIGN U24204 ( .B(clk), .A(\g.we_clk [8570]));
Q_ASSIGN U24205 ( .B(clk), .A(\g.we_clk [8569]));
Q_ASSIGN U24206 ( .B(clk), .A(\g.we_clk [8568]));
Q_ASSIGN U24207 ( .B(clk), .A(\g.we_clk [8567]));
Q_ASSIGN U24208 ( .B(clk), .A(\g.we_clk [8566]));
Q_ASSIGN U24209 ( .B(clk), .A(\g.we_clk [8565]));
Q_ASSIGN U24210 ( .B(clk), .A(\g.we_clk [8564]));
Q_ASSIGN U24211 ( .B(clk), .A(\g.we_clk [8563]));
Q_ASSIGN U24212 ( .B(clk), .A(\g.we_clk [8562]));
Q_ASSIGN U24213 ( .B(clk), .A(\g.we_clk [8561]));
Q_ASSIGN U24214 ( .B(clk), .A(\g.we_clk [8560]));
Q_ASSIGN U24215 ( .B(clk), .A(\g.we_clk [8559]));
Q_ASSIGN U24216 ( .B(clk), .A(\g.we_clk [8558]));
Q_ASSIGN U24217 ( .B(clk), .A(\g.we_clk [8557]));
Q_ASSIGN U24218 ( .B(clk), .A(\g.we_clk [8556]));
Q_ASSIGN U24219 ( .B(clk), .A(\g.we_clk [8555]));
Q_ASSIGN U24220 ( .B(clk), .A(\g.we_clk [8554]));
Q_ASSIGN U24221 ( .B(clk), .A(\g.we_clk [8553]));
Q_ASSIGN U24222 ( .B(clk), .A(\g.we_clk [8552]));
Q_ASSIGN U24223 ( .B(clk), .A(\g.we_clk [8551]));
Q_ASSIGN U24224 ( .B(clk), .A(\g.we_clk [8550]));
Q_ASSIGN U24225 ( .B(clk), .A(\g.we_clk [8549]));
Q_ASSIGN U24226 ( .B(clk), .A(\g.we_clk [8548]));
Q_ASSIGN U24227 ( .B(clk), .A(\g.we_clk [8547]));
Q_ASSIGN U24228 ( .B(clk), .A(\g.we_clk [8546]));
Q_ASSIGN U24229 ( .B(clk), .A(\g.we_clk [8545]));
Q_ASSIGN U24230 ( .B(clk), .A(\g.we_clk [8544]));
Q_ASSIGN U24231 ( .B(clk), .A(\g.we_clk [8543]));
Q_ASSIGN U24232 ( .B(clk), .A(\g.we_clk [8542]));
Q_ASSIGN U24233 ( .B(clk), .A(\g.we_clk [8541]));
Q_ASSIGN U24234 ( .B(clk), .A(\g.we_clk [8540]));
Q_ASSIGN U24235 ( .B(clk), .A(\g.we_clk [8539]));
Q_ASSIGN U24236 ( .B(clk), .A(\g.we_clk [8538]));
Q_ASSIGN U24237 ( .B(clk), .A(\g.we_clk [8537]));
Q_ASSIGN U24238 ( .B(clk), .A(\g.we_clk [8536]));
Q_ASSIGN U24239 ( .B(clk), .A(\g.we_clk [8535]));
Q_ASSIGN U24240 ( .B(clk), .A(\g.we_clk [8534]));
Q_ASSIGN U24241 ( .B(clk), .A(\g.we_clk [8533]));
Q_ASSIGN U24242 ( .B(clk), .A(\g.we_clk [8532]));
Q_ASSIGN U24243 ( .B(clk), .A(\g.we_clk [8531]));
Q_ASSIGN U24244 ( .B(clk), .A(\g.we_clk [8530]));
Q_ASSIGN U24245 ( .B(clk), .A(\g.we_clk [8529]));
Q_ASSIGN U24246 ( .B(clk), .A(\g.we_clk [8528]));
Q_ASSIGN U24247 ( .B(clk), .A(\g.we_clk [8527]));
Q_ASSIGN U24248 ( .B(clk), .A(\g.we_clk [8526]));
Q_ASSIGN U24249 ( .B(clk), .A(\g.we_clk [8525]));
Q_ASSIGN U24250 ( .B(clk), .A(\g.we_clk [8524]));
Q_ASSIGN U24251 ( .B(clk), .A(\g.we_clk [8523]));
Q_ASSIGN U24252 ( .B(clk), .A(\g.we_clk [8522]));
Q_ASSIGN U24253 ( .B(clk), .A(\g.we_clk [8521]));
Q_ASSIGN U24254 ( .B(clk), .A(\g.we_clk [8520]));
Q_ASSIGN U24255 ( .B(clk), .A(\g.we_clk [8519]));
Q_ASSIGN U24256 ( .B(clk), .A(\g.we_clk [8518]));
Q_ASSIGN U24257 ( .B(clk), .A(\g.we_clk [8517]));
Q_ASSIGN U24258 ( .B(clk), .A(\g.we_clk [8516]));
Q_ASSIGN U24259 ( .B(clk), .A(\g.we_clk [8515]));
Q_ASSIGN U24260 ( .B(clk), .A(\g.we_clk [8514]));
Q_ASSIGN U24261 ( .B(clk), .A(\g.we_clk [8513]));
Q_ASSIGN U24262 ( .B(clk), .A(\g.we_clk [8512]));
Q_ASSIGN U24263 ( .B(clk), .A(\g.we_clk [8511]));
Q_ASSIGN U24264 ( .B(clk), .A(\g.we_clk [8510]));
Q_ASSIGN U24265 ( .B(clk), .A(\g.we_clk [8509]));
Q_ASSIGN U24266 ( .B(clk), .A(\g.we_clk [8508]));
Q_ASSIGN U24267 ( .B(clk), .A(\g.we_clk [8507]));
Q_ASSIGN U24268 ( .B(clk), .A(\g.we_clk [8506]));
Q_ASSIGN U24269 ( .B(clk), .A(\g.we_clk [8505]));
Q_ASSIGN U24270 ( .B(clk), .A(\g.we_clk [8504]));
Q_ASSIGN U24271 ( .B(clk), .A(\g.we_clk [8503]));
Q_ASSIGN U24272 ( .B(clk), .A(\g.we_clk [8502]));
Q_ASSIGN U24273 ( .B(clk), .A(\g.we_clk [8501]));
Q_ASSIGN U24274 ( .B(clk), .A(\g.we_clk [8500]));
Q_ASSIGN U24275 ( .B(clk), .A(\g.we_clk [8499]));
Q_ASSIGN U24276 ( .B(clk), .A(\g.we_clk [8498]));
Q_ASSIGN U24277 ( .B(clk), .A(\g.we_clk [8497]));
Q_ASSIGN U24278 ( .B(clk), .A(\g.we_clk [8496]));
Q_ASSIGN U24279 ( .B(clk), .A(\g.we_clk [8495]));
Q_ASSIGN U24280 ( .B(clk), .A(\g.we_clk [8494]));
Q_ASSIGN U24281 ( .B(clk), .A(\g.we_clk [8493]));
Q_ASSIGN U24282 ( .B(clk), .A(\g.we_clk [8492]));
Q_ASSIGN U24283 ( .B(clk), .A(\g.we_clk [8491]));
Q_ASSIGN U24284 ( .B(clk), .A(\g.we_clk [8490]));
Q_ASSIGN U24285 ( .B(clk), .A(\g.we_clk [8489]));
Q_ASSIGN U24286 ( .B(clk), .A(\g.we_clk [8488]));
Q_ASSIGN U24287 ( .B(clk), .A(\g.we_clk [8487]));
Q_ASSIGN U24288 ( .B(clk), .A(\g.we_clk [8486]));
Q_ASSIGN U24289 ( .B(clk), .A(\g.we_clk [8485]));
Q_ASSIGN U24290 ( .B(clk), .A(\g.we_clk [8484]));
Q_ASSIGN U24291 ( .B(clk), .A(\g.we_clk [8483]));
Q_ASSIGN U24292 ( .B(clk), .A(\g.we_clk [8482]));
Q_ASSIGN U24293 ( .B(clk), .A(\g.we_clk [8481]));
Q_ASSIGN U24294 ( .B(clk), .A(\g.we_clk [8480]));
Q_ASSIGN U24295 ( .B(clk), .A(\g.we_clk [8479]));
Q_ASSIGN U24296 ( .B(clk), .A(\g.we_clk [8478]));
Q_ASSIGN U24297 ( .B(clk), .A(\g.we_clk [8477]));
Q_ASSIGN U24298 ( .B(clk), .A(\g.we_clk [8476]));
Q_ASSIGN U24299 ( .B(clk), .A(\g.we_clk [8475]));
Q_ASSIGN U24300 ( .B(clk), .A(\g.we_clk [8474]));
Q_ASSIGN U24301 ( .B(clk), .A(\g.we_clk [8473]));
Q_ASSIGN U24302 ( .B(clk), .A(\g.we_clk [8472]));
Q_ASSIGN U24303 ( .B(clk), .A(\g.we_clk [8471]));
Q_ASSIGN U24304 ( .B(clk), .A(\g.we_clk [8470]));
Q_ASSIGN U24305 ( .B(clk), .A(\g.we_clk [8469]));
Q_ASSIGN U24306 ( .B(clk), .A(\g.we_clk [8468]));
Q_ASSIGN U24307 ( .B(clk), .A(\g.we_clk [8467]));
Q_ASSIGN U24308 ( .B(clk), .A(\g.we_clk [8466]));
Q_ASSIGN U24309 ( .B(clk), .A(\g.we_clk [8465]));
Q_ASSIGN U24310 ( .B(clk), .A(\g.we_clk [8464]));
Q_ASSIGN U24311 ( .B(clk), .A(\g.we_clk [8463]));
Q_ASSIGN U24312 ( .B(clk), .A(\g.we_clk [8462]));
Q_ASSIGN U24313 ( .B(clk), .A(\g.we_clk [8461]));
Q_ASSIGN U24314 ( .B(clk), .A(\g.we_clk [8460]));
Q_ASSIGN U24315 ( .B(clk), .A(\g.we_clk [8459]));
Q_ASSIGN U24316 ( .B(clk), .A(\g.we_clk [8458]));
Q_ASSIGN U24317 ( .B(clk), .A(\g.we_clk [8457]));
Q_ASSIGN U24318 ( .B(clk), .A(\g.we_clk [8456]));
Q_ASSIGN U24319 ( .B(clk), .A(\g.we_clk [8455]));
Q_ASSIGN U24320 ( .B(clk), .A(\g.we_clk [8454]));
Q_ASSIGN U24321 ( .B(clk), .A(\g.we_clk [8453]));
Q_ASSIGN U24322 ( .B(clk), .A(\g.we_clk [8452]));
Q_ASSIGN U24323 ( .B(clk), .A(\g.we_clk [8451]));
Q_ASSIGN U24324 ( .B(clk), .A(\g.we_clk [8450]));
Q_ASSIGN U24325 ( .B(clk), .A(\g.we_clk [8449]));
Q_ASSIGN U24326 ( .B(clk), .A(\g.we_clk [8448]));
Q_ASSIGN U24327 ( .B(clk), .A(\g.we_clk [8447]));
Q_ASSIGN U24328 ( .B(clk), .A(\g.we_clk [8446]));
Q_ASSIGN U24329 ( .B(clk), .A(\g.we_clk [8445]));
Q_ASSIGN U24330 ( .B(clk), .A(\g.we_clk [8444]));
Q_ASSIGN U24331 ( .B(clk), .A(\g.we_clk [8443]));
Q_ASSIGN U24332 ( .B(clk), .A(\g.we_clk [8442]));
Q_ASSIGN U24333 ( .B(clk), .A(\g.we_clk [8441]));
Q_ASSIGN U24334 ( .B(clk), .A(\g.we_clk [8440]));
Q_ASSIGN U24335 ( .B(clk), .A(\g.we_clk [8439]));
Q_ASSIGN U24336 ( .B(clk), .A(\g.we_clk [8438]));
Q_ASSIGN U24337 ( .B(clk), .A(\g.we_clk [8437]));
Q_ASSIGN U24338 ( .B(clk), .A(\g.we_clk [8436]));
Q_ASSIGN U24339 ( .B(clk), .A(\g.we_clk [8435]));
Q_ASSIGN U24340 ( .B(clk), .A(\g.we_clk [8434]));
Q_ASSIGN U24341 ( .B(clk), .A(\g.we_clk [8433]));
Q_ASSIGN U24342 ( .B(clk), .A(\g.we_clk [8432]));
Q_ASSIGN U24343 ( .B(clk), .A(\g.we_clk [8431]));
Q_ASSIGN U24344 ( .B(clk), .A(\g.we_clk [8430]));
Q_ASSIGN U24345 ( .B(clk), .A(\g.we_clk [8429]));
Q_ASSIGN U24346 ( .B(clk), .A(\g.we_clk [8428]));
Q_ASSIGN U24347 ( .B(clk), .A(\g.we_clk [8427]));
Q_ASSIGN U24348 ( .B(clk), .A(\g.we_clk [8426]));
Q_ASSIGN U24349 ( .B(clk), .A(\g.we_clk [8425]));
Q_ASSIGN U24350 ( .B(clk), .A(\g.we_clk [8424]));
Q_ASSIGN U24351 ( .B(clk), .A(\g.we_clk [8423]));
Q_ASSIGN U24352 ( .B(clk), .A(\g.we_clk [8422]));
Q_ASSIGN U24353 ( .B(clk), .A(\g.we_clk [8421]));
Q_ASSIGN U24354 ( .B(clk), .A(\g.we_clk [8420]));
Q_ASSIGN U24355 ( .B(clk), .A(\g.we_clk [8419]));
Q_ASSIGN U24356 ( .B(clk), .A(\g.we_clk [8418]));
Q_ASSIGN U24357 ( .B(clk), .A(\g.we_clk [8417]));
Q_ASSIGN U24358 ( .B(clk), .A(\g.we_clk [8416]));
Q_ASSIGN U24359 ( .B(clk), .A(\g.we_clk [8415]));
Q_ASSIGN U24360 ( .B(clk), .A(\g.we_clk [8414]));
Q_ASSIGN U24361 ( .B(clk), .A(\g.we_clk [8413]));
Q_ASSIGN U24362 ( .B(clk), .A(\g.we_clk [8412]));
Q_ASSIGN U24363 ( .B(clk), .A(\g.we_clk [8411]));
Q_ASSIGN U24364 ( .B(clk), .A(\g.we_clk [8410]));
Q_ASSIGN U24365 ( .B(clk), .A(\g.we_clk [8409]));
Q_ASSIGN U24366 ( .B(clk), .A(\g.we_clk [8408]));
Q_ASSIGN U24367 ( .B(clk), .A(\g.we_clk [8407]));
Q_ASSIGN U24368 ( .B(clk), .A(\g.we_clk [8406]));
Q_ASSIGN U24369 ( .B(clk), .A(\g.we_clk [8405]));
Q_ASSIGN U24370 ( .B(clk), .A(\g.we_clk [8404]));
Q_ASSIGN U24371 ( .B(clk), .A(\g.we_clk [8403]));
Q_ASSIGN U24372 ( .B(clk), .A(\g.we_clk [8402]));
Q_ASSIGN U24373 ( .B(clk), .A(\g.we_clk [8401]));
Q_ASSIGN U24374 ( .B(clk), .A(\g.we_clk [8400]));
Q_ASSIGN U24375 ( .B(clk), .A(\g.we_clk [8399]));
Q_ASSIGN U24376 ( .B(clk), .A(\g.we_clk [8398]));
Q_ASSIGN U24377 ( .B(clk), .A(\g.we_clk [8397]));
Q_ASSIGN U24378 ( .B(clk), .A(\g.we_clk [8396]));
Q_ASSIGN U24379 ( .B(clk), .A(\g.we_clk [8395]));
Q_ASSIGN U24380 ( .B(clk), .A(\g.we_clk [8394]));
Q_ASSIGN U24381 ( .B(clk), .A(\g.we_clk [8393]));
Q_ASSIGN U24382 ( .B(clk), .A(\g.we_clk [8392]));
Q_ASSIGN U24383 ( .B(clk), .A(\g.we_clk [8391]));
Q_ASSIGN U24384 ( .B(clk), .A(\g.we_clk [8390]));
Q_ASSIGN U24385 ( .B(clk), .A(\g.we_clk [8389]));
Q_ASSIGN U24386 ( .B(clk), .A(\g.we_clk [8388]));
Q_ASSIGN U24387 ( .B(clk), .A(\g.we_clk [8387]));
Q_ASSIGN U24388 ( .B(clk), .A(\g.we_clk [8386]));
Q_ASSIGN U24389 ( .B(clk), .A(\g.we_clk [8385]));
Q_ASSIGN U24390 ( .B(clk), .A(\g.we_clk [8384]));
Q_ASSIGN U24391 ( .B(clk), .A(\g.we_clk [8383]));
Q_ASSIGN U24392 ( .B(clk), .A(\g.we_clk [8382]));
Q_ASSIGN U24393 ( .B(clk), .A(\g.we_clk [8381]));
Q_ASSIGN U24394 ( .B(clk), .A(\g.we_clk [8380]));
Q_ASSIGN U24395 ( .B(clk), .A(\g.we_clk [8379]));
Q_ASSIGN U24396 ( .B(clk), .A(\g.we_clk [8378]));
Q_ASSIGN U24397 ( .B(clk), .A(\g.we_clk [8377]));
Q_ASSIGN U24398 ( .B(clk), .A(\g.we_clk [8376]));
Q_ASSIGN U24399 ( .B(clk), .A(\g.we_clk [8375]));
Q_ASSIGN U24400 ( .B(clk), .A(\g.we_clk [8374]));
Q_ASSIGN U24401 ( .B(clk), .A(\g.we_clk [8373]));
Q_ASSIGN U24402 ( .B(clk), .A(\g.we_clk [8372]));
Q_ASSIGN U24403 ( .B(clk), .A(\g.we_clk [8371]));
Q_ASSIGN U24404 ( .B(clk), .A(\g.we_clk [8370]));
Q_ASSIGN U24405 ( .B(clk), .A(\g.we_clk [8369]));
Q_ASSIGN U24406 ( .B(clk), .A(\g.we_clk [8368]));
Q_ASSIGN U24407 ( .B(clk), .A(\g.we_clk [8367]));
Q_ASSIGN U24408 ( .B(clk), .A(\g.we_clk [8366]));
Q_ASSIGN U24409 ( .B(clk), .A(\g.we_clk [8365]));
Q_ASSIGN U24410 ( .B(clk), .A(\g.we_clk [8364]));
Q_ASSIGN U24411 ( .B(clk), .A(\g.we_clk [8363]));
Q_ASSIGN U24412 ( .B(clk), .A(\g.we_clk [8362]));
Q_ASSIGN U24413 ( .B(clk), .A(\g.we_clk [8361]));
Q_ASSIGN U24414 ( .B(clk), .A(\g.we_clk [8360]));
Q_ASSIGN U24415 ( .B(clk), .A(\g.we_clk [8359]));
Q_ASSIGN U24416 ( .B(clk), .A(\g.we_clk [8358]));
Q_ASSIGN U24417 ( .B(clk), .A(\g.we_clk [8357]));
Q_ASSIGN U24418 ( .B(clk), .A(\g.we_clk [8356]));
Q_ASSIGN U24419 ( .B(clk), .A(\g.we_clk [8355]));
Q_ASSIGN U24420 ( .B(clk), .A(\g.we_clk [8354]));
Q_ASSIGN U24421 ( .B(clk), .A(\g.we_clk [8353]));
Q_ASSIGN U24422 ( .B(clk), .A(\g.we_clk [8352]));
Q_ASSIGN U24423 ( .B(clk), .A(\g.we_clk [8351]));
Q_ASSIGN U24424 ( .B(clk), .A(\g.we_clk [8350]));
Q_ASSIGN U24425 ( .B(clk), .A(\g.we_clk [8349]));
Q_ASSIGN U24426 ( .B(clk), .A(\g.we_clk [8348]));
Q_ASSIGN U24427 ( .B(clk), .A(\g.we_clk [8347]));
Q_ASSIGN U24428 ( .B(clk), .A(\g.we_clk [8346]));
Q_ASSIGN U24429 ( .B(clk), .A(\g.we_clk [8345]));
Q_ASSIGN U24430 ( .B(clk), .A(\g.we_clk [8344]));
Q_ASSIGN U24431 ( .B(clk), .A(\g.we_clk [8343]));
Q_ASSIGN U24432 ( .B(clk), .A(\g.we_clk [8342]));
Q_ASSIGN U24433 ( .B(clk), .A(\g.we_clk [8341]));
Q_ASSIGN U24434 ( .B(clk), .A(\g.we_clk [8340]));
Q_ASSIGN U24435 ( .B(clk), .A(\g.we_clk [8339]));
Q_ASSIGN U24436 ( .B(clk), .A(\g.we_clk [8338]));
Q_ASSIGN U24437 ( .B(clk), .A(\g.we_clk [8337]));
Q_ASSIGN U24438 ( .B(clk), .A(\g.we_clk [8336]));
Q_ASSIGN U24439 ( .B(clk), .A(\g.we_clk [8335]));
Q_ASSIGN U24440 ( .B(clk), .A(\g.we_clk [8334]));
Q_ASSIGN U24441 ( .B(clk), .A(\g.we_clk [8333]));
Q_ASSIGN U24442 ( .B(clk), .A(\g.we_clk [8332]));
Q_ASSIGN U24443 ( .B(clk), .A(\g.we_clk [8331]));
Q_ASSIGN U24444 ( .B(clk), .A(\g.we_clk [8330]));
Q_ASSIGN U24445 ( .B(clk), .A(\g.we_clk [8329]));
Q_ASSIGN U24446 ( .B(clk), .A(\g.we_clk [8328]));
Q_ASSIGN U24447 ( .B(clk), .A(\g.we_clk [8327]));
Q_ASSIGN U24448 ( .B(clk), .A(\g.we_clk [8326]));
Q_ASSIGN U24449 ( .B(clk), .A(\g.we_clk [8325]));
Q_ASSIGN U24450 ( .B(clk), .A(\g.we_clk [8324]));
Q_ASSIGN U24451 ( .B(clk), .A(\g.we_clk [8323]));
Q_ASSIGN U24452 ( .B(clk), .A(\g.we_clk [8322]));
Q_ASSIGN U24453 ( .B(clk), .A(\g.we_clk [8321]));
Q_ASSIGN U24454 ( .B(clk), .A(\g.we_clk [8320]));
Q_ASSIGN U24455 ( .B(clk), .A(\g.we_clk [8319]));
Q_ASSIGN U24456 ( .B(clk), .A(\g.we_clk [8318]));
Q_ASSIGN U24457 ( .B(clk), .A(\g.we_clk [8317]));
Q_ASSIGN U24458 ( .B(clk), .A(\g.we_clk [8316]));
Q_ASSIGN U24459 ( .B(clk), .A(\g.we_clk [8315]));
Q_ASSIGN U24460 ( .B(clk), .A(\g.we_clk [8314]));
Q_ASSIGN U24461 ( .B(clk), .A(\g.we_clk [8313]));
Q_ASSIGN U24462 ( .B(clk), .A(\g.we_clk [8312]));
Q_ASSIGN U24463 ( .B(clk), .A(\g.we_clk [8311]));
Q_ASSIGN U24464 ( .B(clk), .A(\g.we_clk [8310]));
Q_ASSIGN U24465 ( .B(clk), .A(\g.we_clk [8309]));
Q_ASSIGN U24466 ( .B(clk), .A(\g.we_clk [8308]));
Q_ASSIGN U24467 ( .B(clk), .A(\g.we_clk [8307]));
Q_ASSIGN U24468 ( .B(clk), .A(\g.we_clk [8306]));
Q_ASSIGN U24469 ( .B(clk), .A(\g.we_clk [8305]));
Q_ASSIGN U24470 ( .B(clk), .A(\g.we_clk [8304]));
Q_ASSIGN U24471 ( .B(clk), .A(\g.we_clk [8303]));
Q_ASSIGN U24472 ( .B(clk), .A(\g.we_clk [8302]));
Q_ASSIGN U24473 ( .B(clk), .A(\g.we_clk [8301]));
Q_ASSIGN U24474 ( .B(clk), .A(\g.we_clk [8300]));
Q_ASSIGN U24475 ( .B(clk), .A(\g.we_clk [8299]));
Q_ASSIGN U24476 ( .B(clk), .A(\g.we_clk [8298]));
Q_ASSIGN U24477 ( .B(clk), .A(\g.we_clk [8297]));
Q_ASSIGN U24478 ( .B(clk), .A(\g.we_clk [8296]));
Q_ASSIGN U24479 ( .B(clk), .A(\g.we_clk [8295]));
Q_ASSIGN U24480 ( .B(clk), .A(\g.we_clk [8294]));
Q_ASSIGN U24481 ( .B(clk), .A(\g.we_clk [8293]));
Q_ASSIGN U24482 ( .B(clk), .A(\g.we_clk [8292]));
Q_ASSIGN U24483 ( .B(clk), .A(\g.we_clk [8291]));
Q_ASSIGN U24484 ( .B(clk), .A(\g.we_clk [8290]));
Q_ASSIGN U24485 ( .B(clk), .A(\g.we_clk [8289]));
Q_ASSIGN U24486 ( .B(clk), .A(\g.we_clk [8288]));
Q_ASSIGN U24487 ( .B(clk), .A(\g.we_clk [8287]));
Q_ASSIGN U24488 ( .B(clk), .A(\g.we_clk [8286]));
Q_ASSIGN U24489 ( .B(clk), .A(\g.we_clk [8285]));
Q_ASSIGN U24490 ( .B(clk), .A(\g.we_clk [8284]));
Q_ASSIGN U24491 ( .B(clk), .A(\g.we_clk [8283]));
Q_ASSIGN U24492 ( .B(clk), .A(\g.we_clk [8282]));
Q_ASSIGN U24493 ( .B(clk), .A(\g.we_clk [8281]));
Q_ASSIGN U24494 ( .B(clk), .A(\g.we_clk [8280]));
Q_ASSIGN U24495 ( .B(clk), .A(\g.we_clk [8279]));
Q_ASSIGN U24496 ( .B(clk), .A(\g.we_clk [8278]));
Q_ASSIGN U24497 ( .B(clk), .A(\g.we_clk [8277]));
Q_ASSIGN U24498 ( .B(clk), .A(\g.we_clk [8276]));
Q_ASSIGN U24499 ( .B(clk), .A(\g.we_clk [8275]));
Q_ASSIGN U24500 ( .B(clk), .A(\g.we_clk [8274]));
Q_ASSIGN U24501 ( .B(clk), .A(\g.we_clk [8273]));
Q_ASSIGN U24502 ( .B(clk), .A(\g.we_clk [8272]));
Q_ASSIGN U24503 ( .B(clk), .A(\g.we_clk [8271]));
Q_ASSIGN U24504 ( .B(clk), .A(\g.we_clk [8270]));
Q_ASSIGN U24505 ( .B(clk), .A(\g.we_clk [8269]));
Q_ASSIGN U24506 ( .B(clk), .A(\g.we_clk [8268]));
Q_ASSIGN U24507 ( .B(clk), .A(\g.we_clk [8267]));
Q_ASSIGN U24508 ( .B(clk), .A(\g.we_clk [8266]));
Q_ASSIGN U24509 ( .B(clk), .A(\g.we_clk [8265]));
Q_ASSIGN U24510 ( .B(clk), .A(\g.we_clk [8264]));
Q_ASSIGN U24511 ( .B(clk), .A(\g.we_clk [8263]));
Q_ASSIGN U24512 ( .B(clk), .A(\g.we_clk [8262]));
Q_ASSIGN U24513 ( .B(clk), .A(\g.we_clk [8261]));
Q_ASSIGN U24514 ( .B(clk), .A(\g.we_clk [8260]));
Q_ASSIGN U24515 ( .B(clk), .A(\g.we_clk [8259]));
Q_ASSIGN U24516 ( .B(clk), .A(\g.we_clk [8258]));
Q_ASSIGN U24517 ( .B(clk), .A(\g.we_clk [8257]));
Q_ASSIGN U24518 ( .B(clk), .A(\g.we_clk [8256]));
Q_ASSIGN U24519 ( .B(clk), .A(\g.we_clk [8255]));
Q_ASSIGN U24520 ( .B(clk), .A(\g.we_clk [8254]));
Q_ASSIGN U24521 ( .B(clk), .A(\g.we_clk [8253]));
Q_ASSIGN U24522 ( .B(clk), .A(\g.we_clk [8252]));
Q_ASSIGN U24523 ( .B(clk), .A(\g.we_clk [8251]));
Q_ASSIGN U24524 ( .B(clk), .A(\g.we_clk [8250]));
Q_ASSIGN U24525 ( .B(clk), .A(\g.we_clk [8249]));
Q_ASSIGN U24526 ( .B(clk), .A(\g.we_clk [8248]));
Q_ASSIGN U24527 ( .B(clk), .A(\g.we_clk [8247]));
Q_ASSIGN U24528 ( .B(clk), .A(\g.we_clk [8246]));
Q_ASSIGN U24529 ( .B(clk), .A(\g.we_clk [8245]));
Q_ASSIGN U24530 ( .B(clk), .A(\g.we_clk [8244]));
Q_ASSIGN U24531 ( .B(clk), .A(\g.we_clk [8243]));
Q_ASSIGN U24532 ( .B(clk), .A(\g.we_clk [8242]));
Q_ASSIGN U24533 ( .B(clk), .A(\g.we_clk [8241]));
Q_ASSIGN U24534 ( .B(clk), .A(\g.we_clk [8240]));
Q_ASSIGN U24535 ( .B(clk), .A(\g.we_clk [8239]));
Q_ASSIGN U24536 ( .B(clk), .A(\g.we_clk [8238]));
Q_ASSIGN U24537 ( .B(clk), .A(\g.we_clk [8237]));
Q_ASSIGN U24538 ( .B(clk), .A(\g.we_clk [8236]));
Q_ASSIGN U24539 ( .B(clk), .A(\g.we_clk [8235]));
Q_ASSIGN U24540 ( .B(clk), .A(\g.we_clk [8234]));
Q_ASSIGN U24541 ( .B(clk), .A(\g.we_clk [8233]));
Q_ASSIGN U24542 ( .B(clk), .A(\g.we_clk [8232]));
Q_ASSIGN U24543 ( .B(clk), .A(\g.we_clk [8231]));
Q_ASSIGN U24544 ( .B(clk), .A(\g.we_clk [8230]));
Q_ASSIGN U24545 ( .B(clk), .A(\g.we_clk [8229]));
Q_ASSIGN U24546 ( .B(clk), .A(\g.we_clk [8228]));
Q_ASSIGN U24547 ( .B(clk), .A(\g.we_clk [8227]));
Q_ASSIGN U24548 ( .B(clk), .A(\g.we_clk [8226]));
Q_ASSIGN U24549 ( .B(clk), .A(\g.we_clk [8225]));
Q_ASSIGN U24550 ( .B(clk), .A(\g.we_clk [8224]));
Q_ASSIGN U24551 ( .B(clk), .A(\g.we_clk [8223]));
Q_ASSIGN U24552 ( .B(clk), .A(\g.we_clk [8222]));
Q_ASSIGN U24553 ( .B(clk), .A(\g.we_clk [8221]));
Q_ASSIGN U24554 ( .B(clk), .A(\g.we_clk [8220]));
Q_ASSIGN U24555 ( .B(clk), .A(\g.we_clk [8219]));
Q_ASSIGN U24556 ( .B(clk), .A(\g.we_clk [8218]));
Q_ASSIGN U24557 ( .B(clk), .A(\g.we_clk [8217]));
Q_ASSIGN U24558 ( .B(clk), .A(\g.we_clk [8216]));
Q_ASSIGN U24559 ( .B(clk), .A(\g.we_clk [8215]));
Q_ASSIGN U24560 ( .B(clk), .A(\g.we_clk [8214]));
Q_ASSIGN U24561 ( .B(clk), .A(\g.we_clk [8213]));
Q_ASSIGN U24562 ( .B(clk), .A(\g.we_clk [8212]));
Q_ASSIGN U24563 ( .B(clk), .A(\g.we_clk [8211]));
Q_ASSIGN U24564 ( .B(clk), .A(\g.we_clk [8210]));
Q_ASSIGN U24565 ( .B(clk), .A(\g.we_clk [8209]));
Q_ASSIGN U24566 ( .B(clk), .A(\g.we_clk [8208]));
Q_ASSIGN U24567 ( .B(clk), .A(\g.we_clk [8207]));
Q_ASSIGN U24568 ( .B(clk), .A(\g.we_clk [8206]));
Q_ASSIGN U24569 ( .B(clk), .A(\g.we_clk [8205]));
Q_ASSIGN U24570 ( .B(clk), .A(\g.we_clk [8204]));
Q_ASSIGN U24571 ( .B(clk), .A(\g.we_clk [8203]));
Q_ASSIGN U24572 ( .B(clk), .A(\g.we_clk [8202]));
Q_ASSIGN U24573 ( .B(clk), .A(\g.we_clk [8201]));
Q_ASSIGN U24574 ( .B(clk), .A(\g.we_clk [8200]));
Q_ASSIGN U24575 ( .B(clk), .A(\g.we_clk [8199]));
Q_ASSIGN U24576 ( .B(clk), .A(\g.we_clk [8198]));
Q_ASSIGN U24577 ( .B(clk), .A(\g.we_clk [8197]));
Q_ASSIGN U24578 ( .B(clk), .A(\g.we_clk [8196]));
Q_ASSIGN U24579 ( .B(clk), .A(\g.we_clk [8195]));
Q_ASSIGN U24580 ( .B(clk), .A(\g.we_clk [8194]));
Q_ASSIGN U24581 ( .B(clk), .A(\g.we_clk [8193]));
Q_ASSIGN U24582 ( .B(clk), .A(\g.we_clk [8192]));
Q_ASSIGN U24583 ( .B(clk), .A(\g.we_clk [8191]));
Q_ASSIGN U24584 ( .B(clk), .A(\g.we_clk [8190]));
Q_ASSIGN U24585 ( .B(clk), .A(\g.we_clk [8189]));
Q_ASSIGN U24586 ( .B(clk), .A(\g.we_clk [8188]));
Q_ASSIGN U24587 ( .B(clk), .A(\g.we_clk [8187]));
Q_ASSIGN U24588 ( .B(clk), .A(\g.we_clk [8186]));
Q_ASSIGN U24589 ( .B(clk), .A(\g.we_clk [8185]));
Q_ASSIGN U24590 ( .B(clk), .A(\g.we_clk [8184]));
Q_ASSIGN U24591 ( .B(clk), .A(\g.we_clk [8183]));
Q_ASSIGN U24592 ( .B(clk), .A(\g.we_clk [8182]));
Q_ASSIGN U24593 ( .B(clk), .A(\g.we_clk [8181]));
Q_ASSIGN U24594 ( .B(clk), .A(\g.we_clk [8180]));
Q_ASSIGN U24595 ( .B(clk), .A(\g.we_clk [8179]));
Q_ASSIGN U24596 ( .B(clk), .A(\g.we_clk [8178]));
Q_ASSIGN U24597 ( .B(clk), .A(\g.we_clk [8177]));
Q_ASSIGN U24598 ( .B(clk), .A(\g.we_clk [8176]));
Q_ASSIGN U24599 ( .B(clk), .A(\g.we_clk [8175]));
Q_ASSIGN U24600 ( .B(clk), .A(\g.we_clk [8174]));
Q_ASSIGN U24601 ( .B(clk), .A(\g.we_clk [8173]));
Q_ASSIGN U24602 ( .B(clk), .A(\g.we_clk [8172]));
Q_ASSIGN U24603 ( .B(clk), .A(\g.we_clk [8171]));
Q_ASSIGN U24604 ( .B(clk), .A(\g.we_clk [8170]));
Q_ASSIGN U24605 ( .B(clk), .A(\g.we_clk [8169]));
Q_ASSIGN U24606 ( .B(clk), .A(\g.we_clk [8168]));
Q_ASSIGN U24607 ( .B(clk), .A(\g.we_clk [8167]));
Q_ASSIGN U24608 ( .B(clk), .A(\g.we_clk [8166]));
Q_ASSIGN U24609 ( .B(clk), .A(\g.we_clk [8165]));
Q_ASSIGN U24610 ( .B(clk), .A(\g.we_clk [8164]));
Q_ASSIGN U24611 ( .B(clk), .A(\g.we_clk [8163]));
Q_ASSIGN U24612 ( .B(clk), .A(\g.we_clk [8162]));
Q_ASSIGN U24613 ( .B(clk), .A(\g.we_clk [8161]));
Q_ASSIGN U24614 ( .B(clk), .A(\g.we_clk [8160]));
Q_ASSIGN U24615 ( .B(clk), .A(\g.we_clk [8159]));
Q_ASSIGN U24616 ( .B(clk), .A(\g.we_clk [8158]));
Q_ASSIGN U24617 ( .B(clk), .A(\g.we_clk [8157]));
Q_ASSIGN U24618 ( .B(clk), .A(\g.we_clk [8156]));
Q_ASSIGN U24619 ( .B(clk), .A(\g.we_clk [8155]));
Q_ASSIGN U24620 ( .B(clk), .A(\g.we_clk [8154]));
Q_ASSIGN U24621 ( .B(clk), .A(\g.we_clk [8153]));
Q_ASSIGN U24622 ( .B(clk), .A(\g.we_clk [8152]));
Q_ASSIGN U24623 ( .B(clk), .A(\g.we_clk [8151]));
Q_ASSIGN U24624 ( .B(clk), .A(\g.we_clk [8150]));
Q_ASSIGN U24625 ( .B(clk), .A(\g.we_clk [8149]));
Q_ASSIGN U24626 ( .B(clk), .A(\g.we_clk [8148]));
Q_ASSIGN U24627 ( .B(clk), .A(\g.we_clk [8147]));
Q_ASSIGN U24628 ( .B(clk), .A(\g.we_clk [8146]));
Q_ASSIGN U24629 ( .B(clk), .A(\g.we_clk [8145]));
Q_ASSIGN U24630 ( .B(clk), .A(\g.we_clk [8144]));
Q_ASSIGN U24631 ( .B(clk), .A(\g.we_clk [8143]));
Q_ASSIGN U24632 ( .B(clk), .A(\g.we_clk [8142]));
Q_ASSIGN U24633 ( .B(clk), .A(\g.we_clk [8141]));
Q_ASSIGN U24634 ( .B(clk), .A(\g.we_clk [8140]));
Q_ASSIGN U24635 ( .B(clk), .A(\g.we_clk [8139]));
Q_ASSIGN U24636 ( .B(clk), .A(\g.we_clk [8138]));
Q_ASSIGN U24637 ( .B(clk), .A(\g.we_clk [8137]));
Q_ASSIGN U24638 ( .B(clk), .A(\g.we_clk [8136]));
Q_ASSIGN U24639 ( .B(clk), .A(\g.we_clk [8135]));
Q_ASSIGN U24640 ( .B(clk), .A(\g.we_clk [8134]));
Q_ASSIGN U24641 ( .B(clk), .A(\g.we_clk [8133]));
Q_ASSIGN U24642 ( .B(clk), .A(\g.we_clk [8132]));
Q_ASSIGN U24643 ( .B(clk), .A(\g.we_clk [8131]));
Q_ASSIGN U24644 ( .B(clk), .A(\g.we_clk [8130]));
Q_ASSIGN U24645 ( .B(clk), .A(\g.we_clk [8129]));
Q_ASSIGN U24646 ( .B(clk), .A(\g.we_clk [8128]));
Q_ASSIGN U24647 ( .B(clk), .A(\g.we_clk [8127]));
Q_ASSIGN U24648 ( .B(clk), .A(\g.we_clk [8126]));
Q_ASSIGN U24649 ( .B(clk), .A(\g.we_clk [8125]));
Q_ASSIGN U24650 ( .B(clk), .A(\g.we_clk [8124]));
Q_ASSIGN U24651 ( .B(clk), .A(\g.we_clk [8123]));
Q_ASSIGN U24652 ( .B(clk), .A(\g.we_clk [8122]));
Q_ASSIGN U24653 ( .B(clk), .A(\g.we_clk [8121]));
Q_ASSIGN U24654 ( .B(clk), .A(\g.we_clk [8120]));
Q_ASSIGN U24655 ( .B(clk), .A(\g.we_clk [8119]));
Q_ASSIGN U24656 ( .B(clk), .A(\g.we_clk [8118]));
Q_ASSIGN U24657 ( .B(clk), .A(\g.we_clk [8117]));
Q_ASSIGN U24658 ( .B(clk), .A(\g.we_clk [8116]));
Q_ASSIGN U24659 ( .B(clk), .A(\g.we_clk [8115]));
Q_ASSIGN U24660 ( .B(clk), .A(\g.we_clk [8114]));
Q_ASSIGN U24661 ( .B(clk), .A(\g.we_clk [8113]));
Q_ASSIGN U24662 ( .B(clk), .A(\g.we_clk [8112]));
Q_ASSIGN U24663 ( .B(clk), .A(\g.we_clk [8111]));
Q_ASSIGN U24664 ( .B(clk), .A(\g.we_clk [8110]));
Q_ASSIGN U24665 ( .B(clk), .A(\g.we_clk [8109]));
Q_ASSIGN U24666 ( .B(clk), .A(\g.we_clk [8108]));
Q_ASSIGN U24667 ( .B(clk), .A(\g.we_clk [8107]));
Q_ASSIGN U24668 ( .B(clk), .A(\g.we_clk [8106]));
Q_ASSIGN U24669 ( .B(clk), .A(\g.we_clk [8105]));
Q_ASSIGN U24670 ( .B(clk), .A(\g.we_clk [8104]));
Q_ASSIGN U24671 ( .B(clk), .A(\g.we_clk [8103]));
Q_ASSIGN U24672 ( .B(clk), .A(\g.we_clk [8102]));
Q_ASSIGN U24673 ( .B(clk), .A(\g.we_clk [8101]));
Q_ASSIGN U24674 ( .B(clk), .A(\g.we_clk [8100]));
Q_ASSIGN U24675 ( .B(clk), .A(\g.we_clk [8099]));
Q_ASSIGN U24676 ( .B(clk), .A(\g.we_clk [8098]));
Q_ASSIGN U24677 ( .B(clk), .A(\g.we_clk [8097]));
Q_ASSIGN U24678 ( .B(clk), .A(\g.we_clk [8096]));
Q_ASSIGN U24679 ( .B(clk), .A(\g.we_clk [8095]));
Q_ASSIGN U24680 ( .B(clk), .A(\g.we_clk [8094]));
Q_ASSIGN U24681 ( .B(clk), .A(\g.we_clk [8093]));
Q_ASSIGN U24682 ( .B(clk), .A(\g.we_clk [8092]));
Q_ASSIGN U24683 ( .B(clk), .A(\g.we_clk [8091]));
Q_ASSIGN U24684 ( .B(clk), .A(\g.we_clk [8090]));
Q_ASSIGN U24685 ( .B(clk), .A(\g.we_clk [8089]));
Q_ASSIGN U24686 ( .B(clk), .A(\g.we_clk [8088]));
Q_ASSIGN U24687 ( .B(clk), .A(\g.we_clk [8087]));
Q_ASSIGN U24688 ( .B(clk), .A(\g.we_clk [8086]));
Q_ASSIGN U24689 ( .B(clk), .A(\g.we_clk [8085]));
Q_ASSIGN U24690 ( .B(clk), .A(\g.we_clk [8084]));
Q_ASSIGN U24691 ( .B(clk), .A(\g.we_clk [8083]));
Q_ASSIGN U24692 ( .B(clk), .A(\g.we_clk [8082]));
Q_ASSIGN U24693 ( .B(clk), .A(\g.we_clk [8081]));
Q_ASSIGN U24694 ( .B(clk), .A(\g.we_clk [8080]));
Q_ASSIGN U24695 ( .B(clk), .A(\g.we_clk [8079]));
Q_ASSIGN U24696 ( .B(clk), .A(\g.we_clk [8078]));
Q_ASSIGN U24697 ( .B(clk), .A(\g.we_clk [8077]));
Q_ASSIGN U24698 ( .B(clk), .A(\g.we_clk [8076]));
Q_ASSIGN U24699 ( .B(clk), .A(\g.we_clk [8075]));
Q_ASSIGN U24700 ( .B(clk), .A(\g.we_clk [8074]));
Q_ASSIGN U24701 ( .B(clk), .A(\g.we_clk [8073]));
Q_ASSIGN U24702 ( .B(clk), .A(\g.we_clk [8072]));
Q_ASSIGN U24703 ( .B(clk), .A(\g.we_clk [8071]));
Q_ASSIGN U24704 ( .B(clk), .A(\g.we_clk [8070]));
Q_ASSIGN U24705 ( .B(clk), .A(\g.we_clk [8069]));
Q_ASSIGN U24706 ( .B(clk), .A(\g.we_clk [8068]));
Q_ASSIGN U24707 ( .B(clk), .A(\g.we_clk [8067]));
Q_ASSIGN U24708 ( .B(clk), .A(\g.we_clk [8066]));
Q_ASSIGN U24709 ( .B(clk), .A(\g.we_clk [8065]));
Q_ASSIGN U24710 ( .B(clk), .A(\g.we_clk [8064]));
Q_ASSIGN U24711 ( .B(clk), .A(\g.we_clk [8063]));
Q_ASSIGN U24712 ( .B(clk), .A(\g.we_clk [8062]));
Q_ASSIGN U24713 ( .B(clk), .A(\g.we_clk [8061]));
Q_ASSIGN U24714 ( .B(clk), .A(\g.we_clk [8060]));
Q_ASSIGN U24715 ( .B(clk), .A(\g.we_clk [8059]));
Q_ASSIGN U24716 ( .B(clk), .A(\g.we_clk [8058]));
Q_ASSIGN U24717 ( .B(clk), .A(\g.we_clk [8057]));
Q_ASSIGN U24718 ( .B(clk), .A(\g.we_clk [8056]));
Q_ASSIGN U24719 ( .B(clk), .A(\g.we_clk [8055]));
Q_ASSIGN U24720 ( .B(clk), .A(\g.we_clk [8054]));
Q_ASSIGN U24721 ( .B(clk), .A(\g.we_clk [8053]));
Q_ASSIGN U24722 ( .B(clk), .A(\g.we_clk [8052]));
Q_ASSIGN U24723 ( .B(clk), .A(\g.we_clk [8051]));
Q_ASSIGN U24724 ( .B(clk), .A(\g.we_clk [8050]));
Q_ASSIGN U24725 ( .B(clk), .A(\g.we_clk [8049]));
Q_ASSIGN U24726 ( .B(clk), .A(\g.we_clk [8048]));
Q_ASSIGN U24727 ( .B(clk), .A(\g.we_clk [8047]));
Q_ASSIGN U24728 ( .B(clk), .A(\g.we_clk [8046]));
Q_ASSIGN U24729 ( .B(clk), .A(\g.we_clk [8045]));
Q_ASSIGN U24730 ( .B(clk), .A(\g.we_clk [8044]));
Q_ASSIGN U24731 ( .B(clk), .A(\g.we_clk [8043]));
Q_ASSIGN U24732 ( .B(clk), .A(\g.we_clk [8042]));
Q_ASSIGN U24733 ( .B(clk), .A(\g.we_clk [8041]));
Q_ASSIGN U24734 ( .B(clk), .A(\g.we_clk [8040]));
Q_ASSIGN U24735 ( .B(clk), .A(\g.we_clk [8039]));
Q_ASSIGN U24736 ( .B(clk), .A(\g.we_clk [8038]));
Q_ASSIGN U24737 ( .B(clk), .A(\g.we_clk [8037]));
Q_ASSIGN U24738 ( .B(clk), .A(\g.we_clk [8036]));
Q_ASSIGN U24739 ( .B(clk), .A(\g.we_clk [8035]));
Q_ASSIGN U24740 ( .B(clk), .A(\g.we_clk [8034]));
Q_ASSIGN U24741 ( .B(clk), .A(\g.we_clk [8033]));
Q_ASSIGN U24742 ( .B(clk), .A(\g.we_clk [8032]));
Q_ASSIGN U24743 ( .B(clk), .A(\g.we_clk [8031]));
Q_ASSIGN U24744 ( .B(clk), .A(\g.we_clk [8030]));
Q_ASSIGN U24745 ( .B(clk), .A(\g.we_clk [8029]));
Q_ASSIGN U24746 ( .B(clk), .A(\g.we_clk [8028]));
Q_ASSIGN U24747 ( .B(clk), .A(\g.we_clk [8027]));
Q_ASSIGN U24748 ( .B(clk), .A(\g.we_clk [8026]));
Q_ASSIGN U24749 ( .B(clk), .A(\g.we_clk [8025]));
Q_ASSIGN U24750 ( .B(clk), .A(\g.we_clk [8024]));
Q_ASSIGN U24751 ( .B(clk), .A(\g.we_clk [8023]));
Q_ASSIGN U24752 ( .B(clk), .A(\g.we_clk [8022]));
Q_ASSIGN U24753 ( .B(clk), .A(\g.we_clk [8021]));
Q_ASSIGN U24754 ( .B(clk), .A(\g.we_clk [8020]));
Q_ASSIGN U24755 ( .B(clk), .A(\g.we_clk [8019]));
Q_ASSIGN U24756 ( .B(clk), .A(\g.we_clk [8018]));
Q_ASSIGN U24757 ( .B(clk), .A(\g.we_clk [8017]));
Q_ASSIGN U24758 ( .B(clk), .A(\g.we_clk [8016]));
Q_ASSIGN U24759 ( .B(clk), .A(\g.we_clk [8015]));
Q_ASSIGN U24760 ( .B(clk), .A(\g.we_clk [8014]));
Q_ASSIGN U24761 ( .B(clk), .A(\g.we_clk [8013]));
Q_ASSIGN U24762 ( .B(clk), .A(\g.we_clk [8012]));
Q_ASSIGN U24763 ( .B(clk), .A(\g.we_clk [8011]));
Q_ASSIGN U24764 ( .B(clk), .A(\g.we_clk [8010]));
Q_ASSIGN U24765 ( .B(clk), .A(\g.we_clk [8009]));
Q_ASSIGN U24766 ( .B(clk), .A(\g.we_clk [8008]));
Q_ASSIGN U24767 ( .B(clk), .A(\g.we_clk [8007]));
Q_ASSIGN U24768 ( .B(clk), .A(\g.we_clk [8006]));
Q_ASSIGN U24769 ( .B(clk), .A(\g.we_clk [8005]));
Q_ASSIGN U24770 ( .B(clk), .A(\g.we_clk [8004]));
Q_ASSIGN U24771 ( .B(clk), .A(\g.we_clk [8003]));
Q_ASSIGN U24772 ( .B(clk), .A(\g.we_clk [8002]));
Q_ASSIGN U24773 ( .B(clk), .A(\g.we_clk [8001]));
Q_ASSIGN U24774 ( .B(clk), .A(\g.we_clk [8000]));
Q_ASSIGN U24775 ( .B(clk), .A(\g.we_clk [7999]));
Q_ASSIGN U24776 ( .B(clk), .A(\g.we_clk [7998]));
Q_ASSIGN U24777 ( .B(clk), .A(\g.we_clk [7997]));
Q_ASSIGN U24778 ( .B(clk), .A(\g.we_clk [7996]));
Q_ASSIGN U24779 ( .B(clk), .A(\g.we_clk [7995]));
Q_ASSIGN U24780 ( .B(clk), .A(\g.we_clk [7994]));
Q_ASSIGN U24781 ( .B(clk), .A(\g.we_clk [7993]));
Q_ASSIGN U24782 ( .B(clk), .A(\g.we_clk [7992]));
Q_ASSIGN U24783 ( .B(clk), .A(\g.we_clk [7991]));
Q_ASSIGN U24784 ( .B(clk), .A(\g.we_clk [7990]));
Q_ASSIGN U24785 ( .B(clk), .A(\g.we_clk [7989]));
Q_ASSIGN U24786 ( .B(clk), .A(\g.we_clk [7988]));
Q_ASSIGN U24787 ( .B(clk), .A(\g.we_clk [7987]));
Q_ASSIGN U24788 ( .B(clk), .A(\g.we_clk [7986]));
Q_ASSIGN U24789 ( .B(clk), .A(\g.we_clk [7985]));
Q_ASSIGN U24790 ( .B(clk), .A(\g.we_clk [7984]));
Q_ASSIGN U24791 ( .B(clk), .A(\g.we_clk [7983]));
Q_ASSIGN U24792 ( .B(clk), .A(\g.we_clk [7982]));
Q_ASSIGN U24793 ( .B(clk), .A(\g.we_clk [7981]));
Q_ASSIGN U24794 ( .B(clk), .A(\g.we_clk [7980]));
Q_ASSIGN U24795 ( .B(clk), .A(\g.we_clk [7979]));
Q_ASSIGN U24796 ( .B(clk), .A(\g.we_clk [7978]));
Q_ASSIGN U24797 ( .B(clk), .A(\g.we_clk [7977]));
Q_ASSIGN U24798 ( .B(clk), .A(\g.we_clk [7976]));
Q_ASSIGN U24799 ( .B(clk), .A(\g.we_clk [7975]));
Q_ASSIGN U24800 ( .B(clk), .A(\g.we_clk [7974]));
Q_ASSIGN U24801 ( .B(clk), .A(\g.we_clk [7973]));
Q_ASSIGN U24802 ( .B(clk), .A(\g.we_clk [7972]));
Q_ASSIGN U24803 ( .B(clk), .A(\g.we_clk [7971]));
Q_ASSIGN U24804 ( .B(clk), .A(\g.we_clk [7970]));
Q_ASSIGN U24805 ( .B(clk), .A(\g.we_clk [7969]));
Q_ASSIGN U24806 ( .B(clk), .A(\g.we_clk [7968]));
Q_ASSIGN U24807 ( .B(clk), .A(\g.we_clk [7967]));
Q_ASSIGN U24808 ( .B(clk), .A(\g.we_clk [7966]));
Q_ASSIGN U24809 ( .B(clk), .A(\g.we_clk [7965]));
Q_ASSIGN U24810 ( .B(clk), .A(\g.we_clk [7964]));
Q_ASSIGN U24811 ( .B(clk), .A(\g.we_clk [7963]));
Q_ASSIGN U24812 ( .B(clk), .A(\g.we_clk [7962]));
Q_ASSIGN U24813 ( .B(clk), .A(\g.we_clk [7961]));
Q_ASSIGN U24814 ( .B(clk), .A(\g.we_clk [7960]));
Q_ASSIGN U24815 ( .B(clk), .A(\g.we_clk [7959]));
Q_ASSIGN U24816 ( .B(clk), .A(\g.we_clk [7958]));
Q_ASSIGN U24817 ( .B(clk), .A(\g.we_clk [7957]));
Q_ASSIGN U24818 ( .B(clk), .A(\g.we_clk [7956]));
Q_ASSIGN U24819 ( .B(clk), .A(\g.we_clk [7955]));
Q_ASSIGN U24820 ( .B(clk), .A(\g.we_clk [7954]));
Q_ASSIGN U24821 ( .B(clk), .A(\g.we_clk [7953]));
Q_ASSIGN U24822 ( .B(clk), .A(\g.we_clk [7952]));
Q_ASSIGN U24823 ( .B(clk), .A(\g.we_clk [7951]));
Q_ASSIGN U24824 ( .B(clk), .A(\g.we_clk [7950]));
Q_ASSIGN U24825 ( .B(clk), .A(\g.we_clk [7949]));
Q_ASSIGN U24826 ( .B(clk), .A(\g.we_clk [7948]));
Q_ASSIGN U24827 ( .B(clk), .A(\g.we_clk [7947]));
Q_ASSIGN U24828 ( .B(clk), .A(\g.we_clk [7946]));
Q_ASSIGN U24829 ( .B(clk), .A(\g.we_clk [7945]));
Q_ASSIGN U24830 ( .B(clk), .A(\g.we_clk [7944]));
Q_ASSIGN U24831 ( .B(clk), .A(\g.we_clk [7943]));
Q_ASSIGN U24832 ( .B(clk), .A(\g.we_clk [7942]));
Q_ASSIGN U24833 ( .B(clk), .A(\g.we_clk [7941]));
Q_ASSIGN U24834 ( .B(clk), .A(\g.we_clk [7940]));
Q_ASSIGN U24835 ( .B(clk), .A(\g.we_clk [7939]));
Q_ASSIGN U24836 ( .B(clk), .A(\g.we_clk [7938]));
Q_ASSIGN U24837 ( .B(clk), .A(\g.we_clk [7937]));
Q_ASSIGN U24838 ( .B(clk), .A(\g.we_clk [7936]));
Q_ASSIGN U24839 ( .B(clk), .A(\g.we_clk [7935]));
Q_ASSIGN U24840 ( .B(clk), .A(\g.we_clk [7934]));
Q_ASSIGN U24841 ( .B(clk), .A(\g.we_clk [7933]));
Q_ASSIGN U24842 ( .B(clk), .A(\g.we_clk [7932]));
Q_ASSIGN U24843 ( .B(clk), .A(\g.we_clk [7931]));
Q_ASSIGN U24844 ( .B(clk), .A(\g.we_clk [7930]));
Q_ASSIGN U24845 ( .B(clk), .A(\g.we_clk [7929]));
Q_ASSIGN U24846 ( .B(clk), .A(\g.we_clk [7928]));
Q_ASSIGN U24847 ( .B(clk), .A(\g.we_clk [7927]));
Q_ASSIGN U24848 ( .B(clk), .A(\g.we_clk [7926]));
Q_ASSIGN U24849 ( .B(clk), .A(\g.we_clk [7925]));
Q_ASSIGN U24850 ( .B(clk), .A(\g.we_clk [7924]));
Q_ASSIGN U24851 ( .B(clk), .A(\g.we_clk [7923]));
Q_ASSIGN U24852 ( .B(clk), .A(\g.we_clk [7922]));
Q_ASSIGN U24853 ( .B(clk), .A(\g.we_clk [7921]));
Q_ASSIGN U24854 ( .B(clk), .A(\g.we_clk [7920]));
Q_ASSIGN U24855 ( .B(clk), .A(\g.we_clk [7919]));
Q_ASSIGN U24856 ( .B(clk), .A(\g.we_clk [7918]));
Q_ASSIGN U24857 ( .B(clk), .A(\g.we_clk [7917]));
Q_ASSIGN U24858 ( .B(clk), .A(\g.we_clk [7916]));
Q_ASSIGN U24859 ( .B(clk), .A(\g.we_clk [7915]));
Q_ASSIGN U24860 ( .B(clk), .A(\g.we_clk [7914]));
Q_ASSIGN U24861 ( .B(clk), .A(\g.we_clk [7913]));
Q_ASSIGN U24862 ( .B(clk), .A(\g.we_clk [7912]));
Q_ASSIGN U24863 ( .B(clk), .A(\g.we_clk [7911]));
Q_ASSIGN U24864 ( .B(clk), .A(\g.we_clk [7910]));
Q_ASSIGN U24865 ( .B(clk), .A(\g.we_clk [7909]));
Q_ASSIGN U24866 ( .B(clk), .A(\g.we_clk [7908]));
Q_ASSIGN U24867 ( .B(clk), .A(\g.we_clk [7907]));
Q_ASSIGN U24868 ( .B(clk), .A(\g.we_clk [7906]));
Q_ASSIGN U24869 ( .B(clk), .A(\g.we_clk [7905]));
Q_ASSIGN U24870 ( .B(clk), .A(\g.we_clk [7904]));
Q_ASSIGN U24871 ( .B(clk), .A(\g.we_clk [7903]));
Q_ASSIGN U24872 ( .B(clk), .A(\g.we_clk [7902]));
Q_ASSIGN U24873 ( .B(clk), .A(\g.we_clk [7901]));
Q_ASSIGN U24874 ( .B(clk), .A(\g.we_clk [7900]));
Q_ASSIGN U24875 ( .B(clk), .A(\g.we_clk [7899]));
Q_ASSIGN U24876 ( .B(clk), .A(\g.we_clk [7898]));
Q_ASSIGN U24877 ( .B(clk), .A(\g.we_clk [7897]));
Q_ASSIGN U24878 ( .B(clk), .A(\g.we_clk [7896]));
Q_ASSIGN U24879 ( .B(clk), .A(\g.we_clk [7895]));
Q_ASSIGN U24880 ( .B(clk), .A(\g.we_clk [7894]));
Q_ASSIGN U24881 ( .B(clk), .A(\g.we_clk [7893]));
Q_ASSIGN U24882 ( .B(clk), .A(\g.we_clk [7892]));
Q_ASSIGN U24883 ( .B(clk), .A(\g.we_clk [7891]));
Q_ASSIGN U24884 ( .B(clk), .A(\g.we_clk [7890]));
Q_ASSIGN U24885 ( .B(clk), .A(\g.we_clk [7889]));
Q_ASSIGN U24886 ( .B(clk), .A(\g.we_clk [7888]));
Q_ASSIGN U24887 ( .B(clk), .A(\g.we_clk [7887]));
Q_ASSIGN U24888 ( .B(clk), .A(\g.we_clk [7886]));
Q_ASSIGN U24889 ( .B(clk), .A(\g.we_clk [7885]));
Q_ASSIGN U24890 ( .B(clk), .A(\g.we_clk [7884]));
Q_ASSIGN U24891 ( .B(clk), .A(\g.we_clk [7883]));
Q_ASSIGN U24892 ( .B(clk), .A(\g.we_clk [7882]));
Q_ASSIGN U24893 ( .B(clk), .A(\g.we_clk [7881]));
Q_ASSIGN U24894 ( .B(clk), .A(\g.we_clk [7880]));
Q_ASSIGN U24895 ( .B(clk), .A(\g.we_clk [7879]));
Q_ASSIGN U24896 ( .B(clk), .A(\g.we_clk [7878]));
Q_ASSIGN U24897 ( .B(clk), .A(\g.we_clk [7877]));
Q_ASSIGN U24898 ( .B(clk), .A(\g.we_clk [7876]));
Q_ASSIGN U24899 ( .B(clk), .A(\g.we_clk [7875]));
Q_ASSIGN U24900 ( .B(clk), .A(\g.we_clk [7874]));
Q_ASSIGN U24901 ( .B(clk), .A(\g.we_clk [7873]));
Q_ASSIGN U24902 ( .B(clk), .A(\g.we_clk [7872]));
Q_ASSIGN U24903 ( .B(clk), .A(\g.we_clk [7871]));
Q_ASSIGN U24904 ( .B(clk), .A(\g.we_clk [7870]));
Q_ASSIGN U24905 ( .B(clk), .A(\g.we_clk [7869]));
Q_ASSIGN U24906 ( .B(clk), .A(\g.we_clk [7868]));
Q_ASSIGN U24907 ( .B(clk), .A(\g.we_clk [7867]));
Q_ASSIGN U24908 ( .B(clk), .A(\g.we_clk [7866]));
Q_ASSIGN U24909 ( .B(clk), .A(\g.we_clk [7865]));
Q_ASSIGN U24910 ( .B(clk), .A(\g.we_clk [7864]));
Q_ASSIGN U24911 ( .B(clk), .A(\g.we_clk [7863]));
Q_ASSIGN U24912 ( .B(clk), .A(\g.we_clk [7862]));
Q_ASSIGN U24913 ( .B(clk), .A(\g.we_clk [7861]));
Q_ASSIGN U24914 ( .B(clk), .A(\g.we_clk [7860]));
Q_ASSIGN U24915 ( .B(clk), .A(\g.we_clk [7859]));
Q_ASSIGN U24916 ( .B(clk), .A(\g.we_clk [7858]));
Q_ASSIGN U24917 ( .B(clk), .A(\g.we_clk [7857]));
Q_ASSIGN U24918 ( .B(clk), .A(\g.we_clk [7856]));
Q_ASSIGN U24919 ( .B(clk), .A(\g.we_clk [7855]));
Q_ASSIGN U24920 ( .B(clk), .A(\g.we_clk [7854]));
Q_ASSIGN U24921 ( .B(clk), .A(\g.we_clk [7853]));
Q_ASSIGN U24922 ( .B(clk), .A(\g.we_clk [7852]));
Q_ASSIGN U24923 ( .B(clk), .A(\g.we_clk [7851]));
Q_ASSIGN U24924 ( .B(clk), .A(\g.we_clk [7850]));
Q_ASSIGN U24925 ( .B(clk), .A(\g.we_clk [7849]));
Q_ASSIGN U24926 ( .B(clk), .A(\g.we_clk [7848]));
Q_ASSIGN U24927 ( .B(clk), .A(\g.we_clk [7847]));
Q_ASSIGN U24928 ( .B(clk), .A(\g.we_clk [7846]));
Q_ASSIGN U24929 ( .B(clk), .A(\g.we_clk [7845]));
Q_ASSIGN U24930 ( .B(clk), .A(\g.we_clk [7844]));
Q_ASSIGN U24931 ( .B(clk), .A(\g.we_clk [7843]));
Q_ASSIGN U24932 ( .B(clk), .A(\g.we_clk [7842]));
Q_ASSIGN U24933 ( .B(clk), .A(\g.we_clk [7841]));
Q_ASSIGN U24934 ( .B(clk), .A(\g.we_clk [7840]));
Q_ASSIGN U24935 ( .B(clk), .A(\g.we_clk [7839]));
Q_ASSIGN U24936 ( .B(clk), .A(\g.we_clk [7838]));
Q_ASSIGN U24937 ( .B(clk), .A(\g.we_clk [7837]));
Q_ASSIGN U24938 ( .B(clk), .A(\g.we_clk [7836]));
Q_ASSIGN U24939 ( .B(clk), .A(\g.we_clk [7835]));
Q_ASSIGN U24940 ( .B(clk), .A(\g.we_clk [7834]));
Q_ASSIGN U24941 ( .B(clk), .A(\g.we_clk [7833]));
Q_ASSIGN U24942 ( .B(clk), .A(\g.we_clk [7832]));
Q_ASSIGN U24943 ( .B(clk), .A(\g.we_clk [7831]));
Q_ASSIGN U24944 ( .B(clk), .A(\g.we_clk [7830]));
Q_ASSIGN U24945 ( .B(clk), .A(\g.we_clk [7829]));
Q_ASSIGN U24946 ( .B(clk), .A(\g.we_clk [7828]));
Q_ASSIGN U24947 ( .B(clk), .A(\g.we_clk [7827]));
Q_ASSIGN U24948 ( .B(clk), .A(\g.we_clk [7826]));
Q_ASSIGN U24949 ( .B(clk), .A(\g.we_clk [7825]));
Q_ASSIGN U24950 ( .B(clk), .A(\g.we_clk [7824]));
Q_ASSIGN U24951 ( .B(clk), .A(\g.we_clk [7823]));
Q_ASSIGN U24952 ( .B(clk), .A(\g.we_clk [7822]));
Q_ASSIGN U24953 ( .B(clk), .A(\g.we_clk [7821]));
Q_ASSIGN U24954 ( .B(clk), .A(\g.we_clk [7820]));
Q_ASSIGN U24955 ( .B(clk), .A(\g.we_clk [7819]));
Q_ASSIGN U24956 ( .B(clk), .A(\g.we_clk [7818]));
Q_ASSIGN U24957 ( .B(clk), .A(\g.we_clk [7817]));
Q_ASSIGN U24958 ( .B(clk), .A(\g.we_clk [7816]));
Q_ASSIGN U24959 ( .B(clk), .A(\g.we_clk [7815]));
Q_ASSIGN U24960 ( .B(clk), .A(\g.we_clk [7814]));
Q_ASSIGN U24961 ( .B(clk), .A(\g.we_clk [7813]));
Q_ASSIGN U24962 ( .B(clk), .A(\g.we_clk [7812]));
Q_ASSIGN U24963 ( .B(clk), .A(\g.we_clk [7811]));
Q_ASSIGN U24964 ( .B(clk), .A(\g.we_clk [7810]));
Q_ASSIGN U24965 ( .B(clk), .A(\g.we_clk [7809]));
Q_ASSIGN U24966 ( .B(clk), .A(\g.we_clk [7808]));
Q_ASSIGN U24967 ( .B(clk), .A(\g.we_clk [7807]));
Q_ASSIGN U24968 ( .B(clk), .A(\g.we_clk [7806]));
Q_ASSIGN U24969 ( .B(clk), .A(\g.we_clk [7805]));
Q_ASSIGN U24970 ( .B(clk), .A(\g.we_clk [7804]));
Q_ASSIGN U24971 ( .B(clk), .A(\g.we_clk [7803]));
Q_ASSIGN U24972 ( .B(clk), .A(\g.we_clk [7802]));
Q_ASSIGN U24973 ( .B(clk), .A(\g.we_clk [7801]));
Q_ASSIGN U24974 ( .B(clk), .A(\g.we_clk [7800]));
Q_ASSIGN U24975 ( .B(clk), .A(\g.we_clk [7799]));
Q_ASSIGN U24976 ( .B(clk), .A(\g.we_clk [7798]));
Q_ASSIGN U24977 ( .B(clk), .A(\g.we_clk [7797]));
Q_ASSIGN U24978 ( .B(clk), .A(\g.we_clk [7796]));
Q_ASSIGN U24979 ( .B(clk), .A(\g.we_clk [7795]));
Q_ASSIGN U24980 ( .B(clk), .A(\g.we_clk [7794]));
Q_ASSIGN U24981 ( .B(clk), .A(\g.we_clk [7793]));
Q_ASSIGN U24982 ( .B(clk), .A(\g.we_clk [7792]));
Q_ASSIGN U24983 ( .B(clk), .A(\g.we_clk [7791]));
Q_ASSIGN U24984 ( .B(clk), .A(\g.we_clk [7790]));
Q_ASSIGN U24985 ( .B(clk), .A(\g.we_clk [7789]));
Q_ASSIGN U24986 ( .B(clk), .A(\g.we_clk [7788]));
Q_ASSIGN U24987 ( .B(clk), .A(\g.we_clk [7787]));
Q_ASSIGN U24988 ( .B(clk), .A(\g.we_clk [7786]));
Q_ASSIGN U24989 ( .B(clk), .A(\g.we_clk [7785]));
Q_ASSIGN U24990 ( .B(clk), .A(\g.we_clk [7784]));
Q_ASSIGN U24991 ( .B(clk), .A(\g.we_clk [7783]));
Q_ASSIGN U24992 ( .B(clk), .A(\g.we_clk [7782]));
Q_ASSIGN U24993 ( .B(clk), .A(\g.we_clk [7781]));
Q_ASSIGN U24994 ( .B(clk), .A(\g.we_clk [7780]));
Q_ASSIGN U24995 ( .B(clk), .A(\g.we_clk [7779]));
Q_ASSIGN U24996 ( .B(clk), .A(\g.we_clk [7778]));
Q_ASSIGN U24997 ( .B(clk), .A(\g.we_clk [7777]));
Q_ASSIGN U24998 ( .B(clk), .A(\g.we_clk [7776]));
Q_ASSIGN U24999 ( .B(clk), .A(\g.we_clk [7775]));
Q_ASSIGN U25000 ( .B(clk), .A(\g.we_clk [7774]));
Q_ASSIGN U25001 ( .B(clk), .A(\g.we_clk [7773]));
Q_ASSIGN U25002 ( .B(clk), .A(\g.we_clk [7772]));
Q_ASSIGN U25003 ( .B(clk), .A(\g.we_clk [7771]));
Q_ASSIGN U25004 ( .B(clk), .A(\g.we_clk [7770]));
Q_ASSIGN U25005 ( .B(clk), .A(\g.we_clk [7769]));
Q_ASSIGN U25006 ( .B(clk), .A(\g.we_clk [7768]));
Q_ASSIGN U25007 ( .B(clk), .A(\g.we_clk [7767]));
Q_ASSIGN U25008 ( .B(clk), .A(\g.we_clk [7766]));
Q_ASSIGN U25009 ( .B(clk), .A(\g.we_clk [7765]));
Q_ASSIGN U25010 ( .B(clk), .A(\g.we_clk [7764]));
Q_ASSIGN U25011 ( .B(clk), .A(\g.we_clk [7763]));
Q_ASSIGN U25012 ( .B(clk), .A(\g.we_clk [7762]));
Q_ASSIGN U25013 ( .B(clk), .A(\g.we_clk [7761]));
Q_ASSIGN U25014 ( .B(clk), .A(\g.we_clk [7760]));
Q_ASSIGN U25015 ( .B(clk), .A(\g.we_clk [7759]));
Q_ASSIGN U25016 ( .B(clk), .A(\g.we_clk [7758]));
Q_ASSIGN U25017 ( .B(clk), .A(\g.we_clk [7757]));
Q_ASSIGN U25018 ( .B(clk), .A(\g.we_clk [7756]));
Q_ASSIGN U25019 ( .B(clk), .A(\g.we_clk [7755]));
Q_ASSIGN U25020 ( .B(clk), .A(\g.we_clk [7754]));
Q_ASSIGN U25021 ( .B(clk), .A(\g.we_clk [7753]));
Q_ASSIGN U25022 ( .B(clk), .A(\g.we_clk [7752]));
Q_ASSIGN U25023 ( .B(clk), .A(\g.we_clk [7751]));
Q_ASSIGN U25024 ( .B(clk), .A(\g.we_clk [7750]));
Q_ASSIGN U25025 ( .B(clk), .A(\g.we_clk [7749]));
Q_ASSIGN U25026 ( .B(clk), .A(\g.we_clk [7748]));
Q_ASSIGN U25027 ( .B(clk), .A(\g.we_clk [7747]));
Q_ASSIGN U25028 ( .B(clk), .A(\g.we_clk [7746]));
Q_ASSIGN U25029 ( .B(clk), .A(\g.we_clk [7745]));
Q_ASSIGN U25030 ( .B(clk), .A(\g.we_clk [7744]));
Q_ASSIGN U25031 ( .B(clk), .A(\g.we_clk [7743]));
Q_ASSIGN U25032 ( .B(clk), .A(\g.we_clk [7742]));
Q_ASSIGN U25033 ( .B(clk), .A(\g.we_clk [7741]));
Q_ASSIGN U25034 ( .B(clk), .A(\g.we_clk [7740]));
Q_ASSIGN U25035 ( .B(clk), .A(\g.we_clk [7739]));
Q_ASSIGN U25036 ( .B(clk), .A(\g.we_clk [7738]));
Q_ASSIGN U25037 ( .B(clk), .A(\g.we_clk [7737]));
Q_ASSIGN U25038 ( .B(clk), .A(\g.we_clk [7736]));
Q_ASSIGN U25039 ( .B(clk), .A(\g.we_clk [7735]));
Q_ASSIGN U25040 ( .B(clk), .A(\g.we_clk [7734]));
Q_ASSIGN U25041 ( .B(clk), .A(\g.we_clk [7733]));
Q_ASSIGN U25042 ( .B(clk), .A(\g.we_clk [7732]));
Q_ASSIGN U25043 ( .B(clk), .A(\g.we_clk [7731]));
Q_ASSIGN U25044 ( .B(clk), .A(\g.we_clk [7730]));
Q_ASSIGN U25045 ( .B(clk), .A(\g.we_clk [7729]));
Q_ASSIGN U25046 ( .B(clk), .A(\g.we_clk [7728]));
Q_ASSIGN U25047 ( .B(clk), .A(\g.we_clk [7727]));
Q_ASSIGN U25048 ( .B(clk), .A(\g.we_clk [7726]));
Q_ASSIGN U25049 ( .B(clk), .A(\g.we_clk [7725]));
Q_ASSIGN U25050 ( .B(clk), .A(\g.we_clk [7724]));
Q_ASSIGN U25051 ( .B(clk), .A(\g.we_clk [7723]));
Q_ASSIGN U25052 ( .B(clk), .A(\g.we_clk [7722]));
Q_ASSIGN U25053 ( .B(clk), .A(\g.we_clk [7721]));
Q_ASSIGN U25054 ( .B(clk), .A(\g.we_clk [7720]));
Q_ASSIGN U25055 ( .B(clk), .A(\g.we_clk [7719]));
Q_ASSIGN U25056 ( .B(clk), .A(\g.we_clk [7718]));
Q_ASSIGN U25057 ( .B(clk), .A(\g.we_clk [7717]));
Q_ASSIGN U25058 ( .B(clk), .A(\g.we_clk [7716]));
Q_ASSIGN U25059 ( .B(clk), .A(\g.we_clk [7715]));
Q_ASSIGN U25060 ( .B(clk), .A(\g.we_clk [7714]));
Q_ASSIGN U25061 ( .B(clk), .A(\g.we_clk [7713]));
Q_ASSIGN U25062 ( .B(clk), .A(\g.we_clk [7712]));
Q_ASSIGN U25063 ( .B(clk), .A(\g.we_clk [7711]));
Q_ASSIGN U25064 ( .B(clk), .A(\g.we_clk [7710]));
Q_ASSIGN U25065 ( .B(clk), .A(\g.we_clk [7709]));
Q_ASSIGN U25066 ( .B(clk), .A(\g.we_clk [7708]));
Q_ASSIGN U25067 ( .B(clk), .A(\g.we_clk [7707]));
Q_ASSIGN U25068 ( .B(clk), .A(\g.we_clk [7706]));
Q_ASSIGN U25069 ( .B(clk), .A(\g.we_clk [7705]));
Q_ASSIGN U25070 ( .B(clk), .A(\g.we_clk [7704]));
Q_ASSIGN U25071 ( .B(clk), .A(\g.we_clk [7703]));
Q_ASSIGN U25072 ( .B(clk), .A(\g.we_clk [7702]));
Q_ASSIGN U25073 ( .B(clk), .A(\g.we_clk [7701]));
Q_ASSIGN U25074 ( .B(clk), .A(\g.we_clk [7700]));
Q_ASSIGN U25075 ( .B(clk), .A(\g.we_clk [7699]));
Q_ASSIGN U25076 ( .B(clk), .A(\g.we_clk [7698]));
Q_ASSIGN U25077 ( .B(clk), .A(\g.we_clk [7697]));
Q_ASSIGN U25078 ( .B(clk), .A(\g.we_clk [7696]));
Q_ASSIGN U25079 ( .B(clk), .A(\g.we_clk [7695]));
Q_ASSIGN U25080 ( .B(clk), .A(\g.we_clk [7694]));
Q_ASSIGN U25081 ( .B(clk), .A(\g.we_clk [7693]));
Q_ASSIGN U25082 ( .B(clk), .A(\g.we_clk [7692]));
Q_ASSIGN U25083 ( .B(clk), .A(\g.we_clk [7691]));
Q_ASSIGN U25084 ( .B(clk), .A(\g.we_clk [7690]));
Q_ASSIGN U25085 ( .B(clk), .A(\g.we_clk [7689]));
Q_ASSIGN U25086 ( .B(clk), .A(\g.we_clk [7688]));
Q_ASSIGN U25087 ( .B(clk), .A(\g.we_clk [7687]));
Q_ASSIGN U25088 ( .B(clk), .A(\g.we_clk [7686]));
Q_ASSIGN U25089 ( .B(clk), .A(\g.we_clk [7685]));
Q_ASSIGN U25090 ( .B(clk), .A(\g.we_clk [7684]));
Q_ASSIGN U25091 ( .B(clk), .A(\g.we_clk [7683]));
Q_ASSIGN U25092 ( .B(clk), .A(\g.we_clk [7682]));
Q_ASSIGN U25093 ( .B(clk), .A(\g.we_clk [7681]));
Q_ASSIGN U25094 ( .B(clk), .A(\g.we_clk [7680]));
Q_ASSIGN U25095 ( .B(clk), .A(\g.we_clk [7679]));
Q_ASSIGN U25096 ( .B(clk), .A(\g.we_clk [7678]));
Q_ASSIGN U25097 ( .B(clk), .A(\g.we_clk [7677]));
Q_ASSIGN U25098 ( .B(clk), .A(\g.we_clk [7676]));
Q_ASSIGN U25099 ( .B(clk), .A(\g.we_clk [7675]));
Q_ASSIGN U25100 ( .B(clk), .A(\g.we_clk [7674]));
Q_ASSIGN U25101 ( .B(clk), .A(\g.we_clk [7673]));
Q_ASSIGN U25102 ( .B(clk), .A(\g.we_clk [7672]));
Q_ASSIGN U25103 ( .B(clk), .A(\g.we_clk [7671]));
Q_ASSIGN U25104 ( .B(clk), .A(\g.we_clk [7670]));
Q_ASSIGN U25105 ( .B(clk), .A(\g.we_clk [7669]));
Q_ASSIGN U25106 ( .B(clk), .A(\g.we_clk [7668]));
Q_ASSIGN U25107 ( .B(clk), .A(\g.we_clk [7667]));
Q_ASSIGN U25108 ( .B(clk), .A(\g.we_clk [7666]));
Q_ASSIGN U25109 ( .B(clk), .A(\g.we_clk [7665]));
Q_ASSIGN U25110 ( .B(clk), .A(\g.we_clk [7664]));
Q_ASSIGN U25111 ( .B(clk), .A(\g.we_clk [7663]));
Q_ASSIGN U25112 ( .B(clk), .A(\g.we_clk [7662]));
Q_ASSIGN U25113 ( .B(clk), .A(\g.we_clk [7661]));
Q_ASSIGN U25114 ( .B(clk), .A(\g.we_clk [7660]));
Q_ASSIGN U25115 ( .B(clk), .A(\g.we_clk [7659]));
Q_ASSIGN U25116 ( .B(clk), .A(\g.we_clk [7658]));
Q_ASSIGN U25117 ( .B(clk), .A(\g.we_clk [7657]));
Q_ASSIGN U25118 ( .B(clk), .A(\g.we_clk [7656]));
Q_ASSIGN U25119 ( .B(clk), .A(\g.we_clk [7655]));
Q_ASSIGN U25120 ( .B(clk), .A(\g.we_clk [7654]));
Q_ASSIGN U25121 ( .B(clk), .A(\g.we_clk [7653]));
Q_ASSIGN U25122 ( .B(clk), .A(\g.we_clk [7652]));
Q_ASSIGN U25123 ( .B(clk), .A(\g.we_clk [7651]));
Q_ASSIGN U25124 ( .B(clk), .A(\g.we_clk [7650]));
Q_ASSIGN U25125 ( .B(clk), .A(\g.we_clk [7649]));
Q_ASSIGN U25126 ( .B(clk), .A(\g.we_clk [7648]));
Q_ASSIGN U25127 ( .B(clk), .A(\g.we_clk [7647]));
Q_ASSIGN U25128 ( .B(clk), .A(\g.we_clk [7646]));
Q_ASSIGN U25129 ( .B(clk), .A(\g.we_clk [7645]));
Q_ASSIGN U25130 ( .B(clk), .A(\g.we_clk [7644]));
Q_ASSIGN U25131 ( .B(clk), .A(\g.we_clk [7643]));
Q_ASSIGN U25132 ( .B(clk), .A(\g.we_clk [7642]));
Q_ASSIGN U25133 ( .B(clk), .A(\g.we_clk [7641]));
Q_ASSIGN U25134 ( .B(clk), .A(\g.we_clk [7640]));
Q_ASSIGN U25135 ( .B(clk), .A(\g.we_clk [7639]));
Q_ASSIGN U25136 ( .B(clk), .A(\g.we_clk [7638]));
Q_ASSIGN U25137 ( .B(clk), .A(\g.we_clk [7637]));
Q_ASSIGN U25138 ( .B(clk), .A(\g.we_clk [7636]));
Q_ASSIGN U25139 ( .B(clk), .A(\g.we_clk [7635]));
Q_ASSIGN U25140 ( .B(clk), .A(\g.we_clk [7634]));
Q_ASSIGN U25141 ( .B(clk), .A(\g.we_clk [7633]));
Q_ASSIGN U25142 ( .B(clk), .A(\g.we_clk [7632]));
Q_ASSIGN U25143 ( .B(clk), .A(\g.we_clk [7631]));
Q_ASSIGN U25144 ( .B(clk), .A(\g.we_clk [7630]));
Q_ASSIGN U25145 ( .B(clk), .A(\g.we_clk [7629]));
Q_ASSIGN U25146 ( .B(clk), .A(\g.we_clk [7628]));
Q_ASSIGN U25147 ( .B(clk), .A(\g.we_clk [7627]));
Q_ASSIGN U25148 ( .B(clk), .A(\g.we_clk [7626]));
Q_ASSIGN U25149 ( .B(clk), .A(\g.we_clk [7625]));
Q_ASSIGN U25150 ( .B(clk), .A(\g.we_clk [7624]));
Q_ASSIGN U25151 ( .B(clk), .A(\g.we_clk [7623]));
Q_ASSIGN U25152 ( .B(clk), .A(\g.we_clk [7622]));
Q_ASSIGN U25153 ( .B(clk), .A(\g.we_clk [7621]));
Q_ASSIGN U25154 ( .B(clk), .A(\g.we_clk [7620]));
Q_ASSIGN U25155 ( .B(clk), .A(\g.we_clk [7619]));
Q_ASSIGN U25156 ( .B(clk), .A(\g.we_clk [7618]));
Q_ASSIGN U25157 ( .B(clk), .A(\g.we_clk [7617]));
Q_ASSIGN U25158 ( .B(clk), .A(\g.we_clk [7616]));
Q_ASSIGN U25159 ( .B(clk), .A(\g.we_clk [7615]));
Q_ASSIGN U25160 ( .B(clk), .A(\g.we_clk [7614]));
Q_ASSIGN U25161 ( .B(clk), .A(\g.we_clk [7613]));
Q_ASSIGN U25162 ( .B(clk), .A(\g.we_clk [7612]));
Q_ASSIGN U25163 ( .B(clk), .A(\g.we_clk [7611]));
Q_ASSIGN U25164 ( .B(clk), .A(\g.we_clk [7610]));
Q_ASSIGN U25165 ( .B(clk), .A(\g.we_clk [7609]));
Q_ASSIGN U25166 ( .B(clk), .A(\g.we_clk [7608]));
Q_ASSIGN U25167 ( .B(clk), .A(\g.we_clk [7607]));
Q_ASSIGN U25168 ( .B(clk), .A(\g.we_clk [7606]));
Q_ASSIGN U25169 ( .B(clk), .A(\g.we_clk [7605]));
Q_ASSIGN U25170 ( .B(clk), .A(\g.we_clk [7604]));
Q_ASSIGN U25171 ( .B(clk), .A(\g.we_clk [7603]));
Q_ASSIGN U25172 ( .B(clk), .A(\g.we_clk [7602]));
Q_ASSIGN U25173 ( .B(clk), .A(\g.we_clk [7601]));
Q_ASSIGN U25174 ( .B(clk), .A(\g.we_clk [7600]));
Q_ASSIGN U25175 ( .B(clk), .A(\g.we_clk [7599]));
Q_ASSIGN U25176 ( .B(clk), .A(\g.we_clk [7598]));
Q_ASSIGN U25177 ( .B(clk), .A(\g.we_clk [7597]));
Q_ASSIGN U25178 ( .B(clk), .A(\g.we_clk [7596]));
Q_ASSIGN U25179 ( .B(clk), .A(\g.we_clk [7595]));
Q_ASSIGN U25180 ( .B(clk), .A(\g.we_clk [7594]));
Q_ASSIGN U25181 ( .B(clk), .A(\g.we_clk [7593]));
Q_ASSIGN U25182 ( .B(clk), .A(\g.we_clk [7592]));
Q_ASSIGN U25183 ( .B(clk), .A(\g.we_clk [7591]));
Q_ASSIGN U25184 ( .B(clk), .A(\g.we_clk [7590]));
Q_ASSIGN U25185 ( .B(clk), .A(\g.we_clk [7589]));
Q_ASSIGN U25186 ( .B(clk), .A(\g.we_clk [7588]));
Q_ASSIGN U25187 ( .B(clk), .A(\g.we_clk [7587]));
Q_ASSIGN U25188 ( .B(clk), .A(\g.we_clk [7586]));
Q_ASSIGN U25189 ( .B(clk), .A(\g.we_clk [7585]));
Q_ASSIGN U25190 ( .B(clk), .A(\g.we_clk [7584]));
Q_ASSIGN U25191 ( .B(clk), .A(\g.we_clk [7583]));
Q_ASSIGN U25192 ( .B(clk), .A(\g.we_clk [7582]));
Q_ASSIGN U25193 ( .B(clk), .A(\g.we_clk [7581]));
Q_ASSIGN U25194 ( .B(clk), .A(\g.we_clk [7580]));
Q_ASSIGN U25195 ( .B(clk), .A(\g.we_clk [7579]));
Q_ASSIGN U25196 ( .B(clk), .A(\g.we_clk [7578]));
Q_ASSIGN U25197 ( .B(clk), .A(\g.we_clk [7577]));
Q_ASSIGN U25198 ( .B(clk), .A(\g.we_clk [7576]));
Q_ASSIGN U25199 ( .B(clk), .A(\g.we_clk [7575]));
Q_ASSIGN U25200 ( .B(clk), .A(\g.we_clk [7574]));
Q_ASSIGN U25201 ( .B(clk), .A(\g.we_clk [7573]));
Q_ASSIGN U25202 ( .B(clk), .A(\g.we_clk [7572]));
Q_ASSIGN U25203 ( .B(clk), .A(\g.we_clk [7571]));
Q_ASSIGN U25204 ( .B(clk), .A(\g.we_clk [7570]));
Q_ASSIGN U25205 ( .B(clk), .A(\g.we_clk [7569]));
Q_ASSIGN U25206 ( .B(clk), .A(\g.we_clk [7568]));
Q_ASSIGN U25207 ( .B(clk), .A(\g.we_clk [7567]));
Q_ASSIGN U25208 ( .B(clk), .A(\g.we_clk [7566]));
Q_ASSIGN U25209 ( .B(clk), .A(\g.we_clk [7565]));
Q_ASSIGN U25210 ( .B(clk), .A(\g.we_clk [7564]));
Q_ASSIGN U25211 ( .B(clk), .A(\g.we_clk [7563]));
Q_ASSIGN U25212 ( .B(clk), .A(\g.we_clk [7562]));
Q_ASSIGN U25213 ( .B(clk), .A(\g.we_clk [7561]));
Q_ASSIGN U25214 ( .B(clk), .A(\g.we_clk [7560]));
Q_ASSIGN U25215 ( .B(clk), .A(\g.we_clk [7559]));
Q_ASSIGN U25216 ( .B(clk), .A(\g.we_clk [7558]));
Q_ASSIGN U25217 ( .B(clk), .A(\g.we_clk [7557]));
Q_ASSIGN U25218 ( .B(clk), .A(\g.we_clk [7556]));
Q_ASSIGN U25219 ( .B(clk), .A(\g.we_clk [7555]));
Q_ASSIGN U25220 ( .B(clk), .A(\g.we_clk [7554]));
Q_ASSIGN U25221 ( .B(clk), .A(\g.we_clk [7553]));
Q_ASSIGN U25222 ( .B(clk), .A(\g.we_clk [7552]));
Q_ASSIGN U25223 ( .B(clk), .A(\g.we_clk [7551]));
Q_ASSIGN U25224 ( .B(clk), .A(\g.we_clk [7550]));
Q_ASSIGN U25225 ( .B(clk), .A(\g.we_clk [7549]));
Q_ASSIGN U25226 ( .B(clk), .A(\g.we_clk [7548]));
Q_ASSIGN U25227 ( .B(clk), .A(\g.we_clk [7547]));
Q_ASSIGN U25228 ( .B(clk), .A(\g.we_clk [7546]));
Q_ASSIGN U25229 ( .B(clk), .A(\g.we_clk [7545]));
Q_ASSIGN U25230 ( .B(clk), .A(\g.we_clk [7544]));
Q_ASSIGN U25231 ( .B(clk), .A(\g.we_clk [7543]));
Q_ASSIGN U25232 ( .B(clk), .A(\g.we_clk [7542]));
Q_ASSIGN U25233 ( .B(clk), .A(\g.we_clk [7541]));
Q_ASSIGN U25234 ( .B(clk), .A(\g.we_clk [7540]));
Q_ASSIGN U25235 ( .B(clk), .A(\g.we_clk [7539]));
Q_ASSIGN U25236 ( .B(clk), .A(\g.we_clk [7538]));
Q_ASSIGN U25237 ( .B(clk), .A(\g.we_clk [7537]));
Q_ASSIGN U25238 ( .B(clk), .A(\g.we_clk [7536]));
Q_ASSIGN U25239 ( .B(clk), .A(\g.we_clk [7535]));
Q_ASSIGN U25240 ( .B(clk), .A(\g.we_clk [7534]));
Q_ASSIGN U25241 ( .B(clk), .A(\g.we_clk [7533]));
Q_ASSIGN U25242 ( .B(clk), .A(\g.we_clk [7532]));
Q_ASSIGN U25243 ( .B(clk), .A(\g.we_clk [7531]));
Q_ASSIGN U25244 ( .B(clk), .A(\g.we_clk [7530]));
Q_ASSIGN U25245 ( .B(clk), .A(\g.we_clk [7529]));
Q_ASSIGN U25246 ( .B(clk), .A(\g.we_clk [7528]));
Q_ASSIGN U25247 ( .B(clk), .A(\g.we_clk [7527]));
Q_ASSIGN U25248 ( .B(clk), .A(\g.we_clk [7526]));
Q_ASSIGN U25249 ( .B(clk), .A(\g.we_clk [7525]));
Q_ASSIGN U25250 ( .B(clk), .A(\g.we_clk [7524]));
Q_ASSIGN U25251 ( .B(clk), .A(\g.we_clk [7523]));
Q_ASSIGN U25252 ( .B(clk), .A(\g.we_clk [7522]));
Q_ASSIGN U25253 ( .B(clk), .A(\g.we_clk [7521]));
Q_ASSIGN U25254 ( .B(clk), .A(\g.we_clk [7520]));
Q_ASSIGN U25255 ( .B(clk), .A(\g.we_clk [7519]));
Q_ASSIGN U25256 ( .B(clk), .A(\g.we_clk [7518]));
Q_ASSIGN U25257 ( .B(clk), .A(\g.we_clk [7517]));
Q_ASSIGN U25258 ( .B(clk), .A(\g.we_clk [7516]));
Q_ASSIGN U25259 ( .B(clk), .A(\g.we_clk [7515]));
Q_ASSIGN U25260 ( .B(clk), .A(\g.we_clk [7514]));
Q_ASSIGN U25261 ( .B(clk), .A(\g.we_clk [7513]));
Q_ASSIGN U25262 ( .B(clk), .A(\g.we_clk [7512]));
Q_ASSIGN U25263 ( .B(clk), .A(\g.we_clk [7511]));
Q_ASSIGN U25264 ( .B(clk), .A(\g.we_clk [7510]));
Q_ASSIGN U25265 ( .B(clk), .A(\g.we_clk [7509]));
Q_ASSIGN U25266 ( .B(clk), .A(\g.we_clk [7508]));
Q_ASSIGN U25267 ( .B(clk), .A(\g.we_clk [7507]));
Q_ASSIGN U25268 ( .B(clk), .A(\g.we_clk [7506]));
Q_ASSIGN U25269 ( .B(clk), .A(\g.we_clk [7505]));
Q_ASSIGN U25270 ( .B(clk), .A(\g.we_clk [7504]));
Q_ASSIGN U25271 ( .B(clk), .A(\g.we_clk [7503]));
Q_ASSIGN U25272 ( .B(clk), .A(\g.we_clk [7502]));
Q_ASSIGN U25273 ( .B(clk), .A(\g.we_clk [7501]));
Q_ASSIGN U25274 ( .B(clk), .A(\g.we_clk [7500]));
Q_ASSIGN U25275 ( .B(clk), .A(\g.we_clk [7499]));
Q_ASSIGN U25276 ( .B(clk), .A(\g.we_clk [7498]));
Q_ASSIGN U25277 ( .B(clk), .A(\g.we_clk [7497]));
Q_ASSIGN U25278 ( .B(clk), .A(\g.we_clk [7496]));
Q_ASSIGN U25279 ( .B(clk), .A(\g.we_clk [7495]));
Q_ASSIGN U25280 ( .B(clk), .A(\g.we_clk [7494]));
Q_ASSIGN U25281 ( .B(clk), .A(\g.we_clk [7493]));
Q_ASSIGN U25282 ( .B(clk), .A(\g.we_clk [7492]));
Q_ASSIGN U25283 ( .B(clk), .A(\g.we_clk [7491]));
Q_ASSIGN U25284 ( .B(clk), .A(\g.we_clk [7490]));
Q_ASSIGN U25285 ( .B(clk), .A(\g.we_clk [7489]));
Q_ASSIGN U25286 ( .B(clk), .A(\g.we_clk [7488]));
Q_ASSIGN U25287 ( .B(clk), .A(\g.we_clk [7487]));
Q_ASSIGN U25288 ( .B(clk), .A(\g.we_clk [7486]));
Q_ASSIGN U25289 ( .B(clk), .A(\g.we_clk [7485]));
Q_ASSIGN U25290 ( .B(clk), .A(\g.we_clk [7484]));
Q_ASSIGN U25291 ( .B(clk), .A(\g.we_clk [7483]));
Q_ASSIGN U25292 ( .B(clk), .A(\g.we_clk [7482]));
Q_ASSIGN U25293 ( .B(clk), .A(\g.we_clk [7481]));
Q_ASSIGN U25294 ( .B(clk), .A(\g.we_clk [7480]));
Q_ASSIGN U25295 ( .B(clk), .A(\g.we_clk [7479]));
Q_ASSIGN U25296 ( .B(clk), .A(\g.we_clk [7478]));
Q_ASSIGN U25297 ( .B(clk), .A(\g.we_clk [7477]));
Q_ASSIGN U25298 ( .B(clk), .A(\g.we_clk [7476]));
Q_ASSIGN U25299 ( .B(clk), .A(\g.we_clk [7475]));
Q_ASSIGN U25300 ( .B(clk), .A(\g.we_clk [7474]));
Q_ASSIGN U25301 ( .B(clk), .A(\g.we_clk [7473]));
Q_ASSIGN U25302 ( .B(clk), .A(\g.we_clk [7472]));
Q_ASSIGN U25303 ( .B(clk), .A(\g.we_clk [7471]));
Q_ASSIGN U25304 ( .B(clk), .A(\g.we_clk [7470]));
Q_ASSIGN U25305 ( .B(clk), .A(\g.we_clk [7469]));
Q_ASSIGN U25306 ( .B(clk), .A(\g.we_clk [7468]));
Q_ASSIGN U25307 ( .B(clk), .A(\g.we_clk [7467]));
Q_ASSIGN U25308 ( .B(clk), .A(\g.we_clk [7466]));
Q_ASSIGN U25309 ( .B(clk), .A(\g.we_clk [7465]));
Q_ASSIGN U25310 ( .B(clk), .A(\g.we_clk [7464]));
Q_ASSIGN U25311 ( .B(clk), .A(\g.we_clk [7463]));
Q_ASSIGN U25312 ( .B(clk), .A(\g.we_clk [7462]));
Q_ASSIGN U25313 ( .B(clk), .A(\g.we_clk [7461]));
Q_ASSIGN U25314 ( .B(clk), .A(\g.we_clk [7460]));
Q_ASSIGN U25315 ( .B(clk), .A(\g.we_clk [7459]));
Q_ASSIGN U25316 ( .B(clk), .A(\g.we_clk [7458]));
Q_ASSIGN U25317 ( .B(clk), .A(\g.we_clk [7457]));
Q_ASSIGN U25318 ( .B(clk), .A(\g.we_clk [7456]));
Q_ASSIGN U25319 ( .B(clk), .A(\g.we_clk [7455]));
Q_ASSIGN U25320 ( .B(clk), .A(\g.we_clk [7454]));
Q_ASSIGN U25321 ( .B(clk), .A(\g.we_clk [7453]));
Q_ASSIGN U25322 ( .B(clk), .A(\g.we_clk [7452]));
Q_ASSIGN U25323 ( .B(clk), .A(\g.we_clk [7451]));
Q_ASSIGN U25324 ( .B(clk), .A(\g.we_clk [7450]));
Q_ASSIGN U25325 ( .B(clk), .A(\g.we_clk [7449]));
Q_ASSIGN U25326 ( .B(clk), .A(\g.we_clk [7448]));
Q_ASSIGN U25327 ( .B(clk), .A(\g.we_clk [7447]));
Q_ASSIGN U25328 ( .B(clk), .A(\g.we_clk [7446]));
Q_ASSIGN U25329 ( .B(clk), .A(\g.we_clk [7445]));
Q_ASSIGN U25330 ( .B(clk), .A(\g.we_clk [7444]));
Q_ASSIGN U25331 ( .B(clk), .A(\g.we_clk [7443]));
Q_ASSIGN U25332 ( .B(clk), .A(\g.we_clk [7442]));
Q_ASSIGN U25333 ( .B(clk), .A(\g.we_clk [7441]));
Q_ASSIGN U25334 ( .B(clk), .A(\g.we_clk [7440]));
Q_ASSIGN U25335 ( .B(clk), .A(\g.we_clk [7439]));
Q_ASSIGN U25336 ( .B(clk), .A(\g.we_clk [7438]));
Q_ASSIGN U25337 ( .B(clk), .A(\g.we_clk [7437]));
Q_ASSIGN U25338 ( .B(clk), .A(\g.we_clk [7436]));
Q_ASSIGN U25339 ( .B(clk), .A(\g.we_clk [7435]));
Q_ASSIGN U25340 ( .B(clk), .A(\g.we_clk [7434]));
Q_ASSIGN U25341 ( .B(clk), .A(\g.we_clk [7433]));
Q_ASSIGN U25342 ( .B(clk), .A(\g.we_clk [7432]));
Q_ASSIGN U25343 ( .B(clk), .A(\g.we_clk [7431]));
Q_ASSIGN U25344 ( .B(clk), .A(\g.we_clk [7430]));
Q_ASSIGN U25345 ( .B(clk), .A(\g.we_clk [7429]));
Q_ASSIGN U25346 ( .B(clk), .A(\g.we_clk [7428]));
Q_ASSIGN U25347 ( .B(clk), .A(\g.we_clk [7427]));
Q_ASSIGN U25348 ( .B(clk), .A(\g.we_clk [7426]));
Q_ASSIGN U25349 ( .B(clk), .A(\g.we_clk [7425]));
Q_ASSIGN U25350 ( .B(clk), .A(\g.we_clk [7424]));
Q_ASSIGN U25351 ( .B(clk), .A(\g.we_clk [7423]));
Q_ASSIGN U25352 ( .B(clk), .A(\g.we_clk [7422]));
Q_ASSIGN U25353 ( .B(clk), .A(\g.we_clk [7421]));
Q_ASSIGN U25354 ( .B(clk), .A(\g.we_clk [7420]));
Q_ASSIGN U25355 ( .B(clk), .A(\g.we_clk [7419]));
Q_ASSIGN U25356 ( .B(clk), .A(\g.we_clk [7418]));
Q_ASSIGN U25357 ( .B(clk), .A(\g.we_clk [7417]));
Q_ASSIGN U25358 ( .B(clk), .A(\g.we_clk [7416]));
Q_ASSIGN U25359 ( .B(clk), .A(\g.we_clk [7415]));
Q_ASSIGN U25360 ( .B(clk), .A(\g.we_clk [7414]));
Q_ASSIGN U25361 ( .B(clk), .A(\g.we_clk [7413]));
Q_ASSIGN U25362 ( .B(clk), .A(\g.we_clk [7412]));
Q_ASSIGN U25363 ( .B(clk), .A(\g.we_clk [7411]));
Q_ASSIGN U25364 ( .B(clk), .A(\g.we_clk [7410]));
Q_ASSIGN U25365 ( .B(clk), .A(\g.we_clk [7409]));
Q_ASSIGN U25366 ( .B(clk), .A(\g.we_clk [7408]));
Q_ASSIGN U25367 ( .B(clk), .A(\g.we_clk [7407]));
Q_ASSIGN U25368 ( .B(clk), .A(\g.we_clk [7406]));
Q_ASSIGN U25369 ( .B(clk), .A(\g.we_clk [7405]));
Q_ASSIGN U25370 ( .B(clk), .A(\g.we_clk [7404]));
Q_ASSIGN U25371 ( .B(clk), .A(\g.we_clk [7403]));
Q_ASSIGN U25372 ( .B(clk), .A(\g.we_clk [7402]));
Q_ASSIGN U25373 ( .B(clk), .A(\g.we_clk [7401]));
Q_ASSIGN U25374 ( .B(clk), .A(\g.we_clk [7400]));
Q_ASSIGN U25375 ( .B(clk), .A(\g.we_clk [7399]));
Q_ASSIGN U25376 ( .B(clk), .A(\g.we_clk [7398]));
Q_ASSIGN U25377 ( .B(clk), .A(\g.we_clk [7397]));
Q_ASSIGN U25378 ( .B(clk), .A(\g.we_clk [7396]));
Q_ASSIGN U25379 ( .B(clk), .A(\g.we_clk [7395]));
Q_ASSIGN U25380 ( .B(clk), .A(\g.we_clk [7394]));
Q_ASSIGN U25381 ( .B(clk), .A(\g.we_clk [7393]));
Q_ASSIGN U25382 ( .B(clk), .A(\g.we_clk [7392]));
Q_ASSIGN U25383 ( .B(clk), .A(\g.we_clk [7391]));
Q_ASSIGN U25384 ( .B(clk), .A(\g.we_clk [7390]));
Q_ASSIGN U25385 ( .B(clk), .A(\g.we_clk [7389]));
Q_ASSIGN U25386 ( .B(clk), .A(\g.we_clk [7388]));
Q_ASSIGN U25387 ( .B(clk), .A(\g.we_clk [7387]));
Q_ASSIGN U25388 ( .B(clk), .A(\g.we_clk [7386]));
Q_ASSIGN U25389 ( .B(clk), .A(\g.we_clk [7385]));
Q_ASSIGN U25390 ( .B(clk), .A(\g.we_clk [7384]));
Q_ASSIGN U25391 ( .B(clk), .A(\g.we_clk [7383]));
Q_ASSIGN U25392 ( .B(clk), .A(\g.we_clk [7382]));
Q_ASSIGN U25393 ( .B(clk), .A(\g.we_clk [7381]));
Q_ASSIGN U25394 ( .B(clk), .A(\g.we_clk [7380]));
Q_ASSIGN U25395 ( .B(clk), .A(\g.we_clk [7379]));
Q_ASSIGN U25396 ( .B(clk), .A(\g.we_clk [7378]));
Q_ASSIGN U25397 ( .B(clk), .A(\g.we_clk [7377]));
Q_ASSIGN U25398 ( .B(clk), .A(\g.we_clk [7376]));
Q_ASSIGN U25399 ( .B(clk), .A(\g.we_clk [7375]));
Q_ASSIGN U25400 ( .B(clk), .A(\g.we_clk [7374]));
Q_ASSIGN U25401 ( .B(clk), .A(\g.we_clk [7373]));
Q_ASSIGN U25402 ( .B(clk), .A(\g.we_clk [7372]));
Q_ASSIGN U25403 ( .B(clk), .A(\g.we_clk [7371]));
Q_ASSIGN U25404 ( .B(clk), .A(\g.we_clk [7370]));
Q_ASSIGN U25405 ( .B(clk), .A(\g.we_clk [7369]));
Q_ASSIGN U25406 ( .B(clk), .A(\g.we_clk [7368]));
Q_ASSIGN U25407 ( .B(clk), .A(\g.we_clk [7367]));
Q_ASSIGN U25408 ( .B(clk), .A(\g.we_clk [7366]));
Q_ASSIGN U25409 ( .B(clk), .A(\g.we_clk [7365]));
Q_ASSIGN U25410 ( .B(clk), .A(\g.we_clk [7364]));
Q_ASSIGN U25411 ( .B(clk), .A(\g.we_clk [7363]));
Q_ASSIGN U25412 ( .B(clk), .A(\g.we_clk [7362]));
Q_ASSIGN U25413 ( .B(clk), .A(\g.we_clk [7361]));
Q_ASSIGN U25414 ( .B(clk), .A(\g.we_clk [7360]));
Q_ASSIGN U25415 ( .B(clk), .A(\g.we_clk [7359]));
Q_ASSIGN U25416 ( .B(clk), .A(\g.we_clk [7358]));
Q_ASSIGN U25417 ( .B(clk), .A(\g.we_clk [7357]));
Q_ASSIGN U25418 ( .B(clk), .A(\g.we_clk [7356]));
Q_ASSIGN U25419 ( .B(clk), .A(\g.we_clk [7355]));
Q_ASSIGN U25420 ( .B(clk), .A(\g.we_clk [7354]));
Q_ASSIGN U25421 ( .B(clk), .A(\g.we_clk [7353]));
Q_ASSIGN U25422 ( .B(clk), .A(\g.we_clk [7352]));
Q_ASSIGN U25423 ( .B(clk), .A(\g.we_clk [7351]));
Q_ASSIGN U25424 ( .B(clk), .A(\g.we_clk [7350]));
Q_ASSIGN U25425 ( .B(clk), .A(\g.we_clk [7349]));
Q_ASSIGN U25426 ( .B(clk), .A(\g.we_clk [7348]));
Q_ASSIGN U25427 ( .B(clk), .A(\g.we_clk [7347]));
Q_ASSIGN U25428 ( .B(clk), .A(\g.we_clk [7346]));
Q_ASSIGN U25429 ( .B(clk), .A(\g.we_clk [7345]));
Q_ASSIGN U25430 ( .B(clk), .A(\g.we_clk [7344]));
Q_ASSIGN U25431 ( .B(clk), .A(\g.we_clk [7343]));
Q_ASSIGN U25432 ( .B(clk), .A(\g.we_clk [7342]));
Q_ASSIGN U25433 ( .B(clk), .A(\g.we_clk [7341]));
Q_ASSIGN U25434 ( .B(clk), .A(\g.we_clk [7340]));
Q_ASSIGN U25435 ( .B(clk), .A(\g.we_clk [7339]));
Q_ASSIGN U25436 ( .B(clk), .A(\g.we_clk [7338]));
Q_ASSIGN U25437 ( .B(clk), .A(\g.we_clk [7337]));
Q_ASSIGN U25438 ( .B(clk), .A(\g.we_clk [7336]));
Q_ASSIGN U25439 ( .B(clk), .A(\g.we_clk [7335]));
Q_ASSIGN U25440 ( .B(clk), .A(\g.we_clk [7334]));
Q_ASSIGN U25441 ( .B(clk), .A(\g.we_clk [7333]));
Q_ASSIGN U25442 ( .B(clk), .A(\g.we_clk [7332]));
Q_ASSIGN U25443 ( .B(clk), .A(\g.we_clk [7331]));
Q_ASSIGN U25444 ( .B(clk), .A(\g.we_clk [7330]));
Q_ASSIGN U25445 ( .B(clk), .A(\g.we_clk [7329]));
Q_ASSIGN U25446 ( .B(clk), .A(\g.we_clk [7328]));
Q_ASSIGN U25447 ( .B(clk), .A(\g.we_clk [7327]));
Q_ASSIGN U25448 ( .B(clk), .A(\g.we_clk [7326]));
Q_ASSIGN U25449 ( .B(clk), .A(\g.we_clk [7325]));
Q_ASSIGN U25450 ( .B(clk), .A(\g.we_clk [7324]));
Q_ASSIGN U25451 ( .B(clk), .A(\g.we_clk [7323]));
Q_ASSIGN U25452 ( .B(clk), .A(\g.we_clk [7322]));
Q_ASSIGN U25453 ( .B(clk), .A(\g.we_clk [7321]));
Q_ASSIGN U25454 ( .B(clk), .A(\g.we_clk [7320]));
Q_ASSIGN U25455 ( .B(clk), .A(\g.we_clk [7319]));
Q_ASSIGN U25456 ( .B(clk), .A(\g.we_clk [7318]));
Q_ASSIGN U25457 ( .B(clk), .A(\g.we_clk [7317]));
Q_ASSIGN U25458 ( .B(clk), .A(\g.we_clk [7316]));
Q_ASSIGN U25459 ( .B(clk), .A(\g.we_clk [7315]));
Q_ASSIGN U25460 ( .B(clk), .A(\g.we_clk [7314]));
Q_ASSIGN U25461 ( .B(clk), .A(\g.we_clk [7313]));
Q_ASSIGN U25462 ( .B(clk), .A(\g.we_clk [7312]));
Q_ASSIGN U25463 ( .B(clk), .A(\g.we_clk [7311]));
Q_ASSIGN U25464 ( .B(clk), .A(\g.we_clk [7310]));
Q_ASSIGN U25465 ( .B(clk), .A(\g.we_clk [7309]));
Q_ASSIGN U25466 ( .B(clk), .A(\g.we_clk [7308]));
Q_ASSIGN U25467 ( .B(clk), .A(\g.we_clk [7307]));
Q_ASSIGN U25468 ( .B(clk), .A(\g.we_clk [7306]));
Q_ASSIGN U25469 ( .B(clk), .A(\g.we_clk [7305]));
Q_ASSIGN U25470 ( .B(clk), .A(\g.we_clk [7304]));
Q_ASSIGN U25471 ( .B(clk), .A(\g.we_clk [7303]));
Q_ASSIGN U25472 ( .B(clk), .A(\g.we_clk [7302]));
Q_ASSIGN U25473 ( .B(clk), .A(\g.we_clk [7301]));
Q_ASSIGN U25474 ( .B(clk), .A(\g.we_clk [7300]));
Q_ASSIGN U25475 ( .B(clk), .A(\g.we_clk [7299]));
Q_ASSIGN U25476 ( .B(clk), .A(\g.we_clk [7298]));
Q_ASSIGN U25477 ( .B(clk), .A(\g.we_clk [7297]));
Q_ASSIGN U25478 ( .B(clk), .A(\g.we_clk [7296]));
Q_ASSIGN U25479 ( .B(clk), .A(\g.we_clk [7295]));
Q_ASSIGN U25480 ( .B(clk), .A(\g.we_clk [7294]));
Q_ASSIGN U25481 ( .B(clk), .A(\g.we_clk [7293]));
Q_ASSIGN U25482 ( .B(clk), .A(\g.we_clk [7292]));
Q_ASSIGN U25483 ( .B(clk), .A(\g.we_clk [7291]));
Q_ASSIGN U25484 ( .B(clk), .A(\g.we_clk [7290]));
Q_ASSIGN U25485 ( .B(clk), .A(\g.we_clk [7289]));
Q_ASSIGN U25486 ( .B(clk), .A(\g.we_clk [7288]));
Q_ASSIGN U25487 ( .B(clk), .A(\g.we_clk [7287]));
Q_ASSIGN U25488 ( .B(clk), .A(\g.we_clk [7286]));
Q_ASSIGN U25489 ( .B(clk), .A(\g.we_clk [7285]));
Q_ASSIGN U25490 ( .B(clk), .A(\g.we_clk [7284]));
Q_ASSIGN U25491 ( .B(clk), .A(\g.we_clk [7283]));
Q_ASSIGN U25492 ( .B(clk), .A(\g.we_clk [7282]));
Q_ASSIGN U25493 ( .B(clk), .A(\g.we_clk [7281]));
Q_ASSIGN U25494 ( .B(clk), .A(\g.we_clk [7280]));
Q_ASSIGN U25495 ( .B(clk), .A(\g.we_clk [7279]));
Q_ASSIGN U25496 ( .B(clk), .A(\g.we_clk [7278]));
Q_ASSIGN U25497 ( .B(clk), .A(\g.we_clk [7277]));
Q_ASSIGN U25498 ( .B(clk), .A(\g.we_clk [7276]));
Q_ASSIGN U25499 ( .B(clk), .A(\g.we_clk [7275]));
Q_ASSIGN U25500 ( .B(clk), .A(\g.we_clk [7274]));
Q_ASSIGN U25501 ( .B(clk), .A(\g.we_clk [7273]));
Q_ASSIGN U25502 ( .B(clk), .A(\g.we_clk [7272]));
Q_ASSIGN U25503 ( .B(clk), .A(\g.we_clk [7271]));
Q_ASSIGN U25504 ( .B(clk), .A(\g.we_clk [7270]));
Q_ASSIGN U25505 ( .B(clk), .A(\g.we_clk [7269]));
Q_ASSIGN U25506 ( .B(clk), .A(\g.we_clk [7268]));
Q_ASSIGN U25507 ( .B(clk), .A(\g.we_clk [7267]));
Q_ASSIGN U25508 ( .B(clk), .A(\g.we_clk [7266]));
Q_ASSIGN U25509 ( .B(clk), .A(\g.we_clk [7265]));
Q_ASSIGN U25510 ( .B(clk), .A(\g.we_clk [7264]));
Q_ASSIGN U25511 ( .B(clk), .A(\g.we_clk [7263]));
Q_ASSIGN U25512 ( .B(clk), .A(\g.we_clk [7262]));
Q_ASSIGN U25513 ( .B(clk), .A(\g.we_clk [7261]));
Q_ASSIGN U25514 ( .B(clk), .A(\g.we_clk [7260]));
Q_ASSIGN U25515 ( .B(clk), .A(\g.we_clk [7259]));
Q_ASSIGN U25516 ( .B(clk), .A(\g.we_clk [7258]));
Q_ASSIGN U25517 ( .B(clk), .A(\g.we_clk [7257]));
Q_ASSIGN U25518 ( .B(clk), .A(\g.we_clk [7256]));
Q_ASSIGN U25519 ( .B(clk), .A(\g.we_clk [7255]));
Q_ASSIGN U25520 ( .B(clk), .A(\g.we_clk [7254]));
Q_ASSIGN U25521 ( .B(clk), .A(\g.we_clk [7253]));
Q_ASSIGN U25522 ( .B(clk), .A(\g.we_clk [7252]));
Q_ASSIGN U25523 ( .B(clk), .A(\g.we_clk [7251]));
Q_ASSIGN U25524 ( .B(clk), .A(\g.we_clk [7250]));
Q_ASSIGN U25525 ( .B(clk), .A(\g.we_clk [7249]));
Q_ASSIGN U25526 ( .B(clk), .A(\g.we_clk [7248]));
Q_ASSIGN U25527 ( .B(clk), .A(\g.we_clk [7247]));
Q_ASSIGN U25528 ( .B(clk), .A(\g.we_clk [7246]));
Q_ASSIGN U25529 ( .B(clk), .A(\g.we_clk [7245]));
Q_ASSIGN U25530 ( .B(clk), .A(\g.we_clk [7244]));
Q_ASSIGN U25531 ( .B(clk), .A(\g.we_clk [7243]));
Q_ASSIGN U25532 ( .B(clk), .A(\g.we_clk [7242]));
Q_ASSIGN U25533 ( .B(clk), .A(\g.we_clk [7241]));
Q_ASSIGN U25534 ( .B(clk), .A(\g.we_clk [7240]));
Q_ASSIGN U25535 ( .B(clk), .A(\g.we_clk [7239]));
Q_ASSIGN U25536 ( .B(clk), .A(\g.we_clk [7238]));
Q_ASSIGN U25537 ( .B(clk), .A(\g.we_clk [7237]));
Q_ASSIGN U25538 ( .B(clk), .A(\g.we_clk [7236]));
Q_ASSIGN U25539 ( .B(clk), .A(\g.we_clk [7235]));
Q_ASSIGN U25540 ( .B(clk), .A(\g.we_clk [7234]));
Q_ASSIGN U25541 ( .B(clk), .A(\g.we_clk [7233]));
Q_ASSIGN U25542 ( .B(clk), .A(\g.we_clk [7232]));
Q_ASSIGN U25543 ( .B(clk), .A(\g.we_clk [7231]));
Q_ASSIGN U25544 ( .B(clk), .A(\g.we_clk [7230]));
Q_ASSIGN U25545 ( .B(clk), .A(\g.we_clk [7229]));
Q_ASSIGN U25546 ( .B(clk), .A(\g.we_clk [7228]));
Q_ASSIGN U25547 ( .B(clk), .A(\g.we_clk [7227]));
Q_ASSIGN U25548 ( .B(clk), .A(\g.we_clk [7226]));
Q_ASSIGN U25549 ( .B(clk), .A(\g.we_clk [7225]));
Q_ASSIGN U25550 ( .B(clk), .A(\g.we_clk [7224]));
Q_ASSIGN U25551 ( .B(clk), .A(\g.we_clk [7223]));
Q_ASSIGN U25552 ( .B(clk), .A(\g.we_clk [7222]));
Q_ASSIGN U25553 ( .B(clk), .A(\g.we_clk [7221]));
Q_ASSIGN U25554 ( .B(clk), .A(\g.we_clk [7220]));
Q_ASSIGN U25555 ( .B(clk), .A(\g.we_clk [7219]));
Q_ASSIGN U25556 ( .B(clk), .A(\g.we_clk [7218]));
Q_ASSIGN U25557 ( .B(clk), .A(\g.we_clk [7217]));
Q_ASSIGN U25558 ( .B(clk), .A(\g.we_clk [7216]));
Q_ASSIGN U25559 ( .B(clk), .A(\g.we_clk [7215]));
Q_ASSIGN U25560 ( .B(clk), .A(\g.we_clk [7214]));
Q_ASSIGN U25561 ( .B(clk), .A(\g.we_clk [7213]));
Q_ASSIGN U25562 ( .B(clk), .A(\g.we_clk [7212]));
Q_ASSIGN U25563 ( .B(clk), .A(\g.we_clk [7211]));
Q_ASSIGN U25564 ( .B(clk), .A(\g.we_clk [7210]));
Q_ASSIGN U25565 ( .B(clk), .A(\g.we_clk [7209]));
Q_ASSIGN U25566 ( .B(clk), .A(\g.we_clk [7208]));
Q_ASSIGN U25567 ( .B(clk), .A(\g.we_clk [7207]));
Q_ASSIGN U25568 ( .B(clk), .A(\g.we_clk [7206]));
Q_ASSIGN U25569 ( .B(clk), .A(\g.we_clk [7205]));
Q_ASSIGN U25570 ( .B(clk), .A(\g.we_clk [7204]));
Q_ASSIGN U25571 ( .B(clk), .A(\g.we_clk [7203]));
Q_ASSIGN U25572 ( .B(clk), .A(\g.we_clk [7202]));
Q_ASSIGN U25573 ( .B(clk), .A(\g.we_clk [7201]));
Q_ASSIGN U25574 ( .B(clk), .A(\g.we_clk [7200]));
Q_ASSIGN U25575 ( .B(clk), .A(\g.we_clk [7199]));
Q_ASSIGN U25576 ( .B(clk), .A(\g.we_clk [7198]));
Q_ASSIGN U25577 ( .B(clk), .A(\g.we_clk [7197]));
Q_ASSIGN U25578 ( .B(clk), .A(\g.we_clk [7196]));
Q_ASSIGN U25579 ( .B(clk), .A(\g.we_clk [7195]));
Q_ASSIGN U25580 ( .B(clk), .A(\g.we_clk [7194]));
Q_ASSIGN U25581 ( .B(clk), .A(\g.we_clk [7193]));
Q_ASSIGN U25582 ( .B(clk), .A(\g.we_clk [7192]));
Q_ASSIGN U25583 ( .B(clk), .A(\g.we_clk [7191]));
Q_ASSIGN U25584 ( .B(clk), .A(\g.we_clk [7190]));
Q_ASSIGN U25585 ( .B(clk), .A(\g.we_clk [7189]));
Q_ASSIGN U25586 ( .B(clk), .A(\g.we_clk [7188]));
Q_ASSIGN U25587 ( .B(clk), .A(\g.we_clk [7187]));
Q_ASSIGN U25588 ( .B(clk), .A(\g.we_clk [7186]));
Q_ASSIGN U25589 ( .B(clk), .A(\g.we_clk [7185]));
Q_ASSIGN U25590 ( .B(clk), .A(\g.we_clk [7184]));
Q_ASSIGN U25591 ( .B(clk), .A(\g.we_clk [7183]));
Q_ASSIGN U25592 ( .B(clk), .A(\g.we_clk [7182]));
Q_ASSIGN U25593 ( .B(clk), .A(\g.we_clk [7181]));
Q_ASSIGN U25594 ( .B(clk), .A(\g.we_clk [7180]));
Q_ASSIGN U25595 ( .B(clk), .A(\g.we_clk [7179]));
Q_ASSIGN U25596 ( .B(clk), .A(\g.we_clk [7178]));
Q_ASSIGN U25597 ( .B(clk), .A(\g.we_clk [7177]));
Q_ASSIGN U25598 ( .B(clk), .A(\g.we_clk [7176]));
Q_ASSIGN U25599 ( .B(clk), .A(\g.we_clk [7175]));
Q_ASSIGN U25600 ( .B(clk), .A(\g.we_clk [7174]));
Q_ASSIGN U25601 ( .B(clk), .A(\g.we_clk [7173]));
Q_ASSIGN U25602 ( .B(clk), .A(\g.we_clk [7172]));
Q_ASSIGN U25603 ( .B(clk), .A(\g.we_clk [7171]));
Q_ASSIGN U25604 ( .B(clk), .A(\g.we_clk [7170]));
Q_ASSIGN U25605 ( .B(clk), .A(\g.we_clk [7169]));
Q_ASSIGN U25606 ( .B(clk), .A(\g.we_clk [7168]));
Q_ASSIGN U25607 ( .B(clk), .A(\g.we_clk [7167]));
Q_ASSIGN U25608 ( .B(clk), .A(\g.we_clk [7166]));
Q_ASSIGN U25609 ( .B(clk), .A(\g.we_clk [7165]));
Q_ASSIGN U25610 ( .B(clk), .A(\g.we_clk [7164]));
Q_ASSIGN U25611 ( .B(clk), .A(\g.we_clk [7163]));
Q_ASSIGN U25612 ( .B(clk), .A(\g.we_clk [7162]));
Q_ASSIGN U25613 ( .B(clk), .A(\g.we_clk [7161]));
Q_ASSIGN U25614 ( .B(clk), .A(\g.we_clk [7160]));
Q_ASSIGN U25615 ( .B(clk), .A(\g.we_clk [7159]));
Q_ASSIGN U25616 ( .B(clk), .A(\g.we_clk [7158]));
Q_ASSIGN U25617 ( .B(clk), .A(\g.we_clk [7157]));
Q_ASSIGN U25618 ( .B(clk), .A(\g.we_clk [7156]));
Q_ASSIGN U25619 ( .B(clk), .A(\g.we_clk [7155]));
Q_ASSIGN U25620 ( .B(clk), .A(\g.we_clk [7154]));
Q_ASSIGN U25621 ( .B(clk), .A(\g.we_clk [7153]));
Q_ASSIGN U25622 ( .B(clk), .A(\g.we_clk [7152]));
Q_ASSIGN U25623 ( .B(clk), .A(\g.we_clk [7151]));
Q_ASSIGN U25624 ( .B(clk), .A(\g.we_clk [7150]));
Q_ASSIGN U25625 ( .B(clk), .A(\g.we_clk [7149]));
Q_ASSIGN U25626 ( .B(clk), .A(\g.we_clk [7148]));
Q_ASSIGN U25627 ( .B(clk), .A(\g.we_clk [7147]));
Q_ASSIGN U25628 ( .B(clk), .A(\g.we_clk [7146]));
Q_ASSIGN U25629 ( .B(clk), .A(\g.we_clk [7145]));
Q_ASSIGN U25630 ( .B(clk), .A(\g.we_clk [7144]));
Q_ASSIGN U25631 ( .B(clk), .A(\g.we_clk [7143]));
Q_ASSIGN U25632 ( .B(clk), .A(\g.we_clk [7142]));
Q_ASSIGN U25633 ( .B(clk), .A(\g.we_clk [7141]));
Q_ASSIGN U25634 ( .B(clk), .A(\g.we_clk [7140]));
Q_ASSIGN U25635 ( .B(clk), .A(\g.we_clk [7139]));
Q_ASSIGN U25636 ( .B(clk), .A(\g.we_clk [7138]));
Q_ASSIGN U25637 ( .B(clk), .A(\g.we_clk [7137]));
Q_ASSIGN U25638 ( .B(clk), .A(\g.we_clk [7136]));
Q_ASSIGN U25639 ( .B(clk), .A(\g.we_clk [7135]));
Q_ASSIGN U25640 ( .B(clk), .A(\g.we_clk [7134]));
Q_ASSIGN U25641 ( .B(clk), .A(\g.we_clk [7133]));
Q_ASSIGN U25642 ( .B(clk), .A(\g.we_clk [7132]));
Q_ASSIGN U25643 ( .B(clk), .A(\g.we_clk [7131]));
Q_ASSIGN U25644 ( .B(clk), .A(\g.we_clk [7130]));
Q_ASSIGN U25645 ( .B(clk), .A(\g.we_clk [7129]));
Q_ASSIGN U25646 ( .B(clk), .A(\g.we_clk [7128]));
Q_ASSIGN U25647 ( .B(clk), .A(\g.we_clk [7127]));
Q_ASSIGN U25648 ( .B(clk), .A(\g.we_clk [7126]));
Q_ASSIGN U25649 ( .B(clk), .A(\g.we_clk [7125]));
Q_ASSIGN U25650 ( .B(clk), .A(\g.we_clk [7124]));
Q_ASSIGN U25651 ( .B(clk), .A(\g.we_clk [7123]));
Q_ASSIGN U25652 ( .B(clk), .A(\g.we_clk [7122]));
Q_ASSIGN U25653 ( .B(clk), .A(\g.we_clk [7121]));
Q_ASSIGN U25654 ( .B(clk), .A(\g.we_clk [7120]));
Q_ASSIGN U25655 ( .B(clk), .A(\g.we_clk [7119]));
Q_ASSIGN U25656 ( .B(clk), .A(\g.we_clk [7118]));
Q_ASSIGN U25657 ( .B(clk), .A(\g.we_clk [7117]));
Q_ASSIGN U25658 ( .B(clk), .A(\g.we_clk [7116]));
Q_ASSIGN U25659 ( .B(clk), .A(\g.we_clk [7115]));
Q_ASSIGN U25660 ( .B(clk), .A(\g.we_clk [7114]));
Q_ASSIGN U25661 ( .B(clk), .A(\g.we_clk [7113]));
Q_ASSIGN U25662 ( .B(clk), .A(\g.we_clk [7112]));
Q_ASSIGN U25663 ( .B(clk), .A(\g.we_clk [7111]));
Q_ASSIGN U25664 ( .B(clk), .A(\g.we_clk [7110]));
Q_ASSIGN U25665 ( .B(clk), .A(\g.we_clk [7109]));
Q_ASSIGN U25666 ( .B(clk), .A(\g.we_clk [7108]));
Q_ASSIGN U25667 ( .B(clk), .A(\g.we_clk [7107]));
Q_ASSIGN U25668 ( .B(clk), .A(\g.we_clk [7106]));
Q_ASSIGN U25669 ( .B(clk), .A(\g.we_clk [7105]));
Q_ASSIGN U25670 ( .B(clk), .A(\g.we_clk [7104]));
Q_ASSIGN U25671 ( .B(clk), .A(\g.we_clk [7103]));
Q_ASSIGN U25672 ( .B(clk), .A(\g.we_clk [7102]));
Q_ASSIGN U25673 ( .B(clk), .A(\g.we_clk [7101]));
Q_ASSIGN U25674 ( .B(clk), .A(\g.we_clk [7100]));
Q_ASSIGN U25675 ( .B(clk), .A(\g.we_clk [7099]));
Q_ASSIGN U25676 ( .B(clk), .A(\g.we_clk [7098]));
Q_ASSIGN U25677 ( .B(clk), .A(\g.we_clk [7097]));
Q_ASSIGN U25678 ( .B(clk), .A(\g.we_clk [7096]));
Q_ASSIGN U25679 ( .B(clk), .A(\g.we_clk [7095]));
Q_ASSIGN U25680 ( .B(clk), .A(\g.we_clk [7094]));
Q_ASSIGN U25681 ( .B(clk), .A(\g.we_clk [7093]));
Q_ASSIGN U25682 ( .B(clk), .A(\g.we_clk [7092]));
Q_ASSIGN U25683 ( .B(clk), .A(\g.we_clk [7091]));
Q_ASSIGN U25684 ( .B(clk), .A(\g.we_clk [7090]));
Q_ASSIGN U25685 ( .B(clk), .A(\g.we_clk [7089]));
Q_ASSIGN U25686 ( .B(clk), .A(\g.we_clk [7088]));
Q_ASSIGN U25687 ( .B(clk), .A(\g.we_clk [7087]));
Q_ASSIGN U25688 ( .B(clk), .A(\g.we_clk [7086]));
Q_ASSIGN U25689 ( .B(clk), .A(\g.we_clk [7085]));
Q_ASSIGN U25690 ( .B(clk), .A(\g.we_clk [7084]));
Q_ASSIGN U25691 ( .B(clk), .A(\g.we_clk [7083]));
Q_ASSIGN U25692 ( .B(clk), .A(\g.we_clk [7082]));
Q_ASSIGN U25693 ( .B(clk), .A(\g.we_clk [7081]));
Q_ASSIGN U25694 ( .B(clk), .A(\g.we_clk [7080]));
Q_ASSIGN U25695 ( .B(clk), .A(\g.we_clk [7079]));
Q_ASSIGN U25696 ( .B(clk), .A(\g.we_clk [7078]));
Q_ASSIGN U25697 ( .B(clk), .A(\g.we_clk [7077]));
Q_ASSIGN U25698 ( .B(clk), .A(\g.we_clk [7076]));
Q_ASSIGN U25699 ( .B(clk), .A(\g.we_clk [7075]));
Q_ASSIGN U25700 ( .B(clk), .A(\g.we_clk [7074]));
Q_ASSIGN U25701 ( .B(clk), .A(\g.we_clk [7073]));
Q_ASSIGN U25702 ( .B(clk), .A(\g.we_clk [7072]));
Q_ASSIGN U25703 ( .B(clk), .A(\g.we_clk [7071]));
Q_ASSIGN U25704 ( .B(clk), .A(\g.we_clk [7070]));
Q_ASSIGN U25705 ( .B(clk), .A(\g.we_clk [7069]));
Q_ASSIGN U25706 ( .B(clk), .A(\g.we_clk [7068]));
Q_ASSIGN U25707 ( .B(clk), .A(\g.we_clk [7067]));
Q_ASSIGN U25708 ( .B(clk), .A(\g.we_clk [7066]));
Q_ASSIGN U25709 ( .B(clk), .A(\g.we_clk [7065]));
Q_ASSIGN U25710 ( .B(clk), .A(\g.we_clk [7064]));
Q_ASSIGN U25711 ( .B(clk), .A(\g.we_clk [7063]));
Q_ASSIGN U25712 ( .B(clk), .A(\g.we_clk [7062]));
Q_ASSIGN U25713 ( .B(clk), .A(\g.we_clk [7061]));
Q_ASSIGN U25714 ( .B(clk), .A(\g.we_clk [7060]));
Q_ASSIGN U25715 ( .B(clk), .A(\g.we_clk [7059]));
Q_ASSIGN U25716 ( .B(clk), .A(\g.we_clk [7058]));
Q_ASSIGN U25717 ( .B(clk), .A(\g.we_clk [7057]));
Q_ASSIGN U25718 ( .B(clk), .A(\g.we_clk [7056]));
Q_ASSIGN U25719 ( .B(clk), .A(\g.we_clk [7055]));
Q_ASSIGN U25720 ( .B(clk), .A(\g.we_clk [7054]));
Q_ASSIGN U25721 ( .B(clk), .A(\g.we_clk [7053]));
Q_ASSIGN U25722 ( .B(clk), .A(\g.we_clk [7052]));
Q_ASSIGN U25723 ( .B(clk), .A(\g.we_clk [7051]));
Q_ASSIGN U25724 ( .B(clk), .A(\g.we_clk [7050]));
Q_ASSIGN U25725 ( .B(clk), .A(\g.we_clk [7049]));
Q_ASSIGN U25726 ( .B(clk), .A(\g.we_clk [7048]));
Q_ASSIGN U25727 ( .B(clk), .A(\g.we_clk [7047]));
Q_ASSIGN U25728 ( .B(clk), .A(\g.we_clk [7046]));
Q_ASSIGN U25729 ( .B(clk), .A(\g.we_clk [7045]));
Q_ASSIGN U25730 ( .B(clk), .A(\g.we_clk [7044]));
Q_ASSIGN U25731 ( .B(clk), .A(\g.we_clk [7043]));
Q_ASSIGN U25732 ( .B(clk), .A(\g.we_clk [7042]));
Q_ASSIGN U25733 ( .B(clk), .A(\g.we_clk [7041]));
Q_ASSIGN U25734 ( .B(clk), .A(\g.we_clk [7040]));
Q_ASSIGN U25735 ( .B(clk), .A(\g.we_clk [7039]));
Q_ASSIGN U25736 ( .B(clk), .A(\g.we_clk [7038]));
Q_ASSIGN U25737 ( .B(clk), .A(\g.we_clk [7037]));
Q_ASSIGN U25738 ( .B(clk), .A(\g.we_clk [7036]));
Q_ASSIGN U25739 ( .B(clk), .A(\g.we_clk [7035]));
Q_ASSIGN U25740 ( .B(clk), .A(\g.we_clk [7034]));
Q_ASSIGN U25741 ( .B(clk), .A(\g.we_clk [7033]));
Q_ASSIGN U25742 ( .B(clk), .A(\g.we_clk [7032]));
Q_ASSIGN U25743 ( .B(clk), .A(\g.we_clk [7031]));
Q_ASSIGN U25744 ( .B(clk), .A(\g.we_clk [7030]));
Q_ASSIGN U25745 ( .B(clk), .A(\g.we_clk [7029]));
Q_ASSIGN U25746 ( .B(clk), .A(\g.we_clk [7028]));
Q_ASSIGN U25747 ( .B(clk), .A(\g.we_clk [7027]));
Q_ASSIGN U25748 ( .B(clk), .A(\g.we_clk [7026]));
Q_ASSIGN U25749 ( .B(clk), .A(\g.we_clk [7025]));
Q_ASSIGN U25750 ( .B(clk), .A(\g.we_clk [7024]));
Q_ASSIGN U25751 ( .B(clk), .A(\g.we_clk [7023]));
Q_ASSIGN U25752 ( .B(clk), .A(\g.we_clk [7022]));
Q_ASSIGN U25753 ( .B(clk), .A(\g.we_clk [7021]));
Q_ASSIGN U25754 ( .B(clk), .A(\g.we_clk [7020]));
Q_ASSIGN U25755 ( .B(clk), .A(\g.we_clk [7019]));
Q_ASSIGN U25756 ( .B(clk), .A(\g.we_clk [7018]));
Q_ASSIGN U25757 ( .B(clk), .A(\g.we_clk [7017]));
Q_ASSIGN U25758 ( .B(clk), .A(\g.we_clk [7016]));
Q_ASSIGN U25759 ( .B(clk), .A(\g.we_clk [7015]));
Q_ASSIGN U25760 ( .B(clk), .A(\g.we_clk [7014]));
Q_ASSIGN U25761 ( .B(clk), .A(\g.we_clk [7013]));
Q_ASSIGN U25762 ( .B(clk), .A(\g.we_clk [7012]));
Q_ASSIGN U25763 ( .B(clk), .A(\g.we_clk [7011]));
Q_ASSIGN U25764 ( .B(clk), .A(\g.we_clk [7010]));
Q_ASSIGN U25765 ( .B(clk), .A(\g.we_clk [7009]));
Q_ASSIGN U25766 ( .B(clk), .A(\g.we_clk [7008]));
Q_ASSIGN U25767 ( .B(clk), .A(\g.we_clk [7007]));
Q_ASSIGN U25768 ( .B(clk), .A(\g.we_clk [7006]));
Q_ASSIGN U25769 ( .B(clk), .A(\g.we_clk [7005]));
Q_ASSIGN U25770 ( .B(clk), .A(\g.we_clk [7004]));
Q_ASSIGN U25771 ( .B(clk), .A(\g.we_clk [7003]));
Q_ASSIGN U25772 ( .B(clk), .A(\g.we_clk [7002]));
Q_ASSIGN U25773 ( .B(clk), .A(\g.we_clk [7001]));
Q_ASSIGN U25774 ( .B(clk), .A(\g.we_clk [7000]));
Q_ASSIGN U25775 ( .B(clk), .A(\g.we_clk [6999]));
Q_ASSIGN U25776 ( .B(clk), .A(\g.we_clk [6998]));
Q_ASSIGN U25777 ( .B(clk), .A(\g.we_clk [6997]));
Q_ASSIGN U25778 ( .B(clk), .A(\g.we_clk [6996]));
Q_ASSIGN U25779 ( .B(clk), .A(\g.we_clk [6995]));
Q_ASSIGN U25780 ( .B(clk), .A(\g.we_clk [6994]));
Q_ASSIGN U25781 ( .B(clk), .A(\g.we_clk [6993]));
Q_ASSIGN U25782 ( .B(clk), .A(\g.we_clk [6992]));
Q_ASSIGN U25783 ( .B(clk), .A(\g.we_clk [6991]));
Q_ASSIGN U25784 ( .B(clk), .A(\g.we_clk [6990]));
Q_ASSIGN U25785 ( .B(clk), .A(\g.we_clk [6989]));
Q_ASSIGN U25786 ( .B(clk), .A(\g.we_clk [6988]));
Q_ASSIGN U25787 ( .B(clk), .A(\g.we_clk [6987]));
Q_ASSIGN U25788 ( .B(clk), .A(\g.we_clk [6986]));
Q_ASSIGN U25789 ( .B(clk), .A(\g.we_clk [6985]));
Q_ASSIGN U25790 ( .B(clk), .A(\g.we_clk [6984]));
Q_ASSIGN U25791 ( .B(clk), .A(\g.we_clk [6983]));
Q_ASSIGN U25792 ( .B(clk), .A(\g.we_clk [6982]));
Q_ASSIGN U25793 ( .B(clk), .A(\g.we_clk [6981]));
Q_ASSIGN U25794 ( .B(clk), .A(\g.we_clk [6980]));
Q_ASSIGN U25795 ( .B(clk), .A(\g.we_clk [6979]));
Q_ASSIGN U25796 ( .B(clk), .A(\g.we_clk [6978]));
Q_ASSIGN U25797 ( .B(clk), .A(\g.we_clk [6977]));
Q_ASSIGN U25798 ( .B(clk), .A(\g.we_clk [6976]));
Q_ASSIGN U25799 ( .B(clk), .A(\g.we_clk [6975]));
Q_ASSIGN U25800 ( .B(clk), .A(\g.we_clk [6974]));
Q_ASSIGN U25801 ( .B(clk), .A(\g.we_clk [6973]));
Q_ASSIGN U25802 ( .B(clk), .A(\g.we_clk [6972]));
Q_ASSIGN U25803 ( .B(clk), .A(\g.we_clk [6971]));
Q_ASSIGN U25804 ( .B(clk), .A(\g.we_clk [6970]));
Q_ASSIGN U25805 ( .B(clk), .A(\g.we_clk [6969]));
Q_ASSIGN U25806 ( .B(clk), .A(\g.we_clk [6968]));
Q_ASSIGN U25807 ( .B(clk), .A(\g.we_clk [6967]));
Q_ASSIGN U25808 ( .B(clk), .A(\g.we_clk [6966]));
Q_ASSIGN U25809 ( .B(clk), .A(\g.we_clk [6965]));
Q_ASSIGN U25810 ( .B(clk), .A(\g.we_clk [6964]));
Q_ASSIGN U25811 ( .B(clk), .A(\g.we_clk [6963]));
Q_ASSIGN U25812 ( .B(clk), .A(\g.we_clk [6962]));
Q_ASSIGN U25813 ( .B(clk), .A(\g.we_clk [6961]));
Q_ASSIGN U25814 ( .B(clk), .A(\g.we_clk [6960]));
Q_ASSIGN U25815 ( .B(clk), .A(\g.we_clk [6959]));
Q_ASSIGN U25816 ( .B(clk), .A(\g.we_clk [6958]));
Q_ASSIGN U25817 ( .B(clk), .A(\g.we_clk [6957]));
Q_ASSIGN U25818 ( .B(clk), .A(\g.we_clk [6956]));
Q_ASSIGN U25819 ( .B(clk), .A(\g.we_clk [6955]));
Q_ASSIGN U25820 ( .B(clk), .A(\g.we_clk [6954]));
Q_ASSIGN U25821 ( .B(clk), .A(\g.we_clk [6953]));
Q_ASSIGN U25822 ( .B(clk), .A(\g.we_clk [6952]));
Q_ASSIGN U25823 ( .B(clk), .A(\g.we_clk [6951]));
Q_ASSIGN U25824 ( .B(clk), .A(\g.we_clk [6950]));
Q_ASSIGN U25825 ( .B(clk), .A(\g.we_clk [6949]));
Q_ASSIGN U25826 ( .B(clk), .A(\g.we_clk [6948]));
Q_ASSIGN U25827 ( .B(clk), .A(\g.we_clk [6947]));
Q_ASSIGN U25828 ( .B(clk), .A(\g.we_clk [6946]));
Q_ASSIGN U25829 ( .B(clk), .A(\g.we_clk [6945]));
Q_ASSIGN U25830 ( .B(clk), .A(\g.we_clk [6944]));
Q_ASSIGN U25831 ( .B(clk), .A(\g.we_clk [6943]));
Q_ASSIGN U25832 ( .B(clk), .A(\g.we_clk [6942]));
Q_ASSIGN U25833 ( .B(clk), .A(\g.we_clk [6941]));
Q_ASSIGN U25834 ( .B(clk), .A(\g.we_clk [6940]));
Q_ASSIGN U25835 ( .B(clk), .A(\g.we_clk [6939]));
Q_ASSIGN U25836 ( .B(clk), .A(\g.we_clk [6938]));
Q_ASSIGN U25837 ( .B(clk), .A(\g.we_clk [6937]));
Q_ASSIGN U25838 ( .B(clk), .A(\g.we_clk [6936]));
Q_ASSIGN U25839 ( .B(clk), .A(\g.we_clk [6935]));
Q_ASSIGN U25840 ( .B(clk), .A(\g.we_clk [6934]));
Q_ASSIGN U25841 ( .B(clk), .A(\g.we_clk [6933]));
Q_ASSIGN U25842 ( .B(clk), .A(\g.we_clk [6932]));
Q_ASSIGN U25843 ( .B(clk), .A(\g.we_clk [6931]));
Q_ASSIGN U25844 ( .B(clk), .A(\g.we_clk [6930]));
Q_ASSIGN U25845 ( .B(clk), .A(\g.we_clk [6929]));
Q_ASSIGN U25846 ( .B(clk), .A(\g.we_clk [6928]));
Q_ASSIGN U25847 ( .B(clk), .A(\g.we_clk [6927]));
Q_ASSIGN U25848 ( .B(clk), .A(\g.we_clk [6926]));
Q_ASSIGN U25849 ( .B(clk), .A(\g.we_clk [6925]));
Q_ASSIGN U25850 ( .B(clk), .A(\g.we_clk [6924]));
Q_ASSIGN U25851 ( .B(clk), .A(\g.we_clk [6923]));
Q_ASSIGN U25852 ( .B(clk), .A(\g.we_clk [6922]));
Q_ASSIGN U25853 ( .B(clk), .A(\g.we_clk [6921]));
Q_ASSIGN U25854 ( .B(clk), .A(\g.we_clk [6920]));
Q_ASSIGN U25855 ( .B(clk), .A(\g.we_clk [6919]));
Q_ASSIGN U25856 ( .B(clk), .A(\g.we_clk [6918]));
Q_ASSIGN U25857 ( .B(clk), .A(\g.we_clk [6917]));
Q_ASSIGN U25858 ( .B(clk), .A(\g.we_clk [6916]));
Q_ASSIGN U25859 ( .B(clk), .A(\g.we_clk [6915]));
Q_ASSIGN U25860 ( .B(clk), .A(\g.we_clk [6914]));
Q_ASSIGN U25861 ( .B(clk), .A(\g.we_clk [6913]));
Q_ASSIGN U25862 ( .B(clk), .A(\g.we_clk [6912]));
Q_ASSIGN U25863 ( .B(clk), .A(\g.we_clk [6911]));
Q_ASSIGN U25864 ( .B(clk), .A(\g.we_clk [6910]));
Q_ASSIGN U25865 ( .B(clk), .A(\g.we_clk [6909]));
Q_ASSIGN U25866 ( .B(clk), .A(\g.we_clk [6908]));
Q_ASSIGN U25867 ( .B(clk), .A(\g.we_clk [6907]));
Q_ASSIGN U25868 ( .B(clk), .A(\g.we_clk [6906]));
Q_ASSIGN U25869 ( .B(clk), .A(\g.we_clk [6905]));
Q_ASSIGN U25870 ( .B(clk), .A(\g.we_clk [6904]));
Q_ASSIGN U25871 ( .B(clk), .A(\g.we_clk [6903]));
Q_ASSIGN U25872 ( .B(clk), .A(\g.we_clk [6902]));
Q_ASSIGN U25873 ( .B(clk), .A(\g.we_clk [6901]));
Q_ASSIGN U25874 ( .B(clk), .A(\g.we_clk [6900]));
Q_ASSIGN U25875 ( .B(clk), .A(\g.we_clk [6899]));
Q_ASSIGN U25876 ( .B(clk), .A(\g.we_clk [6898]));
Q_ASSIGN U25877 ( .B(clk), .A(\g.we_clk [6897]));
Q_ASSIGN U25878 ( .B(clk), .A(\g.we_clk [6896]));
Q_ASSIGN U25879 ( .B(clk), .A(\g.we_clk [6895]));
Q_ASSIGN U25880 ( .B(clk), .A(\g.we_clk [6894]));
Q_ASSIGN U25881 ( .B(clk), .A(\g.we_clk [6893]));
Q_ASSIGN U25882 ( .B(clk), .A(\g.we_clk [6892]));
Q_ASSIGN U25883 ( .B(clk), .A(\g.we_clk [6891]));
Q_ASSIGN U25884 ( .B(clk), .A(\g.we_clk [6890]));
Q_ASSIGN U25885 ( .B(clk), .A(\g.we_clk [6889]));
Q_ASSIGN U25886 ( .B(clk), .A(\g.we_clk [6888]));
Q_ASSIGN U25887 ( .B(clk), .A(\g.we_clk [6887]));
Q_ASSIGN U25888 ( .B(clk), .A(\g.we_clk [6886]));
Q_ASSIGN U25889 ( .B(clk), .A(\g.we_clk [6885]));
Q_ASSIGN U25890 ( .B(clk), .A(\g.we_clk [6884]));
Q_ASSIGN U25891 ( .B(clk), .A(\g.we_clk [6883]));
Q_ASSIGN U25892 ( .B(clk), .A(\g.we_clk [6882]));
Q_ASSIGN U25893 ( .B(clk), .A(\g.we_clk [6881]));
Q_ASSIGN U25894 ( .B(clk), .A(\g.we_clk [6880]));
Q_ASSIGN U25895 ( .B(clk), .A(\g.we_clk [6879]));
Q_ASSIGN U25896 ( .B(clk), .A(\g.we_clk [6878]));
Q_ASSIGN U25897 ( .B(clk), .A(\g.we_clk [6877]));
Q_ASSIGN U25898 ( .B(clk), .A(\g.we_clk [6876]));
Q_ASSIGN U25899 ( .B(clk), .A(\g.we_clk [6875]));
Q_ASSIGN U25900 ( .B(clk), .A(\g.we_clk [6874]));
Q_ASSIGN U25901 ( .B(clk), .A(\g.we_clk [6873]));
Q_ASSIGN U25902 ( .B(clk), .A(\g.we_clk [6872]));
Q_ASSIGN U25903 ( .B(clk), .A(\g.we_clk [6871]));
Q_ASSIGN U25904 ( .B(clk), .A(\g.we_clk [6870]));
Q_ASSIGN U25905 ( .B(clk), .A(\g.we_clk [6869]));
Q_ASSIGN U25906 ( .B(clk), .A(\g.we_clk [6868]));
Q_ASSIGN U25907 ( .B(clk), .A(\g.we_clk [6867]));
Q_ASSIGN U25908 ( .B(clk), .A(\g.we_clk [6866]));
Q_ASSIGN U25909 ( .B(clk), .A(\g.we_clk [6865]));
Q_ASSIGN U25910 ( .B(clk), .A(\g.we_clk [6864]));
Q_ASSIGN U25911 ( .B(clk), .A(\g.we_clk [6863]));
Q_ASSIGN U25912 ( .B(clk), .A(\g.we_clk [6862]));
Q_ASSIGN U25913 ( .B(clk), .A(\g.we_clk [6861]));
Q_ASSIGN U25914 ( .B(clk), .A(\g.we_clk [6860]));
Q_ASSIGN U25915 ( .B(clk), .A(\g.we_clk [6859]));
Q_ASSIGN U25916 ( .B(clk), .A(\g.we_clk [6858]));
Q_ASSIGN U25917 ( .B(clk), .A(\g.we_clk [6857]));
Q_ASSIGN U25918 ( .B(clk), .A(\g.we_clk [6856]));
Q_ASSIGN U25919 ( .B(clk), .A(\g.we_clk [6855]));
Q_ASSIGN U25920 ( .B(clk), .A(\g.we_clk [6854]));
Q_ASSIGN U25921 ( .B(clk), .A(\g.we_clk [6853]));
Q_ASSIGN U25922 ( .B(clk), .A(\g.we_clk [6852]));
Q_ASSIGN U25923 ( .B(clk), .A(\g.we_clk [6851]));
Q_ASSIGN U25924 ( .B(clk), .A(\g.we_clk [6850]));
Q_ASSIGN U25925 ( .B(clk), .A(\g.we_clk [6849]));
Q_ASSIGN U25926 ( .B(clk), .A(\g.we_clk [6848]));
Q_ASSIGN U25927 ( .B(clk), .A(\g.we_clk [6847]));
Q_ASSIGN U25928 ( .B(clk), .A(\g.we_clk [6846]));
Q_ASSIGN U25929 ( .B(clk), .A(\g.we_clk [6845]));
Q_ASSIGN U25930 ( .B(clk), .A(\g.we_clk [6844]));
Q_ASSIGN U25931 ( .B(clk), .A(\g.we_clk [6843]));
Q_ASSIGN U25932 ( .B(clk), .A(\g.we_clk [6842]));
Q_ASSIGN U25933 ( .B(clk), .A(\g.we_clk [6841]));
Q_ASSIGN U25934 ( .B(clk), .A(\g.we_clk [6840]));
Q_ASSIGN U25935 ( .B(clk), .A(\g.we_clk [6839]));
Q_ASSIGN U25936 ( .B(clk), .A(\g.we_clk [6838]));
Q_ASSIGN U25937 ( .B(clk), .A(\g.we_clk [6837]));
Q_ASSIGN U25938 ( .B(clk), .A(\g.we_clk [6836]));
Q_ASSIGN U25939 ( .B(clk), .A(\g.we_clk [6835]));
Q_ASSIGN U25940 ( .B(clk), .A(\g.we_clk [6834]));
Q_ASSIGN U25941 ( .B(clk), .A(\g.we_clk [6833]));
Q_ASSIGN U25942 ( .B(clk), .A(\g.we_clk [6832]));
Q_ASSIGN U25943 ( .B(clk), .A(\g.we_clk [6831]));
Q_ASSIGN U25944 ( .B(clk), .A(\g.we_clk [6830]));
Q_ASSIGN U25945 ( .B(clk), .A(\g.we_clk [6829]));
Q_ASSIGN U25946 ( .B(clk), .A(\g.we_clk [6828]));
Q_ASSIGN U25947 ( .B(clk), .A(\g.we_clk [6827]));
Q_ASSIGN U25948 ( .B(clk), .A(\g.we_clk [6826]));
Q_ASSIGN U25949 ( .B(clk), .A(\g.we_clk [6825]));
Q_ASSIGN U25950 ( .B(clk), .A(\g.we_clk [6824]));
Q_ASSIGN U25951 ( .B(clk), .A(\g.we_clk [6823]));
Q_ASSIGN U25952 ( .B(clk), .A(\g.we_clk [6822]));
Q_ASSIGN U25953 ( .B(clk), .A(\g.we_clk [6821]));
Q_ASSIGN U25954 ( .B(clk), .A(\g.we_clk [6820]));
Q_ASSIGN U25955 ( .B(clk), .A(\g.we_clk [6819]));
Q_ASSIGN U25956 ( .B(clk), .A(\g.we_clk [6818]));
Q_ASSIGN U25957 ( .B(clk), .A(\g.we_clk [6817]));
Q_ASSIGN U25958 ( .B(clk), .A(\g.we_clk [6816]));
Q_ASSIGN U25959 ( .B(clk), .A(\g.we_clk [6815]));
Q_ASSIGN U25960 ( .B(clk), .A(\g.we_clk [6814]));
Q_ASSIGN U25961 ( .B(clk), .A(\g.we_clk [6813]));
Q_ASSIGN U25962 ( .B(clk), .A(\g.we_clk [6812]));
Q_ASSIGN U25963 ( .B(clk), .A(\g.we_clk [6811]));
Q_ASSIGN U25964 ( .B(clk), .A(\g.we_clk [6810]));
Q_ASSIGN U25965 ( .B(clk), .A(\g.we_clk [6809]));
Q_ASSIGN U25966 ( .B(clk), .A(\g.we_clk [6808]));
Q_ASSIGN U25967 ( .B(clk), .A(\g.we_clk [6807]));
Q_ASSIGN U25968 ( .B(clk), .A(\g.we_clk [6806]));
Q_ASSIGN U25969 ( .B(clk), .A(\g.we_clk [6805]));
Q_ASSIGN U25970 ( .B(clk), .A(\g.we_clk [6804]));
Q_ASSIGN U25971 ( .B(clk), .A(\g.we_clk [6803]));
Q_ASSIGN U25972 ( .B(clk), .A(\g.we_clk [6802]));
Q_ASSIGN U25973 ( .B(clk), .A(\g.we_clk [6801]));
Q_ASSIGN U25974 ( .B(clk), .A(\g.we_clk [6800]));
Q_ASSIGN U25975 ( .B(clk), .A(\g.we_clk [6799]));
Q_ASSIGN U25976 ( .B(clk), .A(\g.we_clk [6798]));
Q_ASSIGN U25977 ( .B(clk), .A(\g.we_clk [6797]));
Q_ASSIGN U25978 ( .B(clk), .A(\g.we_clk [6796]));
Q_ASSIGN U25979 ( .B(clk), .A(\g.we_clk [6795]));
Q_ASSIGN U25980 ( .B(clk), .A(\g.we_clk [6794]));
Q_ASSIGN U25981 ( .B(clk), .A(\g.we_clk [6793]));
Q_ASSIGN U25982 ( .B(clk), .A(\g.we_clk [6792]));
Q_ASSIGN U25983 ( .B(clk), .A(\g.we_clk [6791]));
Q_ASSIGN U25984 ( .B(clk), .A(\g.we_clk [6790]));
Q_ASSIGN U25985 ( .B(clk), .A(\g.we_clk [6789]));
Q_ASSIGN U25986 ( .B(clk), .A(\g.we_clk [6788]));
Q_ASSIGN U25987 ( .B(clk), .A(\g.we_clk [6787]));
Q_ASSIGN U25988 ( .B(clk), .A(\g.we_clk [6786]));
Q_ASSIGN U25989 ( .B(clk), .A(\g.we_clk [6785]));
Q_ASSIGN U25990 ( .B(clk), .A(\g.we_clk [6784]));
Q_ASSIGN U25991 ( .B(clk), .A(\g.we_clk [6783]));
Q_ASSIGN U25992 ( .B(clk), .A(\g.we_clk [6782]));
Q_ASSIGN U25993 ( .B(clk), .A(\g.we_clk [6781]));
Q_ASSIGN U25994 ( .B(clk), .A(\g.we_clk [6780]));
Q_ASSIGN U25995 ( .B(clk), .A(\g.we_clk [6779]));
Q_ASSIGN U25996 ( .B(clk), .A(\g.we_clk [6778]));
Q_ASSIGN U25997 ( .B(clk), .A(\g.we_clk [6777]));
Q_ASSIGN U25998 ( .B(clk), .A(\g.we_clk [6776]));
Q_ASSIGN U25999 ( .B(clk), .A(\g.we_clk [6775]));
Q_ASSIGN U26000 ( .B(clk), .A(\g.we_clk [6774]));
Q_ASSIGN U26001 ( .B(clk), .A(\g.we_clk [6773]));
Q_ASSIGN U26002 ( .B(clk), .A(\g.we_clk [6772]));
Q_ASSIGN U26003 ( .B(clk), .A(\g.we_clk [6771]));
Q_ASSIGN U26004 ( .B(clk), .A(\g.we_clk [6770]));
Q_ASSIGN U26005 ( .B(clk), .A(\g.we_clk [6769]));
Q_ASSIGN U26006 ( .B(clk), .A(\g.we_clk [6768]));
Q_ASSIGN U26007 ( .B(clk), .A(\g.we_clk [6767]));
Q_ASSIGN U26008 ( .B(clk), .A(\g.we_clk [6766]));
Q_ASSIGN U26009 ( .B(clk), .A(\g.we_clk [6765]));
Q_ASSIGN U26010 ( .B(clk), .A(\g.we_clk [6764]));
Q_ASSIGN U26011 ( .B(clk), .A(\g.we_clk [6763]));
Q_ASSIGN U26012 ( .B(clk), .A(\g.we_clk [6762]));
Q_ASSIGN U26013 ( .B(clk), .A(\g.we_clk [6761]));
Q_ASSIGN U26014 ( .B(clk), .A(\g.we_clk [6760]));
Q_ASSIGN U26015 ( .B(clk), .A(\g.we_clk [6759]));
Q_ASSIGN U26016 ( .B(clk), .A(\g.we_clk [6758]));
Q_ASSIGN U26017 ( .B(clk), .A(\g.we_clk [6757]));
Q_ASSIGN U26018 ( .B(clk), .A(\g.we_clk [6756]));
Q_ASSIGN U26019 ( .B(clk), .A(\g.we_clk [6755]));
Q_ASSIGN U26020 ( .B(clk), .A(\g.we_clk [6754]));
Q_ASSIGN U26021 ( .B(clk), .A(\g.we_clk [6753]));
Q_ASSIGN U26022 ( .B(clk), .A(\g.we_clk [6752]));
Q_ASSIGN U26023 ( .B(clk), .A(\g.we_clk [6751]));
Q_ASSIGN U26024 ( .B(clk), .A(\g.we_clk [6750]));
Q_ASSIGN U26025 ( .B(clk), .A(\g.we_clk [6749]));
Q_ASSIGN U26026 ( .B(clk), .A(\g.we_clk [6748]));
Q_ASSIGN U26027 ( .B(clk), .A(\g.we_clk [6747]));
Q_ASSIGN U26028 ( .B(clk), .A(\g.we_clk [6746]));
Q_ASSIGN U26029 ( .B(clk), .A(\g.we_clk [6745]));
Q_ASSIGN U26030 ( .B(clk), .A(\g.we_clk [6744]));
Q_ASSIGN U26031 ( .B(clk), .A(\g.we_clk [6743]));
Q_ASSIGN U26032 ( .B(clk), .A(\g.we_clk [6742]));
Q_ASSIGN U26033 ( .B(clk), .A(\g.we_clk [6741]));
Q_ASSIGN U26034 ( .B(clk), .A(\g.we_clk [6740]));
Q_ASSIGN U26035 ( .B(clk), .A(\g.we_clk [6739]));
Q_ASSIGN U26036 ( .B(clk), .A(\g.we_clk [6738]));
Q_ASSIGN U26037 ( .B(clk), .A(\g.we_clk [6737]));
Q_ASSIGN U26038 ( .B(clk), .A(\g.we_clk [6736]));
Q_ASSIGN U26039 ( .B(clk), .A(\g.we_clk [6735]));
Q_ASSIGN U26040 ( .B(clk), .A(\g.we_clk [6734]));
Q_ASSIGN U26041 ( .B(clk), .A(\g.we_clk [6733]));
Q_ASSIGN U26042 ( .B(clk), .A(\g.we_clk [6732]));
Q_ASSIGN U26043 ( .B(clk), .A(\g.we_clk [6731]));
Q_ASSIGN U26044 ( .B(clk), .A(\g.we_clk [6730]));
Q_ASSIGN U26045 ( .B(clk), .A(\g.we_clk [6729]));
Q_ASSIGN U26046 ( .B(clk), .A(\g.we_clk [6728]));
Q_ASSIGN U26047 ( .B(clk), .A(\g.we_clk [6727]));
Q_ASSIGN U26048 ( .B(clk), .A(\g.we_clk [6726]));
Q_ASSIGN U26049 ( .B(clk), .A(\g.we_clk [6725]));
Q_ASSIGN U26050 ( .B(clk), .A(\g.we_clk [6724]));
Q_ASSIGN U26051 ( .B(clk), .A(\g.we_clk [6723]));
Q_ASSIGN U26052 ( .B(clk), .A(\g.we_clk [6722]));
Q_ASSIGN U26053 ( .B(clk), .A(\g.we_clk [6721]));
Q_ASSIGN U26054 ( .B(clk), .A(\g.we_clk [6720]));
Q_ASSIGN U26055 ( .B(clk), .A(\g.we_clk [6719]));
Q_ASSIGN U26056 ( .B(clk), .A(\g.we_clk [6718]));
Q_ASSIGN U26057 ( .B(clk), .A(\g.we_clk [6717]));
Q_ASSIGN U26058 ( .B(clk), .A(\g.we_clk [6716]));
Q_ASSIGN U26059 ( .B(clk), .A(\g.we_clk [6715]));
Q_ASSIGN U26060 ( .B(clk), .A(\g.we_clk [6714]));
Q_ASSIGN U26061 ( .B(clk), .A(\g.we_clk [6713]));
Q_ASSIGN U26062 ( .B(clk), .A(\g.we_clk [6712]));
Q_ASSIGN U26063 ( .B(clk), .A(\g.we_clk [6711]));
Q_ASSIGN U26064 ( .B(clk), .A(\g.we_clk [6710]));
Q_ASSIGN U26065 ( .B(clk), .A(\g.we_clk [6709]));
Q_ASSIGN U26066 ( .B(clk), .A(\g.we_clk [6708]));
Q_ASSIGN U26067 ( .B(clk), .A(\g.we_clk [6707]));
Q_ASSIGN U26068 ( .B(clk), .A(\g.we_clk [6706]));
Q_ASSIGN U26069 ( .B(clk), .A(\g.we_clk [6705]));
Q_ASSIGN U26070 ( .B(clk), .A(\g.we_clk [6704]));
Q_ASSIGN U26071 ( .B(clk), .A(\g.we_clk [6703]));
Q_ASSIGN U26072 ( .B(clk), .A(\g.we_clk [6702]));
Q_ASSIGN U26073 ( .B(clk), .A(\g.we_clk [6701]));
Q_ASSIGN U26074 ( .B(clk), .A(\g.we_clk [6700]));
Q_ASSIGN U26075 ( .B(clk), .A(\g.we_clk [6699]));
Q_ASSIGN U26076 ( .B(clk), .A(\g.we_clk [6698]));
Q_ASSIGN U26077 ( .B(clk), .A(\g.we_clk [6697]));
Q_ASSIGN U26078 ( .B(clk), .A(\g.we_clk [6696]));
Q_ASSIGN U26079 ( .B(clk), .A(\g.we_clk [6695]));
Q_ASSIGN U26080 ( .B(clk), .A(\g.we_clk [6694]));
Q_ASSIGN U26081 ( .B(clk), .A(\g.we_clk [6693]));
Q_ASSIGN U26082 ( .B(clk), .A(\g.we_clk [6692]));
Q_ASSIGN U26083 ( .B(clk), .A(\g.we_clk [6691]));
Q_ASSIGN U26084 ( .B(clk), .A(\g.we_clk [6690]));
Q_ASSIGN U26085 ( .B(clk), .A(\g.we_clk [6689]));
Q_ASSIGN U26086 ( .B(clk), .A(\g.we_clk [6688]));
Q_ASSIGN U26087 ( .B(clk), .A(\g.we_clk [6687]));
Q_ASSIGN U26088 ( .B(clk), .A(\g.we_clk [6686]));
Q_ASSIGN U26089 ( .B(clk), .A(\g.we_clk [6685]));
Q_ASSIGN U26090 ( .B(clk), .A(\g.we_clk [6684]));
Q_ASSIGN U26091 ( .B(clk), .A(\g.we_clk [6683]));
Q_ASSIGN U26092 ( .B(clk), .A(\g.we_clk [6682]));
Q_ASSIGN U26093 ( .B(clk), .A(\g.we_clk [6681]));
Q_ASSIGN U26094 ( .B(clk), .A(\g.we_clk [6680]));
Q_ASSIGN U26095 ( .B(clk), .A(\g.we_clk [6679]));
Q_ASSIGN U26096 ( .B(clk), .A(\g.we_clk [6678]));
Q_ASSIGN U26097 ( .B(clk), .A(\g.we_clk [6677]));
Q_ASSIGN U26098 ( .B(clk), .A(\g.we_clk [6676]));
Q_ASSIGN U26099 ( .B(clk), .A(\g.we_clk [6675]));
Q_ASSIGN U26100 ( .B(clk), .A(\g.we_clk [6674]));
Q_ASSIGN U26101 ( .B(clk), .A(\g.we_clk [6673]));
Q_ASSIGN U26102 ( .B(clk), .A(\g.we_clk [6672]));
Q_ASSIGN U26103 ( .B(clk), .A(\g.we_clk [6671]));
Q_ASSIGN U26104 ( .B(clk), .A(\g.we_clk [6670]));
Q_ASSIGN U26105 ( .B(clk), .A(\g.we_clk [6669]));
Q_ASSIGN U26106 ( .B(clk), .A(\g.we_clk [6668]));
Q_ASSIGN U26107 ( .B(clk), .A(\g.we_clk [6667]));
Q_ASSIGN U26108 ( .B(clk), .A(\g.we_clk [6666]));
Q_ASSIGN U26109 ( .B(clk), .A(\g.we_clk [6665]));
Q_ASSIGN U26110 ( .B(clk), .A(\g.we_clk [6664]));
Q_ASSIGN U26111 ( .B(clk), .A(\g.we_clk [6663]));
Q_ASSIGN U26112 ( .B(clk), .A(\g.we_clk [6662]));
Q_ASSIGN U26113 ( .B(clk), .A(\g.we_clk [6661]));
Q_ASSIGN U26114 ( .B(clk), .A(\g.we_clk [6660]));
Q_ASSIGN U26115 ( .B(clk), .A(\g.we_clk [6659]));
Q_ASSIGN U26116 ( .B(clk), .A(\g.we_clk [6658]));
Q_ASSIGN U26117 ( .B(clk), .A(\g.we_clk [6657]));
Q_ASSIGN U26118 ( .B(clk), .A(\g.we_clk [6656]));
Q_ASSIGN U26119 ( .B(clk), .A(\g.we_clk [6655]));
Q_ASSIGN U26120 ( .B(clk), .A(\g.we_clk [6654]));
Q_ASSIGN U26121 ( .B(clk), .A(\g.we_clk [6653]));
Q_ASSIGN U26122 ( .B(clk), .A(\g.we_clk [6652]));
Q_ASSIGN U26123 ( .B(clk), .A(\g.we_clk [6651]));
Q_ASSIGN U26124 ( .B(clk), .A(\g.we_clk [6650]));
Q_ASSIGN U26125 ( .B(clk), .A(\g.we_clk [6649]));
Q_ASSIGN U26126 ( .B(clk), .A(\g.we_clk [6648]));
Q_ASSIGN U26127 ( .B(clk), .A(\g.we_clk [6647]));
Q_ASSIGN U26128 ( .B(clk), .A(\g.we_clk [6646]));
Q_ASSIGN U26129 ( .B(clk), .A(\g.we_clk [6645]));
Q_ASSIGN U26130 ( .B(clk), .A(\g.we_clk [6644]));
Q_ASSIGN U26131 ( .B(clk), .A(\g.we_clk [6643]));
Q_ASSIGN U26132 ( .B(clk), .A(\g.we_clk [6642]));
Q_ASSIGN U26133 ( .B(clk), .A(\g.we_clk [6641]));
Q_ASSIGN U26134 ( .B(clk), .A(\g.we_clk [6640]));
Q_ASSIGN U26135 ( .B(clk), .A(\g.we_clk [6639]));
Q_ASSIGN U26136 ( .B(clk), .A(\g.we_clk [6638]));
Q_ASSIGN U26137 ( .B(clk), .A(\g.we_clk [6637]));
Q_ASSIGN U26138 ( .B(clk), .A(\g.we_clk [6636]));
Q_ASSIGN U26139 ( .B(clk), .A(\g.we_clk [6635]));
Q_ASSIGN U26140 ( .B(clk), .A(\g.we_clk [6634]));
Q_ASSIGN U26141 ( .B(clk), .A(\g.we_clk [6633]));
Q_ASSIGN U26142 ( .B(clk), .A(\g.we_clk [6632]));
Q_ASSIGN U26143 ( .B(clk), .A(\g.we_clk [6631]));
Q_ASSIGN U26144 ( .B(clk), .A(\g.we_clk [6630]));
Q_ASSIGN U26145 ( .B(clk), .A(\g.we_clk [6629]));
Q_ASSIGN U26146 ( .B(clk), .A(\g.we_clk [6628]));
Q_ASSIGN U26147 ( .B(clk), .A(\g.we_clk [6627]));
Q_ASSIGN U26148 ( .B(clk), .A(\g.we_clk [6626]));
Q_ASSIGN U26149 ( .B(clk), .A(\g.we_clk [6625]));
Q_ASSIGN U26150 ( .B(clk), .A(\g.we_clk [6624]));
Q_ASSIGN U26151 ( .B(clk), .A(\g.we_clk [6623]));
Q_ASSIGN U26152 ( .B(clk), .A(\g.we_clk [6622]));
Q_ASSIGN U26153 ( .B(clk), .A(\g.we_clk [6621]));
Q_ASSIGN U26154 ( .B(clk), .A(\g.we_clk [6620]));
Q_ASSIGN U26155 ( .B(clk), .A(\g.we_clk [6619]));
Q_ASSIGN U26156 ( .B(clk), .A(\g.we_clk [6618]));
Q_ASSIGN U26157 ( .B(clk), .A(\g.we_clk [6617]));
Q_ASSIGN U26158 ( .B(clk), .A(\g.we_clk [6616]));
Q_ASSIGN U26159 ( .B(clk), .A(\g.we_clk [6615]));
Q_ASSIGN U26160 ( .B(clk), .A(\g.we_clk [6614]));
Q_ASSIGN U26161 ( .B(clk), .A(\g.we_clk [6613]));
Q_ASSIGN U26162 ( .B(clk), .A(\g.we_clk [6612]));
Q_ASSIGN U26163 ( .B(clk), .A(\g.we_clk [6611]));
Q_ASSIGN U26164 ( .B(clk), .A(\g.we_clk [6610]));
Q_ASSIGN U26165 ( .B(clk), .A(\g.we_clk [6609]));
Q_ASSIGN U26166 ( .B(clk), .A(\g.we_clk [6608]));
Q_ASSIGN U26167 ( .B(clk), .A(\g.we_clk [6607]));
Q_ASSIGN U26168 ( .B(clk), .A(\g.we_clk [6606]));
Q_ASSIGN U26169 ( .B(clk), .A(\g.we_clk [6605]));
Q_ASSIGN U26170 ( .B(clk), .A(\g.we_clk [6604]));
Q_ASSIGN U26171 ( .B(clk), .A(\g.we_clk [6603]));
Q_ASSIGN U26172 ( .B(clk), .A(\g.we_clk [6602]));
Q_ASSIGN U26173 ( .B(clk), .A(\g.we_clk [6601]));
Q_ASSIGN U26174 ( .B(clk), .A(\g.we_clk [6600]));
Q_ASSIGN U26175 ( .B(clk), .A(\g.we_clk [6599]));
Q_ASSIGN U26176 ( .B(clk), .A(\g.we_clk [6598]));
Q_ASSIGN U26177 ( .B(clk), .A(\g.we_clk [6597]));
Q_ASSIGN U26178 ( .B(clk), .A(\g.we_clk [6596]));
Q_ASSIGN U26179 ( .B(clk), .A(\g.we_clk [6595]));
Q_ASSIGN U26180 ( .B(clk), .A(\g.we_clk [6594]));
Q_ASSIGN U26181 ( .B(clk), .A(\g.we_clk [6593]));
Q_ASSIGN U26182 ( .B(clk), .A(\g.we_clk [6592]));
Q_ASSIGN U26183 ( .B(clk), .A(\g.we_clk [6591]));
Q_ASSIGN U26184 ( .B(clk), .A(\g.we_clk [6590]));
Q_ASSIGN U26185 ( .B(clk), .A(\g.we_clk [6589]));
Q_ASSIGN U26186 ( .B(clk), .A(\g.we_clk [6588]));
Q_ASSIGN U26187 ( .B(clk), .A(\g.we_clk [6587]));
Q_ASSIGN U26188 ( .B(clk), .A(\g.we_clk [6586]));
Q_ASSIGN U26189 ( .B(clk), .A(\g.we_clk [6585]));
Q_ASSIGN U26190 ( .B(clk), .A(\g.we_clk [6584]));
Q_ASSIGN U26191 ( .B(clk), .A(\g.we_clk [6583]));
Q_ASSIGN U26192 ( .B(clk), .A(\g.we_clk [6582]));
Q_ASSIGN U26193 ( .B(clk), .A(\g.we_clk [6581]));
Q_ASSIGN U26194 ( .B(clk), .A(\g.we_clk [6580]));
Q_ASSIGN U26195 ( .B(clk), .A(\g.we_clk [6579]));
Q_ASSIGN U26196 ( .B(clk), .A(\g.we_clk [6578]));
Q_ASSIGN U26197 ( .B(clk), .A(\g.we_clk [6577]));
Q_ASSIGN U26198 ( .B(clk), .A(\g.we_clk [6576]));
Q_ASSIGN U26199 ( .B(clk), .A(\g.we_clk [6575]));
Q_ASSIGN U26200 ( .B(clk), .A(\g.we_clk [6574]));
Q_ASSIGN U26201 ( .B(clk), .A(\g.we_clk [6573]));
Q_ASSIGN U26202 ( .B(clk), .A(\g.we_clk [6572]));
Q_ASSIGN U26203 ( .B(clk), .A(\g.we_clk [6571]));
Q_ASSIGN U26204 ( .B(clk), .A(\g.we_clk [6570]));
Q_ASSIGN U26205 ( .B(clk), .A(\g.we_clk [6569]));
Q_ASSIGN U26206 ( .B(clk), .A(\g.we_clk [6568]));
Q_ASSIGN U26207 ( .B(clk), .A(\g.we_clk [6567]));
Q_ASSIGN U26208 ( .B(clk), .A(\g.we_clk [6566]));
Q_ASSIGN U26209 ( .B(clk), .A(\g.we_clk [6565]));
Q_ASSIGN U26210 ( .B(clk), .A(\g.we_clk [6564]));
Q_ASSIGN U26211 ( .B(clk), .A(\g.we_clk [6563]));
Q_ASSIGN U26212 ( .B(clk), .A(\g.we_clk [6562]));
Q_ASSIGN U26213 ( .B(clk), .A(\g.we_clk [6561]));
Q_ASSIGN U26214 ( .B(clk), .A(\g.we_clk [6560]));
Q_ASSIGN U26215 ( .B(clk), .A(\g.we_clk [6559]));
Q_ASSIGN U26216 ( .B(clk), .A(\g.we_clk [6558]));
Q_ASSIGN U26217 ( .B(clk), .A(\g.we_clk [6557]));
Q_ASSIGN U26218 ( .B(clk), .A(\g.we_clk [6556]));
Q_ASSIGN U26219 ( .B(clk), .A(\g.we_clk [6555]));
Q_ASSIGN U26220 ( .B(clk), .A(\g.we_clk [6554]));
Q_ASSIGN U26221 ( .B(clk), .A(\g.we_clk [6553]));
Q_ASSIGN U26222 ( .B(clk), .A(\g.we_clk [6552]));
Q_ASSIGN U26223 ( .B(clk), .A(\g.we_clk [6551]));
Q_ASSIGN U26224 ( .B(clk), .A(\g.we_clk [6550]));
Q_ASSIGN U26225 ( .B(clk), .A(\g.we_clk [6549]));
Q_ASSIGN U26226 ( .B(clk), .A(\g.we_clk [6548]));
Q_ASSIGN U26227 ( .B(clk), .A(\g.we_clk [6547]));
Q_ASSIGN U26228 ( .B(clk), .A(\g.we_clk [6546]));
Q_ASSIGN U26229 ( .B(clk), .A(\g.we_clk [6545]));
Q_ASSIGN U26230 ( .B(clk), .A(\g.we_clk [6544]));
Q_ASSIGN U26231 ( .B(clk), .A(\g.we_clk [6543]));
Q_ASSIGN U26232 ( .B(clk), .A(\g.we_clk [6542]));
Q_ASSIGN U26233 ( .B(clk), .A(\g.we_clk [6541]));
Q_ASSIGN U26234 ( .B(clk), .A(\g.we_clk [6540]));
Q_ASSIGN U26235 ( .B(clk), .A(\g.we_clk [6539]));
Q_ASSIGN U26236 ( .B(clk), .A(\g.we_clk [6538]));
Q_ASSIGN U26237 ( .B(clk), .A(\g.we_clk [6537]));
Q_ASSIGN U26238 ( .B(clk), .A(\g.we_clk [6536]));
Q_ASSIGN U26239 ( .B(clk), .A(\g.we_clk [6535]));
Q_ASSIGN U26240 ( .B(clk), .A(\g.we_clk [6534]));
Q_ASSIGN U26241 ( .B(clk), .A(\g.we_clk [6533]));
Q_ASSIGN U26242 ( .B(clk), .A(\g.we_clk [6532]));
Q_ASSIGN U26243 ( .B(clk), .A(\g.we_clk [6531]));
Q_ASSIGN U26244 ( .B(clk), .A(\g.we_clk [6530]));
Q_ASSIGN U26245 ( .B(clk), .A(\g.we_clk [6529]));
Q_ASSIGN U26246 ( .B(clk), .A(\g.we_clk [6528]));
Q_ASSIGN U26247 ( .B(clk), .A(\g.we_clk [6527]));
Q_ASSIGN U26248 ( .B(clk), .A(\g.we_clk [6526]));
Q_ASSIGN U26249 ( .B(clk), .A(\g.we_clk [6525]));
Q_ASSIGN U26250 ( .B(clk), .A(\g.we_clk [6524]));
Q_ASSIGN U26251 ( .B(clk), .A(\g.we_clk [6523]));
Q_ASSIGN U26252 ( .B(clk), .A(\g.we_clk [6522]));
Q_ASSIGN U26253 ( .B(clk), .A(\g.we_clk [6521]));
Q_ASSIGN U26254 ( .B(clk), .A(\g.we_clk [6520]));
Q_ASSIGN U26255 ( .B(clk), .A(\g.we_clk [6519]));
Q_ASSIGN U26256 ( .B(clk), .A(\g.we_clk [6518]));
Q_ASSIGN U26257 ( .B(clk), .A(\g.we_clk [6517]));
Q_ASSIGN U26258 ( .B(clk), .A(\g.we_clk [6516]));
Q_ASSIGN U26259 ( .B(clk), .A(\g.we_clk [6515]));
Q_ASSIGN U26260 ( .B(clk), .A(\g.we_clk [6514]));
Q_ASSIGN U26261 ( .B(clk), .A(\g.we_clk [6513]));
Q_ASSIGN U26262 ( .B(clk), .A(\g.we_clk [6512]));
Q_ASSIGN U26263 ( .B(clk), .A(\g.we_clk [6511]));
Q_ASSIGN U26264 ( .B(clk), .A(\g.we_clk [6510]));
Q_ASSIGN U26265 ( .B(clk), .A(\g.we_clk [6509]));
Q_ASSIGN U26266 ( .B(clk), .A(\g.we_clk [6508]));
Q_ASSIGN U26267 ( .B(clk), .A(\g.we_clk [6507]));
Q_ASSIGN U26268 ( .B(clk), .A(\g.we_clk [6506]));
Q_ASSIGN U26269 ( .B(clk), .A(\g.we_clk [6505]));
Q_ASSIGN U26270 ( .B(clk), .A(\g.we_clk [6504]));
Q_ASSIGN U26271 ( .B(clk), .A(\g.we_clk [6503]));
Q_ASSIGN U26272 ( .B(clk), .A(\g.we_clk [6502]));
Q_ASSIGN U26273 ( .B(clk), .A(\g.we_clk [6501]));
Q_ASSIGN U26274 ( .B(clk), .A(\g.we_clk [6500]));
Q_ASSIGN U26275 ( .B(clk), .A(\g.we_clk [6499]));
Q_ASSIGN U26276 ( .B(clk), .A(\g.we_clk [6498]));
Q_ASSIGN U26277 ( .B(clk), .A(\g.we_clk [6497]));
Q_ASSIGN U26278 ( .B(clk), .A(\g.we_clk [6496]));
Q_ASSIGN U26279 ( .B(clk), .A(\g.we_clk [6495]));
Q_ASSIGN U26280 ( .B(clk), .A(\g.we_clk [6494]));
Q_ASSIGN U26281 ( .B(clk), .A(\g.we_clk [6493]));
Q_ASSIGN U26282 ( .B(clk), .A(\g.we_clk [6492]));
Q_ASSIGN U26283 ( .B(clk), .A(\g.we_clk [6491]));
Q_ASSIGN U26284 ( .B(clk), .A(\g.we_clk [6490]));
Q_ASSIGN U26285 ( .B(clk), .A(\g.we_clk [6489]));
Q_ASSIGN U26286 ( .B(clk), .A(\g.we_clk [6488]));
Q_ASSIGN U26287 ( .B(clk), .A(\g.we_clk [6487]));
Q_ASSIGN U26288 ( .B(clk), .A(\g.we_clk [6486]));
Q_ASSIGN U26289 ( .B(clk), .A(\g.we_clk [6485]));
Q_ASSIGN U26290 ( .B(clk), .A(\g.we_clk [6484]));
Q_ASSIGN U26291 ( .B(clk), .A(\g.we_clk [6483]));
Q_ASSIGN U26292 ( .B(clk), .A(\g.we_clk [6482]));
Q_ASSIGN U26293 ( .B(clk), .A(\g.we_clk [6481]));
Q_ASSIGN U26294 ( .B(clk), .A(\g.we_clk [6480]));
Q_ASSIGN U26295 ( .B(clk), .A(\g.we_clk [6479]));
Q_ASSIGN U26296 ( .B(clk), .A(\g.we_clk [6478]));
Q_ASSIGN U26297 ( .B(clk), .A(\g.we_clk [6477]));
Q_ASSIGN U26298 ( .B(clk), .A(\g.we_clk [6476]));
Q_ASSIGN U26299 ( .B(clk), .A(\g.we_clk [6475]));
Q_ASSIGN U26300 ( .B(clk), .A(\g.we_clk [6474]));
Q_ASSIGN U26301 ( .B(clk), .A(\g.we_clk [6473]));
Q_ASSIGN U26302 ( .B(clk), .A(\g.we_clk [6472]));
Q_ASSIGN U26303 ( .B(clk), .A(\g.we_clk [6471]));
Q_ASSIGN U26304 ( .B(clk), .A(\g.we_clk [6470]));
Q_ASSIGN U26305 ( .B(clk), .A(\g.we_clk [6469]));
Q_ASSIGN U26306 ( .B(clk), .A(\g.we_clk [6468]));
Q_ASSIGN U26307 ( .B(clk), .A(\g.we_clk [6467]));
Q_ASSIGN U26308 ( .B(clk), .A(\g.we_clk [6466]));
Q_ASSIGN U26309 ( .B(clk), .A(\g.we_clk [6465]));
Q_ASSIGN U26310 ( .B(clk), .A(\g.we_clk [6464]));
Q_ASSIGN U26311 ( .B(clk), .A(\g.we_clk [6463]));
Q_ASSIGN U26312 ( .B(clk), .A(\g.we_clk [6462]));
Q_ASSIGN U26313 ( .B(clk), .A(\g.we_clk [6461]));
Q_ASSIGN U26314 ( .B(clk), .A(\g.we_clk [6460]));
Q_ASSIGN U26315 ( .B(clk), .A(\g.we_clk [6459]));
Q_ASSIGN U26316 ( .B(clk), .A(\g.we_clk [6458]));
Q_ASSIGN U26317 ( .B(clk), .A(\g.we_clk [6457]));
Q_ASSIGN U26318 ( .B(clk), .A(\g.we_clk [6456]));
Q_ASSIGN U26319 ( .B(clk), .A(\g.we_clk [6455]));
Q_ASSIGN U26320 ( .B(clk), .A(\g.we_clk [6454]));
Q_ASSIGN U26321 ( .B(clk), .A(\g.we_clk [6453]));
Q_ASSIGN U26322 ( .B(clk), .A(\g.we_clk [6452]));
Q_ASSIGN U26323 ( .B(clk), .A(\g.we_clk [6451]));
Q_ASSIGN U26324 ( .B(clk), .A(\g.we_clk [6450]));
Q_ASSIGN U26325 ( .B(clk), .A(\g.we_clk [6449]));
Q_ASSIGN U26326 ( .B(clk), .A(\g.we_clk [6448]));
Q_ASSIGN U26327 ( .B(clk), .A(\g.we_clk [6447]));
Q_ASSIGN U26328 ( .B(clk), .A(\g.we_clk [6446]));
Q_ASSIGN U26329 ( .B(clk), .A(\g.we_clk [6445]));
Q_ASSIGN U26330 ( .B(clk), .A(\g.we_clk [6444]));
Q_ASSIGN U26331 ( .B(clk), .A(\g.we_clk [6443]));
Q_ASSIGN U26332 ( .B(clk), .A(\g.we_clk [6442]));
Q_ASSIGN U26333 ( .B(clk), .A(\g.we_clk [6441]));
Q_ASSIGN U26334 ( .B(clk), .A(\g.we_clk [6440]));
Q_ASSIGN U26335 ( .B(clk), .A(\g.we_clk [6439]));
Q_ASSIGN U26336 ( .B(clk), .A(\g.we_clk [6438]));
Q_ASSIGN U26337 ( .B(clk), .A(\g.we_clk [6437]));
Q_ASSIGN U26338 ( .B(clk), .A(\g.we_clk [6436]));
Q_ASSIGN U26339 ( .B(clk), .A(\g.we_clk [6435]));
Q_ASSIGN U26340 ( .B(clk), .A(\g.we_clk [6434]));
Q_ASSIGN U26341 ( .B(clk), .A(\g.we_clk [6433]));
Q_ASSIGN U26342 ( .B(clk), .A(\g.we_clk [6432]));
Q_ASSIGN U26343 ( .B(clk), .A(\g.we_clk [6431]));
Q_ASSIGN U26344 ( .B(clk), .A(\g.we_clk [6430]));
Q_ASSIGN U26345 ( .B(clk), .A(\g.we_clk [6429]));
Q_ASSIGN U26346 ( .B(clk), .A(\g.we_clk [6428]));
Q_ASSIGN U26347 ( .B(clk), .A(\g.we_clk [6427]));
Q_ASSIGN U26348 ( .B(clk), .A(\g.we_clk [6426]));
Q_ASSIGN U26349 ( .B(clk), .A(\g.we_clk [6425]));
Q_ASSIGN U26350 ( .B(clk), .A(\g.we_clk [6424]));
Q_ASSIGN U26351 ( .B(clk), .A(\g.we_clk [6423]));
Q_ASSIGN U26352 ( .B(clk), .A(\g.we_clk [6422]));
Q_ASSIGN U26353 ( .B(clk), .A(\g.we_clk [6421]));
Q_ASSIGN U26354 ( .B(clk), .A(\g.we_clk [6420]));
Q_ASSIGN U26355 ( .B(clk), .A(\g.we_clk [6419]));
Q_ASSIGN U26356 ( .B(clk), .A(\g.we_clk [6418]));
Q_ASSIGN U26357 ( .B(clk), .A(\g.we_clk [6417]));
Q_ASSIGN U26358 ( .B(clk), .A(\g.we_clk [6416]));
Q_ASSIGN U26359 ( .B(clk), .A(\g.we_clk [6415]));
Q_ASSIGN U26360 ( .B(clk), .A(\g.we_clk [6414]));
Q_ASSIGN U26361 ( .B(clk), .A(\g.we_clk [6413]));
Q_ASSIGN U26362 ( .B(clk), .A(\g.we_clk [6412]));
Q_ASSIGN U26363 ( .B(clk), .A(\g.we_clk [6411]));
Q_ASSIGN U26364 ( .B(clk), .A(\g.we_clk [6410]));
Q_ASSIGN U26365 ( .B(clk), .A(\g.we_clk [6409]));
Q_ASSIGN U26366 ( .B(clk), .A(\g.we_clk [6408]));
Q_ASSIGN U26367 ( .B(clk), .A(\g.we_clk [6407]));
Q_ASSIGN U26368 ( .B(clk), .A(\g.we_clk [6406]));
Q_ASSIGN U26369 ( .B(clk), .A(\g.we_clk [6405]));
Q_ASSIGN U26370 ( .B(clk), .A(\g.we_clk [6404]));
Q_ASSIGN U26371 ( .B(clk), .A(\g.we_clk [6403]));
Q_ASSIGN U26372 ( .B(clk), .A(\g.we_clk [6402]));
Q_ASSIGN U26373 ( .B(clk), .A(\g.we_clk [6401]));
Q_ASSIGN U26374 ( .B(clk), .A(\g.we_clk [6400]));
Q_ASSIGN U26375 ( .B(clk), .A(\g.we_clk [6399]));
Q_ASSIGN U26376 ( .B(clk), .A(\g.we_clk [6398]));
Q_ASSIGN U26377 ( .B(clk), .A(\g.we_clk [6397]));
Q_ASSIGN U26378 ( .B(clk), .A(\g.we_clk [6396]));
Q_ASSIGN U26379 ( .B(clk), .A(\g.we_clk [6395]));
Q_ASSIGN U26380 ( .B(clk), .A(\g.we_clk [6394]));
Q_ASSIGN U26381 ( .B(clk), .A(\g.we_clk [6393]));
Q_ASSIGN U26382 ( .B(clk), .A(\g.we_clk [6392]));
Q_ASSIGN U26383 ( .B(clk), .A(\g.we_clk [6391]));
Q_ASSIGN U26384 ( .B(clk), .A(\g.we_clk [6390]));
Q_ASSIGN U26385 ( .B(clk), .A(\g.we_clk [6389]));
Q_ASSIGN U26386 ( .B(clk), .A(\g.we_clk [6388]));
Q_ASSIGN U26387 ( .B(clk), .A(\g.we_clk [6387]));
Q_ASSIGN U26388 ( .B(clk), .A(\g.we_clk [6386]));
Q_ASSIGN U26389 ( .B(clk), .A(\g.we_clk [6385]));
Q_ASSIGN U26390 ( .B(clk), .A(\g.we_clk [6384]));
Q_ASSIGN U26391 ( .B(clk), .A(\g.we_clk [6383]));
Q_ASSIGN U26392 ( .B(clk), .A(\g.we_clk [6382]));
Q_ASSIGN U26393 ( .B(clk), .A(\g.we_clk [6381]));
Q_ASSIGN U26394 ( .B(clk), .A(\g.we_clk [6380]));
Q_ASSIGN U26395 ( .B(clk), .A(\g.we_clk [6379]));
Q_ASSIGN U26396 ( .B(clk), .A(\g.we_clk [6378]));
Q_ASSIGN U26397 ( .B(clk), .A(\g.we_clk [6377]));
Q_ASSIGN U26398 ( .B(clk), .A(\g.we_clk [6376]));
Q_ASSIGN U26399 ( .B(clk), .A(\g.we_clk [6375]));
Q_ASSIGN U26400 ( .B(clk), .A(\g.we_clk [6374]));
Q_ASSIGN U26401 ( .B(clk), .A(\g.we_clk [6373]));
Q_ASSIGN U26402 ( .B(clk), .A(\g.we_clk [6372]));
Q_ASSIGN U26403 ( .B(clk), .A(\g.we_clk [6371]));
Q_ASSIGN U26404 ( .B(clk), .A(\g.we_clk [6370]));
Q_ASSIGN U26405 ( .B(clk), .A(\g.we_clk [6369]));
Q_ASSIGN U26406 ( .B(clk), .A(\g.we_clk [6368]));
Q_ASSIGN U26407 ( .B(clk), .A(\g.we_clk [6367]));
Q_ASSIGN U26408 ( .B(clk), .A(\g.we_clk [6366]));
Q_ASSIGN U26409 ( .B(clk), .A(\g.we_clk [6365]));
Q_ASSIGN U26410 ( .B(clk), .A(\g.we_clk [6364]));
Q_ASSIGN U26411 ( .B(clk), .A(\g.we_clk [6363]));
Q_ASSIGN U26412 ( .B(clk), .A(\g.we_clk [6362]));
Q_ASSIGN U26413 ( .B(clk), .A(\g.we_clk [6361]));
Q_ASSIGN U26414 ( .B(clk), .A(\g.we_clk [6360]));
Q_ASSIGN U26415 ( .B(clk), .A(\g.we_clk [6359]));
Q_ASSIGN U26416 ( .B(clk), .A(\g.we_clk [6358]));
Q_ASSIGN U26417 ( .B(clk), .A(\g.we_clk [6357]));
Q_ASSIGN U26418 ( .B(clk), .A(\g.we_clk [6356]));
Q_ASSIGN U26419 ( .B(clk), .A(\g.we_clk [6355]));
Q_ASSIGN U26420 ( .B(clk), .A(\g.we_clk [6354]));
Q_ASSIGN U26421 ( .B(clk), .A(\g.we_clk [6353]));
Q_ASSIGN U26422 ( .B(clk), .A(\g.we_clk [6352]));
Q_ASSIGN U26423 ( .B(clk), .A(\g.we_clk [6351]));
Q_ASSIGN U26424 ( .B(clk), .A(\g.we_clk [6350]));
Q_ASSIGN U26425 ( .B(clk), .A(\g.we_clk [6349]));
Q_ASSIGN U26426 ( .B(clk), .A(\g.we_clk [6348]));
Q_ASSIGN U26427 ( .B(clk), .A(\g.we_clk [6347]));
Q_ASSIGN U26428 ( .B(clk), .A(\g.we_clk [6346]));
Q_ASSIGN U26429 ( .B(clk), .A(\g.we_clk [6345]));
Q_ASSIGN U26430 ( .B(clk), .A(\g.we_clk [6344]));
Q_ASSIGN U26431 ( .B(clk), .A(\g.we_clk [6343]));
Q_ASSIGN U26432 ( .B(clk), .A(\g.we_clk [6342]));
Q_ASSIGN U26433 ( .B(clk), .A(\g.we_clk [6341]));
Q_ASSIGN U26434 ( .B(clk), .A(\g.we_clk [6340]));
Q_ASSIGN U26435 ( .B(clk), .A(\g.we_clk [6339]));
Q_ASSIGN U26436 ( .B(clk), .A(\g.we_clk [6338]));
Q_ASSIGN U26437 ( .B(clk), .A(\g.we_clk [6337]));
Q_ASSIGN U26438 ( .B(clk), .A(\g.we_clk [6336]));
Q_ASSIGN U26439 ( .B(clk), .A(\g.we_clk [6335]));
Q_ASSIGN U26440 ( .B(clk), .A(\g.we_clk [6334]));
Q_ASSIGN U26441 ( .B(clk), .A(\g.we_clk [6333]));
Q_ASSIGN U26442 ( .B(clk), .A(\g.we_clk [6332]));
Q_ASSIGN U26443 ( .B(clk), .A(\g.we_clk [6331]));
Q_ASSIGN U26444 ( .B(clk), .A(\g.we_clk [6330]));
Q_ASSIGN U26445 ( .B(clk), .A(\g.we_clk [6329]));
Q_ASSIGN U26446 ( .B(clk), .A(\g.we_clk [6328]));
Q_ASSIGN U26447 ( .B(clk), .A(\g.we_clk [6327]));
Q_ASSIGN U26448 ( .B(clk), .A(\g.we_clk [6326]));
Q_ASSIGN U26449 ( .B(clk), .A(\g.we_clk [6325]));
Q_ASSIGN U26450 ( .B(clk), .A(\g.we_clk [6324]));
Q_ASSIGN U26451 ( .B(clk), .A(\g.we_clk [6323]));
Q_ASSIGN U26452 ( .B(clk), .A(\g.we_clk [6322]));
Q_ASSIGN U26453 ( .B(clk), .A(\g.we_clk [6321]));
Q_ASSIGN U26454 ( .B(clk), .A(\g.we_clk [6320]));
Q_ASSIGN U26455 ( .B(clk), .A(\g.we_clk [6319]));
Q_ASSIGN U26456 ( .B(clk), .A(\g.we_clk [6318]));
Q_ASSIGN U26457 ( .B(clk), .A(\g.we_clk [6317]));
Q_ASSIGN U26458 ( .B(clk), .A(\g.we_clk [6316]));
Q_ASSIGN U26459 ( .B(clk), .A(\g.we_clk [6315]));
Q_ASSIGN U26460 ( .B(clk), .A(\g.we_clk [6314]));
Q_ASSIGN U26461 ( .B(clk), .A(\g.we_clk [6313]));
Q_ASSIGN U26462 ( .B(clk), .A(\g.we_clk [6312]));
Q_ASSIGN U26463 ( .B(clk), .A(\g.we_clk [6311]));
Q_ASSIGN U26464 ( .B(clk), .A(\g.we_clk [6310]));
Q_ASSIGN U26465 ( .B(clk), .A(\g.we_clk [6309]));
Q_ASSIGN U26466 ( .B(clk), .A(\g.we_clk [6308]));
Q_ASSIGN U26467 ( .B(clk), .A(\g.we_clk [6307]));
Q_ASSIGN U26468 ( .B(clk), .A(\g.we_clk [6306]));
Q_ASSIGN U26469 ( .B(clk), .A(\g.we_clk [6305]));
Q_ASSIGN U26470 ( .B(clk), .A(\g.we_clk [6304]));
Q_ASSIGN U26471 ( .B(clk), .A(\g.we_clk [6303]));
Q_ASSIGN U26472 ( .B(clk), .A(\g.we_clk [6302]));
Q_ASSIGN U26473 ( .B(clk), .A(\g.we_clk [6301]));
Q_ASSIGN U26474 ( .B(clk), .A(\g.we_clk [6300]));
Q_ASSIGN U26475 ( .B(clk), .A(\g.we_clk [6299]));
Q_ASSIGN U26476 ( .B(clk), .A(\g.we_clk [6298]));
Q_ASSIGN U26477 ( .B(clk), .A(\g.we_clk [6297]));
Q_ASSIGN U26478 ( .B(clk), .A(\g.we_clk [6296]));
Q_ASSIGN U26479 ( .B(clk), .A(\g.we_clk [6295]));
Q_ASSIGN U26480 ( .B(clk), .A(\g.we_clk [6294]));
Q_ASSIGN U26481 ( .B(clk), .A(\g.we_clk [6293]));
Q_ASSIGN U26482 ( .B(clk), .A(\g.we_clk [6292]));
Q_ASSIGN U26483 ( .B(clk), .A(\g.we_clk [6291]));
Q_ASSIGN U26484 ( .B(clk), .A(\g.we_clk [6290]));
Q_ASSIGN U26485 ( .B(clk), .A(\g.we_clk [6289]));
Q_ASSIGN U26486 ( .B(clk), .A(\g.we_clk [6288]));
Q_ASSIGN U26487 ( .B(clk), .A(\g.we_clk [6287]));
Q_ASSIGN U26488 ( .B(clk), .A(\g.we_clk [6286]));
Q_ASSIGN U26489 ( .B(clk), .A(\g.we_clk [6285]));
Q_ASSIGN U26490 ( .B(clk), .A(\g.we_clk [6284]));
Q_ASSIGN U26491 ( .B(clk), .A(\g.we_clk [6283]));
Q_ASSIGN U26492 ( .B(clk), .A(\g.we_clk [6282]));
Q_ASSIGN U26493 ( .B(clk), .A(\g.we_clk [6281]));
Q_ASSIGN U26494 ( .B(clk), .A(\g.we_clk [6280]));
Q_ASSIGN U26495 ( .B(clk), .A(\g.we_clk [6279]));
Q_ASSIGN U26496 ( .B(clk), .A(\g.we_clk [6278]));
Q_ASSIGN U26497 ( .B(clk), .A(\g.we_clk [6277]));
Q_ASSIGN U26498 ( .B(clk), .A(\g.we_clk [6276]));
Q_ASSIGN U26499 ( .B(clk), .A(\g.we_clk [6275]));
Q_ASSIGN U26500 ( .B(clk), .A(\g.we_clk [6274]));
Q_ASSIGN U26501 ( .B(clk), .A(\g.we_clk [6273]));
Q_ASSIGN U26502 ( .B(clk), .A(\g.we_clk [6272]));
Q_ASSIGN U26503 ( .B(clk), .A(\g.we_clk [6271]));
Q_ASSIGN U26504 ( .B(clk), .A(\g.we_clk [6270]));
Q_ASSIGN U26505 ( .B(clk), .A(\g.we_clk [6269]));
Q_ASSIGN U26506 ( .B(clk), .A(\g.we_clk [6268]));
Q_ASSIGN U26507 ( .B(clk), .A(\g.we_clk [6267]));
Q_ASSIGN U26508 ( .B(clk), .A(\g.we_clk [6266]));
Q_ASSIGN U26509 ( .B(clk), .A(\g.we_clk [6265]));
Q_ASSIGN U26510 ( .B(clk), .A(\g.we_clk [6264]));
Q_ASSIGN U26511 ( .B(clk), .A(\g.we_clk [6263]));
Q_ASSIGN U26512 ( .B(clk), .A(\g.we_clk [6262]));
Q_ASSIGN U26513 ( .B(clk), .A(\g.we_clk [6261]));
Q_ASSIGN U26514 ( .B(clk), .A(\g.we_clk [6260]));
Q_ASSIGN U26515 ( .B(clk), .A(\g.we_clk [6259]));
Q_ASSIGN U26516 ( .B(clk), .A(\g.we_clk [6258]));
Q_ASSIGN U26517 ( .B(clk), .A(\g.we_clk [6257]));
Q_ASSIGN U26518 ( .B(clk), .A(\g.we_clk [6256]));
Q_ASSIGN U26519 ( .B(clk), .A(\g.we_clk [6255]));
Q_ASSIGN U26520 ( .B(clk), .A(\g.we_clk [6254]));
Q_ASSIGN U26521 ( .B(clk), .A(\g.we_clk [6253]));
Q_ASSIGN U26522 ( .B(clk), .A(\g.we_clk [6252]));
Q_ASSIGN U26523 ( .B(clk), .A(\g.we_clk [6251]));
Q_ASSIGN U26524 ( .B(clk), .A(\g.we_clk [6250]));
Q_ASSIGN U26525 ( .B(clk), .A(\g.we_clk [6249]));
Q_ASSIGN U26526 ( .B(clk), .A(\g.we_clk [6248]));
Q_ASSIGN U26527 ( .B(clk), .A(\g.we_clk [6247]));
Q_ASSIGN U26528 ( .B(clk), .A(\g.we_clk [6246]));
Q_ASSIGN U26529 ( .B(clk), .A(\g.we_clk [6245]));
Q_ASSIGN U26530 ( .B(clk), .A(\g.we_clk [6244]));
Q_ASSIGN U26531 ( .B(clk), .A(\g.we_clk [6243]));
Q_ASSIGN U26532 ( .B(clk), .A(\g.we_clk [6242]));
Q_ASSIGN U26533 ( .B(clk), .A(\g.we_clk [6241]));
Q_ASSIGN U26534 ( .B(clk), .A(\g.we_clk [6240]));
Q_ASSIGN U26535 ( .B(clk), .A(\g.we_clk [6239]));
Q_ASSIGN U26536 ( .B(clk), .A(\g.we_clk [6238]));
Q_ASSIGN U26537 ( .B(clk), .A(\g.we_clk [6237]));
Q_ASSIGN U26538 ( .B(clk), .A(\g.we_clk [6236]));
Q_ASSIGN U26539 ( .B(clk), .A(\g.we_clk [6235]));
Q_ASSIGN U26540 ( .B(clk), .A(\g.we_clk [6234]));
Q_ASSIGN U26541 ( .B(clk), .A(\g.we_clk [6233]));
Q_ASSIGN U26542 ( .B(clk), .A(\g.we_clk [6232]));
Q_ASSIGN U26543 ( .B(clk), .A(\g.we_clk [6231]));
Q_ASSIGN U26544 ( .B(clk), .A(\g.we_clk [6230]));
Q_ASSIGN U26545 ( .B(clk), .A(\g.we_clk [6229]));
Q_ASSIGN U26546 ( .B(clk), .A(\g.we_clk [6228]));
Q_ASSIGN U26547 ( .B(clk), .A(\g.we_clk [6227]));
Q_ASSIGN U26548 ( .B(clk), .A(\g.we_clk [6226]));
Q_ASSIGN U26549 ( .B(clk), .A(\g.we_clk [6225]));
Q_ASSIGN U26550 ( .B(clk), .A(\g.we_clk [6224]));
Q_ASSIGN U26551 ( .B(clk), .A(\g.we_clk [6223]));
Q_ASSIGN U26552 ( .B(clk), .A(\g.we_clk [6222]));
Q_ASSIGN U26553 ( .B(clk), .A(\g.we_clk [6221]));
Q_ASSIGN U26554 ( .B(clk), .A(\g.we_clk [6220]));
Q_ASSIGN U26555 ( .B(clk), .A(\g.we_clk [6219]));
Q_ASSIGN U26556 ( .B(clk), .A(\g.we_clk [6218]));
Q_ASSIGN U26557 ( .B(clk), .A(\g.we_clk [6217]));
Q_ASSIGN U26558 ( .B(clk), .A(\g.we_clk [6216]));
Q_ASSIGN U26559 ( .B(clk), .A(\g.we_clk [6215]));
Q_ASSIGN U26560 ( .B(clk), .A(\g.we_clk [6214]));
Q_ASSIGN U26561 ( .B(clk), .A(\g.we_clk [6213]));
Q_ASSIGN U26562 ( .B(clk), .A(\g.we_clk [6212]));
Q_ASSIGN U26563 ( .B(clk), .A(\g.we_clk [6211]));
Q_ASSIGN U26564 ( .B(clk), .A(\g.we_clk [6210]));
Q_ASSIGN U26565 ( .B(clk), .A(\g.we_clk [6209]));
Q_ASSIGN U26566 ( .B(clk), .A(\g.we_clk [6208]));
Q_ASSIGN U26567 ( .B(clk), .A(\g.we_clk [6207]));
Q_ASSIGN U26568 ( .B(clk), .A(\g.we_clk [6206]));
Q_ASSIGN U26569 ( .B(clk), .A(\g.we_clk [6205]));
Q_ASSIGN U26570 ( .B(clk), .A(\g.we_clk [6204]));
Q_ASSIGN U26571 ( .B(clk), .A(\g.we_clk [6203]));
Q_ASSIGN U26572 ( .B(clk), .A(\g.we_clk [6202]));
Q_ASSIGN U26573 ( .B(clk), .A(\g.we_clk [6201]));
Q_ASSIGN U26574 ( .B(clk), .A(\g.we_clk [6200]));
Q_ASSIGN U26575 ( .B(clk), .A(\g.we_clk [6199]));
Q_ASSIGN U26576 ( .B(clk), .A(\g.we_clk [6198]));
Q_ASSIGN U26577 ( .B(clk), .A(\g.we_clk [6197]));
Q_ASSIGN U26578 ( .B(clk), .A(\g.we_clk [6196]));
Q_ASSIGN U26579 ( .B(clk), .A(\g.we_clk [6195]));
Q_ASSIGN U26580 ( .B(clk), .A(\g.we_clk [6194]));
Q_ASSIGN U26581 ( .B(clk), .A(\g.we_clk [6193]));
Q_ASSIGN U26582 ( .B(clk), .A(\g.we_clk [6192]));
Q_ASSIGN U26583 ( .B(clk), .A(\g.we_clk [6191]));
Q_ASSIGN U26584 ( .B(clk), .A(\g.we_clk [6190]));
Q_ASSIGN U26585 ( .B(clk), .A(\g.we_clk [6189]));
Q_ASSIGN U26586 ( .B(clk), .A(\g.we_clk [6188]));
Q_ASSIGN U26587 ( .B(clk), .A(\g.we_clk [6187]));
Q_ASSIGN U26588 ( .B(clk), .A(\g.we_clk [6186]));
Q_ASSIGN U26589 ( .B(clk), .A(\g.we_clk [6185]));
Q_ASSIGN U26590 ( .B(clk), .A(\g.we_clk [6184]));
Q_ASSIGN U26591 ( .B(clk), .A(\g.we_clk [6183]));
Q_ASSIGN U26592 ( .B(clk), .A(\g.we_clk [6182]));
Q_ASSIGN U26593 ( .B(clk), .A(\g.we_clk [6181]));
Q_ASSIGN U26594 ( .B(clk), .A(\g.we_clk [6180]));
Q_ASSIGN U26595 ( .B(clk), .A(\g.we_clk [6179]));
Q_ASSIGN U26596 ( .B(clk), .A(\g.we_clk [6178]));
Q_ASSIGN U26597 ( .B(clk), .A(\g.we_clk [6177]));
Q_ASSIGN U26598 ( .B(clk), .A(\g.we_clk [6176]));
Q_ASSIGN U26599 ( .B(clk), .A(\g.we_clk [6175]));
Q_ASSIGN U26600 ( .B(clk), .A(\g.we_clk [6174]));
Q_ASSIGN U26601 ( .B(clk), .A(\g.we_clk [6173]));
Q_ASSIGN U26602 ( .B(clk), .A(\g.we_clk [6172]));
Q_ASSIGN U26603 ( .B(clk), .A(\g.we_clk [6171]));
Q_ASSIGN U26604 ( .B(clk), .A(\g.we_clk [6170]));
Q_ASSIGN U26605 ( .B(clk), .A(\g.we_clk [6169]));
Q_ASSIGN U26606 ( .B(clk), .A(\g.we_clk [6168]));
Q_ASSIGN U26607 ( .B(clk), .A(\g.we_clk [6167]));
Q_ASSIGN U26608 ( .B(clk), .A(\g.we_clk [6166]));
Q_ASSIGN U26609 ( .B(clk), .A(\g.we_clk [6165]));
Q_ASSIGN U26610 ( .B(clk), .A(\g.we_clk [6164]));
Q_ASSIGN U26611 ( .B(clk), .A(\g.we_clk [6163]));
Q_ASSIGN U26612 ( .B(clk), .A(\g.we_clk [6162]));
Q_ASSIGN U26613 ( .B(clk), .A(\g.we_clk [6161]));
Q_ASSIGN U26614 ( .B(clk), .A(\g.we_clk [6160]));
Q_ASSIGN U26615 ( .B(clk), .A(\g.we_clk [6159]));
Q_ASSIGN U26616 ( .B(clk), .A(\g.we_clk [6158]));
Q_ASSIGN U26617 ( .B(clk), .A(\g.we_clk [6157]));
Q_ASSIGN U26618 ( .B(clk), .A(\g.we_clk [6156]));
Q_ASSIGN U26619 ( .B(clk), .A(\g.we_clk [6155]));
Q_ASSIGN U26620 ( .B(clk), .A(\g.we_clk [6154]));
Q_ASSIGN U26621 ( .B(clk), .A(\g.we_clk [6153]));
Q_ASSIGN U26622 ( .B(clk), .A(\g.we_clk [6152]));
Q_ASSIGN U26623 ( .B(clk), .A(\g.we_clk [6151]));
Q_ASSIGN U26624 ( .B(clk), .A(\g.we_clk [6150]));
Q_ASSIGN U26625 ( .B(clk), .A(\g.we_clk [6149]));
Q_ASSIGN U26626 ( .B(clk), .A(\g.we_clk [6148]));
Q_ASSIGN U26627 ( .B(clk), .A(\g.we_clk [6147]));
Q_ASSIGN U26628 ( .B(clk), .A(\g.we_clk [6146]));
Q_ASSIGN U26629 ( .B(clk), .A(\g.we_clk [6145]));
Q_ASSIGN U26630 ( .B(clk), .A(\g.we_clk [6144]));
Q_ASSIGN U26631 ( .B(clk), .A(\g.we_clk [6143]));
Q_ASSIGN U26632 ( .B(clk), .A(\g.we_clk [6142]));
Q_ASSIGN U26633 ( .B(clk), .A(\g.we_clk [6141]));
Q_ASSIGN U26634 ( .B(clk), .A(\g.we_clk [6140]));
Q_ASSIGN U26635 ( .B(clk), .A(\g.we_clk [6139]));
Q_ASSIGN U26636 ( .B(clk), .A(\g.we_clk [6138]));
Q_ASSIGN U26637 ( .B(clk), .A(\g.we_clk [6137]));
Q_ASSIGN U26638 ( .B(clk), .A(\g.we_clk [6136]));
Q_ASSIGN U26639 ( .B(clk), .A(\g.we_clk [6135]));
Q_ASSIGN U26640 ( .B(clk), .A(\g.we_clk [6134]));
Q_ASSIGN U26641 ( .B(clk), .A(\g.we_clk [6133]));
Q_ASSIGN U26642 ( .B(clk), .A(\g.we_clk [6132]));
Q_ASSIGN U26643 ( .B(clk), .A(\g.we_clk [6131]));
Q_ASSIGN U26644 ( .B(clk), .A(\g.we_clk [6130]));
Q_ASSIGN U26645 ( .B(clk), .A(\g.we_clk [6129]));
Q_ASSIGN U26646 ( .B(clk), .A(\g.we_clk [6128]));
Q_ASSIGN U26647 ( .B(clk), .A(\g.we_clk [6127]));
Q_ASSIGN U26648 ( .B(clk), .A(\g.we_clk [6126]));
Q_ASSIGN U26649 ( .B(clk), .A(\g.we_clk [6125]));
Q_ASSIGN U26650 ( .B(clk), .A(\g.we_clk [6124]));
Q_ASSIGN U26651 ( .B(clk), .A(\g.we_clk [6123]));
Q_ASSIGN U26652 ( .B(clk), .A(\g.we_clk [6122]));
Q_ASSIGN U26653 ( .B(clk), .A(\g.we_clk [6121]));
Q_ASSIGN U26654 ( .B(clk), .A(\g.we_clk [6120]));
Q_ASSIGN U26655 ( .B(clk), .A(\g.we_clk [6119]));
Q_ASSIGN U26656 ( .B(clk), .A(\g.we_clk [6118]));
Q_ASSIGN U26657 ( .B(clk), .A(\g.we_clk [6117]));
Q_ASSIGN U26658 ( .B(clk), .A(\g.we_clk [6116]));
Q_ASSIGN U26659 ( .B(clk), .A(\g.we_clk [6115]));
Q_ASSIGN U26660 ( .B(clk), .A(\g.we_clk [6114]));
Q_ASSIGN U26661 ( .B(clk), .A(\g.we_clk [6113]));
Q_ASSIGN U26662 ( .B(clk), .A(\g.we_clk [6112]));
Q_ASSIGN U26663 ( .B(clk), .A(\g.we_clk [6111]));
Q_ASSIGN U26664 ( .B(clk), .A(\g.we_clk [6110]));
Q_ASSIGN U26665 ( .B(clk), .A(\g.we_clk [6109]));
Q_ASSIGN U26666 ( .B(clk), .A(\g.we_clk [6108]));
Q_ASSIGN U26667 ( .B(clk), .A(\g.we_clk [6107]));
Q_ASSIGN U26668 ( .B(clk), .A(\g.we_clk [6106]));
Q_ASSIGN U26669 ( .B(clk), .A(\g.we_clk [6105]));
Q_ASSIGN U26670 ( .B(clk), .A(\g.we_clk [6104]));
Q_ASSIGN U26671 ( .B(clk), .A(\g.we_clk [6103]));
Q_ASSIGN U26672 ( .B(clk), .A(\g.we_clk [6102]));
Q_ASSIGN U26673 ( .B(clk), .A(\g.we_clk [6101]));
Q_ASSIGN U26674 ( .B(clk), .A(\g.we_clk [6100]));
Q_ASSIGN U26675 ( .B(clk), .A(\g.we_clk [6099]));
Q_ASSIGN U26676 ( .B(clk), .A(\g.we_clk [6098]));
Q_ASSIGN U26677 ( .B(clk), .A(\g.we_clk [6097]));
Q_ASSIGN U26678 ( .B(clk), .A(\g.we_clk [6096]));
Q_ASSIGN U26679 ( .B(clk), .A(\g.we_clk [6095]));
Q_ASSIGN U26680 ( .B(clk), .A(\g.we_clk [6094]));
Q_ASSIGN U26681 ( .B(clk), .A(\g.we_clk [6093]));
Q_ASSIGN U26682 ( .B(clk), .A(\g.we_clk [6092]));
Q_ASSIGN U26683 ( .B(clk), .A(\g.we_clk [6091]));
Q_ASSIGN U26684 ( .B(clk), .A(\g.we_clk [6090]));
Q_ASSIGN U26685 ( .B(clk), .A(\g.we_clk [6089]));
Q_ASSIGN U26686 ( .B(clk), .A(\g.we_clk [6088]));
Q_ASSIGN U26687 ( .B(clk), .A(\g.we_clk [6087]));
Q_ASSIGN U26688 ( .B(clk), .A(\g.we_clk [6086]));
Q_ASSIGN U26689 ( .B(clk), .A(\g.we_clk [6085]));
Q_ASSIGN U26690 ( .B(clk), .A(\g.we_clk [6084]));
Q_ASSIGN U26691 ( .B(clk), .A(\g.we_clk [6083]));
Q_ASSIGN U26692 ( .B(clk), .A(\g.we_clk [6082]));
Q_ASSIGN U26693 ( .B(clk), .A(\g.we_clk [6081]));
Q_ASSIGN U26694 ( .B(clk), .A(\g.we_clk [6080]));
Q_ASSIGN U26695 ( .B(clk), .A(\g.we_clk [6079]));
Q_ASSIGN U26696 ( .B(clk), .A(\g.we_clk [6078]));
Q_ASSIGN U26697 ( .B(clk), .A(\g.we_clk [6077]));
Q_ASSIGN U26698 ( .B(clk), .A(\g.we_clk [6076]));
Q_ASSIGN U26699 ( .B(clk), .A(\g.we_clk [6075]));
Q_ASSIGN U26700 ( .B(clk), .A(\g.we_clk [6074]));
Q_ASSIGN U26701 ( .B(clk), .A(\g.we_clk [6073]));
Q_ASSIGN U26702 ( .B(clk), .A(\g.we_clk [6072]));
Q_ASSIGN U26703 ( .B(clk), .A(\g.we_clk [6071]));
Q_ASSIGN U26704 ( .B(clk), .A(\g.we_clk [6070]));
Q_ASSIGN U26705 ( .B(clk), .A(\g.we_clk [6069]));
Q_ASSIGN U26706 ( .B(clk), .A(\g.we_clk [6068]));
Q_ASSIGN U26707 ( .B(clk), .A(\g.we_clk [6067]));
Q_ASSIGN U26708 ( .B(clk), .A(\g.we_clk [6066]));
Q_ASSIGN U26709 ( .B(clk), .A(\g.we_clk [6065]));
Q_ASSIGN U26710 ( .B(clk), .A(\g.we_clk [6064]));
Q_ASSIGN U26711 ( .B(clk), .A(\g.we_clk [6063]));
Q_ASSIGN U26712 ( .B(clk), .A(\g.we_clk [6062]));
Q_ASSIGN U26713 ( .B(clk), .A(\g.we_clk [6061]));
Q_ASSIGN U26714 ( .B(clk), .A(\g.we_clk [6060]));
Q_ASSIGN U26715 ( .B(clk), .A(\g.we_clk [6059]));
Q_ASSIGN U26716 ( .B(clk), .A(\g.we_clk [6058]));
Q_ASSIGN U26717 ( .B(clk), .A(\g.we_clk [6057]));
Q_ASSIGN U26718 ( .B(clk), .A(\g.we_clk [6056]));
Q_ASSIGN U26719 ( .B(clk), .A(\g.we_clk [6055]));
Q_ASSIGN U26720 ( .B(clk), .A(\g.we_clk [6054]));
Q_ASSIGN U26721 ( .B(clk), .A(\g.we_clk [6053]));
Q_ASSIGN U26722 ( .B(clk), .A(\g.we_clk [6052]));
Q_ASSIGN U26723 ( .B(clk), .A(\g.we_clk [6051]));
Q_ASSIGN U26724 ( .B(clk), .A(\g.we_clk [6050]));
Q_ASSIGN U26725 ( .B(clk), .A(\g.we_clk [6049]));
Q_ASSIGN U26726 ( .B(clk), .A(\g.we_clk [6048]));
Q_ASSIGN U26727 ( .B(clk), .A(\g.we_clk [6047]));
Q_ASSIGN U26728 ( .B(clk), .A(\g.we_clk [6046]));
Q_ASSIGN U26729 ( .B(clk), .A(\g.we_clk [6045]));
Q_ASSIGN U26730 ( .B(clk), .A(\g.we_clk [6044]));
Q_ASSIGN U26731 ( .B(clk), .A(\g.we_clk [6043]));
Q_ASSIGN U26732 ( .B(clk), .A(\g.we_clk [6042]));
Q_ASSIGN U26733 ( .B(clk), .A(\g.we_clk [6041]));
Q_ASSIGN U26734 ( .B(clk), .A(\g.we_clk [6040]));
Q_ASSIGN U26735 ( .B(clk), .A(\g.we_clk [6039]));
Q_ASSIGN U26736 ( .B(clk), .A(\g.we_clk [6038]));
Q_ASSIGN U26737 ( .B(clk), .A(\g.we_clk [6037]));
Q_ASSIGN U26738 ( .B(clk), .A(\g.we_clk [6036]));
Q_ASSIGN U26739 ( .B(clk), .A(\g.we_clk [6035]));
Q_ASSIGN U26740 ( .B(clk), .A(\g.we_clk [6034]));
Q_ASSIGN U26741 ( .B(clk), .A(\g.we_clk [6033]));
Q_ASSIGN U26742 ( .B(clk), .A(\g.we_clk [6032]));
Q_ASSIGN U26743 ( .B(clk), .A(\g.we_clk [6031]));
Q_ASSIGN U26744 ( .B(clk), .A(\g.we_clk [6030]));
Q_ASSIGN U26745 ( .B(clk), .A(\g.we_clk [6029]));
Q_ASSIGN U26746 ( .B(clk), .A(\g.we_clk [6028]));
Q_ASSIGN U26747 ( .B(clk), .A(\g.we_clk [6027]));
Q_ASSIGN U26748 ( .B(clk), .A(\g.we_clk [6026]));
Q_ASSIGN U26749 ( .B(clk), .A(\g.we_clk [6025]));
Q_ASSIGN U26750 ( .B(clk), .A(\g.we_clk [6024]));
Q_ASSIGN U26751 ( .B(clk), .A(\g.we_clk [6023]));
Q_ASSIGN U26752 ( .B(clk), .A(\g.we_clk [6022]));
Q_ASSIGN U26753 ( .B(clk), .A(\g.we_clk [6021]));
Q_ASSIGN U26754 ( .B(clk), .A(\g.we_clk [6020]));
Q_ASSIGN U26755 ( .B(clk), .A(\g.we_clk [6019]));
Q_ASSIGN U26756 ( .B(clk), .A(\g.we_clk [6018]));
Q_ASSIGN U26757 ( .B(clk), .A(\g.we_clk [6017]));
Q_ASSIGN U26758 ( .B(clk), .A(\g.we_clk [6016]));
Q_ASSIGN U26759 ( .B(clk), .A(\g.we_clk [6015]));
Q_ASSIGN U26760 ( .B(clk), .A(\g.we_clk [6014]));
Q_ASSIGN U26761 ( .B(clk), .A(\g.we_clk [6013]));
Q_ASSIGN U26762 ( .B(clk), .A(\g.we_clk [6012]));
Q_ASSIGN U26763 ( .B(clk), .A(\g.we_clk [6011]));
Q_ASSIGN U26764 ( .B(clk), .A(\g.we_clk [6010]));
Q_ASSIGN U26765 ( .B(clk), .A(\g.we_clk [6009]));
Q_ASSIGN U26766 ( .B(clk), .A(\g.we_clk [6008]));
Q_ASSIGN U26767 ( .B(clk), .A(\g.we_clk [6007]));
Q_ASSIGN U26768 ( .B(clk), .A(\g.we_clk [6006]));
Q_ASSIGN U26769 ( .B(clk), .A(\g.we_clk [6005]));
Q_ASSIGN U26770 ( .B(clk), .A(\g.we_clk [6004]));
Q_ASSIGN U26771 ( .B(clk), .A(\g.we_clk [6003]));
Q_ASSIGN U26772 ( .B(clk), .A(\g.we_clk [6002]));
Q_ASSIGN U26773 ( .B(clk), .A(\g.we_clk [6001]));
Q_ASSIGN U26774 ( .B(clk), .A(\g.we_clk [6000]));
Q_ASSIGN U26775 ( .B(clk), .A(\g.we_clk [5999]));
Q_ASSIGN U26776 ( .B(clk), .A(\g.we_clk [5998]));
Q_ASSIGN U26777 ( .B(clk), .A(\g.we_clk [5997]));
Q_ASSIGN U26778 ( .B(clk), .A(\g.we_clk [5996]));
Q_ASSIGN U26779 ( .B(clk), .A(\g.we_clk [5995]));
Q_ASSIGN U26780 ( .B(clk), .A(\g.we_clk [5994]));
Q_ASSIGN U26781 ( .B(clk), .A(\g.we_clk [5993]));
Q_ASSIGN U26782 ( .B(clk), .A(\g.we_clk [5992]));
Q_ASSIGN U26783 ( .B(clk), .A(\g.we_clk [5991]));
Q_ASSIGN U26784 ( .B(clk), .A(\g.we_clk [5990]));
Q_ASSIGN U26785 ( .B(clk), .A(\g.we_clk [5989]));
Q_ASSIGN U26786 ( .B(clk), .A(\g.we_clk [5988]));
Q_ASSIGN U26787 ( .B(clk), .A(\g.we_clk [5987]));
Q_ASSIGN U26788 ( .B(clk), .A(\g.we_clk [5986]));
Q_ASSIGN U26789 ( .B(clk), .A(\g.we_clk [5985]));
Q_ASSIGN U26790 ( .B(clk), .A(\g.we_clk [5984]));
Q_ASSIGN U26791 ( .B(clk), .A(\g.we_clk [5983]));
Q_ASSIGN U26792 ( .B(clk), .A(\g.we_clk [5982]));
Q_ASSIGN U26793 ( .B(clk), .A(\g.we_clk [5981]));
Q_ASSIGN U26794 ( .B(clk), .A(\g.we_clk [5980]));
Q_ASSIGN U26795 ( .B(clk), .A(\g.we_clk [5979]));
Q_ASSIGN U26796 ( .B(clk), .A(\g.we_clk [5978]));
Q_ASSIGN U26797 ( .B(clk), .A(\g.we_clk [5977]));
Q_ASSIGN U26798 ( .B(clk), .A(\g.we_clk [5976]));
Q_ASSIGN U26799 ( .B(clk), .A(\g.we_clk [5975]));
Q_ASSIGN U26800 ( .B(clk), .A(\g.we_clk [5974]));
Q_ASSIGN U26801 ( .B(clk), .A(\g.we_clk [5973]));
Q_ASSIGN U26802 ( .B(clk), .A(\g.we_clk [5972]));
Q_ASSIGN U26803 ( .B(clk), .A(\g.we_clk [5971]));
Q_ASSIGN U26804 ( .B(clk), .A(\g.we_clk [5970]));
Q_ASSIGN U26805 ( .B(clk), .A(\g.we_clk [5969]));
Q_ASSIGN U26806 ( .B(clk), .A(\g.we_clk [5968]));
Q_ASSIGN U26807 ( .B(clk), .A(\g.we_clk [5967]));
Q_ASSIGN U26808 ( .B(clk), .A(\g.we_clk [5966]));
Q_ASSIGN U26809 ( .B(clk), .A(\g.we_clk [5965]));
Q_ASSIGN U26810 ( .B(clk), .A(\g.we_clk [5964]));
Q_ASSIGN U26811 ( .B(clk), .A(\g.we_clk [5963]));
Q_ASSIGN U26812 ( .B(clk), .A(\g.we_clk [5962]));
Q_ASSIGN U26813 ( .B(clk), .A(\g.we_clk [5961]));
Q_ASSIGN U26814 ( .B(clk), .A(\g.we_clk [5960]));
Q_ASSIGN U26815 ( .B(clk), .A(\g.we_clk [5959]));
Q_ASSIGN U26816 ( .B(clk), .A(\g.we_clk [5958]));
Q_ASSIGN U26817 ( .B(clk), .A(\g.we_clk [5957]));
Q_ASSIGN U26818 ( .B(clk), .A(\g.we_clk [5956]));
Q_ASSIGN U26819 ( .B(clk), .A(\g.we_clk [5955]));
Q_ASSIGN U26820 ( .B(clk), .A(\g.we_clk [5954]));
Q_ASSIGN U26821 ( .B(clk), .A(\g.we_clk [5953]));
Q_ASSIGN U26822 ( .B(clk), .A(\g.we_clk [5952]));
Q_ASSIGN U26823 ( .B(clk), .A(\g.we_clk [5951]));
Q_ASSIGN U26824 ( .B(clk), .A(\g.we_clk [5950]));
Q_ASSIGN U26825 ( .B(clk), .A(\g.we_clk [5949]));
Q_ASSIGN U26826 ( .B(clk), .A(\g.we_clk [5948]));
Q_ASSIGN U26827 ( .B(clk), .A(\g.we_clk [5947]));
Q_ASSIGN U26828 ( .B(clk), .A(\g.we_clk [5946]));
Q_ASSIGN U26829 ( .B(clk), .A(\g.we_clk [5945]));
Q_ASSIGN U26830 ( .B(clk), .A(\g.we_clk [5944]));
Q_ASSIGN U26831 ( .B(clk), .A(\g.we_clk [5943]));
Q_ASSIGN U26832 ( .B(clk), .A(\g.we_clk [5942]));
Q_ASSIGN U26833 ( .B(clk), .A(\g.we_clk [5941]));
Q_ASSIGN U26834 ( .B(clk), .A(\g.we_clk [5940]));
Q_ASSIGN U26835 ( .B(clk), .A(\g.we_clk [5939]));
Q_ASSIGN U26836 ( .B(clk), .A(\g.we_clk [5938]));
Q_ASSIGN U26837 ( .B(clk), .A(\g.we_clk [5937]));
Q_ASSIGN U26838 ( .B(clk), .A(\g.we_clk [5936]));
Q_ASSIGN U26839 ( .B(clk), .A(\g.we_clk [5935]));
Q_ASSIGN U26840 ( .B(clk), .A(\g.we_clk [5934]));
Q_ASSIGN U26841 ( .B(clk), .A(\g.we_clk [5933]));
Q_ASSIGN U26842 ( .B(clk), .A(\g.we_clk [5932]));
Q_ASSIGN U26843 ( .B(clk), .A(\g.we_clk [5931]));
Q_ASSIGN U26844 ( .B(clk), .A(\g.we_clk [5930]));
Q_ASSIGN U26845 ( .B(clk), .A(\g.we_clk [5929]));
Q_ASSIGN U26846 ( .B(clk), .A(\g.we_clk [5928]));
Q_ASSIGN U26847 ( .B(clk), .A(\g.we_clk [5927]));
Q_ASSIGN U26848 ( .B(clk), .A(\g.we_clk [5926]));
Q_ASSIGN U26849 ( .B(clk), .A(\g.we_clk [5925]));
Q_ASSIGN U26850 ( .B(clk), .A(\g.we_clk [5924]));
Q_ASSIGN U26851 ( .B(clk), .A(\g.we_clk [5923]));
Q_ASSIGN U26852 ( .B(clk), .A(\g.we_clk [5922]));
Q_ASSIGN U26853 ( .B(clk), .A(\g.we_clk [5921]));
Q_ASSIGN U26854 ( .B(clk), .A(\g.we_clk [5920]));
Q_ASSIGN U26855 ( .B(clk), .A(\g.we_clk [5919]));
Q_ASSIGN U26856 ( .B(clk), .A(\g.we_clk [5918]));
Q_ASSIGN U26857 ( .B(clk), .A(\g.we_clk [5917]));
Q_ASSIGN U26858 ( .B(clk), .A(\g.we_clk [5916]));
Q_ASSIGN U26859 ( .B(clk), .A(\g.we_clk [5915]));
Q_ASSIGN U26860 ( .B(clk), .A(\g.we_clk [5914]));
Q_ASSIGN U26861 ( .B(clk), .A(\g.we_clk [5913]));
Q_ASSIGN U26862 ( .B(clk), .A(\g.we_clk [5912]));
Q_ASSIGN U26863 ( .B(clk), .A(\g.we_clk [5911]));
Q_ASSIGN U26864 ( .B(clk), .A(\g.we_clk [5910]));
Q_ASSIGN U26865 ( .B(clk), .A(\g.we_clk [5909]));
Q_ASSIGN U26866 ( .B(clk), .A(\g.we_clk [5908]));
Q_ASSIGN U26867 ( .B(clk), .A(\g.we_clk [5907]));
Q_ASSIGN U26868 ( .B(clk), .A(\g.we_clk [5906]));
Q_ASSIGN U26869 ( .B(clk), .A(\g.we_clk [5905]));
Q_ASSIGN U26870 ( .B(clk), .A(\g.we_clk [5904]));
Q_ASSIGN U26871 ( .B(clk), .A(\g.we_clk [5903]));
Q_ASSIGN U26872 ( .B(clk), .A(\g.we_clk [5902]));
Q_ASSIGN U26873 ( .B(clk), .A(\g.we_clk [5901]));
Q_ASSIGN U26874 ( .B(clk), .A(\g.we_clk [5900]));
Q_ASSIGN U26875 ( .B(clk), .A(\g.we_clk [5899]));
Q_ASSIGN U26876 ( .B(clk), .A(\g.we_clk [5898]));
Q_ASSIGN U26877 ( .B(clk), .A(\g.we_clk [5897]));
Q_ASSIGN U26878 ( .B(clk), .A(\g.we_clk [5896]));
Q_ASSIGN U26879 ( .B(clk), .A(\g.we_clk [5895]));
Q_ASSIGN U26880 ( .B(clk), .A(\g.we_clk [5894]));
Q_ASSIGN U26881 ( .B(clk), .A(\g.we_clk [5893]));
Q_ASSIGN U26882 ( .B(clk), .A(\g.we_clk [5892]));
Q_ASSIGN U26883 ( .B(clk), .A(\g.we_clk [5891]));
Q_ASSIGN U26884 ( .B(clk), .A(\g.we_clk [5890]));
Q_ASSIGN U26885 ( .B(clk), .A(\g.we_clk [5889]));
Q_ASSIGN U26886 ( .B(clk), .A(\g.we_clk [5888]));
Q_ASSIGN U26887 ( .B(clk), .A(\g.we_clk [5887]));
Q_ASSIGN U26888 ( .B(clk), .A(\g.we_clk [5886]));
Q_ASSIGN U26889 ( .B(clk), .A(\g.we_clk [5885]));
Q_ASSIGN U26890 ( .B(clk), .A(\g.we_clk [5884]));
Q_ASSIGN U26891 ( .B(clk), .A(\g.we_clk [5883]));
Q_ASSIGN U26892 ( .B(clk), .A(\g.we_clk [5882]));
Q_ASSIGN U26893 ( .B(clk), .A(\g.we_clk [5881]));
Q_ASSIGN U26894 ( .B(clk), .A(\g.we_clk [5880]));
Q_ASSIGN U26895 ( .B(clk), .A(\g.we_clk [5879]));
Q_ASSIGN U26896 ( .B(clk), .A(\g.we_clk [5878]));
Q_ASSIGN U26897 ( .B(clk), .A(\g.we_clk [5877]));
Q_ASSIGN U26898 ( .B(clk), .A(\g.we_clk [5876]));
Q_ASSIGN U26899 ( .B(clk), .A(\g.we_clk [5875]));
Q_ASSIGN U26900 ( .B(clk), .A(\g.we_clk [5874]));
Q_ASSIGN U26901 ( .B(clk), .A(\g.we_clk [5873]));
Q_ASSIGN U26902 ( .B(clk), .A(\g.we_clk [5872]));
Q_ASSIGN U26903 ( .B(clk), .A(\g.we_clk [5871]));
Q_ASSIGN U26904 ( .B(clk), .A(\g.we_clk [5870]));
Q_ASSIGN U26905 ( .B(clk), .A(\g.we_clk [5869]));
Q_ASSIGN U26906 ( .B(clk), .A(\g.we_clk [5868]));
Q_ASSIGN U26907 ( .B(clk), .A(\g.we_clk [5867]));
Q_ASSIGN U26908 ( .B(clk), .A(\g.we_clk [5866]));
Q_ASSIGN U26909 ( .B(clk), .A(\g.we_clk [5865]));
Q_ASSIGN U26910 ( .B(clk), .A(\g.we_clk [5864]));
Q_ASSIGN U26911 ( .B(clk), .A(\g.we_clk [5863]));
Q_ASSIGN U26912 ( .B(clk), .A(\g.we_clk [5862]));
Q_ASSIGN U26913 ( .B(clk), .A(\g.we_clk [5861]));
Q_ASSIGN U26914 ( .B(clk), .A(\g.we_clk [5860]));
Q_ASSIGN U26915 ( .B(clk), .A(\g.we_clk [5859]));
Q_ASSIGN U26916 ( .B(clk), .A(\g.we_clk [5858]));
Q_ASSIGN U26917 ( .B(clk), .A(\g.we_clk [5857]));
Q_ASSIGN U26918 ( .B(clk), .A(\g.we_clk [5856]));
Q_ASSIGN U26919 ( .B(clk), .A(\g.we_clk [5855]));
Q_ASSIGN U26920 ( .B(clk), .A(\g.we_clk [5854]));
Q_ASSIGN U26921 ( .B(clk), .A(\g.we_clk [5853]));
Q_ASSIGN U26922 ( .B(clk), .A(\g.we_clk [5852]));
Q_ASSIGN U26923 ( .B(clk), .A(\g.we_clk [5851]));
Q_ASSIGN U26924 ( .B(clk), .A(\g.we_clk [5850]));
Q_ASSIGN U26925 ( .B(clk), .A(\g.we_clk [5849]));
Q_ASSIGN U26926 ( .B(clk), .A(\g.we_clk [5848]));
Q_ASSIGN U26927 ( .B(clk), .A(\g.we_clk [5847]));
Q_ASSIGN U26928 ( .B(clk), .A(\g.we_clk [5846]));
Q_ASSIGN U26929 ( .B(clk), .A(\g.we_clk [5845]));
Q_ASSIGN U26930 ( .B(clk), .A(\g.we_clk [5844]));
Q_ASSIGN U26931 ( .B(clk), .A(\g.we_clk [5843]));
Q_ASSIGN U26932 ( .B(clk), .A(\g.we_clk [5842]));
Q_ASSIGN U26933 ( .B(clk), .A(\g.we_clk [5841]));
Q_ASSIGN U26934 ( .B(clk), .A(\g.we_clk [5840]));
Q_ASSIGN U26935 ( .B(clk), .A(\g.we_clk [5839]));
Q_ASSIGN U26936 ( .B(clk), .A(\g.we_clk [5838]));
Q_ASSIGN U26937 ( .B(clk), .A(\g.we_clk [5837]));
Q_ASSIGN U26938 ( .B(clk), .A(\g.we_clk [5836]));
Q_ASSIGN U26939 ( .B(clk), .A(\g.we_clk [5835]));
Q_ASSIGN U26940 ( .B(clk), .A(\g.we_clk [5834]));
Q_ASSIGN U26941 ( .B(clk), .A(\g.we_clk [5833]));
Q_ASSIGN U26942 ( .B(clk), .A(\g.we_clk [5832]));
Q_ASSIGN U26943 ( .B(clk), .A(\g.we_clk [5831]));
Q_ASSIGN U26944 ( .B(clk), .A(\g.we_clk [5830]));
Q_ASSIGN U26945 ( .B(clk), .A(\g.we_clk [5829]));
Q_ASSIGN U26946 ( .B(clk), .A(\g.we_clk [5828]));
Q_ASSIGN U26947 ( .B(clk), .A(\g.we_clk [5827]));
Q_ASSIGN U26948 ( .B(clk), .A(\g.we_clk [5826]));
Q_ASSIGN U26949 ( .B(clk), .A(\g.we_clk [5825]));
Q_ASSIGN U26950 ( .B(clk), .A(\g.we_clk [5824]));
Q_ASSIGN U26951 ( .B(clk), .A(\g.we_clk [5823]));
Q_ASSIGN U26952 ( .B(clk), .A(\g.we_clk [5822]));
Q_ASSIGN U26953 ( .B(clk), .A(\g.we_clk [5821]));
Q_ASSIGN U26954 ( .B(clk), .A(\g.we_clk [5820]));
Q_ASSIGN U26955 ( .B(clk), .A(\g.we_clk [5819]));
Q_ASSIGN U26956 ( .B(clk), .A(\g.we_clk [5818]));
Q_ASSIGN U26957 ( .B(clk), .A(\g.we_clk [5817]));
Q_ASSIGN U26958 ( .B(clk), .A(\g.we_clk [5816]));
Q_ASSIGN U26959 ( .B(clk), .A(\g.we_clk [5815]));
Q_ASSIGN U26960 ( .B(clk), .A(\g.we_clk [5814]));
Q_ASSIGN U26961 ( .B(clk), .A(\g.we_clk [5813]));
Q_ASSIGN U26962 ( .B(clk), .A(\g.we_clk [5812]));
Q_ASSIGN U26963 ( .B(clk), .A(\g.we_clk [5811]));
Q_ASSIGN U26964 ( .B(clk), .A(\g.we_clk [5810]));
Q_ASSIGN U26965 ( .B(clk), .A(\g.we_clk [5809]));
Q_ASSIGN U26966 ( .B(clk), .A(\g.we_clk [5808]));
Q_ASSIGN U26967 ( .B(clk), .A(\g.we_clk [5807]));
Q_ASSIGN U26968 ( .B(clk), .A(\g.we_clk [5806]));
Q_ASSIGN U26969 ( .B(clk), .A(\g.we_clk [5805]));
Q_ASSIGN U26970 ( .B(clk), .A(\g.we_clk [5804]));
Q_ASSIGN U26971 ( .B(clk), .A(\g.we_clk [5803]));
Q_ASSIGN U26972 ( .B(clk), .A(\g.we_clk [5802]));
Q_ASSIGN U26973 ( .B(clk), .A(\g.we_clk [5801]));
Q_ASSIGN U26974 ( .B(clk), .A(\g.we_clk [5800]));
Q_ASSIGN U26975 ( .B(clk), .A(\g.we_clk [5799]));
Q_ASSIGN U26976 ( .B(clk), .A(\g.we_clk [5798]));
Q_ASSIGN U26977 ( .B(clk), .A(\g.we_clk [5797]));
Q_ASSIGN U26978 ( .B(clk), .A(\g.we_clk [5796]));
Q_ASSIGN U26979 ( .B(clk), .A(\g.we_clk [5795]));
Q_ASSIGN U26980 ( .B(clk), .A(\g.we_clk [5794]));
Q_ASSIGN U26981 ( .B(clk), .A(\g.we_clk [5793]));
Q_ASSIGN U26982 ( .B(clk), .A(\g.we_clk [5792]));
Q_ASSIGN U26983 ( .B(clk), .A(\g.we_clk [5791]));
Q_ASSIGN U26984 ( .B(clk), .A(\g.we_clk [5790]));
Q_ASSIGN U26985 ( .B(clk), .A(\g.we_clk [5789]));
Q_ASSIGN U26986 ( .B(clk), .A(\g.we_clk [5788]));
Q_ASSIGN U26987 ( .B(clk), .A(\g.we_clk [5787]));
Q_ASSIGN U26988 ( .B(clk), .A(\g.we_clk [5786]));
Q_ASSIGN U26989 ( .B(clk), .A(\g.we_clk [5785]));
Q_ASSIGN U26990 ( .B(clk), .A(\g.we_clk [5784]));
Q_ASSIGN U26991 ( .B(clk), .A(\g.we_clk [5783]));
Q_ASSIGN U26992 ( .B(clk), .A(\g.we_clk [5782]));
Q_ASSIGN U26993 ( .B(clk), .A(\g.we_clk [5781]));
Q_ASSIGN U26994 ( .B(clk), .A(\g.we_clk [5780]));
Q_ASSIGN U26995 ( .B(clk), .A(\g.we_clk [5779]));
Q_ASSIGN U26996 ( .B(clk), .A(\g.we_clk [5778]));
Q_ASSIGN U26997 ( .B(clk), .A(\g.we_clk [5777]));
Q_ASSIGN U26998 ( .B(clk), .A(\g.we_clk [5776]));
Q_ASSIGN U26999 ( .B(clk), .A(\g.we_clk [5775]));
Q_ASSIGN U27000 ( .B(clk), .A(\g.we_clk [5774]));
Q_ASSIGN U27001 ( .B(clk), .A(\g.we_clk [5773]));
Q_ASSIGN U27002 ( .B(clk), .A(\g.we_clk [5772]));
Q_ASSIGN U27003 ( .B(clk), .A(\g.we_clk [5771]));
Q_ASSIGN U27004 ( .B(clk), .A(\g.we_clk [5770]));
Q_ASSIGN U27005 ( .B(clk), .A(\g.we_clk [5769]));
Q_ASSIGN U27006 ( .B(clk), .A(\g.we_clk [5768]));
Q_ASSIGN U27007 ( .B(clk), .A(\g.we_clk [5767]));
Q_ASSIGN U27008 ( .B(clk), .A(\g.we_clk [5766]));
Q_ASSIGN U27009 ( .B(clk), .A(\g.we_clk [5765]));
Q_ASSIGN U27010 ( .B(clk), .A(\g.we_clk [5764]));
Q_ASSIGN U27011 ( .B(clk), .A(\g.we_clk [5763]));
Q_ASSIGN U27012 ( .B(clk), .A(\g.we_clk [5762]));
Q_ASSIGN U27013 ( .B(clk), .A(\g.we_clk [5761]));
Q_ASSIGN U27014 ( .B(clk), .A(\g.we_clk [5760]));
Q_ASSIGN U27015 ( .B(clk), .A(\g.we_clk [5759]));
Q_ASSIGN U27016 ( .B(clk), .A(\g.we_clk [5758]));
Q_ASSIGN U27017 ( .B(clk), .A(\g.we_clk [5757]));
Q_ASSIGN U27018 ( .B(clk), .A(\g.we_clk [5756]));
Q_ASSIGN U27019 ( .B(clk), .A(\g.we_clk [5755]));
Q_ASSIGN U27020 ( .B(clk), .A(\g.we_clk [5754]));
Q_ASSIGN U27021 ( .B(clk), .A(\g.we_clk [5753]));
Q_ASSIGN U27022 ( .B(clk), .A(\g.we_clk [5752]));
Q_ASSIGN U27023 ( .B(clk), .A(\g.we_clk [5751]));
Q_ASSIGN U27024 ( .B(clk), .A(\g.we_clk [5750]));
Q_ASSIGN U27025 ( .B(clk), .A(\g.we_clk [5749]));
Q_ASSIGN U27026 ( .B(clk), .A(\g.we_clk [5748]));
Q_ASSIGN U27027 ( .B(clk), .A(\g.we_clk [5747]));
Q_ASSIGN U27028 ( .B(clk), .A(\g.we_clk [5746]));
Q_ASSIGN U27029 ( .B(clk), .A(\g.we_clk [5745]));
Q_ASSIGN U27030 ( .B(clk), .A(\g.we_clk [5744]));
Q_ASSIGN U27031 ( .B(clk), .A(\g.we_clk [5743]));
Q_ASSIGN U27032 ( .B(clk), .A(\g.we_clk [5742]));
Q_ASSIGN U27033 ( .B(clk), .A(\g.we_clk [5741]));
Q_ASSIGN U27034 ( .B(clk), .A(\g.we_clk [5740]));
Q_ASSIGN U27035 ( .B(clk), .A(\g.we_clk [5739]));
Q_ASSIGN U27036 ( .B(clk), .A(\g.we_clk [5738]));
Q_ASSIGN U27037 ( .B(clk), .A(\g.we_clk [5737]));
Q_ASSIGN U27038 ( .B(clk), .A(\g.we_clk [5736]));
Q_ASSIGN U27039 ( .B(clk), .A(\g.we_clk [5735]));
Q_ASSIGN U27040 ( .B(clk), .A(\g.we_clk [5734]));
Q_ASSIGN U27041 ( .B(clk), .A(\g.we_clk [5733]));
Q_ASSIGN U27042 ( .B(clk), .A(\g.we_clk [5732]));
Q_ASSIGN U27043 ( .B(clk), .A(\g.we_clk [5731]));
Q_ASSIGN U27044 ( .B(clk), .A(\g.we_clk [5730]));
Q_ASSIGN U27045 ( .B(clk), .A(\g.we_clk [5729]));
Q_ASSIGN U27046 ( .B(clk), .A(\g.we_clk [5728]));
Q_ASSIGN U27047 ( .B(clk), .A(\g.we_clk [5727]));
Q_ASSIGN U27048 ( .B(clk), .A(\g.we_clk [5726]));
Q_ASSIGN U27049 ( .B(clk), .A(\g.we_clk [5725]));
Q_ASSIGN U27050 ( .B(clk), .A(\g.we_clk [5724]));
Q_ASSIGN U27051 ( .B(clk), .A(\g.we_clk [5723]));
Q_ASSIGN U27052 ( .B(clk), .A(\g.we_clk [5722]));
Q_ASSIGN U27053 ( .B(clk), .A(\g.we_clk [5721]));
Q_ASSIGN U27054 ( .B(clk), .A(\g.we_clk [5720]));
Q_ASSIGN U27055 ( .B(clk), .A(\g.we_clk [5719]));
Q_ASSIGN U27056 ( .B(clk), .A(\g.we_clk [5718]));
Q_ASSIGN U27057 ( .B(clk), .A(\g.we_clk [5717]));
Q_ASSIGN U27058 ( .B(clk), .A(\g.we_clk [5716]));
Q_ASSIGN U27059 ( .B(clk), .A(\g.we_clk [5715]));
Q_ASSIGN U27060 ( .B(clk), .A(\g.we_clk [5714]));
Q_ASSIGN U27061 ( .B(clk), .A(\g.we_clk [5713]));
Q_ASSIGN U27062 ( .B(clk), .A(\g.we_clk [5712]));
Q_ASSIGN U27063 ( .B(clk), .A(\g.we_clk [5711]));
Q_ASSIGN U27064 ( .B(clk), .A(\g.we_clk [5710]));
Q_ASSIGN U27065 ( .B(clk), .A(\g.we_clk [5709]));
Q_ASSIGN U27066 ( .B(clk), .A(\g.we_clk [5708]));
Q_ASSIGN U27067 ( .B(clk), .A(\g.we_clk [5707]));
Q_ASSIGN U27068 ( .B(clk), .A(\g.we_clk [5706]));
Q_ASSIGN U27069 ( .B(clk), .A(\g.we_clk [5705]));
Q_ASSIGN U27070 ( .B(clk), .A(\g.we_clk [5704]));
Q_ASSIGN U27071 ( .B(clk), .A(\g.we_clk [5703]));
Q_ASSIGN U27072 ( .B(clk), .A(\g.we_clk [5702]));
Q_ASSIGN U27073 ( .B(clk), .A(\g.we_clk [5701]));
Q_ASSIGN U27074 ( .B(clk), .A(\g.we_clk [5700]));
Q_ASSIGN U27075 ( .B(clk), .A(\g.we_clk [5699]));
Q_ASSIGN U27076 ( .B(clk), .A(\g.we_clk [5698]));
Q_ASSIGN U27077 ( .B(clk), .A(\g.we_clk [5697]));
Q_ASSIGN U27078 ( .B(clk), .A(\g.we_clk [5696]));
Q_ASSIGN U27079 ( .B(clk), .A(\g.we_clk [5695]));
Q_ASSIGN U27080 ( .B(clk), .A(\g.we_clk [5694]));
Q_ASSIGN U27081 ( .B(clk), .A(\g.we_clk [5693]));
Q_ASSIGN U27082 ( .B(clk), .A(\g.we_clk [5692]));
Q_ASSIGN U27083 ( .B(clk), .A(\g.we_clk [5691]));
Q_ASSIGN U27084 ( .B(clk), .A(\g.we_clk [5690]));
Q_ASSIGN U27085 ( .B(clk), .A(\g.we_clk [5689]));
Q_ASSIGN U27086 ( .B(clk), .A(\g.we_clk [5688]));
Q_ASSIGN U27087 ( .B(clk), .A(\g.we_clk [5687]));
Q_ASSIGN U27088 ( .B(clk), .A(\g.we_clk [5686]));
Q_ASSIGN U27089 ( .B(clk), .A(\g.we_clk [5685]));
Q_ASSIGN U27090 ( .B(clk), .A(\g.we_clk [5684]));
Q_ASSIGN U27091 ( .B(clk), .A(\g.we_clk [5683]));
Q_ASSIGN U27092 ( .B(clk), .A(\g.we_clk [5682]));
Q_ASSIGN U27093 ( .B(clk), .A(\g.we_clk [5681]));
Q_ASSIGN U27094 ( .B(clk), .A(\g.we_clk [5680]));
Q_ASSIGN U27095 ( .B(clk), .A(\g.we_clk [5679]));
Q_ASSIGN U27096 ( .B(clk), .A(\g.we_clk [5678]));
Q_ASSIGN U27097 ( .B(clk), .A(\g.we_clk [5677]));
Q_ASSIGN U27098 ( .B(clk), .A(\g.we_clk [5676]));
Q_ASSIGN U27099 ( .B(clk), .A(\g.we_clk [5675]));
Q_ASSIGN U27100 ( .B(clk), .A(\g.we_clk [5674]));
Q_ASSIGN U27101 ( .B(clk), .A(\g.we_clk [5673]));
Q_ASSIGN U27102 ( .B(clk), .A(\g.we_clk [5672]));
Q_ASSIGN U27103 ( .B(clk), .A(\g.we_clk [5671]));
Q_ASSIGN U27104 ( .B(clk), .A(\g.we_clk [5670]));
Q_ASSIGN U27105 ( .B(clk), .A(\g.we_clk [5669]));
Q_ASSIGN U27106 ( .B(clk), .A(\g.we_clk [5668]));
Q_ASSIGN U27107 ( .B(clk), .A(\g.we_clk [5667]));
Q_ASSIGN U27108 ( .B(clk), .A(\g.we_clk [5666]));
Q_ASSIGN U27109 ( .B(clk), .A(\g.we_clk [5665]));
Q_ASSIGN U27110 ( .B(clk), .A(\g.we_clk [5664]));
Q_ASSIGN U27111 ( .B(clk), .A(\g.we_clk [5663]));
Q_ASSIGN U27112 ( .B(clk), .A(\g.we_clk [5662]));
Q_ASSIGN U27113 ( .B(clk), .A(\g.we_clk [5661]));
Q_ASSIGN U27114 ( .B(clk), .A(\g.we_clk [5660]));
Q_ASSIGN U27115 ( .B(clk), .A(\g.we_clk [5659]));
Q_ASSIGN U27116 ( .B(clk), .A(\g.we_clk [5658]));
Q_ASSIGN U27117 ( .B(clk), .A(\g.we_clk [5657]));
Q_ASSIGN U27118 ( .B(clk), .A(\g.we_clk [5656]));
Q_ASSIGN U27119 ( .B(clk), .A(\g.we_clk [5655]));
Q_ASSIGN U27120 ( .B(clk), .A(\g.we_clk [5654]));
Q_ASSIGN U27121 ( .B(clk), .A(\g.we_clk [5653]));
Q_ASSIGN U27122 ( .B(clk), .A(\g.we_clk [5652]));
Q_ASSIGN U27123 ( .B(clk), .A(\g.we_clk [5651]));
Q_ASSIGN U27124 ( .B(clk), .A(\g.we_clk [5650]));
Q_ASSIGN U27125 ( .B(clk), .A(\g.we_clk [5649]));
Q_ASSIGN U27126 ( .B(clk), .A(\g.we_clk [5648]));
Q_ASSIGN U27127 ( .B(clk), .A(\g.we_clk [5647]));
Q_ASSIGN U27128 ( .B(clk), .A(\g.we_clk [5646]));
Q_ASSIGN U27129 ( .B(clk), .A(\g.we_clk [5645]));
Q_ASSIGN U27130 ( .B(clk), .A(\g.we_clk [5644]));
Q_ASSIGN U27131 ( .B(clk), .A(\g.we_clk [5643]));
Q_ASSIGN U27132 ( .B(clk), .A(\g.we_clk [5642]));
Q_ASSIGN U27133 ( .B(clk), .A(\g.we_clk [5641]));
Q_ASSIGN U27134 ( .B(clk), .A(\g.we_clk [5640]));
Q_ASSIGN U27135 ( .B(clk), .A(\g.we_clk [5639]));
Q_ASSIGN U27136 ( .B(clk), .A(\g.we_clk [5638]));
Q_ASSIGN U27137 ( .B(clk), .A(\g.we_clk [5637]));
Q_ASSIGN U27138 ( .B(clk), .A(\g.we_clk [5636]));
Q_ASSIGN U27139 ( .B(clk), .A(\g.we_clk [5635]));
Q_ASSIGN U27140 ( .B(clk), .A(\g.we_clk [5634]));
Q_ASSIGN U27141 ( .B(clk), .A(\g.we_clk [5633]));
Q_ASSIGN U27142 ( .B(clk), .A(\g.we_clk [5632]));
Q_ASSIGN U27143 ( .B(clk), .A(\g.we_clk [5631]));
Q_ASSIGN U27144 ( .B(clk), .A(\g.we_clk [5630]));
Q_ASSIGN U27145 ( .B(clk), .A(\g.we_clk [5629]));
Q_ASSIGN U27146 ( .B(clk), .A(\g.we_clk [5628]));
Q_ASSIGN U27147 ( .B(clk), .A(\g.we_clk [5627]));
Q_ASSIGN U27148 ( .B(clk), .A(\g.we_clk [5626]));
Q_ASSIGN U27149 ( .B(clk), .A(\g.we_clk [5625]));
Q_ASSIGN U27150 ( .B(clk), .A(\g.we_clk [5624]));
Q_ASSIGN U27151 ( .B(clk), .A(\g.we_clk [5623]));
Q_ASSIGN U27152 ( .B(clk), .A(\g.we_clk [5622]));
Q_ASSIGN U27153 ( .B(clk), .A(\g.we_clk [5621]));
Q_ASSIGN U27154 ( .B(clk), .A(\g.we_clk [5620]));
Q_ASSIGN U27155 ( .B(clk), .A(\g.we_clk [5619]));
Q_ASSIGN U27156 ( .B(clk), .A(\g.we_clk [5618]));
Q_ASSIGN U27157 ( .B(clk), .A(\g.we_clk [5617]));
Q_ASSIGN U27158 ( .B(clk), .A(\g.we_clk [5616]));
Q_ASSIGN U27159 ( .B(clk), .A(\g.we_clk [5615]));
Q_ASSIGN U27160 ( .B(clk), .A(\g.we_clk [5614]));
Q_ASSIGN U27161 ( .B(clk), .A(\g.we_clk [5613]));
Q_ASSIGN U27162 ( .B(clk), .A(\g.we_clk [5612]));
Q_ASSIGN U27163 ( .B(clk), .A(\g.we_clk [5611]));
Q_ASSIGN U27164 ( .B(clk), .A(\g.we_clk [5610]));
Q_ASSIGN U27165 ( .B(clk), .A(\g.we_clk [5609]));
Q_ASSIGN U27166 ( .B(clk), .A(\g.we_clk [5608]));
Q_ASSIGN U27167 ( .B(clk), .A(\g.we_clk [5607]));
Q_ASSIGN U27168 ( .B(clk), .A(\g.we_clk [5606]));
Q_ASSIGN U27169 ( .B(clk), .A(\g.we_clk [5605]));
Q_ASSIGN U27170 ( .B(clk), .A(\g.we_clk [5604]));
Q_ASSIGN U27171 ( .B(clk), .A(\g.we_clk [5603]));
Q_ASSIGN U27172 ( .B(clk), .A(\g.we_clk [5602]));
Q_ASSIGN U27173 ( .B(clk), .A(\g.we_clk [5601]));
Q_ASSIGN U27174 ( .B(clk), .A(\g.we_clk [5600]));
Q_ASSIGN U27175 ( .B(clk), .A(\g.we_clk [5599]));
Q_ASSIGN U27176 ( .B(clk), .A(\g.we_clk [5598]));
Q_ASSIGN U27177 ( .B(clk), .A(\g.we_clk [5597]));
Q_ASSIGN U27178 ( .B(clk), .A(\g.we_clk [5596]));
Q_ASSIGN U27179 ( .B(clk), .A(\g.we_clk [5595]));
Q_ASSIGN U27180 ( .B(clk), .A(\g.we_clk [5594]));
Q_ASSIGN U27181 ( .B(clk), .A(\g.we_clk [5593]));
Q_ASSIGN U27182 ( .B(clk), .A(\g.we_clk [5592]));
Q_ASSIGN U27183 ( .B(clk), .A(\g.we_clk [5591]));
Q_ASSIGN U27184 ( .B(clk), .A(\g.we_clk [5590]));
Q_ASSIGN U27185 ( .B(clk), .A(\g.we_clk [5589]));
Q_ASSIGN U27186 ( .B(clk), .A(\g.we_clk [5588]));
Q_ASSIGN U27187 ( .B(clk), .A(\g.we_clk [5587]));
Q_ASSIGN U27188 ( .B(clk), .A(\g.we_clk [5586]));
Q_ASSIGN U27189 ( .B(clk), .A(\g.we_clk [5585]));
Q_ASSIGN U27190 ( .B(clk), .A(\g.we_clk [5584]));
Q_ASSIGN U27191 ( .B(clk), .A(\g.we_clk [5583]));
Q_ASSIGN U27192 ( .B(clk), .A(\g.we_clk [5582]));
Q_ASSIGN U27193 ( .B(clk), .A(\g.we_clk [5581]));
Q_ASSIGN U27194 ( .B(clk), .A(\g.we_clk [5580]));
Q_ASSIGN U27195 ( .B(clk), .A(\g.we_clk [5579]));
Q_ASSIGN U27196 ( .B(clk), .A(\g.we_clk [5578]));
Q_ASSIGN U27197 ( .B(clk), .A(\g.we_clk [5577]));
Q_ASSIGN U27198 ( .B(clk), .A(\g.we_clk [5576]));
Q_ASSIGN U27199 ( .B(clk), .A(\g.we_clk [5575]));
Q_ASSIGN U27200 ( .B(clk), .A(\g.we_clk [5574]));
Q_ASSIGN U27201 ( .B(clk), .A(\g.we_clk [5573]));
Q_ASSIGN U27202 ( .B(clk), .A(\g.we_clk [5572]));
Q_ASSIGN U27203 ( .B(clk), .A(\g.we_clk [5571]));
Q_ASSIGN U27204 ( .B(clk), .A(\g.we_clk [5570]));
Q_ASSIGN U27205 ( .B(clk), .A(\g.we_clk [5569]));
Q_ASSIGN U27206 ( .B(clk), .A(\g.we_clk [5568]));
Q_ASSIGN U27207 ( .B(clk), .A(\g.we_clk [5567]));
Q_ASSIGN U27208 ( .B(clk), .A(\g.we_clk [5566]));
Q_ASSIGN U27209 ( .B(clk), .A(\g.we_clk [5565]));
Q_ASSIGN U27210 ( .B(clk), .A(\g.we_clk [5564]));
Q_ASSIGN U27211 ( .B(clk), .A(\g.we_clk [5563]));
Q_ASSIGN U27212 ( .B(clk), .A(\g.we_clk [5562]));
Q_ASSIGN U27213 ( .B(clk), .A(\g.we_clk [5561]));
Q_ASSIGN U27214 ( .B(clk), .A(\g.we_clk [5560]));
Q_ASSIGN U27215 ( .B(clk), .A(\g.we_clk [5559]));
Q_ASSIGN U27216 ( .B(clk), .A(\g.we_clk [5558]));
Q_ASSIGN U27217 ( .B(clk), .A(\g.we_clk [5557]));
Q_ASSIGN U27218 ( .B(clk), .A(\g.we_clk [5556]));
Q_ASSIGN U27219 ( .B(clk), .A(\g.we_clk [5555]));
Q_ASSIGN U27220 ( .B(clk), .A(\g.we_clk [5554]));
Q_ASSIGN U27221 ( .B(clk), .A(\g.we_clk [5553]));
Q_ASSIGN U27222 ( .B(clk), .A(\g.we_clk [5552]));
Q_ASSIGN U27223 ( .B(clk), .A(\g.we_clk [5551]));
Q_ASSIGN U27224 ( .B(clk), .A(\g.we_clk [5550]));
Q_ASSIGN U27225 ( .B(clk), .A(\g.we_clk [5549]));
Q_ASSIGN U27226 ( .B(clk), .A(\g.we_clk [5548]));
Q_ASSIGN U27227 ( .B(clk), .A(\g.we_clk [5547]));
Q_ASSIGN U27228 ( .B(clk), .A(\g.we_clk [5546]));
Q_ASSIGN U27229 ( .B(clk), .A(\g.we_clk [5545]));
Q_ASSIGN U27230 ( .B(clk), .A(\g.we_clk [5544]));
Q_ASSIGN U27231 ( .B(clk), .A(\g.we_clk [5543]));
Q_ASSIGN U27232 ( .B(clk), .A(\g.we_clk [5542]));
Q_ASSIGN U27233 ( .B(clk), .A(\g.we_clk [5541]));
Q_ASSIGN U27234 ( .B(clk), .A(\g.we_clk [5540]));
Q_ASSIGN U27235 ( .B(clk), .A(\g.we_clk [5539]));
Q_ASSIGN U27236 ( .B(clk), .A(\g.we_clk [5538]));
Q_ASSIGN U27237 ( .B(clk), .A(\g.we_clk [5537]));
Q_ASSIGN U27238 ( .B(clk), .A(\g.we_clk [5536]));
Q_ASSIGN U27239 ( .B(clk), .A(\g.we_clk [5535]));
Q_ASSIGN U27240 ( .B(clk), .A(\g.we_clk [5534]));
Q_ASSIGN U27241 ( .B(clk), .A(\g.we_clk [5533]));
Q_ASSIGN U27242 ( .B(clk), .A(\g.we_clk [5532]));
Q_ASSIGN U27243 ( .B(clk), .A(\g.we_clk [5531]));
Q_ASSIGN U27244 ( .B(clk), .A(\g.we_clk [5530]));
Q_ASSIGN U27245 ( .B(clk), .A(\g.we_clk [5529]));
Q_ASSIGN U27246 ( .B(clk), .A(\g.we_clk [5528]));
Q_ASSIGN U27247 ( .B(clk), .A(\g.we_clk [5527]));
Q_ASSIGN U27248 ( .B(clk), .A(\g.we_clk [5526]));
Q_ASSIGN U27249 ( .B(clk), .A(\g.we_clk [5525]));
Q_ASSIGN U27250 ( .B(clk), .A(\g.we_clk [5524]));
Q_ASSIGN U27251 ( .B(clk), .A(\g.we_clk [5523]));
Q_ASSIGN U27252 ( .B(clk), .A(\g.we_clk [5522]));
Q_ASSIGN U27253 ( .B(clk), .A(\g.we_clk [5521]));
Q_ASSIGN U27254 ( .B(clk), .A(\g.we_clk [5520]));
Q_ASSIGN U27255 ( .B(clk), .A(\g.we_clk [5519]));
Q_ASSIGN U27256 ( .B(clk), .A(\g.we_clk [5518]));
Q_ASSIGN U27257 ( .B(clk), .A(\g.we_clk [5517]));
Q_ASSIGN U27258 ( .B(clk), .A(\g.we_clk [5516]));
Q_ASSIGN U27259 ( .B(clk), .A(\g.we_clk [5515]));
Q_ASSIGN U27260 ( .B(clk), .A(\g.we_clk [5514]));
Q_ASSIGN U27261 ( .B(clk), .A(\g.we_clk [5513]));
Q_ASSIGN U27262 ( .B(clk), .A(\g.we_clk [5512]));
Q_ASSIGN U27263 ( .B(clk), .A(\g.we_clk [5511]));
Q_ASSIGN U27264 ( .B(clk), .A(\g.we_clk [5510]));
Q_ASSIGN U27265 ( .B(clk), .A(\g.we_clk [5509]));
Q_ASSIGN U27266 ( .B(clk), .A(\g.we_clk [5508]));
Q_ASSIGN U27267 ( .B(clk), .A(\g.we_clk [5507]));
Q_ASSIGN U27268 ( .B(clk), .A(\g.we_clk [5506]));
Q_ASSIGN U27269 ( .B(clk), .A(\g.we_clk [5505]));
Q_ASSIGN U27270 ( .B(clk), .A(\g.we_clk [5504]));
Q_ASSIGN U27271 ( .B(clk), .A(\g.we_clk [5503]));
Q_ASSIGN U27272 ( .B(clk), .A(\g.we_clk [5502]));
Q_ASSIGN U27273 ( .B(clk), .A(\g.we_clk [5501]));
Q_ASSIGN U27274 ( .B(clk), .A(\g.we_clk [5500]));
Q_ASSIGN U27275 ( .B(clk), .A(\g.we_clk [5499]));
Q_ASSIGN U27276 ( .B(clk), .A(\g.we_clk [5498]));
Q_ASSIGN U27277 ( .B(clk), .A(\g.we_clk [5497]));
Q_ASSIGN U27278 ( .B(clk), .A(\g.we_clk [5496]));
Q_ASSIGN U27279 ( .B(clk), .A(\g.we_clk [5495]));
Q_ASSIGN U27280 ( .B(clk), .A(\g.we_clk [5494]));
Q_ASSIGN U27281 ( .B(clk), .A(\g.we_clk [5493]));
Q_ASSIGN U27282 ( .B(clk), .A(\g.we_clk [5492]));
Q_ASSIGN U27283 ( .B(clk), .A(\g.we_clk [5491]));
Q_ASSIGN U27284 ( .B(clk), .A(\g.we_clk [5490]));
Q_ASSIGN U27285 ( .B(clk), .A(\g.we_clk [5489]));
Q_ASSIGN U27286 ( .B(clk), .A(\g.we_clk [5488]));
Q_ASSIGN U27287 ( .B(clk), .A(\g.we_clk [5487]));
Q_ASSIGN U27288 ( .B(clk), .A(\g.we_clk [5486]));
Q_ASSIGN U27289 ( .B(clk), .A(\g.we_clk [5485]));
Q_ASSIGN U27290 ( .B(clk), .A(\g.we_clk [5484]));
Q_ASSIGN U27291 ( .B(clk), .A(\g.we_clk [5483]));
Q_ASSIGN U27292 ( .B(clk), .A(\g.we_clk [5482]));
Q_ASSIGN U27293 ( .B(clk), .A(\g.we_clk [5481]));
Q_ASSIGN U27294 ( .B(clk), .A(\g.we_clk [5480]));
Q_ASSIGN U27295 ( .B(clk), .A(\g.we_clk [5479]));
Q_ASSIGN U27296 ( .B(clk), .A(\g.we_clk [5478]));
Q_ASSIGN U27297 ( .B(clk), .A(\g.we_clk [5477]));
Q_ASSIGN U27298 ( .B(clk), .A(\g.we_clk [5476]));
Q_ASSIGN U27299 ( .B(clk), .A(\g.we_clk [5475]));
Q_ASSIGN U27300 ( .B(clk), .A(\g.we_clk [5474]));
Q_ASSIGN U27301 ( .B(clk), .A(\g.we_clk [5473]));
Q_ASSIGN U27302 ( .B(clk), .A(\g.we_clk [5472]));
Q_ASSIGN U27303 ( .B(clk), .A(\g.we_clk [5471]));
Q_ASSIGN U27304 ( .B(clk), .A(\g.we_clk [5470]));
Q_ASSIGN U27305 ( .B(clk), .A(\g.we_clk [5469]));
Q_ASSIGN U27306 ( .B(clk), .A(\g.we_clk [5468]));
Q_ASSIGN U27307 ( .B(clk), .A(\g.we_clk [5467]));
Q_ASSIGN U27308 ( .B(clk), .A(\g.we_clk [5466]));
Q_ASSIGN U27309 ( .B(clk), .A(\g.we_clk [5465]));
Q_ASSIGN U27310 ( .B(clk), .A(\g.we_clk [5464]));
Q_ASSIGN U27311 ( .B(clk), .A(\g.we_clk [5463]));
Q_ASSIGN U27312 ( .B(clk), .A(\g.we_clk [5462]));
Q_ASSIGN U27313 ( .B(clk), .A(\g.we_clk [5461]));
Q_ASSIGN U27314 ( .B(clk), .A(\g.we_clk [5460]));
Q_ASSIGN U27315 ( .B(clk), .A(\g.we_clk [5459]));
Q_ASSIGN U27316 ( .B(clk), .A(\g.we_clk [5458]));
Q_ASSIGN U27317 ( .B(clk), .A(\g.we_clk [5457]));
Q_ASSIGN U27318 ( .B(clk), .A(\g.we_clk [5456]));
Q_ASSIGN U27319 ( .B(clk), .A(\g.we_clk [5455]));
Q_ASSIGN U27320 ( .B(clk), .A(\g.we_clk [5454]));
Q_ASSIGN U27321 ( .B(clk), .A(\g.we_clk [5453]));
Q_ASSIGN U27322 ( .B(clk), .A(\g.we_clk [5452]));
Q_ASSIGN U27323 ( .B(clk), .A(\g.we_clk [5451]));
Q_ASSIGN U27324 ( .B(clk), .A(\g.we_clk [5450]));
Q_ASSIGN U27325 ( .B(clk), .A(\g.we_clk [5449]));
Q_ASSIGN U27326 ( .B(clk), .A(\g.we_clk [5448]));
Q_ASSIGN U27327 ( .B(clk), .A(\g.we_clk [5447]));
Q_ASSIGN U27328 ( .B(clk), .A(\g.we_clk [5446]));
Q_ASSIGN U27329 ( .B(clk), .A(\g.we_clk [5445]));
Q_ASSIGN U27330 ( .B(clk), .A(\g.we_clk [5444]));
Q_ASSIGN U27331 ( .B(clk), .A(\g.we_clk [5443]));
Q_ASSIGN U27332 ( .B(clk), .A(\g.we_clk [5442]));
Q_ASSIGN U27333 ( .B(clk), .A(\g.we_clk [5441]));
Q_ASSIGN U27334 ( .B(clk), .A(\g.we_clk [5440]));
Q_ASSIGN U27335 ( .B(clk), .A(\g.we_clk [5439]));
Q_ASSIGN U27336 ( .B(clk), .A(\g.we_clk [5438]));
Q_ASSIGN U27337 ( .B(clk), .A(\g.we_clk [5437]));
Q_ASSIGN U27338 ( .B(clk), .A(\g.we_clk [5436]));
Q_ASSIGN U27339 ( .B(clk), .A(\g.we_clk [5435]));
Q_ASSIGN U27340 ( .B(clk), .A(\g.we_clk [5434]));
Q_ASSIGN U27341 ( .B(clk), .A(\g.we_clk [5433]));
Q_ASSIGN U27342 ( .B(clk), .A(\g.we_clk [5432]));
Q_ASSIGN U27343 ( .B(clk), .A(\g.we_clk [5431]));
Q_ASSIGN U27344 ( .B(clk), .A(\g.we_clk [5430]));
Q_ASSIGN U27345 ( .B(clk), .A(\g.we_clk [5429]));
Q_ASSIGN U27346 ( .B(clk), .A(\g.we_clk [5428]));
Q_ASSIGN U27347 ( .B(clk), .A(\g.we_clk [5427]));
Q_ASSIGN U27348 ( .B(clk), .A(\g.we_clk [5426]));
Q_ASSIGN U27349 ( .B(clk), .A(\g.we_clk [5425]));
Q_ASSIGN U27350 ( .B(clk), .A(\g.we_clk [5424]));
Q_ASSIGN U27351 ( .B(clk), .A(\g.we_clk [5423]));
Q_ASSIGN U27352 ( .B(clk), .A(\g.we_clk [5422]));
Q_ASSIGN U27353 ( .B(clk), .A(\g.we_clk [5421]));
Q_ASSIGN U27354 ( .B(clk), .A(\g.we_clk [5420]));
Q_ASSIGN U27355 ( .B(clk), .A(\g.we_clk [5419]));
Q_ASSIGN U27356 ( .B(clk), .A(\g.we_clk [5418]));
Q_ASSIGN U27357 ( .B(clk), .A(\g.we_clk [5417]));
Q_ASSIGN U27358 ( .B(clk), .A(\g.we_clk [5416]));
Q_ASSIGN U27359 ( .B(clk), .A(\g.we_clk [5415]));
Q_ASSIGN U27360 ( .B(clk), .A(\g.we_clk [5414]));
Q_ASSIGN U27361 ( .B(clk), .A(\g.we_clk [5413]));
Q_ASSIGN U27362 ( .B(clk), .A(\g.we_clk [5412]));
Q_ASSIGN U27363 ( .B(clk), .A(\g.we_clk [5411]));
Q_ASSIGN U27364 ( .B(clk), .A(\g.we_clk [5410]));
Q_ASSIGN U27365 ( .B(clk), .A(\g.we_clk [5409]));
Q_ASSIGN U27366 ( .B(clk), .A(\g.we_clk [5408]));
Q_ASSIGN U27367 ( .B(clk), .A(\g.we_clk [5407]));
Q_ASSIGN U27368 ( .B(clk), .A(\g.we_clk [5406]));
Q_ASSIGN U27369 ( .B(clk), .A(\g.we_clk [5405]));
Q_ASSIGN U27370 ( .B(clk), .A(\g.we_clk [5404]));
Q_ASSIGN U27371 ( .B(clk), .A(\g.we_clk [5403]));
Q_ASSIGN U27372 ( .B(clk), .A(\g.we_clk [5402]));
Q_ASSIGN U27373 ( .B(clk), .A(\g.we_clk [5401]));
Q_ASSIGN U27374 ( .B(clk), .A(\g.we_clk [5400]));
Q_ASSIGN U27375 ( .B(clk), .A(\g.we_clk [5399]));
Q_ASSIGN U27376 ( .B(clk), .A(\g.we_clk [5398]));
Q_ASSIGN U27377 ( .B(clk), .A(\g.we_clk [5397]));
Q_ASSIGN U27378 ( .B(clk), .A(\g.we_clk [5396]));
Q_ASSIGN U27379 ( .B(clk), .A(\g.we_clk [5395]));
Q_ASSIGN U27380 ( .B(clk), .A(\g.we_clk [5394]));
Q_ASSIGN U27381 ( .B(clk), .A(\g.we_clk [5393]));
Q_ASSIGN U27382 ( .B(clk), .A(\g.we_clk [5392]));
Q_ASSIGN U27383 ( .B(clk), .A(\g.we_clk [5391]));
Q_ASSIGN U27384 ( .B(clk), .A(\g.we_clk [5390]));
Q_ASSIGN U27385 ( .B(clk), .A(\g.we_clk [5389]));
Q_ASSIGN U27386 ( .B(clk), .A(\g.we_clk [5388]));
Q_ASSIGN U27387 ( .B(clk), .A(\g.we_clk [5387]));
Q_ASSIGN U27388 ( .B(clk), .A(\g.we_clk [5386]));
Q_ASSIGN U27389 ( .B(clk), .A(\g.we_clk [5385]));
Q_ASSIGN U27390 ( .B(clk), .A(\g.we_clk [5384]));
Q_ASSIGN U27391 ( .B(clk), .A(\g.we_clk [5383]));
Q_ASSIGN U27392 ( .B(clk), .A(\g.we_clk [5382]));
Q_ASSIGN U27393 ( .B(clk), .A(\g.we_clk [5381]));
Q_ASSIGN U27394 ( .B(clk), .A(\g.we_clk [5380]));
Q_ASSIGN U27395 ( .B(clk), .A(\g.we_clk [5379]));
Q_ASSIGN U27396 ( .B(clk), .A(\g.we_clk [5378]));
Q_ASSIGN U27397 ( .B(clk), .A(\g.we_clk [5377]));
Q_ASSIGN U27398 ( .B(clk), .A(\g.we_clk [5376]));
Q_ASSIGN U27399 ( .B(clk), .A(\g.we_clk [5375]));
Q_ASSIGN U27400 ( .B(clk), .A(\g.we_clk [5374]));
Q_ASSIGN U27401 ( .B(clk), .A(\g.we_clk [5373]));
Q_ASSIGN U27402 ( .B(clk), .A(\g.we_clk [5372]));
Q_ASSIGN U27403 ( .B(clk), .A(\g.we_clk [5371]));
Q_ASSIGN U27404 ( .B(clk), .A(\g.we_clk [5370]));
Q_ASSIGN U27405 ( .B(clk), .A(\g.we_clk [5369]));
Q_ASSIGN U27406 ( .B(clk), .A(\g.we_clk [5368]));
Q_ASSIGN U27407 ( .B(clk), .A(\g.we_clk [5367]));
Q_ASSIGN U27408 ( .B(clk), .A(\g.we_clk [5366]));
Q_ASSIGN U27409 ( .B(clk), .A(\g.we_clk [5365]));
Q_ASSIGN U27410 ( .B(clk), .A(\g.we_clk [5364]));
Q_ASSIGN U27411 ( .B(clk), .A(\g.we_clk [5363]));
Q_ASSIGN U27412 ( .B(clk), .A(\g.we_clk [5362]));
Q_ASSIGN U27413 ( .B(clk), .A(\g.we_clk [5361]));
Q_ASSIGN U27414 ( .B(clk), .A(\g.we_clk [5360]));
Q_ASSIGN U27415 ( .B(clk), .A(\g.we_clk [5359]));
Q_ASSIGN U27416 ( .B(clk), .A(\g.we_clk [5358]));
Q_ASSIGN U27417 ( .B(clk), .A(\g.we_clk [5357]));
Q_ASSIGN U27418 ( .B(clk), .A(\g.we_clk [5356]));
Q_ASSIGN U27419 ( .B(clk), .A(\g.we_clk [5355]));
Q_ASSIGN U27420 ( .B(clk), .A(\g.we_clk [5354]));
Q_ASSIGN U27421 ( .B(clk), .A(\g.we_clk [5353]));
Q_ASSIGN U27422 ( .B(clk), .A(\g.we_clk [5352]));
Q_ASSIGN U27423 ( .B(clk), .A(\g.we_clk [5351]));
Q_ASSIGN U27424 ( .B(clk), .A(\g.we_clk [5350]));
Q_ASSIGN U27425 ( .B(clk), .A(\g.we_clk [5349]));
Q_ASSIGN U27426 ( .B(clk), .A(\g.we_clk [5348]));
Q_ASSIGN U27427 ( .B(clk), .A(\g.we_clk [5347]));
Q_ASSIGN U27428 ( .B(clk), .A(\g.we_clk [5346]));
Q_ASSIGN U27429 ( .B(clk), .A(\g.we_clk [5345]));
Q_ASSIGN U27430 ( .B(clk), .A(\g.we_clk [5344]));
Q_ASSIGN U27431 ( .B(clk), .A(\g.we_clk [5343]));
Q_ASSIGN U27432 ( .B(clk), .A(\g.we_clk [5342]));
Q_ASSIGN U27433 ( .B(clk), .A(\g.we_clk [5341]));
Q_ASSIGN U27434 ( .B(clk), .A(\g.we_clk [5340]));
Q_ASSIGN U27435 ( .B(clk), .A(\g.we_clk [5339]));
Q_ASSIGN U27436 ( .B(clk), .A(\g.we_clk [5338]));
Q_ASSIGN U27437 ( .B(clk), .A(\g.we_clk [5337]));
Q_ASSIGN U27438 ( .B(clk), .A(\g.we_clk [5336]));
Q_ASSIGN U27439 ( .B(clk), .A(\g.we_clk [5335]));
Q_ASSIGN U27440 ( .B(clk), .A(\g.we_clk [5334]));
Q_ASSIGN U27441 ( .B(clk), .A(\g.we_clk [5333]));
Q_ASSIGN U27442 ( .B(clk), .A(\g.we_clk [5332]));
Q_ASSIGN U27443 ( .B(clk), .A(\g.we_clk [5331]));
Q_ASSIGN U27444 ( .B(clk), .A(\g.we_clk [5330]));
Q_ASSIGN U27445 ( .B(clk), .A(\g.we_clk [5329]));
Q_ASSIGN U27446 ( .B(clk), .A(\g.we_clk [5328]));
Q_ASSIGN U27447 ( .B(clk), .A(\g.we_clk [5327]));
Q_ASSIGN U27448 ( .B(clk), .A(\g.we_clk [5326]));
Q_ASSIGN U27449 ( .B(clk), .A(\g.we_clk [5325]));
Q_ASSIGN U27450 ( .B(clk), .A(\g.we_clk [5324]));
Q_ASSIGN U27451 ( .B(clk), .A(\g.we_clk [5323]));
Q_ASSIGN U27452 ( .B(clk), .A(\g.we_clk [5322]));
Q_ASSIGN U27453 ( .B(clk), .A(\g.we_clk [5321]));
Q_ASSIGN U27454 ( .B(clk), .A(\g.we_clk [5320]));
Q_ASSIGN U27455 ( .B(clk), .A(\g.we_clk [5319]));
Q_ASSIGN U27456 ( .B(clk), .A(\g.we_clk [5318]));
Q_ASSIGN U27457 ( .B(clk), .A(\g.we_clk [5317]));
Q_ASSIGN U27458 ( .B(clk), .A(\g.we_clk [5316]));
Q_ASSIGN U27459 ( .B(clk), .A(\g.we_clk [5315]));
Q_ASSIGN U27460 ( .B(clk), .A(\g.we_clk [5314]));
Q_ASSIGN U27461 ( .B(clk), .A(\g.we_clk [5313]));
Q_ASSIGN U27462 ( .B(clk), .A(\g.we_clk [5312]));
Q_ASSIGN U27463 ( .B(clk), .A(\g.we_clk [5311]));
Q_ASSIGN U27464 ( .B(clk), .A(\g.we_clk [5310]));
Q_ASSIGN U27465 ( .B(clk), .A(\g.we_clk [5309]));
Q_ASSIGN U27466 ( .B(clk), .A(\g.we_clk [5308]));
Q_ASSIGN U27467 ( .B(clk), .A(\g.we_clk [5307]));
Q_ASSIGN U27468 ( .B(clk), .A(\g.we_clk [5306]));
Q_ASSIGN U27469 ( .B(clk), .A(\g.we_clk [5305]));
Q_ASSIGN U27470 ( .B(clk), .A(\g.we_clk [5304]));
Q_ASSIGN U27471 ( .B(clk), .A(\g.we_clk [5303]));
Q_ASSIGN U27472 ( .B(clk), .A(\g.we_clk [5302]));
Q_ASSIGN U27473 ( .B(clk), .A(\g.we_clk [5301]));
Q_ASSIGN U27474 ( .B(clk), .A(\g.we_clk [5300]));
Q_ASSIGN U27475 ( .B(clk), .A(\g.we_clk [5299]));
Q_ASSIGN U27476 ( .B(clk), .A(\g.we_clk [5298]));
Q_ASSIGN U27477 ( .B(clk), .A(\g.we_clk [5297]));
Q_ASSIGN U27478 ( .B(clk), .A(\g.we_clk [5296]));
Q_ASSIGN U27479 ( .B(clk), .A(\g.we_clk [5295]));
Q_ASSIGN U27480 ( .B(clk), .A(\g.we_clk [5294]));
Q_ASSIGN U27481 ( .B(clk), .A(\g.we_clk [5293]));
Q_ASSIGN U27482 ( .B(clk), .A(\g.we_clk [5292]));
Q_ASSIGN U27483 ( .B(clk), .A(\g.we_clk [5291]));
Q_ASSIGN U27484 ( .B(clk), .A(\g.we_clk [5290]));
Q_ASSIGN U27485 ( .B(clk), .A(\g.we_clk [5289]));
Q_ASSIGN U27486 ( .B(clk), .A(\g.we_clk [5288]));
Q_ASSIGN U27487 ( .B(clk), .A(\g.we_clk [5287]));
Q_ASSIGN U27488 ( .B(clk), .A(\g.we_clk [5286]));
Q_ASSIGN U27489 ( .B(clk), .A(\g.we_clk [5285]));
Q_ASSIGN U27490 ( .B(clk), .A(\g.we_clk [5284]));
Q_ASSIGN U27491 ( .B(clk), .A(\g.we_clk [5283]));
Q_ASSIGN U27492 ( .B(clk), .A(\g.we_clk [5282]));
Q_ASSIGN U27493 ( .B(clk), .A(\g.we_clk [5281]));
Q_ASSIGN U27494 ( .B(clk), .A(\g.we_clk [5280]));
Q_ASSIGN U27495 ( .B(clk), .A(\g.we_clk [5279]));
Q_ASSIGN U27496 ( .B(clk), .A(\g.we_clk [5278]));
Q_ASSIGN U27497 ( .B(clk), .A(\g.we_clk [5277]));
Q_ASSIGN U27498 ( .B(clk), .A(\g.we_clk [5276]));
Q_ASSIGN U27499 ( .B(clk), .A(\g.we_clk [5275]));
Q_ASSIGN U27500 ( .B(clk), .A(\g.we_clk [5274]));
Q_ASSIGN U27501 ( .B(clk), .A(\g.we_clk [5273]));
Q_ASSIGN U27502 ( .B(clk), .A(\g.we_clk [5272]));
Q_ASSIGN U27503 ( .B(clk), .A(\g.we_clk [5271]));
Q_ASSIGN U27504 ( .B(clk), .A(\g.we_clk [5270]));
Q_ASSIGN U27505 ( .B(clk), .A(\g.we_clk [5269]));
Q_ASSIGN U27506 ( .B(clk), .A(\g.we_clk [5268]));
Q_ASSIGN U27507 ( .B(clk), .A(\g.we_clk [5267]));
Q_ASSIGN U27508 ( .B(clk), .A(\g.we_clk [5266]));
Q_ASSIGN U27509 ( .B(clk), .A(\g.we_clk [5265]));
Q_ASSIGN U27510 ( .B(clk), .A(\g.we_clk [5264]));
Q_ASSIGN U27511 ( .B(clk), .A(\g.we_clk [5263]));
Q_ASSIGN U27512 ( .B(clk), .A(\g.we_clk [5262]));
Q_ASSIGN U27513 ( .B(clk), .A(\g.we_clk [5261]));
Q_ASSIGN U27514 ( .B(clk), .A(\g.we_clk [5260]));
Q_ASSIGN U27515 ( .B(clk), .A(\g.we_clk [5259]));
Q_ASSIGN U27516 ( .B(clk), .A(\g.we_clk [5258]));
Q_ASSIGN U27517 ( .B(clk), .A(\g.we_clk [5257]));
Q_ASSIGN U27518 ( .B(clk), .A(\g.we_clk [5256]));
Q_ASSIGN U27519 ( .B(clk), .A(\g.we_clk [5255]));
Q_ASSIGN U27520 ( .B(clk), .A(\g.we_clk [5254]));
Q_ASSIGN U27521 ( .B(clk), .A(\g.we_clk [5253]));
Q_ASSIGN U27522 ( .B(clk), .A(\g.we_clk [5252]));
Q_ASSIGN U27523 ( .B(clk), .A(\g.we_clk [5251]));
Q_ASSIGN U27524 ( .B(clk), .A(\g.we_clk [5250]));
Q_ASSIGN U27525 ( .B(clk), .A(\g.we_clk [5249]));
Q_ASSIGN U27526 ( .B(clk), .A(\g.we_clk [5248]));
Q_ASSIGN U27527 ( .B(clk), .A(\g.we_clk [5247]));
Q_ASSIGN U27528 ( .B(clk), .A(\g.we_clk [5246]));
Q_ASSIGN U27529 ( .B(clk), .A(\g.we_clk [5245]));
Q_ASSIGN U27530 ( .B(clk), .A(\g.we_clk [5244]));
Q_ASSIGN U27531 ( .B(clk), .A(\g.we_clk [5243]));
Q_ASSIGN U27532 ( .B(clk), .A(\g.we_clk [5242]));
Q_ASSIGN U27533 ( .B(clk), .A(\g.we_clk [5241]));
Q_ASSIGN U27534 ( .B(clk), .A(\g.we_clk [5240]));
Q_ASSIGN U27535 ( .B(clk), .A(\g.we_clk [5239]));
Q_ASSIGN U27536 ( .B(clk), .A(\g.we_clk [5238]));
Q_ASSIGN U27537 ( .B(clk), .A(\g.we_clk [5237]));
Q_ASSIGN U27538 ( .B(clk), .A(\g.we_clk [5236]));
Q_ASSIGN U27539 ( .B(clk), .A(\g.we_clk [5235]));
Q_ASSIGN U27540 ( .B(clk), .A(\g.we_clk [5234]));
Q_ASSIGN U27541 ( .B(clk), .A(\g.we_clk [5233]));
Q_ASSIGN U27542 ( .B(clk), .A(\g.we_clk [5232]));
Q_ASSIGN U27543 ( .B(clk), .A(\g.we_clk [5231]));
Q_ASSIGN U27544 ( .B(clk), .A(\g.we_clk [5230]));
Q_ASSIGN U27545 ( .B(clk), .A(\g.we_clk [5229]));
Q_ASSIGN U27546 ( .B(clk), .A(\g.we_clk [5228]));
Q_ASSIGN U27547 ( .B(clk), .A(\g.we_clk [5227]));
Q_ASSIGN U27548 ( .B(clk), .A(\g.we_clk [5226]));
Q_ASSIGN U27549 ( .B(clk), .A(\g.we_clk [5225]));
Q_ASSIGN U27550 ( .B(clk), .A(\g.we_clk [5224]));
Q_ASSIGN U27551 ( .B(clk), .A(\g.we_clk [5223]));
Q_ASSIGN U27552 ( .B(clk), .A(\g.we_clk [5222]));
Q_ASSIGN U27553 ( .B(clk), .A(\g.we_clk [5221]));
Q_ASSIGN U27554 ( .B(clk), .A(\g.we_clk [5220]));
Q_ASSIGN U27555 ( .B(clk), .A(\g.we_clk [5219]));
Q_ASSIGN U27556 ( .B(clk), .A(\g.we_clk [5218]));
Q_ASSIGN U27557 ( .B(clk), .A(\g.we_clk [5217]));
Q_ASSIGN U27558 ( .B(clk), .A(\g.we_clk [5216]));
Q_ASSIGN U27559 ( .B(clk), .A(\g.we_clk [5215]));
Q_ASSIGN U27560 ( .B(clk), .A(\g.we_clk [5214]));
Q_ASSIGN U27561 ( .B(clk), .A(\g.we_clk [5213]));
Q_ASSIGN U27562 ( .B(clk), .A(\g.we_clk [5212]));
Q_ASSIGN U27563 ( .B(clk), .A(\g.we_clk [5211]));
Q_ASSIGN U27564 ( .B(clk), .A(\g.we_clk [5210]));
Q_ASSIGN U27565 ( .B(clk), .A(\g.we_clk [5209]));
Q_ASSIGN U27566 ( .B(clk), .A(\g.we_clk [5208]));
Q_ASSIGN U27567 ( .B(clk), .A(\g.we_clk [5207]));
Q_ASSIGN U27568 ( .B(clk), .A(\g.we_clk [5206]));
Q_ASSIGN U27569 ( .B(clk), .A(\g.we_clk [5205]));
Q_ASSIGN U27570 ( .B(clk), .A(\g.we_clk [5204]));
Q_ASSIGN U27571 ( .B(clk), .A(\g.we_clk [5203]));
Q_ASSIGN U27572 ( .B(clk), .A(\g.we_clk [5202]));
Q_ASSIGN U27573 ( .B(clk), .A(\g.we_clk [5201]));
Q_ASSIGN U27574 ( .B(clk), .A(\g.we_clk [5200]));
Q_ASSIGN U27575 ( .B(clk), .A(\g.we_clk [5199]));
Q_ASSIGN U27576 ( .B(clk), .A(\g.we_clk [5198]));
Q_ASSIGN U27577 ( .B(clk), .A(\g.we_clk [5197]));
Q_ASSIGN U27578 ( .B(clk), .A(\g.we_clk [5196]));
Q_ASSIGN U27579 ( .B(clk), .A(\g.we_clk [5195]));
Q_ASSIGN U27580 ( .B(clk), .A(\g.we_clk [5194]));
Q_ASSIGN U27581 ( .B(clk), .A(\g.we_clk [5193]));
Q_ASSIGN U27582 ( .B(clk), .A(\g.we_clk [5192]));
Q_ASSIGN U27583 ( .B(clk), .A(\g.we_clk [5191]));
Q_ASSIGN U27584 ( .B(clk), .A(\g.we_clk [5190]));
Q_ASSIGN U27585 ( .B(clk), .A(\g.we_clk [5189]));
Q_ASSIGN U27586 ( .B(clk), .A(\g.we_clk [5188]));
Q_ASSIGN U27587 ( .B(clk), .A(\g.we_clk [5187]));
Q_ASSIGN U27588 ( .B(clk), .A(\g.we_clk [5186]));
Q_ASSIGN U27589 ( .B(clk), .A(\g.we_clk [5185]));
Q_ASSIGN U27590 ( .B(clk), .A(\g.we_clk [5184]));
Q_ASSIGN U27591 ( .B(clk), .A(\g.we_clk [5183]));
Q_ASSIGN U27592 ( .B(clk), .A(\g.we_clk [5182]));
Q_ASSIGN U27593 ( .B(clk), .A(\g.we_clk [5181]));
Q_ASSIGN U27594 ( .B(clk), .A(\g.we_clk [5180]));
Q_ASSIGN U27595 ( .B(clk), .A(\g.we_clk [5179]));
Q_ASSIGN U27596 ( .B(clk), .A(\g.we_clk [5178]));
Q_ASSIGN U27597 ( .B(clk), .A(\g.we_clk [5177]));
Q_ASSIGN U27598 ( .B(clk), .A(\g.we_clk [5176]));
Q_ASSIGN U27599 ( .B(clk), .A(\g.we_clk [5175]));
Q_ASSIGN U27600 ( .B(clk), .A(\g.we_clk [5174]));
Q_ASSIGN U27601 ( .B(clk), .A(\g.we_clk [5173]));
Q_ASSIGN U27602 ( .B(clk), .A(\g.we_clk [5172]));
Q_ASSIGN U27603 ( .B(clk), .A(\g.we_clk [5171]));
Q_ASSIGN U27604 ( .B(clk), .A(\g.we_clk [5170]));
Q_ASSIGN U27605 ( .B(clk), .A(\g.we_clk [5169]));
Q_ASSIGN U27606 ( .B(clk), .A(\g.we_clk [5168]));
Q_ASSIGN U27607 ( .B(clk), .A(\g.we_clk [5167]));
Q_ASSIGN U27608 ( .B(clk), .A(\g.we_clk [5166]));
Q_ASSIGN U27609 ( .B(clk), .A(\g.we_clk [5165]));
Q_ASSIGN U27610 ( .B(clk), .A(\g.we_clk [5164]));
Q_ASSIGN U27611 ( .B(clk), .A(\g.we_clk [5163]));
Q_ASSIGN U27612 ( .B(clk), .A(\g.we_clk [5162]));
Q_ASSIGN U27613 ( .B(clk), .A(\g.we_clk [5161]));
Q_ASSIGN U27614 ( .B(clk), .A(\g.we_clk [5160]));
Q_ASSIGN U27615 ( .B(clk), .A(\g.we_clk [5159]));
Q_ASSIGN U27616 ( .B(clk), .A(\g.we_clk [5158]));
Q_ASSIGN U27617 ( .B(clk), .A(\g.we_clk [5157]));
Q_ASSIGN U27618 ( .B(clk), .A(\g.we_clk [5156]));
Q_ASSIGN U27619 ( .B(clk), .A(\g.we_clk [5155]));
Q_ASSIGN U27620 ( .B(clk), .A(\g.we_clk [5154]));
Q_ASSIGN U27621 ( .B(clk), .A(\g.we_clk [5153]));
Q_ASSIGN U27622 ( .B(clk), .A(\g.we_clk [5152]));
Q_ASSIGN U27623 ( .B(clk), .A(\g.we_clk [5151]));
Q_ASSIGN U27624 ( .B(clk), .A(\g.we_clk [5150]));
Q_ASSIGN U27625 ( .B(clk), .A(\g.we_clk [5149]));
Q_ASSIGN U27626 ( .B(clk), .A(\g.we_clk [5148]));
Q_ASSIGN U27627 ( .B(clk), .A(\g.we_clk [5147]));
Q_ASSIGN U27628 ( .B(clk), .A(\g.we_clk [5146]));
Q_ASSIGN U27629 ( .B(clk), .A(\g.we_clk [5145]));
Q_ASSIGN U27630 ( .B(clk), .A(\g.we_clk [5144]));
Q_ASSIGN U27631 ( .B(clk), .A(\g.we_clk [5143]));
Q_ASSIGN U27632 ( .B(clk), .A(\g.we_clk [5142]));
Q_ASSIGN U27633 ( .B(clk), .A(\g.we_clk [5141]));
Q_ASSIGN U27634 ( .B(clk), .A(\g.we_clk [5140]));
Q_ASSIGN U27635 ( .B(clk), .A(\g.we_clk [5139]));
Q_ASSIGN U27636 ( .B(clk), .A(\g.we_clk [5138]));
Q_ASSIGN U27637 ( .B(clk), .A(\g.we_clk [5137]));
Q_ASSIGN U27638 ( .B(clk), .A(\g.we_clk [5136]));
Q_ASSIGN U27639 ( .B(clk), .A(\g.we_clk [5135]));
Q_ASSIGN U27640 ( .B(clk), .A(\g.we_clk [5134]));
Q_ASSIGN U27641 ( .B(clk), .A(\g.we_clk [5133]));
Q_ASSIGN U27642 ( .B(clk), .A(\g.we_clk [5132]));
Q_ASSIGN U27643 ( .B(clk), .A(\g.we_clk [5131]));
Q_ASSIGN U27644 ( .B(clk), .A(\g.we_clk [5130]));
Q_ASSIGN U27645 ( .B(clk), .A(\g.we_clk [5129]));
Q_ASSIGN U27646 ( .B(clk), .A(\g.we_clk [5128]));
Q_ASSIGN U27647 ( .B(clk), .A(\g.we_clk [5127]));
Q_ASSIGN U27648 ( .B(clk), .A(\g.we_clk [5126]));
Q_ASSIGN U27649 ( .B(clk), .A(\g.we_clk [5125]));
Q_ASSIGN U27650 ( .B(clk), .A(\g.we_clk [5124]));
Q_ASSIGN U27651 ( .B(clk), .A(\g.we_clk [5123]));
Q_ASSIGN U27652 ( .B(clk), .A(\g.we_clk [5122]));
Q_ASSIGN U27653 ( .B(clk), .A(\g.we_clk [5121]));
Q_ASSIGN U27654 ( .B(clk), .A(\g.we_clk [5120]));
Q_ASSIGN U27655 ( .B(clk), .A(\g.we_clk [5119]));
Q_ASSIGN U27656 ( .B(clk), .A(\g.we_clk [5118]));
Q_ASSIGN U27657 ( .B(clk), .A(\g.we_clk [5117]));
Q_ASSIGN U27658 ( .B(clk), .A(\g.we_clk [5116]));
Q_ASSIGN U27659 ( .B(clk), .A(\g.we_clk [5115]));
Q_ASSIGN U27660 ( .B(clk), .A(\g.we_clk [5114]));
Q_ASSIGN U27661 ( .B(clk), .A(\g.we_clk [5113]));
Q_ASSIGN U27662 ( .B(clk), .A(\g.we_clk [5112]));
Q_ASSIGN U27663 ( .B(clk), .A(\g.we_clk [5111]));
Q_ASSIGN U27664 ( .B(clk), .A(\g.we_clk [5110]));
Q_ASSIGN U27665 ( .B(clk), .A(\g.we_clk [5109]));
Q_ASSIGN U27666 ( .B(clk), .A(\g.we_clk [5108]));
Q_ASSIGN U27667 ( .B(clk), .A(\g.we_clk [5107]));
Q_ASSIGN U27668 ( .B(clk), .A(\g.we_clk [5106]));
Q_ASSIGN U27669 ( .B(clk), .A(\g.we_clk [5105]));
Q_ASSIGN U27670 ( .B(clk), .A(\g.we_clk [5104]));
Q_ASSIGN U27671 ( .B(clk), .A(\g.we_clk [5103]));
Q_ASSIGN U27672 ( .B(clk), .A(\g.we_clk [5102]));
Q_ASSIGN U27673 ( .B(clk), .A(\g.we_clk [5101]));
Q_ASSIGN U27674 ( .B(clk), .A(\g.we_clk [5100]));
Q_ASSIGN U27675 ( .B(clk), .A(\g.we_clk [5099]));
Q_ASSIGN U27676 ( .B(clk), .A(\g.we_clk [5098]));
Q_ASSIGN U27677 ( .B(clk), .A(\g.we_clk [5097]));
Q_ASSIGN U27678 ( .B(clk), .A(\g.we_clk [5096]));
Q_ASSIGN U27679 ( .B(clk), .A(\g.we_clk [5095]));
Q_ASSIGN U27680 ( .B(clk), .A(\g.we_clk [5094]));
Q_ASSIGN U27681 ( .B(clk), .A(\g.we_clk [5093]));
Q_ASSIGN U27682 ( .B(clk), .A(\g.we_clk [5092]));
Q_ASSIGN U27683 ( .B(clk), .A(\g.we_clk [5091]));
Q_ASSIGN U27684 ( .B(clk), .A(\g.we_clk [5090]));
Q_ASSIGN U27685 ( .B(clk), .A(\g.we_clk [5089]));
Q_ASSIGN U27686 ( .B(clk), .A(\g.we_clk [5088]));
Q_ASSIGN U27687 ( .B(clk), .A(\g.we_clk [5087]));
Q_ASSIGN U27688 ( .B(clk), .A(\g.we_clk [5086]));
Q_ASSIGN U27689 ( .B(clk), .A(\g.we_clk [5085]));
Q_ASSIGN U27690 ( .B(clk), .A(\g.we_clk [5084]));
Q_ASSIGN U27691 ( .B(clk), .A(\g.we_clk [5083]));
Q_ASSIGN U27692 ( .B(clk), .A(\g.we_clk [5082]));
Q_ASSIGN U27693 ( .B(clk), .A(\g.we_clk [5081]));
Q_ASSIGN U27694 ( .B(clk), .A(\g.we_clk [5080]));
Q_ASSIGN U27695 ( .B(clk), .A(\g.we_clk [5079]));
Q_ASSIGN U27696 ( .B(clk), .A(\g.we_clk [5078]));
Q_ASSIGN U27697 ( .B(clk), .A(\g.we_clk [5077]));
Q_ASSIGN U27698 ( .B(clk), .A(\g.we_clk [5076]));
Q_ASSIGN U27699 ( .B(clk), .A(\g.we_clk [5075]));
Q_ASSIGN U27700 ( .B(clk), .A(\g.we_clk [5074]));
Q_ASSIGN U27701 ( .B(clk), .A(\g.we_clk [5073]));
Q_ASSIGN U27702 ( .B(clk), .A(\g.we_clk [5072]));
Q_ASSIGN U27703 ( .B(clk), .A(\g.we_clk [5071]));
Q_ASSIGN U27704 ( .B(clk), .A(\g.we_clk [5070]));
Q_ASSIGN U27705 ( .B(clk), .A(\g.we_clk [5069]));
Q_ASSIGN U27706 ( .B(clk), .A(\g.we_clk [5068]));
Q_ASSIGN U27707 ( .B(clk), .A(\g.we_clk [5067]));
Q_ASSIGN U27708 ( .B(clk), .A(\g.we_clk [5066]));
Q_ASSIGN U27709 ( .B(clk), .A(\g.we_clk [5065]));
Q_ASSIGN U27710 ( .B(clk), .A(\g.we_clk [5064]));
Q_ASSIGN U27711 ( .B(clk), .A(\g.we_clk [5063]));
Q_ASSIGN U27712 ( .B(clk), .A(\g.we_clk [5062]));
Q_ASSIGN U27713 ( .B(clk), .A(\g.we_clk [5061]));
Q_ASSIGN U27714 ( .B(clk), .A(\g.we_clk [5060]));
Q_ASSIGN U27715 ( .B(clk), .A(\g.we_clk [5059]));
Q_ASSIGN U27716 ( .B(clk), .A(\g.we_clk [5058]));
Q_ASSIGN U27717 ( .B(clk), .A(\g.we_clk [5057]));
Q_ASSIGN U27718 ( .B(clk), .A(\g.we_clk [5056]));
Q_ASSIGN U27719 ( .B(clk), .A(\g.we_clk [5055]));
Q_ASSIGN U27720 ( .B(clk), .A(\g.we_clk [5054]));
Q_ASSIGN U27721 ( .B(clk), .A(\g.we_clk [5053]));
Q_ASSIGN U27722 ( .B(clk), .A(\g.we_clk [5052]));
Q_ASSIGN U27723 ( .B(clk), .A(\g.we_clk [5051]));
Q_ASSIGN U27724 ( .B(clk), .A(\g.we_clk [5050]));
Q_ASSIGN U27725 ( .B(clk), .A(\g.we_clk [5049]));
Q_ASSIGN U27726 ( .B(clk), .A(\g.we_clk [5048]));
Q_ASSIGN U27727 ( .B(clk), .A(\g.we_clk [5047]));
Q_ASSIGN U27728 ( .B(clk), .A(\g.we_clk [5046]));
Q_ASSIGN U27729 ( .B(clk), .A(\g.we_clk [5045]));
Q_ASSIGN U27730 ( .B(clk), .A(\g.we_clk [5044]));
Q_ASSIGN U27731 ( .B(clk), .A(\g.we_clk [5043]));
Q_ASSIGN U27732 ( .B(clk), .A(\g.we_clk [5042]));
Q_ASSIGN U27733 ( .B(clk), .A(\g.we_clk [5041]));
Q_ASSIGN U27734 ( .B(clk), .A(\g.we_clk [5040]));
Q_ASSIGN U27735 ( .B(clk), .A(\g.we_clk [5039]));
Q_ASSIGN U27736 ( .B(clk), .A(\g.we_clk [5038]));
Q_ASSIGN U27737 ( .B(clk), .A(\g.we_clk [5037]));
Q_ASSIGN U27738 ( .B(clk), .A(\g.we_clk [5036]));
Q_ASSIGN U27739 ( .B(clk), .A(\g.we_clk [5035]));
Q_ASSIGN U27740 ( .B(clk), .A(\g.we_clk [5034]));
Q_ASSIGN U27741 ( .B(clk), .A(\g.we_clk [5033]));
Q_ASSIGN U27742 ( .B(clk), .A(\g.we_clk [5032]));
Q_ASSIGN U27743 ( .B(clk), .A(\g.we_clk [5031]));
Q_ASSIGN U27744 ( .B(clk), .A(\g.we_clk [5030]));
Q_ASSIGN U27745 ( .B(clk), .A(\g.we_clk [5029]));
Q_ASSIGN U27746 ( .B(clk), .A(\g.we_clk [5028]));
Q_ASSIGN U27747 ( .B(clk), .A(\g.we_clk [5027]));
Q_ASSIGN U27748 ( .B(clk), .A(\g.we_clk [5026]));
Q_ASSIGN U27749 ( .B(clk), .A(\g.we_clk [5025]));
Q_ASSIGN U27750 ( .B(clk), .A(\g.we_clk [5024]));
Q_ASSIGN U27751 ( .B(clk), .A(\g.we_clk [5023]));
Q_ASSIGN U27752 ( .B(clk), .A(\g.we_clk [5022]));
Q_ASSIGN U27753 ( .B(clk), .A(\g.we_clk [5021]));
Q_ASSIGN U27754 ( .B(clk), .A(\g.we_clk [5020]));
Q_ASSIGN U27755 ( .B(clk), .A(\g.we_clk [5019]));
Q_ASSIGN U27756 ( .B(clk), .A(\g.we_clk [5018]));
Q_ASSIGN U27757 ( .B(clk), .A(\g.we_clk [5017]));
Q_ASSIGN U27758 ( .B(clk), .A(\g.we_clk [5016]));
Q_ASSIGN U27759 ( .B(clk), .A(\g.we_clk [5015]));
Q_ASSIGN U27760 ( .B(clk), .A(\g.we_clk [5014]));
Q_ASSIGN U27761 ( .B(clk), .A(\g.we_clk [5013]));
Q_ASSIGN U27762 ( .B(clk), .A(\g.we_clk [5012]));
Q_ASSIGN U27763 ( .B(clk), .A(\g.we_clk [5011]));
Q_ASSIGN U27764 ( .B(clk), .A(\g.we_clk [5010]));
Q_ASSIGN U27765 ( .B(clk), .A(\g.we_clk [5009]));
Q_ASSIGN U27766 ( .B(clk), .A(\g.we_clk [5008]));
Q_ASSIGN U27767 ( .B(clk), .A(\g.we_clk [5007]));
Q_ASSIGN U27768 ( .B(clk), .A(\g.we_clk [5006]));
Q_ASSIGN U27769 ( .B(clk), .A(\g.we_clk [5005]));
Q_ASSIGN U27770 ( .B(clk), .A(\g.we_clk [5004]));
Q_ASSIGN U27771 ( .B(clk), .A(\g.we_clk [5003]));
Q_ASSIGN U27772 ( .B(clk), .A(\g.we_clk [5002]));
Q_ASSIGN U27773 ( .B(clk), .A(\g.we_clk [5001]));
Q_ASSIGN U27774 ( .B(clk), .A(\g.we_clk [5000]));
Q_ASSIGN U27775 ( .B(clk), .A(\g.we_clk [4999]));
Q_ASSIGN U27776 ( .B(clk), .A(\g.we_clk [4998]));
Q_ASSIGN U27777 ( .B(clk), .A(\g.we_clk [4997]));
Q_ASSIGN U27778 ( .B(clk), .A(\g.we_clk [4996]));
Q_ASSIGN U27779 ( .B(clk), .A(\g.we_clk [4995]));
Q_ASSIGN U27780 ( .B(clk), .A(\g.we_clk [4994]));
Q_ASSIGN U27781 ( .B(clk), .A(\g.we_clk [4993]));
Q_ASSIGN U27782 ( .B(clk), .A(\g.we_clk [4992]));
Q_ASSIGN U27783 ( .B(clk), .A(\g.we_clk [4991]));
Q_ASSIGN U27784 ( .B(clk), .A(\g.we_clk [4990]));
Q_ASSIGN U27785 ( .B(clk), .A(\g.we_clk [4989]));
Q_ASSIGN U27786 ( .B(clk), .A(\g.we_clk [4988]));
Q_ASSIGN U27787 ( .B(clk), .A(\g.we_clk [4987]));
Q_ASSIGN U27788 ( .B(clk), .A(\g.we_clk [4986]));
Q_ASSIGN U27789 ( .B(clk), .A(\g.we_clk [4985]));
Q_ASSIGN U27790 ( .B(clk), .A(\g.we_clk [4984]));
Q_ASSIGN U27791 ( .B(clk), .A(\g.we_clk [4983]));
Q_ASSIGN U27792 ( .B(clk), .A(\g.we_clk [4982]));
Q_ASSIGN U27793 ( .B(clk), .A(\g.we_clk [4981]));
Q_ASSIGN U27794 ( .B(clk), .A(\g.we_clk [4980]));
Q_ASSIGN U27795 ( .B(clk), .A(\g.we_clk [4979]));
Q_ASSIGN U27796 ( .B(clk), .A(\g.we_clk [4978]));
Q_ASSIGN U27797 ( .B(clk), .A(\g.we_clk [4977]));
Q_ASSIGN U27798 ( .B(clk), .A(\g.we_clk [4976]));
Q_ASSIGN U27799 ( .B(clk), .A(\g.we_clk [4975]));
Q_ASSIGN U27800 ( .B(clk), .A(\g.we_clk [4974]));
Q_ASSIGN U27801 ( .B(clk), .A(\g.we_clk [4973]));
Q_ASSIGN U27802 ( .B(clk), .A(\g.we_clk [4972]));
Q_ASSIGN U27803 ( .B(clk), .A(\g.we_clk [4971]));
Q_ASSIGN U27804 ( .B(clk), .A(\g.we_clk [4970]));
Q_ASSIGN U27805 ( .B(clk), .A(\g.we_clk [4969]));
Q_ASSIGN U27806 ( .B(clk), .A(\g.we_clk [4968]));
Q_ASSIGN U27807 ( .B(clk), .A(\g.we_clk [4967]));
Q_ASSIGN U27808 ( .B(clk), .A(\g.we_clk [4966]));
Q_ASSIGN U27809 ( .B(clk), .A(\g.we_clk [4965]));
Q_ASSIGN U27810 ( .B(clk), .A(\g.we_clk [4964]));
Q_ASSIGN U27811 ( .B(clk), .A(\g.we_clk [4963]));
Q_ASSIGN U27812 ( .B(clk), .A(\g.we_clk [4962]));
Q_ASSIGN U27813 ( .B(clk), .A(\g.we_clk [4961]));
Q_ASSIGN U27814 ( .B(clk), .A(\g.we_clk [4960]));
Q_ASSIGN U27815 ( .B(clk), .A(\g.we_clk [4959]));
Q_ASSIGN U27816 ( .B(clk), .A(\g.we_clk [4958]));
Q_ASSIGN U27817 ( .B(clk), .A(\g.we_clk [4957]));
Q_ASSIGN U27818 ( .B(clk), .A(\g.we_clk [4956]));
Q_ASSIGN U27819 ( .B(clk), .A(\g.we_clk [4955]));
Q_ASSIGN U27820 ( .B(clk), .A(\g.we_clk [4954]));
Q_ASSIGN U27821 ( .B(clk), .A(\g.we_clk [4953]));
Q_ASSIGN U27822 ( .B(clk), .A(\g.we_clk [4952]));
Q_ASSIGN U27823 ( .B(clk), .A(\g.we_clk [4951]));
Q_ASSIGN U27824 ( .B(clk), .A(\g.we_clk [4950]));
Q_ASSIGN U27825 ( .B(clk), .A(\g.we_clk [4949]));
Q_ASSIGN U27826 ( .B(clk), .A(\g.we_clk [4948]));
Q_ASSIGN U27827 ( .B(clk), .A(\g.we_clk [4947]));
Q_ASSIGN U27828 ( .B(clk), .A(\g.we_clk [4946]));
Q_ASSIGN U27829 ( .B(clk), .A(\g.we_clk [4945]));
Q_ASSIGN U27830 ( .B(clk), .A(\g.we_clk [4944]));
Q_ASSIGN U27831 ( .B(clk), .A(\g.we_clk [4943]));
Q_ASSIGN U27832 ( .B(clk), .A(\g.we_clk [4942]));
Q_ASSIGN U27833 ( .B(clk), .A(\g.we_clk [4941]));
Q_ASSIGN U27834 ( .B(clk), .A(\g.we_clk [4940]));
Q_ASSIGN U27835 ( .B(clk), .A(\g.we_clk [4939]));
Q_ASSIGN U27836 ( .B(clk), .A(\g.we_clk [4938]));
Q_ASSIGN U27837 ( .B(clk), .A(\g.we_clk [4937]));
Q_ASSIGN U27838 ( .B(clk), .A(\g.we_clk [4936]));
Q_ASSIGN U27839 ( .B(clk), .A(\g.we_clk [4935]));
Q_ASSIGN U27840 ( .B(clk), .A(\g.we_clk [4934]));
Q_ASSIGN U27841 ( .B(clk), .A(\g.we_clk [4933]));
Q_ASSIGN U27842 ( .B(clk), .A(\g.we_clk [4932]));
Q_ASSIGN U27843 ( .B(clk), .A(\g.we_clk [4931]));
Q_ASSIGN U27844 ( .B(clk), .A(\g.we_clk [4930]));
Q_ASSIGN U27845 ( .B(clk), .A(\g.we_clk [4929]));
Q_ASSIGN U27846 ( .B(clk), .A(\g.we_clk [4928]));
Q_ASSIGN U27847 ( .B(clk), .A(\g.we_clk [4927]));
Q_ASSIGN U27848 ( .B(clk), .A(\g.we_clk [4926]));
Q_ASSIGN U27849 ( .B(clk), .A(\g.we_clk [4925]));
Q_ASSIGN U27850 ( .B(clk), .A(\g.we_clk [4924]));
Q_ASSIGN U27851 ( .B(clk), .A(\g.we_clk [4923]));
Q_ASSIGN U27852 ( .B(clk), .A(\g.we_clk [4922]));
Q_ASSIGN U27853 ( .B(clk), .A(\g.we_clk [4921]));
Q_ASSIGN U27854 ( .B(clk), .A(\g.we_clk [4920]));
Q_ASSIGN U27855 ( .B(clk), .A(\g.we_clk [4919]));
Q_ASSIGN U27856 ( .B(clk), .A(\g.we_clk [4918]));
Q_ASSIGN U27857 ( .B(clk), .A(\g.we_clk [4917]));
Q_ASSIGN U27858 ( .B(clk), .A(\g.we_clk [4916]));
Q_ASSIGN U27859 ( .B(clk), .A(\g.we_clk [4915]));
Q_ASSIGN U27860 ( .B(clk), .A(\g.we_clk [4914]));
Q_ASSIGN U27861 ( .B(clk), .A(\g.we_clk [4913]));
Q_ASSIGN U27862 ( .B(clk), .A(\g.we_clk [4912]));
Q_ASSIGN U27863 ( .B(clk), .A(\g.we_clk [4911]));
Q_ASSIGN U27864 ( .B(clk), .A(\g.we_clk [4910]));
Q_ASSIGN U27865 ( .B(clk), .A(\g.we_clk [4909]));
Q_ASSIGN U27866 ( .B(clk), .A(\g.we_clk [4908]));
Q_ASSIGN U27867 ( .B(clk), .A(\g.we_clk [4907]));
Q_ASSIGN U27868 ( .B(clk), .A(\g.we_clk [4906]));
Q_ASSIGN U27869 ( .B(clk), .A(\g.we_clk [4905]));
Q_ASSIGN U27870 ( .B(clk), .A(\g.we_clk [4904]));
Q_ASSIGN U27871 ( .B(clk), .A(\g.we_clk [4903]));
Q_ASSIGN U27872 ( .B(clk), .A(\g.we_clk [4902]));
Q_ASSIGN U27873 ( .B(clk), .A(\g.we_clk [4901]));
Q_ASSIGN U27874 ( .B(clk), .A(\g.we_clk [4900]));
Q_ASSIGN U27875 ( .B(clk), .A(\g.we_clk [4899]));
Q_ASSIGN U27876 ( .B(clk), .A(\g.we_clk [4898]));
Q_ASSIGN U27877 ( .B(clk), .A(\g.we_clk [4897]));
Q_ASSIGN U27878 ( .B(clk), .A(\g.we_clk [4896]));
Q_ASSIGN U27879 ( .B(clk), .A(\g.we_clk [4895]));
Q_ASSIGN U27880 ( .B(clk), .A(\g.we_clk [4894]));
Q_ASSIGN U27881 ( .B(clk), .A(\g.we_clk [4893]));
Q_ASSIGN U27882 ( .B(clk), .A(\g.we_clk [4892]));
Q_ASSIGN U27883 ( .B(clk), .A(\g.we_clk [4891]));
Q_ASSIGN U27884 ( .B(clk), .A(\g.we_clk [4890]));
Q_ASSIGN U27885 ( .B(clk), .A(\g.we_clk [4889]));
Q_ASSIGN U27886 ( .B(clk), .A(\g.we_clk [4888]));
Q_ASSIGN U27887 ( .B(clk), .A(\g.we_clk [4887]));
Q_ASSIGN U27888 ( .B(clk), .A(\g.we_clk [4886]));
Q_ASSIGN U27889 ( .B(clk), .A(\g.we_clk [4885]));
Q_ASSIGN U27890 ( .B(clk), .A(\g.we_clk [4884]));
Q_ASSIGN U27891 ( .B(clk), .A(\g.we_clk [4883]));
Q_ASSIGN U27892 ( .B(clk), .A(\g.we_clk [4882]));
Q_ASSIGN U27893 ( .B(clk), .A(\g.we_clk [4881]));
Q_ASSIGN U27894 ( .B(clk), .A(\g.we_clk [4880]));
Q_ASSIGN U27895 ( .B(clk), .A(\g.we_clk [4879]));
Q_ASSIGN U27896 ( .B(clk), .A(\g.we_clk [4878]));
Q_ASSIGN U27897 ( .B(clk), .A(\g.we_clk [4877]));
Q_ASSIGN U27898 ( .B(clk), .A(\g.we_clk [4876]));
Q_ASSIGN U27899 ( .B(clk), .A(\g.we_clk [4875]));
Q_ASSIGN U27900 ( .B(clk), .A(\g.we_clk [4874]));
Q_ASSIGN U27901 ( .B(clk), .A(\g.we_clk [4873]));
Q_ASSIGN U27902 ( .B(clk), .A(\g.we_clk [4872]));
Q_ASSIGN U27903 ( .B(clk), .A(\g.we_clk [4871]));
Q_ASSIGN U27904 ( .B(clk), .A(\g.we_clk [4870]));
Q_ASSIGN U27905 ( .B(clk), .A(\g.we_clk [4869]));
Q_ASSIGN U27906 ( .B(clk), .A(\g.we_clk [4868]));
Q_ASSIGN U27907 ( .B(clk), .A(\g.we_clk [4867]));
Q_ASSIGN U27908 ( .B(clk), .A(\g.we_clk [4866]));
Q_ASSIGN U27909 ( .B(clk), .A(\g.we_clk [4865]));
Q_ASSIGN U27910 ( .B(clk), .A(\g.we_clk [4864]));
Q_ASSIGN U27911 ( .B(clk), .A(\g.we_clk [4863]));
Q_ASSIGN U27912 ( .B(clk), .A(\g.we_clk [4862]));
Q_ASSIGN U27913 ( .B(clk), .A(\g.we_clk [4861]));
Q_ASSIGN U27914 ( .B(clk), .A(\g.we_clk [4860]));
Q_ASSIGN U27915 ( .B(clk), .A(\g.we_clk [4859]));
Q_ASSIGN U27916 ( .B(clk), .A(\g.we_clk [4858]));
Q_ASSIGN U27917 ( .B(clk), .A(\g.we_clk [4857]));
Q_ASSIGN U27918 ( .B(clk), .A(\g.we_clk [4856]));
Q_ASSIGN U27919 ( .B(clk), .A(\g.we_clk [4855]));
Q_ASSIGN U27920 ( .B(clk), .A(\g.we_clk [4854]));
Q_ASSIGN U27921 ( .B(clk), .A(\g.we_clk [4853]));
Q_ASSIGN U27922 ( .B(clk), .A(\g.we_clk [4852]));
Q_ASSIGN U27923 ( .B(clk), .A(\g.we_clk [4851]));
Q_ASSIGN U27924 ( .B(clk), .A(\g.we_clk [4850]));
Q_ASSIGN U27925 ( .B(clk), .A(\g.we_clk [4849]));
Q_ASSIGN U27926 ( .B(clk), .A(\g.we_clk [4848]));
Q_ASSIGN U27927 ( .B(clk), .A(\g.we_clk [4847]));
Q_ASSIGN U27928 ( .B(clk), .A(\g.we_clk [4846]));
Q_ASSIGN U27929 ( .B(clk), .A(\g.we_clk [4845]));
Q_ASSIGN U27930 ( .B(clk), .A(\g.we_clk [4844]));
Q_ASSIGN U27931 ( .B(clk), .A(\g.we_clk [4843]));
Q_ASSIGN U27932 ( .B(clk), .A(\g.we_clk [4842]));
Q_ASSIGN U27933 ( .B(clk), .A(\g.we_clk [4841]));
Q_ASSIGN U27934 ( .B(clk), .A(\g.we_clk [4840]));
Q_ASSIGN U27935 ( .B(clk), .A(\g.we_clk [4839]));
Q_ASSIGN U27936 ( .B(clk), .A(\g.we_clk [4838]));
Q_ASSIGN U27937 ( .B(clk), .A(\g.we_clk [4837]));
Q_ASSIGN U27938 ( .B(clk), .A(\g.we_clk [4836]));
Q_ASSIGN U27939 ( .B(clk), .A(\g.we_clk [4835]));
Q_ASSIGN U27940 ( .B(clk), .A(\g.we_clk [4834]));
Q_ASSIGN U27941 ( .B(clk), .A(\g.we_clk [4833]));
Q_ASSIGN U27942 ( .B(clk), .A(\g.we_clk [4832]));
Q_ASSIGN U27943 ( .B(clk), .A(\g.we_clk [4831]));
Q_ASSIGN U27944 ( .B(clk), .A(\g.we_clk [4830]));
Q_ASSIGN U27945 ( .B(clk), .A(\g.we_clk [4829]));
Q_ASSIGN U27946 ( .B(clk), .A(\g.we_clk [4828]));
Q_ASSIGN U27947 ( .B(clk), .A(\g.we_clk [4827]));
Q_ASSIGN U27948 ( .B(clk), .A(\g.we_clk [4826]));
Q_ASSIGN U27949 ( .B(clk), .A(\g.we_clk [4825]));
Q_ASSIGN U27950 ( .B(clk), .A(\g.we_clk [4824]));
Q_ASSIGN U27951 ( .B(clk), .A(\g.we_clk [4823]));
Q_ASSIGN U27952 ( .B(clk), .A(\g.we_clk [4822]));
Q_ASSIGN U27953 ( .B(clk), .A(\g.we_clk [4821]));
Q_ASSIGN U27954 ( .B(clk), .A(\g.we_clk [4820]));
Q_ASSIGN U27955 ( .B(clk), .A(\g.we_clk [4819]));
Q_ASSIGN U27956 ( .B(clk), .A(\g.we_clk [4818]));
Q_ASSIGN U27957 ( .B(clk), .A(\g.we_clk [4817]));
Q_ASSIGN U27958 ( .B(clk), .A(\g.we_clk [4816]));
Q_ASSIGN U27959 ( .B(clk), .A(\g.we_clk [4815]));
Q_ASSIGN U27960 ( .B(clk), .A(\g.we_clk [4814]));
Q_ASSIGN U27961 ( .B(clk), .A(\g.we_clk [4813]));
Q_ASSIGN U27962 ( .B(clk), .A(\g.we_clk [4812]));
Q_ASSIGN U27963 ( .B(clk), .A(\g.we_clk [4811]));
Q_ASSIGN U27964 ( .B(clk), .A(\g.we_clk [4810]));
Q_ASSIGN U27965 ( .B(clk), .A(\g.we_clk [4809]));
Q_ASSIGN U27966 ( .B(clk), .A(\g.we_clk [4808]));
Q_ASSIGN U27967 ( .B(clk), .A(\g.we_clk [4807]));
Q_ASSIGN U27968 ( .B(clk), .A(\g.we_clk [4806]));
Q_ASSIGN U27969 ( .B(clk), .A(\g.we_clk [4805]));
Q_ASSIGN U27970 ( .B(clk), .A(\g.we_clk [4804]));
Q_ASSIGN U27971 ( .B(clk), .A(\g.we_clk [4803]));
Q_ASSIGN U27972 ( .B(clk), .A(\g.we_clk [4802]));
Q_ASSIGN U27973 ( .B(clk), .A(\g.we_clk [4801]));
Q_ASSIGN U27974 ( .B(clk), .A(\g.we_clk [4800]));
Q_ASSIGN U27975 ( .B(clk), .A(\g.we_clk [4799]));
Q_ASSIGN U27976 ( .B(clk), .A(\g.we_clk [4798]));
Q_ASSIGN U27977 ( .B(clk), .A(\g.we_clk [4797]));
Q_ASSIGN U27978 ( .B(clk), .A(\g.we_clk [4796]));
Q_ASSIGN U27979 ( .B(clk), .A(\g.we_clk [4795]));
Q_ASSIGN U27980 ( .B(clk), .A(\g.we_clk [4794]));
Q_ASSIGN U27981 ( .B(clk), .A(\g.we_clk [4793]));
Q_ASSIGN U27982 ( .B(clk), .A(\g.we_clk [4792]));
Q_ASSIGN U27983 ( .B(clk), .A(\g.we_clk [4791]));
Q_ASSIGN U27984 ( .B(clk), .A(\g.we_clk [4790]));
Q_ASSIGN U27985 ( .B(clk), .A(\g.we_clk [4789]));
Q_ASSIGN U27986 ( .B(clk), .A(\g.we_clk [4788]));
Q_ASSIGN U27987 ( .B(clk), .A(\g.we_clk [4787]));
Q_ASSIGN U27988 ( .B(clk), .A(\g.we_clk [4786]));
Q_ASSIGN U27989 ( .B(clk), .A(\g.we_clk [4785]));
Q_ASSIGN U27990 ( .B(clk), .A(\g.we_clk [4784]));
Q_ASSIGN U27991 ( .B(clk), .A(\g.we_clk [4783]));
Q_ASSIGN U27992 ( .B(clk), .A(\g.we_clk [4782]));
Q_ASSIGN U27993 ( .B(clk), .A(\g.we_clk [4781]));
Q_ASSIGN U27994 ( .B(clk), .A(\g.we_clk [4780]));
Q_ASSIGN U27995 ( .B(clk), .A(\g.we_clk [4779]));
Q_ASSIGN U27996 ( .B(clk), .A(\g.we_clk [4778]));
Q_ASSIGN U27997 ( .B(clk), .A(\g.we_clk [4777]));
Q_ASSIGN U27998 ( .B(clk), .A(\g.we_clk [4776]));
Q_ASSIGN U27999 ( .B(clk), .A(\g.we_clk [4775]));
Q_ASSIGN U28000 ( .B(clk), .A(\g.we_clk [4774]));
Q_ASSIGN U28001 ( .B(clk), .A(\g.we_clk [4773]));
Q_ASSIGN U28002 ( .B(clk), .A(\g.we_clk [4772]));
Q_ASSIGN U28003 ( .B(clk), .A(\g.we_clk [4771]));
Q_ASSIGN U28004 ( .B(clk), .A(\g.we_clk [4770]));
Q_ASSIGN U28005 ( .B(clk), .A(\g.we_clk [4769]));
Q_ASSIGN U28006 ( .B(clk), .A(\g.we_clk [4768]));
Q_ASSIGN U28007 ( .B(clk), .A(\g.we_clk [4767]));
Q_ASSIGN U28008 ( .B(clk), .A(\g.we_clk [4766]));
Q_ASSIGN U28009 ( .B(clk), .A(\g.we_clk [4765]));
Q_ASSIGN U28010 ( .B(clk), .A(\g.we_clk [4764]));
Q_ASSIGN U28011 ( .B(clk), .A(\g.we_clk [4763]));
Q_ASSIGN U28012 ( .B(clk), .A(\g.we_clk [4762]));
Q_ASSIGN U28013 ( .B(clk), .A(\g.we_clk [4761]));
Q_ASSIGN U28014 ( .B(clk), .A(\g.we_clk [4760]));
Q_ASSIGN U28015 ( .B(clk), .A(\g.we_clk [4759]));
Q_ASSIGN U28016 ( .B(clk), .A(\g.we_clk [4758]));
Q_ASSIGN U28017 ( .B(clk), .A(\g.we_clk [4757]));
Q_ASSIGN U28018 ( .B(clk), .A(\g.we_clk [4756]));
Q_ASSIGN U28019 ( .B(clk), .A(\g.we_clk [4755]));
Q_ASSIGN U28020 ( .B(clk), .A(\g.we_clk [4754]));
Q_ASSIGN U28021 ( .B(clk), .A(\g.we_clk [4753]));
Q_ASSIGN U28022 ( .B(clk), .A(\g.we_clk [4752]));
Q_ASSIGN U28023 ( .B(clk), .A(\g.we_clk [4751]));
Q_ASSIGN U28024 ( .B(clk), .A(\g.we_clk [4750]));
Q_ASSIGN U28025 ( .B(clk), .A(\g.we_clk [4749]));
Q_ASSIGN U28026 ( .B(clk), .A(\g.we_clk [4748]));
Q_ASSIGN U28027 ( .B(clk), .A(\g.we_clk [4747]));
Q_ASSIGN U28028 ( .B(clk), .A(\g.we_clk [4746]));
Q_ASSIGN U28029 ( .B(clk), .A(\g.we_clk [4745]));
Q_ASSIGN U28030 ( .B(clk), .A(\g.we_clk [4744]));
Q_ASSIGN U28031 ( .B(clk), .A(\g.we_clk [4743]));
Q_ASSIGN U28032 ( .B(clk), .A(\g.we_clk [4742]));
Q_ASSIGN U28033 ( .B(clk), .A(\g.we_clk [4741]));
Q_ASSIGN U28034 ( .B(clk), .A(\g.we_clk [4740]));
Q_ASSIGN U28035 ( .B(clk), .A(\g.we_clk [4739]));
Q_ASSIGN U28036 ( .B(clk), .A(\g.we_clk [4738]));
Q_ASSIGN U28037 ( .B(clk), .A(\g.we_clk [4737]));
Q_ASSIGN U28038 ( .B(clk), .A(\g.we_clk [4736]));
Q_ASSIGN U28039 ( .B(clk), .A(\g.we_clk [4735]));
Q_ASSIGN U28040 ( .B(clk), .A(\g.we_clk [4734]));
Q_ASSIGN U28041 ( .B(clk), .A(\g.we_clk [4733]));
Q_ASSIGN U28042 ( .B(clk), .A(\g.we_clk [4732]));
Q_ASSIGN U28043 ( .B(clk), .A(\g.we_clk [4731]));
Q_ASSIGN U28044 ( .B(clk), .A(\g.we_clk [4730]));
Q_ASSIGN U28045 ( .B(clk), .A(\g.we_clk [4729]));
Q_ASSIGN U28046 ( .B(clk), .A(\g.we_clk [4728]));
Q_ASSIGN U28047 ( .B(clk), .A(\g.we_clk [4727]));
Q_ASSIGN U28048 ( .B(clk), .A(\g.we_clk [4726]));
Q_ASSIGN U28049 ( .B(clk), .A(\g.we_clk [4725]));
Q_ASSIGN U28050 ( .B(clk), .A(\g.we_clk [4724]));
Q_ASSIGN U28051 ( .B(clk), .A(\g.we_clk [4723]));
Q_ASSIGN U28052 ( .B(clk), .A(\g.we_clk [4722]));
Q_ASSIGN U28053 ( .B(clk), .A(\g.we_clk [4721]));
Q_ASSIGN U28054 ( .B(clk), .A(\g.we_clk [4720]));
Q_ASSIGN U28055 ( .B(clk), .A(\g.we_clk [4719]));
Q_ASSIGN U28056 ( .B(clk), .A(\g.we_clk [4718]));
Q_ASSIGN U28057 ( .B(clk), .A(\g.we_clk [4717]));
Q_ASSIGN U28058 ( .B(clk), .A(\g.we_clk [4716]));
Q_ASSIGN U28059 ( .B(clk), .A(\g.we_clk [4715]));
Q_ASSIGN U28060 ( .B(clk), .A(\g.we_clk [4714]));
Q_ASSIGN U28061 ( .B(clk), .A(\g.we_clk [4713]));
Q_ASSIGN U28062 ( .B(clk), .A(\g.we_clk [4712]));
Q_ASSIGN U28063 ( .B(clk), .A(\g.we_clk [4711]));
Q_ASSIGN U28064 ( .B(clk), .A(\g.we_clk [4710]));
Q_ASSIGN U28065 ( .B(clk), .A(\g.we_clk [4709]));
Q_ASSIGN U28066 ( .B(clk), .A(\g.we_clk [4708]));
Q_ASSIGN U28067 ( .B(clk), .A(\g.we_clk [4707]));
Q_ASSIGN U28068 ( .B(clk), .A(\g.we_clk [4706]));
Q_ASSIGN U28069 ( .B(clk), .A(\g.we_clk [4705]));
Q_ASSIGN U28070 ( .B(clk), .A(\g.we_clk [4704]));
Q_ASSIGN U28071 ( .B(clk), .A(\g.we_clk [4703]));
Q_ASSIGN U28072 ( .B(clk), .A(\g.we_clk [4702]));
Q_ASSIGN U28073 ( .B(clk), .A(\g.we_clk [4701]));
Q_ASSIGN U28074 ( .B(clk), .A(\g.we_clk [4700]));
Q_ASSIGN U28075 ( .B(clk), .A(\g.we_clk [4699]));
Q_ASSIGN U28076 ( .B(clk), .A(\g.we_clk [4698]));
Q_ASSIGN U28077 ( .B(clk), .A(\g.we_clk [4697]));
Q_ASSIGN U28078 ( .B(clk), .A(\g.we_clk [4696]));
Q_ASSIGN U28079 ( .B(clk), .A(\g.we_clk [4695]));
Q_ASSIGN U28080 ( .B(clk), .A(\g.we_clk [4694]));
Q_ASSIGN U28081 ( .B(clk), .A(\g.we_clk [4693]));
Q_ASSIGN U28082 ( .B(clk), .A(\g.we_clk [4692]));
Q_ASSIGN U28083 ( .B(clk), .A(\g.we_clk [4691]));
Q_ASSIGN U28084 ( .B(clk), .A(\g.we_clk [4690]));
Q_ASSIGN U28085 ( .B(clk), .A(\g.we_clk [4689]));
Q_ASSIGN U28086 ( .B(clk), .A(\g.we_clk [4688]));
Q_ASSIGN U28087 ( .B(clk), .A(\g.we_clk [4687]));
Q_ASSIGN U28088 ( .B(clk), .A(\g.we_clk [4686]));
Q_ASSIGN U28089 ( .B(clk), .A(\g.we_clk [4685]));
Q_ASSIGN U28090 ( .B(clk), .A(\g.we_clk [4684]));
Q_ASSIGN U28091 ( .B(clk), .A(\g.we_clk [4683]));
Q_ASSIGN U28092 ( .B(clk), .A(\g.we_clk [4682]));
Q_ASSIGN U28093 ( .B(clk), .A(\g.we_clk [4681]));
Q_ASSIGN U28094 ( .B(clk), .A(\g.we_clk [4680]));
Q_ASSIGN U28095 ( .B(clk), .A(\g.we_clk [4679]));
Q_ASSIGN U28096 ( .B(clk), .A(\g.we_clk [4678]));
Q_ASSIGN U28097 ( .B(clk), .A(\g.we_clk [4677]));
Q_ASSIGN U28098 ( .B(clk), .A(\g.we_clk [4676]));
Q_ASSIGN U28099 ( .B(clk), .A(\g.we_clk [4675]));
Q_ASSIGN U28100 ( .B(clk), .A(\g.we_clk [4674]));
Q_ASSIGN U28101 ( .B(clk), .A(\g.we_clk [4673]));
Q_ASSIGN U28102 ( .B(clk), .A(\g.we_clk [4672]));
Q_ASSIGN U28103 ( .B(clk), .A(\g.we_clk [4671]));
Q_ASSIGN U28104 ( .B(clk), .A(\g.we_clk [4670]));
Q_ASSIGN U28105 ( .B(clk), .A(\g.we_clk [4669]));
Q_ASSIGN U28106 ( .B(clk), .A(\g.we_clk [4668]));
Q_ASSIGN U28107 ( .B(clk), .A(\g.we_clk [4667]));
Q_ASSIGN U28108 ( .B(clk), .A(\g.we_clk [4666]));
Q_ASSIGN U28109 ( .B(clk), .A(\g.we_clk [4665]));
Q_ASSIGN U28110 ( .B(clk), .A(\g.we_clk [4664]));
Q_ASSIGN U28111 ( .B(clk), .A(\g.we_clk [4663]));
Q_ASSIGN U28112 ( .B(clk), .A(\g.we_clk [4662]));
Q_ASSIGN U28113 ( .B(clk), .A(\g.we_clk [4661]));
Q_ASSIGN U28114 ( .B(clk), .A(\g.we_clk [4660]));
Q_ASSIGN U28115 ( .B(clk), .A(\g.we_clk [4659]));
Q_ASSIGN U28116 ( .B(clk), .A(\g.we_clk [4658]));
Q_ASSIGN U28117 ( .B(clk), .A(\g.we_clk [4657]));
Q_ASSIGN U28118 ( .B(clk), .A(\g.we_clk [4656]));
Q_ASSIGN U28119 ( .B(clk), .A(\g.we_clk [4655]));
Q_ASSIGN U28120 ( .B(clk), .A(\g.we_clk [4654]));
Q_ASSIGN U28121 ( .B(clk), .A(\g.we_clk [4653]));
Q_ASSIGN U28122 ( .B(clk), .A(\g.we_clk [4652]));
Q_ASSIGN U28123 ( .B(clk), .A(\g.we_clk [4651]));
Q_ASSIGN U28124 ( .B(clk), .A(\g.we_clk [4650]));
Q_ASSIGN U28125 ( .B(clk), .A(\g.we_clk [4649]));
Q_ASSIGN U28126 ( .B(clk), .A(\g.we_clk [4648]));
Q_ASSIGN U28127 ( .B(clk), .A(\g.we_clk [4647]));
Q_ASSIGN U28128 ( .B(clk), .A(\g.we_clk [4646]));
Q_ASSIGN U28129 ( .B(clk), .A(\g.we_clk [4645]));
Q_ASSIGN U28130 ( .B(clk), .A(\g.we_clk [4644]));
Q_ASSIGN U28131 ( .B(clk), .A(\g.we_clk [4643]));
Q_ASSIGN U28132 ( .B(clk), .A(\g.we_clk [4642]));
Q_ASSIGN U28133 ( .B(clk), .A(\g.we_clk [4641]));
Q_ASSIGN U28134 ( .B(clk), .A(\g.we_clk [4640]));
Q_ASSIGN U28135 ( .B(clk), .A(\g.we_clk [4639]));
Q_ASSIGN U28136 ( .B(clk), .A(\g.we_clk [4638]));
Q_ASSIGN U28137 ( .B(clk), .A(\g.we_clk [4637]));
Q_ASSIGN U28138 ( .B(clk), .A(\g.we_clk [4636]));
Q_ASSIGN U28139 ( .B(clk), .A(\g.we_clk [4635]));
Q_ASSIGN U28140 ( .B(clk), .A(\g.we_clk [4634]));
Q_ASSIGN U28141 ( .B(clk), .A(\g.we_clk [4633]));
Q_ASSIGN U28142 ( .B(clk), .A(\g.we_clk [4632]));
Q_ASSIGN U28143 ( .B(clk), .A(\g.we_clk [4631]));
Q_ASSIGN U28144 ( .B(clk), .A(\g.we_clk [4630]));
Q_ASSIGN U28145 ( .B(clk), .A(\g.we_clk [4629]));
Q_ASSIGN U28146 ( .B(clk), .A(\g.we_clk [4628]));
Q_ASSIGN U28147 ( .B(clk), .A(\g.we_clk [4627]));
Q_ASSIGN U28148 ( .B(clk), .A(\g.we_clk [4626]));
Q_ASSIGN U28149 ( .B(clk), .A(\g.we_clk [4625]));
Q_ASSIGN U28150 ( .B(clk), .A(\g.we_clk [4624]));
Q_ASSIGN U28151 ( .B(clk), .A(\g.we_clk [4623]));
Q_ASSIGN U28152 ( .B(clk), .A(\g.we_clk [4622]));
Q_ASSIGN U28153 ( .B(clk), .A(\g.we_clk [4621]));
Q_ASSIGN U28154 ( .B(clk), .A(\g.we_clk [4620]));
Q_ASSIGN U28155 ( .B(clk), .A(\g.we_clk [4619]));
Q_ASSIGN U28156 ( .B(clk), .A(\g.we_clk [4618]));
Q_ASSIGN U28157 ( .B(clk), .A(\g.we_clk [4617]));
Q_ASSIGN U28158 ( .B(clk), .A(\g.we_clk [4616]));
Q_ASSIGN U28159 ( .B(clk), .A(\g.we_clk [4615]));
Q_ASSIGN U28160 ( .B(clk), .A(\g.we_clk [4614]));
Q_ASSIGN U28161 ( .B(clk), .A(\g.we_clk [4613]));
Q_ASSIGN U28162 ( .B(clk), .A(\g.we_clk [4612]));
Q_ASSIGN U28163 ( .B(clk), .A(\g.we_clk [4611]));
Q_ASSIGN U28164 ( .B(clk), .A(\g.we_clk [4610]));
Q_ASSIGN U28165 ( .B(clk), .A(\g.we_clk [4609]));
Q_ASSIGN U28166 ( .B(clk), .A(\g.we_clk [4608]));
Q_ASSIGN U28167 ( .B(clk), .A(\g.we_clk [4607]));
Q_ASSIGN U28168 ( .B(clk), .A(\g.we_clk [4606]));
Q_ASSIGN U28169 ( .B(clk), .A(\g.we_clk [4605]));
Q_ASSIGN U28170 ( .B(clk), .A(\g.we_clk [4604]));
Q_ASSIGN U28171 ( .B(clk), .A(\g.we_clk [4603]));
Q_ASSIGN U28172 ( .B(clk), .A(\g.we_clk [4602]));
Q_ASSIGN U28173 ( .B(clk), .A(\g.we_clk [4601]));
Q_ASSIGN U28174 ( .B(clk), .A(\g.we_clk [4600]));
Q_ASSIGN U28175 ( .B(clk), .A(\g.we_clk [4599]));
Q_ASSIGN U28176 ( .B(clk), .A(\g.we_clk [4598]));
Q_ASSIGN U28177 ( .B(clk), .A(\g.we_clk [4597]));
Q_ASSIGN U28178 ( .B(clk), .A(\g.we_clk [4596]));
Q_ASSIGN U28179 ( .B(clk), .A(\g.we_clk [4595]));
Q_ASSIGN U28180 ( .B(clk), .A(\g.we_clk [4594]));
Q_ASSIGN U28181 ( .B(clk), .A(\g.we_clk [4593]));
Q_ASSIGN U28182 ( .B(clk), .A(\g.we_clk [4592]));
Q_ASSIGN U28183 ( .B(clk), .A(\g.we_clk [4591]));
Q_ASSIGN U28184 ( .B(clk), .A(\g.we_clk [4590]));
Q_ASSIGN U28185 ( .B(clk), .A(\g.we_clk [4589]));
Q_ASSIGN U28186 ( .B(clk), .A(\g.we_clk [4588]));
Q_ASSIGN U28187 ( .B(clk), .A(\g.we_clk [4587]));
Q_ASSIGN U28188 ( .B(clk), .A(\g.we_clk [4586]));
Q_ASSIGN U28189 ( .B(clk), .A(\g.we_clk [4585]));
Q_ASSIGN U28190 ( .B(clk), .A(\g.we_clk [4584]));
Q_ASSIGN U28191 ( .B(clk), .A(\g.we_clk [4583]));
Q_ASSIGN U28192 ( .B(clk), .A(\g.we_clk [4582]));
Q_ASSIGN U28193 ( .B(clk), .A(\g.we_clk [4581]));
Q_ASSIGN U28194 ( .B(clk), .A(\g.we_clk [4580]));
Q_ASSIGN U28195 ( .B(clk), .A(\g.we_clk [4579]));
Q_ASSIGN U28196 ( .B(clk), .A(\g.we_clk [4578]));
Q_ASSIGN U28197 ( .B(clk), .A(\g.we_clk [4577]));
Q_ASSIGN U28198 ( .B(clk), .A(\g.we_clk [4576]));
Q_ASSIGN U28199 ( .B(clk), .A(\g.we_clk [4575]));
Q_ASSIGN U28200 ( .B(clk), .A(\g.we_clk [4574]));
Q_ASSIGN U28201 ( .B(clk), .A(\g.we_clk [4573]));
Q_ASSIGN U28202 ( .B(clk), .A(\g.we_clk [4572]));
Q_ASSIGN U28203 ( .B(clk), .A(\g.we_clk [4571]));
Q_ASSIGN U28204 ( .B(clk), .A(\g.we_clk [4570]));
Q_ASSIGN U28205 ( .B(clk), .A(\g.we_clk [4569]));
Q_ASSIGN U28206 ( .B(clk), .A(\g.we_clk [4568]));
Q_ASSIGN U28207 ( .B(clk), .A(\g.we_clk [4567]));
Q_ASSIGN U28208 ( .B(clk), .A(\g.we_clk [4566]));
Q_ASSIGN U28209 ( .B(clk), .A(\g.we_clk [4565]));
Q_ASSIGN U28210 ( .B(clk), .A(\g.we_clk [4564]));
Q_ASSIGN U28211 ( .B(clk), .A(\g.we_clk [4563]));
Q_ASSIGN U28212 ( .B(clk), .A(\g.we_clk [4562]));
Q_ASSIGN U28213 ( .B(clk), .A(\g.we_clk [4561]));
Q_ASSIGN U28214 ( .B(clk), .A(\g.we_clk [4560]));
Q_ASSIGN U28215 ( .B(clk), .A(\g.we_clk [4559]));
Q_ASSIGN U28216 ( .B(clk), .A(\g.we_clk [4558]));
Q_ASSIGN U28217 ( .B(clk), .A(\g.we_clk [4557]));
Q_ASSIGN U28218 ( .B(clk), .A(\g.we_clk [4556]));
Q_ASSIGN U28219 ( .B(clk), .A(\g.we_clk [4555]));
Q_ASSIGN U28220 ( .B(clk), .A(\g.we_clk [4554]));
Q_ASSIGN U28221 ( .B(clk), .A(\g.we_clk [4553]));
Q_ASSIGN U28222 ( .B(clk), .A(\g.we_clk [4552]));
Q_ASSIGN U28223 ( .B(clk), .A(\g.we_clk [4551]));
Q_ASSIGN U28224 ( .B(clk), .A(\g.we_clk [4550]));
Q_ASSIGN U28225 ( .B(clk), .A(\g.we_clk [4549]));
Q_ASSIGN U28226 ( .B(clk), .A(\g.we_clk [4548]));
Q_ASSIGN U28227 ( .B(clk), .A(\g.we_clk [4547]));
Q_ASSIGN U28228 ( .B(clk), .A(\g.we_clk [4546]));
Q_ASSIGN U28229 ( .B(clk), .A(\g.we_clk [4545]));
Q_ASSIGN U28230 ( .B(clk), .A(\g.we_clk [4544]));
Q_ASSIGN U28231 ( .B(clk), .A(\g.we_clk [4543]));
Q_ASSIGN U28232 ( .B(clk), .A(\g.we_clk [4542]));
Q_ASSIGN U28233 ( .B(clk), .A(\g.we_clk [4541]));
Q_ASSIGN U28234 ( .B(clk), .A(\g.we_clk [4540]));
Q_ASSIGN U28235 ( .B(clk), .A(\g.we_clk [4539]));
Q_ASSIGN U28236 ( .B(clk), .A(\g.we_clk [4538]));
Q_ASSIGN U28237 ( .B(clk), .A(\g.we_clk [4537]));
Q_ASSIGN U28238 ( .B(clk), .A(\g.we_clk [4536]));
Q_ASSIGN U28239 ( .B(clk), .A(\g.we_clk [4535]));
Q_ASSIGN U28240 ( .B(clk), .A(\g.we_clk [4534]));
Q_ASSIGN U28241 ( .B(clk), .A(\g.we_clk [4533]));
Q_ASSIGN U28242 ( .B(clk), .A(\g.we_clk [4532]));
Q_ASSIGN U28243 ( .B(clk), .A(\g.we_clk [4531]));
Q_ASSIGN U28244 ( .B(clk), .A(\g.we_clk [4530]));
Q_ASSIGN U28245 ( .B(clk), .A(\g.we_clk [4529]));
Q_ASSIGN U28246 ( .B(clk), .A(\g.we_clk [4528]));
Q_ASSIGN U28247 ( .B(clk), .A(\g.we_clk [4527]));
Q_ASSIGN U28248 ( .B(clk), .A(\g.we_clk [4526]));
Q_ASSIGN U28249 ( .B(clk), .A(\g.we_clk [4525]));
Q_ASSIGN U28250 ( .B(clk), .A(\g.we_clk [4524]));
Q_ASSIGN U28251 ( .B(clk), .A(\g.we_clk [4523]));
Q_ASSIGN U28252 ( .B(clk), .A(\g.we_clk [4522]));
Q_ASSIGN U28253 ( .B(clk), .A(\g.we_clk [4521]));
Q_ASSIGN U28254 ( .B(clk), .A(\g.we_clk [4520]));
Q_ASSIGN U28255 ( .B(clk), .A(\g.we_clk [4519]));
Q_ASSIGN U28256 ( .B(clk), .A(\g.we_clk [4518]));
Q_ASSIGN U28257 ( .B(clk), .A(\g.we_clk [4517]));
Q_ASSIGN U28258 ( .B(clk), .A(\g.we_clk [4516]));
Q_ASSIGN U28259 ( .B(clk), .A(\g.we_clk [4515]));
Q_ASSIGN U28260 ( .B(clk), .A(\g.we_clk [4514]));
Q_ASSIGN U28261 ( .B(clk), .A(\g.we_clk [4513]));
Q_ASSIGN U28262 ( .B(clk), .A(\g.we_clk [4512]));
Q_ASSIGN U28263 ( .B(clk), .A(\g.we_clk [4511]));
Q_ASSIGN U28264 ( .B(clk), .A(\g.we_clk [4510]));
Q_ASSIGN U28265 ( .B(clk), .A(\g.we_clk [4509]));
Q_ASSIGN U28266 ( .B(clk), .A(\g.we_clk [4508]));
Q_ASSIGN U28267 ( .B(clk), .A(\g.we_clk [4507]));
Q_ASSIGN U28268 ( .B(clk), .A(\g.we_clk [4506]));
Q_ASSIGN U28269 ( .B(clk), .A(\g.we_clk [4505]));
Q_ASSIGN U28270 ( .B(clk), .A(\g.we_clk [4504]));
Q_ASSIGN U28271 ( .B(clk), .A(\g.we_clk [4503]));
Q_ASSIGN U28272 ( .B(clk), .A(\g.we_clk [4502]));
Q_ASSIGN U28273 ( .B(clk), .A(\g.we_clk [4501]));
Q_ASSIGN U28274 ( .B(clk), .A(\g.we_clk [4500]));
Q_ASSIGN U28275 ( .B(clk), .A(\g.we_clk [4499]));
Q_ASSIGN U28276 ( .B(clk), .A(\g.we_clk [4498]));
Q_ASSIGN U28277 ( .B(clk), .A(\g.we_clk [4497]));
Q_ASSIGN U28278 ( .B(clk), .A(\g.we_clk [4496]));
Q_ASSIGN U28279 ( .B(clk), .A(\g.we_clk [4495]));
Q_ASSIGN U28280 ( .B(clk), .A(\g.we_clk [4494]));
Q_ASSIGN U28281 ( .B(clk), .A(\g.we_clk [4493]));
Q_ASSIGN U28282 ( .B(clk), .A(\g.we_clk [4492]));
Q_ASSIGN U28283 ( .B(clk), .A(\g.we_clk [4491]));
Q_ASSIGN U28284 ( .B(clk), .A(\g.we_clk [4490]));
Q_ASSIGN U28285 ( .B(clk), .A(\g.we_clk [4489]));
Q_ASSIGN U28286 ( .B(clk), .A(\g.we_clk [4488]));
Q_ASSIGN U28287 ( .B(clk), .A(\g.we_clk [4487]));
Q_ASSIGN U28288 ( .B(clk), .A(\g.we_clk [4486]));
Q_ASSIGN U28289 ( .B(clk), .A(\g.we_clk [4485]));
Q_ASSIGN U28290 ( .B(clk), .A(\g.we_clk [4484]));
Q_ASSIGN U28291 ( .B(clk), .A(\g.we_clk [4483]));
Q_ASSIGN U28292 ( .B(clk), .A(\g.we_clk [4482]));
Q_ASSIGN U28293 ( .B(clk), .A(\g.we_clk [4481]));
Q_ASSIGN U28294 ( .B(clk), .A(\g.we_clk [4480]));
Q_ASSIGN U28295 ( .B(clk), .A(\g.we_clk [4479]));
Q_ASSIGN U28296 ( .B(clk), .A(\g.we_clk [4478]));
Q_ASSIGN U28297 ( .B(clk), .A(\g.we_clk [4477]));
Q_ASSIGN U28298 ( .B(clk), .A(\g.we_clk [4476]));
Q_ASSIGN U28299 ( .B(clk), .A(\g.we_clk [4475]));
Q_ASSIGN U28300 ( .B(clk), .A(\g.we_clk [4474]));
Q_ASSIGN U28301 ( .B(clk), .A(\g.we_clk [4473]));
Q_ASSIGN U28302 ( .B(clk), .A(\g.we_clk [4472]));
Q_ASSIGN U28303 ( .B(clk), .A(\g.we_clk [4471]));
Q_ASSIGN U28304 ( .B(clk), .A(\g.we_clk [4470]));
Q_ASSIGN U28305 ( .B(clk), .A(\g.we_clk [4469]));
Q_ASSIGN U28306 ( .B(clk), .A(\g.we_clk [4468]));
Q_ASSIGN U28307 ( .B(clk), .A(\g.we_clk [4467]));
Q_ASSIGN U28308 ( .B(clk), .A(\g.we_clk [4466]));
Q_ASSIGN U28309 ( .B(clk), .A(\g.we_clk [4465]));
Q_ASSIGN U28310 ( .B(clk), .A(\g.we_clk [4464]));
Q_ASSIGN U28311 ( .B(clk), .A(\g.we_clk [4463]));
Q_ASSIGN U28312 ( .B(clk), .A(\g.we_clk [4462]));
Q_ASSIGN U28313 ( .B(clk), .A(\g.we_clk [4461]));
Q_ASSIGN U28314 ( .B(clk), .A(\g.we_clk [4460]));
Q_ASSIGN U28315 ( .B(clk), .A(\g.we_clk [4459]));
Q_ASSIGN U28316 ( .B(clk), .A(\g.we_clk [4458]));
Q_ASSIGN U28317 ( .B(clk), .A(\g.we_clk [4457]));
Q_ASSIGN U28318 ( .B(clk), .A(\g.we_clk [4456]));
Q_ASSIGN U28319 ( .B(clk), .A(\g.we_clk [4455]));
Q_ASSIGN U28320 ( .B(clk), .A(\g.we_clk [4454]));
Q_ASSIGN U28321 ( .B(clk), .A(\g.we_clk [4453]));
Q_ASSIGN U28322 ( .B(clk), .A(\g.we_clk [4452]));
Q_ASSIGN U28323 ( .B(clk), .A(\g.we_clk [4451]));
Q_ASSIGN U28324 ( .B(clk), .A(\g.we_clk [4450]));
Q_ASSIGN U28325 ( .B(clk), .A(\g.we_clk [4449]));
Q_ASSIGN U28326 ( .B(clk), .A(\g.we_clk [4448]));
Q_ASSIGN U28327 ( .B(clk), .A(\g.we_clk [4447]));
Q_ASSIGN U28328 ( .B(clk), .A(\g.we_clk [4446]));
Q_ASSIGN U28329 ( .B(clk), .A(\g.we_clk [4445]));
Q_ASSIGN U28330 ( .B(clk), .A(\g.we_clk [4444]));
Q_ASSIGN U28331 ( .B(clk), .A(\g.we_clk [4443]));
Q_ASSIGN U28332 ( .B(clk), .A(\g.we_clk [4442]));
Q_ASSIGN U28333 ( .B(clk), .A(\g.we_clk [4441]));
Q_ASSIGN U28334 ( .B(clk), .A(\g.we_clk [4440]));
Q_ASSIGN U28335 ( .B(clk), .A(\g.we_clk [4439]));
Q_ASSIGN U28336 ( .B(clk), .A(\g.we_clk [4438]));
Q_ASSIGN U28337 ( .B(clk), .A(\g.we_clk [4437]));
Q_ASSIGN U28338 ( .B(clk), .A(\g.we_clk [4436]));
Q_ASSIGN U28339 ( .B(clk), .A(\g.we_clk [4435]));
Q_ASSIGN U28340 ( .B(clk), .A(\g.we_clk [4434]));
Q_ASSIGN U28341 ( .B(clk), .A(\g.we_clk [4433]));
Q_ASSIGN U28342 ( .B(clk), .A(\g.we_clk [4432]));
Q_ASSIGN U28343 ( .B(clk), .A(\g.we_clk [4431]));
Q_ASSIGN U28344 ( .B(clk), .A(\g.we_clk [4430]));
Q_ASSIGN U28345 ( .B(clk), .A(\g.we_clk [4429]));
Q_ASSIGN U28346 ( .B(clk), .A(\g.we_clk [4428]));
Q_ASSIGN U28347 ( .B(clk), .A(\g.we_clk [4427]));
Q_ASSIGN U28348 ( .B(clk), .A(\g.we_clk [4426]));
Q_ASSIGN U28349 ( .B(clk), .A(\g.we_clk [4425]));
Q_ASSIGN U28350 ( .B(clk), .A(\g.we_clk [4424]));
Q_ASSIGN U28351 ( .B(clk), .A(\g.we_clk [4423]));
Q_ASSIGN U28352 ( .B(clk), .A(\g.we_clk [4422]));
Q_ASSIGN U28353 ( .B(clk), .A(\g.we_clk [4421]));
Q_ASSIGN U28354 ( .B(clk), .A(\g.we_clk [4420]));
Q_ASSIGN U28355 ( .B(clk), .A(\g.we_clk [4419]));
Q_ASSIGN U28356 ( .B(clk), .A(\g.we_clk [4418]));
Q_ASSIGN U28357 ( .B(clk), .A(\g.we_clk [4417]));
Q_ASSIGN U28358 ( .B(clk), .A(\g.we_clk [4416]));
Q_ASSIGN U28359 ( .B(clk), .A(\g.we_clk [4415]));
Q_ASSIGN U28360 ( .B(clk), .A(\g.we_clk [4414]));
Q_ASSIGN U28361 ( .B(clk), .A(\g.we_clk [4413]));
Q_ASSIGN U28362 ( .B(clk), .A(\g.we_clk [4412]));
Q_ASSIGN U28363 ( .B(clk), .A(\g.we_clk [4411]));
Q_ASSIGN U28364 ( .B(clk), .A(\g.we_clk [4410]));
Q_ASSIGN U28365 ( .B(clk), .A(\g.we_clk [4409]));
Q_ASSIGN U28366 ( .B(clk), .A(\g.we_clk [4408]));
Q_ASSIGN U28367 ( .B(clk), .A(\g.we_clk [4407]));
Q_ASSIGN U28368 ( .B(clk), .A(\g.we_clk [4406]));
Q_ASSIGN U28369 ( .B(clk), .A(\g.we_clk [4405]));
Q_ASSIGN U28370 ( .B(clk), .A(\g.we_clk [4404]));
Q_ASSIGN U28371 ( .B(clk), .A(\g.we_clk [4403]));
Q_ASSIGN U28372 ( .B(clk), .A(\g.we_clk [4402]));
Q_ASSIGN U28373 ( .B(clk), .A(\g.we_clk [4401]));
Q_ASSIGN U28374 ( .B(clk), .A(\g.we_clk [4400]));
Q_ASSIGN U28375 ( .B(clk), .A(\g.we_clk [4399]));
Q_ASSIGN U28376 ( .B(clk), .A(\g.we_clk [4398]));
Q_ASSIGN U28377 ( .B(clk), .A(\g.we_clk [4397]));
Q_ASSIGN U28378 ( .B(clk), .A(\g.we_clk [4396]));
Q_ASSIGN U28379 ( .B(clk), .A(\g.we_clk [4395]));
Q_ASSIGN U28380 ( .B(clk), .A(\g.we_clk [4394]));
Q_ASSIGN U28381 ( .B(clk), .A(\g.we_clk [4393]));
Q_ASSIGN U28382 ( .B(clk), .A(\g.we_clk [4392]));
Q_ASSIGN U28383 ( .B(clk), .A(\g.we_clk [4391]));
Q_ASSIGN U28384 ( .B(clk), .A(\g.we_clk [4390]));
Q_ASSIGN U28385 ( .B(clk), .A(\g.we_clk [4389]));
Q_ASSIGN U28386 ( .B(clk), .A(\g.we_clk [4388]));
Q_ASSIGN U28387 ( .B(clk), .A(\g.we_clk [4387]));
Q_ASSIGN U28388 ( .B(clk), .A(\g.we_clk [4386]));
Q_ASSIGN U28389 ( .B(clk), .A(\g.we_clk [4385]));
Q_ASSIGN U28390 ( .B(clk), .A(\g.we_clk [4384]));
Q_ASSIGN U28391 ( .B(clk), .A(\g.we_clk [4383]));
Q_ASSIGN U28392 ( .B(clk), .A(\g.we_clk [4382]));
Q_ASSIGN U28393 ( .B(clk), .A(\g.we_clk [4381]));
Q_ASSIGN U28394 ( .B(clk), .A(\g.we_clk [4380]));
Q_ASSIGN U28395 ( .B(clk), .A(\g.we_clk [4379]));
Q_ASSIGN U28396 ( .B(clk), .A(\g.we_clk [4378]));
Q_ASSIGN U28397 ( .B(clk), .A(\g.we_clk [4377]));
Q_ASSIGN U28398 ( .B(clk), .A(\g.we_clk [4376]));
Q_ASSIGN U28399 ( .B(clk), .A(\g.we_clk [4375]));
Q_ASSIGN U28400 ( .B(clk), .A(\g.we_clk [4374]));
Q_ASSIGN U28401 ( .B(clk), .A(\g.we_clk [4373]));
Q_ASSIGN U28402 ( .B(clk), .A(\g.we_clk [4372]));
Q_ASSIGN U28403 ( .B(clk), .A(\g.we_clk [4371]));
Q_ASSIGN U28404 ( .B(clk), .A(\g.we_clk [4370]));
Q_ASSIGN U28405 ( .B(clk), .A(\g.we_clk [4369]));
Q_ASSIGN U28406 ( .B(clk), .A(\g.we_clk [4368]));
Q_ASSIGN U28407 ( .B(clk), .A(\g.we_clk [4367]));
Q_ASSIGN U28408 ( .B(clk), .A(\g.we_clk [4366]));
Q_ASSIGN U28409 ( .B(clk), .A(\g.we_clk [4365]));
Q_ASSIGN U28410 ( .B(clk), .A(\g.we_clk [4364]));
Q_ASSIGN U28411 ( .B(clk), .A(\g.we_clk [4363]));
Q_ASSIGN U28412 ( .B(clk), .A(\g.we_clk [4362]));
Q_ASSIGN U28413 ( .B(clk), .A(\g.we_clk [4361]));
Q_ASSIGN U28414 ( .B(clk), .A(\g.we_clk [4360]));
Q_ASSIGN U28415 ( .B(clk), .A(\g.we_clk [4359]));
Q_ASSIGN U28416 ( .B(clk), .A(\g.we_clk [4358]));
Q_ASSIGN U28417 ( .B(clk), .A(\g.we_clk [4357]));
Q_ASSIGN U28418 ( .B(clk), .A(\g.we_clk [4356]));
Q_ASSIGN U28419 ( .B(clk), .A(\g.we_clk [4355]));
Q_ASSIGN U28420 ( .B(clk), .A(\g.we_clk [4354]));
Q_ASSIGN U28421 ( .B(clk), .A(\g.we_clk [4353]));
Q_ASSIGN U28422 ( .B(clk), .A(\g.we_clk [4352]));
Q_ASSIGN U28423 ( .B(clk), .A(\g.we_clk [4351]));
Q_ASSIGN U28424 ( .B(clk), .A(\g.we_clk [4350]));
Q_ASSIGN U28425 ( .B(clk), .A(\g.we_clk [4349]));
Q_ASSIGN U28426 ( .B(clk), .A(\g.we_clk [4348]));
Q_ASSIGN U28427 ( .B(clk), .A(\g.we_clk [4347]));
Q_ASSIGN U28428 ( .B(clk), .A(\g.we_clk [4346]));
Q_ASSIGN U28429 ( .B(clk), .A(\g.we_clk [4345]));
Q_ASSIGN U28430 ( .B(clk), .A(\g.we_clk [4344]));
Q_ASSIGN U28431 ( .B(clk), .A(\g.we_clk [4343]));
Q_ASSIGN U28432 ( .B(clk), .A(\g.we_clk [4342]));
Q_ASSIGN U28433 ( .B(clk), .A(\g.we_clk [4341]));
Q_ASSIGN U28434 ( .B(clk), .A(\g.we_clk [4340]));
Q_ASSIGN U28435 ( .B(clk), .A(\g.we_clk [4339]));
Q_ASSIGN U28436 ( .B(clk), .A(\g.we_clk [4338]));
Q_ASSIGN U28437 ( .B(clk), .A(\g.we_clk [4337]));
Q_ASSIGN U28438 ( .B(clk), .A(\g.we_clk [4336]));
Q_ASSIGN U28439 ( .B(clk), .A(\g.we_clk [4335]));
Q_ASSIGN U28440 ( .B(clk), .A(\g.we_clk [4334]));
Q_ASSIGN U28441 ( .B(clk), .A(\g.we_clk [4333]));
Q_ASSIGN U28442 ( .B(clk), .A(\g.we_clk [4332]));
Q_ASSIGN U28443 ( .B(clk), .A(\g.we_clk [4331]));
Q_ASSIGN U28444 ( .B(clk), .A(\g.we_clk [4330]));
Q_ASSIGN U28445 ( .B(clk), .A(\g.we_clk [4329]));
Q_ASSIGN U28446 ( .B(clk), .A(\g.we_clk [4328]));
Q_ASSIGN U28447 ( .B(clk), .A(\g.we_clk [4327]));
Q_ASSIGN U28448 ( .B(clk), .A(\g.we_clk [4326]));
Q_ASSIGN U28449 ( .B(clk), .A(\g.we_clk [4325]));
Q_ASSIGN U28450 ( .B(clk), .A(\g.we_clk [4324]));
Q_ASSIGN U28451 ( .B(clk), .A(\g.we_clk [4323]));
Q_ASSIGN U28452 ( .B(clk), .A(\g.we_clk [4322]));
Q_ASSIGN U28453 ( .B(clk), .A(\g.we_clk [4321]));
Q_ASSIGN U28454 ( .B(clk), .A(\g.we_clk [4320]));
Q_ASSIGN U28455 ( .B(clk), .A(\g.we_clk [4319]));
Q_ASSIGN U28456 ( .B(clk), .A(\g.we_clk [4318]));
Q_ASSIGN U28457 ( .B(clk), .A(\g.we_clk [4317]));
Q_ASSIGN U28458 ( .B(clk), .A(\g.we_clk [4316]));
Q_ASSIGN U28459 ( .B(clk), .A(\g.we_clk [4315]));
Q_ASSIGN U28460 ( .B(clk), .A(\g.we_clk [4314]));
Q_ASSIGN U28461 ( .B(clk), .A(\g.we_clk [4313]));
Q_ASSIGN U28462 ( .B(clk), .A(\g.we_clk [4312]));
Q_ASSIGN U28463 ( .B(clk), .A(\g.we_clk [4311]));
Q_ASSIGN U28464 ( .B(clk), .A(\g.we_clk [4310]));
Q_ASSIGN U28465 ( .B(clk), .A(\g.we_clk [4309]));
Q_ASSIGN U28466 ( .B(clk), .A(\g.we_clk [4308]));
Q_ASSIGN U28467 ( .B(clk), .A(\g.we_clk [4307]));
Q_ASSIGN U28468 ( .B(clk), .A(\g.we_clk [4306]));
Q_ASSIGN U28469 ( .B(clk), .A(\g.we_clk [4305]));
Q_ASSIGN U28470 ( .B(clk), .A(\g.we_clk [4304]));
Q_ASSIGN U28471 ( .B(clk), .A(\g.we_clk [4303]));
Q_ASSIGN U28472 ( .B(clk), .A(\g.we_clk [4302]));
Q_ASSIGN U28473 ( .B(clk), .A(\g.we_clk [4301]));
Q_ASSIGN U28474 ( .B(clk), .A(\g.we_clk [4300]));
Q_ASSIGN U28475 ( .B(clk), .A(\g.we_clk [4299]));
Q_ASSIGN U28476 ( .B(clk), .A(\g.we_clk [4298]));
Q_ASSIGN U28477 ( .B(clk), .A(\g.we_clk [4297]));
Q_ASSIGN U28478 ( .B(clk), .A(\g.we_clk [4296]));
Q_ASSIGN U28479 ( .B(clk), .A(\g.we_clk [4295]));
Q_ASSIGN U28480 ( .B(clk), .A(\g.we_clk [4294]));
Q_ASSIGN U28481 ( .B(clk), .A(\g.we_clk [4293]));
Q_ASSIGN U28482 ( .B(clk), .A(\g.we_clk [4292]));
Q_ASSIGN U28483 ( .B(clk), .A(\g.we_clk [4291]));
Q_ASSIGN U28484 ( .B(clk), .A(\g.we_clk [4290]));
Q_ASSIGN U28485 ( .B(clk), .A(\g.we_clk [4289]));
Q_ASSIGN U28486 ( .B(clk), .A(\g.we_clk [4288]));
Q_ASSIGN U28487 ( .B(clk), .A(\g.we_clk [4287]));
Q_ASSIGN U28488 ( .B(clk), .A(\g.we_clk [4286]));
Q_ASSIGN U28489 ( .B(clk), .A(\g.we_clk [4285]));
Q_ASSIGN U28490 ( .B(clk), .A(\g.we_clk [4284]));
Q_ASSIGN U28491 ( .B(clk), .A(\g.we_clk [4283]));
Q_ASSIGN U28492 ( .B(clk), .A(\g.we_clk [4282]));
Q_ASSIGN U28493 ( .B(clk), .A(\g.we_clk [4281]));
Q_ASSIGN U28494 ( .B(clk), .A(\g.we_clk [4280]));
Q_ASSIGN U28495 ( .B(clk), .A(\g.we_clk [4279]));
Q_ASSIGN U28496 ( .B(clk), .A(\g.we_clk [4278]));
Q_ASSIGN U28497 ( .B(clk), .A(\g.we_clk [4277]));
Q_ASSIGN U28498 ( .B(clk), .A(\g.we_clk [4276]));
Q_ASSIGN U28499 ( .B(clk), .A(\g.we_clk [4275]));
Q_ASSIGN U28500 ( .B(clk), .A(\g.we_clk [4274]));
Q_ASSIGN U28501 ( .B(clk), .A(\g.we_clk [4273]));
Q_ASSIGN U28502 ( .B(clk), .A(\g.we_clk [4272]));
Q_ASSIGN U28503 ( .B(clk), .A(\g.we_clk [4271]));
Q_ASSIGN U28504 ( .B(clk), .A(\g.we_clk [4270]));
Q_ASSIGN U28505 ( .B(clk), .A(\g.we_clk [4269]));
Q_ASSIGN U28506 ( .B(clk), .A(\g.we_clk [4268]));
Q_ASSIGN U28507 ( .B(clk), .A(\g.we_clk [4267]));
Q_ASSIGN U28508 ( .B(clk), .A(\g.we_clk [4266]));
Q_ASSIGN U28509 ( .B(clk), .A(\g.we_clk [4265]));
Q_ASSIGN U28510 ( .B(clk), .A(\g.we_clk [4264]));
Q_ASSIGN U28511 ( .B(clk), .A(\g.we_clk [4263]));
Q_ASSIGN U28512 ( .B(clk), .A(\g.we_clk [4262]));
Q_ASSIGN U28513 ( .B(clk), .A(\g.we_clk [4261]));
Q_ASSIGN U28514 ( .B(clk), .A(\g.we_clk [4260]));
Q_ASSIGN U28515 ( .B(clk), .A(\g.we_clk [4259]));
Q_ASSIGN U28516 ( .B(clk), .A(\g.we_clk [4258]));
Q_ASSIGN U28517 ( .B(clk), .A(\g.we_clk [4257]));
Q_ASSIGN U28518 ( .B(clk), .A(\g.we_clk [4256]));
Q_ASSIGN U28519 ( .B(clk), .A(\g.we_clk [4255]));
Q_ASSIGN U28520 ( .B(clk), .A(\g.we_clk [4254]));
Q_ASSIGN U28521 ( .B(clk), .A(\g.we_clk [4253]));
Q_ASSIGN U28522 ( .B(clk), .A(\g.we_clk [4252]));
Q_ASSIGN U28523 ( .B(clk), .A(\g.we_clk [4251]));
Q_ASSIGN U28524 ( .B(clk), .A(\g.we_clk [4250]));
Q_ASSIGN U28525 ( .B(clk), .A(\g.we_clk [4249]));
Q_ASSIGN U28526 ( .B(clk), .A(\g.we_clk [4248]));
Q_ASSIGN U28527 ( .B(clk), .A(\g.we_clk [4247]));
Q_ASSIGN U28528 ( .B(clk), .A(\g.we_clk [4246]));
Q_ASSIGN U28529 ( .B(clk), .A(\g.we_clk [4245]));
Q_ASSIGN U28530 ( .B(clk), .A(\g.we_clk [4244]));
Q_ASSIGN U28531 ( .B(clk), .A(\g.we_clk [4243]));
Q_ASSIGN U28532 ( .B(clk), .A(\g.we_clk [4242]));
Q_ASSIGN U28533 ( .B(clk), .A(\g.we_clk [4241]));
Q_ASSIGN U28534 ( .B(clk), .A(\g.we_clk [4240]));
Q_ASSIGN U28535 ( .B(clk), .A(\g.we_clk [4239]));
Q_ASSIGN U28536 ( .B(clk), .A(\g.we_clk [4238]));
Q_ASSIGN U28537 ( .B(clk), .A(\g.we_clk [4237]));
Q_ASSIGN U28538 ( .B(clk), .A(\g.we_clk [4236]));
Q_ASSIGN U28539 ( .B(clk), .A(\g.we_clk [4235]));
Q_ASSIGN U28540 ( .B(clk), .A(\g.we_clk [4234]));
Q_ASSIGN U28541 ( .B(clk), .A(\g.we_clk [4233]));
Q_ASSIGN U28542 ( .B(clk), .A(\g.we_clk [4232]));
Q_ASSIGN U28543 ( .B(clk), .A(\g.we_clk [4231]));
Q_ASSIGN U28544 ( .B(clk), .A(\g.we_clk [4230]));
Q_ASSIGN U28545 ( .B(clk), .A(\g.we_clk [4229]));
Q_ASSIGN U28546 ( .B(clk), .A(\g.we_clk [4228]));
Q_ASSIGN U28547 ( .B(clk), .A(\g.we_clk [4227]));
Q_ASSIGN U28548 ( .B(clk), .A(\g.we_clk [4226]));
Q_ASSIGN U28549 ( .B(clk), .A(\g.we_clk [4225]));
Q_ASSIGN U28550 ( .B(clk), .A(\g.we_clk [4224]));
Q_ASSIGN U28551 ( .B(clk), .A(\g.we_clk [4223]));
Q_ASSIGN U28552 ( .B(clk), .A(\g.we_clk [4222]));
Q_ASSIGN U28553 ( .B(clk), .A(\g.we_clk [4221]));
Q_ASSIGN U28554 ( .B(clk), .A(\g.we_clk [4220]));
Q_ASSIGN U28555 ( .B(clk), .A(\g.we_clk [4219]));
Q_ASSIGN U28556 ( .B(clk), .A(\g.we_clk [4218]));
Q_ASSIGN U28557 ( .B(clk), .A(\g.we_clk [4217]));
Q_ASSIGN U28558 ( .B(clk), .A(\g.we_clk [4216]));
Q_ASSIGN U28559 ( .B(clk), .A(\g.we_clk [4215]));
Q_ASSIGN U28560 ( .B(clk), .A(\g.we_clk [4214]));
Q_ASSIGN U28561 ( .B(clk), .A(\g.we_clk [4213]));
Q_ASSIGN U28562 ( .B(clk), .A(\g.we_clk [4212]));
Q_ASSIGN U28563 ( .B(clk), .A(\g.we_clk [4211]));
Q_ASSIGN U28564 ( .B(clk), .A(\g.we_clk [4210]));
Q_ASSIGN U28565 ( .B(clk), .A(\g.we_clk [4209]));
Q_ASSIGN U28566 ( .B(clk), .A(\g.we_clk [4208]));
Q_ASSIGN U28567 ( .B(clk), .A(\g.we_clk [4207]));
Q_ASSIGN U28568 ( .B(clk), .A(\g.we_clk [4206]));
Q_ASSIGN U28569 ( .B(clk), .A(\g.we_clk [4205]));
Q_ASSIGN U28570 ( .B(clk), .A(\g.we_clk [4204]));
Q_ASSIGN U28571 ( .B(clk), .A(\g.we_clk [4203]));
Q_ASSIGN U28572 ( .B(clk), .A(\g.we_clk [4202]));
Q_ASSIGN U28573 ( .B(clk), .A(\g.we_clk [4201]));
Q_ASSIGN U28574 ( .B(clk), .A(\g.we_clk [4200]));
Q_ASSIGN U28575 ( .B(clk), .A(\g.we_clk [4199]));
Q_ASSIGN U28576 ( .B(clk), .A(\g.we_clk [4198]));
Q_ASSIGN U28577 ( .B(clk), .A(\g.we_clk [4197]));
Q_ASSIGN U28578 ( .B(clk), .A(\g.we_clk [4196]));
Q_ASSIGN U28579 ( .B(clk), .A(\g.we_clk [4195]));
Q_ASSIGN U28580 ( .B(clk), .A(\g.we_clk [4194]));
Q_ASSIGN U28581 ( .B(clk), .A(\g.we_clk [4193]));
Q_ASSIGN U28582 ( .B(clk), .A(\g.we_clk [4192]));
Q_ASSIGN U28583 ( .B(clk), .A(\g.we_clk [4191]));
Q_ASSIGN U28584 ( .B(clk), .A(\g.we_clk [4190]));
Q_ASSIGN U28585 ( .B(clk), .A(\g.we_clk [4189]));
Q_ASSIGN U28586 ( .B(clk), .A(\g.we_clk [4188]));
Q_ASSIGN U28587 ( .B(clk), .A(\g.we_clk [4187]));
Q_ASSIGN U28588 ( .B(clk), .A(\g.we_clk [4186]));
Q_ASSIGN U28589 ( .B(clk), .A(\g.we_clk [4185]));
Q_ASSIGN U28590 ( .B(clk), .A(\g.we_clk [4184]));
Q_ASSIGN U28591 ( .B(clk), .A(\g.we_clk [4183]));
Q_ASSIGN U28592 ( .B(clk), .A(\g.we_clk [4182]));
Q_ASSIGN U28593 ( .B(clk), .A(\g.we_clk [4181]));
Q_ASSIGN U28594 ( .B(clk), .A(\g.we_clk [4180]));
Q_ASSIGN U28595 ( .B(clk), .A(\g.we_clk [4179]));
Q_ASSIGN U28596 ( .B(clk), .A(\g.we_clk [4178]));
Q_ASSIGN U28597 ( .B(clk), .A(\g.we_clk [4177]));
Q_ASSIGN U28598 ( .B(clk), .A(\g.we_clk [4176]));
Q_ASSIGN U28599 ( .B(clk), .A(\g.we_clk [4175]));
Q_ASSIGN U28600 ( .B(clk), .A(\g.we_clk [4174]));
Q_ASSIGN U28601 ( .B(clk), .A(\g.we_clk [4173]));
Q_ASSIGN U28602 ( .B(clk), .A(\g.we_clk [4172]));
Q_ASSIGN U28603 ( .B(clk), .A(\g.we_clk [4171]));
Q_ASSIGN U28604 ( .B(clk), .A(\g.we_clk [4170]));
Q_ASSIGN U28605 ( .B(clk), .A(\g.we_clk [4169]));
Q_ASSIGN U28606 ( .B(clk), .A(\g.we_clk [4168]));
Q_ASSIGN U28607 ( .B(clk), .A(\g.we_clk [4167]));
Q_ASSIGN U28608 ( .B(clk), .A(\g.we_clk [4166]));
Q_ASSIGN U28609 ( .B(clk), .A(\g.we_clk [4165]));
Q_ASSIGN U28610 ( .B(clk), .A(\g.we_clk [4164]));
Q_ASSIGN U28611 ( .B(clk), .A(\g.we_clk [4163]));
Q_ASSIGN U28612 ( .B(clk), .A(\g.we_clk [4162]));
Q_ASSIGN U28613 ( .B(clk), .A(\g.we_clk [4161]));
Q_ASSIGN U28614 ( .B(clk), .A(\g.we_clk [4160]));
Q_ASSIGN U28615 ( .B(clk), .A(\g.we_clk [4159]));
Q_ASSIGN U28616 ( .B(clk), .A(\g.we_clk [4158]));
Q_ASSIGN U28617 ( .B(clk), .A(\g.we_clk [4157]));
Q_ASSIGN U28618 ( .B(clk), .A(\g.we_clk [4156]));
Q_ASSIGN U28619 ( .B(clk), .A(\g.we_clk [4155]));
Q_ASSIGN U28620 ( .B(clk), .A(\g.we_clk [4154]));
Q_ASSIGN U28621 ( .B(clk), .A(\g.we_clk [4153]));
Q_ASSIGN U28622 ( .B(clk), .A(\g.we_clk [4152]));
Q_ASSIGN U28623 ( .B(clk), .A(\g.we_clk [4151]));
Q_ASSIGN U28624 ( .B(clk), .A(\g.we_clk [4150]));
Q_ASSIGN U28625 ( .B(clk), .A(\g.we_clk [4149]));
Q_ASSIGN U28626 ( .B(clk), .A(\g.we_clk [4148]));
Q_ASSIGN U28627 ( .B(clk), .A(\g.we_clk [4147]));
Q_ASSIGN U28628 ( .B(clk), .A(\g.we_clk [4146]));
Q_ASSIGN U28629 ( .B(clk), .A(\g.we_clk [4145]));
Q_ASSIGN U28630 ( .B(clk), .A(\g.we_clk [4144]));
Q_ASSIGN U28631 ( .B(clk), .A(\g.we_clk [4143]));
Q_ASSIGN U28632 ( .B(clk), .A(\g.we_clk [4142]));
Q_ASSIGN U28633 ( .B(clk), .A(\g.we_clk [4141]));
Q_ASSIGN U28634 ( .B(clk), .A(\g.we_clk [4140]));
Q_ASSIGN U28635 ( .B(clk), .A(\g.we_clk [4139]));
Q_ASSIGN U28636 ( .B(clk), .A(\g.we_clk [4138]));
Q_ASSIGN U28637 ( .B(clk), .A(\g.we_clk [4137]));
Q_ASSIGN U28638 ( .B(clk), .A(\g.we_clk [4136]));
Q_ASSIGN U28639 ( .B(clk), .A(\g.we_clk [4135]));
Q_ASSIGN U28640 ( .B(clk), .A(\g.we_clk [4134]));
Q_ASSIGN U28641 ( .B(clk), .A(\g.we_clk [4133]));
Q_ASSIGN U28642 ( .B(clk), .A(\g.we_clk [4132]));
Q_ASSIGN U28643 ( .B(clk), .A(\g.we_clk [4131]));
Q_ASSIGN U28644 ( .B(clk), .A(\g.we_clk [4130]));
Q_ASSIGN U28645 ( .B(clk), .A(\g.we_clk [4129]));
Q_ASSIGN U28646 ( .B(clk), .A(\g.we_clk [4128]));
Q_ASSIGN U28647 ( .B(clk), .A(\g.we_clk [4127]));
Q_ASSIGN U28648 ( .B(clk), .A(\g.we_clk [4126]));
Q_ASSIGN U28649 ( .B(clk), .A(\g.we_clk [4125]));
Q_ASSIGN U28650 ( .B(clk), .A(\g.we_clk [4124]));
Q_ASSIGN U28651 ( .B(clk), .A(\g.we_clk [4123]));
Q_ASSIGN U28652 ( .B(clk), .A(\g.we_clk [4122]));
Q_ASSIGN U28653 ( .B(clk), .A(\g.we_clk [4121]));
Q_ASSIGN U28654 ( .B(clk), .A(\g.we_clk [4120]));
Q_ASSIGN U28655 ( .B(clk), .A(\g.we_clk [4119]));
Q_ASSIGN U28656 ( .B(clk), .A(\g.we_clk [4118]));
Q_ASSIGN U28657 ( .B(clk), .A(\g.we_clk [4117]));
Q_ASSIGN U28658 ( .B(clk), .A(\g.we_clk [4116]));
Q_ASSIGN U28659 ( .B(clk), .A(\g.we_clk [4115]));
Q_ASSIGN U28660 ( .B(clk), .A(\g.we_clk [4114]));
Q_ASSIGN U28661 ( .B(clk), .A(\g.we_clk [4113]));
Q_ASSIGN U28662 ( .B(clk), .A(\g.we_clk [4112]));
Q_ASSIGN U28663 ( .B(clk), .A(\g.we_clk [4111]));
Q_ASSIGN U28664 ( .B(clk), .A(\g.we_clk [4110]));
Q_ASSIGN U28665 ( .B(clk), .A(\g.we_clk [4109]));
Q_ASSIGN U28666 ( .B(clk), .A(\g.we_clk [4108]));
Q_ASSIGN U28667 ( .B(clk), .A(\g.we_clk [4107]));
Q_ASSIGN U28668 ( .B(clk), .A(\g.we_clk [4106]));
Q_ASSIGN U28669 ( .B(clk), .A(\g.we_clk [4105]));
Q_ASSIGN U28670 ( .B(clk), .A(\g.we_clk [4104]));
Q_ASSIGN U28671 ( .B(clk), .A(\g.we_clk [4103]));
Q_ASSIGN U28672 ( .B(clk), .A(\g.we_clk [4102]));
Q_ASSIGN U28673 ( .B(clk), .A(\g.we_clk [4101]));
Q_ASSIGN U28674 ( .B(clk), .A(\g.we_clk [4100]));
Q_ASSIGN U28675 ( .B(clk), .A(\g.we_clk [4099]));
Q_ASSIGN U28676 ( .B(clk), .A(\g.we_clk [4098]));
Q_ASSIGN U28677 ( .B(clk), .A(\g.we_clk [4097]));
Q_ASSIGN U28678 ( .B(clk), .A(\g.we_clk [4096]));
Q_ASSIGN U28679 ( .B(clk), .A(\g.we_clk [4095]));
Q_ASSIGN U28680 ( .B(clk), .A(\g.we_clk [4094]));
Q_ASSIGN U28681 ( .B(clk), .A(\g.we_clk [4093]));
Q_ASSIGN U28682 ( .B(clk), .A(\g.we_clk [4092]));
Q_ASSIGN U28683 ( .B(clk), .A(\g.we_clk [4091]));
Q_ASSIGN U28684 ( .B(clk), .A(\g.we_clk [4090]));
Q_ASSIGN U28685 ( .B(clk), .A(\g.we_clk [4089]));
Q_ASSIGN U28686 ( .B(clk), .A(\g.we_clk [4088]));
Q_ASSIGN U28687 ( .B(clk), .A(\g.we_clk [4087]));
Q_ASSIGN U28688 ( .B(clk), .A(\g.we_clk [4086]));
Q_ASSIGN U28689 ( .B(clk), .A(\g.we_clk [4085]));
Q_ASSIGN U28690 ( .B(clk), .A(\g.we_clk [4084]));
Q_ASSIGN U28691 ( .B(clk), .A(\g.we_clk [4083]));
Q_ASSIGN U28692 ( .B(clk), .A(\g.we_clk [4082]));
Q_ASSIGN U28693 ( .B(clk), .A(\g.we_clk [4081]));
Q_ASSIGN U28694 ( .B(clk), .A(\g.we_clk [4080]));
Q_ASSIGN U28695 ( .B(clk), .A(\g.we_clk [4079]));
Q_ASSIGN U28696 ( .B(clk), .A(\g.we_clk [4078]));
Q_ASSIGN U28697 ( .B(clk), .A(\g.we_clk [4077]));
Q_ASSIGN U28698 ( .B(clk), .A(\g.we_clk [4076]));
Q_ASSIGN U28699 ( .B(clk), .A(\g.we_clk [4075]));
Q_ASSIGN U28700 ( .B(clk), .A(\g.we_clk [4074]));
Q_ASSIGN U28701 ( .B(clk), .A(\g.we_clk [4073]));
Q_ASSIGN U28702 ( .B(clk), .A(\g.we_clk [4072]));
Q_ASSIGN U28703 ( .B(clk), .A(\g.we_clk [4071]));
Q_ASSIGN U28704 ( .B(clk), .A(\g.we_clk [4070]));
Q_ASSIGN U28705 ( .B(clk), .A(\g.we_clk [4069]));
Q_ASSIGN U28706 ( .B(clk), .A(\g.we_clk [4068]));
Q_ASSIGN U28707 ( .B(clk), .A(\g.we_clk [4067]));
Q_ASSIGN U28708 ( .B(clk), .A(\g.we_clk [4066]));
Q_ASSIGN U28709 ( .B(clk), .A(\g.we_clk [4065]));
Q_ASSIGN U28710 ( .B(clk), .A(\g.we_clk [4064]));
Q_ASSIGN U28711 ( .B(clk), .A(\g.we_clk [4063]));
Q_ASSIGN U28712 ( .B(clk), .A(\g.we_clk [4062]));
Q_ASSIGN U28713 ( .B(clk), .A(\g.we_clk [4061]));
Q_ASSIGN U28714 ( .B(clk), .A(\g.we_clk [4060]));
Q_ASSIGN U28715 ( .B(clk), .A(\g.we_clk [4059]));
Q_ASSIGN U28716 ( .B(clk), .A(\g.we_clk [4058]));
Q_ASSIGN U28717 ( .B(clk), .A(\g.we_clk [4057]));
Q_ASSIGN U28718 ( .B(clk), .A(\g.we_clk [4056]));
Q_ASSIGN U28719 ( .B(clk), .A(\g.we_clk [4055]));
Q_ASSIGN U28720 ( .B(clk), .A(\g.we_clk [4054]));
Q_ASSIGN U28721 ( .B(clk), .A(\g.we_clk [4053]));
Q_ASSIGN U28722 ( .B(clk), .A(\g.we_clk [4052]));
Q_ASSIGN U28723 ( .B(clk), .A(\g.we_clk [4051]));
Q_ASSIGN U28724 ( .B(clk), .A(\g.we_clk [4050]));
Q_ASSIGN U28725 ( .B(clk), .A(\g.we_clk [4049]));
Q_ASSIGN U28726 ( .B(clk), .A(\g.we_clk [4048]));
Q_ASSIGN U28727 ( .B(clk), .A(\g.we_clk [4047]));
Q_ASSIGN U28728 ( .B(clk), .A(\g.we_clk [4046]));
Q_ASSIGN U28729 ( .B(clk), .A(\g.we_clk [4045]));
Q_ASSIGN U28730 ( .B(clk), .A(\g.we_clk [4044]));
Q_ASSIGN U28731 ( .B(clk), .A(\g.we_clk [4043]));
Q_ASSIGN U28732 ( .B(clk), .A(\g.we_clk [4042]));
Q_ASSIGN U28733 ( .B(clk), .A(\g.we_clk [4041]));
Q_ASSIGN U28734 ( .B(clk), .A(\g.we_clk [4040]));
Q_ASSIGN U28735 ( .B(clk), .A(\g.we_clk [4039]));
Q_ASSIGN U28736 ( .B(clk), .A(\g.we_clk [4038]));
Q_ASSIGN U28737 ( .B(clk), .A(\g.we_clk [4037]));
Q_ASSIGN U28738 ( .B(clk), .A(\g.we_clk [4036]));
Q_ASSIGN U28739 ( .B(clk), .A(\g.we_clk [4035]));
Q_ASSIGN U28740 ( .B(clk), .A(\g.we_clk [4034]));
Q_ASSIGN U28741 ( .B(clk), .A(\g.we_clk [4033]));
Q_ASSIGN U28742 ( .B(clk), .A(\g.we_clk [4032]));
Q_ASSIGN U28743 ( .B(clk), .A(\g.we_clk [4031]));
Q_ASSIGN U28744 ( .B(clk), .A(\g.we_clk [4030]));
Q_ASSIGN U28745 ( .B(clk), .A(\g.we_clk [4029]));
Q_ASSIGN U28746 ( .B(clk), .A(\g.we_clk [4028]));
Q_ASSIGN U28747 ( .B(clk), .A(\g.we_clk [4027]));
Q_ASSIGN U28748 ( .B(clk), .A(\g.we_clk [4026]));
Q_ASSIGN U28749 ( .B(clk), .A(\g.we_clk [4025]));
Q_ASSIGN U28750 ( .B(clk), .A(\g.we_clk [4024]));
Q_ASSIGN U28751 ( .B(clk), .A(\g.we_clk [4023]));
Q_ASSIGN U28752 ( .B(clk), .A(\g.we_clk [4022]));
Q_ASSIGN U28753 ( .B(clk), .A(\g.we_clk [4021]));
Q_ASSIGN U28754 ( .B(clk), .A(\g.we_clk [4020]));
Q_ASSIGN U28755 ( .B(clk), .A(\g.we_clk [4019]));
Q_ASSIGN U28756 ( .B(clk), .A(\g.we_clk [4018]));
Q_ASSIGN U28757 ( .B(clk), .A(\g.we_clk [4017]));
Q_ASSIGN U28758 ( .B(clk), .A(\g.we_clk [4016]));
Q_ASSIGN U28759 ( .B(clk), .A(\g.we_clk [4015]));
Q_ASSIGN U28760 ( .B(clk), .A(\g.we_clk [4014]));
Q_ASSIGN U28761 ( .B(clk), .A(\g.we_clk [4013]));
Q_ASSIGN U28762 ( .B(clk), .A(\g.we_clk [4012]));
Q_ASSIGN U28763 ( .B(clk), .A(\g.we_clk [4011]));
Q_ASSIGN U28764 ( .B(clk), .A(\g.we_clk [4010]));
Q_ASSIGN U28765 ( .B(clk), .A(\g.we_clk [4009]));
Q_ASSIGN U28766 ( .B(clk), .A(\g.we_clk [4008]));
Q_ASSIGN U28767 ( .B(clk), .A(\g.we_clk [4007]));
Q_ASSIGN U28768 ( .B(clk), .A(\g.we_clk [4006]));
Q_ASSIGN U28769 ( .B(clk), .A(\g.we_clk [4005]));
Q_ASSIGN U28770 ( .B(clk), .A(\g.we_clk [4004]));
Q_ASSIGN U28771 ( .B(clk), .A(\g.we_clk [4003]));
Q_ASSIGN U28772 ( .B(clk), .A(\g.we_clk [4002]));
Q_ASSIGN U28773 ( .B(clk), .A(\g.we_clk [4001]));
Q_ASSIGN U28774 ( .B(clk), .A(\g.we_clk [4000]));
Q_ASSIGN U28775 ( .B(clk), .A(\g.we_clk [3999]));
Q_ASSIGN U28776 ( .B(clk), .A(\g.we_clk [3998]));
Q_ASSIGN U28777 ( .B(clk), .A(\g.we_clk [3997]));
Q_ASSIGN U28778 ( .B(clk), .A(\g.we_clk [3996]));
Q_ASSIGN U28779 ( .B(clk), .A(\g.we_clk [3995]));
Q_ASSIGN U28780 ( .B(clk), .A(\g.we_clk [3994]));
Q_ASSIGN U28781 ( .B(clk), .A(\g.we_clk [3993]));
Q_ASSIGN U28782 ( .B(clk), .A(\g.we_clk [3992]));
Q_ASSIGN U28783 ( .B(clk), .A(\g.we_clk [3991]));
Q_ASSIGN U28784 ( .B(clk), .A(\g.we_clk [3990]));
Q_ASSIGN U28785 ( .B(clk), .A(\g.we_clk [3989]));
Q_ASSIGN U28786 ( .B(clk), .A(\g.we_clk [3988]));
Q_ASSIGN U28787 ( .B(clk), .A(\g.we_clk [3987]));
Q_ASSIGN U28788 ( .B(clk), .A(\g.we_clk [3986]));
Q_ASSIGN U28789 ( .B(clk), .A(\g.we_clk [3985]));
Q_ASSIGN U28790 ( .B(clk), .A(\g.we_clk [3984]));
Q_ASSIGN U28791 ( .B(clk), .A(\g.we_clk [3983]));
Q_ASSIGN U28792 ( .B(clk), .A(\g.we_clk [3982]));
Q_ASSIGN U28793 ( .B(clk), .A(\g.we_clk [3981]));
Q_ASSIGN U28794 ( .B(clk), .A(\g.we_clk [3980]));
Q_ASSIGN U28795 ( .B(clk), .A(\g.we_clk [3979]));
Q_ASSIGN U28796 ( .B(clk), .A(\g.we_clk [3978]));
Q_ASSIGN U28797 ( .B(clk), .A(\g.we_clk [3977]));
Q_ASSIGN U28798 ( .B(clk), .A(\g.we_clk [3976]));
Q_ASSIGN U28799 ( .B(clk), .A(\g.we_clk [3975]));
Q_ASSIGN U28800 ( .B(clk), .A(\g.we_clk [3974]));
Q_ASSIGN U28801 ( .B(clk), .A(\g.we_clk [3973]));
Q_ASSIGN U28802 ( .B(clk), .A(\g.we_clk [3972]));
Q_ASSIGN U28803 ( .B(clk), .A(\g.we_clk [3971]));
Q_ASSIGN U28804 ( .B(clk), .A(\g.we_clk [3970]));
Q_ASSIGN U28805 ( .B(clk), .A(\g.we_clk [3969]));
Q_ASSIGN U28806 ( .B(clk), .A(\g.we_clk [3968]));
Q_ASSIGN U28807 ( .B(clk), .A(\g.we_clk [3967]));
Q_ASSIGN U28808 ( .B(clk), .A(\g.we_clk [3966]));
Q_ASSIGN U28809 ( .B(clk), .A(\g.we_clk [3965]));
Q_ASSIGN U28810 ( .B(clk), .A(\g.we_clk [3964]));
Q_ASSIGN U28811 ( .B(clk), .A(\g.we_clk [3963]));
Q_ASSIGN U28812 ( .B(clk), .A(\g.we_clk [3962]));
Q_ASSIGN U28813 ( .B(clk), .A(\g.we_clk [3961]));
Q_ASSIGN U28814 ( .B(clk), .A(\g.we_clk [3960]));
Q_ASSIGN U28815 ( .B(clk), .A(\g.we_clk [3959]));
Q_ASSIGN U28816 ( .B(clk), .A(\g.we_clk [3958]));
Q_ASSIGN U28817 ( .B(clk), .A(\g.we_clk [3957]));
Q_ASSIGN U28818 ( .B(clk), .A(\g.we_clk [3956]));
Q_ASSIGN U28819 ( .B(clk), .A(\g.we_clk [3955]));
Q_ASSIGN U28820 ( .B(clk), .A(\g.we_clk [3954]));
Q_ASSIGN U28821 ( .B(clk), .A(\g.we_clk [3953]));
Q_ASSIGN U28822 ( .B(clk), .A(\g.we_clk [3952]));
Q_ASSIGN U28823 ( .B(clk), .A(\g.we_clk [3951]));
Q_ASSIGN U28824 ( .B(clk), .A(\g.we_clk [3950]));
Q_ASSIGN U28825 ( .B(clk), .A(\g.we_clk [3949]));
Q_ASSIGN U28826 ( .B(clk), .A(\g.we_clk [3948]));
Q_ASSIGN U28827 ( .B(clk), .A(\g.we_clk [3947]));
Q_ASSIGN U28828 ( .B(clk), .A(\g.we_clk [3946]));
Q_ASSIGN U28829 ( .B(clk), .A(\g.we_clk [3945]));
Q_ASSIGN U28830 ( .B(clk), .A(\g.we_clk [3944]));
Q_ASSIGN U28831 ( .B(clk), .A(\g.we_clk [3943]));
Q_ASSIGN U28832 ( .B(clk), .A(\g.we_clk [3942]));
Q_ASSIGN U28833 ( .B(clk), .A(\g.we_clk [3941]));
Q_ASSIGN U28834 ( .B(clk), .A(\g.we_clk [3940]));
Q_ASSIGN U28835 ( .B(clk), .A(\g.we_clk [3939]));
Q_ASSIGN U28836 ( .B(clk), .A(\g.we_clk [3938]));
Q_ASSIGN U28837 ( .B(clk), .A(\g.we_clk [3937]));
Q_ASSIGN U28838 ( .B(clk), .A(\g.we_clk [3936]));
Q_ASSIGN U28839 ( .B(clk), .A(\g.we_clk [3935]));
Q_ASSIGN U28840 ( .B(clk), .A(\g.we_clk [3934]));
Q_ASSIGN U28841 ( .B(clk), .A(\g.we_clk [3933]));
Q_ASSIGN U28842 ( .B(clk), .A(\g.we_clk [3932]));
Q_ASSIGN U28843 ( .B(clk), .A(\g.we_clk [3931]));
Q_ASSIGN U28844 ( .B(clk), .A(\g.we_clk [3930]));
Q_ASSIGN U28845 ( .B(clk), .A(\g.we_clk [3929]));
Q_ASSIGN U28846 ( .B(clk), .A(\g.we_clk [3928]));
Q_ASSIGN U28847 ( .B(clk), .A(\g.we_clk [3927]));
Q_ASSIGN U28848 ( .B(clk), .A(\g.we_clk [3926]));
Q_ASSIGN U28849 ( .B(clk), .A(\g.we_clk [3925]));
Q_ASSIGN U28850 ( .B(clk), .A(\g.we_clk [3924]));
Q_ASSIGN U28851 ( .B(clk), .A(\g.we_clk [3923]));
Q_ASSIGN U28852 ( .B(clk), .A(\g.we_clk [3922]));
Q_ASSIGN U28853 ( .B(clk), .A(\g.we_clk [3921]));
Q_ASSIGN U28854 ( .B(clk), .A(\g.we_clk [3920]));
Q_ASSIGN U28855 ( .B(clk), .A(\g.we_clk [3919]));
Q_ASSIGN U28856 ( .B(clk), .A(\g.we_clk [3918]));
Q_ASSIGN U28857 ( .B(clk), .A(\g.we_clk [3917]));
Q_ASSIGN U28858 ( .B(clk), .A(\g.we_clk [3916]));
Q_ASSIGN U28859 ( .B(clk), .A(\g.we_clk [3915]));
Q_ASSIGN U28860 ( .B(clk), .A(\g.we_clk [3914]));
Q_ASSIGN U28861 ( .B(clk), .A(\g.we_clk [3913]));
Q_ASSIGN U28862 ( .B(clk), .A(\g.we_clk [3912]));
Q_ASSIGN U28863 ( .B(clk), .A(\g.we_clk [3911]));
Q_ASSIGN U28864 ( .B(clk), .A(\g.we_clk [3910]));
Q_ASSIGN U28865 ( .B(clk), .A(\g.we_clk [3909]));
Q_ASSIGN U28866 ( .B(clk), .A(\g.we_clk [3908]));
Q_ASSIGN U28867 ( .B(clk), .A(\g.we_clk [3907]));
Q_ASSIGN U28868 ( .B(clk), .A(\g.we_clk [3906]));
Q_ASSIGN U28869 ( .B(clk), .A(\g.we_clk [3905]));
Q_ASSIGN U28870 ( .B(clk), .A(\g.we_clk [3904]));
Q_ASSIGN U28871 ( .B(clk), .A(\g.we_clk [3903]));
Q_ASSIGN U28872 ( .B(clk), .A(\g.we_clk [3902]));
Q_ASSIGN U28873 ( .B(clk), .A(\g.we_clk [3901]));
Q_ASSIGN U28874 ( .B(clk), .A(\g.we_clk [3900]));
Q_ASSIGN U28875 ( .B(clk), .A(\g.we_clk [3899]));
Q_ASSIGN U28876 ( .B(clk), .A(\g.we_clk [3898]));
Q_ASSIGN U28877 ( .B(clk), .A(\g.we_clk [3897]));
Q_ASSIGN U28878 ( .B(clk), .A(\g.we_clk [3896]));
Q_ASSIGN U28879 ( .B(clk), .A(\g.we_clk [3895]));
Q_ASSIGN U28880 ( .B(clk), .A(\g.we_clk [3894]));
Q_ASSIGN U28881 ( .B(clk), .A(\g.we_clk [3893]));
Q_ASSIGN U28882 ( .B(clk), .A(\g.we_clk [3892]));
Q_ASSIGN U28883 ( .B(clk), .A(\g.we_clk [3891]));
Q_ASSIGN U28884 ( .B(clk), .A(\g.we_clk [3890]));
Q_ASSIGN U28885 ( .B(clk), .A(\g.we_clk [3889]));
Q_ASSIGN U28886 ( .B(clk), .A(\g.we_clk [3888]));
Q_ASSIGN U28887 ( .B(clk), .A(\g.we_clk [3887]));
Q_ASSIGN U28888 ( .B(clk), .A(\g.we_clk [3886]));
Q_ASSIGN U28889 ( .B(clk), .A(\g.we_clk [3885]));
Q_ASSIGN U28890 ( .B(clk), .A(\g.we_clk [3884]));
Q_ASSIGN U28891 ( .B(clk), .A(\g.we_clk [3883]));
Q_ASSIGN U28892 ( .B(clk), .A(\g.we_clk [3882]));
Q_ASSIGN U28893 ( .B(clk), .A(\g.we_clk [3881]));
Q_ASSIGN U28894 ( .B(clk), .A(\g.we_clk [3880]));
Q_ASSIGN U28895 ( .B(clk), .A(\g.we_clk [3879]));
Q_ASSIGN U28896 ( .B(clk), .A(\g.we_clk [3878]));
Q_ASSIGN U28897 ( .B(clk), .A(\g.we_clk [3877]));
Q_ASSIGN U28898 ( .B(clk), .A(\g.we_clk [3876]));
Q_ASSIGN U28899 ( .B(clk), .A(\g.we_clk [3875]));
Q_ASSIGN U28900 ( .B(clk), .A(\g.we_clk [3874]));
Q_ASSIGN U28901 ( .B(clk), .A(\g.we_clk [3873]));
Q_ASSIGN U28902 ( .B(clk), .A(\g.we_clk [3872]));
Q_ASSIGN U28903 ( .B(clk), .A(\g.we_clk [3871]));
Q_ASSIGN U28904 ( .B(clk), .A(\g.we_clk [3870]));
Q_ASSIGN U28905 ( .B(clk), .A(\g.we_clk [3869]));
Q_ASSIGN U28906 ( .B(clk), .A(\g.we_clk [3868]));
Q_ASSIGN U28907 ( .B(clk), .A(\g.we_clk [3867]));
Q_ASSIGN U28908 ( .B(clk), .A(\g.we_clk [3866]));
Q_ASSIGN U28909 ( .B(clk), .A(\g.we_clk [3865]));
Q_ASSIGN U28910 ( .B(clk), .A(\g.we_clk [3864]));
Q_ASSIGN U28911 ( .B(clk), .A(\g.we_clk [3863]));
Q_ASSIGN U28912 ( .B(clk), .A(\g.we_clk [3862]));
Q_ASSIGN U28913 ( .B(clk), .A(\g.we_clk [3861]));
Q_ASSIGN U28914 ( .B(clk), .A(\g.we_clk [3860]));
Q_ASSIGN U28915 ( .B(clk), .A(\g.we_clk [3859]));
Q_ASSIGN U28916 ( .B(clk), .A(\g.we_clk [3858]));
Q_ASSIGN U28917 ( .B(clk), .A(\g.we_clk [3857]));
Q_ASSIGN U28918 ( .B(clk), .A(\g.we_clk [3856]));
Q_ASSIGN U28919 ( .B(clk), .A(\g.we_clk [3855]));
Q_ASSIGN U28920 ( .B(clk), .A(\g.we_clk [3854]));
Q_ASSIGN U28921 ( .B(clk), .A(\g.we_clk [3853]));
Q_ASSIGN U28922 ( .B(clk), .A(\g.we_clk [3852]));
Q_ASSIGN U28923 ( .B(clk), .A(\g.we_clk [3851]));
Q_ASSIGN U28924 ( .B(clk), .A(\g.we_clk [3850]));
Q_ASSIGN U28925 ( .B(clk), .A(\g.we_clk [3849]));
Q_ASSIGN U28926 ( .B(clk), .A(\g.we_clk [3848]));
Q_ASSIGN U28927 ( .B(clk), .A(\g.we_clk [3847]));
Q_ASSIGN U28928 ( .B(clk), .A(\g.we_clk [3846]));
Q_ASSIGN U28929 ( .B(clk), .A(\g.we_clk [3845]));
Q_ASSIGN U28930 ( .B(clk), .A(\g.we_clk [3844]));
Q_ASSIGN U28931 ( .B(clk), .A(\g.we_clk [3843]));
Q_ASSIGN U28932 ( .B(clk), .A(\g.we_clk [3842]));
Q_ASSIGN U28933 ( .B(clk), .A(\g.we_clk [3841]));
Q_ASSIGN U28934 ( .B(clk), .A(\g.we_clk [3840]));
Q_ASSIGN U28935 ( .B(clk), .A(\g.we_clk [3839]));
Q_ASSIGN U28936 ( .B(clk), .A(\g.we_clk [3838]));
Q_ASSIGN U28937 ( .B(clk), .A(\g.we_clk [3837]));
Q_ASSIGN U28938 ( .B(clk), .A(\g.we_clk [3836]));
Q_ASSIGN U28939 ( .B(clk), .A(\g.we_clk [3835]));
Q_ASSIGN U28940 ( .B(clk), .A(\g.we_clk [3834]));
Q_ASSIGN U28941 ( .B(clk), .A(\g.we_clk [3833]));
Q_ASSIGN U28942 ( .B(clk), .A(\g.we_clk [3832]));
Q_ASSIGN U28943 ( .B(clk), .A(\g.we_clk [3831]));
Q_ASSIGN U28944 ( .B(clk), .A(\g.we_clk [3830]));
Q_ASSIGN U28945 ( .B(clk), .A(\g.we_clk [3829]));
Q_ASSIGN U28946 ( .B(clk), .A(\g.we_clk [3828]));
Q_ASSIGN U28947 ( .B(clk), .A(\g.we_clk [3827]));
Q_ASSIGN U28948 ( .B(clk), .A(\g.we_clk [3826]));
Q_ASSIGN U28949 ( .B(clk), .A(\g.we_clk [3825]));
Q_ASSIGN U28950 ( .B(clk), .A(\g.we_clk [3824]));
Q_ASSIGN U28951 ( .B(clk), .A(\g.we_clk [3823]));
Q_ASSIGN U28952 ( .B(clk), .A(\g.we_clk [3822]));
Q_ASSIGN U28953 ( .B(clk), .A(\g.we_clk [3821]));
Q_ASSIGN U28954 ( .B(clk), .A(\g.we_clk [3820]));
Q_ASSIGN U28955 ( .B(clk), .A(\g.we_clk [3819]));
Q_ASSIGN U28956 ( .B(clk), .A(\g.we_clk [3818]));
Q_ASSIGN U28957 ( .B(clk), .A(\g.we_clk [3817]));
Q_ASSIGN U28958 ( .B(clk), .A(\g.we_clk [3816]));
Q_ASSIGN U28959 ( .B(clk), .A(\g.we_clk [3815]));
Q_ASSIGN U28960 ( .B(clk), .A(\g.we_clk [3814]));
Q_ASSIGN U28961 ( .B(clk), .A(\g.we_clk [3813]));
Q_ASSIGN U28962 ( .B(clk), .A(\g.we_clk [3812]));
Q_ASSIGN U28963 ( .B(clk), .A(\g.we_clk [3811]));
Q_ASSIGN U28964 ( .B(clk), .A(\g.we_clk [3810]));
Q_ASSIGN U28965 ( .B(clk), .A(\g.we_clk [3809]));
Q_ASSIGN U28966 ( .B(clk), .A(\g.we_clk [3808]));
Q_ASSIGN U28967 ( .B(clk), .A(\g.we_clk [3807]));
Q_ASSIGN U28968 ( .B(clk), .A(\g.we_clk [3806]));
Q_ASSIGN U28969 ( .B(clk), .A(\g.we_clk [3805]));
Q_ASSIGN U28970 ( .B(clk), .A(\g.we_clk [3804]));
Q_ASSIGN U28971 ( .B(clk), .A(\g.we_clk [3803]));
Q_ASSIGN U28972 ( .B(clk), .A(\g.we_clk [3802]));
Q_ASSIGN U28973 ( .B(clk), .A(\g.we_clk [3801]));
Q_ASSIGN U28974 ( .B(clk), .A(\g.we_clk [3800]));
Q_ASSIGN U28975 ( .B(clk), .A(\g.we_clk [3799]));
Q_ASSIGN U28976 ( .B(clk), .A(\g.we_clk [3798]));
Q_ASSIGN U28977 ( .B(clk), .A(\g.we_clk [3797]));
Q_ASSIGN U28978 ( .B(clk), .A(\g.we_clk [3796]));
Q_ASSIGN U28979 ( .B(clk), .A(\g.we_clk [3795]));
Q_ASSIGN U28980 ( .B(clk), .A(\g.we_clk [3794]));
Q_ASSIGN U28981 ( .B(clk), .A(\g.we_clk [3793]));
Q_ASSIGN U28982 ( .B(clk), .A(\g.we_clk [3792]));
Q_ASSIGN U28983 ( .B(clk), .A(\g.we_clk [3791]));
Q_ASSIGN U28984 ( .B(clk), .A(\g.we_clk [3790]));
Q_ASSIGN U28985 ( .B(clk), .A(\g.we_clk [3789]));
Q_ASSIGN U28986 ( .B(clk), .A(\g.we_clk [3788]));
Q_ASSIGN U28987 ( .B(clk), .A(\g.we_clk [3787]));
Q_ASSIGN U28988 ( .B(clk), .A(\g.we_clk [3786]));
Q_ASSIGN U28989 ( .B(clk), .A(\g.we_clk [3785]));
Q_ASSIGN U28990 ( .B(clk), .A(\g.we_clk [3784]));
Q_ASSIGN U28991 ( .B(clk), .A(\g.we_clk [3783]));
Q_ASSIGN U28992 ( .B(clk), .A(\g.we_clk [3782]));
Q_ASSIGN U28993 ( .B(clk), .A(\g.we_clk [3781]));
Q_ASSIGN U28994 ( .B(clk), .A(\g.we_clk [3780]));
Q_ASSIGN U28995 ( .B(clk), .A(\g.we_clk [3779]));
Q_ASSIGN U28996 ( .B(clk), .A(\g.we_clk [3778]));
Q_ASSIGN U28997 ( .B(clk), .A(\g.we_clk [3777]));
Q_ASSIGN U28998 ( .B(clk), .A(\g.we_clk [3776]));
Q_ASSIGN U28999 ( .B(clk), .A(\g.we_clk [3775]));
Q_ASSIGN U29000 ( .B(clk), .A(\g.we_clk [3774]));
Q_ASSIGN U29001 ( .B(clk), .A(\g.we_clk [3773]));
Q_ASSIGN U29002 ( .B(clk), .A(\g.we_clk [3772]));
Q_ASSIGN U29003 ( .B(clk), .A(\g.we_clk [3771]));
Q_ASSIGN U29004 ( .B(clk), .A(\g.we_clk [3770]));
Q_ASSIGN U29005 ( .B(clk), .A(\g.we_clk [3769]));
Q_ASSIGN U29006 ( .B(clk), .A(\g.we_clk [3768]));
Q_ASSIGN U29007 ( .B(clk), .A(\g.we_clk [3767]));
Q_ASSIGN U29008 ( .B(clk), .A(\g.we_clk [3766]));
Q_ASSIGN U29009 ( .B(clk), .A(\g.we_clk [3765]));
Q_ASSIGN U29010 ( .B(clk), .A(\g.we_clk [3764]));
Q_ASSIGN U29011 ( .B(clk), .A(\g.we_clk [3763]));
Q_ASSIGN U29012 ( .B(clk), .A(\g.we_clk [3762]));
Q_ASSIGN U29013 ( .B(clk), .A(\g.we_clk [3761]));
Q_ASSIGN U29014 ( .B(clk), .A(\g.we_clk [3760]));
Q_ASSIGN U29015 ( .B(clk), .A(\g.we_clk [3759]));
Q_ASSIGN U29016 ( .B(clk), .A(\g.we_clk [3758]));
Q_ASSIGN U29017 ( .B(clk), .A(\g.we_clk [3757]));
Q_ASSIGN U29018 ( .B(clk), .A(\g.we_clk [3756]));
Q_ASSIGN U29019 ( .B(clk), .A(\g.we_clk [3755]));
Q_ASSIGN U29020 ( .B(clk), .A(\g.we_clk [3754]));
Q_ASSIGN U29021 ( .B(clk), .A(\g.we_clk [3753]));
Q_ASSIGN U29022 ( .B(clk), .A(\g.we_clk [3752]));
Q_ASSIGN U29023 ( .B(clk), .A(\g.we_clk [3751]));
Q_ASSIGN U29024 ( .B(clk), .A(\g.we_clk [3750]));
Q_ASSIGN U29025 ( .B(clk), .A(\g.we_clk [3749]));
Q_ASSIGN U29026 ( .B(clk), .A(\g.we_clk [3748]));
Q_ASSIGN U29027 ( .B(clk), .A(\g.we_clk [3747]));
Q_ASSIGN U29028 ( .B(clk), .A(\g.we_clk [3746]));
Q_ASSIGN U29029 ( .B(clk), .A(\g.we_clk [3745]));
Q_ASSIGN U29030 ( .B(clk), .A(\g.we_clk [3744]));
Q_ASSIGN U29031 ( .B(clk), .A(\g.we_clk [3743]));
Q_ASSIGN U29032 ( .B(clk), .A(\g.we_clk [3742]));
Q_ASSIGN U29033 ( .B(clk), .A(\g.we_clk [3741]));
Q_ASSIGN U29034 ( .B(clk), .A(\g.we_clk [3740]));
Q_ASSIGN U29035 ( .B(clk), .A(\g.we_clk [3739]));
Q_ASSIGN U29036 ( .B(clk), .A(\g.we_clk [3738]));
Q_ASSIGN U29037 ( .B(clk), .A(\g.we_clk [3737]));
Q_ASSIGN U29038 ( .B(clk), .A(\g.we_clk [3736]));
Q_ASSIGN U29039 ( .B(clk), .A(\g.we_clk [3735]));
Q_ASSIGN U29040 ( .B(clk), .A(\g.we_clk [3734]));
Q_ASSIGN U29041 ( .B(clk), .A(\g.we_clk [3733]));
Q_ASSIGN U29042 ( .B(clk), .A(\g.we_clk [3732]));
Q_ASSIGN U29043 ( .B(clk), .A(\g.we_clk [3731]));
Q_ASSIGN U29044 ( .B(clk), .A(\g.we_clk [3730]));
Q_ASSIGN U29045 ( .B(clk), .A(\g.we_clk [3729]));
Q_ASSIGN U29046 ( .B(clk), .A(\g.we_clk [3728]));
Q_ASSIGN U29047 ( .B(clk), .A(\g.we_clk [3727]));
Q_ASSIGN U29048 ( .B(clk), .A(\g.we_clk [3726]));
Q_ASSIGN U29049 ( .B(clk), .A(\g.we_clk [3725]));
Q_ASSIGN U29050 ( .B(clk), .A(\g.we_clk [3724]));
Q_ASSIGN U29051 ( .B(clk), .A(\g.we_clk [3723]));
Q_ASSIGN U29052 ( .B(clk), .A(\g.we_clk [3722]));
Q_ASSIGN U29053 ( .B(clk), .A(\g.we_clk [3721]));
Q_ASSIGN U29054 ( .B(clk), .A(\g.we_clk [3720]));
Q_ASSIGN U29055 ( .B(clk), .A(\g.we_clk [3719]));
Q_ASSIGN U29056 ( .B(clk), .A(\g.we_clk [3718]));
Q_ASSIGN U29057 ( .B(clk), .A(\g.we_clk [3717]));
Q_ASSIGN U29058 ( .B(clk), .A(\g.we_clk [3716]));
Q_ASSIGN U29059 ( .B(clk), .A(\g.we_clk [3715]));
Q_ASSIGN U29060 ( .B(clk), .A(\g.we_clk [3714]));
Q_ASSIGN U29061 ( .B(clk), .A(\g.we_clk [3713]));
Q_ASSIGN U29062 ( .B(clk), .A(\g.we_clk [3712]));
Q_ASSIGN U29063 ( .B(clk), .A(\g.we_clk [3711]));
Q_ASSIGN U29064 ( .B(clk), .A(\g.we_clk [3710]));
Q_ASSIGN U29065 ( .B(clk), .A(\g.we_clk [3709]));
Q_ASSIGN U29066 ( .B(clk), .A(\g.we_clk [3708]));
Q_ASSIGN U29067 ( .B(clk), .A(\g.we_clk [3707]));
Q_ASSIGN U29068 ( .B(clk), .A(\g.we_clk [3706]));
Q_ASSIGN U29069 ( .B(clk), .A(\g.we_clk [3705]));
Q_ASSIGN U29070 ( .B(clk), .A(\g.we_clk [3704]));
Q_ASSIGN U29071 ( .B(clk), .A(\g.we_clk [3703]));
Q_ASSIGN U29072 ( .B(clk), .A(\g.we_clk [3702]));
Q_ASSIGN U29073 ( .B(clk), .A(\g.we_clk [3701]));
Q_ASSIGN U29074 ( .B(clk), .A(\g.we_clk [3700]));
Q_ASSIGN U29075 ( .B(clk), .A(\g.we_clk [3699]));
Q_ASSIGN U29076 ( .B(clk), .A(\g.we_clk [3698]));
Q_ASSIGN U29077 ( .B(clk), .A(\g.we_clk [3697]));
Q_ASSIGN U29078 ( .B(clk), .A(\g.we_clk [3696]));
Q_ASSIGN U29079 ( .B(clk), .A(\g.we_clk [3695]));
Q_ASSIGN U29080 ( .B(clk), .A(\g.we_clk [3694]));
Q_ASSIGN U29081 ( .B(clk), .A(\g.we_clk [3693]));
Q_ASSIGN U29082 ( .B(clk), .A(\g.we_clk [3692]));
Q_ASSIGN U29083 ( .B(clk), .A(\g.we_clk [3691]));
Q_ASSIGN U29084 ( .B(clk), .A(\g.we_clk [3690]));
Q_ASSIGN U29085 ( .B(clk), .A(\g.we_clk [3689]));
Q_ASSIGN U29086 ( .B(clk), .A(\g.we_clk [3688]));
Q_ASSIGN U29087 ( .B(clk), .A(\g.we_clk [3687]));
Q_ASSIGN U29088 ( .B(clk), .A(\g.we_clk [3686]));
Q_ASSIGN U29089 ( .B(clk), .A(\g.we_clk [3685]));
Q_ASSIGN U29090 ( .B(clk), .A(\g.we_clk [3684]));
Q_ASSIGN U29091 ( .B(clk), .A(\g.we_clk [3683]));
Q_ASSIGN U29092 ( .B(clk), .A(\g.we_clk [3682]));
Q_ASSIGN U29093 ( .B(clk), .A(\g.we_clk [3681]));
Q_ASSIGN U29094 ( .B(clk), .A(\g.we_clk [3680]));
Q_ASSIGN U29095 ( .B(clk), .A(\g.we_clk [3679]));
Q_ASSIGN U29096 ( .B(clk), .A(\g.we_clk [3678]));
Q_ASSIGN U29097 ( .B(clk), .A(\g.we_clk [3677]));
Q_ASSIGN U29098 ( .B(clk), .A(\g.we_clk [3676]));
Q_ASSIGN U29099 ( .B(clk), .A(\g.we_clk [3675]));
Q_ASSIGN U29100 ( .B(clk), .A(\g.we_clk [3674]));
Q_ASSIGN U29101 ( .B(clk), .A(\g.we_clk [3673]));
Q_ASSIGN U29102 ( .B(clk), .A(\g.we_clk [3672]));
Q_ASSIGN U29103 ( .B(clk), .A(\g.we_clk [3671]));
Q_ASSIGN U29104 ( .B(clk), .A(\g.we_clk [3670]));
Q_ASSIGN U29105 ( .B(clk), .A(\g.we_clk [3669]));
Q_ASSIGN U29106 ( .B(clk), .A(\g.we_clk [3668]));
Q_ASSIGN U29107 ( .B(clk), .A(\g.we_clk [3667]));
Q_ASSIGN U29108 ( .B(clk), .A(\g.we_clk [3666]));
Q_ASSIGN U29109 ( .B(clk), .A(\g.we_clk [3665]));
Q_ASSIGN U29110 ( .B(clk), .A(\g.we_clk [3664]));
Q_ASSIGN U29111 ( .B(clk), .A(\g.we_clk [3663]));
Q_ASSIGN U29112 ( .B(clk), .A(\g.we_clk [3662]));
Q_ASSIGN U29113 ( .B(clk), .A(\g.we_clk [3661]));
Q_ASSIGN U29114 ( .B(clk), .A(\g.we_clk [3660]));
Q_ASSIGN U29115 ( .B(clk), .A(\g.we_clk [3659]));
Q_ASSIGN U29116 ( .B(clk), .A(\g.we_clk [3658]));
Q_ASSIGN U29117 ( .B(clk), .A(\g.we_clk [3657]));
Q_ASSIGN U29118 ( .B(clk), .A(\g.we_clk [3656]));
Q_ASSIGN U29119 ( .B(clk), .A(\g.we_clk [3655]));
Q_ASSIGN U29120 ( .B(clk), .A(\g.we_clk [3654]));
Q_ASSIGN U29121 ( .B(clk), .A(\g.we_clk [3653]));
Q_ASSIGN U29122 ( .B(clk), .A(\g.we_clk [3652]));
Q_ASSIGN U29123 ( .B(clk), .A(\g.we_clk [3651]));
Q_ASSIGN U29124 ( .B(clk), .A(\g.we_clk [3650]));
Q_ASSIGN U29125 ( .B(clk), .A(\g.we_clk [3649]));
Q_ASSIGN U29126 ( .B(clk), .A(\g.we_clk [3648]));
Q_ASSIGN U29127 ( .B(clk), .A(\g.we_clk [3647]));
Q_ASSIGN U29128 ( .B(clk), .A(\g.we_clk [3646]));
Q_ASSIGN U29129 ( .B(clk), .A(\g.we_clk [3645]));
Q_ASSIGN U29130 ( .B(clk), .A(\g.we_clk [3644]));
Q_ASSIGN U29131 ( .B(clk), .A(\g.we_clk [3643]));
Q_ASSIGN U29132 ( .B(clk), .A(\g.we_clk [3642]));
Q_ASSIGN U29133 ( .B(clk), .A(\g.we_clk [3641]));
Q_ASSIGN U29134 ( .B(clk), .A(\g.we_clk [3640]));
Q_ASSIGN U29135 ( .B(clk), .A(\g.we_clk [3639]));
Q_ASSIGN U29136 ( .B(clk), .A(\g.we_clk [3638]));
Q_ASSIGN U29137 ( .B(clk), .A(\g.we_clk [3637]));
Q_ASSIGN U29138 ( .B(clk), .A(\g.we_clk [3636]));
Q_ASSIGN U29139 ( .B(clk), .A(\g.we_clk [3635]));
Q_ASSIGN U29140 ( .B(clk), .A(\g.we_clk [3634]));
Q_ASSIGN U29141 ( .B(clk), .A(\g.we_clk [3633]));
Q_ASSIGN U29142 ( .B(clk), .A(\g.we_clk [3632]));
Q_ASSIGN U29143 ( .B(clk), .A(\g.we_clk [3631]));
Q_ASSIGN U29144 ( .B(clk), .A(\g.we_clk [3630]));
Q_ASSIGN U29145 ( .B(clk), .A(\g.we_clk [3629]));
Q_ASSIGN U29146 ( .B(clk), .A(\g.we_clk [3628]));
Q_ASSIGN U29147 ( .B(clk), .A(\g.we_clk [3627]));
Q_ASSIGN U29148 ( .B(clk), .A(\g.we_clk [3626]));
Q_ASSIGN U29149 ( .B(clk), .A(\g.we_clk [3625]));
Q_ASSIGN U29150 ( .B(clk), .A(\g.we_clk [3624]));
Q_ASSIGN U29151 ( .B(clk), .A(\g.we_clk [3623]));
Q_ASSIGN U29152 ( .B(clk), .A(\g.we_clk [3622]));
Q_ASSIGN U29153 ( .B(clk), .A(\g.we_clk [3621]));
Q_ASSIGN U29154 ( .B(clk), .A(\g.we_clk [3620]));
Q_ASSIGN U29155 ( .B(clk), .A(\g.we_clk [3619]));
Q_ASSIGN U29156 ( .B(clk), .A(\g.we_clk [3618]));
Q_ASSIGN U29157 ( .B(clk), .A(\g.we_clk [3617]));
Q_ASSIGN U29158 ( .B(clk), .A(\g.we_clk [3616]));
Q_ASSIGN U29159 ( .B(clk), .A(\g.we_clk [3615]));
Q_ASSIGN U29160 ( .B(clk), .A(\g.we_clk [3614]));
Q_ASSIGN U29161 ( .B(clk), .A(\g.we_clk [3613]));
Q_ASSIGN U29162 ( .B(clk), .A(\g.we_clk [3612]));
Q_ASSIGN U29163 ( .B(clk), .A(\g.we_clk [3611]));
Q_ASSIGN U29164 ( .B(clk), .A(\g.we_clk [3610]));
Q_ASSIGN U29165 ( .B(clk), .A(\g.we_clk [3609]));
Q_ASSIGN U29166 ( .B(clk), .A(\g.we_clk [3608]));
Q_ASSIGN U29167 ( .B(clk), .A(\g.we_clk [3607]));
Q_ASSIGN U29168 ( .B(clk), .A(\g.we_clk [3606]));
Q_ASSIGN U29169 ( .B(clk), .A(\g.we_clk [3605]));
Q_ASSIGN U29170 ( .B(clk), .A(\g.we_clk [3604]));
Q_ASSIGN U29171 ( .B(clk), .A(\g.we_clk [3603]));
Q_ASSIGN U29172 ( .B(clk), .A(\g.we_clk [3602]));
Q_ASSIGN U29173 ( .B(clk), .A(\g.we_clk [3601]));
Q_ASSIGN U29174 ( .B(clk), .A(\g.we_clk [3600]));
Q_ASSIGN U29175 ( .B(clk), .A(\g.we_clk [3599]));
Q_ASSIGN U29176 ( .B(clk), .A(\g.we_clk [3598]));
Q_ASSIGN U29177 ( .B(clk), .A(\g.we_clk [3597]));
Q_ASSIGN U29178 ( .B(clk), .A(\g.we_clk [3596]));
Q_ASSIGN U29179 ( .B(clk), .A(\g.we_clk [3595]));
Q_ASSIGN U29180 ( .B(clk), .A(\g.we_clk [3594]));
Q_ASSIGN U29181 ( .B(clk), .A(\g.we_clk [3593]));
Q_ASSIGN U29182 ( .B(clk), .A(\g.we_clk [3592]));
Q_ASSIGN U29183 ( .B(clk), .A(\g.we_clk [3591]));
Q_ASSIGN U29184 ( .B(clk), .A(\g.we_clk [3590]));
Q_ASSIGN U29185 ( .B(clk), .A(\g.we_clk [3589]));
Q_ASSIGN U29186 ( .B(clk), .A(\g.we_clk [3588]));
Q_ASSIGN U29187 ( .B(clk), .A(\g.we_clk [3587]));
Q_ASSIGN U29188 ( .B(clk), .A(\g.we_clk [3586]));
Q_ASSIGN U29189 ( .B(clk), .A(\g.we_clk [3585]));
Q_ASSIGN U29190 ( .B(clk), .A(\g.we_clk [3584]));
Q_ASSIGN U29191 ( .B(clk), .A(\g.we_clk [3583]));
Q_ASSIGN U29192 ( .B(clk), .A(\g.we_clk [3582]));
Q_ASSIGN U29193 ( .B(clk), .A(\g.we_clk [3581]));
Q_ASSIGN U29194 ( .B(clk), .A(\g.we_clk [3580]));
Q_ASSIGN U29195 ( .B(clk), .A(\g.we_clk [3579]));
Q_ASSIGN U29196 ( .B(clk), .A(\g.we_clk [3578]));
Q_ASSIGN U29197 ( .B(clk), .A(\g.we_clk [3577]));
Q_ASSIGN U29198 ( .B(clk), .A(\g.we_clk [3576]));
Q_ASSIGN U29199 ( .B(clk), .A(\g.we_clk [3575]));
Q_ASSIGN U29200 ( .B(clk), .A(\g.we_clk [3574]));
Q_ASSIGN U29201 ( .B(clk), .A(\g.we_clk [3573]));
Q_ASSIGN U29202 ( .B(clk), .A(\g.we_clk [3572]));
Q_ASSIGN U29203 ( .B(clk), .A(\g.we_clk [3571]));
Q_ASSIGN U29204 ( .B(clk), .A(\g.we_clk [3570]));
Q_ASSIGN U29205 ( .B(clk), .A(\g.we_clk [3569]));
Q_ASSIGN U29206 ( .B(clk), .A(\g.we_clk [3568]));
Q_ASSIGN U29207 ( .B(clk), .A(\g.we_clk [3567]));
Q_ASSIGN U29208 ( .B(clk), .A(\g.we_clk [3566]));
Q_ASSIGN U29209 ( .B(clk), .A(\g.we_clk [3565]));
Q_ASSIGN U29210 ( .B(clk), .A(\g.we_clk [3564]));
Q_ASSIGN U29211 ( .B(clk), .A(\g.we_clk [3563]));
Q_ASSIGN U29212 ( .B(clk), .A(\g.we_clk [3562]));
Q_ASSIGN U29213 ( .B(clk), .A(\g.we_clk [3561]));
Q_ASSIGN U29214 ( .B(clk), .A(\g.we_clk [3560]));
Q_ASSIGN U29215 ( .B(clk), .A(\g.we_clk [3559]));
Q_ASSIGN U29216 ( .B(clk), .A(\g.we_clk [3558]));
Q_ASSIGN U29217 ( .B(clk), .A(\g.we_clk [3557]));
Q_ASSIGN U29218 ( .B(clk), .A(\g.we_clk [3556]));
Q_ASSIGN U29219 ( .B(clk), .A(\g.we_clk [3555]));
Q_ASSIGN U29220 ( .B(clk), .A(\g.we_clk [3554]));
Q_ASSIGN U29221 ( .B(clk), .A(\g.we_clk [3553]));
Q_ASSIGN U29222 ( .B(clk), .A(\g.we_clk [3552]));
Q_ASSIGN U29223 ( .B(clk), .A(\g.we_clk [3551]));
Q_ASSIGN U29224 ( .B(clk), .A(\g.we_clk [3550]));
Q_ASSIGN U29225 ( .B(clk), .A(\g.we_clk [3549]));
Q_ASSIGN U29226 ( .B(clk), .A(\g.we_clk [3548]));
Q_ASSIGN U29227 ( .B(clk), .A(\g.we_clk [3547]));
Q_ASSIGN U29228 ( .B(clk), .A(\g.we_clk [3546]));
Q_ASSIGN U29229 ( .B(clk), .A(\g.we_clk [3545]));
Q_ASSIGN U29230 ( .B(clk), .A(\g.we_clk [3544]));
Q_ASSIGN U29231 ( .B(clk), .A(\g.we_clk [3543]));
Q_ASSIGN U29232 ( .B(clk), .A(\g.we_clk [3542]));
Q_ASSIGN U29233 ( .B(clk), .A(\g.we_clk [3541]));
Q_ASSIGN U29234 ( .B(clk), .A(\g.we_clk [3540]));
Q_ASSIGN U29235 ( .B(clk), .A(\g.we_clk [3539]));
Q_ASSIGN U29236 ( .B(clk), .A(\g.we_clk [3538]));
Q_ASSIGN U29237 ( .B(clk), .A(\g.we_clk [3537]));
Q_ASSIGN U29238 ( .B(clk), .A(\g.we_clk [3536]));
Q_ASSIGN U29239 ( .B(clk), .A(\g.we_clk [3535]));
Q_ASSIGN U29240 ( .B(clk), .A(\g.we_clk [3534]));
Q_ASSIGN U29241 ( .B(clk), .A(\g.we_clk [3533]));
Q_ASSIGN U29242 ( .B(clk), .A(\g.we_clk [3532]));
Q_ASSIGN U29243 ( .B(clk), .A(\g.we_clk [3531]));
Q_ASSIGN U29244 ( .B(clk), .A(\g.we_clk [3530]));
Q_ASSIGN U29245 ( .B(clk), .A(\g.we_clk [3529]));
Q_ASSIGN U29246 ( .B(clk), .A(\g.we_clk [3528]));
Q_ASSIGN U29247 ( .B(clk), .A(\g.we_clk [3527]));
Q_ASSIGN U29248 ( .B(clk), .A(\g.we_clk [3526]));
Q_ASSIGN U29249 ( .B(clk), .A(\g.we_clk [3525]));
Q_ASSIGN U29250 ( .B(clk), .A(\g.we_clk [3524]));
Q_ASSIGN U29251 ( .B(clk), .A(\g.we_clk [3523]));
Q_ASSIGN U29252 ( .B(clk), .A(\g.we_clk [3522]));
Q_ASSIGN U29253 ( .B(clk), .A(\g.we_clk [3521]));
Q_ASSIGN U29254 ( .B(clk), .A(\g.we_clk [3520]));
Q_ASSIGN U29255 ( .B(clk), .A(\g.we_clk [3519]));
Q_ASSIGN U29256 ( .B(clk), .A(\g.we_clk [3518]));
Q_ASSIGN U29257 ( .B(clk), .A(\g.we_clk [3517]));
Q_ASSIGN U29258 ( .B(clk), .A(\g.we_clk [3516]));
Q_ASSIGN U29259 ( .B(clk), .A(\g.we_clk [3515]));
Q_ASSIGN U29260 ( .B(clk), .A(\g.we_clk [3514]));
Q_ASSIGN U29261 ( .B(clk), .A(\g.we_clk [3513]));
Q_ASSIGN U29262 ( .B(clk), .A(\g.we_clk [3512]));
Q_ASSIGN U29263 ( .B(clk), .A(\g.we_clk [3511]));
Q_ASSIGN U29264 ( .B(clk), .A(\g.we_clk [3510]));
Q_ASSIGN U29265 ( .B(clk), .A(\g.we_clk [3509]));
Q_ASSIGN U29266 ( .B(clk), .A(\g.we_clk [3508]));
Q_ASSIGN U29267 ( .B(clk), .A(\g.we_clk [3507]));
Q_ASSIGN U29268 ( .B(clk), .A(\g.we_clk [3506]));
Q_ASSIGN U29269 ( .B(clk), .A(\g.we_clk [3505]));
Q_ASSIGN U29270 ( .B(clk), .A(\g.we_clk [3504]));
Q_ASSIGN U29271 ( .B(clk), .A(\g.we_clk [3503]));
Q_ASSIGN U29272 ( .B(clk), .A(\g.we_clk [3502]));
Q_ASSIGN U29273 ( .B(clk), .A(\g.we_clk [3501]));
Q_ASSIGN U29274 ( .B(clk), .A(\g.we_clk [3500]));
Q_ASSIGN U29275 ( .B(clk), .A(\g.we_clk [3499]));
Q_ASSIGN U29276 ( .B(clk), .A(\g.we_clk [3498]));
Q_ASSIGN U29277 ( .B(clk), .A(\g.we_clk [3497]));
Q_ASSIGN U29278 ( .B(clk), .A(\g.we_clk [3496]));
Q_ASSIGN U29279 ( .B(clk), .A(\g.we_clk [3495]));
Q_ASSIGN U29280 ( .B(clk), .A(\g.we_clk [3494]));
Q_ASSIGN U29281 ( .B(clk), .A(\g.we_clk [3493]));
Q_ASSIGN U29282 ( .B(clk), .A(\g.we_clk [3492]));
Q_ASSIGN U29283 ( .B(clk), .A(\g.we_clk [3491]));
Q_ASSIGN U29284 ( .B(clk), .A(\g.we_clk [3490]));
Q_ASSIGN U29285 ( .B(clk), .A(\g.we_clk [3489]));
Q_ASSIGN U29286 ( .B(clk), .A(\g.we_clk [3488]));
Q_ASSIGN U29287 ( .B(clk), .A(\g.we_clk [3487]));
Q_ASSIGN U29288 ( .B(clk), .A(\g.we_clk [3486]));
Q_ASSIGN U29289 ( .B(clk), .A(\g.we_clk [3485]));
Q_ASSIGN U29290 ( .B(clk), .A(\g.we_clk [3484]));
Q_ASSIGN U29291 ( .B(clk), .A(\g.we_clk [3483]));
Q_ASSIGN U29292 ( .B(clk), .A(\g.we_clk [3482]));
Q_ASSIGN U29293 ( .B(clk), .A(\g.we_clk [3481]));
Q_ASSIGN U29294 ( .B(clk), .A(\g.we_clk [3480]));
Q_ASSIGN U29295 ( .B(clk), .A(\g.we_clk [3479]));
Q_ASSIGN U29296 ( .B(clk), .A(\g.we_clk [3478]));
Q_ASSIGN U29297 ( .B(clk), .A(\g.we_clk [3477]));
Q_ASSIGN U29298 ( .B(clk), .A(\g.we_clk [3476]));
Q_ASSIGN U29299 ( .B(clk), .A(\g.we_clk [3475]));
Q_ASSIGN U29300 ( .B(clk), .A(\g.we_clk [3474]));
Q_ASSIGN U29301 ( .B(clk), .A(\g.we_clk [3473]));
Q_ASSIGN U29302 ( .B(clk), .A(\g.we_clk [3472]));
Q_ASSIGN U29303 ( .B(clk), .A(\g.we_clk [3471]));
Q_ASSIGN U29304 ( .B(clk), .A(\g.we_clk [3470]));
Q_ASSIGN U29305 ( .B(clk), .A(\g.we_clk [3469]));
Q_ASSIGN U29306 ( .B(clk), .A(\g.we_clk [3468]));
Q_ASSIGN U29307 ( .B(clk), .A(\g.we_clk [3467]));
Q_ASSIGN U29308 ( .B(clk), .A(\g.we_clk [3466]));
Q_ASSIGN U29309 ( .B(clk), .A(\g.we_clk [3465]));
Q_ASSIGN U29310 ( .B(clk), .A(\g.we_clk [3464]));
Q_ASSIGN U29311 ( .B(clk), .A(\g.we_clk [3463]));
Q_ASSIGN U29312 ( .B(clk), .A(\g.we_clk [3462]));
Q_ASSIGN U29313 ( .B(clk), .A(\g.we_clk [3461]));
Q_ASSIGN U29314 ( .B(clk), .A(\g.we_clk [3460]));
Q_ASSIGN U29315 ( .B(clk), .A(\g.we_clk [3459]));
Q_ASSIGN U29316 ( .B(clk), .A(\g.we_clk [3458]));
Q_ASSIGN U29317 ( .B(clk), .A(\g.we_clk [3457]));
Q_ASSIGN U29318 ( .B(clk), .A(\g.we_clk [3456]));
Q_ASSIGN U29319 ( .B(clk), .A(\g.we_clk [3455]));
Q_ASSIGN U29320 ( .B(clk), .A(\g.we_clk [3454]));
Q_ASSIGN U29321 ( .B(clk), .A(\g.we_clk [3453]));
Q_ASSIGN U29322 ( .B(clk), .A(\g.we_clk [3452]));
Q_ASSIGN U29323 ( .B(clk), .A(\g.we_clk [3451]));
Q_ASSIGN U29324 ( .B(clk), .A(\g.we_clk [3450]));
Q_ASSIGN U29325 ( .B(clk), .A(\g.we_clk [3449]));
Q_ASSIGN U29326 ( .B(clk), .A(\g.we_clk [3448]));
Q_ASSIGN U29327 ( .B(clk), .A(\g.we_clk [3447]));
Q_ASSIGN U29328 ( .B(clk), .A(\g.we_clk [3446]));
Q_ASSIGN U29329 ( .B(clk), .A(\g.we_clk [3445]));
Q_ASSIGN U29330 ( .B(clk), .A(\g.we_clk [3444]));
Q_ASSIGN U29331 ( .B(clk), .A(\g.we_clk [3443]));
Q_ASSIGN U29332 ( .B(clk), .A(\g.we_clk [3442]));
Q_ASSIGN U29333 ( .B(clk), .A(\g.we_clk [3441]));
Q_ASSIGN U29334 ( .B(clk), .A(\g.we_clk [3440]));
Q_ASSIGN U29335 ( .B(clk), .A(\g.we_clk [3439]));
Q_ASSIGN U29336 ( .B(clk), .A(\g.we_clk [3438]));
Q_ASSIGN U29337 ( .B(clk), .A(\g.we_clk [3437]));
Q_ASSIGN U29338 ( .B(clk), .A(\g.we_clk [3436]));
Q_ASSIGN U29339 ( .B(clk), .A(\g.we_clk [3435]));
Q_ASSIGN U29340 ( .B(clk), .A(\g.we_clk [3434]));
Q_ASSIGN U29341 ( .B(clk), .A(\g.we_clk [3433]));
Q_ASSIGN U29342 ( .B(clk), .A(\g.we_clk [3432]));
Q_ASSIGN U29343 ( .B(clk), .A(\g.we_clk [3431]));
Q_ASSIGN U29344 ( .B(clk), .A(\g.we_clk [3430]));
Q_ASSIGN U29345 ( .B(clk), .A(\g.we_clk [3429]));
Q_ASSIGN U29346 ( .B(clk), .A(\g.we_clk [3428]));
Q_ASSIGN U29347 ( .B(clk), .A(\g.we_clk [3427]));
Q_ASSIGN U29348 ( .B(clk), .A(\g.we_clk [3426]));
Q_ASSIGN U29349 ( .B(clk), .A(\g.we_clk [3425]));
Q_ASSIGN U29350 ( .B(clk), .A(\g.we_clk [3424]));
Q_ASSIGN U29351 ( .B(clk), .A(\g.we_clk [3423]));
Q_ASSIGN U29352 ( .B(clk), .A(\g.we_clk [3422]));
Q_ASSIGN U29353 ( .B(clk), .A(\g.we_clk [3421]));
Q_ASSIGN U29354 ( .B(clk), .A(\g.we_clk [3420]));
Q_ASSIGN U29355 ( .B(clk), .A(\g.we_clk [3419]));
Q_ASSIGN U29356 ( .B(clk), .A(\g.we_clk [3418]));
Q_ASSIGN U29357 ( .B(clk), .A(\g.we_clk [3417]));
Q_ASSIGN U29358 ( .B(clk), .A(\g.we_clk [3416]));
Q_ASSIGN U29359 ( .B(clk), .A(\g.we_clk [3415]));
Q_ASSIGN U29360 ( .B(clk), .A(\g.we_clk [3414]));
Q_ASSIGN U29361 ( .B(clk), .A(\g.we_clk [3413]));
Q_ASSIGN U29362 ( .B(clk), .A(\g.we_clk [3412]));
Q_ASSIGN U29363 ( .B(clk), .A(\g.we_clk [3411]));
Q_ASSIGN U29364 ( .B(clk), .A(\g.we_clk [3410]));
Q_ASSIGN U29365 ( .B(clk), .A(\g.we_clk [3409]));
Q_ASSIGN U29366 ( .B(clk), .A(\g.we_clk [3408]));
Q_ASSIGN U29367 ( .B(clk), .A(\g.we_clk [3407]));
Q_ASSIGN U29368 ( .B(clk), .A(\g.we_clk [3406]));
Q_ASSIGN U29369 ( .B(clk), .A(\g.we_clk [3405]));
Q_ASSIGN U29370 ( .B(clk), .A(\g.we_clk [3404]));
Q_ASSIGN U29371 ( .B(clk), .A(\g.we_clk [3403]));
Q_ASSIGN U29372 ( .B(clk), .A(\g.we_clk [3402]));
Q_ASSIGN U29373 ( .B(clk), .A(\g.we_clk [3401]));
Q_ASSIGN U29374 ( .B(clk), .A(\g.we_clk [3400]));
Q_ASSIGN U29375 ( .B(clk), .A(\g.we_clk [3399]));
Q_ASSIGN U29376 ( .B(clk), .A(\g.we_clk [3398]));
Q_ASSIGN U29377 ( .B(clk), .A(\g.we_clk [3397]));
Q_ASSIGN U29378 ( .B(clk), .A(\g.we_clk [3396]));
Q_ASSIGN U29379 ( .B(clk), .A(\g.we_clk [3395]));
Q_ASSIGN U29380 ( .B(clk), .A(\g.we_clk [3394]));
Q_ASSIGN U29381 ( .B(clk), .A(\g.we_clk [3393]));
Q_ASSIGN U29382 ( .B(clk), .A(\g.we_clk [3392]));
Q_ASSIGN U29383 ( .B(clk), .A(\g.we_clk [3391]));
Q_ASSIGN U29384 ( .B(clk), .A(\g.we_clk [3390]));
Q_ASSIGN U29385 ( .B(clk), .A(\g.we_clk [3389]));
Q_ASSIGN U29386 ( .B(clk), .A(\g.we_clk [3388]));
Q_ASSIGN U29387 ( .B(clk), .A(\g.we_clk [3387]));
Q_ASSIGN U29388 ( .B(clk), .A(\g.we_clk [3386]));
Q_ASSIGN U29389 ( .B(clk), .A(\g.we_clk [3385]));
Q_ASSIGN U29390 ( .B(clk), .A(\g.we_clk [3384]));
Q_ASSIGN U29391 ( .B(clk), .A(\g.we_clk [3383]));
Q_ASSIGN U29392 ( .B(clk), .A(\g.we_clk [3382]));
Q_ASSIGN U29393 ( .B(clk), .A(\g.we_clk [3381]));
Q_ASSIGN U29394 ( .B(clk), .A(\g.we_clk [3380]));
Q_ASSIGN U29395 ( .B(clk), .A(\g.we_clk [3379]));
Q_ASSIGN U29396 ( .B(clk), .A(\g.we_clk [3378]));
Q_ASSIGN U29397 ( .B(clk), .A(\g.we_clk [3377]));
Q_ASSIGN U29398 ( .B(clk), .A(\g.we_clk [3376]));
Q_ASSIGN U29399 ( .B(clk), .A(\g.we_clk [3375]));
Q_ASSIGN U29400 ( .B(clk), .A(\g.we_clk [3374]));
Q_ASSIGN U29401 ( .B(clk), .A(\g.we_clk [3373]));
Q_ASSIGN U29402 ( .B(clk), .A(\g.we_clk [3372]));
Q_ASSIGN U29403 ( .B(clk), .A(\g.we_clk [3371]));
Q_ASSIGN U29404 ( .B(clk), .A(\g.we_clk [3370]));
Q_ASSIGN U29405 ( .B(clk), .A(\g.we_clk [3369]));
Q_ASSIGN U29406 ( .B(clk), .A(\g.we_clk [3368]));
Q_ASSIGN U29407 ( .B(clk), .A(\g.we_clk [3367]));
Q_ASSIGN U29408 ( .B(clk), .A(\g.we_clk [3366]));
Q_ASSIGN U29409 ( .B(clk), .A(\g.we_clk [3365]));
Q_ASSIGN U29410 ( .B(clk), .A(\g.we_clk [3364]));
Q_ASSIGN U29411 ( .B(clk), .A(\g.we_clk [3363]));
Q_ASSIGN U29412 ( .B(clk), .A(\g.we_clk [3362]));
Q_ASSIGN U29413 ( .B(clk), .A(\g.we_clk [3361]));
Q_ASSIGN U29414 ( .B(clk), .A(\g.we_clk [3360]));
Q_ASSIGN U29415 ( .B(clk), .A(\g.we_clk [3359]));
Q_ASSIGN U29416 ( .B(clk), .A(\g.we_clk [3358]));
Q_ASSIGN U29417 ( .B(clk), .A(\g.we_clk [3357]));
Q_ASSIGN U29418 ( .B(clk), .A(\g.we_clk [3356]));
Q_ASSIGN U29419 ( .B(clk), .A(\g.we_clk [3355]));
Q_ASSIGN U29420 ( .B(clk), .A(\g.we_clk [3354]));
Q_ASSIGN U29421 ( .B(clk), .A(\g.we_clk [3353]));
Q_ASSIGN U29422 ( .B(clk), .A(\g.we_clk [3352]));
Q_ASSIGN U29423 ( .B(clk), .A(\g.we_clk [3351]));
Q_ASSIGN U29424 ( .B(clk), .A(\g.we_clk [3350]));
Q_ASSIGN U29425 ( .B(clk), .A(\g.we_clk [3349]));
Q_ASSIGN U29426 ( .B(clk), .A(\g.we_clk [3348]));
Q_ASSIGN U29427 ( .B(clk), .A(\g.we_clk [3347]));
Q_ASSIGN U29428 ( .B(clk), .A(\g.we_clk [3346]));
Q_ASSIGN U29429 ( .B(clk), .A(\g.we_clk [3345]));
Q_ASSIGN U29430 ( .B(clk), .A(\g.we_clk [3344]));
Q_ASSIGN U29431 ( .B(clk), .A(\g.we_clk [3343]));
Q_ASSIGN U29432 ( .B(clk), .A(\g.we_clk [3342]));
Q_ASSIGN U29433 ( .B(clk), .A(\g.we_clk [3341]));
Q_ASSIGN U29434 ( .B(clk), .A(\g.we_clk [3340]));
Q_ASSIGN U29435 ( .B(clk), .A(\g.we_clk [3339]));
Q_ASSIGN U29436 ( .B(clk), .A(\g.we_clk [3338]));
Q_ASSIGN U29437 ( .B(clk), .A(\g.we_clk [3337]));
Q_ASSIGN U29438 ( .B(clk), .A(\g.we_clk [3336]));
Q_ASSIGN U29439 ( .B(clk), .A(\g.we_clk [3335]));
Q_ASSIGN U29440 ( .B(clk), .A(\g.we_clk [3334]));
Q_ASSIGN U29441 ( .B(clk), .A(\g.we_clk [3333]));
Q_ASSIGN U29442 ( .B(clk), .A(\g.we_clk [3332]));
Q_ASSIGN U29443 ( .B(clk), .A(\g.we_clk [3331]));
Q_ASSIGN U29444 ( .B(clk), .A(\g.we_clk [3330]));
Q_ASSIGN U29445 ( .B(clk), .A(\g.we_clk [3329]));
Q_ASSIGN U29446 ( .B(clk), .A(\g.we_clk [3328]));
Q_ASSIGN U29447 ( .B(clk), .A(\g.we_clk [3327]));
Q_ASSIGN U29448 ( .B(clk), .A(\g.we_clk [3326]));
Q_ASSIGN U29449 ( .B(clk), .A(\g.we_clk [3325]));
Q_ASSIGN U29450 ( .B(clk), .A(\g.we_clk [3324]));
Q_ASSIGN U29451 ( .B(clk), .A(\g.we_clk [3323]));
Q_ASSIGN U29452 ( .B(clk), .A(\g.we_clk [3322]));
Q_ASSIGN U29453 ( .B(clk), .A(\g.we_clk [3321]));
Q_ASSIGN U29454 ( .B(clk), .A(\g.we_clk [3320]));
Q_ASSIGN U29455 ( .B(clk), .A(\g.we_clk [3319]));
Q_ASSIGN U29456 ( .B(clk), .A(\g.we_clk [3318]));
Q_ASSIGN U29457 ( .B(clk), .A(\g.we_clk [3317]));
Q_ASSIGN U29458 ( .B(clk), .A(\g.we_clk [3316]));
Q_ASSIGN U29459 ( .B(clk), .A(\g.we_clk [3315]));
Q_ASSIGN U29460 ( .B(clk), .A(\g.we_clk [3314]));
Q_ASSIGN U29461 ( .B(clk), .A(\g.we_clk [3313]));
Q_ASSIGN U29462 ( .B(clk), .A(\g.we_clk [3312]));
Q_ASSIGN U29463 ( .B(clk), .A(\g.we_clk [3311]));
Q_ASSIGN U29464 ( .B(clk), .A(\g.we_clk [3310]));
Q_ASSIGN U29465 ( .B(clk), .A(\g.we_clk [3309]));
Q_ASSIGN U29466 ( .B(clk), .A(\g.we_clk [3308]));
Q_ASSIGN U29467 ( .B(clk), .A(\g.we_clk [3307]));
Q_ASSIGN U29468 ( .B(clk), .A(\g.we_clk [3306]));
Q_ASSIGN U29469 ( .B(clk), .A(\g.we_clk [3305]));
Q_ASSIGN U29470 ( .B(clk), .A(\g.we_clk [3304]));
Q_ASSIGN U29471 ( .B(clk), .A(\g.we_clk [3303]));
Q_ASSIGN U29472 ( .B(clk), .A(\g.we_clk [3302]));
Q_ASSIGN U29473 ( .B(clk), .A(\g.we_clk [3301]));
Q_ASSIGN U29474 ( .B(clk), .A(\g.we_clk [3300]));
Q_ASSIGN U29475 ( .B(clk), .A(\g.we_clk [3299]));
Q_ASSIGN U29476 ( .B(clk), .A(\g.we_clk [3298]));
Q_ASSIGN U29477 ( .B(clk), .A(\g.we_clk [3297]));
Q_ASSIGN U29478 ( .B(clk), .A(\g.we_clk [3296]));
Q_ASSIGN U29479 ( .B(clk), .A(\g.we_clk [3295]));
Q_ASSIGN U29480 ( .B(clk), .A(\g.we_clk [3294]));
Q_ASSIGN U29481 ( .B(clk), .A(\g.we_clk [3293]));
Q_ASSIGN U29482 ( .B(clk), .A(\g.we_clk [3292]));
Q_ASSIGN U29483 ( .B(clk), .A(\g.we_clk [3291]));
Q_ASSIGN U29484 ( .B(clk), .A(\g.we_clk [3290]));
Q_ASSIGN U29485 ( .B(clk), .A(\g.we_clk [3289]));
Q_ASSIGN U29486 ( .B(clk), .A(\g.we_clk [3288]));
Q_ASSIGN U29487 ( .B(clk), .A(\g.we_clk [3287]));
Q_ASSIGN U29488 ( .B(clk), .A(\g.we_clk [3286]));
Q_ASSIGN U29489 ( .B(clk), .A(\g.we_clk [3285]));
Q_ASSIGN U29490 ( .B(clk), .A(\g.we_clk [3284]));
Q_ASSIGN U29491 ( .B(clk), .A(\g.we_clk [3283]));
Q_ASSIGN U29492 ( .B(clk), .A(\g.we_clk [3282]));
Q_ASSIGN U29493 ( .B(clk), .A(\g.we_clk [3281]));
Q_ASSIGN U29494 ( .B(clk), .A(\g.we_clk [3280]));
Q_ASSIGN U29495 ( .B(clk), .A(\g.we_clk [3279]));
Q_ASSIGN U29496 ( .B(clk), .A(\g.we_clk [3278]));
Q_ASSIGN U29497 ( .B(clk), .A(\g.we_clk [3277]));
Q_ASSIGN U29498 ( .B(clk), .A(\g.we_clk [3276]));
Q_ASSIGN U29499 ( .B(clk), .A(\g.we_clk [3275]));
Q_ASSIGN U29500 ( .B(clk), .A(\g.we_clk [3274]));
Q_ASSIGN U29501 ( .B(clk), .A(\g.we_clk [3273]));
Q_ASSIGN U29502 ( .B(clk), .A(\g.we_clk [3272]));
Q_ASSIGN U29503 ( .B(clk), .A(\g.we_clk [3271]));
Q_ASSIGN U29504 ( .B(clk), .A(\g.we_clk [3270]));
Q_ASSIGN U29505 ( .B(clk), .A(\g.we_clk [3269]));
Q_ASSIGN U29506 ( .B(clk), .A(\g.we_clk [3268]));
Q_ASSIGN U29507 ( .B(clk), .A(\g.we_clk [3267]));
Q_ASSIGN U29508 ( .B(clk), .A(\g.we_clk [3266]));
Q_ASSIGN U29509 ( .B(clk), .A(\g.we_clk [3265]));
Q_ASSIGN U29510 ( .B(clk), .A(\g.we_clk [3264]));
Q_ASSIGN U29511 ( .B(clk), .A(\g.we_clk [3263]));
Q_ASSIGN U29512 ( .B(clk), .A(\g.we_clk [3262]));
Q_ASSIGN U29513 ( .B(clk), .A(\g.we_clk [3261]));
Q_ASSIGN U29514 ( .B(clk), .A(\g.we_clk [3260]));
Q_ASSIGN U29515 ( .B(clk), .A(\g.we_clk [3259]));
Q_ASSIGN U29516 ( .B(clk), .A(\g.we_clk [3258]));
Q_ASSIGN U29517 ( .B(clk), .A(\g.we_clk [3257]));
Q_ASSIGN U29518 ( .B(clk), .A(\g.we_clk [3256]));
Q_ASSIGN U29519 ( .B(clk), .A(\g.we_clk [3255]));
Q_ASSIGN U29520 ( .B(clk), .A(\g.we_clk [3254]));
Q_ASSIGN U29521 ( .B(clk), .A(\g.we_clk [3253]));
Q_ASSIGN U29522 ( .B(clk), .A(\g.we_clk [3252]));
Q_ASSIGN U29523 ( .B(clk), .A(\g.we_clk [3251]));
Q_ASSIGN U29524 ( .B(clk), .A(\g.we_clk [3250]));
Q_ASSIGN U29525 ( .B(clk), .A(\g.we_clk [3249]));
Q_ASSIGN U29526 ( .B(clk), .A(\g.we_clk [3248]));
Q_ASSIGN U29527 ( .B(clk), .A(\g.we_clk [3247]));
Q_ASSIGN U29528 ( .B(clk), .A(\g.we_clk [3246]));
Q_ASSIGN U29529 ( .B(clk), .A(\g.we_clk [3245]));
Q_ASSIGN U29530 ( .B(clk), .A(\g.we_clk [3244]));
Q_ASSIGN U29531 ( .B(clk), .A(\g.we_clk [3243]));
Q_ASSIGN U29532 ( .B(clk), .A(\g.we_clk [3242]));
Q_ASSIGN U29533 ( .B(clk), .A(\g.we_clk [3241]));
Q_ASSIGN U29534 ( .B(clk), .A(\g.we_clk [3240]));
Q_ASSIGN U29535 ( .B(clk), .A(\g.we_clk [3239]));
Q_ASSIGN U29536 ( .B(clk), .A(\g.we_clk [3238]));
Q_ASSIGN U29537 ( .B(clk), .A(\g.we_clk [3237]));
Q_ASSIGN U29538 ( .B(clk), .A(\g.we_clk [3236]));
Q_ASSIGN U29539 ( .B(clk), .A(\g.we_clk [3235]));
Q_ASSIGN U29540 ( .B(clk), .A(\g.we_clk [3234]));
Q_ASSIGN U29541 ( .B(clk), .A(\g.we_clk [3233]));
Q_ASSIGN U29542 ( .B(clk), .A(\g.we_clk [3232]));
Q_ASSIGN U29543 ( .B(clk), .A(\g.we_clk [3231]));
Q_ASSIGN U29544 ( .B(clk), .A(\g.we_clk [3230]));
Q_ASSIGN U29545 ( .B(clk), .A(\g.we_clk [3229]));
Q_ASSIGN U29546 ( .B(clk), .A(\g.we_clk [3228]));
Q_ASSIGN U29547 ( .B(clk), .A(\g.we_clk [3227]));
Q_ASSIGN U29548 ( .B(clk), .A(\g.we_clk [3226]));
Q_ASSIGN U29549 ( .B(clk), .A(\g.we_clk [3225]));
Q_ASSIGN U29550 ( .B(clk), .A(\g.we_clk [3224]));
Q_ASSIGN U29551 ( .B(clk), .A(\g.we_clk [3223]));
Q_ASSIGN U29552 ( .B(clk), .A(\g.we_clk [3222]));
Q_ASSIGN U29553 ( .B(clk), .A(\g.we_clk [3221]));
Q_ASSIGN U29554 ( .B(clk), .A(\g.we_clk [3220]));
Q_ASSIGN U29555 ( .B(clk), .A(\g.we_clk [3219]));
Q_ASSIGN U29556 ( .B(clk), .A(\g.we_clk [3218]));
Q_ASSIGN U29557 ( .B(clk), .A(\g.we_clk [3217]));
Q_ASSIGN U29558 ( .B(clk), .A(\g.we_clk [3216]));
Q_ASSIGN U29559 ( .B(clk), .A(\g.we_clk [3215]));
Q_ASSIGN U29560 ( .B(clk), .A(\g.we_clk [3214]));
Q_ASSIGN U29561 ( .B(clk), .A(\g.we_clk [3213]));
Q_ASSIGN U29562 ( .B(clk), .A(\g.we_clk [3212]));
Q_ASSIGN U29563 ( .B(clk), .A(\g.we_clk [3211]));
Q_ASSIGN U29564 ( .B(clk), .A(\g.we_clk [3210]));
Q_ASSIGN U29565 ( .B(clk), .A(\g.we_clk [3209]));
Q_ASSIGN U29566 ( .B(clk), .A(\g.we_clk [3208]));
Q_ASSIGN U29567 ( .B(clk), .A(\g.we_clk [3207]));
Q_ASSIGN U29568 ( .B(clk), .A(\g.we_clk [3206]));
Q_ASSIGN U29569 ( .B(clk), .A(\g.we_clk [3205]));
Q_ASSIGN U29570 ( .B(clk), .A(\g.we_clk [3204]));
Q_ASSIGN U29571 ( .B(clk), .A(\g.we_clk [3203]));
Q_ASSIGN U29572 ( .B(clk), .A(\g.we_clk [3202]));
Q_ASSIGN U29573 ( .B(clk), .A(\g.we_clk [3201]));
Q_ASSIGN U29574 ( .B(clk), .A(\g.we_clk [3200]));
Q_ASSIGN U29575 ( .B(clk), .A(\g.we_clk [3199]));
Q_ASSIGN U29576 ( .B(clk), .A(\g.we_clk [3198]));
Q_ASSIGN U29577 ( .B(clk), .A(\g.we_clk [3197]));
Q_ASSIGN U29578 ( .B(clk), .A(\g.we_clk [3196]));
Q_ASSIGN U29579 ( .B(clk), .A(\g.we_clk [3195]));
Q_ASSIGN U29580 ( .B(clk), .A(\g.we_clk [3194]));
Q_ASSIGN U29581 ( .B(clk), .A(\g.we_clk [3193]));
Q_ASSIGN U29582 ( .B(clk), .A(\g.we_clk [3192]));
Q_ASSIGN U29583 ( .B(clk), .A(\g.we_clk [3191]));
Q_ASSIGN U29584 ( .B(clk), .A(\g.we_clk [3190]));
Q_ASSIGN U29585 ( .B(clk), .A(\g.we_clk [3189]));
Q_ASSIGN U29586 ( .B(clk), .A(\g.we_clk [3188]));
Q_ASSIGN U29587 ( .B(clk), .A(\g.we_clk [3187]));
Q_ASSIGN U29588 ( .B(clk), .A(\g.we_clk [3186]));
Q_ASSIGN U29589 ( .B(clk), .A(\g.we_clk [3185]));
Q_ASSIGN U29590 ( .B(clk), .A(\g.we_clk [3184]));
Q_ASSIGN U29591 ( .B(clk), .A(\g.we_clk [3183]));
Q_ASSIGN U29592 ( .B(clk), .A(\g.we_clk [3182]));
Q_ASSIGN U29593 ( .B(clk), .A(\g.we_clk [3181]));
Q_ASSIGN U29594 ( .B(clk), .A(\g.we_clk [3180]));
Q_ASSIGN U29595 ( .B(clk), .A(\g.we_clk [3179]));
Q_ASSIGN U29596 ( .B(clk), .A(\g.we_clk [3178]));
Q_ASSIGN U29597 ( .B(clk), .A(\g.we_clk [3177]));
Q_ASSIGN U29598 ( .B(clk), .A(\g.we_clk [3176]));
Q_ASSIGN U29599 ( .B(clk), .A(\g.we_clk [3175]));
Q_ASSIGN U29600 ( .B(clk), .A(\g.we_clk [3174]));
Q_ASSIGN U29601 ( .B(clk), .A(\g.we_clk [3173]));
Q_ASSIGN U29602 ( .B(clk), .A(\g.we_clk [3172]));
Q_ASSIGN U29603 ( .B(clk), .A(\g.we_clk [3171]));
Q_ASSIGN U29604 ( .B(clk), .A(\g.we_clk [3170]));
Q_ASSIGN U29605 ( .B(clk), .A(\g.we_clk [3169]));
Q_ASSIGN U29606 ( .B(clk), .A(\g.we_clk [3168]));
Q_ASSIGN U29607 ( .B(clk), .A(\g.we_clk [3167]));
Q_ASSIGN U29608 ( .B(clk), .A(\g.we_clk [3166]));
Q_ASSIGN U29609 ( .B(clk), .A(\g.we_clk [3165]));
Q_ASSIGN U29610 ( .B(clk), .A(\g.we_clk [3164]));
Q_ASSIGN U29611 ( .B(clk), .A(\g.we_clk [3163]));
Q_ASSIGN U29612 ( .B(clk), .A(\g.we_clk [3162]));
Q_ASSIGN U29613 ( .B(clk), .A(\g.we_clk [3161]));
Q_ASSIGN U29614 ( .B(clk), .A(\g.we_clk [3160]));
Q_ASSIGN U29615 ( .B(clk), .A(\g.we_clk [3159]));
Q_ASSIGN U29616 ( .B(clk), .A(\g.we_clk [3158]));
Q_ASSIGN U29617 ( .B(clk), .A(\g.we_clk [3157]));
Q_ASSIGN U29618 ( .B(clk), .A(\g.we_clk [3156]));
Q_ASSIGN U29619 ( .B(clk), .A(\g.we_clk [3155]));
Q_ASSIGN U29620 ( .B(clk), .A(\g.we_clk [3154]));
Q_ASSIGN U29621 ( .B(clk), .A(\g.we_clk [3153]));
Q_ASSIGN U29622 ( .B(clk), .A(\g.we_clk [3152]));
Q_ASSIGN U29623 ( .B(clk), .A(\g.we_clk [3151]));
Q_ASSIGN U29624 ( .B(clk), .A(\g.we_clk [3150]));
Q_ASSIGN U29625 ( .B(clk), .A(\g.we_clk [3149]));
Q_ASSIGN U29626 ( .B(clk), .A(\g.we_clk [3148]));
Q_ASSIGN U29627 ( .B(clk), .A(\g.we_clk [3147]));
Q_ASSIGN U29628 ( .B(clk), .A(\g.we_clk [3146]));
Q_ASSIGN U29629 ( .B(clk), .A(\g.we_clk [3145]));
Q_ASSIGN U29630 ( .B(clk), .A(\g.we_clk [3144]));
Q_ASSIGN U29631 ( .B(clk), .A(\g.we_clk [3143]));
Q_ASSIGN U29632 ( .B(clk), .A(\g.we_clk [3142]));
Q_ASSIGN U29633 ( .B(clk), .A(\g.we_clk [3141]));
Q_ASSIGN U29634 ( .B(clk), .A(\g.we_clk [3140]));
Q_ASSIGN U29635 ( .B(clk), .A(\g.we_clk [3139]));
Q_ASSIGN U29636 ( .B(clk), .A(\g.we_clk [3138]));
Q_ASSIGN U29637 ( .B(clk), .A(\g.we_clk [3137]));
Q_ASSIGN U29638 ( .B(clk), .A(\g.we_clk [3136]));
Q_ASSIGN U29639 ( .B(clk), .A(\g.we_clk [3135]));
Q_ASSIGN U29640 ( .B(clk), .A(\g.we_clk [3134]));
Q_ASSIGN U29641 ( .B(clk), .A(\g.we_clk [3133]));
Q_ASSIGN U29642 ( .B(clk), .A(\g.we_clk [3132]));
Q_ASSIGN U29643 ( .B(clk), .A(\g.we_clk [3131]));
Q_ASSIGN U29644 ( .B(clk), .A(\g.we_clk [3130]));
Q_ASSIGN U29645 ( .B(clk), .A(\g.we_clk [3129]));
Q_ASSIGN U29646 ( .B(clk), .A(\g.we_clk [3128]));
Q_ASSIGN U29647 ( .B(clk), .A(\g.we_clk [3127]));
Q_ASSIGN U29648 ( .B(clk), .A(\g.we_clk [3126]));
Q_ASSIGN U29649 ( .B(clk), .A(\g.we_clk [3125]));
Q_ASSIGN U29650 ( .B(clk), .A(\g.we_clk [3124]));
Q_ASSIGN U29651 ( .B(clk), .A(\g.we_clk [3123]));
Q_ASSIGN U29652 ( .B(clk), .A(\g.we_clk [3122]));
Q_ASSIGN U29653 ( .B(clk), .A(\g.we_clk [3121]));
Q_ASSIGN U29654 ( .B(clk), .A(\g.we_clk [3120]));
Q_ASSIGN U29655 ( .B(clk), .A(\g.we_clk [3119]));
Q_ASSIGN U29656 ( .B(clk), .A(\g.we_clk [3118]));
Q_ASSIGN U29657 ( .B(clk), .A(\g.we_clk [3117]));
Q_ASSIGN U29658 ( .B(clk), .A(\g.we_clk [3116]));
Q_ASSIGN U29659 ( .B(clk), .A(\g.we_clk [3115]));
Q_ASSIGN U29660 ( .B(clk), .A(\g.we_clk [3114]));
Q_ASSIGN U29661 ( .B(clk), .A(\g.we_clk [3113]));
Q_ASSIGN U29662 ( .B(clk), .A(\g.we_clk [3112]));
Q_ASSIGN U29663 ( .B(clk), .A(\g.we_clk [3111]));
Q_ASSIGN U29664 ( .B(clk), .A(\g.we_clk [3110]));
Q_ASSIGN U29665 ( .B(clk), .A(\g.we_clk [3109]));
Q_ASSIGN U29666 ( .B(clk), .A(\g.we_clk [3108]));
Q_ASSIGN U29667 ( .B(clk), .A(\g.we_clk [3107]));
Q_ASSIGN U29668 ( .B(clk), .A(\g.we_clk [3106]));
Q_ASSIGN U29669 ( .B(clk), .A(\g.we_clk [3105]));
Q_ASSIGN U29670 ( .B(clk), .A(\g.we_clk [3104]));
Q_ASSIGN U29671 ( .B(clk), .A(\g.we_clk [3103]));
Q_ASSIGN U29672 ( .B(clk), .A(\g.we_clk [3102]));
Q_ASSIGN U29673 ( .B(clk), .A(\g.we_clk [3101]));
Q_ASSIGN U29674 ( .B(clk), .A(\g.we_clk [3100]));
Q_ASSIGN U29675 ( .B(clk), .A(\g.we_clk [3099]));
Q_ASSIGN U29676 ( .B(clk), .A(\g.we_clk [3098]));
Q_ASSIGN U29677 ( .B(clk), .A(\g.we_clk [3097]));
Q_ASSIGN U29678 ( .B(clk), .A(\g.we_clk [3096]));
Q_ASSIGN U29679 ( .B(clk), .A(\g.we_clk [3095]));
Q_ASSIGN U29680 ( .B(clk), .A(\g.we_clk [3094]));
Q_ASSIGN U29681 ( .B(clk), .A(\g.we_clk [3093]));
Q_ASSIGN U29682 ( .B(clk), .A(\g.we_clk [3092]));
Q_ASSIGN U29683 ( .B(clk), .A(\g.we_clk [3091]));
Q_ASSIGN U29684 ( .B(clk), .A(\g.we_clk [3090]));
Q_ASSIGN U29685 ( .B(clk), .A(\g.we_clk [3089]));
Q_ASSIGN U29686 ( .B(clk), .A(\g.we_clk [3088]));
Q_ASSIGN U29687 ( .B(clk), .A(\g.we_clk [3087]));
Q_ASSIGN U29688 ( .B(clk), .A(\g.we_clk [3086]));
Q_ASSIGN U29689 ( .B(clk), .A(\g.we_clk [3085]));
Q_ASSIGN U29690 ( .B(clk), .A(\g.we_clk [3084]));
Q_ASSIGN U29691 ( .B(clk), .A(\g.we_clk [3083]));
Q_ASSIGN U29692 ( .B(clk), .A(\g.we_clk [3082]));
Q_ASSIGN U29693 ( .B(clk), .A(\g.we_clk [3081]));
Q_ASSIGN U29694 ( .B(clk), .A(\g.we_clk [3080]));
Q_ASSIGN U29695 ( .B(clk), .A(\g.we_clk [3079]));
Q_ASSIGN U29696 ( .B(clk), .A(\g.we_clk [3078]));
Q_ASSIGN U29697 ( .B(clk), .A(\g.we_clk [3077]));
Q_ASSIGN U29698 ( .B(clk), .A(\g.we_clk [3076]));
Q_ASSIGN U29699 ( .B(clk), .A(\g.we_clk [3075]));
Q_ASSIGN U29700 ( .B(clk), .A(\g.we_clk [3074]));
Q_ASSIGN U29701 ( .B(clk), .A(\g.we_clk [3073]));
Q_ASSIGN U29702 ( .B(clk), .A(\g.we_clk [3072]));
Q_ASSIGN U29703 ( .B(clk), .A(\g.we_clk [3071]));
Q_ASSIGN U29704 ( .B(clk), .A(\g.we_clk [3070]));
Q_ASSIGN U29705 ( .B(clk), .A(\g.we_clk [3069]));
Q_ASSIGN U29706 ( .B(clk), .A(\g.we_clk [3068]));
Q_ASSIGN U29707 ( .B(clk), .A(\g.we_clk [3067]));
Q_ASSIGN U29708 ( .B(clk), .A(\g.we_clk [3066]));
Q_ASSIGN U29709 ( .B(clk), .A(\g.we_clk [3065]));
Q_ASSIGN U29710 ( .B(clk), .A(\g.we_clk [3064]));
Q_ASSIGN U29711 ( .B(clk), .A(\g.we_clk [3063]));
Q_ASSIGN U29712 ( .B(clk), .A(\g.we_clk [3062]));
Q_ASSIGN U29713 ( .B(clk), .A(\g.we_clk [3061]));
Q_ASSIGN U29714 ( .B(clk), .A(\g.we_clk [3060]));
Q_ASSIGN U29715 ( .B(clk), .A(\g.we_clk [3059]));
Q_ASSIGN U29716 ( .B(clk), .A(\g.we_clk [3058]));
Q_ASSIGN U29717 ( .B(clk), .A(\g.we_clk [3057]));
Q_ASSIGN U29718 ( .B(clk), .A(\g.we_clk [3056]));
Q_ASSIGN U29719 ( .B(clk), .A(\g.we_clk [3055]));
Q_ASSIGN U29720 ( .B(clk), .A(\g.we_clk [3054]));
Q_ASSIGN U29721 ( .B(clk), .A(\g.we_clk [3053]));
Q_ASSIGN U29722 ( .B(clk), .A(\g.we_clk [3052]));
Q_ASSIGN U29723 ( .B(clk), .A(\g.we_clk [3051]));
Q_ASSIGN U29724 ( .B(clk), .A(\g.we_clk [3050]));
Q_ASSIGN U29725 ( .B(clk), .A(\g.we_clk [3049]));
Q_ASSIGN U29726 ( .B(clk), .A(\g.we_clk [3048]));
Q_ASSIGN U29727 ( .B(clk), .A(\g.we_clk [3047]));
Q_ASSIGN U29728 ( .B(clk), .A(\g.we_clk [3046]));
Q_ASSIGN U29729 ( .B(clk), .A(\g.we_clk [3045]));
Q_ASSIGN U29730 ( .B(clk), .A(\g.we_clk [3044]));
Q_ASSIGN U29731 ( .B(clk), .A(\g.we_clk [3043]));
Q_ASSIGN U29732 ( .B(clk), .A(\g.we_clk [3042]));
Q_ASSIGN U29733 ( .B(clk), .A(\g.we_clk [3041]));
Q_ASSIGN U29734 ( .B(clk), .A(\g.we_clk [3040]));
Q_ASSIGN U29735 ( .B(clk), .A(\g.we_clk [3039]));
Q_ASSIGN U29736 ( .B(clk), .A(\g.we_clk [3038]));
Q_ASSIGN U29737 ( .B(clk), .A(\g.we_clk [3037]));
Q_ASSIGN U29738 ( .B(clk), .A(\g.we_clk [3036]));
Q_ASSIGN U29739 ( .B(clk), .A(\g.we_clk [3035]));
Q_ASSIGN U29740 ( .B(clk), .A(\g.we_clk [3034]));
Q_ASSIGN U29741 ( .B(clk), .A(\g.we_clk [3033]));
Q_ASSIGN U29742 ( .B(clk), .A(\g.we_clk [3032]));
Q_ASSIGN U29743 ( .B(clk), .A(\g.we_clk [3031]));
Q_ASSIGN U29744 ( .B(clk), .A(\g.we_clk [3030]));
Q_ASSIGN U29745 ( .B(clk), .A(\g.we_clk [3029]));
Q_ASSIGN U29746 ( .B(clk), .A(\g.we_clk [3028]));
Q_ASSIGN U29747 ( .B(clk), .A(\g.we_clk [3027]));
Q_ASSIGN U29748 ( .B(clk), .A(\g.we_clk [3026]));
Q_ASSIGN U29749 ( .B(clk), .A(\g.we_clk [3025]));
Q_ASSIGN U29750 ( .B(clk), .A(\g.we_clk [3024]));
Q_ASSIGN U29751 ( .B(clk), .A(\g.we_clk [3023]));
Q_ASSIGN U29752 ( .B(clk), .A(\g.we_clk [3022]));
Q_ASSIGN U29753 ( .B(clk), .A(\g.we_clk [3021]));
Q_ASSIGN U29754 ( .B(clk), .A(\g.we_clk [3020]));
Q_ASSIGN U29755 ( .B(clk), .A(\g.we_clk [3019]));
Q_ASSIGN U29756 ( .B(clk), .A(\g.we_clk [3018]));
Q_ASSIGN U29757 ( .B(clk), .A(\g.we_clk [3017]));
Q_ASSIGN U29758 ( .B(clk), .A(\g.we_clk [3016]));
Q_ASSIGN U29759 ( .B(clk), .A(\g.we_clk [3015]));
Q_ASSIGN U29760 ( .B(clk), .A(\g.we_clk [3014]));
Q_ASSIGN U29761 ( .B(clk), .A(\g.we_clk [3013]));
Q_ASSIGN U29762 ( .B(clk), .A(\g.we_clk [3012]));
Q_ASSIGN U29763 ( .B(clk), .A(\g.we_clk [3011]));
Q_ASSIGN U29764 ( .B(clk), .A(\g.we_clk [3010]));
Q_ASSIGN U29765 ( .B(clk), .A(\g.we_clk [3009]));
Q_ASSIGN U29766 ( .B(clk), .A(\g.we_clk [3008]));
Q_ASSIGN U29767 ( .B(clk), .A(\g.we_clk [3007]));
Q_ASSIGN U29768 ( .B(clk), .A(\g.we_clk [3006]));
Q_ASSIGN U29769 ( .B(clk), .A(\g.we_clk [3005]));
Q_ASSIGN U29770 ( .B(clk), .A(\g.we_clk [3004]));
Q_ASSIGN U29771 ( .B(clk), .A(\g.we_clk [3003]));
Q_ASSIGN U29772 ( .B(clk), .A(\g.we_clk [3002]));
Q_ASSIGN U29773 ( .B(clk), .A(\g.we_clk [3001]));
Q_ASSIGN U29774 ( .B(clk), .A(\g.we_clk [3000]));
Q_ASSIGN U29775 ( .B(clk), .A(\g.we_clk [2999]));
Q_ASSIGN U29776 ( .B(clk), .A(\g.we_clk [2998]));
Q_ASSIGN U29777 ( .B(clk), .A(\g.we_clk [2997]));
Q_ASSIGN U29778 ( .B(clk), .A(\g.we_clk [2996]));
Q_ASSIGN U29779 ( .B(clk), .A(\g.we_clk [2995]));
Q_ASSIGN U29780 ( .B(clk), .A(\g.we_clk [2994]));
Q_ASSIGN U29781 ( .B(clk), .A(\g.we_clk [2993]));
Q_ASSIGN U29782 ( .B(clk), .A(\g.we_clk [2992]));
Q_ASSIGN U29783 ( .B(clk), .A(\g.we_clk [2991]));
Q_ASSIGN U29784 ( .B(clk), .A(\g.we_clk [2990]));
Q_ASSIGN U29785 ( .B(clk), .A(\g.we_clk [2989]));
Q_ASSIGN U29786 ( .B(clk), .A(\g.we_clk [2988]));
Q_ASSIGN U29787 ( .B(clk), .A(\g.we_clk [2987]));
Q_ASSIGN U29788 ( .B(clk), .A(\g.we_clk [2986]));
Q_ASSIGN U29789 ( .B(clk), .A(\g.we_clk [2985]));
Q_ASSIGN U29790 ( .B(clk), .A(\g.we_clk [2984]));
Q_ASSIGN U29791 ( .B(clk), .A(\g.we_clk [2983]));
Q_ASSIGN U29792 ( .B(clk), .A(\g.we_clk [2982]));
Q_ASSIGN U29793 ( .B(clk), .A(\g.we_clk [2981]));
Q_ASSIGN U29794 ( .B(clk), .A(\g.we_clk [2980]));
Q_ASSIGN U29795 ( .B(clk), .A(\g.we_clk [2979]));
Q_ASSIGN U29796 ( .B(clk), .A(\g.we_clk [2978]));
Q_ASSIGN U29797 ( .B(clk), .A(\g.we_clk [2977]));
Q_ASSIGN U29798 ( .B(clk), .A(\g.we_clk [2976]));
Q_ASSIGN U29799 ( .B(clk), .A(\g.we_clk [2975]));
Q_ASSIGN U29800 ( .B(clk), .A(\g.we_clk [2974]));
Q_ASSIGN U29801 ( .B(clk), .A(\g.we_clk [2973]));
Q_ASSIGN U29802 ( .B(clk), .A(\g.we_clk [2972]));
Q_ASSIGN U29803 ( .B(clk), .A(\g.we_clk [2971]));
Q_ASSIGN U29804 ( .B(clk), .A(\g.we_clk [2970]));
Q_ASSIGN U29805 ( .B(clk), .A(\g.we_clk [2969]));
Q_ASSIGN U29806 ( .B(clk), .A(\g.we_clk [2968]));
Q_ASSIGN U29807 ( .B(clk), .A(\g.we_clk [2967]));
Q_ASSIGN U29808 ( .B(clk), .A(\g.we_clk [2966]));
Q_ASSIGN U29809 ( .B(clk), .A(\g.we_clk [2965]));
Q_ASSIGN U29810 ( .B(clk), .A(\g.we_clk [2964]));
Q_ASSIGN U29811 ( .B(clk), .A(\g.we_clk [2963]));
Q_ASSIGN U29812 ( .B(clk), .A(\g.we_clk [2962]));
Q_ASSIGN U29813 ( .B(clk), .A(\g.we_clk [2961]));
Q_ASSIGN U29814 ( .B(clk), .A(\g.we_clk [2960]));
Q_ASSIGN U29815 ( .B(clk), .A(\g.we_clk [2959]));
Q_ASSIGN U29816 ( .B(clk), .A(\g.we_clk [2958]));
Q_ASSIGN U29817 ( .B(clk), .A(\g.we_clk [2957]));
Q_ASSIGN U29818 ( .B(clk), .A(\g.we_clk [2956]));
Q_ASSIGN U29819 ( .B(clk), .A(\g.we_clk [2955]));
Q_ASSIGN U29820 ( .B(clk), .A(\g.we_clk [2954]));
Q_ASSIGN U29821 ( .B(clk), .A(\g.we_clk [2953]));
Q_ASSIGN U29822 ( .B(clk), .A(\g.we_clk [2952]));
Q_ASSIGN U29823 ( .B(clk), .A(\g.we_clk [2951]));
Q_ASSIGN U29824 ( .B(clk), .A(\g.we_clk [2950]));
Q_ASSIGN U29825 ( .B(clk), .A(\g.we_clk [2949]));
Q_ASSIGN U29826 ( .B(clk), .A(\g.we_clk [2948]));
Q_ASSIGN U29827 ( .B(clk), .A(\g.we_clk [2947]));
Q_ASSIGN U29828 ( .B(clk), .A(\g.we_clk [2946]));
Q_ASSIGN U29829 ( .B(clk), .A(\g.we_clk [2945]));
Q_ASSIGN U29830 ( .B(clk), .A(\g.we_clk [2944]));
Q_ASSIGN U29831 ( .B(clk), .A(\g.we_clk [2943]));
Q_ASSIGN U29832 ( .B(clk), .A(\g.we_clk [2942]));
Q_ASSIGN U29833 ( .B(clk), .A(\g.we_clk [2941]));
Q_ASSIGN U29834 ( .B(clk), .A(\g.we_clk [2940]));
Q_ASSIGN U29835 ( .B(clk), .A(\g.we_clk [2939]));
Q_ASSIGN U29836 ( .B(clk), .A(\g.we_clk [2938]));
Q_ASSIGN U29837 ( .B(clk), .A(\g.we_clk [2937]));
Q_ASSIGN U29838 ( .B(clk), .A(\g.we_clk [2936]));
Q_ASSIGN U29839 ( .B(clk), .A(\g.we_clk [2935]));
Q_ASSIGN U29840 ( .B(clk), .A(\g.we_clk [2934]));
Q_ASSIGN U29841 ( .B(clk), .A(\g.we_clk [2933]));
Q_ASSIGN U29842 ( .B(clk), .A(\g.we_clk [2932]));
Q_ASSIGN U29843 ( .B(clk), .A(\g.we_clk [2931]));
Q_ASSIGN U29844 ( .B(clk), .A(\g.we_clk [2930]));
Q_ASSIGN U29845 ( .B(clk), .A(\g.we_clk [2929]));
Q_ASSIGN U29846 ( .B(clk), .A(\g.we_clk [2928]));
Q_ASSIGN U29847 ( .B(clk), .A(\g.we_clk [2927]));
Q_ASSIGN U29848 ( .B(clk), .A(\g.we_clk [2926]));
Q_ASSIGN U29849 ( .B(clk), .A(\g.we_clk [2925]));
Q_ASSIGN U29850 ( .B(clk), .A(\g.we_clk [2924]));
Q_ASSIGN U29851 ( .B(clk), .A(\g.we_clk [2923]));
Q_ASSIGN U29852 ( .B(clk), .A(\g.we_clk [2922]));
Q_ASSIGN U29853 ( .B(clk), .A(\g.we_clk [2921]));
Q_ASSIGN U29854 ( .B(clk), .A(\g.we_clk [2920]));
Q_ASSIGN U29855 ( .B(clk), .A(\g.we_clk [2919]));
Q_ASSIGN U29856 ( .B(clk), .A(\g.we_clk [2918]));
Q_ASSIGN U29857 ( .B(clk), .A(\g.we_clk [2917]));
Q_ASSIGN U29858 ( .B(clk), .A(\g.we_clk [2916]));
Q_ASSIGN U29859 ( .B(clk), .A(\g.we_clk [2915]));
Q_ASSIGN U29860 ( .B(clk), .A(\g.we_clk [2914]));
Q_ASSIGN U29861 ( .B(clk), .A(\g.we_clk [2913]));
Q_ASSIGN U29862 ( .B(clk), .A(\g.we_clk [2912]));
Q_ASSIGN U29863 ( .B(clk), .A(\g.we_clk [2911]));
Q_ASSIGN U29864 ( .B(clk), .A(\g.we_clk [2910]));
Q_ASSIGN U29865 ( .B(clk), .A(\g.we_clk [2909]));
Q_ASSIGN U29866 ( .B(clk), .A(\g.we_clk [2908]));
Q_ASSIGN U29867 ( .B(clk), .A(\g.we_clk [2907]));
Q_ASSIGN U29868 ( .B(clk), .A(\g.we_clk [2906]));
Q_ASSIGN U29869 ( .B(clk), .A(\g.we_clk [2905]));
Q_ASSIGN U29870 ( .B(clk), .A(\g.we_clk [2904]));
Q_ASSIGN U29871 ( .B(clk), .A(\g.we_clk [2903]));
Q_ASSIGN U29872 ( .B(clk), .A(\g.we_clk [2902]));
Q_ASSIGN U29873 ( .B(clk), .A(\g.we_clk [2901]));
Q_ASSIGN U29874 ( .B(clk), .A(\g.we_clk [2900]));
Q_ASSIGN U29875 ( .B(clk), .A(\g.we_clk [2899]));
Q_ASSIGN U29876 ( .B(clk), .A(\g.we_clk [2898]));
Q_ASSIGN U29877 ( .B(clk), .A(\g.we_clk [2897]));
Q_ASSIGN U29878 ( .B(clk), .A(\g.we_clk [2896]));
Q_ASSIGN U29879 ( .B(clk), .A(\g.we_clk [2895]));
Q_ASSIGN U29880 ( .B(clk), .A(\g.we_clk [2894]));
Q_ASSIGN U29881 ( .B(clk), .A(\g.we_clk [2893]));
Q_ASSIGN U29882 ( .B(clk), .A(\g.we_clk [2892]));
Q_ASSIGN U29883 ( .B(clk), .A(\g.we_clk [2891]));
Q_ASSIGN U29884 ( .B(clk), .A(\g.we_clk [2890]));
Q_ASSIGN U29885 ( .B(clk), .A(\g.we_clk [2889]));
Q_ASSIGN U29886 ( .B(clk), .A(\g.we_clk [2888]));
Q_ASSIGN U29887 ( .B(clk), .A(\g.we_clk [2887]));
Q_ASSIGN U29888 ( .B(clk), .A(\g.we_clk [2886]));
Q_ASSIGN U29889 ( .B(clk), .A(\g.we_clk [2885]));
Q_ASSIGN U29890 ( .B(clk), .A(\g.we_clk [2884]));
Q_ASSIGN U29891 ( .B(clk), .A(\g.we_clk [2883]));
Q_ASSIGN U29892 ( .B(clk), .A(\g.we_clk [2882]));
Q_ASSIGN U29893 ( .B(clk), .A(\g.we_clk [2881]));
Q_ASSIGN U29894 ( .B(clk), .A(\g.we_clk [2880]));
Q_ASSIGN U29895 ( .B(clk), .A(\g.we_clk [2879]));
Q_ASSIGN U29896 ( .B(clk), .A(\g.we_clk [2878]));
Q_ASSIGN U29897 ( .B(clk), .A(\g.we_clk [2877]));
Q_ASSIGN U29898 ( .B(clk), .A(\g.we_clk [2876]));
Q_ASSIGN U29899 ( .B(clk), .A(\g.we_clk [2875]));
Q_ASSIGN U29900 ( .B(clk), .A(\g.we_clk [2874]));
Q_ASSIGN U29901 ( .B(clk), .A(\g.we_clk [2873]));
Q_ASSIGN U29902 ( .B(clk), .A(\g.we_clk [2872]));
Q_ASSIGN U29903 ( .B(clk), .A(\g.we_clk [2871]));
Q_ASSIGN U29904 ( .B(clk), .A(\g.we_clk [2870]));
Q_ASSIGN U29905 ( .B(clk), .A(\g.we_clk [2869]));
Q_ASSIGN U29906 ( .B(clk), .A(\g.we_clk [2868]));
Q_ASSIGN U29907 ( .B(clk), .A(\g.we_clk [2867]));
Q_ASSIGN U29908 ( .B(clk), .A(\g.we_clk [2866]));
Q_ASSIGN U29909 ( .B(clk), .A(\g.we_clk [2865]));
Q_ASSIGN U29910 ( .B(clk), .A(\g.we_clk [2864]));
Q_ASSIGN U29911 ( .B(clk), .A(\g.we_clk [2863]));
Q_ASSIGN U29912 ( .B(clk), .A(\g.we_clk [2862]));
Q_ASSIGN U29913 ( .B(clk), .A(\g.we_clk [2861]));
Q_ASSIGN U29914 ( .B(clk), .A(\g.we_clk [2860]));
Q_ASSIGN U29915 ( .B(clk), .A(\g.we_clk [2859]));
Q_ASSIGN U29916 ( .B(clk), .A(\g.we_clk [2858]));
Q_ASSIGN U29917 ( .B(clk), .A(\g.we_clk [2857]));
Q_ASSIGN U29918 ( .B(clk), .A(\g.we_clk [2856]));
Q_ASSIGN U29919 ( .B(clk), .A(\g.we_clk [2855]));
Q_ASSIGN U29920 ( .B(clk), .A(\g.we_clk [2854]));
Q_ASSIGN U29921 ( .B(clk), .A(\g.we_clk [2853]));
Q_ASSIGN U29922 ( .B(clk), .A(\g.we_clk [2852]));
Q_ASSIGN U29923 ( .B(clk), .A(\g.we_clk [2851]));
Q_ASSIGN U29924 ( .B(clk), .A(\g.we_clk [2850]));
Q_ASSIGN U29925 ( .B(clk), .A(\g.we_clk [2849]));
Q_ASSIGN U29926 ( .B(clk), .A(\g.we_clk [2848]));
Q_ASSIGN U29927 ( .B(clk), .A(\g.we_clk [2847]));
Q_ASSIGN U29928 ( .B(clk), .A(\g.we_clk [2846]));
Q_ASSIGN U29929 ( .B(clk), .A(\g.we_clk [2845]));
Q_ASSIGN U29930 ( .B(clk), .A(\g.we_clk [2844]));
Q_ASSIGN U29931 ( .B(clk), .A(\g.we_clk [2843]));
Q_ASSIGN U29932 ( .B(clk), .A(\g.we_clk [2842]));
Q_ASSIGN U29933 ( .B(clk), .A(\g.we_clk [2841]));
Q_ASSIGN U29934 ( .B(clk), .A(\g.we_clk [2840]));
Q_ASSIGN U29935 ( .B(clk), .A(\g.we_clk [2839]));
Q_ASSIGN U29936 ( .B(clk), .A(\g.we_clk [2838]));
Q_ASSIGN U29937 ( .B(clk), .A(\g.we_clk [2837]));
Q_ASSIGN U29938 ( .B(clk), .A(\g.we_clk [2836]));
Q_ASSIGN U29939 ( .B(clk), .A(\g.we_clk [2835]));
Q_ASSIGN U29940 ( .B(clk), .A(\g.we_clk [2834]));
Q_ASSIGN U29941 ( .B(clk), .A(\g.we_clk [2833]));
Q_ASSIGN U29942 ( .B(clk), .A(\g.we_clk [2832]));
Q_ASSIGN U29943 ( .B(clk), .A(\g.we_clk [2831]));
Q_ASSIGN U29944 ( .B(clk), .A(\g.we_clk [2830]));
Q_ASSIGN U29945 ( .B(clk), .A(\g.we_clk [2829]));
Q_ASSIGN U29946 ( .B(clk), .A(\g.we_clk [2828]));
Q_ASSIGN U29947 ( .B(clk), .A(\g.we_clk [2827]));
Q_ASSIGN U29948 ( .B(clk), .A(\g.we_clk [2826]));
Q_ASSIGN U29949 ( .B(clk), .A(\g.we_clk [2825]));
Q_ASSIGN U29950 ( .B(clk), .A(\g.we_clk [2824]));
Q_ASSIGN U29951 ( .B(clk), .A(\g.we_clk [2823]));
Q_ASSIGN U29952 ( .B(clk), .A(\g.we_clk [2822]));
Q_ASSIGN U29953 ( .B(clk), .A(\g.we_clk [2821]));
Q_ASSIGN U29954 ( .B(clk), .A(\g.we_clk [2820]));
Q_ASSIGN U29955 ( .B(clk), .A(\g.we_clk [2819]));
Q_ASSIGN U29956 ( .B(clk), .A(\g.we_clk [2818]));
Q_ASSIGN U29957 ( .B(clk), .A(\g.we_clk [2817]));
Q_ASSIGN U29958 ( .B(clk), .A(\g.we_clk [2816]));
Q_ASSIGN U29959 ( .B(clk), .A(\g.we_clk [2815]));
Q_ASSIGN U29960 ( .B(clk), .A(\g.we_clk [2814]));
Q_ASSIGN U29961 ( .B(clk), .A(\g.we_clk [2813]));
Q_ASSIGN U29962 ( .B(clk), .A(\g.we_clk [2812]));
Q_ASSIGN U29963 ( .B(clk), .A(\g.we_clk [2811]));
Q_ASSIGN U29964 ( .B(clk), .A(\g.we_clk [2810]));
Q_ASSIGN U29965 ( .B(clk), .A(\g.we_clk [2809]));
Q_ASSIGN U29966 ( .B(clk), .A(\g.we_clk [2808]));
Q_ASSIGN U29967 ( .B(clk), .A(\g.we_clk [2807]));
Q_ASSIGN U29968 ( .B(clk), .A(\g.we_clk [2806]));
Q_ASSIGN U29969 ( .B(clk), .A(\g.we_clk [2805]));
Q_ASSIGN U29970 ( .B(clk), .A(\g.we_clk [2804]));
Q_ASSIGN U29971 ( .B(clk), .A(\g.we_clk [2803]));
Q_ASSIGN U29972 ( .B(clk), .A(\g.we_clk [2802]));
Q_ASSIGN U29973 ( .B(clk), .A(\g.we_clk [2801]));
Q_ASSIGN U29974 ( .B(clk), .A(\g.we_clk [2800]));
Q_ASSIGN U29975 ( .B(clk), .A(\g.we_clk [2799]));
Q_ASSIGN U29976 ( .B(clk), .A(\g.we_clk [2798]));
Q_ASSIGN U29977 ( .B(clk), .A(\g.we_clk [2797]));
Q_ASSIGN U29978 ( .B(clk), .A(\g.we_clk [2796]));
Q_ASSIGN U29979 ( .B(clk), .A(\g.we_clk [2795]));
Q_ASSIGN U29980 ( .B(clk), .A(\g.we_clk [2794]));
Q_ASSIGN U29981 ( .B(clk), .A(\g.we_clk [2793]));
Q_ASSIGN U29982 ( .B(clk), .A(\g.we_clk [2792]));
Q_ASSIGN U29983 ( .B(clk), .A(\g.we_clk [2791]));
Q_ASSIGN U29984 ( .B(clk), .A(\g.we_clk [2790]));
Q_ASSIGN U29985 ( .B(clk), .A(\g.we_clk [2789]));
Q_ASSIGN U29986 ( .B(clk), .A(\g.we_clk [2788]));
Q_ASSIGN U29987 ( .B(clk), .A(\g.we_clk [2787]));
Q_ASSIGN U29988 ( .B(clk), .A(\g.we_clk [2786]));
Q_ASSIGN U29989 ( .B(clk), .A(\g.we_clk [2785]));
Q_ASSIGN U29990 ( .B(clk), .A(\g.we_clk [2784]));
Q_ASSIGN U29991 ( .B(clk), .A(\g.we_clk [2783]));
Q_ASSIGN U29992 ( .B(clk), .A(\g.we_clk [2782]));
Q_ASSIGN U29993 ( .B(clk), .A(\g.we_clk [2781]));
Q_ASSIGN U29994 ( .B(clk), .A(\g.we_clk [2780]));
Q_ASSIGN U29995 ( .B(clk), .A(\g.we_clk [2779]));
Q_ASSIGN U29996 ( .B(clk), .A(\g.we_clk [2778]));
Q_ASSIGN U29997 ( .B(clk), .A(\g.we_clk [2777]));
Q_ASSIGN U29998 ( .B(clk), .A(\g.we_clk [2776]));
Q_ASSIGN U29999 ( .B(clk), .A(\g.we_clk [2775]));
Q_ASSIGN U30000 ( .B(clk), .A(\g.we_clk [2774]));
Q_ASSIGN U30001 ( .B(clk), .A(\g.we_clk [2773]));
Q_ASSIGN U30002 ( .B(clk), .A(\g.we_clk [2772]));
Q_ASSIGN U30003 ( .B(clk), .A(\g.we_clk [2771]));
Q_ASSIGN U30004 ( .B(clk), .A(\g.we_clk [2770]));
Q_ASSIGN U30005 ( .B(clk), .A(\g.we_clk [2769]));
Q_ASSIGN U30006 ( .B(clk), .A(\g.we_clk [2768]));
Q_ASSIGN U30007 ( .B(clk), .A(\g.we_clk [2767]));
Q_ASSIGN U30008 ( .B(clk), .A(\g.we_clk [2766]));
Q_ASSIGN U30009 ( .B(clk), .A(\g.we_clk [2765]));
Q_ASSIGN U30010 ( .B(clk), .A(\g.we_clk [2764]));
Q_ASSIGN U30011 ( .B(clk), .A(\g.we_clk [2763]));
Q_ASSIGN U30012 ( .B(clk), .A(\g.we_clk [2762]));
Q_ASSIGN U30013 ( .B(clk), .A(\g.we_clk [2761]));
Q_ASSIGN U30014 ( .B(clk), .A(\g.we_clk [2760]));
Q_ASSIGN U30015 ( .B(clk), .A(\g.we_clk [2759]));
Q_ASSIGN U30016 ( .B(clk), .A(\g.we_clk [2758]));
Q_ASSIGN U30017 ( .B(clk), .A(\g.we_clk [2757]));
Q_ASSIGN U30018 ( .B(clk), .A(\g.we_clk [2756]));
Q_ASSIGN U30019 ( .B(clk), .A(\g.we_clk [2755]));
Q_ASSIGN U30020 ( .B(clk), .A(\g.we_clk [2754]));
Q_ASSIGN U30021 ( .B(clk), .A(\g.we_clk [2753]));
Q_ASSIGN U30022 ( .B(clk), .A(\g.we_clk [2752]));
Q_ASSIGN U30023 ( .B(clk), .A(\g.we_clk [2751]));
Q_ASSIGN U30024 ( .B(clk), .A(\g.we_clk [2750]));
Q_ASSIGN U30025 ( .B(clk), .A(\g.we_clk [2749]));
Q_ASSIGN U30026 ( .B(clk), .A(\g.we_clk [2748]));
Q_ASSIGN U30027 ( .B(clk), .A(\g.we_clk [2747]));
Q_ASSIGN U30028 ( .B(clk), .A(\g.we_clk [2746]));
Q_ASSIGN U30029 ( .B(clk), .A(\g.we_clk [2745]));
Q_ASSIGN U30030 ( .B(clk), .A(\g.we_clk [2744]));
Q_ASSIGN U30031 ( .B(clk), .A(\g.we_clk [2743]));
Q_ASSIGN U30032 ( .B(clk), .A(\g.we_clk [2742]));
Q_ASSIGN U30033 ( .B(clk), .A(\g.we_clk [2741]));
Q_ASSIGN U30034 ( .B(clk), .A(\g.we_clk [2740]));
Q_ASSIGN U30035 ( .B(clk), .A(\g.we_clk [2739]));
Q_ASSIGN U30036 ( .B(clk), .A(\g.we_clk [2738]));
Q_ASSIGN U30037 ( .B(clk), .A(\g.we_clk [2737]));
Q_ASSIGN U30038 ( .B(clk), .A(\g.we_clk [2736]));
Q_ASSIGN U30039 ( .B(clk), .A(\g.we_clk [2735]));
Q_ASSIGN U30040 ( .B(clk), .A(\g.we_clk [2734]));
Q_ASSIGN U30041 ( .B(clk), .A(\g.we_clk [2733]));
Q_ASSIGN U30042 ( .B(clk), .A(\g.we_clk [2732]));
Q_ASSIGN U30043 ( .B(clk), .A(\g.we_clk [2731]));
Q_ASSIGN U30044 ( .B(clk), .A(\g.we_clk [2730]));
Q_ASSIGN U30045 ( .B(clk), .A(\g.we_clk [2729]));
Q_ASSIGN U30046 ( .B(clk), .A(\g.we_clk [2728]));
Q_ASSIGN U30047 ( .B(clk), .A(\g.we_clk [2727]));
Q_ASSIGN U30048 ( .B(clk), .A(\g.we_clk [2726]));
Q_ASSIGN U30049 ( .B(clk), .A(\g.we_clk [2725]));
Q_ASSIGN U30050 ( .B(clk), .A(\g.we_clk [2724]));
Q_ASSIGN U30051 ( .B(clk), .A(\g.we_clk [2723]));
Q_ASSIGN U30052 ( .B(clk), .A(\g.we_clk [2722]));
Q_ASSIGN U30053 ( .B(clk), .A(\g.we_clk [2721]));
Q_ASSIGN U30054 ( .B(clk), .A(\g.we_clk [2720]));
Q_ASSIGN U30055 ( .B(clk), .A(\g.we_clk [2719]));
Q_ASSIGN U30056 ( .B(clk), .A(\g.we_clk [2718]));
Q_ASSIGN U30057 ( .B(clk), .A(\g.we_clk [2717]));
Q_ASSIGN U30058 ( .B(clk), .A(\g.we_clk [2716]));
Q_ASSIGN U30059 ( .B(clk), .A(\g.we_clk [2715]));
Q_ASSIGN U30060 ( .B(clk), .A(\g.we_clk [2714]));
Q_ASSIGN U30061 ( .B(clk), .A(\g.we_clk [2713]));
Q_ASSIGN U30062 ( .B(clk), .A(\g.we_clk [2712]));
Q_ASSIGN U30063 ( .B(clk), .A(\g.we_clk [2711]));
Q_ASSIGN U30064 ( .B(clk), .A(\g.we_clk [2710]));
Q_ASSIGN U30065 ( .B(clk), .A(\g.we_clk [2709]));
Q_ASSIGN U30066 ( .B(clk), .A(\g.we_clk [2708]));
Q_ASSIGN U30067 ( .B(clk), .A(\g.we_clk [2707]));
Q_ASSIGN U30068 ( .B(clk), .A(\g.we_clk [2706]));
Q_ASSIGN U30069 ( .B(clk), .A(\g.we_clk [2705]));
Q_ASSIGN U30070 ( .B(clk), .A(\g.we_clk [2704]));
Q_ASSIGN U30071 ( .B(clk), .A(\g.we_clk [2703]));
Q_ASSIGN U30072 ( .B(clk), .A(\g.we_clk [2702]));
Q_ASSIGN U30073 ( .B(clk), .A(\g.we_clk [2701]));
Q_ASSIGN U30074 ( .B(clk), .A(\g.we_clk [2700]));
Q_ASSIGN U30075 ( .B(clk), .A(\g.we_clk [2699]));
Q_ASSIGN U30076 ( .B(clk), .A(\g.we_clk [2698]));
Q_ASSIGN U30077 ( .B(clk), .A(\g.we_clk [2697]));
Q_ASSIGN U30078 ( .B(clk), .A(\g.we_clk [2696]));
Q_ASSIGN U30079 ( .B(clk), .A(\g.we_clk [2695]));
Q_ASSIGN U30080 ( .B(clk), .A(\g.we_clk [2694]));
Q_ASSIGN U30081 ( .B(clk), .A(\g.we_clk [2693]));
Q_ASSIGN U30082 ( .B(clk), .A(\g.we_clk [2692]));
Q_ASSIGN U30083 ( .B(clk), .A(\g.we_clk [2691]));
Q_ASSIGN U30084 ( .B(clk), .A(\g.we_clk [2690]));
Q_ASSIGN U30085 ( .B(clk), .A(\g.we_clk [2689]));
Q_ASSIGN U30086 ( .B(clk), .A(\g.we_clk [2688]));
Q_ASSIGN U30087 ( .B(clk), .A(\g.we_clk [2687]));
Q_ASSIGN U30088 ( .B(clk), .A(\g.we_clk [2686]));
Q_ASSIGN U30089 ( .B(clk), .A(\g.we_clk [2685]));
Q_ASSIGN U30090 ( .B(clk), .A(\g.we_clk [2684]));
Q_ASSIGN U30091 ( .B(clk), .A(\g.we_clk [2683]));
Q_ASSIGN U30092 ( .B(clk), .A(\g.we_clk [2682]));
Q_ASSIGN U30093 ( .B(clk), .A(\g.we_clk [2681]));
Q_ASSIGN U30094 ( .B(clk), .A(\g.we_clk [2680]));
Q_ASSIGN U30095 ( .B(clk), .A(\g.we_clk [2679]));
Q_ASSIGN U30096 ( .B(clk), .A(\g.we_clk [2678]));
Q_ASSIGN U30097 ( .B(clk), .A(\g.we_clk [2677]));
Q_ASSIGN U30098 ( .B(clk), .A(\g.we_clk [2676]));
Q_ASSIGN U30099 ( .B(clk), .A(\g.we_clk [2675]));
Q_ASSIGN U30100 ( .B(clk), .A(\g.we_clk [2674]));
Q_ASSIGN U30101 ( .B(clk), .A(\g.we_clk [2673]));
Q_ASSIGN U30102 ( .B(clk), .A(\g.we_clk [2672]));
Q_ASSIGN U30103 ( .B(clk), .A(\g.we_clk [2671]));
Q_ASSIGN U30104 ( .B(clk), .A(\g.we_clk [2670]));
Q_ASSIGN U30105 ( .B(clk), .A(\g.we_clk [2669]));
Q_ASSIGN U30106 ( .B(clk), .A(\g.we_clk [2668]));
Q_ASSIGN U30107 ( .B(clk), .A(\g.we_clk [2667]));
Q_ASSIGN U30108 ( .B(clk), .A(\g.we_clk [2666]));
Q_ASSIGN U30109 ( .B(clk), .A(\g.we_clk [2665]));
Q_ASSIGN U30110 ( .B(clk), .A(\g.we_clk [2664]));
Q_ASSIGN U30111 ( .B(clk), .A(\g.we_clk [2663]));
Q_ASSIGN U30112 ( .B(clk), .A(\g.we_clk [2662]));
Q_ASSIGN U30113 ( .B(clk), .A(\g.we_clk [2661]));
Q_ASSIGN U30114 ( .B(clk), .A(\g.we_clk [2660]));
Q_ASSIGN U30115 ( .B(clk), .A(\g.we_clk [2659]));
Q_ASSIGN U30116 ( .B(clk), .A(\g.we_clk [2658]));
Q_ASSIGN U30117 ( .B(clk), .A(\g.we_clk [2657]));
Q_ASSIGN U30118 ( .B(clk), .A(\g.we_clk [2656]));
Q_ASSIGN U30119 ( .B(clk), .A(\g.we_clk [2655]));
Q_ASSIGN U30120 ( .B(clk), .A(\g.we_clk [2654]));
Q_ASSIGN U30121 ( .B(clk), .A(\g.we_clk [2653]));
Q_ASSIGN U30122 ( .B(clk), .A(\g.we_clk [2652]));
Q_ASSIGN U30123 ( .B(clk), .A(\g.we_clk [2651]));
Q_ASSIGN U30124 ( .B(clk), .A(\g.we_clk [2650]));
Q_ASSIGN U30125 ( .B(clk), .A(\g.we_clk [2649]));
Q_ASSIGN U30126 ( .B(clk), .A(\g.we_clk [2648]));
Q_ASSIGN U30127 ( .B(clk), .A(\g.we_clk [2647]));
Q_ASSIGN U30128 ( .B(clk), .A(\g.we_clk [2646]));
Q_ASSIGN U30129 ( .B(clk), .A(\g.we_clk [2645]));
Q_ASSIGN U30130 ( .B(clk), .A(\g.we_clk [2644]));
Q_ASSIGN U30131 ( .B(clk), .A(\g.we_clk [2643]));
Q_ASSIGN U30132 ( .B(clk), .A(\g.we_clk [2642]));
Q_ASSIGN U30133 ( .B(clk), .A(\g.we_clk [2641]));
Q_ASSIGN U30134 ( .B(clk), .A(\g.we_clk [2640]));
Q_ASSIGN U30135 ( .B(clk), .A(\g.we_clk [2639]));
Q_ASSIGN U30136 ( .B(clk), .A(\g.we_clk [2638]));
Q_ASSIGN U30137 ( .B(clk), .A(\g.we_clk [2637]));
Q_ASSIGN U30138 ( .B(clk), .A(\g.we_clk [2636]));
Q_ASSIGN U30139 ( .B(clk), .A(\g.we_clk [2635]));
Q_ASSIGN U30140 ( .B(clk), .A(\g.we_clk [2634]));
Q_ASSIGN U30141 ( .B(clk), .A(\g.we_clk [2633]));
Q_ASSIGN U30142 ( .B(clk), .A(\g.we_clk [2632]));
Q_ASSIGN U30143 ( .B(clk), .A(\g.we_clk [2631]));
Q_ASSIGN U30144 ( .B(clk), .A(\g.we_clk [2630]));
Q_ASSIGN U30145 ( .B(clk), .A(\g.we_clk [2629]));
Q_ASSIGN U30146 ( .B(clk), .A(\g.we_clk [2628]));
Q_ASSIGN U30147 ( .B(clk), .A(\g.we_clk [2627]));
Q_ASSIGN U30148 ( .B(clk), .A(\g.we_clk [2626]));
Q_ASSIGN U30149 ( .B(clk), .A(\g.we_clk [2625]));
Q_ASSIGN U30150 ( .B(clk), .A(\g.we_clk [2624]));
Q_ASSIGN U30151 ( .B(clk), .A(\g.we_clk [2623]));
Q_ASSIGN U30152 ( .B(clk), .A(\g.we_clk [2622]));
Q_ASSIGN U30153 ( .B(clk), .A(\g.we_clk [2621]));
Q_ASSIGN U30154 ( .B(clk), .A(\g.we_clk [2620]));
Q_ASSIGN U30155 ( .B(clk), .A(\g.we_clk [2619]));
Q_ASSIGN U30156 ( .B(clk), .A(\g.we_clk [2618]));
Q_ASSIGN U30157 ( .B(clk), .A(\g.we_clk [2617]));
Q_ASSIGN U30158 ( .B(clk), .A(\g.we_clk [2616]));
Q_ASSIGN U30159 ( .B(clk), .A(\g.we_clk [2615]));
Q_ASSIGN U30160 ( .B(clk), .A(\g.we_clk [2614]));
Q_ASSIGN U30161 ( .B(clk), .A(\g.we_clk [2613]));
Q_ASSIGN U30162 ( .B(clk), .A(\g.we_clk [2612]));
Q_ASSIGN U30163 ( .B(clk), .A(\g.we_clk [2611]));
Q_ASSIGN U30164 ( .B(clk), .A(\g.we_clk [2610]));
Q_ASSIGN U30165 ( .B(clk), .A(\g.we_clk [2609]));
Q_ASSIGN U30166 ( .B(clk), .A(\g.we_clk [2608]));
Q_ASSIGN U30167 ( .B(clk), .A(\g.we_clk [2607]));
Q_ASSIGN U30168 ( .B(clk), .A(\g.we_clk [2606]));
Q_ASSIGN U30169 ( .B(clk), .A(\g.we_clk [2605]));
Q_ASSIGN U30170 ( .B(clk), .A(\g.we_clk [2604]));
Q_ASSIGN U30171 ( .B(clk), .A(\g.we_clk [2603]));
Q_ASSIGN U30172 ( .B(clk), .A(\g.we_clk [2602]));
Q_ASSIGN U30173 ( .B(clk), .A(\g.we_clk [2601]));
Q_ASSIGN U30174 ( .B(clk), .A(\g.we_clk [2600]));
Q_ASSIGN U30175 ( .B(clk), .A(\g.we_clk [2599]));
Q_ASSIGN U30176 ( .B(clk), .A(\g.we_clk [2598]));
Q_ASSIGN U30177 ( .B(clk), .A(\g.we_clk [2597]));
Q_ASSIGN U30178 ( .B(clk), .A(\g.we_clk [2596]));
Q_ASSIGN U30179 ( .B(clk), .A(\g.we_clk [2595]));
Q_ASSIGN U30180 ( .B(clk), .A(\g.we_clk [2594]));
Q_ASSIGN U30181 ( .B(clk), .A(\g.we_clk [2593]));
Q_ASSIGN U30182 ( .B(clk), .A(\g.we_clk [2592]));
Q_ASSIGN U30183 ( .B(clk), .A(\g.we_clk [2591]));
Q_ASSIGN U30184 ( .B(clk), .A(\g.we_clk [2590]));
Q_ASSIGN U30185 ( .B(clk), .A(\g.we_clk [2589]));
Q_ASSIGN U30186 ( .B(clk), .A(\g.we_clk [2588]));
Q_ASSIGN U30187 ( .B(clk), .A(\g.we_clk [2587]));
Q_ASSIGN U30188 ( .B(clk), .A(\g.we_clk [2586]));
Q_ASSIGN U30189 ( .B(clk), .A(\g.we_clk [2585]));
Q_ASSIGN U30190 ( .B(clk), .A(\g.we_clk [2584]));
Q_ASSIGN U30191 ( .B(clk), .A(\g.we_clk [2583]));
Q_ASSIGN U30192 ( .B(clk), .A(\g.we_clk [2582]));
Q_ASSIGN U30193 ( .B(clk), .A(\g.we_clk [2581]));
Q_ASSIGN U30194 ( .B(clk), .A(\g.we_clk [2580]));
Q_ASSIGN U30195 ( .B(clk), .A(\g.we_clk [2579]));
Q_ASSIGN U30196 ( .B(clk), .A(\g.we_clk [2578]));
Q_ASSIGN U30197 ( .B(clk), .A(\g.we_clk [2577]));
Q_ASSIGN U30198 ( .B(clk), .A(\g.we_clk [2576]));
Q_ASSIGN U30199 ( .B(clk), .A(\g.we_clk [2575]));
Q_ASSIGN U30200 ( .B(clk), .A(\g.we_clk [2574]));
Q_ASSIGN U30201 ( .B(clk), .A(\g.we_clk [2573]));
Q_ASSIGN U30202 ( .B(clk), .A(\g.we_clk [2572]));
Q_ASSIGN U30203 ( .B(clk), .A(\g.we_clk [2571]));
Q_ASSIGN U30204 ( .B(clk), .A(\g.we_clk [2570]));
Q_ASSIGN U30205 ( .B(clk), .A(\g.we_clk [2569]));
Q_ASSIGN U30206 ( .B(clk), .A(\g.we_clk [2568]));
Q_ASSIGN U30207 ( .B(clk), .A(\g.we_clk [2567]));
Q_ASSIGN U30208 ( .B(clk), .A(\g.we_clk [2566]));
Q_ASSIGN U30209 ( .B(clk), .A(\g.we_clk [2565]));
Q_ASSIGN U30210 ( .B(clk), .A(\g.we_clk [2564]));
Q_ASSIGN U30211 ( .B(clk), .A(\g.we_clk [2563]));
Q_ASSIGN U30212 ( .B(clk), .A(\g.we_clk [2562]));
Q_ASSIGN U30213 ( .B(clk), .A(\g.we_clk [2561]));
Q_ASSIGN U30214 ( .B(clk), .A(\g.we_clk [2560]));
Q_ASSIGN U30215 ( .B(clk), .A(\g.we_clk [2559]));
Q_ASSIGN U30216 ( .B(clk), .A(\g.we_clk [2558]));
Q_ASSIGN U30217 ( .B(clk), .A(\g.we_clk [2557]));
Q_ASSIGN U30218 ( .B(clk), .A(\g.we_clk [2556]));
Q_ASSIGN U30219 ( .B(clk), .A(\g.we_clk [2555]));
Q_ASSIGN U30220 ( .B(clk), .A(\g.we_clk [2554]));
Q_ASSIGN U30221 ( .B(clk), .A(\g.we_clk [2553]));
Q_ASSIGN U30222 ( .B(clk), .A(\g.we_clk [2552]));
Q_ASSIGN U30223 ( .B(clk), .A(\g.we_clk [2551]));
Q_ASSIGN U30224 ( .B(clk), .A(\g.we_clk [2550]));
Q_ASSIGN U30225 ( .B(clk), .A(\g.we_clk [2549]));
Q_ASSIGN U30226 ( .B(clk), .A(\g.we_clk [2548]));
Q_ASSIGN U30227 ( .B(clk), .A(\g.we_clk [2547]));
Q_ASSIGN U30228 ( .B(clk), .A(\g.we_clk [2546]));
Q_ASSIGN U30229 ( .B(clk), .A(\g.we_clk [2545]));
Q_ASSIGN U30230 ( .B(clk), .A(\g.we_clk [2544]));
Q_ASSIGN U30231 ( .B(clk), .A(\g.we_clk [2543]));
Q_ASSIGN U30232 ( .B(clk), .A(\g.we_clk [2542]));
Q_ASSIGN U30233 ( .B(clk), .A(\g.we_clk [2541]));
Q_ASSIGN U30234 ( .B(clk), .A(\g.we_clk [2540]));
Q_ASSIGN U30235 ( .B(clk), .A(\g.we_clk [2539]));
Q_ASSIGN U30236 ( .B(clk), .A(\g.we_clk [2538]));
Q_ASSIGN U30237 ( .B(clk), .A(\g.we_clk [2537]));
Q_ASSIGN U30238 ( .B(clk), .A(\g.we_clk [2536]));
Q_ASSIGN U30239 ( .B(clk), .A(\g.we_clk [2535]));
Q_ASSIGN U30240 ( .B(clk), .A(\g.we_clk [2534]));
Q_ASSIGN U30241 ( .B(clk), .A(\g.we_clk [2533]));
Q_ASSIGN U30242 ( .B(clk), .A(\g.we_clk [2532]));
Q_ASSIGN U30243 ( .B(clk), .A(\g.we_clk [2531]));
Q_ASSIGN U30244 ( .B(clk), .A(\g.we_clk [2530]));
Q_ASSIGN U30245 ( .B(clk), .A(\g.we_clk [2529]));
Q_ASSIGN U30246 ( .B(clk), .A(\g.we_clk [2528]));
Q_ASSIGN U30247 ( .B(clk), .A(\g.we_clk [2527]));
Q_ASSIGN U30248 ( .B(clk), .A(\g.we_clk [2526]));
Q_ASSIGN U30249 ( .B(clk), .A(\g.we_clk [2525]));
Q_ASSIGN U30250 ( .B(clk), .A(\g.we_clk [2524]));
Q_ASSIGN U30251 ( .B(clk), .A(\g.we_clk [2523]));
Q_ASSIGN U30252 ( .B(clk), .A(\g.we_clk [2522]));
Q_ASSIGN U30253 ( .B(clk), .A(\g.we_clk [2521]));
Q_ASSIGN U30254 ( .B(clk), .A(\g.we_clk [2520]));
Q_ASSIGN U30255 ( .B(clk), .A(\g.we_clk [2519]));
Q_ASSIGN U30256 ( .B(clk), .A(\g.we_clk [2518]));
Q_ASSIGN U30257 ( .B(clk), .A(\g.we_clk [2517]));
Q_ASSIGN U30258 ( .B(clk), .A(\g.we_clk [2516]));
Q_ASSIGN U30259 ( .B(clk), .A(\g.we_clk [2515]));
Q_ASSIGN U30260 ( .B(clk), .A(\g.we_clk [2514]));
Q_ASSIGN U30261 ( .B(clk), .A(\g.we_clk [2513]));
Q_ASSIGN U30262 ( .B(clk), .A(\g.we_clk [2512]));
Q_ASSIGN U30263 ( .B(clk), .A(\g.we_clk [2511]));
Q_ASSIGN U30264 ( .B(clk), .A(\g.we_clk [2510]));
Q_ASSIGN U30265 ( .B(clk), .A(\g.we_clk [2509]));
Q_ASSIGN U30266 ( .B(clk), .A(\g.we_clk [2508]));
Q_ASSIGN U30267 ( .B(clk), .A(\g.we_clk [2507]));
Q_ASSIGN U30268 ( .B(clk), .A(\g.we_clk [2506]));
Q_ASSIGN U30269 ( .B(clk), .A(\g.we_clk [2505]));
Q_ASSIGN U30270 ( .B(clk), .A(\g.we_clk [2504]));
Q_ASSIGN U30271 ( .B(clk), .A(\g.we_clk [2503]));
Q_ASSIGN U30272 ( .B(clk), .A(\g.we_clk [2502]));
Q_ASSIGN U30273 ( .B(clk), .A(\g.we_clk [2501]));
Q_ASSIGN U30274 ( .B(clk), .A(\g.we_clk [2500]));
Q_ASSIGN U30275 ( .B(clk), .A(\g.we_clk [2499]));
Q_ASSIGN U30276 ( .B(clk), .A(\g.we_clk [2498]));
Q_ASSIGN U30277 ( .B(clk), .A(\g.we_clk [2497]));
Q_ASSIGN U30278 ( .B(clk), .A(\g.we_clk [2496]));
Q_ASSIGN U30279 ( .B(clk), .A(\g.we_clk [2495]));
Q_ASSIGN U30280 ( .B(clk), .A(\g.we_clk [2494]));
Q_ASSIGN U30281 ( .B(clk), .A(\g.we_clk [2493]));
Q_ASSIGN U30282 ( .B(clk), .A(\g.we_clk [2492]));
Q_ASSIGN U30283 ( .B(clk), .A(\g.we_clk [2491]));
Q_ASSIGN U30284 ( .B(clk), .A(\g.we_clk [2490]));
Q_ASSIGN U30285 ( .B(clk), .A(\g.we_clk [2489]));
Q_ASSIGN U30286 ( .B(clk), .A(\g.we_clk [2488]));
Q_ASSIGN U30287 ( .B(clk), .A(\g.we_clk [2487]));
Q_ASSIGN U30288 ( .B(clk), .A(\g.we_clk [2486]));
Q_ASSIGN U30289 ( .B(clk), .A(\g.we_clk [2485]));
Q_ASSIGN U30290 ( .B(clk), .A(\g.we_clk [2484]));
Q_ASSIGN U30291 ( .B(clk), .A(\g.we_clk [2483]));
Q_ASSIGN U30292 ( .B(clk), .A(\g.we_clk [2482]));
Q_ASSIGN U30293 ( .B(clk), .A(\g.we_clk [2481]));
Q_ASSIGN U30294 ( .B(clk), .A(\g.we_clk [2480]));
Q_ASSIGN U30295 ( .B(clk), .A(\g.we_clk [2479]));
Q_ASSIGN U30296 ( .B(clk), .A(\g.we_clk [2478]));
Q_ASSIGN U30297 ( .B(clk), .A(\g.we_clk [2477]));
Q_ASSIGN U30298 ( .B(clk), .A(\g.we_clk [2476]));
Q_ASSIGN U30299 ( .B(clk), .A(\g.we_clk [2475]));
Q_ASSIGN U30300 ( .B(clk), .A(\g.we_clk [2474]));
Q_ASSIGN U30301 ( .B(clk), .A(\g.we_clk [2473]));
Q_ASSIGN U30302 ( .B(clk), .A(\g.we_clk [2472]));
Q_ASSIGN U30303 ( .B(clk), .A(\g.we_clk [2471]));
Q_ASSIGN U30304 ( .B(clk), .A(\g.we_clk [2470]));
Q_ASSIGN U30305 ( .B(clk), .A(\g.we_clk [2469]));
Q_ASSIGN U30306 ( .B(clk), .A(\g.we_clk [2468]));
Q_ASSIGN U30307 ( .B(clk), .A(\g.we_clk [2467]));
Q_ASSIGN U30308 ( .B(clk), .A(\g.we_clk [2466]));
Q_ASSIGN U30309 ( .B(clk), .A(\g.we_clk [2465]));
Q_ASSIGN U30310 ( .B(clk), .A(\g.we_clk [2464]));
Q_ASSIGN U30311 ( .B(clk), .A(\g.we_clk [2463]));
Q_ASSIGN U30312 ( .B(clk), .A(\g.we_clk [2462]));
Q_ASSIGN U30313 ( .B(clk), .A(\g.we_clk [2461]));
Q_ASSIGN U30314 ( .B(clk), .A(\g.we_clk [2460]));
Q_ASSIGN U30315 ( .B(clk), .A(\g.we_clk [2459]));
Q_ASSIGN U30316 ( .B(clk), .A(\g.we_clk [2458]));
Q_ASSIGN U30317 ( .B(clk), .A(\g.we_clk [2457]));
Q_ASSIGN U30318 ( .B(clk), .A(\g.we_clk [2456]));
Q_ASSIGN U30319 ( .B(clk), .A(\g.we_clk [2455]));
Q_ASSIGN U30320 ( .B(clk), .A(\g.we_clk [2454]));
Q_ASSIGN U30321 ( .B(clk), .A(\g.we_clk [2453]));
Q_ASSIGN U30322 ( .B(clk), .A(\g.we_clk [2452]));
Q_ASSIGN U30323 ( .B(clk), .A(\g.we_clk [2451]));
Q_ASSIGN U30324 ( .B(clk), .A(\g.we_clk [2450]));
Q_ASSIGN U30325 ( .B(clk), .A(\g.we_clk [2449]));
Q_ASSIGN U30326 ( .B(clk), .A(\g.we_clk [2448]));
Q_ASSIGN U30327 ( .B(clk), .A(\g.we_clk [2447]));
Q_ASSIGN U30328 ( .B(clk), .A(\g.we_clk [2446]));
Q_ASSIGN U30329 ( .B(clk), .A(\g.we_clk [2445]));
Q_ASSIGN U30330 ( .B(clk), .A(\g.we_clk [2444]));
Q_ASSIGN U30331 ( .B(clk), .A(\g.we_clk [2443]));
Q_ASSIGN U30332 ( .B(clk), .A(\g.we_clk [2442]));
Q_ASSIGN U30333 ( .B(clk), .A(\g.we_clk [2441]));
Q_ASSIGN U30334 ( .B(clk), .A(\g.we_clk [2440]));
Q_ASSIGN U30335 ( .B(clk), .A(\g.we_clk [2439]));
Q_ASSIGN U30336 ( .B(clk), .A(\g.we_clk [2438]));
Q_ASSIGN U30337 ( .B(clk), .A(\g.we_clk [2437]));
Q_ASSIGN U30338 ( .B(clk), .A(\g.we_clk [2436]));
Q_ASSIGN U30339 ( .B(clk), .A(\g.we_clk [2435]));
Q_ASSIGN U30340 ( .B(clk), .A(\g.we_clk [2434]));
Q_ASSIGN U30341 ( .B(clk), .A(\g.we_clk [2433]));
Q_ASSIGN U30342 ( .B(clk), .A(\g.we_clk [2432]));
Q_ASSIGN U30343 ( .B(clk), .A(\g.we_clk [2431]));
Q_ASSIGN U30344 ( .B(clk), .A(\g.we_clk [2430]));
Q_ASSIGN U30345 ( .B(clk), .A(\g.we_clk [2429]));
Q_ASSIGN U30346 ( .B(clk), .A(\g.we_clk [2428]));
Q_ASSIGN U30347 ( .B(clk), .A(\g.we_clk [2427]));
Q_ASSIGN U30348 ( .B(clk), .A(\g.we_clk [2426]));
Q_ASSIGN U30349 ( .B(clk), .A(\g.we_clk [2425]));
Q_ASSIGN U30350 ( .B(clk), .A(\g.we_clk [2424]));
Q_ASSIGN U30351 ( .B(clk), .A(\g.we_clk [2423]));
Q_ASSIGN U30352 ( .B(clk), .A(\g.we_clk [2422]));
Q_ASSIGN U30353 ( .B(clk), .A(\g.we_clk [2421]));
Q_ASSIGN U30354 ( .B(clk), .A(\g.we_clk [2420]));
Q_ASSIGN U30355 ( .B(clk), .A(\g.we_clk [2419]));
Q_ASSIGN U30356 ( .B(clk), .A(\g.we_clk [2418]));
Q_ASSIGN U30357 ( .B(clk), .A(\g.we_clk [2417]));
Q_ASSIGN U30358 ( .B(clk), .A(\g.we_clk [2416]));
Q_ASSIGN U30359 ( .B(clk), .A(\g.we_clk [2415]));
Q_ASSIGN U30360 ( .B(clk), .A(\g.we_clk [2414]));
Q_ASSIGN U30361 ( .B(clk), .A(\g.we_clk [2413]));
Q_ASSIGN U30362 ( .B(clk), .A(\g.we_clk [2412]));
Q_ASSIGN U30363 ( .B(clk), .A(\g.we_clk [2411]));
Q_ASSIGN U30364 ( .B(clk), .A(\g.we_clk [2410]));
Q_ASSIGN U30365 ( .B(clk), .A(\g.we_clk [2409]));
Q_ASSIGN U30366 ( .B(clk), .A(\g.we_clk [2408]));
Q_ASSIGN U30367 ( .B(clk), .A(\g.we_clk [2407]));
Q_ASSIGN U30368 ( .B(clk), .A(\g.we_clk [2406]));
Q_ASSIGN U30369 ( .B(clk), .A(\g.we_clk [2405]));
Q_ASSIGN U30370 ( .B(clk), .A(\g.we_clk [2404]));
Q_ASSIGN U30371 ( .B(clk), .A(\g.we_clk [2403]));
Q_ASSIGN U30372 ( .B(clk), .A(\g.we_clk [2402]));
Q_ASSIGN U30373 ( .B(clk), .A(\g.we_clk [2401]));
Q_ASSIGN U30374 ( .B(clk), .A(\g.we_clk [2400]));
Q_ASSIGN U30375 ( .B(clk), .A(\g.we_clk [2399]));
Q_ASSIGN U30376 ( .B(clk), .A(\g.we_clk [2398]));
Q_ASSIGN U30377 ( .B(clk), .A(\g.we_clk [2397]));
Q_ASSIGN U30378 ( .B(clk), .A(\g.we_clk [2396]));
Q_ASSIGN U30379 ( .B(clk), .A(\g.we_clk [2395]));
Q_ASSIGN U30380 ( .B(clk), .A(\g.we_clk [2394]));
Q_ASSIGN U30381 ( .B(clk), .A(\g.we_clk [2393]));
Q_ASSIGN U30382 ( .B(clk), .A(\g.we_clk [2392]));
Q_ASSIGN U30383 ( .B(clk), .A(\g.we_clk [2391]));
Q_ASSIGN U30384 ( .B(clk), .A(\g.we_clk [2390]));
Q_ASSIGN U30385 ( .B(clk), .A(\g.we_clk [2389]));
Q_ASSIGN U30386 ( .B(clk), .A(\g.we_clk [2388]));
Q_ASSIGN U30387 ( .B(clk), .A(\g.we_clk [2387]));
Q_ASSIGN U30388 ( .B(clk), .A(\g.we_clk [2386]));
Q_ASSIGN U30389 ( .B(clk), .A(\g.we_clk [2385]));
Q_ASSIGN U30390 ( .B(clk), .A(\g.we_clk [2384]));
Q_ASSIGN U30391 ( .B(clk), .A(\g.we_clk [2383]));
Q_ASSIGN U30392 ( .B(clk), .A(\g.we_clk [2382]));
Q_ASSIGN U30393 ( .B(clk), .A(\g.we_clk [2381]));
Q_ASSIGN U30394 ( .B(clk), .A(\g.we_clk [2380]));
Q_ASSIGN U30395 ( .B(clk), .A(\g.we_clk [2379]));
Q_ASSIGN U30396 ( .B(clk), .A(\g.we_clk [2378]));
Q_ASSIGN U30397 ( .B(clk), .A(\g.we_clk [2377]));
Q_ASSIGN U30398 ( .B(clk), .A(\g.we_clk [2376]));
Q_ASSIGN U30399 ( .B(clk), .A(\g.we_clk [2375]));
Q_ASSIGN U30400 ( .B(clk), .A(\g.we_clk [2374]));
Q_ASSIGN U30401 ( .B(clk), .A(\g.we_clk [2373]));
Q_ASSIGN U30402 ( .B(clk), .A(\g.we_clk [2372]));
Q_ASSIGN U30403 ( .B(clk), .A(\g.we_clk [2371]));
Q_ASSIGN U30404 ( .B(clk), .A(\g.we_clk [2370]));
Q_ASSIGN U30405 ( .B(clk), .A(\g.we_clk [2369]));
Q_ASSIGN U30406 ( .B(clk), .A(\g.we_clk [2368]));
Q_ASSIGN U30407 ( .B(clk), .A(\g.we_clk [2367]));
Q_ASSIGN U30408 ( .B(clk), .A(\g.we_clk [2366]));
Q_ASSIGN U30409 ( .B(clk), .A(\g.we_clk [2365]));
Q_ASSIGN U30410 ( .B(clk), .A(\g.we_clk [2364]));
Q_ASSIGN U30411 ( .B(clk), .A(\g.we_clk [2363]));
Q_ASSIGN U30412 ( .B(clk), .A(\g.we_clk [2362]));
Q_ASSIGN U30413 ( .B(clk), .A(\g.we_clk [2361]));
Q_ASSIGN U30414 ( .B(clk), .A(\g.we_clk [2360]));
Q_ASSIGN U30415 ( .B(clk), .A(\g.we_clk [2359]));
Q_ASSIGN U30416 ( .B(clk), .A(\g.we_clk [2358]));
Q_ASSIGN U30417 ( .B(clk), .A(\g.we_clk [2357]));
Q_ASSIGN U30418 ( .B(clk), .A(\g.we_clk [2356]));
Q_ASSIGN U30419 ( .B(clk), .A(\g.we_clk [2355]));
Q_ASSIGN U30420 ( .B(clk), .A(\g.we_clk [2354]));
Q_ASSIGN U30421 ( .B(clk), .A(\g.we_clk [2353]));
Q_ASSIGN U30422 ( .B(clk), .A(\g.we_clk [2352]));
Q_ASSIGN U30423 ( .B(clk), .A(\g.we_clk [2351]));
Q_ASSIGN U30424 ( .B(clk), .A(\g.we_clk [2350]));
Q_ASSIGN U30425 ( .B(clk), .A(\g.we_clk [2349]));
Q_ASSIGN U30426 ( .B(clk), .A(\g.we_clk [2348]));
Q_ASSIGN U30427 ( .B(clk), .A(\g.we_clk [2347]));
Q_ASSIGN U30428 ( .B(clk), .A(\g.we_clk [2346]));
Q_ASSIGN U30429 ( .B(clk), .A(\g.we_clk [2345]));
Q_ASSIGN U30430 ( .B(clk), .A(\g.we_clk [2344]));
Q_ASSIGN U30431 ( .B(clk), .A(\g.we_clk [2343]));
Q_ASSIGN U30432 ( .B(clk), .A(\g.we_clk [2342]));
Q_ASSIGN U30433 ( .B(clk), .A(\g.we_clk [2341]));
Q_ASSIGN U30434 ( .B(clk), .A(\g.we_clk [2340]));
Q_ASSIGN U30435 ( .B(clk), .A(\g.we_clk [2339]));
Q_ASSIGN U30436 ( .B(clk), .A(\g.we_clk [2338]));
Q_ASSIGN U30437 ( .B(clk), .A(\g.we_clk [2337]));
Q_ASSIGN U30438 ( .B(clk), .A(\g.we_clk [2336]));
Q_ASSIGN U30439 ( .B(clk), .A(\g.we_clk [2335]));
Q_ASSIGN U30440 ( .B(clk), .A(\g.we_clk [2334]));
Q_ASSIGN U30441 ( .B(clk), .A(\g.we_clk [2333]));
Q_ASSIGN U30442 ( .B(clk), .A(\g.we_clk [2332]));
Q_ASSIGN U30443 ( .B(clk), .A(\g.we_clk [2331]));
Q_ASSIGN U30444 ( .B(clk), .A(\g.we_clk [2330]));
Q_ASSIGN U30445 ( .B(clk), .A(\g.we_clk [2329]));
Q_ASSIGN U30446 ( .B(clk), .A(\g.we_clk [2328]));
Q_ASSIGN U30447 ( .B(clk), .A(\g.we_clk [2327]));
Q_ASSIGN U30448 ( .B(clk), .A(\g.we_clk [2326]));
Q_ASSIGN U30449 ( .B(clk), .A(\g.we_clk [2325]));
Q_ASSIGN U30450 ( .B(clk), .A(\g.we_clk [2324]));
Q_ASSIGN U30451 ( .B(clk), .A(\g.we_clk [2323]));
Q_ASSIGN U30452 ( .B(clk), .A(\g.we_clk [2322]));
Q_ASSIGN U30453 ( .B(clk), .A(\g.we_clk [2321]));
Q_ASSIGN U30454 ( .B(clk), .A(\g.we_clk [2320]));
Q_ASSIGN U30455 ( .B(clk), .A(\g.we_clk [2319]));
Q_ASSIGN U30456 ( .B(clk), .A(\g.we_clk [2318]));
Q_ASSIGN U30457 ( .B(clk), .A(\g.we_clk [2317]));
Q_ASSIGN U30458 ( .B(clk), .A(\g.we_clk [2316]));
Q_ASSIGN U30459 ( .B(clk), .A(\g.we_clk [2315]));
Q_ASSIGN U30460 ( .B(clk), .A(\g.we_clk [2314]));
Q_ASSIGN U30461 ( .B(clk), .A(\g.we_clk [2313]));
Q_ASSIGN U30462 ( .B(clk), .A(\g.we_clk [2312]));
Q_ASSIGN U30463 ( .B(clk), .A(\g.we_clk [2311]));
Q_ASSIGN U30464 ( .B(clk), .A(\g.we_clk [2310]));
Q_ASSIGN U30465 ( .B(clk), .A(\g.we_clk [2309]));
Q_ASSIGN U30466 ( .B(clk), .A(\g.we_clk [2308]));
Q_ASSIGN U30467 ( .B(clk), .A(\g.we_clk [2307]));
Q_ASSIGN U30468 ( .B(clk), .A(\g.we_clk [2306]));
Q_ASSIGN U30469 ( .B(clk), .A(\g.we_clk [2305]));
Q_ASSIGN U30470 ( .B(clk), .A(\g.we_clk [2304]));
Q_ASSIGN U30471 ( .B(clk), .A(\g.we_clk [2303]));
Q_ASSIGN U30472 ( .B(clk), .A(\g.we_clk [2302]));
Q_ASSIGN U30473 ( .B(clk), .A(\g.we_clk [2301]));
Q_ASSIGN U30474 ( .B(clk), .A(\g.we_clk [2300]));
Q_ASSIGN U30475 ( .B(clk), .A(\g.we_clk [2299]));
Q_ASSIGN U30476 ( .B(clk), .A(\g.we_clk [2298]));
Q_ASSIGN U30477 ( .B(clk), .A(\g.we_clk [2297]));
Q_ASSIGN U30478 ( .B(clk), .A(\g.we_clk [2296]));
Q_ASSIGN U30479 ( .B(clk), .A(\g.we_clk [2295]));
Q_ASSIGN U30480 ( .B(clk), .A(\g.we_clk [2294]));
Q_ASSIGN U30481 ( .B(clk), .A(\g.we_clk [2293]));
Q_ASSIGN U30482 ( .B(clk), .A(\g.we_clk [2292]));
Q_ASSIGN U30483 ( .B(clk), .A(\g.we_clk [2291]));
Q_ASSIGN U30484 ( .B(clk), .A(\g.we_clk [2290]));
Q_ASSIGN U30485 ( .B(clk), .A(\g.we_clk [2289]));
Q_ASSIGN U30486 ( .B(clk), .A(\g.we_clk [2288]));
Q_ASSIGN U30487 ( .B(clk), .A(\g.we_clk [2287]));
Q_ASSIGN U30488 ( .B(clk), .A(\g.we_clk [2286]));
Q_ASSIGN U30489 ( .B(clk), .A(\g.we_clk [2285]));
Q_ASSIGN U30490 ( .B(clk), .A(\g.we_clk [2284]));
Q_ASSIGN U30491 ( .B(clk), .A(\g.we_clk [2283]));
Q_ASSIGN U30492 ( .B(clk), .A(\g.we_clk [2282]));
Q_ASSIGN U30493 ( .B(clk), .A(\g.we_clk [2281]));
Q_ASSIGN U30494 ( .B(clk), .A(\g.we_clk [2280]));
Q_ASSIGN U30495 ( .B(clk), .A(\g.we_clk [2279]));
Q_ASSIGN U30496 ( .B(clk), .A(\g.we_clk [2278]));
Q_ASSIGN U30497 ( .B(clk), .A(\g.we_clk [2277]));
Q_ASSIGN U30498 ( .B(clk), .A(\g.we_clk [2276]));
Q_ASSIGN U30499 ( .B(clk), .A(\g.we_clk [2275]));
Q_ASSIGN U30500 ( .B(clk), .A(\g.we_clk [2274]));
Q_ASSIGN U30501 ( .B(clk), .A(\g.we_clk [2273]));
Q_ASSIGN U30502 ( .B(clk), .A(\g.we_clk [2272]));
Q_ASSIGN U30503 ( .B(clk), .A(\g.we_clk [2271]));
Q_ASSIGN U30504 ( .B(clk), .A(\g.we_clk [2270]));
Q_ASSIGN U30505 ( .B(clk), .A(\g.we_clk [2269]));
Q_ASSIGN U30506 ( .B(clk), .A(\g.we_clk [2268]));
Q_ASSIGN U30507 ( .B(clk), .A(\g.we_clk [2267]));
Q_ASSIGN U30508 ( .B(clk), .A(\g.we_clk [2266]));
Q_ASSIGN U30509 ( .B(clk), .A(\g.we_clk [2265]));
Q_ASSIGN U30510 ( .B(clk), .A(\g.we_clk [2264]));
Q_ASSIGN U30511 ( .B(clk), .A(\g.we_clk [2263]));
Q_ASSIGN U30512 ( .B(clk), .A(\g.we_clk [2262]));
Q_ASSIGN U30513 ( .B(clk), .A(\g.we_clk [2261]));
Q_ASSIGN U30514 ( .B(clk), .A(\g.we_clk [2260]));
Q_ASSIGN U30515 ( .B(clk), .A(\g.we_clk [2259]));
Q_ASSIGN U30516 ( .B(clk), .A(\g.we_clk [2258]));
Q_ASSIGN U30517 ( .B(clk), .A(\g.we_clk [2257]));
Q_ASSIGN U30518 ( .B(clk), .A(\g.we_clk [2256]));
Q_ASSIGN U30519 ( .B(clk), .A(\g.we_clk [2255]));
Q_ASSIGN U30520 ( .B(clk), .A(\g.we_clk [2254]));
Q_ASSIGN U30521 ( .B(clk), .A(\g.we_clk [2253]));
Q_ASSIGN U30522 ( .B(clk), .A(\g.we_clk [2252]));
Q_ASSIGN U30523 ( .B(clk), .A(\g.we_clk [2251]));
Q_ASSIGN U30524 ( .B(clk), .A(\g.we_clk [2250]));
Q_ASSIGN U30525 ( .B(clk), .A(\g.we_clk [2249]));
Q_ASSIGN U30526 ( .B(clk), .A(\g.we_clk [2248]));
Q_ASSIGN U30527 ( .B(clk), .A(\g.we_clk [2247]));
Q_ASSIGN U30528 ( .B(clk), .A(\g.we_clk [2246]));
Q_ASSIGN U30529 ( .B(clk), .A(\g.we_clk [2245]));
Q_ASSIGN U30530 ( .B(clk), .A(\g.we_clk [2244]));
Q_ASSIGN U30531 ( .B(clk), .A(\g.we_clk [2243]));
Q_ASSIGN U30532 ( .B(clk), .A(\g.we_clk [2242]));
Q_ASSIGN U30533 ( .B(clk), .A(\g.we_clk [2241]));
Q_ASSIGN U30534 ( .B(clk), .A(\g.we_clk [2240]));
Q_ASSIGN U30535 ( .B(clk), .A(\g.we_clk [2239]));
Q_ASSIGN U30536 ( .B(clk), .A(\g.we_clk [2238]));
Q_ASSIGN U30537 ( .B(clk), .A(\g.we_clk [2237]));
Q_ASSIGN U30538 ( .B(clk), .A(\g.we_clk [2236]));
Q_ASSIGN U30539 ( .B(clk), .A(\g.we_clk [2235]));
Q_ASSIGN U30540 ( .B(clk), .A(\g.we_clk [2234]));
Q_ASSIGN U30541 ( .B(clk), .A(\g.we_clk [2233]));
Q_ASSIGN U30542 ( .B(clk), .A(\g.we_clk [2232]));
Q_ASSIGN U30543 ( .B(clk), .A(\g.we_clk [2231]));
Q_ASSIGN U30544 ( .B(clk), .A(\g.we_clk [2230]));
Q_ASSIGN U30545 ( .B(clk), .A(\g.we_clk [2229]));
Q_ASSIGN U30546 ( .B(clk), .A(\g.we_clk [2228]));
Q_ASSIGN U30547 ( .B(clk), .A(\g.we_clk [2227]));
Q_ASSIGN U30548 ( .B(clk), .A(\g.we_clk [2226]));
Q_ASSIGN U30549 ( .B(clk), .A(\g.we_clk [2225]));
Q_ASSIGN U30550 ( .B(clk), .A(\g.we_clk [2224]));
Q_ASSIGN U30551 ( .B(clk), .A(\g.we_clk [2223]));
Q_ASSIGN U30552 ( .B(clk), .A(\g.we_clk [2222]));
Q_ASSIGN U30553 ( .B(clk), .A(\g.we_clk [2221]));
Q_ASSIGN U30554 ( .B(clk), .A(\g.we_clk [2220]));
Q_ASSIGN U30555 ( .B(clk), .A(\g.we_clk [2219]));
Q_ASSIGN U30556 ( .B(clk), .A(\g.we_clk [2218]));
Q_ASSIGN U30557 ( .B(clk), .A(\g.we_clk [2217]));
Q_ASSIGN U30558 ( .B(clk), .A(\g.we_clk [2216]));
Q_ASSIGN U30559 ( .B(clk), .A(\g.we_clk [2215]));
Q_ASSIGN U30560 ( .B(clk), .A(\g.we_clk [2214]));
Q_ASSIGN U30561 ( .B(clk), .A(\g.we_clk [2213]));
Q_ASSIGN U30562 ( .B(clk), .A(\g.we_clk [2212]));
Q_ASSIGN U30563 ( .B(clk), .A(\g.we_clk [2211]));
Q_ASSIGN U30564 ( .B(clk), .A(\g.we_clk [2210]));
Q_ASSIGN U30565 ( .B(clk), .A(\g.we_clk [2209]));
Q_ASSIGN U30566 ( .B(clk), .A(\g.we_clk [2208]));
Q_ASSIGN U30567 ( .B(clk), .A(\g.we_clk [2207]));
Q_ASSIGN U30568 ( .B(clk), .A(\g.we_clk [2206]));
Q_ASSIGN U30569 ( .B(clk), .A(\g.we_clk [2205]));
Q_ASSIGN U30570 ( .B(clk), .A(\g.we_clk [2204]));
Q_ASSIGN U30571 ( .B(clk), .A(\g.we_clk [2203]));
Q_ASSIGN U30572 ( .B(clk), .A(\g.we_clk [2202]));
Q_ASSIGN U30573 ( .B(clk), .A(\g.we_clk [2201]));
Q_ASSIGN U30574 ( .B(clk), .A(\g.we_clk [2200]));
Q_ASSIGN U30575 ( .B(clk), .A(\g.we_clk [2199]));
Q_ASSIGN U30576 ( .B(clk), .A(\g.we_clk [2198]));
Q_ASSIGN U30577 ( .B(clk), .A(\g.we_clk [2197]));
Q_ASSIGN U30578 ( .B(clk), .A(\g.we_clk [2196]));
Q_ASSIGN U30579 ( .B(clk), .A(\g.we_clk [2195]));
Q_ASSIGN U30580 ( .B(clk), .A(\g.we_clk [2194]));
Q_ASSIGN U30581 ( .B(clk), .A(\g.we_clk [2193]));
Q_ASSIGN U30582 ( .B(clk), .A(\g.we_clk [2192]));
Q_ASSIGN U30583 ( .B(clk), .A(\g.we_clk [2191]));
Q_ASSIGN U30584 ( .B(clk), .A(\g.we_clk [2190]));
Q_ASSIGN U30585 ( .B(clk), .A(\g.we_clk [2189]));
Q_ASSIGN U30586 ( .B(clk), .A(\g.we_clk [2188]));
Q_ASSIGN U30587 ( .B(clk), .A(\g.we_clk [2187]));
Q_ASSIGN U30588 ( .B(clk), .A(\g.we_clk [2186]));
Q_ASSIGN U30589 ( .B(clk), .A(\g.we_clk [2185]));
Q_ASSIGN U30590 ( .B(clk), .A(\g.we_clk [2184]));
Q_ASSIGN U30591 ( .B(clk), .A(\g.we_clk [2183]));
Q_ASSIGN U30592 ( .B(clk), .A(\g.we_clk [2182]));
Q_ASSIGN U30593 ( .B(clk), .A(\g.we_clk [2181]));
Q_ASSIGN U30594 ( .B(clk), .A(\g.we_clk [2180]));
Q_ASSIGN U30595 ( .B(clk), .A(\g.we_clk [2179]));
Q_ASSIGN U30596 ( .B(clk), .A(\g.we_clk [2178]));
Q_ASSIGN U30597 ( .B(clk), .A(\g.we_clk [2177]));
Q_ASSIGN U30598 ( .B(clk), .A(\g.we_clk [2176]));
Q_ASSIGN U30599 ( .B(clk), .A(\g.we_clk [2175]));
Q_ASSIGN U30600 ( .B(clk), .A(\g.we_clk [2174]));
Q_ASSIGN U30601 ( .B(clk), .A(\g.we_clk [2173]));
Q_ASSIGN U30602 ( .B(clk), .A(\g.we_clk [2172]));
Q_ASSIGN U30603 ( .B(clk), .A(\g.we_clk [2171]));
Q_ASSIGN U30604 ( .B(clk), .A(\g.we_clk [2170]));
Q_ASSIGN U30605 ( .B(clk), .A(\g.we_clk [2169]));
Q_ASSIGN U30606 ( .B(clk), .A(\g.we_clk [2168]));
Q_ASSIGN U30607 ( .B(clk), .A(\g.we_clk [2167]));
Q_ASSIGN U30608 ( .B(clk), .A(\g.we_clk [2166]));
Q_ASSIGN U30609 ( .B(clk), .A(\g.we_clk [2165]));
Q_ASSIGN U30610 ( .B(clk), .A(\g.we_clk [2164]));
Q_ASSIGN U30611 ( .B(clk), .A(\g.we_clk [2163]));
Q_ASSIGN U30612 ( .B(clk), .A(\g.we_clk [2162]));
Q_ASSIGN U30613 ( .B(clk), .A(\g.we_clk [2161]));
Q_ASSIGN U30614 ( .B(clk), .A(\g.we_clk [2160]));
Q_ASSIGN U30615 ( .B(clk), .A(\g.we_clk [2159]));
Q_ASSIGN U30616 ( .B(clk), .A(\g.we_clk [2158]));
Q_ASSIGN U30617 ( .B(clk), .A(\g.we_clk [2157]));
Q_ASSIGN U30618 ( .B(clk), .A(\g.we_clk [2156]));
Q_ASSIGN U30619 ( .B(clk), .A(\g.we_clk [2155]));
Q_ASSIGN U30620 ( .B(clk), .A(\g.we_clk [2154]));
Q_ASSIGN U30621 ( .B(clk), .A(\g.we_clk [2153]));
Q_ASSIGN U30622 ( .B(clk), .A(\g.we_clk [2152]));
Q_ASSIGN U30623 ( .B(clk), .A(\g.we_clk [2151]));
Q_ASSIGN U30624 ( .B(clk), .A(\g.we_clk [2150]));
Q_ASSIGN U30625 ( .B(clk), .A(\g.we_clk [2149]));
Q_ASSIGN U30626 ( .B(clk), .A(\g.we_clk [2148]));
Q_ASSIGN U30627 ( .B(clk), .A(\g.we_clk [2147]));
Q_ASSIGN U30628 ( .B(clk), .A(\g.we_clk [2146]));
Q_ASSIGN U30629 ( .B(clk), .A(\g.we_clk [2145]));
Q_ASSIGN U30630 ( .B(clk), .A(\g.we_clk [2144]));
Q_ASSIGN U30631 ( .B(clk), .A(\g.we_clk [2143]));
Q_ASSIGN U30632 ( .B(clk), .A(\g.we_clk [2142]));
Q_ASSIGN U30633 ( .B(clk), .A(\g.we_clk [2141]));
Q_ASSIGN U30634 ( .B(clk), .A(\g.we_clk [2140]));
Q_ASSIGN U30635 ( .B(clk), .A(\g.we_clk [2139]));
Q_ASSIGN U30636 ( .B(clk), .A(\g.we_clk [2138]));
Q_ASSIGN U30637 ( .B(clk), .A(\g.we_clk [2137]));
Q_ASSIGN U30638 ( .B(clk), .A(\g.we_clk [2136]));
Q_ASSIGN U30639 ( .B(clk), .A(\g.we_clk [2135]));
Q_ASSIGN U30640 ( .B(clk), .A(\g.we_clk [2134]));
Q_ASSIGN U30641 ( .B(clk), .A(\g.we_clk [2133]));
Q_ASSIGN U30642 ( .B(clk), .A(\g.we_clk [2132]));
Q_ASSIGN U30643 ( .B(clk), .A(\g.we_clk [2131]));
Q_ASSIGN U30644 ( .B(clk), .A(\g.we_clk [2130]));
Q_ASSIGN U30645 ( .B(clk), .A(\g.we_clk [2129]));
Q_ASSIGN U30646 ( .B(clk), .A(\g.we_clk [2128]));
Q_ASSIGN U30647 ( .B(clk), .A(\g.we_clk [2127]));
Q_ASSIGN U30648 ( .B(clk), .A(\g.we_clk [2126]));
Q_ASSIGN U30649 ( .B(clk), .A(\g.we_clk [2125]));
Q_ASSIGN U30650 ( .B(clk), .A(\g.we_clk [2124]));
Q_ASSIGN U30651 ( .B(clk), .A(\g.we_clk [2123]));
Q_ASSIGN U30652 ( .B(clk), .A(\g.we_clk [2122]));
Q_ASSIGN U30653 ( .B(clk), .A(\g.we_clk [2121]));
Q_ASSIGN U30654 ( .B(clk), .A(\g.we_clk [2120]));
Q_ASSIGN U30655 ( .B(clk), .A(\g.we_clk [2119]));
Q_ASSIGN U30656 ( .B(clk), .A(\g.we_clk [2118]));
Q_ASSIGN U30657 ( .B(clk), .A(\g.we_clk [2117]));
Q_ASSIGN U30658 ( .B(clk), .A(\g.we_clk [2116]));
Q_ASSIGN U30659 ( .B(clk), .A(\g.we_clk [2115]));
Q_ASSIGN U30660 ( .B(clk), .A(\g.we_clk [2114]));
Q_ASSIGN U30661 ( .B(clk), .A(\g.we_clk [2113]));
Q_ASSIGN U30662 ( .B(clk), .A(\g.we_clk [2112]));
Q_ASSIGN U30663 ( .B(clk), .A(\g.we_clk [2111]));
Q_ASSIGN U30664 ( .B(clk), .A(\g.we_clk [2110]));
Q_ASSIGN U30665 ( .B(clk), .A(\g.we_clk [2109]));
Q_ASSIGN U30666 ( .B(clk), .A(\g.we_clk [2108]));
Q_ASSIGN U30667 ( .B(clk), .A(\g.we_clk [2107]));
Q_ASSIGN U30668 ( .B(clk), .A(\g.we_clk [2106]));
Q_ASSIGN U30669 ( .B(clk), .A(\g.we_clk [2105]));
Q_ASSIGN U30670 ( .B(clk), .A(\g.we_clk [2104]));
Q_ASSIGN U30671 ( .B(clk), .A(\g.we_clk [2103]));
Q_ASSIGN U30672 ( .B(clk), .A(\g.we_clk [2102]));
Q_ASSIGN U30673 ( .B(clk), .A(\g.we_clk [2101]));
Q_ASSIGN U30674 ( .B(clk), .A(\g.we_clk [2100]));
Q_ASSIGN U30675 ( .B(clk), .A(\g.we_clk [2099]));
Q_ASSIGN U30676 ( .B(clk), .A(\g.we_clk [2098]));
Q_ASSIGN U30677 ( .B(clk), .A(\g.we_clk [2097]));
Q_ASSIGN U30678 ( .B(clk), .A(\g.we_clk [2096]));
Q_ASSIGN U30679 ( .B(clk), .A(\g.we_clk [2095]));
Q_ASSIGN U30680 ( .B(clk), .A(\g.we_clk [2094]));
Q_ASSIGN U30681 ( .B(clk), .A(\g.we_clk [2093]));
Q_ASSIGN U30682 ( .B(clk), .A(\g.we_clk [2092]));
Q_ASSIGN U30683 ( .B(clk), .A(\g.we_clk [2091]));
Q_ASSIGN U30684 ( .B(clk), .A(\g.we_clk [2090]));
Q_ASSIGN U30685 ( .B(clk), .A(\g.we_clk [2089]));
Q_ASSIGN U30686 ( .B(clk), .A(\g.we_clk [2088]));
Q_ASSIGN U30687 ( .B(clk), .A(\g.we_clk [2087]));
Q_ASSIGN U30688 ( .B(clk), .A(\g.we_clk [2086]));
Q_ASSIGN U30689 ( .B(clk), .A(\g.we_clk [2085]));
Q_ASSIGN U30690 ( .B(clk), .A(\g.we_clk [2084]));
Q_ASSIGN U30691 ( .B(clk), .A(\g.we_clk [2083]));
Q_ASSIGN U30692 ( .B(clk), .A(\g.we_clk [2082]));
Q_ASSIGN U30693 ( .B(clk), .A(\g.we_clk [2081]));
Q_ASSIGN U30694 ( .B(clk), .A(\g.we_clk [2080]));
Q_ASSIGN U30695 ( .B(clk), .A(\g.we_clk [2079]));
Q_ASSIGN U30696 ( .B(clk), .A(\g.we_clk [2078]));
Q_ASSIGN U30697 ( .B(clk), .A(\g.we_clk [2077]));
Q_ASSIGN U30698 ( .B(clk), .A(\g.we_clk [2076]));
Q_ASSIGN U30699 ( .B(clk), .A(\g.we_clk [2075]));
Q_ASSIGN U30700 ( .B(clk), .A(\g.we_clk [2074]));
Q_ASSIGN U30701 ( .B(clk), .A(\g.we_clk [2073]));
Q_ASSIGN U30702 ( .B(clk), .A(\g.we_clk [2072]));
Q_ASSIGN U30703 ( .B(clk), .A(\g.we_clk [2071]));
Q_ASSIGN U30704 ( .B(clk), .A(\g.we_clk [2070]));
Q_ASSIGN U30705 ( .B(clk), .A(\g.we_clk [2069]));
Q_ASSIGN U30706 ( .B(clk), .A(\g.we_clk [2068]));
Q_ASSIGN U30707 ( .B(clk), .A(\g.we_clk [2067]));
Q_ASSIGN U30708 ( .B(clk), .A(\g.we_clk [2066]));
Q_ASSIGN U30709 ( .B(clk), .A(\g.we_clk [2065]));
Q_ASSIGN U30710 ( .B(clk), .A(\g.we_clk [2064]));
Q_ASSIGN U30711 ( .B(clk), .A(\g.we_clk [2063]));
Q_ASSIGN U30712 ( .B(clk), .A(\g.we_clk [2062]));
Q_ASSIGN U30713 ( .B(clk), .A(\g.we_clk [2061]));
Q_ASSIGN U30714 ( .B(clk), .A(\g.we_clk [2060]));
Q_ASSIGN U30715 ( .B(clk), .A(\g.we_clk [2059]));
Q_ASSIGN U30716 ( .B(clk), .A(\g.we_clk [2058]));
Q_ASSIGN U30717 ( .B(clk), .A(\g.we_clk [2057]));
Q_ASSIGN U30718 ( .B(clk), .A(\g.we_clk [2056]));
Q_ASSIGN U30719 ( .B(clk), .A(\g.we_clk [2055]));
Q_ASSIGN U30720 ( .B(clk), .A(\g.we_clk [2054]));
Q_ASSIGN U30721 ( .B(clk), .A(\g.we_clk [2053]));
Q_ASSIGN U30722 ( .B(clk), .A(\g.we_clk [2052]));
Q_ASSIGN U30723 ( .B(clk), .A(\g.we_clk [2051]));
Q_ASSIGN U30724 ( .B(clk), .A(\g.we_clk [2050]));
Q_ASSIGN U30725 ( .B(clk), .A(\g.we_clk [2049]));
Q_ASSIGN U30726 ( .B(clk), .A(\g.we_clk [2048]));
Q_ASSIGN U30727 ( .B(clk), .A(\g.we_clk [2047]));
Q_ASSIGN U30728 ( .B(clk), .A(\g.we_clk [2046]));
Q_ASSIGN U30729 ( .B(clk), .A(\g.we_clk [2045]));
Q_ASSIGN U30730 ( .B(clk), .A(\g.we_clk [2044]));
Q_ASSIGN U30731 ( .B(clk), .A(\g.we_clk [2043]));
Q_ASSIGN U30732 ( .B(clk), .A(\g.we_clk [2042]));
Q_ASSIGN U30733 ( .B(clk), .A(\g.we_clk [2041]));
Q_ASSIGN U30734 ( .B(clk), .A(\g.we_clk [2040]));
Q_ASSIGN U30735 ( .B(clk), .A(\g.we_clk [2039]));
Q_ASSIGN U30736 ( .B(clk), .A(\g.we_clk [2038]));
Q_ASSIGN U30737 ( .B(clk), .A(\g.we_clk [2037]));
Q_ASSIGN U30738 ( .B(clk), .A(\g.we_clk [2036]));
Q_ASSIGN U30739 ( .B(clk), .A(\g.we_clk [2035]));
Q_ASSIGN U30740 ( .B(clk), .A(\g.we_clk [2034]));
Q_ASSIGN U30741 ( .B(clk), .A(\g.we_clk [2033]));
Q_ASSIGN U30742 ( .B(clk), .A(\g.we_clk [2032]));
Q_ASSIGN U30743 ( .B(clk), .A(\g.we_clk [2031]));
Q_ASSIGN U30744 ( .B(clk), .A(\g.we_clk [2030]));
Q_ASSIGN U30745 ( .B(clk), .A(\g.we_clk [2029]));
Q_ASSIGN U30746 ( .B(clk), .A(\g.we_clk [2028]));
Q_ASSIGN U30747 ( .B(clk), .A(\g.we_clk [2027]));
Q_ASSIGN U30748 ( .B(clk), .A(\g.we_clk [2026]));
Q_ASSIGN U30749 ( .B(clk), .A(\g.we_clk [2025]));
Q_ASSIGN U30750 ( .B(clk), .A(\g.we_clk [2024]));
Q_ASSIGN U30751 ( .B(clk), .A(\g.we_clk [2023]));
Q_ASSIGN U30752 ( .B(clk), .A(\g.we_clk [2022]));
Q_ASSIGN U30753 ( .B(clk), .A(\g.we_clk [2021]));
Q_ASSIGN U30754 ( .B(clk), .A(\g.we_clk [2020]));
Q_ASSIGN U30755 ( .B(clk), .A(\g.we_clk [2019]));
Q_ASSIGN U30756 ( .B(clk), .A(\g.we_clk [2018]));
Q_ASSIGN U30757 ( .B(clk), .A(\g.we_clk [2017]));
Q_ASSIGN U30758 ( .B(clk), .A(\g.we_clk [2016]));
Q_ASSIGN U30759 ( .B(clk), .A(\g.we_clk [2015]));
Q_ASSIGN U30760 ( .B(clk), .A(\g.we_clk [2014]));
Q_ASSIGN U30761 ( .B(clk), .A(\g.we_clk [2013]));
Q_ASSIGN U30762 ( .B(clk), .A(\g.we_clk [2012]));
Q_ASSIGN U30763 ( .B(clk), .A(\g.we_clk [2011]));
Q_ASSIGN U30764 ( .B(clk), .A(\g.we_clk [2010]));
Q_ASSIGN U30765 ( .B(clk), .A(\g.we_clk [2009]));
Q_ASSIGN U30766 ( .B(clk), .A(\g.we_clk [2008]));
Q_ASSIGN U30767 ( .B(clk), .A(\g.we_clk [2007]));
Q_ASSIGN U30768 ( .B(clk), .A(\g.we_clk [2006]));
Q_ASSIGN U30769 ( .B(clk), .A(\g.we_clk [2005]));
Q_ASSIGN U30770 ( .B(clk), .A(\g.we_clk [2004]));
Q_ASSIGN U30771 ( .B(clk), .A(\g.we_clk [2003]));
Q_ASSIGN U30772 ( .B(clk), .A(\g.we_clk [2002]));
Q_ASSIGN U30773 ( .B(clk), .A(\g.we_clk [2001]));
Q_ASSIGN U30774 ( .B(clk), .A(\g.we_clk [2000]));
Q_ASSIGN U30775 ( .B(clk), .A(\g.we_clk [1999]));
Q_ASSIGN U30776 ( .B(clk), .A(\g.we_clk [1998]));
Q_ASSIGN U30777 ( .B(clk), .A(\g.we_clk [1997]));
Q_ASSIGN U30778 ( .B(clk), .A(\g.we_clk [1996]));
Q_ASSIGN U30779 ( .B(clk), .A(\g.we_clk [1995]));
Q_ASSIGN U30780 ( .B(clk), .A(\g.we_clk [1994]));
Q_ASSIGN U30781 ( .B(clk), .A(\g.we_clk [1993]));
Q_ASSIGN U30782 ( .B(clk), .A(\g.we_clk [1992]));
Q_ASSIGN U30783 ( .B(clk), .A(\g.we_clk [1991]));
Q_ASSIGN U30784 ( .B(clk), .A(\g.we_clk [1990]));
Q_ASSIGN U30785 ( .B(clk), .A(\g.we_clk [1989]));
Q_ASSIGN U30786 ( .B(clk), .A(\g.we_clk [1988]));
Q_ASSIGN U30787 ( .B(clk), .A(\g.we_clk [1987]));
Q_ASSIGN U30788 ( .B(clk), .A(\g.we_clk [1986]));
Q_ASSIGN U30789 ( .B(clk), .A(\g.we_clk [1985]));
Q_ASSIGN U30790 ( .B(clk), .A(\g.we_clk [1984]));
Q_ASSIGN U30791 ( .B(clk), .A(\g.we_clk [1983]));
Q_ASSIGN U30792 ( .B(clk), .A(\g.we_clk [1982]));
Q_ASSIGN U30793 ( .B(clk), .A(\g.we_clk [1981]));
Q_ASSIGN U30794 ( .B(clk), .A(\g.we_clk [1980]));
Q_ASSIGN U30795 ( .B(clk), .A(\g.we_clk [1979]));
Q_ASSIGN U30796 ( .B(clk), .A(\g.we_clk [1978]));
Q_ASSIGN U30797 ( .B(clk), .A(\g.we_clk [1977]));
Q_ASSIGN U30798 ( .B(clk), .A(\g.we_clk [1976]));
Q_ASSIGN U30799 ( .B(clk), .A(\g.we_clk [1975]));
Q_ASSIGN U30800 ( .B(clk), .A(\g.we_clk [1974]));
Q_ASSIGN U30801 ( .B(clk), .A(\g.we_clk [1973]));
Q_ASSIGN U30802 ( .B(clk), .A(\g.we_clk [1972]));
Q_ASSIGN U30803 ( .B(clk), .A(\g.we_clk [1971]));
Q_ASSIGN U30804 ( .B(clk), .A(\g.we_clk [1970]));
Q_ASSIGN U30805 ( .B(clk), .A(\g.we_clk [1969]));
Q_ASSIGN U30806 ( .B(clk), .A(\g.we_clk [1968]));
Q_ASSIGN U30807 ( .B(clk), .A(\g.we_clk [1967]));
Q_ASSIGN U30808 ( .B(clk), .A(\g.we_clk [1966]));
Q_ASSIGN U30809 ( .B(clk), .A(\g.we_clk [1965]));
Q_ASSIGN U30810 ( .B(clk), .A(\g.we_clk [1964]));
Q_ASSIGN U30811 ( .B(clk), .A(\g.we_clk [1963]));
Q_ASSIGN U30812 ( .B(clk), .A(\g.we_clk [1962]));
Q_ASSIGN U30813 ( .B(clk), .A(\g.we_clk [1961]));
Q_ASSIGN U30814 ( .B(clk), .A(\g.we_clk [1960]));
Q_ASSIGN U30815 ( .B(clk), .A(\g.we_clk [1959]));
Q_ASSIGN U30816 ( .B(clk), .A(\g.we_clk [1958]));
Q_ASSIGN U30817 ( .B(clk), .A(\g.we_clk [1957]));
Q_ASSIGN U30818 ( .B(clk), .A(\g.we_clk [1956]));
Q_ASSIGN U30819 ( .B(clk), .A(\g.we_clk [1955]));
Q_ASSIGN U30820 ( .B(clk), .A(\g.we_clk [1954]));
Q_ASSIGN U30821 ( .B(clk), .A(\g.we_clk [1953]));
Q_ASSIGN U30822 ( .B(clk), .A(\g.we_clk [1952]));
Q_ASSIGN U30823 ( .B(clk), .A(\g.we_clk [1951]));
Q_ASSIGN U30824 ( .B(clk), .A(\g.we_clk [1950]));
Q_ASSIGN U30825 ( .B(clk), .A(\g.we_clk [1949]));
Q_ASSIGN U30826 ( .B(clk), .A(\g.we_clk [1948]));
Q_ASSIGN U30827 ( .B(clk), .A(\g.we_clk [1947]));
Q_ASSIGN U30828 ( .B(clk), .A(\g.we_clk [1946]));
Q_ASSIGN U30829 ( .B(clk), .A(\g.we_clk [1945]));
Q_ASSIGN U30830 ( .B(clk), .A(\g.we_clk [1944]));
Q_ASSIGN U30831 ( .B(clk), .A(\g.we_clk [1943]));
Q_ASSIGN U30832 ( .B(clk), .A(\g.we_clk [1942]));
Q_ASSIGN U30833 ( .B(clk), .A(\g.we_clk [1941]));
Q_ASSIGN U30834 ( .B(clk), .A(\g.we_clk [1940]));
Q_ASSIGN U30835 ( .B(clk), .A(\g.we_clk [1939]));
Q_ASSIGN U30836 ( .B(clk), .A(\g.we_clk [1938]));
Q_ASSIGN U30837 ( .B(clk), .A(\g.we_clk [1937]));
Q_ASSIGN U30838 ( .B(clk), .A(\g.we_clk [1936]));
Q_ASSIGN U30839 ( .B(clk), .A(\g.we_clk [1935]));
Q_ASSIGN U30840 ( .B(clk), .A(\g.we_clk [1934]));
Q_ASSIGN U30841 ( .B(clk), .A(\g.we_clk [1933]));
Q_ASSIGN U30842 ( .B(clk), .A(\g.we_clk [1932]));
Q_ASSIGN U30843 ( .B(clk), .A(\g.we_clk [1931]));
Q_ASSIGN U30844 ( .B(clk), .A(\g.we_clk [1930]));
Q_ASSIGN U30845 ( .B(clk), .A(\g.we_clk [1929]));
Q_ASSIGN U30846 ( .B(clk), .A(\g.we_clk [1928]));
Q_ASSIGN U30847 ( .B(clk), .A(\g.we_clk [1927]));
Q_ASSIGN U30848 ( .B(clk), .A(\g.we_clk [1926]));
Q_ASSIGN U30849 ( .B(clk), .A(\g.we_clk [1925]));
Q_ASSIGN U30850 ( .B(clk), .A(\g.we_clk [1924]));
Q_ASSIGN U30851 ( .B(clk), .A(\g.we_clk [1923]));
Q_ASSIGN U30852 ( .B(clk), .A(\g.we_clk [1922]));
Q_ASSIGN U30853 ( .B(clk), .A(\g.we_clk [1921]));
Q_ASSIGN U30854 ( .B(clk), .A(\g.we_clk [1920]));
Q_ASSIGN U30855 ( .B(clk), .A(\g.we_clk [1919]));
Q_ASSIGN U30856 ( .B(clk), .A(\g.we_clk [1918]));
Q_ASSIGN U30857 ( .B(clk), .A(\g.we_clk [1917]));
Q_ASSIGN U30858 ( .B(clk), .A(\g.we_clk [1916]));
Q_ASSIGN U30859 ( .B(clk), .A(\g.we_clk [1915]));
Q_ASSIGN U30860 ( .B(clk), .A(\g.we_clk [1914]));
Q_ASSIGN U30861 ( .B(clk), .A(\g.we_clk [1913]));
Q_ASSIGN U30862 ( .B(clk), .A(\g.we_clk [1912]));
Q_ASSIGN U30863 ( .B(clk), .A(\g.we_clk [1911]));
Q_ASSIGN U30864 ( .B(clk), .A(\g.we_clk [1910]));
Q_ASSIGN U30865 ( .B(clk), .A(\g.we_clk [1909]));
Q_ASSIGN U30866 ( .B(clk), .A(\g.we_clk [1908]));
Q_ASSIGN U30867 ( .B(clk), .A(\g.we_clk [1907]));
Q_ASSIGN U30868 ( .B(clk), .A(\g.we_clk [1906]));
Q_ASSIGN U30869 ( .B(clk), .A(\g.we_clk [1905]));
Q_ASSIGN U30870 ( .B(clk), .A(\g.we_clk [1904]));
Q_ASSIGN U30871 ( .B(clk), .A(\g.we_clk [1903]));
Q_ASSIGN U30872 ( .B(clk), .A(\g.we_clk [1902]));
Q_ASSIGN U30873 ( .B(clk), .A(\g.we_clk [1901]));
Q_ASSIGN U30874 ( .B(clk), .A(\g.we_clk [1900]));
Q_ASSIGN U30875 ( .B(clk), .A(\g.we_clk [1899]));
Q_ASSIGN U30876 ( .B(clk), .A(\g.we_clk [1898]));
Q_ASSIGN U30877 ( .B(clk), .A(\g.we_clk [1897]));
Q_ASSIGN U30878 ( .B(clk), .A(\g.we_clk [1896]));
Q_ASSIGN U30879 ( .B(clk), .A(\g.we_clk [1895]));
Q_ASSIGN U30880 ( .B(clk), .A(\g.we_clk [1894]));
Q_ASSIGN U30881 ( .B(clk), .A(\g.we_clk [1893]));
Q_ASSIGN U30882 ( .B(clk), .A(\g.we_clk [1892]));
Q_ASSIGN U30883 ( .B(clk), .A(\g.we_clk [1891]));
Q_ASSIGN U30884 ( .B(clk), .A(\g.we_clk [1890]));
Q_ASSIGN U30885 ( .B(clk), .A(\g.we_clk [1889]));
Q_ASSIGN U30886 ( .B(clk), .A(\g.we_clk [1888]));
Q_ASSIGN U30887 ( .B(clk), .A(\g.we_clk [1887]));
Q_ASSIGN U30888 ( .B(clk), .A(\g.we_clk [1886]));
Q_ASSIGN U30889 ( .B(clk), .A(\g.we_clk [1885]));
Q_ASSIGN U30890 ( .B(clk), .A(\g.we_clk [1884]));
Q_ASSIGN U30891 ( .B(clk), .A(\g.we_clk [1883]));
Q_ASSIGN U30892 ( .B(clk), .A(\g.we_clk [1882]));
Q_ASSIGN U30893 ( .B(clk), .A(\g.we_clk [1881]));
Q_ASSIGN U30894 ( .B(clk), .A(\g.we_clk [1880]));
Q_ASSIGN U30895 ( .B(clk), .A(\g.we_clk [1879]));
Q_ASSIGN U30896 ( .B(clk), .A(\g.we_clk [1878]));
Q_ASSIGN U30897 ( .B(clk), .A(\g.we_clk [1877]));
Q_ASSIGN U30898 ( .B(clk), .A(\g.we_clk [1876]));
Q_ASSIGN U30899 ( .B(clk), .A(\g.we_clk [1875]));
Q_ASSIGN U30900 ( .B(clk), .A(\g.we_clk [1874]));
Q_ASSIGN U30901 ( .B(clk), .A(\g.we_clk [1873]));
Q_ASSIGN U30902 ( .B(clk), .A(\g.we_clk [1872]));
Q_ASSIGN U30903 ( .B(clk), .A(\g.we_clk [1871]));
Q_ASSIGN U30904 ( .B(clk), .A(\g.we_clk [1870]));
Q_ASSIGN U30905 ( .B(clk), .A(\g.we_clk [1869]));
Q_ASSIGN U30906 ( .B(clk), .A(\g.we_clk [1868]));
Q_ASSIGN U30907 ( .B(clk), .A(\g.we_clk [1867]));
Q_ASSIGN U30908 ( .B(clk), .A(\g.we_clk [1866]));
Q_ASSIGN U30909 ( .B(clk), .A(\g.we_clk [1865]));
Q_ASSIGN U30910 ( .B(clk), .A(\g.we_clk [1864]));
Q_ASSIGN U30911 ( .B(clk), .A(\g.we_clk [1863]));
Q_ASSIGN U30912 ( .B(clk), .A(\g.we_clk [1862]));
Q_ASSIGN U30913 ( .B(clk), .A(\g.we_clk [1861]));
Q_ASSIGN U30914 ( .B(clk), .A(\g.we_clk [1860]));
Q_ASSIGN U30915 ( .B(clk), .A(\g.we_clk [1859]));
Q_ASSIGN U30916 ( .B(clk), .A(\g.we_clk [1858]));
Q_ASSIGN U30917 ( .B(clk), .A(\g.we_clk [1857]));
Q_ASSIGN U30918 ( .B(clk), .A(\g.we_clk [1856]));
Q_ASSIGN U30919 ( .B(clk), .A(\g.we_clk [1855]));
Q_ASSIGN U30920 ( .B(clk), .A(\g.we_clk [1854]));
Q_ASSIGN U30921 ( .B(clk), .A(\g.we_clk [1853]));
Q_ASSIGN U30922 ( .B(clk), .A(\g.we_clk [1852]));
Q_ASSIGN U30923 ( .B(clk), .A(\g.we_clk [1851]));
Q_ASSIGN U30924 ( .B(clk), .A(\g.we_clk [1850]));
Q_ASSIGN U30925 ( .B(clk), .A(\g.we_clk [1849]));
Q_ASSIGN U30926 ( .B(clk), .A(\g.we_clk [1848]));
Q_ASSIGN U30927 ( .B(clk), .A(\g.we_clk [1847]));
Q_ASSIGN U30928 ( .B(clk), .A(\g.we_clk [1846]));
Q_ASSIGN U30929 ( .B(clk), .A(\g.we_clk [1845]));
Q_ASSIGN U30930 ( .B(clk), .A(\g.we_clk [1844]));
Q_ASSIGN U30931 ( .B(clk), .A(\g.we_clk [1843]));
Q_ASSIGN U30932 ( .B(clk), .A(\g.we_clk [1842]));
Q_ASSIGN U30933 ( .B(clk), .A(\g.we_clk [1841]));
Q_ASSIGN U30934 ( .B(clk), .A(\g.we_clk [1840]));
Q_ASSIGN U30935 ( .B(clk), .A(\g.we_clk [1839]));
Q_ASSIGN U30936 ( .B(clk), .A(\g.we_clk [1838]));
Q_ASSIGN U30937 ( .B(clk), .A(\g.we_clk [1837]));
Q_ASSIGN U30938 ( .B(clk), .A(\g.we_clk [1836]));
Q_ASSIGN U30939 ( .B(clk), .A(\g.we_clk [1835]));
Q_ASSIGN U30940 ( .B(clk), .A(\g.we_clk [1834]));
Q_ASSIGN U30941 ( .B(clk), .A(\g.we_clk [1833]));
Q_ASSIGN U30942 ( .B(clk), .A(\g.we_clk [1832]));
Q_ASSIGN U30943 ( .B(clk), .A(\g.we_clk [1831]));
Q_ASSIGN U30944 ( .B(clk), .A(\g.we_clk [1830]));
Q_ASSIGN U30945 ( .B(clk), .A(\g.we_clk [1829]));
Q_ASSIGN U30946 ( .B(clk), .A(\g.we_clk [1828]));
Q_ASSIGN U30947 ( .B(clk), .A(\g.we_clk [1827]));
Q_ASSIGN U30948 ( .B(clk), .A(\g.we_clk [1826]));
Q_ASSIGN U30949 ( .B(clk), .A(\g.we_clk [1825]));
Q_ASSIGN U30950 ( .B(clk), .A(\g.we_clk [1824]));
Q_ASSIGN U30951 ( .B(clk), .A(\g.we_clk [1823]));
Q_ASSIGN U30952 ( .B(clk), .A(\g.we_clk [1822]));
Q_ASSIGN U30953 ( .B(clk), .A(\g.we_clk [1821]));
Q_ASSIGN U30954 ( .B(clk), .A(\g.we_clk [1820]));
Q_ASSIGN U30955 ( .B(clk), .A(\g.we_clk [1819]));
Q_ASSIGN U30956 ( .B(clk), .A(\g.we_clk [1818]));
Q_ASSIGN U30957 ( .B(clk), .A(\g.we_clk [1817]));
Q_ASSIGN U30958 ( .B(clk), .A(\g.we_clk [1816]));
Q_ASSIGN U30959 ( .B(clk), .A(\g.we_clk [1815]));
Q_ASSIGN U30960 ( .B(clk), .A(\g.we_clk [1814]));
Q_ASSIGN U30961 ( .B(clk), .A(\g.we_clk [1813]));
Q_ASSIGN U30962 ( .B(clk), .A(\g.we_clk [1812]));
Q_ASSIGN U30963 ( .B(clk), .A(\g.we_clk [1811]));
Q_ASSIGN U30964 ( .B(clk), .A(\g.we_clk [1810]));
Q_ASSIGN U30965 ( .B(clk), .A(\g.we_clk [1809]));
Q_ASSIGN U30966 ( .B(clk), .A(\g.we_clk [1808]));
Q_ASSIGN U30967 ( .B(clk), .A(\g.we_clk [1807]));
Q_ASSIGN U30968 ( .B(clk), .A(\g.we_clk [1806]));
Q_ASSIGN U30969 ( .B(clk), .A(\g.we_clk [1805]));
Q_ASSIGN U30970 ( .B(clk), .A(\g.we_clk [1804]));
Q_ASSIGN U30971 ( .B(clk), .A(\g.we_clk [1803]));
Q_ASSIGN U30972 ( .B(clk), .A(\g.we_clk [1802]));
Q_ASSIGN U30973 ( .B(clk), .A(\g.we_clk [1801]));
Q_ASSIGN U30974 ( .B(clk), .A(\g.we_clk [1800]));
Q_ASSIGN U30975 ( .B(clk), .A(\g.we_clk [1799]));
Q_ASSIGN U30976 ( .B(clk), .A(\g.we_clk [1798]));
Q_ASSIGN U30977 ( .B(clk), .A(\g.we_clk [1797]));
Q_ASSIGN U30978 ( .B(clk), .A(\g.we_clk [1796]));
Q_ASSIGN U30979 ( .B(clk), .A(\g.we_clk [1795]));
Q_ASSIGN U30980 ( .B(clk), .A(\g.we_clk [1794]));
Q_ASSIGN U30981 ( .B(clk), .A(\g.we_clk [1793]));
Q_ASSIGN U30982 ( .B(clk), .A(\g.we_clk [1792]));
Q_ASSIGN U30983 ( .B(clk), .A(\g.we_clk [1791]));
Q_ASSIGN U30984 ( .B(clk), .A(\g.we_clk [1790]));
Q_ASSIGN U30985 ( .B(clk), .A(\g.we_clk [1789]));
Q_ASSIGN U30986 ( .B(clk), .A(\g.we_clk [1788]));
Q_ASSIGN U30987 ( .B(clk), .A(\g.we_clk [1787]));
Q_ASSIGN U30988 ( .B(clk), .A(\g.we_clk [1786]));
Q_ASSIGN U30989 ( .B(clk), .A(\g.we_clk [1785]));
Q_ASSIGN U30990 ( .B(clk), .A(\g.we_clk [1784]));
Q_ASSIGN U30991 ( .B(clk), .A(\g.we_clk [1783]));
Q_ASSIGN U30992 ( .B(clk), .A(\g.we_clk [1782]));
Q_ASSIGN U30993 ( .B(clk), .A(\g.we_clk [1781]));
Q_ASSIGN U30994 ( .B(clk), .A(\g.we_clk [1780]));
Q_ASSIGN U30995 ( .B(clk), .A(\g.we_clk [1779]));
Q_ASSIGN U30996 ( .B(clk), .A(\g.we_clk [1778]));
Q_ASSIGN U30997 ( .B(clk), .A(\g.we_clk [1777]));
Q_ASSIGN U30998 ( .B(clk), .A(\g.we_clk [1776]));
Q_ASSIGN U30999 ( .B(clk), .A(\g.we_clk [1775]));
Q_ASSIGN U31000 ( .B(clk), .A(\g.we_clk [1774]));
Q_ASSIGN U31001 ( .B(clk), .A(\g.we_clk [1773]));
Q_ASSIGN U31002 ( .B(clk), .A(\g.we_clk [1772]));
Q_ASSIGN U31003 ( .B(clk), .A(\g.we_clk [1771]));
Q_ASSIGN U31004 ( .B(clk), .A(\g.we_clk [1770]));
Q_ASSIGN U31005 ( .B(clk), .A(\g.we_clk [1769]));
Q_ASSIGN U31006 ( .B(clk), .A(\g.we_clk [1768]));
Q_ASSIGN U31007 ( .B(clk), .A(\g.we_clk [1767]));
Q_ASSIGN U31008 ( .B(clk), .A(\g.we_clk [1766]));
Q_ASSIGN U31009 ( .B(clk), .A(\g.we_clk [1765]));
Q_ASSIGN U31010 ( .B(clk), .A(\g.we_clk [1764]));
Q_ASSIGN U31011 ( .B(clk), .A(\g.we_clk [1763]));
Q_ASSIGN U31012 ( .B(clk), .A(\g.we_clk [1762]));
Q_ASSIGN U31013 ( .B(clk), .A(\g.we_clk [1761]));
Q_ASSIGN U31014 ( .B(clk), .A(\g.we_clk [1760]));
Q_ASSIGN U31015 ( .B(clk), .A(\g.we_clk [1759]));
Q_ASSIGN U31016 ( .B(clk), .A(\g.we_clk [1758]));
Q_ASSIGN U31017 ( .B(clk), .A(\g.we_clk [1757]));
Q_ASSIGN U31018 ( .B(clk), .A(\g.we_clk [1756]));
Q_ASSIGN U31019 ( .B(clk), .A(\g.we_clk [1755]));
Q_ASSIGN U31020 ( .B(clk), .A(\g.we_clk [1754]));
Q_ASSIGN U31021 ( .B(clk), .A(\g.we_clk [1753]));
Q_ASSIGN U31022 ( .B(clk), .A(\g.we_clk [1752]));
Q_ASSIGN U31023 ( .B(clk), .A(\g.we_clk [1751]));
Q_ASSIGN U31024 ( .B(clk), .A(\g.we_clk [1750]));
Q_ASSIGN U31025 ( .B(clk), .A(\g.we_clk [1749]));
Q_ASSIGN U31026 ( .B(clk), .A(\g.we_clk [1748]));
Q_ASSIGN U31027 ( .B(clk), .A(\g.we_clk [1747]));
Q_ASSIGN U31028 ( .B(clk), .A(\g.we_clk [1746]));
Q_ASSIGN U31029 ( .B(clk), .A(\g.we_clk [1745]));
Q_ASSIGN U31030 ( .B(clk), .A(\g.we_clk [1744]));
Q_ASSIGN U31031 ( .B(clk), .A(\g.we_clk [1743]));
Q_ASSIGN U31032 ( .B(clk), .A(\g.we_clk [1742]));
Q_ASSIGN U31033 ( .B(clk), .A(\g.we_clk [1741]));
Q_ASSIGN U31034 ( .B(clk), .A(\g.we_clk [1740]));
Q_ASSIGN U31035 ( .B(clk), .A(\g.we_clk [1739]));
Q_ASSIGN U31036 ( .B(clk), .A(\g.we_clk [1738]));
Q_ASSIGN U31037 ( .B(clk), .A(\g.we_clk [1737]));
Q_ASSIGN U31038 ( .B(clk), .A(\g.we_clk [1736]));
Q_ASSIGN U31039 ( .B(clk), .A(\g.we_clk [1735]));
Q_ASSIGN U31040 ( .B(clk), .A(\g.we_clk [1734]));
Q_ASSIGN U31041 ( .B(clk), .A(\g.we_clk [1733]));
Q_ASSIGN U31042 ( .B(clk), .A(\g.we_clk [1732]));
Q_ASSIGN U31043 ( .B(clk), .A(\g.we_clk [1731]));
Q_ASSIGN U31044 ( .B(clk), .A(\g.we_clk [1730]));
Q_ASSIGN U31045 ( .B(clk), .A(\g.we_clk [1729]));
Q_ASSIGN U31046 ( .B(clk), .A(\g.we_clk [1728]));
Q_ASSIGN U31047 ( .B(clk), .A(\g.we_clk [1727]));
Q_ASSIGN U31048 ( .B(clk), .A(\g.we_clk [1726]));
Q_ASSIGN U31049 ( .B(clk), .A(\g.we_clk [1725]));
Q_ASSIGN U31050 ( .B(clk), .A(\g.we_clk [1724]));
Q_ASSIGN U31051 ( .B(clk), .A(\g.we_clk [1723]));
Q_ASSIGN U31052 ( .B(clk), .A(\g.we_clk [1722]));
Q_ASSIGN U31053 ( .B(clk), .A(\g.we_clk [1721]));
Q_ASSIGN U31054 ( .B(clk), .A(\g.we_clk [1720]));
Q_ASSIGN U31055 ( .B(clk), .A(\g.we_clk [1719]));
Q_ASSIGN U31056 ( .B(clk), .A(\g.we_clk [1718]));
Q_ASSIGN U31057 ( .B(clk), .A(\g.we_clk [1717]));
Q_ASSIGN U31058 ( .B(clk), .A(\g.we_clk [1716]));
Q_ASSIGN U31059 ( .B(clk), .A(\g.we_clk [1715]));
Q_ASSIGN U31060 ( .B(clk), .A(\g.we_clk [1714]));
Q_ASSIGN U31061 ( .B(clk), .A(\g.we_clk [1713]));
Q_ASSIGN U31062 ( .B(clk), .A(\g.we_clk [1712]));
Q_ASSIGN U31063 ( .B(clk), .A(\g.we_clk [1711]));
Q_ASSIGN U31064 ( .B(clk), .A(\g.we_clk [1710]));
Q_ASSIGN U31065 ( .B(clk), .A(\g.we_clk [1709]));
Q_ASSIGN U31066 ( .B(clk), .A(\g.we_clk [1708]));
Q_ASSIGN U31067 ( .B(clk), .A(\g.we_clk [1707]));
Q_ASSIGN U31068 ( .B(clk), .A(\g.we_clk [1706]));
Q_ASSIGN U31069 ( .B(clk), .A(\g.we_clk [1705]));
Q_ASSIGN U31070 ( .B(clk), .A(\g.we_clk [1704]));
Q_ASSIGN U31071 ( .B(clk), .A(\g.we_clk [1703]));
Q_ASSIGN U31072 ( .B(clk), .A(\g.we_clk [1702]));
Q_ASSIGN U31073 ( .B(clk), .A(\g.we_clk [1701]));
Q_ASSIGN U31074 ( .B(clk), .A(\g.we_clk [1700]));
Q_ASSIGN U31075 ( .B(clk), .A(\g.we_clk [1699]));
Q_ASSIGN U31076 ( .B(clk), .A(\g.we_clk [1698]));
Q_ASSIGN U31077 ( .B(clk), .A(\g.we_clk [1697]));
Q_ASSIGN U31078 ( .B(clk), .A(\g.we_clk [1696]));
Q_ASSIGN U31079 ( .B(clk), .A(\g.we_clk [1695]));
Q_ASSIGN U31080 ( .B(clk), .A(\g.we_clk [1694]));
Q_ASSIGN U31081 ( .B(clk), .A(\g.we_clk [1693]));
Q_ASSIGN U31082 ( .B(clk), .A(\g.we_clk [1692]));
Q_ASSIGN U31083 ( .B(clk), .A(\g.we_clk [1691]));
Q_ASSIGN U31084 ( .B(clk), .A(\g.we_clk [1690]));
Q_ASSIGN U31085 ( .B(clk), .A(\g.we_clk [1689]));
Q_ASSIGN U31086 ( .B(clk), .A(\g.we_clk [1688]));
Q_ASSIGN U31087 ( .B(clk), .A(\g.we_clk [1687]));
Q_ASSIGN U31088 ( .B(clk), .A(\g.we_clk [1686]));
Q_ASSIGN U31089 ( .B(clk), .A(\g.we_clk [1685]));
Q_ASSIGN U31090 ( .B(clk), .A(\g.we_clk [1684]));
Q_ASSIGN U31091 ( .B(clk), .A(\g.we_clk [1683]));
Q_ASSIGN U31092 ( .B(clk), .A(\g.we_clk [1682]));
Q_ASSIGN U31093 ( .B(clk), .A(\g.we_clk [1681]));
Q_ASSIGN U31094 ( .B(clk), .A(\g.we_clk [1680]));
Q_ASSIGN U31095 ( .B(clk), .A(\g.we_clk [1679]));
Q_ASSIGN U31096 ( .B(clk), .A(\g.we_clk [1678]));
Q_ASSIGN U31097 ( .B(clk), .A(\g.we_clk [1677]));
Q_ASSIGN U31098 ( .B(clk), .A(\g.we_clk [1676]));
Q_ASSIGN U31099 ( .B(clk), .A(\g.we_clk [1675]));
Q_ASSIGN U31100 ( .B(clk), .A(\g.we_clk [1674]));
Q_ASSIGN U31101 ( .B(clk), .A(\g.we_clk [1673]));
Q_ASSIGN U31102 ( .B(clk), .A(\g.we_clk [1672]));
Q_ASSIGN U31103 ( .B(clk), .A(\g.we_clk [1671]));
Q_ASSIGN U31104 ( .B(clk), .A(\g.we_clk [1670]));
Q_ASSIGN U31105 ( .B(clk), .A(\g.we_clk [1669]));
Q_ASSIGN U31106 ( .B(clk), .A(\g.we_clk [1668]));
Q_ASSIGN U31107 ( .B(clk), .A(\g.we_clk [1667]));
Q_ASSIGN U31108 ( .B(clk), .A(\g.we_clk [1666]));
Q_ASSIGN U31109 ( .B(clk), .A(\g.we_clk [1665]));
Q_ASSIGN U31110 ( .B(clk), .A(\g.we_clk [1664]));
Q_ASSIGN U31111 ( .B(clk), .A(\g.we_clk [1663]));
Q_ASSIGN U31112 ( .B(clk), .A(\g.we_clk [1662]));
Q_ASSIGN U31113 ( .B(clk), .A(\g.we_clk [1661]));
Q_ASSIGN U31114 ( .B(clk), .A(\g.we_clk [1660]));
Q_ASSIGN U31115 ( .B(clk), .A(\g.we_clk [1659]));
Q_ASSIGN U31116 ( .B(clk), .A(\g.we_clk [1658]));
Q_ASSIGN U31117 ( .B(clk), .A(\g.we_clk [1657]));
Q_ASSIGN U31118 ( .B(clk), .A(\g.we_clk [1656]));
Q_ASSIGN U31119 ( .B(clk), .A(\g.we_clk [1655]));
Q_ASSIGN U31120 ( .B(clk), .A(\g.we_clk [1654]));
Q_ASSIGN U31121 ( .B(clk), .A(\g.we_clk [1653]));
Q_ASSIGN U31122 ( .B(clk), .A(\g.we_clk [1652]));
Q_ASSIGN U31123 ( .B(clk), .A(\g.we_clk [1651]));
Q_ASSIGN U31124 ( .B(clk), .A(\g.we_clk [1650]));
Q_ASSIGN U31125 ( .B(clk), .A(\g.we_clk [1649]));
Q_ASSIGN U31126 ( .B(clk), .A(\g.we_clk [1648]));
Q_ASSIGN U31127 ( .B(clk), .A(\g.we_clk [1647]));
Q_ASSIGN U31128 ( .B(clk), .A(\g.we_clk [1646]));
Q_ASSIGN U31129 ( .B(clk), .A(\g.we_clk [1645]));
Q_ASSIGN U31130 ( .B(clk), .A(\g.we_clk [1644]));
Q_ASSIGN U31131 ( .B(clk), .A(\g.we_clk [1643]));
Q_ASSIGN U31132 ( .B(clk), .A(\g.we_clk [1642]));
Q_ASSIGN U31133 ( .B(clk), .A(\g.we_clk [1641]));
Q_ASSIGN U31134 ( .B(clk), .A(\g.we_clk [1640]));
Q_ASSIGN U31135 ( .B(clk), .A(\g.we_clk [1639]));
Q_ASSIGN U31136 ( .B(clk), .A(\g.we_clk [1638]));
Q_ASSIGN U31137 ( .B(clk), .A(\g.we_clk [1637]));
Q_ASSIGN U31138 ( .B(clk), .A(\g.we_clk [1636]));
Q_ASSIGN U31139 ( .B(clk), .A(\g.we_clk [1635]));
Q_ASSIGN U31140 ( .B(clk), .A(\g.we_clk [1634]));
Q_ASSIGN U31141 ( .B(clk), .A(\g.we_clk [1633]));
Q_ASSIGN U31142 ( .B(clk), .A(\g.we_clk [1632]));
Q_ASSIGN U31143 ( .B(clk), .A(\g.we_clk [1631]));
Q_ASSIGN U31144 ( .B(clk), .A(\g.we_clk [1630]));
Q_ASSIGN U31145 ( .B(clk), .A(\g.we_clk [1629]));
Q_ASSIGN U31146 ( .B(clk), .A(\g.we_clk [1628]));
Q_ASSIGN U31147 ( .B(clk), .A(\g.we_clk [1627]));
Q_ASSIGN U31148 ( .B(clk), .A(\g.we_clk [1626]));
Q_ASSIGN U31149 ( .B(clk), .A(\g.we_clk [1625]));
Q_ASSIGN U31150 ( .B(clk), .A(\g.we_clk [1624]));
Q_ASSIGN U31151 ( .B(clk), .A(\g.we_clk [1623]));
Q_ASSIGN U31152 ( .B(clk), .A(\g.we_clk [1622]));
Q_ASSIGN U31153 ( .B(clk), .A(\g.we_clk [1621]));
Q_ASSIGN U31154 ( .B(clk), .A(\g.we_clk [1620]));
Q_ASSIGN U31155 ( .B(clk), .A(\g.we_clk [1619]));
Q_ASSIGN U31156 ( .B(clk), .A(\g.we_clk [1618]));
Q_ASSIGN U31157 ( .B(clk), .A(\g.we_clk [1617]));
Q_ASSIGN U31158 ( .B(clk), .A(\g.we_clk [1616]));
Q_ASSIGN U31159 ( .B(clk), .A(\g.we_clk [1615]));
Q_ASSIGN U31160 ( .B(clk), .A(\g.we_clk [1614]));
Q_ASSIGN U31161 ( .B(clk), .A(\g.we_clk [1613]));
Q_ASSIGN U31162 ( .B(clk), .A(\g.we_clk [1612]));
Q_ASSIGN U31163 ( .B(clk), .A(\g.we_clk [1611]));
Q_ASSIGN U31164 ( .B(clk), .A(\g.we_clk [1610]));
Q_ASSIGN U31165 ( .B(clk), .A(\g.we_clk [1609]));
Q_ASSIGN U31166 ( .B(clk), .A(\g.we_clk [1608]));
Q_ASSIGN U31167 ( .B(clk), .A(\g.we_clk [1607]));
Q_ASSIGN U31168 ( .B(clk), .A(\g.we_clk [1606]));
Q_ASSIGN U31169 ( .B(clk), .A(\g.we_clk [1605]));
Q_ASSIGN U31170 ( .B(clk), .A(\g.we_clk [1604]));
Q_ASSIGN U31171 ( .B(clk), .A(\g.we_clk [1603]));
Q_ASSIGN U31172 ( .B(clk), .A(\g.we_clk [1602]));
Q_ASSIGN U31173 ( .B(clk), .A(\g.we_clk [1601]));
Q_ASSIGN U31174 ( .B(clk), .A(\g.we_clk [1600]));
Q_ASSIGN U31175 ( .B(clk), .A(\g.we_clk [1599]));
Q_ASSIGN U31176 ( .B(clk), .A(\g.we_clk [1598]));
Q_ASSIGN U31177 ( .B(clk), .A(\g.we_clk [1597]));
Q_ASSIGN U31178 ( .B(clk), .A(\g.we_clk [1596]));
Q_ASSIGN U31179 ( .B(clk), .A(\g.we_clk [1595]));
Q_ASSIGN U31180 ( .B(clk), .A(\g.we_clk [1594]));
Q_ASSIGN U31181 ( .B(clk), .A(\g.we_clk [1593]));
Q_ASSIGN U31182 ( .B(clk), .A(\g.we_clk [1592]));
Q_ASSIGN U31183 ( .B(clk), .A(\g.we_clk [1591]));
Q_ASSIGN U31184 ( .B(clk), .A(\g.we_clk [1590]));
Q_ASSIGN U31185 ( .B(clk), .A(\g.we_clk [1589]));
Q_ASSIGN U31186 ( .B(clk), .A(\g.we_clk [1588]));
Q_ASSIGN U31187 ( .B(clk), .A(\g.we_clk [1587]));
Q_ASSIGN U31188 ( .B(clk), .A(\g.we_clk [1586]));
Q_ASSIGN U31189 ( .B(clk), .A(\g.we_clk [1585]));
Q_ASSIGN U31190 ( .B(clk), .A(\g.we_clk [1584]));
Q_ASSIGN U31191 ( .B(clk), .A(\g.we_clk [1583]));
Q_ASSIGN U31192 ( .B(clk), .A(\g.we_clk [1582]));
Q_ASSIGN U31193 ( .B(clk), .A(\g.we_clk [1581]));
Q_ASSIGN U31194 ( .B(clk), .A(\g.we_clk [1580]));
Q_ASSIGN U31195 ( .B(clk), .A(\g.we_clk [1579]));
Q_ASSIGN U31196 ( .B(clk), .A(\g.we_clk [1578]));
Q_ASSIGN U31197 ( .B(clk), .A(\g.we_clk [1577]));
Q_ASSIGN U31198 ( .B(clk), .A(\g.we_clk [1576]));
Q_ASSIGN U31199 ( .B(clk), .A(\g.we_clk [1575]));
Q_ASSIGN U31200 ( .B(clk), .A(\g.we_clk [1574]));
Q_ASSIGN U31201 ( .B(clk), .A(\g.we_clk [1573]));
Q_ASSIGN U31202 ( .B(clk), .A(\g.we_clk [1572]));
Q_ASSIGN U31203 ( .B(clk), .A(\g.we_clk [1571]));
Q_ASSIGN U31204 ( .B(clk), .A(\g.we_clk [1570]));
Q_ASSIGN U31205 ( .B(clk), .A(\g.we_clk [1569]));
Q_ASSIGN U31206 ( .B(clk), .A(\g.we_clk [1568]));
Q_ASSIGN U31207 ( .B(clk), .A(\g.we_clk [1567]));
Q_ASSIGN U31208 ( .B(clk), .A(\g.we_clk [1566]));
Q_ASSIGN U31209 ( .B(clk), .A(\g.we_clk [1565]));
Q_ASSIGN U31210 ( .B(clk), .A(\g.we_clk [1564]));
Q_ASSIGN U31211 ( .B(clk), .A(\g.we_clk [1563]));
Q_ASSIGN U31212 ( .B(clk), .A(\g.we_clk [1562]));
Q_ASSIGN U31213 ( .B(clk), .A(\g.we_clk [1561]));
Q_ASSIGN U31214 ( .B(clk), .A(\g.we_clk [1560]));
Q_ASSIGN U31215 ( .B(clk), .A(\g.we_clk [1559]));
Q_ASSIGN U31216 ( .B(clk), .A(\g.we_clk [1558]));
Q_ASSIGN U31217 ( .B(clk), .A(\g.we_clk [1557]));
Q_ASSIGN U31218 ( .B(clk), .A(\g.we_clk [1556]));
Q_ASSIGN U31219 ( .B(clk), .A(\g.we_clk [1555]));
Q_ASSIGN U31220 ( .B(clk), .A(\g.we_clk [1554]));
Q_ASSIGN U31221 ( .B(clk), .A(\g.we_clk [1553]));
Q_ASSIGN U31222 ( .B(clk), .A(\g.we_clk [1552]));
Q_ASSIGN U31223 ( .B(clk), .A(\g.we_clk [1551]));
Q_ASSIGN U31224 ( .B(clk), .A(\g.we_clk [1550]));
Q_ASSIGN U31225 ( .B(clk), .A(\g.we_clk [1549]));
Q_ASSIGN U31226 ( .B(clk), .A(\g.we_clk [1548]));
Q_ASSIGN U31227 ( .B(clk), .A(\g.we_clk [1547]));
Q_ASSIGN U31228 ( .B(clk), .A(\g.we_clk [1546]));
Q_ASSIGN U31229 ( .B(clk), .A(\g.we_clk [1545]));
Q_ASSIGN U31230 ( .B(clk), .A(\g.we_clk [1544]));
Q_ASSIGN U31231 ( .B(clk), .A(\g.we_clk [1543]));
Q_ASSIGN U31232 ( .B(clk), .A(\g.we_clk [1542]));
Q_ASSIGN U31233 ( .B(clk), .A(\g.we_clk [1541]));
Q_ASSIGN U31234 ( .B(clk), .A(\g.we_clk [1540]));
Q_ASSIGN U31235 ( .B(clk), .A(\g.we_clk [1539]));
Q_ASSIGN U31236 ( .B(clk), .A(\g.we_clk [1538]));
Q_ASSIGN U31237 ( .B(clk), .A(\g.we_clk [1537]));
Q_ASSIGN U31238 ( .B(clk), .A(\g.we_clk [1536]));
Q_ASSIGN U31239 ( .B(clk), .A(\g.we_clk [1535]));
Q_ASSIGN U31240 ( .B(clk), .A(\g.we_clk [1534]));
Q_ASSIGN U31241 ( .B(clk), .A(\g.we_clk [1533]));
Q_ASSIGN U31242 ( .B(clk), .A(\g.we_clk [1532]));
Q_ASSIGN U31243 ( .B(clk), .A(\g.we_clk [1531]));
Q_ASSIGN U31244 ( .B(clk), .A(\g.we_clk [1530]));
Q_ASSIGN U31245 ( .B(clk), .A(\g.we_clk [1529]));
Q_ASSIGN U31246 ( .B(clk), .A(\g.we_clk [1528]));
Q_ASSIGN U31247 ( .B(clk), .A(\g.we_clk [1527]));
Q_ASSIGN U31248 ( .B(clk), .A(\g.we_clk [1526]));
Q_ASSIGN U31249 ( .B(clk), .A(\g.we_clk [1525]));
Q_ASSIGN U31250 ( .B(clk), .A(\g.we_clk [1524]));
Q_ASSIGN U31251 ( .B(clk), .A(\g.we_clk [1523]));
Q_ASSIGN U31252 ( .B(clk), .A(\g.we_clk [1522]));
Q_ASSIGN U31253 ( .B(clk), .A(\g.we_clk [1521]));
Q_ASSIGN U31254 ( .B(clk), .A(\g.we_clk [1520]));
Q_ASSIGN U31255 ( .B(clk), .A(\g.we_clk [1519]));
Q_ASSIGN U31256 ( .B(clk), .A(\g.we_clk [1518]));
Q_ASSIGN U31257 ( .B(clk), .A(\g.we_clk [1517]));
Q_ASSIGN U31258 ( .B(clk), .A(\g.we_clk [1516]));
Q_ASSIGN U31259 ( .B(clk), .A(\g.we_clk [1515]));
Q_ASSIGN U31260 ( .B(clk), .A(\g.we_clk [1514]));
Q_ASSIGN U31261 ( .B(clk), .A(\g.we_clk [1513]));
Q_ASSIGN U31262 ( .B(clk), .A(\g.we_clk [1512]));
Q_ASSIGN U31263 ( .B(clk), .A(\g.we_clk [1511]));
Q_ASSIGN U31264 ( .B(clk), .A(\g.we_clk [1510]));
Q_ASSIGN U31265 ( .B(clk), .A(\g.we_clk [1509]));
Q_ASSIGN U31266 ( .B(clk), .A(\g.we_clk [1508]));
Q_ASSIGN U31267 ( .B(clk), .A(\g.we_clk [1507]));
Q_ASSIGN U31268 ( .B(clk), .A(\g.we_clk [1506]));
Q_ASSIGN U31269 ( .B(clk), .A(\g.we_clk [1505]));
Q_ASSIGN U31270 ( .B(clk), .A(\g.we_clk [1504]));
Q_ASSIGN U31271 ( .B(clk), .A(\g.we_clk [1503]));
Q_ASSIGN U31272 ( .B(clk), .A(\g.we_clk [1502]));
Q_ASSIGN U31273 ( .B(clk), .A(\g.we_clk [1501]));
Q_ASSIGN U31274 ( .B(clk), .A(\g.we_clk [1500]));
Q_ASSIGN U31275 ( .B(clk), .A(\g.we_clk [1499]));
Q_ASSIGN U31276 ( .B(clk), .A(\g.we_clk [1498]));
Q_ASSIGN U31277 ( .B(clk), .A(\g.we_clk [1497]));
Q_ASSIGN U31278 ( .B(clk), .A(\g.we_clk [1496]));
Q_ASSIGN U31279 ( .B(clk), .A(\g.we_clk [1495]));
Q_ASSIGN U31280 ( .B(clk), .A(\g.we_clk [1494]));
Q_ASSIGN U31281 ( .B(clk), .A(\g.we_clk [1493]));
Q_ASSIGN U31282 ( .B(clk), .A(\g.we_clk [1492]));
Q_ASSIGN U31283 ( .B(clk), .A(\g.we_clk [1491]));
Q_ASSIGN U31284 ( .B(clk), .A(\g.we_clk [1490]));
Q_ASSIGN U31285 ( .B(clk), .A(\g.we_clk [1489]));
Q_ASSIGN U31286 ( .B(clk), .A(\g.we_clk [1488]));
Q_ASSIGN U31287 ( .B(clk), .A(\g.we_clk [1487]));
Q_ASSIGN U31288 ( .B(clk), .A(\g.we_clk [1486]));
Q_ASSIGN U31289 ( .B(clk), .A(\g.we_clk [1485]));
Q_ASSIGN U31290 ( .B(clk), .A(\g.we_clk [1484]));
Q_ASSIGN U31291 ( .B(clk), .A(\g.we_clk [1483]));
Q_ASSIGN U31292 ( .B(clk), .A(\g.we_clk [1482]));
Q_ASSIGN U31293 ( .B(clk), .A(\g.we_clk [1481]));
Q_ASSIGN U31294 ( .B(clk), .A(\g.we_clk [1480]));
Q_ASSIGN U31295 ( .B(clk), .A(\g.we_clk [1479]));
Q_ASSIGN U31296 ( .B(clk), .A(\g.we_clk [1478]));
Q_ASSIGN U31297 ( .B(clk), .A(\g.we_clk [1477]));
Q_ASSIGN U31298 ( .B(clk), .A(\g.we_clk [1476]));
Q_ASSIGN U31299 ( .B(clk), .A(\g.we_clk [1475]));
Q_ASSIGN U31300 ( .B(clk), .A(\g.we_clk [1474]));
Q_ASSIGN U31301 ( .B(clk), .A(\g.we_clk [1473]));
Q_ASSIGN U31302 ( .B(clk), .A(\g.we_clk [1472]));
Q_ASSIGN U31303 ( .B(clk), .A(\g.we_clk [1471]));
Q_ASSIGN U31304 ( .B(clk), .A(\g.we_clk [1470]));
Q_ASSIGN U31305 ( .B(clk), .A(\g.we_clk [1469]));
Q_ASSIGN U31306 ( .B(clk), .A(\g.we_clk [1468]));
Q_ASSIGN U31307 ( .B(clk), .A(\g.we_clk [1467]));
Q_ASSIGN U31308 ( .B(clk), .A(\g.we_clk [1466]));
Q_ASSIGN U31309 ( .B(clk), .A(\g.we_clk [1465]));
Q_ASSIGN U31310 ( .B(clk), .A(\g.we_clk [1464]));
Q_ASSIGN U31311 ( .B(clk), .A(\g.we_clk [1463]));
Q_ASSIGN U31312 ( .B(clk), .A(\g.we_clk [1462]));
Q_ASSIGN U31313 ( .B(clk), .A(\g.we_clk [1461]));
Q_ASSIGN U31314 ( .B(clk), .A(\g.we_clk [1460]));
Q_ASSIGN U31315 ( .B(clk), .A(\g.we_clk [1459]));
Q_ASSIGN U31316 ( .B(clk), .A(\g.we_clk [1458]));
Q_ASSIGN U31317 ( .B(clk), .A(\g.we_clk [1457]));
Q_ASSIGN U31318 ( .B(clk), .A(\g.we_clk [1456]));
Q_ASSIGN U31319 ( .B(clk), .A(\g.we_clk [1455]));
Q_ASSIGN U31320 ( .B(clk), .A(\g.we_clk [1454]));
Q_ASSIGN U31321 ( .B(clk), .A(\g.we_clk [1453]));
Q_ASSIGN U31322 ( .B(clk), .A(\g.we_clk [1452]));
Q_ASSIGN U31323 ( .B(clk), .A(\g.we_clk [1451]));
Q_ASSIGN U31324 ( .B(clk), .A(\g.we_clk [1450]));
Q_ASSIGN U31325 ( .B(clk), .A(\g.we_clk [1449]));
Q_ASSIGN U31326 ( .B(clk), .A(\g.we_clk [1448]));
Q_ASSIGN U31327 ( .B(clk), .A(\g.we_clk [1447]));
Q_ASSIGN U31328 ( .B(clk), .A(\g.we_clk [1446]));
Q_ASSIGN U31329 ( .B(clk), .A(\g.we_clk [1445]));
Q_ASSIGN U31330 ( .B(clk), .A(\g.we_clk [1444]));
Q_ASSIGN U31331 ( .B(clk), .A(\g.we_clk [1443]));
Q_ASSIGN U31332 ( .B(clk), .A(\g.we_clk [1442]));
Q_ASSIGN U31333 ( .B(clk), .A(\g.we_clk [1441]));
Q_ASSIGN U31334 ( .B(clk), .A(\g.we_clk [1440]));
Q_ASSIGN U31335 ( .B(clk), .A(\g.we_clk [1439]));
Q_ASSIGN U31336 ( .B(clk), .A(\g.we_clk [1438]));
Q_ASSIGN U31337 ( .B(clk), .A(\g.we_clk [1437]));
Q_ASSIGN U31338 ( .B(clk), .A(\g.we_clk [1436]));
Q_ASSIGN U31339 ( .B(clk), .A(\g.we_clk [1435]));
Q_ASSIGN U31340 ( .B(clk), .A(\g.we_clk [1434]));
Q_ASSIGN U31341 ( .B(clk), .A(\g.we_clk [1433]));
Q_ASSIGN U31342 ( .B(clk), .A(\g.we_clk [1432]));
Q_ASSIGN U31343 ( .B(clk), .A(\g.we_clk [1431]));
Q_ASSIGN U31344 ( .B(clk), .A(\g.we_clk [1430]));
Q_ASSIGN U31345 ( .B(clk), .A(\g.we_clk [1429]));
Q_ASSIGN U31346 ( .B(clk), .A(\g.we_clk [1428]));
Q_ASSIGN U31347 ( .B(clk), .A(\g.we_clk [1427]));
Q_ASSIGN U31348 ( .B(clk), .A(\g.we_clk [1426]));
Q_ASSIGN U31349 ( .B(clk), .A(\g.we_clk [1425]));
Q_ASSIGN U31350 ( .B(clk), .A(\g.we_clk [1424]));
Q_ASSIGN U31351 ( .B(clk), .A(\g.we_clk [1423]));
Q_ASSIGN U31352 ( .B(clk), .A(\g.we_clk [1422]));
Q_ASSIGN U31353 ( .B(clk), .A(\g.we_clk [1421]));
Q_ASSIGN U31354 ( .B(clk), .A(\g.we_clk [1420]));
Q_ASSIGN U31355 ( .B(clk), .A(\g.we_clk [1419]));
Q_ASSIGN U31356 ( .B(clk), .A(\g.we_clk [1418]));
Q_ASSIGN U31357 ( .B(clk), .A(\g.we_clk [1417]));
Q_ASSIGN U31358 ( .B(clk), .A(\g.we_clk [1416]));
Q_ASSIGN U31359 ( .B(clk), .A(\g.we_clk [1415]));
Q_ASSIGN U31360 ( .B(clk), .A(\g.we_clk [1414]));
Q_ASSIGN U31361 ( .B(clk), .A(\g.we_clk [1413]));
Q_ASSIGN U31362 ( .B(clk), .A(\g.we_clk [1412]));
Q_ASSIGN U31363 ( .B(clk), .A(\g.we_clk [1411]));
Q_ASSIGN U31364 ( .B(clk), .A(\g.we_clk [1410]));
Q_ASSIGN U31365 ( .B(clk), .A(\g.we_clk [1409]));
Q_ASSIGN U31366 ( .B(clk), .A(\g.we_clk [1408]));
Q_ASSIGN U31367 ( .B(clk), .A(\g.we_clk [1407]));
Q_ASSIGN U31368 ( .B(clk), .A(\g.we_clk [1406]));
Q_ASSIGN U31369 ( .B(clk), .A(\g.we_clk [1405]));
Q_ASSIGN U31370 ( .B(clk), .A(\g.we_clk [1404]));
Q_ASSIGN U31371 ( .B(clk), .A(\g.we_clk [1403]));
Q_ASSIGN U31372 ( .B(clk), .A(\g.we_clk [1402]));
Q_ASSIGN U31373 ( .B(clk), .A(\g.we_clk [1401]));
Q_ASSIGN U31374 ( .B(clk), .A(\g.we_clk [1400]));
Q_ASSIGN U31375 ( .B(clk), .A(\g.we_clk [1399]));
Q_ASSIGN U31376 ( .B(clk), .A(\g.we_clk [1398]));
Q_ASSIGN U31377 ( .B(clk), .A(\g.we_clk [1397]));
Q_ASSIGN U31378 ( .B(clk), .A(\g.we_clk [1396]));
Q_ASSIGN U31379 ( .B(clk), .A(\g.we_clk [1395]));
Q_ASSIGN U31380 ( .B(clk), .A(\g.we_clk [1394]));
Q_ASSIGN U31381 ( .B(clk), .A(\g.we_clk [1393]));
Q_ASSIGN U31382 ( .B(clk), .A(\g.we_clk [1392]));
Q_ASSIGN U31383 ( .B(clk), .A(\g.we_clk [1391]));
Q_ASSIGN U31384 ( .B(clk), .A(\g.we_clk [1390]));
Q_ASSIGN U31385 ( .B(clk), .A(\g.we_clk [1389]));
Q_ASSIGN U31386 ( .B(clk), .A(\g.we_clk [1388]));
Q_ASSIGN U31387 ( .B(clk), .A(\g.we_clk [1387]));
Q_ASSIGN U31388 ( .B(clk), .A(\g.we_clk [1386]));
Q_ASSIGN U31389 ( .B(clk), .A(\g.we_clk [1385]));
Q_ASSIGN U31390 ( .B(clk), .A(\g.we_clk [1384]));
Q_ASSIGN U31391 ( .B(clk), .A(\g.we_clk [1383]));
Q_ASSIGN U31392 ( .B(clk), .A(\g.we_clk [1382]));
Q_ASSIGN U31393 ( .B(clk), .A(\g.we_clk [1381]));
Q_ASSIGN U31394 ( .B(clk), .A(\g.we_clk [1380]));
Q_ASSIGN U31395 ( .B(clk), .A(\g.we_clk [1379]));
Q_ASSIGN U31396 ( .B(clk), .A(\g.we_clk [1378]));
Q_ASSIGN U31397 ( .B(clk), .A(\g.we_clk [1377]));
Q_ASSIGN U31398 ( .B(clk), .A(\g.we_clk [1376]));
Q_ASSIGN U31399 ( .B(clk), .A(\g.we_clk [1375]));
Q_ASSIGN U31400 ( .B(clk), .A(\g.we_clk [1374]));
Q_ASSIGN U31401 ( .B(clk), .A(\g.we_clk [1373]));
Q_ASSIGN U31402 ( .B(clk), .A(\g.we_clk [1372]));
Q_ASSIGN U31403 ( .B(clk), .A(\g.we_clk [1371]));
Q_ASSIGN U31404 ( .B(clk), .A(\g.we_clk [1370]));
Q_ASSIGN U31405 ( .B(clk), .A(\g.we_clk [1369]));
Q_ASSIGN U31406 ( .B(clk), .A(\g.we_clk [1368]));
Q_ASSIGN U31407 ( .B(clk), .A(\g.we_clk [1367]));
Q_ASSIGN U31408 ( .B(clk), .A(\g.we_clk [1366]));
Q_ASSIGN U31409 ( .B(clk), .A(\g.we_clk [1365]));
Q_ASSIGN U31410 ( .B(clk), .A(\g.we_clk [1364]));
Q_ASSIGN U31411 ( .B(clk), .A(\g.we_clk [1363]));
Q_ASSIGN U31412 ( .B(clk), .A(\g.we_clk [1362]));
Q_ASSIGN U31413 ( .B(clk), .A(\g.we_clk [1361]));
Q_ASSIGN U31414 ( .B(clk), .A(\g.we_clk [1360]));
Q_ASSIGN U31415 ( .B(clk), .A(\g.we_clk [1359]));
Q_ASSIGN U31416 ( .B(clk), .A(\g.we_clk [1358]));
Q_ASSIGN U31417 ( .B(clk), .A(\g.we_clk [1357]));
Q_ASSIGN U31418 ( .B(clk), .A(\g.we_clk [1356]));
Q_ASSIGN U31419 ( .B(clk), .A(\g.we_clk [1355]));
Q_ASSIGN U31420 ( .B(clk), .A(\g.we_clk [1354]));
Q_ASSIGN U31421 ( .B(clk), .A(\g.we_clk [1353]));
Q_ASSIGN U31422 ( .B(clk), .A(\g.we_clk [1352]));
Q_ASSIGN U31423 ( .B(clk), .A(\g.we_clk [1351]));
Q_ASSIGN U31424 ( .B(clk), .A(\g.we_clk [1350]));
Q_ASSIGN U31425 ( .B(clk), .A(\g.we_clk [1349]));
Q_ASSIGN U31426 ( .B(clk), .A(\g.we_clk [1348]));
Q_ASSIGN U31427 ( .B(clk), .A(\g.we_clk [1347]));
Q_ASSIGN U31428 ( .B(clk), .A(\g.we_clk [1346]));
Q_ASSIGN U31429 ( .B(clk), .A(\g.we_clk [1345]));
Q_ASSIGN U31430 ( .B(clk), .A(\g.we_clk [1344]));
Q_ASSIGN U31431 ( .B(clk), .A(\g.we_clk [1343]));
Q_ASSIGN U31432 ( .B(clk), .A(\g.we_clk [1342]));
Q_ASSIGN U31433 ( .B(clk), .A(\g.we_clk [1341]));
Q_ASSIGN U31434 ( .B(clk), .A(\g.we_clk [1340]));
Q_ASSIGN U31435 ( .B(clk), .A(\g.we_clk [1339]));
Q_ASSIGN U31436 ( .B(clk), .A(\g.we_clk [1338]));
Q_ASSIGN U31437 ( .B(clk), .A(\g.we_clk [1337]));
Q_ASSIGN U31438 ( .B(clk), .A(\g.we_clk [1336]));
Q_ASSIGN U31439 ( .B(clk), .A(\g.we_clk [1335]));
Q_ASSIGN U31440 ( .B(clk), .A(\g.we_clk [1334]));
Q_ASSIGN U31441 ( .B(clk), .A(\g.we_clk [1333]));
Q_ASSIGN U31442 ( .B(clk), .A(\g.we_clk [1332]));
Q_ASSIGN U31443 ( .B(clk), .A(\g.we_clk [1331]));
Q_ASSIGN U31444 ( .B(clk), .A(\g.we_clk [1330]));
Q_ASSIGN U31445 ( .B(clk), .A(\g.we_clk [1329]));
Q_ASSIGN U31446 ( .B(clk), .A(\g.we_clk [1328]));
Q_ASSIGN U31447 ( .B(clk), .A(\g.we_clk [1327]));
Q_ASSIGN U31448 ( .B(clk), .A(\g.we_clk [1326]));
Q_ASSIGN U31449 ( .B(clk), .A(\g.we_clk [1325]));
Q_ASSIGN U31450 ( .B(clk), .A(\g.we_clk [1324]));
Q_ASSIGN U31451 ( .B(clk), .A(\g.we_clk [1323]));
Q_ASSIGN U31452 ( .B(clk), .A(\g.we_clk [1322]));
Q_ASSIGN U31453 ( .B(clk), .A(\g.we_clk [1321]));
Q_ASSIGN U31454 ( .B(clk), .A(\g.we_clk [1320]));
Q_ASSIGN U31455 ( .B(clk), .A(\g.we_clk [1319]));
Q_ASSIGN U31456 ( .B(clk), .A(\g.we_clk [1318]));
Q_ASSIGN U31457 ( .B(clk), .A(\g.we_clk [1317]));
Q_ASSIGN U31458 ( .B(clk), .A(\g.we_clk [1316]));
Q_ASSIGN U31459 ( .B(clk), .A(\g.we_clk [1315]));
Q_ASSIGN U31460 ( .B(clk), .A(\g.we_clk [1314]));
Q_ASSIGN U31461 ( .B(clk), .A(\g.we_clk [1313]));
Q_ASSIGN U31462 ( .B(clk), .A(\g.we_clk [1312]));
Q_ASSIGN U31463 ( .B(clk), .A(\g.we_clk [1311]));
Q_ASSIGN U31464 ( .B(clk), .A(\g.we_clk [1310]));
Q_ASSIGN U31465 ( .B(clk), .A(\g.we_clk [1309]));
Q_ASSIGN U31466 ( .B(clk), .A(\g.we_clk [1308]));
Q_ASSIGN U31467 ( .B(clk), .A(\g.we_clk [1307]));
Q_ASSIGN U31468 ( .B(clk), .A(\g.we_clk [1306]));
Q_ASSIGN U31469 ( .B(clk), .A(\g.we_clk [1305]));
Q_ASSIGN U31470 ( .B(clk), .A(\g.we_clk [1304]));
Q_ASSIGN U31471 ( .B(clk), .A(\g.we_clk [1303]));
Q_ASSIGN U31472 ( .B(clk), .A(\g.we_clk [1302]));
Q_ASSIGN U31473 ( .B(clk), .A(\g.we_clk [1301]));
Q_ASSIGN U31474 ( .B(clk), .A(\g.we_clk [1300]));
Q_ASSIGN U31475 ( .B(clk), .A(\g.we_clk [1299]));
Q_ASSIGN U31476 ( .B(clk), .A(\g.we_clk [1298]));
Q_ASSIGN U31477 ( .B(clk), .A(\g.we_clk [1297]));
Q_ASSIGN U31478 ( .B(clk), .A(\g.we_clk [1296]));
Q_ASSIGN U31479 ( .B(clk), .A(\g.we_clk [1295]));
Q_ASSIGN U31480 ( .B(clk), .A(\g.we_clk [1294]));
Q_ASSIGN U31481 ( .B(clk), .A(\g.we_clk [1293]));
Q_ASSIGN U31482 ( .B(clk), .A(\g.we_clk [1292]));
Q_ASSIGN U31483 ( .B(clk), .A(\g.we_clk [1291]));
Q_ASSIGN U31484 ( .B(clk), .A(\g.we_clk [1290]));
Q_ASSIGN U31485 ( .B(clk), .A(\g.we_clk [1289]));
Q_ASSIGN U31486 ( .B(clk), .A(\g.we_clk [1288]));
Q_ASSIGN U31487 ( .B(clk), .A(\g.we_clk [1287]));
Q_ASSIGN U31488 ( .B(clk), .A(\g.we_clk [1286]));
Q_ASSIGN U31489 ( .B(clk), .A(\g.we_clk [1285]));
Q_ASSIGN U31490 ( .B(clk), .A(\g.we_clk [1284]));
Q_ASSIGN U31491 ( .B(clk), .A(\g.we_clk [1283]));
Q_ASSIGN U31492 ( .B(clk), .A(\g.we_clk [1282]));
Q_ASSIGN U31493 ( .B(clk), .A(\g.we_clk [1281]));
Q_ASSIGN U31494 ( .B(clk), .A(\g.we_clk [1280]));
Q_ASSIGN U31495 ( .B(clk), .A(\g.we_clk [1279]));
Q_ASSIGN U31496 ( .B(clk), .A(\g.we_clk [1278]));
Q_ASSIGN U31497 ( .B(clk), .A(\g.we_clk [1277]));
Q_ASSIGN U31498 ( .B(clk), .A(\g.we_clk [1276]));
Q_ASSIGN U31499 ( .B(clk), .A(\g.we_clk [1275]));
Q_ASSIGN U31500 ( .B(clk), .A(\g.we_clk [1274]));
Q_ASSIGN U31501 ( .B(clk), .A(\g.we_clk [1273]));
Q_ASSIGN U31502 ( .B(clk), .A(\g.we_clk [1272]));
Q_ASSIGN U31503 ( .B(clk), .A(\g.we_clk [1271]));
Q_ASSIGN U31504 ( .B(clk), .A(\g.we_clk [1270]));
Q_ASSIGN U31505 ( .B(clk), .A(\g.we_clk [1269]));
Q_ASSIGN U31506 ( .B(clk), .A(\g.we_clk [1268]));
Q_ASSIGN U31507 ( .B(clk), .A(\g.we_clk [1267]));
Q_ASSIGN U31508 ( .B(clk), .A(\g.we_clk [1266]));
Q_ASSIGN U31509 ( .B(clk), .A(\g.we_clk [1265]));
Q_ASSIGN U31510 ( .B(clk), .A(\g.we_clk [1264]));
Q_ASSIGN U31511 ( .B(clk), .A(\g.we_clk [1263]));
Q_ASSIGN U31512 ( .B(clk), .A(\g.we_clk [1262]));
Q_ASSIGN U31513 ( .B(clk), .A(\g.we_clk [1261]));
Q_ASSIGN U31514 ( .B(clk), .A(\g.we_clk [1260]));
Q_ASSIGN U31515 ( .B(clk), .A(\g.we_clk [1259]));
Q_ASSIGN U31516 ( .B(clk), .A(\g.we_clk [1258]));
Q_ASSIGN U31517 ( .B(clk), .A(\g.we_clk [1257]));
Q_ASSIGN U31518 ( .B(clk), .A(\g.we_clk [1256]));
Q_ASSIGN U31519 ( .B(clk), .A(\g.we_clk [1255]));
Q_ASSIGN U31520 ( .B(clk), .A(\g.we_clk [1254]));
Q_ASSIGN U31521 ( .B(clk), .A(\g.we_clk [1253]));
Q_ASSIGN U31522 ( .B(clk), .A(\g.we_clk [1252]));
Q_ASSIGN U31523 ( .B(clk), .A(\g.we_clk [1251]));
Q_ASSIGN U31524 ( .B(clk), .A(\g.we_clk [1250]));
Q_ASSIGN U31525 ( .B(clk), .A(\g.we_clk [1249]));
Q_ASSIGN U31526 ( .B(clk), .A(\g.we_clk [1248]));
Q_ASSIGN U31527 ( .B(clk), .A(\g.we_clk [1247]));
Q_ASSIGN U31528 ( .B(clk), .A(\g.we_clk [1246]));
Q_ASSIGN U31529 ( .B(clk), .A(\g.we_clk [1245]));
Q_ASSIGN U31530 ( .B(clk), .A(\g.we_clk [1244]));
Q_ASSIGN U31531 ( .B(clk), .A(\g.we_clk [1243]));
Q_ASSIGN U31532 ( .B(clk), .A(\g.we_clk [1242]));
Q_ASSIGN U31533 ( .B(clk), .A(\g.we_clk [1241]));
Q_ASSIGN U31534 ( .B(clk), .A(\g.we_clk [1240]));
Q_ASSIGN U31535 ( .B(clk), .A(\g.we_clk [1239]));
Q_ASSIGN U31536 ( .B(clk), .A(\g.we_clk [1238]));
Q_ASSIGN U31537 ( .B(clk), .A(\g.we_clk [1237]));
Q_ASSIGN U31538 ( .B(clk), .A(\g.we_clk [1236]));
Q_ASSIGN U31539 ( .B(clk), .A(\g.we_clk [1235]));
Q_ASSIGN U31540 ( .B(clk), .A(\g.we_clk [1234]));
Q_ASSIGN U31541 ( .B(clk), .A(\g.we_clk [1233]));
Q_ASSIGN U31542 ( .B(clk), .A(\g.we_clk [1232]));
Q_ASSIGN U31543 ( .B(clk), .A(\g.we_clk [1231]));
Q_ASSIGN U31544 ( .B(clk), .A(\g.we_clk [1230]));
Q_ASSIGN U31545 ( .B(clk), .A(\g.we_clk [1229]));
Q_ASSIGN U31546 ( .B(clk), .A(\g.we_clk [1228]));
Q_ASSIGN U31547 ( .B(clk), .A(\g.we_clk [1227]));
Q_ASSIGN U31548 ( .B(clk), .A(\g.we_clk [1226]));
Q_ASSIGN U31549 ( .B(clk), .A(\g.we_clk [1225]));
Q_ASSIGN U31550 ( .B(clk), .A(\g.we_clk [1224]));
Q_ASSIGN U31551 ( .B(clk), .A(\g.we_clk [1223]));
Q_ASSIGN U31552 ( .B(clk), .A(\g.we_clk [1222]));
Q_ASSIGN U31553 ( .B(clk), .A(\g.we_clk [1221]));
Q_ASSIGN U31554 ( .B(clk), .A(\g.we_clk [1220]));
Q_ASSIGN U31555 ( .B(clk), .A(\g.we_clk [1219]));
Q_ASSIGN U31556 ( .B(clk), .A(\g.we_clk [1218]));
Q_ASSIGN U31557 ( .B(clk), .A(\g.we_clk [1217]));
Q_ASSIGN U31558 ( .B(clk), .A(\g.we_clk [1216]));
Q_ASSIGN U31559 ( .B(clk), .A(\g.we_clk [1215]));
Q_ASSIGN U31560 ( .B(clk), .A(\g.we_clk [1214]));
Q_ASSIGN U31561 ( .B(clk), .A(\g.we_clk [1213]));
Q_ASSIGN U31562 ( .B(clk), .A(\g.we_clk [1212]));
Q_ASSIGN U31563 ( .B(clk), .A(\g.we_clk [1211]));
Q_ASSIGN U31564 ( .B(clk), .A(\g.we_clk [1210]));
Q_ASSIGN U31565 ( .B(clk), .A(\g.we_clk [1209]));
Q_ASSIGN U31566 ( .B(clk), .A(\g.we_clk [1208]));
Q_ASSIGN U31567 ( .B(clk), .A(\g.we_clk [1207]));
Q_ASSIGN U31568 ( .B(clk), .A(\g.we_clk [1206]));
Q_ASSIGN U31569 ( .B(clk), .A(\g.we_clk [1205]));
Q_ASSIGN U31570 ( .B(clk), .A(\g.we_clk [1204]));
Q_ASSIGN U31571 ( .B(clk), .A(\g.we_clk [1203]));
Q_ASSIGN U31572 ( .B(clk), .A(\g.we_clk [1202]));
Q_ASSIGN U31573 ( .B(clk), .A(\g.we_clk [1201]));
Q_ASSIGN U31574 ( .B(clk), .A(\g.we_clk [1200]));
Q_ASSIGN U31575 ( .B(clk), .A(\g.we_clk [1199]));
Q_ASSIGN U31576 ( .B(clk), .A(\g.we_clk [1198]));
Q_ASSIGN U31577 ( .B(clk), .A(\g.we_clk [1197]));
Q_ASSIGN U31578 ( .B(clk), .A(\g.we_clk [1196]));
Q_ASSIGN U31579 ( .B(clk), .A(\g.we_clk [1195]));
Q_ASSIGN U31580 ( .B(clk), .A(\g.we_clk [1194]));
Q_ASSIGN U31581 ( .B(clk), .A(\g.we_clk [1193]));
Q_ASSIGN U31582 ( .B(clk), .A(\g.we_clk [1192]));
Q_ASSIGN U31583 ( .B(clk), .A(\g.we_clk [1191]));
Q_ASSIGN U31584 ( .B(clk), .A(\g.we_clk [1190]));
Q_ASSIGN U31585 ( .B(clk), .A(\g.we_clk [1189]));
Q_ASSIGN U31586 ( .B(clk), .A(\g.we_clk [1188]));
Q_ASSIGN U31587 ( .B(clk), .A(\g.we_clk [1187]));
Q_ASSIGN U31588 ( .B(clk), .A(\g.we_clk [1186]));
Q_ASSIGN U31589 ( .B(clk), .A(\g.we_clk [1185]));
Q_ASSIGN U31590 ( .B(clk), .A(\g.we_clk [1184]));
Q_ASSIGN U31591 ( .B(clk), .A(\g.we_clk [1183]));
Q_ASSIGN U31592 ( .B(clk), .A(\g.we_clk [1182]));
Q_ASSIGN U31593 ( .B(clk), .A(\g.we_clk [1181]));
Q_ASSIGN U31594 ( .B(clk), .A(\g.we_clk [1180]));
Q_ASSIGN U31595 ( .B(clk), .A(\g.we_clk [1179]));
Q_ASSIGN U31596 ( .B(clk), .A(\g.we_clk [1178]));
Q_ASSIGN U31597 ( .B(clk), .A(\g.we_clk [1177]));
Q_ASSIGN U31598 ( .B(clk), .A(\g.we_clk [1176]));
Q_ASSIGN U31599 ( .B(clk), .A(\g.we_clk [1175]));
Q_ASSIGN U31600 ( .B(clk), .A(\g.we_clk [1174]));
Q_ASSIGN U31601 ( .B(clk), .A(\g.we_clk [1173]));
Q_ASSIGN U31602 ( .B(clk), .A(\g.we_clk [1172]));
Q_ASSIGN U31603 ( .B(clk), .A(\g.we_clk [1171]));
Q_ASSIGN U31604 ( .B(clk), .A(\g.we_clk [1170]));
Q_ASSIGN U31605 ( .B(clk), .A(\g.we_clk [1169]));
Q_ASSIGN U31606 ( .B(clk), .A(\g.we_clk [1168]));
Q_ASSIGN U31607 ( .B(clk), .A(\g.we_clk [1167]));
Q_ASSIGN U31608 ( .B(clk), .A(\g.we_clk [1166]));
Q_ASSIGN U31609 ( .B(clk), .A(\g.we_clk [1165]));
Q_ASSIGN U31610 ( .B(clk), .A(\g.we_clk [1164]));
Q_ASSIGN U31611 ( .B(clk), .A(\g.we_clk [1163]));
Q_ASSIGN U31612 ( .B(clk), .A(\g.we_clk [1162]));
Q_ASSIGN U31613 ( .B(clk), .A(\g.we_clk [1161]));
Q_ASSIGN U31614 ( .B(clk), .A(\g.we_clk [1160]));
Q_ASSIGN U31615 ( .B(clk), .A(\g.we_clk [1159]));
Q_ASSIGN U31616 ( .B(clk), .A(\g.we_clk [1158]));
Q_ASSIGN U31617 ( .B(clk), .A(\g.we_clk [1157]));
Q_ASSIGN U31618 ( .B(clk), .A(\g.we_clk [1156]));
Q_ASSIGN U31619 ( .B(clk), .A(\g.we_clk [1155]));
Q_ASSIGN U31620 ( .B(clk), .A(\g.we_clk [1154]));
Q_ASSIGN U31621 ( .B(clk), .A(\g.we_clk [1153]));
Q_ASSIGN U31622 ( .B(clk), .A(\g.we_clk [1152]));
Q_ASSIGN U31623 ( .B(clk), .A(\g.we_clk [1151]));
Q_ASSIGN U31624 ( .B(clk), .A(\g.we_clk [1150]));
Q_ASSIGN U31625 ( .B(clk), .A(\g.we_clk [1149]));
Q_ASSIGN U31626 ( .B(clk), .A(\g.we_clk [1148]));
Q_ASSIGN U31627 ( .B(clk), .A(\g.we_clk [1147]));
Q_ASSIGN U31628 ( .B(clk), .A(\g.we_clk [1146]));
Q_ASSIGN U31629 ( .B(clk), .A(\g.we_clk [1145]));
Q_ASSIGN U31630 ( .B(clk), .A(\g.we_clk [1144]));
Q_ASSIGN U31631 ( .B(clk), .A(\g.we_clk [1143]));
Q_ASSIGN U31632 ( .B(clk), .A(\g.we_clk [1142]));
Q_ASSIGN U31633 ( .B(clk), .A(\g.we_clk [1141]));
Q_ASSIGN U31634 ( .B(clk), .A(\g.we_clk [1140]));
Q_ASSIGN U31635 ( .B(clk), .A(\g.we_clk [1139]));
Q_ASSIGN U31636 ( .B(clk), .A(\g.we_clk [1138]));
Q_ASSIGN U31637 ( .B(clk), .A(\g.we_clk [1137]));
Q_ASSIGN U31638 ( .B(clk), .A(\g.we_clk [1136]));
Q_ASSIGN U31639 ( .B(clk), .A(\g.we_clk [1135]));
Q_ASSIGN U31640 ( .B(clk), .A(\g.we_clk [1134]));
Q_ASSIGN U31641 ( .B(clk), .A(\g.we_clk [1133]));
Q_ASSIGN U31642 ( .B(clk), .A(\g.we_clk [1132]));
Q_ASSIGN U31643 ( .B(clk), .A(\g.we_clk [1131]));
Q_ASSIGN U31644 ( .B(clk), .A(\g.we_clk [1130]));
Q_ASSIGN U31645 ( .B(clk), .A(\g.we_clk [1129]));
Q_ASSIGN U31646 ( .B(clk), .A(\g.we_clk [1128]));
Q_ASSIGN U31647 ( .B(clk), .A(\g.we_clk [1127]));
Q_ASSIGN U31648 ( .B(clk), .A(\g.we_clk [1126]));
Q_ASSIGN U31649 ( .B(clk), .A(\g.we_clk [1125]));
Q_ASSIGN U31650 ( .B(clk), .A(\g.we_clk [1124]));
Q_ASSIGN U31651 ( .B(clk), .A(\g.we_clk [1123]));
Q_ASSIGN U31652 ( .B(clk), .A(\g.we_clk [1122]));
Q_ASSIGN U31653 ( .B(clk), .A(\g.we_clk [1121]));
Q_ASSIGN U31654 ( .B(clk), .A(\g.we_clk [1120]));
Q_ASSIGN U31655 ( .B(clk), .A(\g.we_clk [1119]));
Q_ASSIGN U31656 ( .B(clk), .A(\g.we_clk [1118]));
Q_ASSIGN U31657 ( .B(clk), .A(\g.we_clk [1117]));
Q_ASSIGN U31658 ( .B(clk), .A(\g.we_clk [1116]));
Q_ASSIGN U31659 ( .B(clk), .A(\g.we_clk [1115]));
Q_ASSIGN U31660 ( .B(clk), .A(\g.we_clk [1114]));
Q_ASSIGN U31661 ( .B(clk), .A(\g.we_clk [1113]));
Q_ASSIGN U31662 ( .B(clk), .A(\g.we_clk [1112]));
Q_ASSIGN U31663 ( .B(clk), .A(\g.we_clk [1111]));
Q_ASSIGN U31664 ( .B(clk), .A(\g.we_clk [1110]));
Q_ASSIGN U31665 ( .B(clk), .A(\g.we_clk [1109]));
Q_ASSIGN U31666 ( .B(clk), .A(\g.we_clk [1108]));
Q_ASSIGN U31667 ( .B(clk), .A(\g.we_clk [1107]));
Q_ASSIGN U31668 ( .B(clk), .A(\g.we_clk [1106]));
Q_ASSIGN U31669 ( .B(clk), .A(\g.we_clk [1105]));
Q_ASSIGN U31670 ( .B(clk), .A(\g.we_clk [1104]));
Q_ASSIGN U31671 ( .B(clk), .A(\g.we_clk [1103]));
Q_ASSIGN U31672 ( .B(clk), .A(\g.we_clk [1102]));
Q_ASSIGN U31673 ( .B(clk), .A(\g.we_clk [1101]));
Q_ASSIGN U31674 ( .B(clk), .A(\g.we_clk [1100]));
Q_ASSIGN U31675 ( .B(clk), .A(\g.we_clk [1099]));
Q_ASSIGN U31676 ( .B(clk), .A(\g.we_clk [1098]));
Q_ASSIGN U31677 ( .B(clk), .A(\g.we_clk [1097]));
Q_ASSIGN U31678 ( .B(clk), .A(\g.we_clk [1096]));
Q_ASSIGN U31679 ( .B(clk), .A(\g.we_clk [1095]));
Q_ASSIGN U31680 ( .B(clk), .A(\g.we_clk [1094]));
Q_ASSIGN U31681 ( .B(clk), .A(\g.we_clk [1093]));
Q_ASSIGN U31682 ( .B(clk), .A(\g.we_clk [1092]));
Q_ASSIGN U31683 ( .B(clk), .A(\g.we_clk [1091]));
Q_ASSIGN U31684 ( .B(clk), .A(\g.we_clk [1090]));
Q_ASSIGN U31685 ( .B(clk), .A(\g.we_clk [1089]));
Q_ASSIGN U31686 ( .B(clk), .A(\g.we_clk [1088]));
Q_ASSIGN U31687 ( .B(clk), .A(\g.we_clk [1087]));
Q_ASSIGN U31688 ( .B(clk), .A(\g.we_clk [1086]));
Q_ASSIGN U31689 ( .B(clk), .A(\g.we_clk [1085]));
Q_ASSIGN U31690 ( .B(clk), .A(\g.we_clk [1084]));
Q_ASSIGN U31691 ( .B(clk), .A(\g.we_clk [1083]));
Q_ASSIGN U31692 ( .B(clk), .A(\g.we_clk [1082]));
Q_ASSIGN U31693 ( .B(clk), .A(\g.we_clk [1081]));
Q_ASSIGN U31694 ( .B(clk), .A(\g.we_clk [1080]));
Q_ASSIGN U31695 ( .B(clk), .A(\g.we_clk [1079]));
Q_ASSIGN U31696 ( .B(clk), .A(\g.we_clk [1078]));
Q_ASSIGN U31697 ( .B(clk), .A(\g.we_clk [1077]));
Q_ASSIGN U31698 ( .B(clk), .A(\g.we_clk [1076]));
Q_ASSIGN U31699 ( .B(clk), .A(\g.we_clk [1075]));
Q_ASSIGN U31700 ( .B(clk), .A(\g.we_clk [1074]));
Q_ASSIGN U31701 ( .B(clk), .A(\g.we_clk [1073]));
Q_ASSIGN U31702 ( .B(clk), .A(\g.we_clk [1072]));
Q_ASSIGN U31703 ( .B(clk), .A(\g.we_clk [1071]));
Q_ASSIGN U31704 ( .B(clk), .A(\g.we_clk [1070]));
Q_ASSIGN U31705 ( .B(clk), .A(\g.we_clk [1069]));
Q_ASSIGN U31706 ( .B(clk), .A(\g.we_clk [1068]));
Q_ASSIGN U31707 ( .B(clk), .A(\g.we_clk [1067]));
Q_ASSIGN U31708 ( .B(clk), .A(\g.we_clk [1066]));
Q_ASSIGN U31709 ( .B(clk), .A(\g.we_clk [1065]));
Q_ASSIGN U31710 ( .B(clk), .A(\g.we_clk [1064]));
Q_ASSIGN U31711 ( .B(clk), .A(\g.we_clk [1063]));
Q_ASSIGN U31712 ( .B(clk), .A(\g.we_clk [1062]));
Q_ASSIGN U31713 ( .B(clk), .A(\g.we_clk [1061]));
Q_ASSIGN U31714 ( .B(clk), .A(\g.we_clk [1060]));
Q_ASSIGN U31715 ( .B(clk), .A(\g.we_clk [1059]));
Q_ASSIGN U31716 ( .B(clk), .A(\g.we_clk [1058]));
Q_ASSIGN U31717 ( .B(clk), .A(\g.we_clk [1057]));
Q_ASSIGN U31718 ( .B(clk), .A(\g.we_clk [1056]));
Q_ASSIGN U31719 ( .B(clk), .A(\g.we_clk [1055]));
Q_ASSIGN U31720 ( .B(clk), .A(\g.we_clk [1054]));
Q_ASSIGN U31721 ( .B(clk), .A(\g.we_clk [1053]));
Q_ASSIGN U31722 ( .B(clk), .A(\g.we_clk [1052]));
Q_ASSIGN U31723 ( .B(clk), .A(\g.we_clk [1051]));
Q_ASSIGN U31724 ( .B(clk), .A(\g.we_clk [1050]));
Q_ASSIGN U31725 ( .B(clk), .A(\g.we_clk [1049]));
Q_ASSIGN U31726 ( .B(clk), .A(\g.we_clk [1048]));
Q_ASSIGN U31727 ( .B(clk), .A(\g.we_clk [1047]));
Q_ASSIGN U31728 ( .B(clk), .A(\g.we_clk [1046]));
Q_ASSIGN U31729 ( .B(clk), .A(\g.we_clk [1045]));
Q_ASSIGN U31730 ( .B(clk), .A(\g.we_clk [1044]));
Q_ASSIGN U31731 ( .B(clk), .A(\g.we_clk [1043]));
Q_ASSIGN U31732 ( .B(clk), .A(\g.we_clk [1042]));
Q_ASSIGN U31733 ( .B(clk), .A(\g.we_clk [1041]));
Q_ASSIGN U31734 ( .B(clk), .A(\g.we_clk [1040]));
Q_ASSIGN U31735 ( .B(clk), .A(\g.we_clk [1039]));
Q_ASSIGN U31736 ( .B(clk), .A(\g.we_clk [1038]));
Q_ASSIGN U31737 ( .B(clk), .A(\g.we_clk [1037]));
Q_ASSIGN U31738 ( .B(clk), .A(\g.we_clk [1036]));
Q_ASSIGN U31739 ( .B(clk), .A(\g.we_clk [1035]));
Q_ASSIGN U31740 ( .B(clk), .A(\g.we_clk [1034]));
Q_ASSIGN U31741 ( .B(clk), .A(\g.we_clk [1033]));
Q_ASSIGN U31742 ( .B(clk), .A(\g.we_clk [1032]));
Q_ASSIGN U31743 ( .B(clk), .A(\g.we_clk [1031]));
Q_ASSIGN U31744 ( .B(clk), .A(\g.we_clk [1030]));
Q_ASSIGN U31745 ( .B(clk), .A(\g.we_clk [1029]));
Q_ASSIGN U31746 ( .B(clk), .A(\g.we_clk [1028]));
Q_ASSIGN U31747 ( .B(clk), .A(\g.we_clk [1027]));
Q_ASSIGN U31748 ( .B(clk), .A(\g.we_clk [1026]));
Q_ASSIGN U31749 ( .B(clk), .A(\g.we_clk [1025]));
Q_ASSIGN U31750 ( .B(clk), .A(\g.we_clk [1024]));
Q_ASSIGN U31751 ( .B(clk), .A(\g.we_clk [1023]));
Q_ASSIGN U31752 ( .B(clk), .A(\g.we_clk [1022]));
Q_ASSIGN U31753 ( .B(clk), .A(\g.we_clk [1021]));
Q_ASSIGN U31754 ( .B(clk), .A(\g.we_clk [1020]));
Q_ASSIGN U31755 ( .B(clk), .A(\g.we_clk [1019]));
Q_ASSIGN U31756 ( .B(clk), .A(\g.we_clk [1018]));
Q_ASSIGN U31757 ( .B(clk), .A(\g.we_clk [1017]));
Q_ASSIGN U31758 ( .B(clk), .A(\g.we_clk [1016]));
Q_ASSIGN U31759 ( .B(clk), .A(\g.we_clk [1015]));
Q_ASSIGN U31760 ( .B(clk), .A(\g.we_clk [1014]));
Q_ASSIGN U31761 ( .B(clk), .A(\g.we_clk [1013]));
Q_ASSIGN U31762 ( .B(clk), .A(\g.we_clk [1012]));
Q_ASSIGN U31763 ( .B(clk), .A(\g.we_clk [1011]));
Q_ASSIGN U31764 ( .B(clk), .A(\g.we_clk [1010]));
Q_ASSIGN U31765 ( .B(clk), .A(\g.we_clk [1009]));
Q_ASSIGN U31766 ( .B(clk), .A(\g.we_clk [1008]));
Q_ASSIGN U31767 ( .B(clk), .A(\g.we_clk [1007]));
Q_ASSIGN U31768 ( .B(clk), .A(\g.we_clk [1006]));
Q_ASSIGN U31769 ( .B(clk), .A(\g.we_clk [1005]));
Q_ASSIGN U31770 ( .B(clk), .A(\g.we_clk [1004]));
Q_ASSIGN U31771 ( .B(clk), .A(\g.we_clk [1003]));
Q_ASSIGN U31772 ( .B(clk), .A(\g.we_clk [1002]));
Q_ASSIGN U31773 ( .B(clk), .A(\g.we_clk [1001]));
Q_ASSIGN U31774 ( .B(clk), .A(\g.we_clk [1000]));
Q_ASSIGN U31775 ( .B(clk), .A(\g.we_clk [999]));
Q_ASSIGN U31776 ( .B(clk), .A(\g.we_clk [998]));
Q_ASSIGN U31777 ( .B(clk), .A(\g.we_clk [997]));
Q_ASSIGN U31778 ( .B(clk), .A(\g.we_clk [996]));
Q_ASSIGN U31779 ( .B(clk), .A(\g.we_clk [995]));
Q_ASSIGN U31780 ( .B(clk), .A(\g.we_clk [994]));
Q_ASSIGN U31781 ( .B(clk), .A(\g.we_clk [993]));
Q_ASSIGN U31782 ( .B(clk), .A(\g.we_clk [992]));
Q_ASSIGN U31783 ( .B(clk), .A(\g.we_clk [991]));
Q_ASSIGN U31784 ( .B(clk), .A(\g.we_clk [990]));
Q_ASSIGN U31785 ( .B(clk), .A(\g.we_clk [989]));
Q_ASSIGN U31786 ( .B(clk), .A(\g.we_clk [988]));
Q_ASSIGN U31787 ( .B(clk), .A(\g.we_clk [987]));
Q_ASSIGN U31788 ( .B(clk), .A(\g.we_clk [986]));
Q_ASSIGN U31789 ( .B(clk), .A(\g.we_clk [985]));
Q_ASSIGN U31790 ( .B(clk), .A(\g.we_clk [984]));
Q_ASSIGN U31791 ( .B(clk), .A(\g.we_clk [983]));
Q_ASSIGN U31792 ( .B(clk), .A(\g.we_clk [982]));
Q_ASSIGN U31793 ( .B(clk), .A(\g.we_clk [981]));
Q_ASSIGN U31794 ( .B(clk), .A(\g.we_clk [980]));
Q_ASSIGN U31795 ( .B(clk), .A(\g.we_clk [979]));
Q_ASSIGN U31796 ( .B(clk), .A(\g.we_clk [978]));
Q_ASSIGN U31797 ( .B(clk), .A(\g.we_clk [977]));
Q_ASSIGN U31798 ( .B(clk), .A(\g.we_clk [976]));
Q_ASSIGN U31799 ( .B(clk), .A(\g.we_clk [975]));
Q_ASSIGN U31800 ( .B(clk), .A(\g.we_clk [974]));
Q_ASSIGN U31801 ( .B(clk), .A(\g.we_clk [973]));
Q_ASSIGN U31802 ( .B(clk), .A(\g.we_clk [972]));
Q_ASSIGN U31803 ( .B(clk), .A(\g.we_clk [971]));
Q_ASSIGN U31804 ( .B(clk), .A(\g.we_clk [970]));
Q_ASSIGN U31805 ( .B(clk), .A(\g.we_clk [969]));
Q_ASSIGN U31806 ( .B(clk), .A(\g.we_clk [968]));
Q_ASSIGN U31807 ( .B(clk), .A(\g.we_clk [967]));
Q_ASSIGN U31808 ( .B(clk), .A(\g.we_clk [966]));
Q_ASSIGN U31809 ( .B(clk), .A(\g.we_clk [965]));
Q_ASSIGN U31810 ( .B(clk), .A(\g.we_clk [964]));
Q_ASSIGN U31811 ( .B(clk), .A(\g.we_clk [963]));
Q_ASSIGN U31812 ( .B(clk), .A(\g.we_clk [962]));
Q_ASSIGN U31813 ( .B(clk), .A(\g.we_clk [961]));
Q_ASSIGN U31814 ( .B(clk), .A(\g.we_clk [960]));
Q_ASSIGN U31815 ( .B(clk), .A(\g.we_clk [959]));
Q_ASSIGN U31816 ( .B(clk), .A(\g.we_clk [958]));
Q_ASSIGN U31817 ( .B(clk), .A(\g.we_clk [957]));
Q_ASSIGN U31818 ( .B(clk), .A(\g.we_clk [956]));
Q_ASSIGN U31819 ( .B(clk), .A(\g.we_clk [955]));
Q_ASSIGN U31820 ( .B(clk), .A(\g.we_clk [954]));
Q_ASSIGN U31821 ( .B(clk), .A(\g.we_clk [953]));
Q_ASSIGN U31822 ( .B(clk), .A(\g.we_clk [952]));
Q_ASSIGN U31823 ( .B(clk), .A(\g.we_clk [951]));
Q_ASSIGN U31824 ( .B(clk), .A(\g.we_clk [950]));
Q_ASSIGN U31825 ( .B(clk), .A(\g.we_clk [949]));
Q_ASSIGN U31826 ( .B(clk), .A(\g.we_clk [948]));
Q_ASSIGN U31827 ( .B(clk), .A(\g.we_clk [947]));
Q_ASSIGN U31828 ( .B(clk), .A(\g.we_clk [946]));
Q_ASSIGN U31829 ( .B(clk), .A(\g.we_clk [945]));
Q_ASSIGN U31830 ( .B(clk), .A(\g.we_clk [944]));
Q_ASSIGN U31831 ( .B(clk), .A(\g.we_clk [943]));
Q_ASSIGN U31832 ( .B(clk), .A(\g.we_clk [942]));
Q_ASSIGN U31833 ( .B(clk), .A(\g.we_clk [941]));
Q_ASSIGN U31834 ( .B(clk), .A(\g.we_clk [940]));
Q_ASSIGN U31835 ( .B(clk), .A(\g.we_clk [939]));
Q_ASSIGN U31836 ( .B(clk), .A(\g.we_clk [938]));
Q_ASSIGN U31837 ( .B(clk), .A(\g.we_clk [937]));
Q_ASSIGN U31838 ( .B(clk), .A(\g.we_clk [936]));
Q_ASSIGN U31839 ( .B(clk), .A(\g.we_clk [935]));
Q_ASSIGN U31840 ( .B(clk), .A(\g.we_clk [934]));
Q_ASSIGN U31841 ( .B(clk), .A(\g.we_clk [933]));
Q_ASSIGN U31842 ( .B(clk), .A(\g.we_clk [932]));
Q_ASSIGN U31843 ( .B(clk), .A(\g.we_clk [931]));
Q_ASSIGN U31844 ( .B(clk), .A(\g.we_clk [930]));
Q_ASSIGN U31845 ( .B(clk), .A(\g.we_clk [929]));
Q_ASSIGN U31846 ( .B(clk), .A(\g.we_clk [928]));
Q_ASSIGN U31847 ( .B(clk), .A(\g.we_clk [927]));
Q_ASSIGN U31848 ( .B(clk), .A(\g.we_clk [926]));
Q_ASSIGN U31849 ( .B(clk), .A(\g.we_clk [925]));
Q_ASSIGN U31850 ( .B(clk), .A(\g.we_clk [924]));
Q_ASSIGN U31851 ( .B(clk), .A(\g.we_clk [923]));
Q_ASSIGN U31852 ( .B(clk), .A(\g.we_clk [922]));
Q_ASSIGN U31853 ( .B(clk), .A(\g.we_clk [921]));
Q_ASSIGN U31854 ( .B(clk), .A(\g.we_clk [920]));
Q_ASSIGN U31855 ( .B(clk), .A(\g.we_clk [919]));
Q_ASSIGN U31856 ( .B(clk), .A(\g.we_clk [918]));
Q_ASSIGN U31857 ( .B(clk), .A(\g.we_clk [917]));
Q_ASSIGN U31858 ( .B(clk), .A(\g.we_clk [916]));
Q_ASSIGN U31859 ( .B(clk), .A(\g.we_clk [915]));
Q_ASSIGN U31860 ( .B(clk), .A(\g.we_clk [914]));
Q_ASSIGN U31861 ( .B(clk), .A(\g.we_clk [913]));
Q_ASSIGN U31862 ( .B(clk), .A(\g.we_clk [912]));
Q_ASSIGN U31863 ( .B(clk), .A(\g.we_clk [911]));
Q_ASSIGN U31864 ( .B(clk), .A(\g.we_clk [910]));
Q_ASSIGN U31865 ( .B(clk), .A(\g.we_clk [909]));
Q_ASSIGN U31866 ( .B(clk), .A(\g.we_clk [908]));
Q_ASSIGN U31867 ( .B(clk), .A(\g.we_clk [907]));
Q_ASSIGN U31868 ( .B(clk), .A(\g.we_clk [906]));
Q_ASSIGN U31869 ( .B(clk), .A(\g.we_clk [905]));
Q_ASSIGN U31870 ( .B(clk), .A(\g.we_clk [904]));
Q_ASSIGN U31871 ( .B(clk), .A(\g.we_clk [903]));
Q_ASSIGN U31872 ( .B(clk), .A(\g.we_clk [902]));
Q_ASSIGN U31873 ( .B(clk), .A(\g.we_clk [901]));
Q_ASSIGN U31874 ( .B(clk), .A(\g.we_clk [900]));
Q_ASSIGN U31875 ( .B(clk), .A(\g.we_clk [899]));
Q_ASSIGN U31876 ( .B(clk), .A(\g.we_clk [898]));
Q_ASSIGN U31877 ( .B(clk), .A(\g.we_clk [897]));
Q_ASSIGN U31878 ( .B(clk), .A(\g.we_clk [896]));
Q_ASSIGN U31879 ( .B(clk), .A(\g.we_clk [895]));
Q_ASSIGN U31880 ( .B(clk), .A(\g.we_clk [894]));
Q_ASSIGN U31881 ( .B(clk), .A(\g.we_clk [893]));
Q_ASSIGN U31882 ( .B(clk), .A(\g.we_clk [892]));
Q_ASSIGN U31883 ( .B(clk), .A(\g.we_clk [891]));
Q_ASSIGN U31884 ( .B(clk), .A(\g.we_clk [890]));
Q_ASSIGN U31885 ( .B(clk), .A(\g.we_clk [889]));
Q_ASSIGN U31886 ( .B(clk), .A(\g.we_clk [888]));
Q_ASSIGN U31887 ( .B(clk), .A(\g.we_clk [887]));
Q_ASSIGN U31888 ( .B(clk), .A(\g.we_clk [886]));
Q_ASSIGN U31889 ( .B(clk), .A(\g.we_clk [885]));
Q_ASSIGN U31890 ( .B(clk), .A(\g.we_clk [884]));
Q_ASSIGN U31891 ( .B(clk), .A(\g.we_clk [883]));
Q_ASSIGN U31892 ( .B(clk), .A(\g.we_clk [882]));
Q_ASSIGN U31893 ( .B(clk), .A(\g.we_clk [881]));
Q_ASSIGN U31894 ( .B(clk), .A(\g.we_clk [880]));
Q_ASSIGN U31895 ( .B(clk), .A(\g.we_clk [879]));
Q_ASSIGN U31896 ( .B(clk), .A(\g.we_clk [878]));
Q_ASSIGN U31897 ( .B(clk), .A(\g.we_clk [877]));
Q_ASSIGN U31898 ( .B(clk), .A(\g.we_clk [876]));
Q_ASSIGN U31899 ( .B(clk), .A(\g.we_clk [875]));
Q_ASSIGN U31900 ( .B(clk), .A(\g.we_clk [874]));
Q_ASSIGN U31901 ( .B(clk), .A(\g.we_clk [873]));
Q_ASSIGN U31902 ( .B(clk), .A(\g.we_clk [872]));
Q_ASSIGN U31903 ( .B(clk), .A(\g.we_clk [871]));
Q_ASSIGN U31904 ( .B(clk), .A(\g.we_clk [870]));
Q_ASSIGN U31905 ( .B(clk), .A(\g.we_clk [869]));
Q_ASSIGN U31906 ( .B(clk), .A(\g.we_clk [868]));
Q_ASSIGN U31907 ( .B(clk), .A(\g.we_clk [867]));
Q_ASSIGN U31908 ( .B(clk), .A(\g.we_clk [866]));
Q_ASSIGN U31909 ( .B(clk), .A(\g.we_clk [865]));
Q_ASSIGN U31910 ( .B(clk), .A(\g.we_clk [864]));
Q_ASSIGN U31911 ( .B(clk), .A(\g.we_clk [863]));
Q_ASSIGN U31912 ( .B(clk), .A(\g.we_clk [862]));
Q_ASSIGN U31913 ( .B(clk), .A(\g.we_clk [861]));
Q_ASSIGN U31914 ( .B(clk), .A(\g.we_clk [860]));
Q_ASSIGN U31915 ( .B(clk), .A(\g.we_clk [859]));
Q_ASSIGN U31916 ( .B(clk), .A(\g.we_clk [858]));
Q_ASSIGN U31917 ( .B(clk), .A(\g.we_clk [857]));
Q_ASSIGN U31918 ( .B(clk), .A(\g.we_clk [856]));
Q_ASSIGN U31919 ( .B(clk), .A(\g.we_clk [855]));
Q_ASSIGN U31920 ( .B(clk), .A(\g.we_clk [854]));
Q_ASSIGN U31921 ( .B(clk), .A(\g.we_clk [853]));
Q_ASSIGN U31922 ( .B(clk), .A(\g.we_clk [852]));
Q_ASSIGN U31923 ( .B(clk), .A(\g.we_clk [851]));
Q_ASSIGN U31924 ( .B(clk), .A(\g.we_clk [850]));
Q_ASSIGN U31925 ( .B(clk), .A(\g.we_clk [849]));
Q_ASSIGN U31926 ( .B(clk), .A(\g.we_clk [848]));
Q_ASSIGN U31927 ( .B(clk), .A(\g.we_clk [847]));
Q_ASSIGN U31928 ( .B(clk), .A(\g.we_clk [846]));
Q_ASSIGN U31929 ( .B(clk), .A(\g.we_clk [845]));
Q_ASSIGN U31930 ( .B(clk), .A(\g.we_clk [844]));
Q_ASSIGN U31931 ( .B(clk), .A(\g.we_clk [843]));
Q_ASSIGN U31932 ( .B(clk), .A(\g.we_clk [842]));
Q_ASSIGN U31933 ( .B(clk), .A(\g.we_clk [841]));
Q_ASSIGN U31934 ( .B(clk), .A(\g.we_clk [840]));
Q_ASSIGN U31935 ( .B(clk), .A(\g.we_clk [839]));
Q_ASSIGN U31936 ( .B(clk), .A(\g.we_clk [838]));
Q_ASSIGN U31937 ( .B(clk), .A(\g.we_clk [837]));
Q_ASSIGN U31938 ( .B(clk), .A(\g.we_clk [836]));
Q_ASSIGN U31939 ( .B(clk), .A(\g.we_clk [835]));
Q_ASSIGN U31940 ( .B(clk), .A(\g.we_clk [834]));
Q_ASSIGN U31941 ( .B(clk), .A(\g.we_clk [833]));
Q_ASSIGN U31942 ( .B(clk), .A(\g.we_clk [832]));
Q_ASSIGN U31943 ( .B(clk), .A(\g.we_clk [831]));
Q_ASSIGN U31944 ( .B(clk), .A(\g.we_clk [830]));
Q_ASSIGN U31945 ( .B(clk), .A(\g.we_clk [829]));
Q_ASSIGN U31946 ( .B(clk), .A(\g.we_clk [828]));
Q_ASSIGN U31947 ( .B(clk), .A(\g.we_clk [827]));
Q_ASSIGN U31948 ( .B(clk), .A(\g.we_clk [826]));
Q_ASSIGN U31949 ( .B(clk), .A(\g.we_clk [825]));
Q_ASSIGN U31950 ( .B(clk), .A(\g.we_clk [824]));
Q_ASSIGN U31951 ( .B(clk), .A(\g.we_clk [823]));
Q_ASSIGN U31952 ( .B(clk), .A(\g.we_clk [822]));
Q_ASSIGN U31953 ( .B(clk), .A(\g.we_clk [821]));
Q_ASSIGN U31954 ( .B(clk), .A(\g.we_clk [820]));
Q_ASSIGN U31955 ( .B(clk), .A(\g.we_clk [819]));
Q_ASSIGN U31956 ( .B(clk), .A(\g.we_clk [818]));
Q_ASSIGN U31957 ( .B(clk), .A(\g.we_clk [817]));
Q_ASSIGN U31958 ( .B(clk), .A(\g.we_clk [816]));
Q_ASSIGN U31959 ( .B(clk), .A(\g.we_clk [815]));
Q_ASSIGN U31960 ( .B(clk), .A(\g.we_clk [814]));
Q_ASSIGN U31961 ( .B(clk), .A(\g.we_clk [813]));
Q_ASSIGN U31962 ( .B(clk), .A(\g.we_clk [812]));
Q_ASSIGN U31963 ( .B(clk), .A(\g.we_clk [811]));
Q_ASSIGN U31964 ( .B(clk), .A(\g.we_clk [810]));
Q_ASSIGN U31965 ( .B(clk), .A(\g.we_clk [809]));
Q_ASSIGN U31966 ( .B(clk), .A(\g.we_clk [808]));
Q_ASSIGN U31967 ( .B(clk), .A(\g.we_clk [807]));
Q_ASSIGN U31968 ( .B(clk), .A(\g.we_clk [806]));
Q_ASSIGN U31969 ( .B(clk), .A(\g.we_clk [805]));
Q_ASSIGN U31970 ( .B(clk), .A(\g.we_clk [804]));
Q_ASSIGN U31971 ( .B(clk), .A(\g.we_clk [803]));
Q_ASSIGN U31972 ( .B(clk), .A(\g.we_clk [802]));
Q_ASSIGN U31973 ( .B(clk), .A(\g.we_clk [801]));
Q_ASSIGN U31974 ( .B(clk), .A(\g.we_clk [800]));
Q_ASSIGN U31975 ( .B(clk), .A(\g.we_clk [799]));
Q_ASSIGN U31976 ( .B(clk), .A(\g.we_clk [798]));
Q_ASSIGN U31977 ( .B(clk), .A(\g.we_clk [797]));
Q_ASSIGN U31978 ( .B(clk), .A(\g.we_clk [796]));
Q_ASSIGN U31979 ( .B(clk), .A(\g.we_clk [795]));
Q_ASSIGN U31980 ( .B(clk), .A(\g.we_clk [794]));
Q_ASSIGN U31981 ( .B(clk), .A(\g.we_clk [793]));
Q_ASSIGN U31982 ( .B(clk), .A(\g.we_clk [792]));
Q_ASSIGN U31983 ( .B(clk), .A(\g.we_clk [791]));
Q_ASSIGN U31984 ( .B(clk), .A(\g.we_clk [790]));
Q_ASSIGN U31985 ( .B(clk), .A(\g.we_clk [789]));
Q_ASSIGN U31986 ( .B(clk), .A(\g.we_clk [788]));
Q_ASSIGN U31987 ( .B(clk), .A(\g.we_clk [787]));
Q_ASSIGN U31988 ( .B(clk), .A(\g.we_clk [786]));
Q_ASSIGN U31989 ( .B(clk), .A(\g.we_clk [785]));
Q_ASSIGN U31990 ( .B(clk), .A(\g.we_clk [784]));
Q_ASSIGN U31991 ( .B(clk), .A(\g.we_clk [783]));
Q_ASSIGN U31992 ( .B(clk), .A(\g.we_clk [782]));
Q_ASSIGN U31993 ( .B(clk), .A(\g.we_clk [781]));
Q_ASSIGN U31994 ( .B(clk), .A(\g.we_clk [780]));
Q_ASSIGN U31995 ( .B(clk), .A(\g.we_clk [779]));
Q_ASSIGN U31996 ( .B(clk), .A(\g.we_clk [778]));
Q_ASSIGN U31997 ( .B(clk), .A(\g.we_clk [777]));
Q_ASSIGN U31998 ( .B(clk), .A(\g.we_clk [776]));
Q_ASSIGN U31999 ( .B(clk), .A(\g.we_clk [775]));
Q_ASSIGN U32000 ( .B(clk), .A(\g.we_clk [774]));
Q_ASSIGN U32001 ( .B(clk), .A(\g.we_clk [773]));
Q_ASSIGN U32002 ( .B(clk), .A(\g.we_clk [772]));
Q_ASSIGN U32003 ( .B(clk), .A(\g.we_clk [771]));
Q_ASSIGN U32004 ( .B(clk), .A(\g.we_clk [770]));
Q_ASSIGN U32005 ( .B(clk), .A(\g.we_clk [769]));
Q_ASSIGN U32006 ( .B(clk), .A(\g.we_clk [768]));
Q_ASSIGN U32007 ( .B(clk), .A(\g.we_clk [767]));
Q_ASSIGN U32008 ( .B(clk), .A(\g.we_clk [766]));
Q_ASSIGN U32009 ( .B(clk), .A(\g.we_clk [765]));
Q_ASSIGN U32010 ( .B(clk), .A(\g.we_clk [764]));
Q_ASSIGN U32011 ( .B(clk), .A(\g.we_clk [763]));
Q_ASSIGN U32012 ( .B(clk), .A(\g.we_clk [762]));
Q_ASSIGN U32013 ( .B(clk), .A(\g.we_clk [761]));
Q_ASSIGN U32014 ( .B(clk), .A(\g.we_clk [760]));
Q_ASSIGN U32015 ( .B(clk), .A(\g.we_clk [759]));
Q_ASSIGN U32016 ( .B(clk), .A(\g.we_clk [758]));
Q_ASSIGN U32017 ( .B(clk), .A(\g.we_clk [757]));
Q_ASSIGN U32018 ( .B(clk), .A(\g.we_clk [756]));
Q_ASSIGN U32019 ( .B(clk), .A(\g.we_clk [755]));
Q_ASSIGN U32020 ( .B(clk), .A(\g.we_clk [754]));
Q_ASSIGN U32021 ( .B(clk), .A(\g.we_clk [753]));
Q_ASSIGN U32022 ( .B(clk), .A(\g.we_clk [752]));
Q_ASSIGN U32023 ( .B(clk), .A(\g.we_clk [751]));
Q_ASSIGN U32024 ( .B(clk), .A(\g.we_clk [750]));
Q_ASSIGN U32025 ( .B(clk), .A(\g.we_clk [749]));
Q_ASSIGN U32026 ( .B(clk), .A(\g.we_clk [748]));
Q_ASSIGN U32027 ( .B(clk), .A(\g.we_clk [747]));
Q_ASSIGN U32028 ( .B(clk), .A(\g.we_clk [746]));
Q_ASSIGN U32029 ( .B(clk), .A(\g.we_clk [745]));
Q_ASSIGN U32030 ( .B(clk), .A(\g.we_clk [744]));
Q_ASSIGN U32031 ( .B(clk), .A(\g.we_clk [743]));
Q_ASSIGN U32032 ( .B(clk), .A(\g.we_clk [742]));
Q_ASSIGN U32033 ( .B(clk), .A(\g.we_clk [741]));
Q_ASSIGN U32034 ( .B(clk), .A(\g.we_clk [740]));
Q_ASSIGN U32035 ( .B(clk), .A(\g.we_clk [739]));
Q_ASSIGN U32036 ( .B(clk), .A(\g.we_clk [738]));
Q_ASSIGN U32037 ( .B(clk), .A(\g.we_clk [737]));
Q_ASSIGN U32038 ( .B(clk), .A(\g.we_clk [736]));
Q_ASSIGN U32039 ( .B(clk), .A(\g.we_clk [735]));
Q_ASSIGN U32040 ( .B(clk), .A(\g.we_clk [734]));
Q_ASSIGN U32041 ( .B(clk), .A(\g.we_clk [733]));
Q_ASSIGN U32042 ( .B(clk), .A(\g.we_clk [732]));
Q_ASSIGN U32043 ( .B(clk), .A(\g.we_clk [731]));
Q_ASSIGN U32044 ( .B(clk), .A(\g.we_clk [730]));
Q_ASSIGN U32045 ( .B(clk), .A(\g.we_clk [729]));
Q_ASSIGN U32046 ( .B(clk), .A(\g.we_clk [728]));
Q_ASSIGN U32047 ( .B(clk), .A(\g.we_clk [727]));
Q_ASSIGN U32048 ( .B(clk), .A(\g.we_clk [726]));
Q_ASSIGN U32049 ( .B(clk), .A(\g.we_clk [725]));
Q_ASSIGN U32050 ( .B(clk), .A(\g.we_clk [724]));
Q_ASSIGN U32051 ( .B(clk), .A(\g.we_clk [723]));
Q_ASSIGN U32052 ( .B(clk), .A(\g.we_clk [722]));
Q_ASSIGN U32053 ( .B(clk), .A(\g.we_clk [721]));
Q_ASSIGN U32054 ( .B(clk), .A(\g.we_clk [720]));
Q_ASSIGN U32055 ( .B(clk), .A(\g.we_clk [719]));
Q_ASSIGN U32056 ( .B(clk), .A(\g.we_clk [718]));
Q_ASSIGN U32057 ( .B(clk), .A(\g.we_clk [717]));
Q_ASSIGN U32058 ( .B(clk), .A(\g.we_clk [716]));
Q_ASSIGN U32059 ( .B(clk), .A(\g.we_clk [715]));
Q_ASSIGN U32060 ( .B(clk), .A(\g.we_clk [714]));
Q_ASSIGN U32061 ( .B(clk), .A(\g.we_clk [713]));
Q_ASSIGN U32062 ( .B(clk), .A(\g.we_clk [712]));
Q_ASSIGN U32063 ( .B(clk), .A(\g.we_clk [711]));
Q_ASSIGN U32064 ( .B(clk), .A(\g.we_clk [710]));
Q_ASSIGN U32065 ( .B(clk), .A(\g.we_clk [709]));
Q_ASSIGN U32066 ( .B(clk), .A(\g.we_clk [708]));
Q_ASSIGN U32067 ( .B(clk), .A(\g.we_clk [707]));
Q_ASSIGN U32068 ( .B(clk), .A(\g.we_clk [706]));
Q_ASSIGN U32069 ( .B(clk), .A(\g.we_clk [705]));
Q_ASSIGN U32070 ( .B(clk), .A(\g.we_clk [704]));
Q_ASSIGN U32071 ( .B(clk), .A(\g.we_clk [703]));
Q_ASSIGN U32072 ( .B(clk), .A(\g.we_clk [702]));
Q_ASSIGN U32073 ( .B(clk), .A(\g.we_clk [701]));
Q_ASSIGN U32074 ( .B(clk), .A(\g.we_clk [700]));
Q_ASSIGN U32075 ( .B(clk), .A(\g.we_clk [699]));
Q_ASSIGN U32076 ( .B(clk), .A(\g.we_clk [698]));
Q_ASSIGN U32077 ( .B(clk), .A(\g.we_clk [697]));
Q_ASSIGN U32078 ( .B(clk), .A(\g.we_clk [696]));
Q_ASSIGN U32079 ( .B(clk), .A(\g.we_clk [695]));
Q_ASSIGN U32080 ( .B(clk), .A(\g.we_clk [694]));
Q_ASSIGN U32081 ( .B(clk), .A(\g.we_clk [693]));
Q_ASSIGN U32082 ( .B(clk), .A(\g.we_clk [692]));
Q_ASSIGN U32083 ( .B(clk), .A(\g.we_clk [691]));
Q_ASSIGN U32084 ( .B(clk), .A(\g.we_clk [690]));
Q_ASSIGN U32085 ( .B(clk), .A(\g.we_clk [689]));
Q_ASSIGN U32086 ( .B(clk), .A(\g.we_clk [688]));
Q_ASSIGN U32087 ( .B(clk), .A(\g.we_clk [687]));
Q_ASSIGN U32088 ( .B(clk), .A(\g.we_clk [686]));
Q_ASSIGN U32089 ( .B(clk), .A(\g.we_clk [685]));
Q_ASSIGN U32090 ( .B(clk), .A(\g.we_clk [684]));
Q_ASSIGN U32091 ( .B(clk), .A(\g.we_clk [683]));
Q_ASSIGN U32092 ( .B(clk), .A(\g.we_clk [682]));
Q_ASSIGN U32093 ( .B(clk), .A(\g.we_clk [681]));
Q_ASSIGN U32094 ( .B(clk), .A(\g.we_clk [680]));
Q_ASSIGN U32095 ( .B(clk), .A(\g.we_clk [679]));
Q_ASSIGN U32096 ( .B(clk), .A(\g.we_clk [678]));
Q_ASSIGN U32097 ( .B(clk), .A(\g.we_clk [677]));
Q_ASSIGN U32098 ( .B(clk), .A(\g.we_clk [676]));
Q_ASSIGN U32099 ( .B(clk), .A(\g.we_clk [675]));
Q_ASSIGN U32100 ( .B(clk), .A(\g.we_clk [674]));
Q_ASSIGN U32101 ( .B(clk), .A(\g.we_clk [673]));
Q_ASSIGN U32102 ( .B(clk), .A(\g.we_clk [672]));
Q_ASSIGN U32103 ( .B(clk), .A(\g.we_clk [671]));
Q_ASSIGN U32104 ( .B(clk), .A(\g.we_clk [670]));
Q_ASSIGN U32105 ( .B(clk), .A(\g.we_clk [669]));
Q_ASSIGN U32106 ( .B(clk), .A(\g.we_clk [668]));
Q_ASSIGN U32107 ( .B(clk), .A(\g.we_clk [667]));
Q_ASSIGN U32108 ( .B(clk), .A(\g.we_clk [666]));
Q_ASSIGN U32109 ( .B(clk), .A(\g.we_clk [665]));
Q_ASSIGN U32110 ( .B(clk), .A(\g.we_clk [664]));
Q_ASSIGN U32111 ( .B(clk), .A(\g.we_clk [663]));
Q_ASSIGN U32112 ( .B(clk), .A(\g.we_clk [662]));
Q_ASSIGN U32113 ( .B(clk), .A(\g.we_clk [661]));
Q_ASSIGN U32114 ( .B(clk), .A(\g.we_clk [660]));
Q_ASSIGN U32115 ( .B(clk), .A(\g.we_clk [659]));
Q_ASSIGN U32116 ( .B(clk), .A(\g.we_clk [658]));
Q_ASSIGN U32117 ( .B(clk), .A(\g.we_clk [657]));
Q_ASSIGN U32118 ( .B(clk), .A(\g.we_clk [656]));
Q_ASSIGN U32119 ( .B(clk), .A(\g.we_clk [655]));
Q_ASSIGN U32120 ( .B(clk), .A(\g.we_clk [654]));
Q_ASSIGN U32121 ( .B(clk), .A(\g.we_clk [653]));
Q_ASSIGN U32122 ( .B(clk), .A(\g.we_clk [652]));
Q_ASSIGN U32123 ( .B(clk), .A(\g.we_clk [651]));
Q_ASSIGN U32124 ( .B(clk), .A(\g.we_clk [650]));
Q_ASSIGN U32125 ( .B(clk), .A(\g.we_clk [649]));
Q_ASSIGN U32126 ( .B(clk), .A(\g.we_clk [648]));
Q_ASSIGN U32127 ( .B(clk), .A(\g.we_clk [647]));
Q_ASSIGN U32128 ( .B(clk), .A(\g.we_clk [646]));
Q_ASSIGN U32129 ( .B(clk), .A(\g.we_clk [645]));
Q_ASSIGN U32130 ( .B(clk), .A(\g.we_clk [644]));
Q_ASSIGN U32131 ( .B(clk), .A(\g.we_clk [643]));
Q_ASSIGN U32132 ( .B(clk), .A(\g.we_clk [642]));
Q_ASSIGN U32133 ( .B(clk), .A(\g.we_clk [641]));
Q_ASSIGN U32134 ( .B(clk), .A(\g.we_clk [640]));
Q_ASSIGN U32135 ( .B(clk), .A(\g.we_clk [639]));
Q_ASSIGN U32136 ( .B(clk), .A(\g.we_clk [638]));
Q_ASSIGN U32137 ( .B(clk), .A(\g.we_clk [637]));
Q_ASSIGN U32138 ( .B(clk), .A(\g.we_clk [636]));
Q_ASSIGN U32139 ( .B(clk), .A(\g.we_clk [635]));
Q_ASSIGN U32140 ( .B(clk), .A(\g.we_clk [634]));
Q_ASSIGN U32141 ( .B(clk), .A(\g.we_clk [633]));
Q_ASSIGN U32142 ( .B(clk), .A(\g.we_clk [632]));
Q_ASSIGN U32143 ( .B(clk), .A(\g.we_clk [631]));
Q_ASSIGN U32144 ( .B(clk), .A(\g.we_clk [630]));
Q_ASSIGN U32145 ( .B(clk), .A(\g.we_clk [629]));
Q_ASSIGN U32146 ( .B(clk), .A(\g.we_clk [628]));
Q_ASSIGN U32147 ( .B(clk), .A(\g.we_clk [627]));
Q_ASSIGN U32148 ( .B(clk), .A(\g.we_clk [626]));
Q_ASSIGN U32149 ( .B(clk), .A(\g.we_clk [625]));
Q_ASSIGN U32150 ( .B(clk), .A(\g.we_clk [624]));
Q_ASSIGN U32151 ( .B(clk), .A(\g.we_clk [623]));
Q_ASSIGN U32152 ( .B(clk), .A(\g.we_clk [622]));
Q_ASSIGN U32153 ( .B(clk), .A(\g.we_clk [621]));
Q_ASSIGN U32154 ( .B(clk), .A(\g.we_clk [620]));
Q_ASSIGN U32155 ( .B(clk), .A(\g.we_clk [619]));
Q_ASSIGN U32156 ( .B(clk), .A(\g.we_clk [618]));
Q_ASSIGN U32157 ( .B(clk), .A(\g.we_clk [617]));
Q_ASSIGN U32158 ( .B(clk), .A(\g.we_clk [616]));
Q_ASSIGN U32159 ( .B(clk), .A(\g.we_clk [615]));
Q_ASSIGN U32160 ( .B(clk), .A(\g.we_clk [614]));
Q_ASSIGN U32161 ( .B(clk), .A(\g.we_clk [613]));
Q_ASSIGN U32162 ( .B(clk), .A(\g.we_clk [612]));
Q_ASSIGN U32163 ( .B(clk), .A(\g.we_clk [611]));
Q_ASSIGN U32164 ( .B(clk), .A(\g.we_clk [610]));
Q_ASSIGN U32165 ( .B(clk), .A(\g.we_clk [609]));
Q_ASSIGN U32166 ( .B(clk), .A(\g.we_clk [608]));
Q_ASSIGN U32167 ( .B(clk), .A(\g.we_clk [607]));
Q_ASSIGN U32168 ( .B(clk), .A(\g.we_clk [606]));
Q_ASSIGN U32169 ( .B(clk), .A(\g.we_clk [605]));
Q_ASSIGN U32170 ( .B(clk), .A(\g.we_clk [604]));
Q_ASSIGN U32171 ( .B(clk), .A(\g.we_clk [603]));
Q_ASSIGN U32172 ( .B(clk), .A(\g.we_clk [602]));
Q_ASSIGN U32173 ( .B(clk), .A(\g.we_clk [601]));
Q_ASSIGN U32174 ( .B(clk), .A(\g.we_clk [600]));
Q_ASSIGN U32175 ( .B(clk), .A(\g.we_clk [599]));
Q_ASSIGN U32176 ( .B(clk), .A(\g.we_clk [598]));
Q_ASSIGN U32177 ( .B(clk), .A(\g.we_clk [597]));
Q_ASSIGN U32178 ( .B(clk), .A(\g.we_clk [596]));
Q_ASSIGN U32179 ( .B(clk), .A(\g.we_clk [595]));
Q_ASSIGN U32180 ( .B(clk), .A(\g.we_clk [594]));
Q_ASSIGN U32181 ( .B(clk), .A(\g.we_clk [593]));
Q_ASSIGN U32182 ( .B(clk), .A(\g.we_clk [592]));
Q_ASSIGN U32183 ( .B(clk), .A(\g.we_clk [591]));
Q_ASSIGN U32184 ( .B(clk), .A(\g.we_clk [590]));
Q_ASSIGN U32185 ( .B(clk), .A(\g.we_clk [589]));
Q_ASSIGN U32186 ( .B(clk), .A(\g.we_clk [588]));
Q_ASSIGN U32187 ( .B(clk), .A(\g.we_clk [587]));
Q_ASSIGN U32188 ( .B(clk), .A(\g.we_clk [586]));
Q_ASSIGN U32189 ( .B(clk), .A(\g.we_clk [585]));
Q_ASSIGN U32190 ( .B(clk), .A(\g.we_clk [584]));
Q_ASSIGN U32191 ( .B(clk), .A(\g.we_clk [583]));
Q_ASSIGN U32192 ( .B(clk), .A(\g.we_clk [582]));
Q_ASSIGN U32193 ( .B(clk), .A(\g.we_clk [581]));
Q_ASSIGN U32194 ( .B(clk), .A(\g.we_clk [580]));
Q_ASSIGN U32195 ( .B(clk), .A(\g.we_clk [579]));
Q_ASSIGN U32196 ( .B(clk), .A(\g.we_clk [578]));
Q_ASSIGN U32197 ( .B(clk), .A(\g.we_clk [577]));
Q_ASSIGN U32198 ( .B(clk), .A(\g.we_clk [576]));
Q_ASSIGN U32199 ( .B(clk), .A(\g.we_clk [575]));
Q_ASSIGN U32200 ( .B(clk), .A(\g.we_clk [574]));
Q_ASSIGN U32201 ( .B(clk), .A(\g.we_clk [573]));
Q_ASSIGN U32202 ( .B(clk), .A(\g.we_clk [572]));
Q_ASSIGN U32203 ( .B(clk), .A(\g.we_clk [571]));
Q_ASSIGN U32204 ( .B(clk), .A(\g.we_clk [570]));
Q_ASSIGN U32205 ( .B(clk), .A(\g.we_clk [569]));
Q_ASSIGN U32206 ( .B(clk), .A(\g.we_clk [568]));
Q_ASSIGN U32207 ( .B(clk), .A(\g.we_clk [567]));
Q_ASSIGN U32208 ( .B(clk), .A(\g.we_clk [566]));
Q_ASSIGN U32209 ( .B(clk), .A(\g.we_clk [565]));
Q_ASSIGN U32210 ( .B(clk), .A(\g.we_clk [564]));
Q_ASSIGN U32211 ( .B(clk), .A(\g.we_clk [563]));
Q_ASSIGN U32212 ( .B(clk), .A(\g.we_clk [562]));
Q_ASSIGN U32213 ( .B(clk), .A(\g.we_clk [561]));
Q_ASSIGN U32214 ( .B(clk), .A(\g.we_clk [560]));
Q_ASSIGN U32215 ( .B(clk), .A(\g.we_clk [559]));
Q_ASSIGN U32216 ( .B(clk), .A(\g.we_clk [558]));
Q_ASSIGN U32217 ( .B(clk), .A(\g.we_clk [557]));
Q_ASSIGN U32218 ( .B(clk), .A(\g.we_clk [556]));
Q_ASSIGN U32219 ( .B(clk), .A(\g.we_clk [555]));
Q_ASSIGN U32220 ( .B(clk), .A(\g.we_clk [554]));
Q_ASSIGN U32221 ( .B(clk), .A(\g.we_clk [553]));
Q_ASSIGN U32222 ( .B(clk), .A(\g.we_clk [552]));
Q_ASSIGN U32223 ( .B(clk), .A(\g.we_clk [551]));
Q_ASSIGN U32224 ( .B(clk), .A(\g.we_clk [550]));
Q_ASSIGN U32225 ( .B(clk), .A(\g.we_clk [549]));
Q_ASSIGN U32226 ( .B(clk), .A(\g.we_clk [548]));
Q_ASSIGN U32227 ( .B(clk), .A(\g.we_clk [547]));
Q_ASSIGN U32228 ( .B(clk), .A(\g.we_clk [546]));
Q_ASSIGN U32229 ( .B(clk), .A(\g.we_clk [545]));
Q_ASSIGN U32230 ( .B(clk), .A(\g.we_clk [544]));
Q_ASSIGN U32231 ( .B(clk), .A(\g.we_clk [543]));
Q_ASSIGN U32232 ( .B(clk), .A(\g.we_clk [542]));
Q_ASSIGN U32233 ( .B(clk), .A(\g.we_clk [541]));
Q_ASSIGN U32234 ( .B(clk), .A(\g.we_clk [540]));
Q_ASSIGN U32235 ( .B(clk), .A(\g.we_clk [539]));
Q_ASSIGN U32236 ( .B(clk), .A(\g.we_clk [538]));
Q_ASSIGN U32237 ( .B(clk), .A(\g.we_clk [537]));
Q_ASSIGN U32238 ( .B(clk), .A(\g.we_clk [536]));
Q_ASSIGN U32239 ( .B(clk), .A(\g.we_clk [535]));
Q_ASSIGN U32240 ( .B(clk), .A(\g.we_clk [534]));
Q_ASSIGN U32241 ( .B(clk), .A(\g.we_clk [533]));
Q_ASSIGN U32242 ( .B(clk), .A(\g.we_clk [532]));
Q_ASSIGN U32243 ( .B(clk), .A(\g.we_clk [531]));
Q_ASSIGN U32244 ( .B(clk), .A(\g.we_clk [530]));
Q_ASSIGN U32245 ( .B(clk), .A(\g.we_clk [529]));
Q_ASSIGN U32246 ( .B(clk), .A(\g.we_clk [528]));
Q_ASSIGN U32247 ( .B(clk), .A(\g.we_clk [527]));
Q_ASSIGN U32248 ( .B(clk), .A(\g.we_clk [526]));
Q_ASSIGN U32249 ( .B(clk), .A(\g.we_clk [525]));
Q_ASSIGN U32250 ( .B(clk), .A(\g.we_clk [524]));
Q_ASSIGN U32251 ( .B(clk), .A(\g.we_clk [523]));
Q_ASSIGN U32252 ( .B(clk), .A(\g.we_clk [522]));
Q_ASSIGN U32253 ( .B(clk), .A(\g.we_clk [521]));
Q_ASSIGN U32254 ( .B(clk), .A(\g.we_clk [520]));
Q_ASSIGN U32255 ( .B(clk), .A(\g.we_clk [519]));
Q_ASSIGN U32256 ( .B(clk), .A(\g.we_clk [518]));
Q_ASSIGN U32257 ( .B(clk), .A(\g.we_clk [517]));
Q_ASSIGN U32258 ( .B(clk), .A(\g.we_clk [516]));
Q_ASSIGN U32259 ( .B(clk), .A(\g.we_clk [515]));
Q_ASSIGN U32260 ( .B(clk), .A(\g.we_clk [514]));
Q_ASSIGN U32261 ( .B(clk), .A(\g.we_clk [513]));
Q_ASSIGN U32262 ( .B(clk), .A(\g.we_clk [512]));
Q_ASSIGN U32263 ( .B(clk), .A(\g.we_clk [511]));
Q_ASSIGN U32264 ( .B(clk), .A(\g.we_clk [510]));
Q_ASSIGN U32265 ( .B(clk), .A(\g.we_clk [509]));
Q_ASSIGN U32266 ( .B(clk), .A(\g.we_clk [508]));
Q_ASSIGN U32267 ( .B(clk), .A(\g.we_clk [507]));
Q_ASSIGN U32268 ( .B(clk), .A(\g.we_clk [506]));
Q_ASSIGN U32269 ( .B(clk), .A(\g.we_clk [505]));
Q_ASSIGN U32270 ( .B(clk), .A(\g.we_clk [504]));
Q_ASSIGN U32271 ( .B(clk), .A(\g.we_clk [503]));
Q_ASSIGN U32272 ( .B(clk), .A(\g.we_clk [502]));
Q_ASSIGN U32273 ( .B(clk), .A(\g.we_clk [501]));
Q_ASSIGN U32274 ( .B(clk), .A(\g.we_clk [500]));
Q_ASSIGN U32275 ( .B(clk), .A(\g.we_clk [499]));
Q_ASSIGN U32276 ( .B(clk), .A(\g.we_clk [498]));
Q_ASSIGN U32277 ( .B(clk), .A(\g.we_clk [497]));
Q_ASSIGN U32278 ( .B(clk), .A(\g.we_clk [496]));
Q_ASSIGN U32279 ( .B(clk), .A(\g.we_clk [495]));
Q_ASSIGN U32280 ( .B(clk), .A(\g.we_clk [494]));
Q_ASSIGN U32281 ( .B(clk), .A(\g.we_clk [493]));
Q_ASSIGN U32282 ( .B(clk), .A(\g.we_clk [492]));
Q_ASSIGN U32283 ( .B(clk), .A(\g.we_clk [491]));
Q_ASSIGN U32284 ( .B(clk), .A(\g.we_clk [490]));
Q_ASSIGN U32285 ( .B(clk), .A(\g.we_clk [489]));
Q_ASSIGN U32286 ( .B(clk), .A(\g.we_clk [488]));
Q_ASSIGN U32287 ( .B(clk), .A(\g.we_clk [487]));
Q_ASSIGN U32288 ( .B(clk), .A(\g.we_clk [486]));
Q_ASSIGN U32289 ( .B(clk), .A(\g.we_clk [485]));
Q_ASSIGN U32290 ( .B(clk), .A(\g.we_clk [484]));
Q_ASSIGN U32291 ( .B(clk), .A(\g.we_clk [483]));
Q_ASSIGN U32292 ( .B(clk), .A(\g.we_clk [482]));
Q_ASSIGN U32293 ( .B(clk), .A(\g.we_clk [481]));
Q_ASSIGN U32294 ( .B(clk), .A(\g.we_clk [480]));
Q_ASSIGN U32295 ( .B(clk), .A(\g.we_clk [479]));
Q_ASSIGN U32296 ( .B(clk), .A(\g.we_clk [478]));
Q_ASSIGN U32297 ( .B(clk), .A(\g.we_clk [477]));
Q_ASSIGN U32298 ( .B(clk), .A(\g.we_clk [476]));
Q_ASSIGN U32299 ( .B(clk), .A(\g.we_clk [475]));
Q_ASSIGN U32300 ( .B(clk), .A(\g.we_clk [474]));
Q_ASSIGN U32301 ( .B(clk), .A(\g.we_clk [473]));
Q_ASSIGN U32302 ( .B(clk), .A(\g.we_clk [472]));
Q_ASSIGN U32303 ( .B(clk), .A(\g.we_clk [471]));
Q_ASSIGN U32304 ( .B(clk), .A(\g.we_clk [470]));
Q_ASSIGN U32305 ( .B(clk), .A(\g.we_clk [469]));
Q_ASSIGN U32306 ( .B(clk), .A(\g.we_clk [468]));
Q_ASSIGN U32307 ( .B(clk), .A(\g.we_clk [467]));
Q_ASSIGN U32308 ( .B(clk), .A(\g.we_clk [466]));
Q_ASSIGN U32309 ( .B(clk), .A(\g.we_clk [465]));
Q_ASSIGN U32310 ( .B(clk), .A(\g.we_clk [464]));
Q_ASSIGN U32311 ( .B(clk), .A(\g.we_clk [463]));
Q_ASSIGN U32312 ( .B(clk), .A(\g.we_clk [462]));
Q_ASSIGN U32313 ( .B(clk), .A(\g.we_clk [461]));
Q_ASSIGN U32314 ( .B(clk), .A(\g.we_clk [460]));
Q_ASSIGN U32315 ( .B(clk), .A(\g.we_clk [459]));
Q_ASSIGN U32316 ( .B(clk), .A(\g.we_clk [458]));
Q_ASSIGN U32317 ( .B(clk), .A(\g.we_clk [457]));
Q_ASSIGN U32318 ( .B(clk), .A(\g.we_clk [456]));
Q_ASSIGN U32319 ( .B(clk), .A(\g.we_clk [455]));
Q_ASSIGN U32320 ( .B(clk), .A(\g.we_clk [454]));
Q_ASSIGN U32321 ( .B(clk), .A(\g.we_clk [453]));
Q_ASSIGN U32322 ( .B(clk), .A(\g.we_clk [452]));
Q_ASSIGN U32323 ( .B(clk), .A(\g.we_clk [451]));
Q_ASSIGN U32324 ( .B(clk), .A(\g.we_clk [450]));
Q_ASSIGN U32325 ( .B(clk), .A(\g.we_clk [449]));
Q_ASSIGN U32326 ( .B(clk), .A(\g.we_clk [448]));
Q_ASSIGN U32327 ( .B(clk), .A(\g.we_clk [447]));
Q_ASSIGN U32328 ( .B(clk), .A(\g.we_clk [446]));
Q_ASSIGN U32329 ( .B(clk), .A(\g.we_clk [445]));
Q_ASSIGN U32330 ( .B(clk), .A(\g.we_clk [444]));
Q_ASSIGN U32331 ( .B(clk), .A(\g.we_clk [443]));
Q_ASSIGN U32332 ( .B(clk), .A(\g.we_clk [442]));
Q_ASSIGN U32333 ( .B(clk), .A(\g.we_clk [441]));
Q_ASSIGN U32334 ( .B(clk), .A(\g.we_clk [440]));
Q_ASSIGN U32335 ( .B(clk), .A(\g.we_clk [439]));
Q_ASSIGN U32336 ( .B(clk), .A(\g.we_clk [438]));
Q_ASSIGN U32337 ( .B(clk), .A(\g.we_clk [437]));
Q_ASSIGN U32338 ( .B(clk), .A(\g.we_clk [436]));
Q_ASSIGN U32339 ( .B(clk), .A(\g.we_clk [435]));
Q_ASSIGN U32340 ( .B(clk), .A(\g.we_clk [434]));
Q_ASSIGN U32341 ( .B(clk), .A(\g.we_clk [433]));
Q_ASSIGN U32342 ( .B(clk), .A(\g.we_clk [432]));
Q_ASSIGN U32343 ( .B(clk), .A(\g.we_clk [431]));
Q_ASSIGN U32344 ( .B(clk), .A(\g.we_clk [430]));
Q_ASSIGN U32345 ( .B(clk), .A(\g.we_clk [429]));
Q_ASSIGN U32346 ( .B(clk), .A(\g.we_clk [428]));
Q_ASSIGN U32347 ( .B(clk), .A(\g.we_clk [427]));
Q_ASSIGN U32348 ( .B(clk), .A(\g.we_clk [426]));
Q_ASSIGN U32349 ( .B(clk), .A(\g.we_clk [425]));
Q_ASSIGN U32350 ( .B(clk), .A(\g.we_clk [424]));
Q_ASSIGN U32351 ( .B(clk), .A(\g.we_clk [423]));
Q_ASSIGN U32352 ( .B(clk), .A(\g.we_clk [422]));
Q_ASSIGN U32353 ( .B(clk), .A(\g.we_clk [421]));
Q_ASSIGN U32354 ( .B(clk), .A(\g.we_clk [420]));
Q_ASSIGN U32355 ( .B(clk), .A(\g.we_clk [419]));
Q_ASSIGN U32356 ( .B(clk), .A(\g.we_clk [418]));
Q_ASSIGN U32357 ( .B(clk), .A(\g.we_clk [417]));
Q_ASSIGN U32358 ( .B(clk), .A(\g.we_clk [416]));
Q_ASSIGN U32359 ( .B(clk), .A(\g.we_clk [415]));
Q_ASSIGN U32360 ( .B(clk), .A(\g.we_clk [414]));
Q_ASSIGN U32361 ( .B(clk), .A(\g.we_clk [413]));
Q_ASSIGN U32362 ( .B(clk), .A(\g.we_clk [412]));
Q_ASSIGN U32363 ( .B(clk), .A(\g.we_clk [411]));
Q_ASSIGN U32364 ( .B(clk), .A(\g.we_clk [410]));
Q_ASSIGN U32365 ( .B(clk), .A(\g.we_clk [409]));
Q_ASSIGN U32366 ( .B(clk), .A(\g.we_clk [408]));
Q_ASSIGN U32367 ( .B(clk), .A(\g.we_clk [407]));
Q_ASSIGN U32368 ( .B(clk), .A(\g.we_clk [406]));
Q_ASSIGN U32369 ( .B(clk), .A(\g.we_clk [405]));
Q_ASSIGN U32370 ( .B(clk), .A(\g.we_clk [404]));
Q_ASSIGN U32371 ( .B(clk), .A(\g.we_clk [403]));
Q_ASSIGN U32372 ( .B(clk), .A(\g.we_clk [402]));
Q_ASSIGN U32373 ( .B(clk), .A(\g.we_clk [401]));
Q_ASSIGN U32374 ( .B(clk), .A(\g.we_clk [400]));
Q_ASSIGN U32375 ( .B(clk), .A(\g.we_clk [399]));
Q_ASSIGN U32376 ( .B(clk), .A(\g.we_clk [398]));
Q_ASSIGN U32377 ( .B(clk), .A(\g.we_clk [397]));
Q_ASSIGN U32378 ( .B(clk), .A(\g.we_clk [396]));
Q_ASSIGN U32379 ( .B(clk), .A(\g.we_clk [395]));
Q_ASSIGN U32380 ( .B(clk), .A(\g.we_clk [394]));
Q_ASSIGN U32381 ( .B(clk), .A(\g.we_clk [393]));
Q_ASSIGN U32382 ( .B(clk), .A(\g.we_clk [392]));
Q_ASSIGN U32383 ( .B(clk), .A(\g.we_clk [391]));
Q_ASSIGN U32384 ( .B(clk), .A(\g.we_clk [390]));
Q_ASSIGN U32385 ( .B(clk), .A(\g.we_clk [389]));
Q_ASSIGN U32386 ( .B(clk), .A(\g.we_clk [388]));
Q_ASSIGN U32387 ( .B(clk), .A(\g.we_clk [387]));
Q_ASSIGN U32388 ( .B(clk), .A(\g.we_clk [386]));
Q_ASSIGN U32389 ( .B(clk), .A(\g.we_clk [385]));
Q_ASSIGN U32390 ( .B(clk), .A(\g.we_clk [384]));
Q_ASSIGN U32391 ( .B(clk), .A(\g.we_clk [383]));
Q_ASSIGN U32392 ( .B(clk), .A(\g.we_clk [382]));
Q_ASSIGN U32393 ( .B(clk), .A(\g.we_clk [381]));
Q_ASSIGN U32394 ( .B(clk), .A(\g.we_clk [380]));
Q_ASSIGN U32395 ( .B(clk), .A(\g.we_clk [379]));
Q_ASSIGN U32396 ( .B(clk), .A(\g.we_clk [378]));
Q_ASSIGN U32397 ( .B(clk), .A(\g.we_clk [377]));
Q_ASSIGN U32398 ( .B(clk), .A(\g.we_clk [376]));
Q_ASSIGN U32399 ( .B(clk), .A(\g.we_clk [375]));
Q_ASSIGN U32400 ( .B(clk), .A(\g.we_clk [374]));
Q_ASSIGN U32401 ( .B(clk), .A(\g.we_clk [373]));
Q_ASSIGN U32402 ( .B(clk), .A(\g.we_clk [372]));
Q_ASSIGN U32403 ( .B(clk), .A(\g.we_clk [371]));
Q_ASSIGN U32404 ( .B(clk), .A(\g.we_clk [370]));
Q_ASSIGN U32405 ( .B(clk), .A(\g.we_clk [369]));
Q_ASSIGN U32406 ( .B(clk), .A(\g.we_clk [368]));
Q_ASSIGN U32407 ( .B(clk), .A(\g.we_clk [367]));
Q_ASSIGN U32408 ( .B(clk), .A(\g.we_clk [366]));
Q_ASSIGN U32409 ( .B(clk), .A(\g.we_clk [365]));
Q_ASSIGN U32410 ( .B(clk), .A(\g.we_clk [364]));
Q_ASSIGN U32411 ( .B(clk), .A(\g.we_clk [363]));
Q_ASSIGN U32412 ( .B(clk), .A(\g.we_clk [362]));
Q_ASSIGN U32413 ( .B(clk), .A(\g.we_clk [361]));
Q_ASSIGN U32414 ( .B(clk), .A(\g.we_clk [360]));
Q_ASSIGN U32415 ( .B(clk), .A(\g.we_clk [359]));
Q_ASSIGN U32416 ( .B(clk), .A(\g.we_clk [358]));
Q_ASSIGN U32417 ( .B(clk), .A(\g.we_clk [357]));
Q_ASSIGN U32418 ( .B(clk), .A(\g.we_clk [356]));
Q_ASSIGN U32419 ( .B(clk), .A(\g.we_clk [355]));
Q_ASSIGN U32420 ( .B(clk), .A(\g.we_clk [354]));
Q_ASSIGN U32421 ( .B(clk), .A(\g.we_clk [353]));
Q_ASSIGN U32422 ( .B(clk), .A(\g.we_clk [352]));
Q_ASSIGN U32423 ( .B(clk), .A(\g.we_clk [351]));
Q_ASSIGN U32424 ( .B(clk), .A(\g.we_clk [350]));
Q_ASSIGN U32425 ( .B(clk), .A(\g.we_clk [349]));
Q_ASSIGN U32426 ( .B(clk), .A(\g.we_clk [348]));
Q_ASSIGN U32427 ( .B(clk), .A(\g.we_clk [347]));
Q_ASSIGN U32428 ( .B(clk), .A(\g.we_clk [346]));
Q_ASSIGN U32429 ( .B(clk), .A(\g.we_clk [345]));
Q_ASSIGN U32430 ( .B(clk), .A(\g.we_clk [344]));
Q_ASSIGN U32431 ( .B(clk), .A(\g.we_clk [343]));
Q_ASSIGN U32432 ( .B(clk), .A(\g.we_clk [342]));
Q_ASSIGN U32433 ( .B(clk), .A(\g.we_clk [341]));
Q_ASSIGN U32434 ( .B(clk), .A(\g.we_clk [340]));
Q_ASSIGN U32435 ( .B(clk), .A(\g.we_clk [339]));
Q_ASSIGN U32436 ( .B(clk), .A(\g.we_clk [338]));
Q_ASSIGN U32437 ( .B(clk), .A(\g.we_clk [337]));
Q_ASSIGN U32438 ( .B(clk), .A(\g.we_clk [336]));
Q_ASSIGN U32439 ( .B(clk), .A(\g.we_clk [335]));
Q_ASSIGN U32440 ( .B(clk), .A(\g.we_clk [334]));
Q_ASSIGN U32441 ( .B(clk), .A(\g.we_clk [333]));
Q_ASSIGN U32442 ( .B(clk), .A(\g.we_clk [332]));
Q_ASSIGN U32443 ( .B(clk), .A(\g.we_clk [331]));
Q_ASSIGN U32444 ( .B(clk), .A(\g.we_clk [330]));
Q_ASSIGN U32445 ( .B(clk), .A(\g.we_clk [329]));
Q_ASSIGN U32446 ( .B(clk), .A(\g.we_clk [328]));
Q_ASSIGN U32447 ( .B(clk), .A(\g.we_clk [327]));
Q_ASSIGN U32448 ( .B(clk), .A(\g.we_clk [326]));
Q_ASSIGN U32449 ( .B(clk), .A(\g.we_clk [325]));
Q_ASSIGN U32450 ( .B(clk), .A(\g.we_clk [324]));
Q_ASSIGN U32451 ( .B(clk), .A(\g.we_clk [323]));
Q_ASSIGN U32452 ( .B(clk), .A(\g.we_clk [322]));
Q_ASSIGN U32453 ( .B(clk), .A(\g.we_clk [321]));
Q_ASSIGN U32454 ( .B(clk), .A(\g.we_clk [320]));
Q_ASSIGN U32455 ( .B(clk), .A(\g.we_clk [319]));
Q_ASSIGN U32456 ( .B(clk), .A(\g.we_clk [318]));
Q_ASSIGN U32457 ( .B(clk), .A(\g.we_clk [317]));
Q_ASSIGN U32458 ( .B(clk), .A(\g.we_clk [316]));
Q_ASSIGN U32459 ( .B(clk), .A(\g.we_clk [315]));
Q_ASSIGN U32460 ( .B(clk), .A(\g.we_clk [314]));
Q_ASSIGN U32461 ( .B(clk), .A(\g.we_clk [313]));
Q_ASSIGN U32462 ( .B(clk), .A(\g.we_clk [312]));
Q_ASSIGN U32463 ( .B(clk), .A(\g.we_clk [311]));
Q_ASSIGN U32464 ( .B(clk), .A(\g.we_clk [310]));
Q_ASSIGN U32465 ( .B(clk), .A(\g.we_clk [309]));
Q_ASSIGN U32466 ( .B(clk), .A(\g.we_clk [308]));
Q_ASSIGN U32467 ( .B(clk), .A(\g.we_clk [307]));
Q_ASSIGN U32468 ( .B(clk), .A(\g.we_clk [306]));
Q_ASSIGN U32469 ( .B(clk), .A(\g.we_clk [305]));
Q_ASSIGN U32470 ( .B(clk), .A(\g.we_clk [304]));
Q_ASSIGN U32471 ( .B(clk), .A(\g.we_clk [303]));
Q_ASSIGN U32472 ( .B(clk), .A(\g.we_clk [302]));
Q_ASSIGN U32473 ( .B(clk), .A(\g.we_clk [301]));
Q_ASSIGN U32474 ( .B(clk), .A(\g.we_clk [300]));
Q_ASSIGN U32475 ( .B(clk), .A(\g.we_clk [299]));
Q_ASSIGN U32476 ( .B(clk), .A(\g.we_clk [298]));
Q_ASSIGN U32477 ( .B(clk), .A(\g.we_clk [297]));
Q_ASSIGN U32478 ( .B(clk), .A(\g.we_clk [296]));
Q_ASSIGN U32479 ( .B(clk), .A(\g.we_clk [295]));
Q_ASSIGN U32480 ( .B(clk), .A(\g.we_clk [294]));
Q_ASSIGN U32481 ( .B(clk), .A(\g.we_clk [293]));
Q_ASSIGN U32482 ( .B(clk), .A(\g.we_clk [292]));
Q_ASSIGN U32483 ( .B(clk), .A(\g.we_clk [291]));
Q_ASSIGN U32484 ( .B(clk), .A(\g.we_clk [290]));
Q_ASSIGN U32485 ( .B(clk), .A(\g.we_clk [289]));
Q_ASSIGN U32486 ( .B(clk), .A(\g.we_clk [288]));
Q_ASSIGN U32487 ( .B(clk), .A(\g.we_clk [287]));
Q_ASSIGN U32488 ( .B(clk), .A(\g.we_clk [286]));
Q_ASSIGN U32489 ( .B(clk), .A(\g.we_clk [285]));
Q_ASSIGN U32490 ( .B(clk), .A(\g.we_clk [284]));
Q_ASSIGN U32491 ( .B(clk), .A(\g.we_clk [283]));
Q_ASSIGN U32492 ( .B(clk), .A(\g.we_clk [282]));
Q_ASSIGN U32493 ( .B(clk), .A(\g.we_clk [281]));
Q_ASSIGN U32494 ( .B(clk), .A(\g.we_clk [280]));
Q_ASSIGN U32495 ( .B(clk), .A(\g.we_clk [279]));
Q_ASSIGN U32496 ( .B(clk), .A(\g.we_clk [278]));
Q_ASSIGN U32497 ( .B(clk), .A(\g.we_clk [277]));
Q_ASSIGN U32498 ( .B(clk), .A(\g.we_clk [276]));
Q_ASSIGN U32499 ( .B(clk), .A(\g.we_clk [275]));
Q_ASSIGN U32500 ( .B(clk), .A(\g.we_clk [274]));
Q_ASSIGN U32501 ( .B(clk), .A(\g.we_clk [273]));
Q_ASSIGN U32502 ( .B(clk), .A(\g.we_clk [272]));
Q_ASSIGN U32503 ( .B(clk), .A(\g.we_clk [271]));
Q_ASSIGN U32504 ( .B(clk), .A(\g.we_clk [270]));
Q_ASSIGN U32505 ( .B(clk), .A(\g.we_clk [269]));
Q_ASSIGN U32506 ( .B(clk), .A(\g.we_clk [268]));
Q_ASSIGN U32507 ( .B(clk), .A(\g.we_clk [267]));
Q_ASSIGN U32508 ( .B(clk), .A(\g.we_clk [266]));
Q_ASSIGN U32509 ( .B(clk), .A(\g.we_clk [265]));
Q_ASSIGN U32510 ( .B(clk), .A(\g.we_clk [264]));
Q_ASSIGN U32511 ( .B(clk), .A(\g.we_clk [263]));
Q_ASSIGN U32512 ( .B(clk), .A(\g.we_clk [262]));
Q_ASSIGN U32513 ( .B(clk), .A(\g.we_clk [261]));
Q_ASSIGN U32514 ( .B(clk), .A(\g.we_clk [260]));
Q_ASSIGN U32515 ( .B(clk), .A(\g.we_clk [259]));
Q_ASSIGN U32516 ( .B(clk), .A(\g.we_clk [258]));
Q_ASSIGN U32517 ( .B(clk), .A(\g.we_clk [257]));
Q_ASSIGN U32518 ( .B(clk), .A(\g.we_clk [256]));
Q_ASSIGN U32519 ( .B(clk), .A(\g.we_clk [255]));
Q_ASSIGN U32520 ( .B(clk), .A(\g.we_clk [254]));
Q_ASSIGN U32521 ( .B(clk), .A(\g.we_clk [253]));
Q_ASSIGN U32522 ( .B(clk), .A(\g.we_clk [252]));
Q_ASSIGN U32523 ( .B(clk), .A(\g.we_clk [251]));
Q_ASSIGN U32524 ( .B(clk), .A(\g.we_clk [250]));
Q_ASSIGN U32525 ( .B(clk), .A(\g.we_clk [249]));
Q_ASSIGN U32526 ( .B(clk), .A(\g.we_clk [248]));
Q_ASSIGN U32527 ( .B(clk), .A(\g.we_clk [247]));
Q_ASSIGN U32528 ( .B(clk), .A(\g.we_clk [246]));
Q_ASSIGN U32529 ( .B(clk), .A(\g.we_clk [245]));
Q_ASSIGN U32530 ( .B(clk), .A(\g.we_clk [244]));
Q_ASSIGN U32531 ( .B(clk), .A(\g.we_clk [243]));
Q_ASSIGN U32532 ( .B(clk), .A(\g.we_clk [242]));
Q_ASSIGN U32533 ( .B(clk), .A(\g.we_clk [241]));
Q_ASSIGN U32534 ( .B(clk), .A(\g.we_clk [240]));
Q_ASSIGN U32535 ( .B(clk), .A(\g.we_clk [239]));
Q_ASSIGN U32536 ( .B(clk), .A(\g.we_clk [238]));
Q_ASSIGN U32537 ( .B(clk), .A(\g.we_clk [237]));
Q_ASSIGN U32538 ( .B(clk), .A(\g.we_clk [236]));
Q_ASSIGN U32539 ( .B(clk), .A(\g.we_clk [235]));
Q_ASSIGN U32540 ( .B(clk), .A(\g.we_clk [234]));
Q_ASSIGN U32541 ( .B(clk), .A(\g.we_clk [233]));
Q_ASSIGN U32542 ( .B(clk), .A(\g.we_clk [232]));
Q_ASSIGN U32543 ( .B(clk), .A(\g.we_clk [231]));
Q_ASSIGN U32544 ( .B(clk), .A(\g.we_clk [230]));
Q_ASSIGN U32545 ( .B(clk), .A(\g.we_clk [229]));
Q_ASSIGN U32546 ( .B(clk), .A(\g.we_clk [228]));
Q_ASSIGN U32547 ( .B(clk), .A(\g.we_clk [227]));
Q_ASSIGN U32548 ( .B(clk), .A(\g.we_clk [226]));
Q_ASSIGN U32549 ( .B(clk), .A(\g.we_clk [225]));
Q_ASSIGN U32550 ( .B(clk), .A(\g.we_clk [224]));
Q_ASSIGN U32551 ( .B(clk), .A(\g.we_clk [223]));
Q_ASSIGN U32552 ( .B(clk), .A(\g.we_clk [222]));
Q_ASSIGN U32553 ( .B(clk), .A(\g.we_clk [221]));
Q_ASSIGN U32554 ( .B(clk), .A(\g.we_clk [220]));
Q_ASSIGN U32555 ( .B(clk), .A(\g.we_clk [219]));
Q_ASSIGN U32556 ( .B(clk), .A(\g.we_clk [218]));
Q_ASSIGN U32557 ( .B(clk), .A(\g.we_clk [217]));
Q_ASSIGN U32558 ( .B(clk), .A(\g.we_clk [216]));
Q_ASSIGN U32559 ( .B(clk), .A(\g.we_clk [215]));
Q_ASSIGN U32560 ( .B(clk), .A(\g.we_clk [214]));
Q_ASSIGN U32561 ( .B(clk), .A(\g.we_clk [213]));
Q_ASSIGN U32562 ( .B(clk), .A(\g.we_clk [212]));
Q_ASSIGN U32563 ( .B(clk), .A(\g.we_clk [211]));
Q_ASSIGN U32564 ( .B(clk), .A(\g.we_clk [210]));
Q_ASSIGN U32565 ( .B(clk), .A(\g.we_clk [209]));
Q_ASSIGN U32566 ( .B(clk), .A(\g.we_clk [208]));
Q_ASSIGN U32567 ( .B(clk), .A(\g.we_clk [207]));
Q_ASSIGN U32568 ( .B(clk), .A(\g.we_clk [206]));
Q_ASSIGN U32569 ( .B(clk), .A(\g.we_clk [205]));
Q_ASSIGN U32570 ( .B(clk), .A(\g.we_clk [204]));
Q_ASSIGN U32571 ( .B(clk), .A(\g.we_clk [203]));
Q_ASSIGN U32572 ( .B(clk), .A(\g.we_clk [202]));
Q_ASSIGN U32573 ( .B(clk), .A(\g.we_clk [201]));
Q_ASSIGN U32574 ( .B(clk), .A(\g.we_clk [200]));
Q_ASSIGN U32575 ( .B(clk), .A(\g.we_clk [199]));
Q_ASSIGN U32576 ( .B(clk), .A(\g.we_clk [198]));
Q_ASSIGN U32577 ( .B(clk), .A(\g.we_clk [197]));
Q_ASSIGN U32578 ( .B(clk), .A(\g.we_clk [196]));
Q_ASSIGN U32579 ( .B(clk), .A(\g.we_clk [195]));
Q_ASSIGN U32580 ( .B(clk), .A(\g.we_clk [194]));
Q_ASSIGN U32581 ( .B(clk), .A(\g.we_clk [193]));
Q_ASSIGN U32582 ( .B(clk), .A(\g.we_clk [192]));
Q_ASSIGN U32583 ( .B(clk), .A(\g.we_clk [191]));
Q_ASSIGN U32584 ( .B(clk), .A(\g.we_clk [190]));
Q_ASSIGN U32585 ( .B(clk), .A(\g.we_clk [189]));
Q_ASSIGN U32586 ( .B(clk), .A(\g.we_clk [188]));
Q_ASSIGN U32587 ( .B(clk), .A(\g.we_clk [187]));
Q_ASSIGN U32588 ( .B(clk), .A(\g.we_clk [186]));
Q_ASSIGN U32589 ( .B(clk), .A(\g.we_clk [185]));
Q_ASSIGN U32590 ( .B(clk), .A(\g.we_clk [184]));
Q_ASSIGN U32591 ( .B(clk), .A(\g.we_clk [183]));
Q_ASSIGN U32592 ( .B(clk), .A(\g.we_clk [182]));
Q_ASSIGN U32593 ( .B(clk), .A(\g.we_clk [181]));
Q_ASSIGN U32594 ( .B(clk), .A(\g.we_clk [180]));
Q_ASSIGN U32595 ( .B(clk), .A(\g.we_clk [179]));
Q_ASSIGN U32596 ( .B(clk), .A(\g.we_clk [178]));
Q_ASSIGN U32597 ( .B(clk), .A(\g.we_clk [177]));
Q_ASSIGN U32598 ( .B(clk), .A(\g.we_clk [176]));
Q_ASSIGN U32599 ( .B(clk), .A(\g.we_clk [175]));
Q_ASSIGN U32600 ( .B(clk), .A(\g.we_clk [174]));
Q_ASSIGN U32601 ( .B(clk), .A(\g.we_clk [173]));
Q_ASSIGN U32602 ( .B(clk), .A(\g.we_clk [172]));
Q_ASSIGN U32603 ( .B(clk), .A(\g.we_clk [171]));
Q_ASSIGN U32604 ( .B(clk), .A(\g.we_clk [170]));
Q_ASSIGN U32605 ( .B(clk), .A(\g.we_clk [169]));
Q_ASSIGN U32606 ( .B(clk), .A(\g.we_clk [168]));
Q_ASSIGN U32607 ( .B(clk), .A(\g.we_clk [167]));
Q_ASSIGN U32608 ( .B(clk), .A(\g.we_clk [166]));
Q_ASSIGN U32609 ( .B(clk), .A(\g.we_clk [165]));
Q_ASSIGN U32610 ( .B(clk), .A(\g.we_clk [164]));
Q_ASSIGN U32611 ( .B(clk), .A(\g.we_clk [163]));
Q_ASSIGN U32612 ( .B(clk), .A(\g.we_clk [162]));
Q_ASSIGN U32613 ( .B(clk), .A(\g.we_clk [161]));
Q_ASSIGN U32614 ( .B(clk), .A(\g.we_clk [160]));
Q_ASSIGN U32615 ( .B(clk), .A(\g.we_clk [159]));
Q_ASSIGN U32616 ( .B(clk), .A(\g.we_clk [158]));
Q_ASSIGN U32617 ( .B(clk), .A(\g.we_clk [157]));
Q_ASSIGN U32618 ( .B(clk), .A(\g.we_clk [156]));
Q_ASSIGN U32619 ( .B(clk), .A(\g.we_clk [155]));
Q_ASSIGN U32620 ( .B(clk), .A(\g.we_clk [154]));
Q_ASSIGN U32621 ( .B(clk), .A(\g.we_clk [153]));
Q_ASSIGN U32622 ( .B(clk), .A(\g.we_clk [152]));
Q_ASSIGN U32623 ( .B(clk), .A(\g.we_clk [151]));
Q_ASSIGN U32624 ( .B(clk), .A(\g.we_clk [150]));
Q_ASSIGN U32625 ( .B(clk), .A(\g.we_clk [149]));
Q_ASSIGN U32626 ( .B(clk), .A(\g.we_clk [148]));
Q_ASSIGN U32627 ( .B(clk), .A(\g.we_clk [147]));
Q_ASSIGN U32628 ( .B(clk), .A(\g.we_clk [146]));
Q_ASSIGN U32629 ( .B(clk), .A(\g.we_clk [145]));
Q_ASSIGN U32630 ( .B(clk), .A(\g.we_clk [144]));
Q_ASSIGN U32631 ( .B(clk), .A(\g.we_clk [143]));
Q_ASSIGN U32632 ( .B(clk), .A(\g.we_clk [142]));
Q_ASSIGN U32633 ( .B(clk), .A(\g.we_clk [141]));
Q_ASSIGN U32634 ( .B(clk), .A(\g.we_clk [140]));
Q_ASSIGN U32635 ( .B(clk), .A(\g.we_clk [139]));
Q_ASSIGN U32636 ( .B(clk), .A(\g.we_clk [138]));
Q_ASSIGN U32637 ( .B(clk), .A(\g.we_clk [137]));
Q_ASSIGN U32638 ( .B(clk), .A(\g.we_clk [136]));
Q_ASSIGN U32639 ( .B(clk), .A(\g.we_clk [135]));
Q_ASSIGN U32640 ( .B(clk), .A(\g.we_clk [134]));
Q_ASSIGN U32641 ( .B(clk), .A(\g.we_clk [133]));
Q_ASSIGN U32642 ( .B(clk), .A(\g.we_clk [132]));
Q_ASSIGN U32643 ( .B(clk), .A(\g.we_clk [131]));
Q_ASSIGN U32644 ( .B(clk), .A(\g.we_clk [130]));
Q_ASSIGN U32645 ( .B(clk), .A(\g.we_clk [129]));
Q_ASSIGN U32646 ( .B(clk), .A(\g.we_clk [128]));
Q_ASSIGN U32647 ( .B(clk), .A(\g.we_clk [127]));
Q_ASSIGN U32648 ( .B(clk), .A(\g.we_clk [126]));
Q_ASSIGN U32649 ( .B(clk), .A(\g.we_clk [125]));
Q_ASSIGN U32650 ( .B(clk), .A(\g.we_clk [124]));
Q_ASSIGN U32651 ( .B(clk), .A(\g.we_clk [123]));
Q_ASSIGN U32652 ( .B(clk), .A(\g.we_clk [122]));
Q_ASSIGN U32653 ( .B(clk), .A(\g.we_clk [121]));
Q_ASSIGN U32654 ( .B(clk), .A(\g.we_clk [120]));
Q_ASSIGN U32655 ( .B(clk), .A(\g.we_clk [119]));
Q_ASSIGN U32656 ( .B(clk), .A(\g.we_clk [118]));
Q_ASSIGN U32657 ( .B(clk), .A(\g.we_clk [117]));
Q_ASSIGN U32658 ( .B(clk), .A(\g.we_clk [116]));
Q_ASSIGN U32659 ( .B(clk), .A(\g.we_clk [115]));
Q_ASSIGN U32660 ( .B(clk), .A(\g.we_clk [114]));
Q_ASSIGN U32661 ( .B(clk), .A(\g.we_clk [113]));
Q_ASSIGN U32662 ( .B(clk), .A(\g.we_clk [112]));
Q_ASSIGN U32663 ( .B(clk), .A(\g.we_clk [111]));
Q_ASSIGN U32664 ( .B(clk), .A(\g.we_clk [110]));
Q_ASSIGN U32665 ( .B(clk), .A(\g.we_clk [109]));
Q_ASSIGN U32666 ( .B(clk), .A(\g.we_clk [108]));
Q_ASSIGN U32667 ( .B(clk), .A(\g.we_clk [107]));
Q_ASSIGN U32668 ( .B(clk), .A(\g.we_clk [106]));
Q_ASSIGN U32669 ( .B(clk), .A(\g.we_clk [105]));
Q_ASSIGN U32670 ( .B(clk), .A(\g.we_clk [104]));
Q_ASSIGN U32671 ( .B(clk), .A(\g.we_clk [103]));
Q_ASSIGN U32672 ( .B(clk), .A(\g.we_clk [102]));
Q_ASSIGN U32673 ( .B(clk), .A(\g.we_clk [101]));
Q_ASSIGN U32674 ( .B(clk), .A(\g.we_clk [100]));
Q_ASSIGN U32675 ( .B(clk), .A(\g.we_clk [99]));
Q_ASSIGN U32676 ( .B(clk), .A(\g.we_clk [98]));
Q_ASSIGN U32677 ( .B(clk), .A(\g.we_clk [97]));
Q_ASSIGN U32678 ( .B(clk), .A(\g.we_clk [96]));
Q_ASSIGN U32679 ( .B(clk), .A(\g.we_clk [95]));
Q_ASSIGN U32680 ( .B(clk), .A(\g.we_clk [94]));
Q_ASSIGN U32681 ( .B(clk), .A(\g.we_clk [93]));
Q_ASSIGN U32682 ( .B(clk), .A(\g.we_clk [92]));
Q_ASSIGN U32683 ( .B(clk), .A(\g.we_clk [91]));
Q_ASSIGN U32684 ( .B(clk), .A(\g.we_clk [90]));
Q_ASSIGN U32685 ( .B(clk), .A(\g.we_clk [89]));
Q_ASSIGN U32686 ( .B(clk), .A(\g.we_clk [88]));
Q_ASSIGN U32687 ( .B(clk), .A(\g.we_clk [87]));
Q_ASSIGN U32688 ( .B(clk), .A(\g.we_clk [86]));
Q_ASSIGN U32689 ( .B(clk), .A(\g.we_clk [85]));
Q_ASSIGN U32690 ( .B(clk), .A(\g.we_clk [84]));
Q_ASSIGN U32691 ( .B(clk), .A(\g.we_clk [83]));
Q_ASSIGN U32692 ( .B(clk), .A(\g.we_clk [82]));
Q_ASSIGN U32693 ( .B(clk), .A(\g.we_clk [81]));
Q_ASSIGN U32694 ( .B(clk), .A(\g.we_clk [80]));
Q_ASSIGN U32695 ( .B(clk), .A(\g.we_clk [79]));
Q_ASSIGN U32696 ( .B(clk), .A(\g.we_clk [78]));
Q_ASSIGN U32697 ( .B(clk), .A(\g.we_clk [77]));
Q_ASSIGN U32698 ( .B(clk), .A(\g.we_clk [76]));
Q_ASSIGN U32699 ( .B(clk), .A(\g.we_clk [75]));
Q_ASSIGN U32700 ( .B(clk), .A(\g.we_clk [74]));
Q_ASSIGN U32701 ( .B(clk), .A(\g.we_clk [73]));
Q_ASSIGN U32702 ( .B(clk), .A(\g.we_clk [72]));
Q_ASSIGN U32703 ( .B(clk), .A(\g.we_clk [71]));
Q_ASSIGN U32704 ( .B(clk), .A(\g.we_clk [70]));
Q_ASSIGN U32705 ( .B(clk), .A(\g.we_clk [69]));
Q_ASSIGN U32706 ( .B(clk), .A(\g.we_clk [68]));
Q_ASSIGN U32707 ( .B(clk), .A(\g.we_clk [67]));
Q_ASSIGN U32708 ( .B(clk), .A(\g.we_clk [66]));
Q_ASSIGN U32709 ( .B(clk), .A(\g.we_clk [65]));
Q_ASSIGN U32710 ( .B(clk), .A(\g.we_clk [64]));
Q_ASSIGN U32711 ( .B(clk), .A(\g.we_clk [63]));
Q_ASSIGN U32712 ( .B(clk), .A(\g.we_clk [62]));
Q_ASSIGN U32713 ( .B(clk), .A(\g.we_clk [61]));
Q_ASSIGN U32714 ( .B(clk), .A(\g.we_clk [60]));
Q_ASSIGN U32715 ( .B(clk), .A(\g.we_clk [59]));
Q_ASSIGN U32716 ( .B(clk), .A(\g.we_clk [58]));
Q_ASSIGN U32717 ( .B(clk), .A(\g.we_clk [57]));
Q_ASSIGN U32718 ( .B(clk), .A(\g.we_clk [56]));
Q_ASSIGN U32719 ( .B(clk), .A(\g.we_clk [55]));
Q_ASSIGN U32720 ( .B(clk), .A(\g.we_clk [54]));
Q_ASSIGN U32721 ( .B(clk), .A(\g.we_clk [53]));
Q_ASSIGN U32722 ( .B(clk), .A(\g.we_clk [52]));
Q_ASSIGN U32723 ( .B(clk), .A(\g.we_clk [51]));
Q_ASSIGN U32724 ( .B(clk), .A(\g.we_clk [50]));
Q_ASSIGN U32725 ( .B(clk), .A(\g.we_clk [49]));
Q_ASSIGN U32726 ( .B(clk), .A(\g.we_clk [48]));
Q_ASSIGN U32727 ( .B(clk), .A(\g.we_clk [47]));
Q_ASSIGN U32728 ( .B(clk), .A(\g.we_clk [46]));
Q_ASSIGN U32729 ( .B(clk), .A(\g.we_clk [45]));
Q_ASSIGN U32730 ( .B(clk), .A(\g.we_clk [44]));
Q_ASSIGN U32731 ( .B(clk), .A(\g.we_clk [43]));
Q_ASSIGN U32732 ( .B(clk), .A(\g.we_clk [42]));
Q_ASSIGN U32733 ( .B(clk), .A(\g.we_clk [41]));
Q_ASSIGN U32734 ( .B(clk), .A(\g.we_clk [40]));
Q_ASSIGN U32735 ( .B(clk), .A(\g.we_clk [39]));
Q_ASSIGN U32736 ( .B(clk), .A(\g.we_clk [38]));
Q_ASSIGN U32737 ( .B(clk), .A(\g.we_clk [37]));
Q_ASSIGN U32738 ( .B(clk), .A(\g.we_clk [36]));
Q_ASSIGN U32739 ( .B(clk), .A(\g.we_clk [35]));
Q_ASSIGN U32740 ( .B(clk), .A(\g.we_clk [34]));
Q_ASSIGN U32741 ( .B(clk), .A(\g.we_clk [33]));
Q_ASSIGN U32742 ( .B(clk), .A(\g.we_clk [32]));
Q_ASSIGN U32743 ( .B(clk), .A(\g.we_clk [31]));
Q_ASSIGN U32744 ( .B(clk), .A(\g.we_clk [30]));
Q_ASSIGN U32745 ( .B(clk), .A(\g.we_clk [29]));
Q_ASSIGN U32746 ( .B(clk), .A(\g.we_clk [28]));
Q_ASSIGN U32747 ( .B(clk), .A(\g.we_clk [27]));
Q_ASSIGN U32748 ( .B(clk), .A(\g.we_clk [26]));
Q_ASSIGN U32749 ( .B(clk), .A(\g.we_clk [25]));
Q_ASSIGN U32750 ( .B(clk), .A(\g.we_clk [24]));
Q_ASSIGN U32751 ( .B(clk), .A(\g.we_clk [23]));
Q_ASSIGN U32752 ( .B(clk), .A(\g.we_clk [22]));
Q_ASSIGN U32753 ( .B(clk), .A(\g.we_clk [21]));
Q_ASSIGN U32754 ( .B(clk), .A(\g.we_clk [20]));
Q_ASSIGN U32755 ( .B(clk), .A(\g.we_clk [19]));
Q_ASSIGN U32756 ( .B(clk), .A(\g.we_clk [18]));
Q_ASSIGN U32757 ( .B(clk), .A(\g.we_clk [17]));
Q_ASSIGN U32758 ( .B(clk), .A(\g.we_clk [16]));
Q_ASSIGN U32759 ( .B(clk), .A(\g.we_clk [15]));
Q_ASSIGN U32760 ( .B(clk), .A(\g.we_clk [14]));
Q_ASSIGN U32761 ( .B(clk), .A(\g.we_clk [13]));
Q_ASSIGN U32762 ( .B(clk), .A(\g.we_clk [12]));
Q_ASSIGN U32763 ( .B(clk), .A(\g.we_clk [11]));
Q_ASSIGN U32764 ( .B(clk), .A(\g.we_clk [10]));
Q_ASSIGN U32765 ( .B(clk), .A(\g.we_clk [9]));
Q_ASSIGN U32766 ( .B(clk), .A(\g.we_clk [8]));
Q_ASSIGN U32767 ( .B(clk), .A(\g.we_clk [7]));
Q_ASSIGN U32768 ( .B(clk), .A(\g.we_clk [6]));
Q_ASSIGN U32769 ( .B(clk), .A(\g.we_clk [5]));
Q_ASSIGN U32770 ( .B(clk), .A(\g.we_clk [4]));
Q_ASSIGN U32771 ( .B(clk), .A(\g.we_clk [3]));
Q_ASSIGN U32772 ( .B(clk), .A(\g.we_clk [2]));
Q_ASSIGN U32773 ( .B(clk), .A(\g.we_clk [1]));
Q_ASSIGN U32774 ( .B(clk), .A(\g.we_clk [0]));
Q_BUF U32775 ( .A(n217), .Z(ro_uncorrectable_ecc_error));
ixc_assign _zz_strnp_10 ( _zy_simnet_ro_uncorrectable_ecc_error_2_w$, n217);
ixc_assign _zz_strnp_9 ( _zy_simnet_bimc_osync_1_w$, bimc_osync);
ixc_assign _zz_strnp_8 ( _zy_simnet_bimc_odat_0_w$, bimc_odat);
Q_INV U32779 ( .A(n216), .Z(web));
Q_AN02 U32780 ( .A0(cs), .A1(we), .Z(n216));
ixc_assign _zz_strnp_7 ( rst_rclk_n, rst_n);
ixc_assign _zz_strnp_6 ( rst_clk_n, rst_n);
ixc_assign _zz_strnp_5 ( bimc_irstn, bimc_rst_n);
ixc_assign _zz_strnp_4 ( bimc_iclk, clk);
Q_FDP0 U32785 ( .CK(clk), .D(\g.din_i [63]), .Q(n215), .QN( ));
Q_FDP0 U32786 ( .CK(clk), .D(\g.din_i [62]), .Q(n214), .QN( ));
Q_FDP0 U32787 ( .CK(clk), .D(\g.din_i [61]), .Q(n213), .QN( ));
Q_FDP0 U32788 ( .CK(clk), .D(\g.din_i [60]), .Q(n212), .QN( ));
Q_FDP0 U32789 ( .CK(clk), .D(\g.din_i [59]), .Q(n211), .QN( ));
Q_FDP0 U32790 ( .CK(clk), .D(\g.din_i [58]), .Q(n210), .QN( ));
Q_FDP0 U32791 ( .CK(clk), .D(\g.din_i [57]), .Q(n209), .QN( ));
Q_FDP0 U32792 ( .CK(clk), .D(\g.din_i [56]), .Q(n208), .QN( ));
Q_FDP0 U32793 ( .CK(clk), .D(\g.din_i [55]), .Q(n207), .QN( ));
Q_FDP0 U32794 ( .CK(clk), .D(\g.din_i [54]), .Q(n206), .QN( ));
Q_FDP0 U32795 ( .CK(clk), .D(\g.din_i [53]), .Q(n205), .QN( ));
Q_FDP0 U32796 ( .CK(clk), .D(\g.din_i [52]), .Q(n204), .QN( ));
Q_FDP0 U32797 ( .CK(clk), .D(\g.din_i [51]), .Q(n203), .QN( ));
Q_FDP0 U32798 ( .CK(clk), .D(\g.din_i [50]), .Q(n202), .QN( ));
Q_FDP0 U32799 ( .CK(clk), .D(\g.din_i [49]), .Q(n201), .QN( ));
Q_FDP0 U32800 ( .CK(clk), .D(\g.din_i [48]), .Q(n200), .QN( ));
Q_FDP0 U32801 ( .CK(clk), .D(\g.din_i [47]), .Q(n199), .QN( ));
Q_FDP0 U32802 ( .CK(clk), .D(\g.din_i [46]), .Q(n198), .QN( ));
Q_FDP0 U32803 ( .CK(clk), .D(\g.din_i [45]), .Q(n197), .QN( ));
Q_FDP0 U32804 ( .CK(clk), .D(\g.din_i [44]), .Q(n196), .QN( ));
Q_FDP0 U32805 ( .CK(clk), .D(\g.din_i [43]), .Q(n195), .QN( ));
Q_FDP0 U32806 ( .CK(clk), .D(\g.din_i [42]), .Q(n194), .QN( ));
Q_FDP0 U32807 ( .CK(clk), .D(\g.din_i [41]), .Q(n193), .QN( ));
Q_FDP0 U32808 ( .CK(clk), .D(\g.din_i [40]), .Q(n192), .QN( ));
Q_FDP0 U32809 ( .CK(clk), .D(\g.din_i [39]), .Q(n191), .QN( ));
Q_FDP0 U32810 ( .CK(clk), .D(\g.din_i [38]), .Q(n190), .QN( ));
Q_FDP0 U32811 ( .CK(clk), .D(\g.din_i [37]), .Q(n189), .QN( ));
Q_FDP0 U32812 ( .CK(clk), .D(\g.din_i [36]), .Q(n188), .QN( ));
Q_FDP0 U32813 ( .CK(clk), .D(\g.din_i [35]), .Q(n187), .QN( ));
Q_FDP0 U32814 ( .CK(clk), .D(\g.din_i [34]), .Q(n186), .QN( ));
Q_FDP0 U32815 ( .CK(clk), .D(\g.din_i [33]), .Q(n185), .QN( ));
Q_FDP0 U32816 ( .CK(clk), .D(\g.din_i [32]), .Q(n184), .QN( ));
Q_FDP0 U32817 ( .CK(clk), .D(\g.din_i [31]), .Q(n183), .QN( ));
Q_FDP0 U32818 ( .CK(clk), .D(\g.din_i [30]), .Q(n182), .QN( ));
Q_FDP0 U32819 ( .CK(clk), .D(\g.din_i [29]), .Q(n181), .QN( ));
Q_FDP0 U32820 ( .CK(clk), .D(\g.din_i [28]), .Q(n180), .QN( ));
Q_FDP0 U32821 ( .CK(clk), .D(\g.din_i [27]), .Q(n179), .QN( ));
Q_FDP0 U32822 ( .CK(clk), .D(\g.din_i [26]), .Q(n178), .QN( ));
Q_FDP0 U32823 ( .CK(clk), .D(\g.din_i [25]), .Q(n177), .QN( ));
Q_FDP0 U32824 ( .CK(clk), .D(\g.din_i [24]), .Q(n176), .QN( ));
Q_FDP0 U32825 ( .CK(clk), .D(\g.din_i [23]), .Q(n175), .QN( ));
Q_FDP0 U32826 ( .CK(clk), .D(\g.din_i [22]), .Q(n174), .QN( ));
Q_FDP0 U32827 ( .CK(clk), .D(\g.din_i [21]), .Q(n173), .QN( ));
Q_FDP0 U32828 ( .CK(clk), .D(\g.din_i [20]), .Q(n172), .QN( ));
Q_FDP0 U32829 ( .CK(clk), .D(\g.din_i [19]), .Q(n171), .QN( ));
Q_FDP0 U32830 ( .CK(clk), .D(\g.din_i [18]), .Q(n170), .QN( ));
Q_FDP0 U32831 ( .CK(clk), .D(\g.din_i [17]), .Q(n169), .QN( ));
Q_FDP0 U32832 ( .CK(clk), .D(\g.din_i [16]), .Q(n168), .QN( ));
Q_FDP0 U32833 ( .CK(clk), .D(\g.din_i [15]), .Q(n167), .QN( ));
Q_FDP0 U32834 ( .CK(clk), .D(\g.din_i [14]), .Q(n166), .QN( ));
Q_FDP0 U32835 ( .CK(clk), .D(\g.din_i [13]), .Q(n165), .QN( ));
Q_FDP0 U32836 ( .CK(clk), .D(\g.din_i [12]), .Q(n164), .QN( ));
Q_FDP0 U32837 ( .CK(clk), .D(\g.din_i [11]), .Q(n163), .QN( ));
Q_FDP0 U32838 ( .CK(clk), .D(\g.din_i [10]), .Q(n162), .QN( ));
Q_FDP0 U32839 ( .CK(clk), .D(\g.din_i [9]), .Q(n161), .QN( ));
Q_FDP0 U32840 ( .CK(clk), .D(\g.din_i [8]), .Q(n160), .QN( ));
Q_FDP0 U32841 ( .CK(clk), .D(\g.din_i [7]), .Q(n159), .QN( ));
Q_FDP0 U32842 ( .CK(clk), .D(\g.din_i [6]), .Q(n158), .QN( ));
Q_FDP0 U32843 ( .CK(clk), .D(\g.din_i [5]), .Q(n157), .QN( ));
Q_FDP0 U32844 ( .CK(clk), .D(\g.din_i [4]), .Q(n156), .QN( ));
Q_FDP0 U32845 ( .CK(clk), .D(\g.din_i [3]), .Q(n155), .QN( ));
Q_FDP0 U32846 ( .CK(clk), .D(\g.din_i [2]), .Q(n154), .QN( ));
Q_FDP0 U32847 ( .CK(clk), .D(\g.din_i [1]), .Q(n153), .QN( ));
Q_FDP0 U32848 ( .CK(clk), .D(\g.din_i [0]), .Q(n152), .QN( ));
Q_FDP0 U32849 ( .CK(clk), .D(add[14]), .Q(n151), .QN( ));
Q_FDP0 U32850 ( .CK(clk), .D(add[13]), .Q(n150), .QN( ));
Q_FDP0 U32851 ( .CK(clk), .D(add[12]), .Q(n149), .QN( ));
Q_FDP0 U32852 ( .CK(clk), .D(add[11]), .Q(n148), .QN( ));
Q_FDP0 U32853 ( .CK(clk), .D(add[10]), .Q(n147), .QN( ));
Q_FDP0 U32854 ( .CK(clk), .D(add[9]), .Q(n146), .QN( ));
Q_FDP0 U32855 ( .CK(clk), .D(add[8]), .Q(n145), .QN( ));
Q_FDP0 U32856 ( .CK(clk), .D(add[7]), .Q(n144), .QN( ));
Q_FDP0 U32857 ( .CK(clk), .D(add[6]), .Q(n143), .QN( ));
Q_FDP0 U32858 ( .CK(clk), .D(add[5]), .Q(n142), .QN( ));
Q_FDP0 U32859 ( .CK(clk), .D(add[4]), .Q(n141), .QN( ));
Q_FDP0 U32860 ( .CK(clk), .D(add[3]), .Q(n140), .QN( ));
Q_FDP0 U32861 ( .CK(clk), .D(add[2]), .Q(n139), .QN( ));
Q_FDP0 U32862 ( .CK(clk), .D(add[1]), .Q(n138), .QN( ));
Q_FDP0 U32863 ( .CK(clk), .D(add[0]), .Q(n137), .QN( ));
Q_AN02 U32864 ( .A0(n132), .A1(n135), .Z(n136));
Q_XOR2 U32865 ( .A0(n131), .A1(n134), .Z(n135));
// pragma CVAINTPROP NET n131 _2_state_ 1
// pragma CVAINTPROP INSTANCE U32865 NOBREAKS 1
Q_FDP0B U32866 ( .D(n131), .QTFCLK( ), .Q(n134));
Q_FDP0 U32867 ( .CK(clk), .D(n216), .Q(n132), .QN( ));
Q_FDP0 U32868 ( .CK(clk), .D(n133), .Q(n131), .QN(n133));
Q_MX02 U32869 ( .S(we), .A0(\g.dout_i [63]), .A1(\g.din_i [63]), .Z(n130));
Q_MX02 U32870 ( .S(we), .A0(\g.dout_i [62]), .A1(\g.din_i [62]), .Z(n129));
Q_MX02 U32871 ( .S(we), .A0(\g.dout_i [61]), .A1(\g.din_i [61]), .Z(n128));
Q_MX02 U32872 ( .S(we), .A0(\g.dout_i [60]), .A1(\g.din_i [60]), .Z(n127));
Q_MX02 U32873 ( .S(we), .A0(\g.dout_i [59]), .A1(\g.din_i [59]), .Z(n126));
Q_MX02 U32874 ( .S(we), .A0(\g.dout_i [58]), .A1(\g.din_i [58]), .Z(n125));
Q_MX02 U32875 ( .S(we), .A0(\g.dout_i [57]), .A1(\g.din_i [57]), .Z(n124));
Q_MX02 U32876 ( .S(we), .A0(\g.dout_i [56]), .A1(\g.din_i [56]), .Z(n123));
Q_MX02 U32877 ( .S(we), .A0(\g.dout_i [55]), .A1(\g.din_i [55]), .Z(n122));
Q_MX02 U32878 ( .S(we), .A0(\g.dout_i [54]), .A1(\g.din_i [54]), .Z(n121));
Q_MX02 U32879 ( .S(we), .A0(\g.dout_i [53]), .A1(\g.din_i [53]), .Z(n120));
Q_MX02 U32880 ( .S(we), .A0(\g.dout_i [52]), .A1(\g.din_i [52]), .Z(n119));
Q_MX02 U32881 ( .S(we), .A0(\g.dout_i [51]), .A1(\g.din_i [51]), .Z(n118));
Q_MX02 U32882 ( .S(we), .A0(\g.dout_i [50]), .A1(\g.din_i [50]), .Z(n117));
Q_MX02 U32883 ( .S(we), .A0(\g.dout_i [49]), .A1(\g.din_i [49]), .Z(n116));
Q_MX02 U32884 ( .S(we), .A0(\g.dout_i [48]), .A1(\g.din_i [48]), .Z(n115));
Q_MX02 U32885 ( .S(we), .A0(\g.dout_i [47]), .A1(\g.din_i [47]), .Z(n114));
Q_MX02 U32886 ( .S(we), .A0(\g.dout_i [46]), .A1(\g.din_i [46]), .Z(n113));
Q_MX02 U32887 ( .S(we), .A0(\g.dout_i [45]), .A1(\g.din_i [45]), .Z(n112));
Q_MX02 U32888 ( .S(we), .A0(\g.dout_i [44]), .A1(\g.din_i [44]), .Z(n111));
Q_MX02 U32889 ( .S(we), .A0(\g.dout_i [43]), .A1(\g.din_i [43]), .Z(n110));
Q_MX02 U32890 ( .S(we), .A0(\g.dout_i [42]), .A1(\g.din_i [42]), .Z(n109));
Q_MX02 U32891 ( .S(we), .A0(\g.dout_i [41]), .A1(\g.din_i [41]), .Z(n108));
Q_MX02 U32892 ( .S(we), .A0(\g.dout_i [40]), .A1(\g.din_i [40]), .Z(n107));
Q_MX02 U32893 ( .S(we), .A0(\g.dout_i [39]), .A1(\g.din_i [39]), .Z(n106));
Q_MX02 U32894 ( .S(we), .A0(\g.dout_i [38]), .A1(\g.din_i [38]), .Z(n105));
Q_MX02 U32895 ( .S(we), .A0(\g.dout_i [37]), .A1(\g.din_i [37]), .Z(n104));
Q_MX02 U32896 ( .S(we), .A0(\g.dout_i [36]), .A1(\g.din_i [36]), .Z(n103));
Q_MX02 U32897 ( .S(we), .A0(\g.dout_i [35]), .A1(\g.din_i [35]), .Z(n102));
Q_MX02 U32898 ( .S(we), .A0(\g.dout_i [34]), .A1(\g.din_i [34]), .Z(n101));
Q_MX02 U32899 ( .S(we), .A0(\g.dout_i [33]), .A1(\g.din_i [33]), .Z(n100));
Q_MX02 U32900 ( .S(we), .A0(\g.dout_i [32]), .A1(\g.din_i [32]), .Z(n99));
Q_MX02 U32901 ( .S(we), .A0(\g.dout_i [31]), .A1(\g.din_i [31]), .Z(n98));
Q_MX02 U32902 ( .S(we), .A0(\g.dout_i [30]), .A1(\g.din_i [30]), .Z(n97));
Q_MX02 U32903 ( .S(we), .A0(\g.dout_i [29]), .A1(\g.din_i [29]), .Z(n96));
Q_MX02 U32904 ( .S(we), .A0(\g.dout_i [28]), .A1(\g.din_i [28]), .Z(n95));
Q_MX02 U32905 ( .S(we), .A0(\g.dout_i [27]), .A1(\g.din_i [27]), .Z(n94));
Q_MX02 U32906 ( .S(we), .A0(\g.dout_i [26]), .A1(\g.din_i [26]), .Z(n93));
Q_MX02 U32907 ( .S(we), .A0(\g.dout_i [25]), .A1(\g.din_i [25]), .Z(n92));
Q_MX02 U32908 ( .S(we), .A0(\g.dout_i [24]), .A1(\g.din_i [24]), .Z(n91));
Q_MX02 U32909 ( .S(we), .A0(\g.dout_i [23]), .A1(\g.din_i [23]), .Z(n90));
Q_MX02 U32910 ( .S(we), .A0(\g.dout_i [22]), .A1(\g.din_i [22]), .Z(n89));
Q_MX02 U32911 ( .S(we), .A0(\g.dout_i [21]), .A1(\g.din_i [21]), .Z(n88));
Q_MX02 U32912 ( .S(we), .A0(\g.dout_i [20]), .A1(\g.din_i [20]), .Z(n87));
Q_MX02 U32913 ( .S(we), .A0(\g.dout_i [19]), .A1(\g.din_i [19]), .Z(n86));
Q_MX02 U32914 ( .S(we), .A0(\g.dout_i [18]), .A1(\g.din_i [18]), .Z(n85));
Q_MX02 U32915 ( .S(we), .A0(\g.dout_i [17]), .A1(\g.din_i [17]), .Z(n84));
Q_MX02 U32916 ( .S(we), .A0(\g.dout_i [16]), .A1(\g.din_i [16]), .Z(n83));
Q_MX02 U32917 ( .S(we), .A0(\g.dout_i [15]), .A1(\g.din_i [15]), .Z(n82));
Q_MX02 U32918 ( .S(we), .A0(\g.dout_i [14]), .A1(\g.din_i [14]), .Z(n81));
Q_MX02 U32919 ( .S(we), .A0(\g.dout_i [13]), .A1(\g.din_i [13]), .Z(n80));
Q_MX02 U32920 ( .S(we), .A0(\g.dout_i [12]), .A1(\g.din_i [12]), .Z(n79));
Q_MX02 U32921 ( .S(we), .A0(\g.dout_i [11]), .A1(\g.din_i [11]), .Z(n78));
Q_MX02 U32922 ( .S(we), .A0(\g.dout_i [10]), .A1(\g.din_i [10]), .Z(n77));
Q_MX02 U32923 ( .S(we), .A0(\g.dout_i [9]), .A1(\g.din_i [9]), .Z(n76));
Q_MX02 U32924 ( .S(we), .A0(\g.dout_i [8]), .A1(\g.din_i [8]), .Z(n75));
Q_MX02 U32925 ( .S(we), .A0(\g.dout_i [7]), .A1(\g.din_i [7]), .Z(n74));
Q_MX02 U32926 ( .S(we), .A0(\g.dout_i [6]), .A1(\g.din_i [6]), .Z(n73));
Q_MX02 U32927 ( .S(we), .A0(\g.dout_i [5]), .A1(\g.din_i [5]), .Z(n72));
Q_MX02 U32928 ( .S(we), .A0(\g.dout_i [4]), .A1(\g.din_i [4]), .Z(n71));
Q_MX02 U32929 ( .S(we), .A0(\g.dout_i [3]), .A1(\g.din_i [3]), .Z(n70));
Q_MX02 U32930 ( .S(we), .A0(\g.dout_i [2]), .A1(\g.din_i [2]), .Z(n69));
Q_MX02 U32931 ( .S(we), .A0(\g.dout_i [1]), .A1(\g.din_i [1]), .Z(n68));
Q_MX02 U32932 ( .S(we), .A0(\g.dout_i [0]), .A1(\g.din_i [0]), .Z(n67));
ixc_assign_64 \g._zz_strnp_0 ( \g.dout_i [63:0], { n66, n65, n64, n63, n62, 
	n61, n60, n59, n58, n57, n56, n55, n54, n53, n52, n51, n50, n49, n48, 
	n47, n46, n45, n44, n43, n42, n41, n40, n39, n38, n37, n36, n35, n34, 
	n33, n32, n31, n30, n29, n28, n27, n26, n25, n24, n23, n22, n21, n20, 
	n19, n18, n17, n16, n15, n14, n13, n12, n11, n10, n9, n8, n7, n6, n5, 
	n4, n3});
ixc_assign \g._zz_strnp_3 ( bimc_osync, bimc_isync);
ixc_assign \g._zz_strnp_2 ( bimc_odat, bimc_idat);
ixc_assign_64 \g._zz_strnp_1 ( dout[63:0], \g.dat_r [63:0]);
Q_MX02 U32937 ( .S(bwe[63]), .A0(\g.dout_i [63]), .A1(din[63]), .Z(\g.din_i [63]));
Q_MX02 U32938 ( .S(bwe[62]), .A0(\g.dout_i [62]), .A1(din[62]), .Z(\g.din_i [62]));
Q_MX02 U32939 ( .S(bwe[61]), .A0(\g.dout_i [61]), .A1(din[61]), .Z(\g.din_i [61]));
Q_MX02 U32940 ( .S(bwe[60]), .A0(\g.dout_i [60]), .A1(din[60]), .Z(\g.din_i [60]));
Q_MX02 U32941 ( .S(bwe[59]), .A0(\g.dout_i [59]), .A1(din[59]), .Z(\g.din_i [59]));
Q_MX02 U32942 ( .S(bwe[58]), .A0(\g.dout_i [58]), .A1(din[58]), .Z(\g.din_i [58]));
Q_MX02 U32943 ( .S(bwe[57]), .A0(\g.dout_i [57]), .A1(din[57]), .Z(\g.din_i [57]));
Q_MX02 U32944 ( .S(bwe[56]), .A0(\g.dout_i [56]), .A1(din[56]), .Z(\g.din_i [56]));
Q_MX02 U32945 ( .S(bwe[55]), .A0(\g.dout_i [55]), .A1(din[55]), .Z(\g.din_i [55]));
Q_MX02 U32946 ( .S(bwe[54]), .A0(\g.dout_i [54]), .A1(din[54]), .Z(\g.din_i [54]));
Q_MX02 U32947 ( .S(bwe[53]), .A0(\g.dout_i [53]), .A1(din[53]), .Z(\g.din_i [53]));
Q_MX02 U32948 ( .S(bwe[52]), .A0(\g.dout_i [52]), .A1(din[52]), .Z(\g.din_i [52]));
Q_MX02 U32949 ( .S(bwe[51]), .A0(\g.dout_i [51]), .A1(din[51]), .Z(\g.din_i [51]));
Q_MX02 U32950 ( .S(bwe[50]), .A0(\g.dout_i [50]), .A1(din[50]), .Z(\g.din_i [50]));
Q_MX02 U32951 ( .S(bwe[49]), .A0(\g.dout_i [49]), .A1(din[49]), .Z(\g.din_i [49]));
Q_MX02 U32952 ( .S(bwe[48]), .A0(\g.dout_i [48]), .A1(din[48]), .Z(\g.din_i [48]));
Q_MX02 U32953 ( .S(bwe[47]), .A0(\g.dout_i [47]), .A1(din[47]), .Z(\g.din_i [47]));
Q_MX02 U32954 ( .S(bwe[46]), .A0(\g.dout_i [46]), .A1(din[46]), .Z(\g.din_i [46]));
Q_MX02 U32955 ( .S(bwe[45]), .A0(\g.dout_i [45]), .A1(din[45]), .Z(\g.din_i [45]));
Q_MX02 U32956 ( .S(bwe[44]), .A0(\g.dout_i [44]), .A1(din[44]), .Z(\g.din_i [44]));
Q_MX02 U32957 ( .S(bwe[43]), .A0(\g.dout_i [43]), .A1(din[43]), .Z(\g.din_i [43]));
Q_MX02 U32958 ( .S(bwe[42]), .A0(\g.dout_i [42]), .A1(din[42]), .Z(\g.din_i [42]));
Q_MX02 U32959 ( .S(bwe[41]), .A0(\g.dout_i [41]), .A1(din[41]), .Z(\g.din_i [41]));
Q_MX02 U32960 ( .S(bwe[40]), .A0(\g.dout_i [40]), .A1(din[40]), .Z(\g.din_i [40]));
Q_MX02 U32961 ( .S(bwe[39]), .A0(\g.dout_i [39]), .A1(din[39]), .Z(\g.din_i [39]));
Q_MX02 U32962 ( .S(bwe[38]), .A0(\g.dout_i [38]), .A1(din[38]), .Z(\g.din_i [38]));
Q_MX02 U32963 ( .S(bwe[37]), .A0(\g.dout_i [37]), .A1(din[37]), .Z(\g.din_i [37]));
Q_MX02 U32964 ( .S(bwe[36]), .A0(\g.dout_i [36]), .A1(din[36]), .Z(\g.din_i [36]));
Q_MX02 U32965 ( .S(bwe[35]), .A0(\g.dout_i [35]), .A1(din[35]), .Z(\g.din_i [35]));
Q_MX02 U32966 ( .S(bwe[34]), .A0(\g.dout_i [34]), .A1(din[34]), .Z(\g.din_i [34]));
Q_MX02 U32967 ( .S(bwe[33]), .A0(\g.dout_i [33]), .A1(din[33]), .Z(\g.din_i [33]));
Q_MX02 U32968 ( .S(bwe[32]), .A0(\g.dout_i [32]), .A1(din[32]), .Z(\g.din_i [32]));
Q_MX02 U32969 ( .S(bwe[31]), .A0(\g.dout_i [31]), .A1(din[31]), .Z(\g.din_i [31]));
Q_MX02 U32970 ( .S(bwe[30]), .A0(\g.dout_i [30]), .A1(din[30]), .Z(\g.din_i [30]));
Q_MX02 U32971 ( .S(bwe[29]), .A0(\g.dout_i [29]), .A1(din[29]), .Z(\g.din_i [29]));
Q_MX02 U32972 ( .S(bwe[28]), .A0(\g.dout_i [28]), .A1(din[28]), .Z(\g.din_i [28]));
Q_MX02 U32973 ( .S(bwe[27]), .A0(\g.dout_i [27]), .A1(din[27]), .Z(\g.din_i [27]));
Q_MX02 U32974 ( .S(bwe[26]), .A0(\g.dout_i [26]), .A1(din[26]), .Z(\g.din_i [26]));
Q_MX02 U32975 ( .S(bwe[25]), .A0(\g.dout_i [25]), .A1(din[25]), .Z(\g.din_i [25]));
Q_MX02 U32976 ( .S(bwe[24]), .A0(\g.dout_i [24]), .A1(din[24]), .Z(\g.din_i [24]));
Q_MX02 U32977 ( .S(bwe[23]), .A0(\g.dout_i [23]), .A1(din[23]), .Z(\g.din_i [23]));
Q_MX02 U32978 ( .S(bwe[22]), .A0(\g.dout_i [22]), .A1(din[22]), .Z(\g.din_i [22]));
Q_MX02 U32979 ( .S(bwe[21]), .A0(\g.dout_i [21]), .A1(din[21]), .Z(\g.din_i [21]));
Q_MX02 U32980 ( .S(bwe[20]), .A0(\g.dout_i [20]), .A1(din[20]), .Z(\g.din_i [20]));
Q_MX02 U32981 ( .S(bwe[19]), .A0(\g.dout_i [19]), .A1(din[19]), .Z(\g.din_i [19]));
Q_MX02 U32982 ( .S(bwe[18]), .A0(\g.dout_i [18]), .A1(din[18]), .Z(\g.din_i [18]));
Q_MX02 U32983 ( .S(bwe[17]), .A0(\g.dout_i [17]), .A1(din[17]), .Z(\g.din_i [17]));
Q_MX02 U32984 ( .S(bwe[16]), .A0(\g.dout_i [16]), .A1(din[16]), .Z(\g.din_i [16]));
Q_MX02 U32985 ( .S(bwe[15]), .A0(\g.dout_i [15]), .A1(din[15]), .Z(\g.din_i [15]));
Q_MX02 U32986 ( .S(bwe[14]), .A0(\g.dout_i [14]), .A1(din[14]), .Z(\g.din_i [14]));
Q_MX02 U32987 ( .S(bwe[13]), .A0(\g.dout_i [13]), .A1(din[13]), .Z(\g.din_i [13]));
Q_MX02 U32988 ( .S(bwe[12]), .A0(\g.dout_i [12]), .A1(din[12]), .Z(\g.din_i [12]));
Q_MX02 U32989 ( .S(bwe[11]), .A0(\g.dout_i [11]), .A1(din[11]), .Z(\g.din_i [11]));
Q_MX02 U32990 ( .S(bwe[10]), .A0(\g.dout_i [10]), .A1(din[10]), .Z(\g.din_i [10]));
Q_MX02 U32991 ( .S(bwe[9]), .A0(\g.dout_i [9]), .A1(din[9]), .Z(\g.din_i [9]));
Q_MX02 U32992 ( .S(bwe[8]), .A0(\g.dout_i [8]), .A1(din[8]), .Z(\g.din_i [8]));
Q_MX02 U32993 ( .S(bwe[7]), .A0(\g.dout_i [7]), .A1(din[7]), .Z(\g.din_i [7]));
Q_MX02 U32994 ( .S(bwe[6]), .A0(\g.dout_i [6]), .A1(din[6]), .Z(\g.din_i [6]));
Q_MX02 U32995 ( .S(bwe[5]), .A0(\g.dout_i [5]), .A1(din[5]), .Z(\g.din_i [5]));
Q_MX02 U32996 ( .S(bwe[4]), .A0(\g.dout_i [4]), .A1(din[4]), .Z(\g.din_i [4]));
Q_MX02 U32997 ( .S(bwe[3]), .A0(\g.dout_i [3]), .A1(din[3]), .Z(\g.din_i [3]));
Q_MX02 U32998 ( .S(bwe[2]), .A0(\g.dout_i [2]), .A1(din[2]), .Z(\g.din_i [2]));
Q_MX02 U32999 ( .S(bwe[1]), .A0(\g.dout_i [1]), .A1(din[1]), .Z(\g.din_i [1]));
Q_MX02 U33000 ( .S(bwe[0]), .A0(\g.dout_i [0]), .A1(din[0]), .Z(\g.din_i [0]));
Q_FDP4EP \g.dat_r_REG[63] ( .CK(clk), .CE(cs), .R(n1), .D(n130), .Q(\g.dat_r [63]));
Q_INV U33002 ( .A(rst_n), .Z(n1));
Q_FDP4EP \g.dat_r_REG[62] ( .CK(clk), .CE(cs), .R(n1), .D(n129), .Q(\g.dat_r [62]));
Q_FDP4EP \g.dat_r_REG[61] ( .CK(clk), .CE(cs), .R(n1), .D(n128), .Q(\g.dat_r [61]));
Q_FDP4EP \g.dat_r_REG[60] ( .CK(clk), .CE(cs), .R(n1), .D(n127), .Q(\g.dat_r [60]));
Q_FDP4EP \g.dat_r_REG[59] ( .CK(clk), .CE(cs), .R(n1), .D(n126), .Q(\g.dat_r [59]));
Q_FDP4EP \g.dat_r_REG[58] ( .CK(clk), .CE(cs), .R(n1), .D(n125), .Q(\g.dat_r [58]));
Q_FDP4EP \g.dat_r_REG[57] ( .CK(clk), .CE(cs), .R(n1), .D(n124), .Q(\g.dat_r [57]));
Q_FDP4EP \g.dat_r_REG[56] ( .CK(clk), .CE(cs), .R(n1), .D(n123), .Q(\g.dat_r [56]));
Q_FDP4EP \g.dat_r_REG[55] ( .CK(clk), .CE(cs), .R(n1), .D(n122), .Q(\g.dat_r [55]));
Q_FDP4EP \g.dat_r_REG[54] ( .CK(clk), .CE(cs), .R(n1), .D(n121), .Q(\g.dat_r [54]));
Q_FDP4EP \g.dat_r_REG[53] ( .CK(clk), .CE(cs), .R(n1), .D(n120), .Q(\g.dat_r [53]));
Q_FDP4EP \g.dat_r_REG[52] ( .CK(clk), .CE(cs), .R(n1), .D(n119), .Q(\g.dat_r [52]));
Q_FDP4EP \g.dat_r_REG[51] ( .CK(clk), .CE(cs), .R(n1), .D(n118), .Q(\g.dat_r [51]));
Q_FDP4EP \g.dat_r_REG[50] ( .CK(clk), .CE(cs), .R(n1), .D(n117), .Q(\g.dat_r [50]));
Q_FDP4EP \g.dat_r_REG[49] ( .CK(clk), .CE(cs), .R(n1), .D(n116), .Q(\g.dat_r [49]));
Q_FDP4EP \g.dat_r_REG[48] ( .CK(clk), .CE(cs), .R(n1), .D(n115), .Q(\g.dat_r [48]));
Q_FDP4EP \g.dat_r_REG[47] ( .CK(clk), .CE(cs), .R(n1), .D(n114), .Q(\g.dat_r [47]));
Q_FDP4EP \g.dat_r_REG[46] ( .CK(clk), .CE(cs), .R(n1), .D(n113), .Q(\g.dat_r [46]));
Q_FDP4EP \g.dat_r_REG[45] ( .CK(clk), .CE(cs), .R(n1), .D(n112), .Q(\g.dat_r [45]));
Q_FDP4EP \g.dat_r_REG[44] ( .CK(clk), .CE(cs), .R(n1), .D(n111), .Q(\g.dat_r [44]));
Q_FDP4EP \g.dat_r_REG[43] ( .CK(clk), .CE(cs), .R(n1), .D(n110), .Q(\g.dat_r [43]));
Q_FDP4EP \g.dat_r_REG[42] ( .CK(clk), .CE(cs), .R(n1), .D(n109), .Q(\g.dat_r [42]));
Q_FDP4EP \g.dat_r_REG[41] ( .CK(clk), .CE(cs), .R(n1), .D(n108), .Q(\g.dat_r [41]));
Q_FDP4EP \g.dat_r_REG[40] ( .CK(clk), .CE(cs), .R(n1), .D(n107), .Q(\g.dat_r [40]));
Q_FDP4EP \g.dat_r_REG[39] ( .CK(clk), .CE(cs), .R(n1), .D(n106), .Q(\g.dat_r [39]));
Q_FDP4EP \g.dat_r_REG[38] ( .CK(clk), .CE(cs), .R(n1), .D(n105), .Q(\g.dat_r [38]));
Q_FDP4EP \g.dat_r_REG[37] ( .CK(clk), .CE(cs), .R(n1), .D(n104), .Q(\g.dat_r [37]));
Q_FDP4EP \g.dat_r_REG[36] ( .CK(clk), .CE(cs), .R(n1), .D(n103), .Q(\g.dat_r [36]));
Q_FDP4EP \g.dat_r_REG[35] ( .CK(clk), .CE(cs), .R(n1), .D(n102), .Q(\g.dat_r [35]));
Q_FDP4EP \g.dat_r_REG[34] ( .CK(clk), .CE(cs), .R(n1), .D(n101), .Q(\g.dat_r [34]));
Q_FDP4EP \g.dat_r_REG[33] ( .CK(clk), .CE(cs), .R(n1), .D(n100), .Q(\g.dat_r [33]));
Q_FDP4EP \g.dat_r_REG[32] ( .CK(clk), .CE(cs), .R(n1), .D(n99), .Q(\g.dat_r [32]));
Q_FDP4EP \g.dat_r_REG[31] ( .CK(clk), .CE(cs), .R(n1), .D(n98), .Q(\g.dat_r [31]));
Q_FDP4EP \g.dat_r_REG[30] ( .CK(clk), .CE(cs), .R(n1), .D(n97), .Q(\g.dat_r [30]));
Q_FDP4EP \g.dat_r_REG[29] ( .CK(clk), .CE(cs), .R(n1), .D(n96), .Q(\g.dat_r [29]));
Q_FDP4EP \g.dat_r_REG[28] ( .CK(clk), .CE(cs), .R(n1), .D(n95), .Q(\g.dat_r [28]));
Q_FDP4EP \g.dat_r_REG[27] ( .CK(clk), .CE(cs), .R(n1), .D(n94), .Q(\g.dat_r [27]));
Q_FDP4EP \g.dat_r_REG[26] ( .CK(clk), .CE(cs), .R(n1), .D(n93), .Q(\g.dat_r [26]));
Q_FDP4EP \g.dat_r_REG[25] ( .CK(clk), .CE(cs), .R(n1), .D(n92), .Q(\g.dat_r [25]));
Q_FDP4EP \g.dat_r_REG[24] ( .CK(clk), .CE(cs), .R(n1), .D(n91), .Q(\g.dat_r [24]));
Q_FDP4EP \g.dat_r_REG[23] ( .CK(clk), .CE(cs), .R(n1), .D(n90), .Q(\g.dat_r [23]));
Q_FDP4EP \g.dat_r_REG[22] ( .CK(clk), .CE(cs), .R(n1), .D(n89), .Q(\g.dat_r [22]));
Q_FDP4EP \g.dat_r_REG[21] ( .CK(clk), .CE(cs), .R(n1), .D(n88), .Q(\g.dat_r [21]));
Q_FDP4EP \g.dat_r_REG[20] ( .CK(clk), .CE(cs), .R(n1), .D(n87), .Q(\g.dat_r [20]));
Q_FDP4EP \g.dat_r_REG[19] ( .CK(clk), .CE(cs), .R(n1), .D(n86), .Q(\g.dat_r [19]));
Q_FDP4EP \g.dat_r_REG[18] ( .CK(clk), .CE(cs), .R(n1), .D(n85), .Q(\g.dat_r [18]));
Q_FDP4EP \g.dat_r_REG[17] ( .CK(clk), .CE(cs), .R(n1), .D(n84), .Q(\g.dat_r [17]));
Q_FDP4EP \g.dat_r_REG[16] ( .CK(clk), .CE(cs), .R(n1), .D(n83), .Q(\g.dat_r [16]));
Q_FDP4EP \g.dat_r_REG[15] ( .CK(clk), .CE(cs), .R(n1), .D(n82), .Q(\g.dat_r [15]));
Q_FDP4EP \g.dat_r_REG[14] ( .CK(clk), .CE(cs), .R(n1), .D(n81), .Q(\g.dat_r [14]));
Q_FDP4EP \g.dat_r_REG[13] ( .CK(clk), .CE(cs), .R(n1), .D(n80), .Q(\g.dat_r [13]));
Q_FDP4EP \g.dat_r_REG[12] ( .CK(clk), .CE(cs), .R(n1), .D(n79), .Q(\g.dat_r [12]));
Q_FDP4EP \g.dat_r_REG[11] ( .CK(clk), .CE(cs), .R(n1), .D(n78), .Q(\g.dat_r [11]));
Q_FDP4EP \g.dat_r_REG[10] ( .CK(clk), .CE(cs), .R(n1), .D(n77), .Q(\g.dat_r [10]));
Q_FDP4EP \g.dat_r_REG[9] ( .CK(clk), .CE(cs), .R(n1), .D(n76), .Q(\g.dat_r [9]));
Q_FDP4EP \g.dat_r_REG[8] ( .CK(clk), .CE(cs), .R(n1), .D(n75), .Q(\g.dat_r [8]));
Q_FDP4EP \g.dat_r_REG[7] ( .CK(clk), .CE(cs), .R(n1), .D(n74), .Q(\g.dat_r [7]));
Q_FDP4EP \g.dat_r_REG[6] ( .CK(clk), .CE(cs), .R(n1), .D(n73), .Q(\g.dat_r [6]));
Q_FDP4EP \g.dat_r_REG[5] ( .CK(clk), .CE(cs), .R(n1), .D(n72), .Q(\g.dat_r [5]));
Q_FDP4EP \g.dat_r_REG[4] ( .CK(clk), .CE(cs), .R(n1), .D(n71), .Q(\g.dat_r [4]));
Q_FDP4EP \g.dat_r_REG[3] ( .CK(clk), .CE(cs), .R(n1), .D(n70), .Q(\g.dat_r [3]));
Q_FDP4EP \g.dat_r_REG[2] ( .CK(clk), .CE(cs), .R(n1), .D(n69), .Q(\g.dat_r [2]));
Q_FDP4EP \g.dat_r_REG[1] ( .CK(clk), .CE(cs), .R(n1), .D(n68), .Q(\g.dat_r [1]));
Q_FDP4EP \g.dat_r_REG[0] ( .CK(clk), .CE(cs), .R(n1), .D(n67), .Q(\g.dat_r [0]));
`ifdef CBV

reg [63:0] \g.mem  [0:32767];
initial begin: U33066
  integer i;
  for (i=0; i<=32767; i=i+1) \g.mem [i] =
`ifdef CBV_MEM_INIT1
  {64{1'b1}};
`else
  64'b0;
`endif
end
reg [63:0] n218;
assign {n66, n65, n64, n63, n62, n61, n60,
n59, n58, n57, n56, n55, n54, n53, n52,
n51, n50, n49, n48, n47, n46, n45, n44,
n43, n42, n41, n40, n39, n38, n37, n36,
n35, n34, n33, n32, n31, n30, n29, n28,
n27, n26, n25, n24, n23, n22, n21, n20,
n19, n18, n17, n16, n15, n14, n13, n12,
n11, n10, n9, n8, n7, n6, n5, n4,
n3} = n218; 
always @(n151 or n150 or n149 or n148 or n147
 or n146 or n145 or n144 or n143 or n142 or n141 or n140 or n139
 or n138 or n137 or n215 or n214 or n213 or n212 or n211 or n210
 or n209 or n208 or n207 or n206 or n205 or n204 or n203 or n202
 or n201 or n200 or n199 or n198 or n197 or n196 or n195 or n194
 or n193 or n192 or n191 or n190 or n189 or n188 or n187 or n186
 or n185 or n184 or n183 or n182 or n181 or n180 or n179 or n178
 or n177 or n176 or n175 or n174 or n173 or n172 or n171 or n170
 or n169 or n168 or n167 or n166 or n165 or n164 or n163 or n162
 or n161 or n160 or n159 or n158 or n157 or n156 or n155 or n154
 or n153 or n152 or n136 or add[14] or add[13] or add[12] or add[11] or add[10]
 or add[9] or add[8] or add[7] or add[6] or add[5] or add[4] or add[3] or add[2]
 or add[1] or add[0])
#0 begin
if (n136)
\g.mem [{n151, n150, n149, n148, n147,
 n146, n145, n144, n143, n142, n141, n140, n139,
 n138, n137}] =
{n215, n214, n213, n212, n211,
 n210, n209, n208, n207, n206, n205, n204, n203,
 n202, n201, n200, n199, n198, n197, n196, n195,
 n194, n193, n192, n191, n190, n189, n188, n187,
 n186, n185, n184, n183, n182, n181, n180, n179,
 n178, n177, n176, n175, n174, n173, n172, n171,
 n170, n169, n168, n167, n166, n165, n164, n163,
 n162, n161, n160, n159, n158, n157, n156, n155,
 n154, n153, n152};
n218 = \g.mem [{add[14], add[13], add[12], add[11], add[10],
 add[9], add[8], add[7], add[6], add[5], add[4], add[3], add[2],
 add[1], add[0]}];
end
`else

MPW32KX64 \g.mem  ( .A14(n151), .A13(n150), .A12(n149), .A11(n148), .A10(n147), .A9(n146),
 .A8(n145), .A7(n144), .A6(n143), .A5(n142), .A4(n141), .A3(n140), .A2(n139), .A1(n138),
 .A0(n137), .DI63(n215), .DI62(n214), .DI61(n213), .DI60(n212), .DI59(n211), .DI58(n210), .DI57(n209),
 .DI56(n208), .DI55(n207), .DI54(n206), .DI53(n205), .DI52(n204), .DI51(n203), .DI50(n202), .DI49(n201),
 .DI48(n200), .DI47(n199), .DI46(n198), .DI45(n197), .DI44(n196), .DI43(n195), .DI42(n194), .DI41(n193),
 .DI40(n192), .DI39(n191), .DI38(n190), .DI37(n189), .DI36(n188), .DI35(n187), .DI34(n186), .DI33(n185),
 .DI32(n184), .DI31(n183), .DI30(n182), .DI29(n181), .DI28(n180), .DI27(n179), .DI26(n178), .DI25(n177),
 .DI24(n176), .DI23(n175), .DI22(n174), .DI21(n173), .DI20(n172), .DI19(n171), .DI18(n170), .DI17(n169),
 .DI16(n168), .DI15(n167), .DI14(n166), .DI13(n165), .DI12(n164), .DI11(n163), .DI10(n162), .DI9(n161),
 .DI8(n160), .DI7(n159), .DI6(n158), .DI5(n157), .DI4(n156), .DI3(n155), .DI2(n154), .DI1(n153),
 .DI0(n152), .WE(n136), .SYNC_IN(n217), .SYNC_OUT(n218));
// pragma CVASTRPROP INSTANCE "\g.mem " HDL_MEMORY_DECL "1 63 0 0 32767"
MPR32KX64 U33067 ( .A14(add[14]), .A13(add[13]), .A12(add[12]), .A11(add[11]), .A10(add[10]), .A9(add[9]),
 .A8(add[8]), .A7(add[7]), .A6(add[6]), .A5(add[5]), .A4(add[4]), .A3(add[3]), .A2(add[2]), .A1(add[1]),
 .A0(add[0]), .SYNC_IN(n218), .DO63(n66), .DO62(n65), .DO61(n64), .DO60(n63), .DO59(n62), .DO58(n61),
 .DO57(n60), .DO56(n59), .DO55(n58), .DO54(n57), .DO53(n56), .DO52(n55), .DO51(n54), .DO50(n53),
 .DO49(n52), .DO48(n51), .DO47(n50), .DO46(n49), .DO45(n48), .DO44(n47), .DO43(n46), .DO42(n45),
 .DO41(n44), .DO40(n43), .DO39(n42), .DO38(n41), .DO37(n40), .DO36(n39), .DO35(n38), .DO34(n37),
 .DO33(n36), .DO32(n35), .DO31(n34), .DO30(n33), .DO29(n32), .DO28(n31), .DO27(n30), .DO26(n29),
 .DO25(n28), .DO24(n27), .DO23(n26), .DO22(n25), .DO21(n24), .DO20(n23), .DO19(n22), .DO18(n21),
 .DO17(n20), .DO16(n19), .DO15(n18), .DO14(n17), .DO13(n16), .DO12(n15), .DO11(n14), .DO10(n13),
 .DO9(n12), .DO8(n11), .DO7(n10), .DO6(n9), .DO5(n8), .DO4(n7), .DO3(n6), .DO2(n5),
 .DO1(n4), .DO0(n3), .SYNC_OUT( ));
`endif
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_1 "0 u_ram  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_0 "-1 g  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "g.u_ram"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "g"
endmodule
`ifdef CBV
`else
`ifdef MPW32KX64_MPR32KX64
`else
module MPW32KX64( A14, A13, A12, A11, A10, A9, A8,
 A7, A6, A5, A4, A3, A2, A1, A0,
 DI63, DI62, DI61, DI60, DI59, DI58, DI57, DI56,
 DI55, DI54, DI53, DI52, DI51, DI50, DI49, DI48,
 DI47, DI46, DI45, DI44, DI43, DI42, DI41, DI40,
 DI39, DI38, DI37, DI36, DI35, DI34, DI33, DI32,
 DI31, DI30, DI29, DI28, DI27, DI26, DI25, DI24,
 DI23, DI22, DI21, DI20, DI19, DI18, DI17, DI16,
 DI15, DI14, DI13, DI12, DI11, DI10, DI9, DI8,
 DI7, DI6, DI5, DI4, DI3, DI2, DI1, DI0,
 WE, SYNC_IN, SYNC_OUT);
input  A14, A13, A12, A11, A10, A9, A8, A7,
 A6, A5, A4, A3, A2, A1, A0, DI63, DI62, DI61,
 DI60, DI59, DI58, DI57, DI56, DI55, DI54, DI53, DI52, DI51,
 DI50, DI49, DI48, DI47, DI46, DI45, DI44, DI43, DI42, DI41,
 DI40, DI39, DI38, DI37, DI36, DI35, DI34, DI33, DI32, DI31,
 DI30, DI29, DI28, DI27, DI26, DI25, DI24, DI23, DI22, DI21,
 DI20, DI19, DI18, DI17, DI16, DI15, DI14, DI13, DI12, DI11,
 DI10, DI9, DI8, DI7, DI6, DI5, DI4, DI3, DI2, DI1,
 DI0, WE, SYNC_IN;
output  SYNC_OUT;
endmodule
`ifdef _MPR32KX64_
`else
module MPR32KX64( A14, A13, A12, A11, A10, A9, A8,
 A7, A6, A5, A4, A3, A2, A1, A0,
 SYNC_IN, DO63, DO62, DO61, DO60, DO59, DO58, DO57,
 DO56, DO55, DO54, DO53, DO52, DO51, DO50, DO49,
 DO48, DO47, DO46, DO45, DO44, DO43, DO42, DO41,
 DO40, DO39, DO38, DO37, DO36, DO35, DO34, DO33,
 DO32, DO31, DO30, DO29, DO28, DO27, DO26, DO25,
 DO24, DO23, DO22, DO21, DO20, DO19, DO18, DO17,
 DO16, DO15, DO14, DO13, DO12, DO11, DO10, DO9,
 DO8, DO7, DO6, DO5, DO4, DO3, DO2, DO1,
 DO0, SYNC_OUT);
input  A14, A13, A12, A11, A10, A9, A8, A7,
 A6, A5, A4, A3, A2, A1, A0, SYNC_IN;
output  DO63, DO62, DO61, DO60, DO59, DO58, DO57, DO56,
 DO55, DO54, DO53, DO52, DO51, DO50, DO49, DO48, DO47, DO46,
 DO45, DO44, DO43, DO42, DO41, DO40, DO39, DO38, DO37, DO36,
 DO35, DO34, DO33, DO32, DO31, DO30, DO29, DO28, DO27, DO26,
 DO25, DO24, DO23, DO22, DO21, DO20, DO19, DO18, DO17, DO16,
 DO15, DO14, DO13, DO12, DO11, DO10, DO9, DO8, DO7, DO6,
 DO5, DO4, DO3, DO2, DO1, DO0, SYNC_OUT;
endmodule
`define _MPR32KX64_
`endif
`define MPW32KX64_MPR32KX64
`endif
`endif
