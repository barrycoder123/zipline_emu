
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module cr_kme_kop_xcm67 ( kme_internal_out_ack, key_tlv_ob_wr, .key_tlv_ob_tlv( {
	\key_tlv_ob_tlv.insert , \key_tlv_ob_tlv.ordern [12], 
	\key_tlv_ob_tlv.ordern [11], \key_tlv_ob_tlv.ordern [10], 
	\key_tlv_ob_tlv.ordern [9], \key_tlv_ob_tlv.ordern [8], 
	\key_tlv_ob_tlv.ordern [7], \key_tlv_ob_tlv.ordern [6], 
	\key_tlv_ob_tlv.ordern [5], \key_tlv_ob_tlv.ordern [4], 
	\key_tlv_ob_tlv.ordern [3], \key_tlv_ob_tlv.ordern [2], 
	\key_tlv_ob_tlv.ordern [1], \key_tlv_ob_tlv.ordern [0], 
	\key_tlv_ob_tlv.typen [7], \key_tlv_ob_tlv.typen [6], 
	\key_tlv_ob_tlv.typen [5], \key_tlv_ob_tlv.typen [4], 
	\key_tlv_ob_tlv.typen [3], \key_tlv_ob_tlv.typen [2], 
	\key_tlv_ob_tlv.typen [1], \key_tlv_ob_tlv.typen [0], 
	\key_tlv_ob_tlv.sot , \key_tlv_ob_tlv.eot , \key_tlv_ob_tlv.tlast , 
	\key_tlv_ob_tlv.tid [0], \key_tlv_ob_tlv.tstrb [7], 
	\key_tlv_ob_tlv.tstrb [6], \key_tlv_ob_tlv.tstrb [5], 
	\key_tlv_ob_tlv.tstrb [4], \key_tlv_ob_tlv.tstrb [3], 
	\key_tlv_ob_tlv.tstrb [2], \key_tlv_ob_tlv.tstrb [1], 
	\key_tlv_ob_tlv.tstrb [0], \key_tlv_ob_tlv.tuser [7], 
	\key_tlv_ob_tlv.tuser [6], \key_tlv_ob_tlv.tuser [5], 
	\key_tlv_ob_tlv.tuser [4], \key_tlv_ob_tlv.tuser [3], 
	\key_tlv_ob_tlv.tuser [2], \key_tlv_ob_tlv.tuser [1], 
	\key_tlv_ob_tlv.tuser [0], \key_tlv_ob_tlv.tdata [63], 
	\key_tlv_ob_tlv.tdata [62], \key_tlv_ob_tlv.tdata [61], 
	\key_tlv_ob_tlv.tdata [60], \key_tlv_ob_tlv.tdata [59], 
	\key_tlv_ob_tlv.tdata [58], \key_tlv_ob_tlv.tdata [57], 
	\key_tlv_ob_tlv.tdata [56], \key_tlv_ob_tlv.tdata [55], 
	\key_tlv_ob_tlv.tdata [54], \key_tlv_ob_tlv.tdata [53], 
	\key_tlv_ob_tlv.tdata [52], \key_tlv_ob_tlv.tdata [51], 
	\key_tlv_ob_tlv.tdata [50], \key_tlv_ob_tlv.tdata [49], 
	\key_tlv_ob_tlv.tdata [48], \key_tlv_ob_tlv.tdata [47], 
	\key_tlv_ob_tlv.tdata [46], \key_tlv_ob_tlv.tdata [45], 
	\key_tlv_ob_tlv.tdata [44], \key_tlv_ob_tlv.tdata [43], 
	\key_tlv_ob_tlv.tdata [42], \key_tlv_ob_tlv.tdata [41], 
	\key_tlv_ob_tlv.tdata [40], \key_tlv_ob_tlv.tdata [39], 
	\key_tlv_ob_tlv.tdata [38], \key_tlv_ob_tlv.tdata [37], 
	\key_tlv_ob_tlv.tdata [36], \key_tlv_ob_tlv.tdata [35], 
	\key_tlv_ob_tlv.tdata [34], \key_tlv_ob_tlv.tdata [33], 
	\key_tlv_ob_tlv.tdata [32], \key_tlv_ob_tlv.tdata [31], 
	\key_tlv_ob_tlv.tdata [30], \key_tlv_ob_tlv.tdata [29], 
	\key_tlv_ob_tlv.tdata [28], \key_tlv_ob_tlv.tdata [27], 
	\key_tlv_ob_tlv.tdata [26], \key_tlv_ob_tlv.tdata [25], 
	\key_tlv_ob_tlv.tdata [24], \key_tlv_ob_tlv.tdata [23], 
	\key_tlv_ob_tlv.tdata [22], \key_tlv_ob_tlv.tdata [21], 
	\key_tlv_ob_tlv.tdata [20], \key_tlv_ob_tlv.tdata [19], 
	\key_tlv_ob_tlv.tdata [18], \key_tlv_ob_tlv.tdata [17], 
	\key_tlv_ob_tlv.tdata [16], \key_tlv_ob_tlv.tdata [15], 
	\key_tlv_ob_tlv.tdata [14], \key_tlv_ob_tlv.tdata [13], 
	\key_tlv_ob_tlv.tdata [12], \key_tlv_ob_tlv.tdata [11], 
	\key_tlv_ob_tlv.tdata [10], \key_tlv_ob_tlv.tdata [9], 
	\key_tlv_ob_tlv.tdata [8], \key_tlv_ob_tlv.tdata [7], 
	\key_tlv_ob_tlv.tdata [6], \key_tlv_ob_tlv.tdata [5], 
	\key_tlv_ob_tlv.tdata [4], \key_tlv_ob_tlv.tdata [3], 
	\key_tlv_ob_tlv.tdata [2], \key_tlv_ob_tlv.tdata [1], 
	\key_tlv_ob_tlv.tdata [0]} ), set_gcm_tag_fail_int, clk, rst_n, 
	scan_en, scan_mode, scan_rst_n, .labels( {\labels[7].guid_size[0] , 
	\labels[7].label_size[5] , \labels[7].label_size[4] , 
	\labels[7].label_size[3] , \labels[7].label_size[2] , 
	\labels[7].label_size[1] , \labels[7].label_size[0] , 
	\labels[7].label[255] , \labels[7].label[254] , 
	\labels[7].label[253] , \labels[7].label[252] , 
	\labels[7].label[251] , \labels[7].label[250] , 
	\labels[7].label[249] , \labels[7].label[248] , 
	\labels[7].label[247] , \labels[7].label[246] , 
	\labels[7].label[245] , \labels[7].label[244] , 
	\labels[7].label[243] , \labels[7].label[242] , 
	\labels[7].label[241] , \labels[7].label[240] , 
	\labels[7].label[239] , \labels[7].label[238] , 
	\labels[7].label[237] , \labels[7].label[236] , 
	\labels[7].label[235] , \labels[7].label[234] , 
	\labels[7].label[233] , \labels[7].label[232] , 
	\labels[7].label[231] , \labels[7].label[230] , 
	\labels[7].label[229] , \labels[7].label[228] , 
	\labels[7].label[227] , \labels[7].label[226] , 
	\labels[7].label[225] , \labels[7].label[224] , 
	\labels[7].label[223] , \labels[7].label[222] , 
	\labels[7].label[221] , \labels[7].label[220] , 
	\labels[7].label[219] , \labels[7].label[218] , 
	\labels[7].label[217] , \labels[7].label[216] , 
	\labels[7].label[215] , \labels[7].label[214] , 
	\labels[7].label[213] , \labels[7].label[212] , 
	\labels[7].label[211] , \labels[7].label[210] , 
	\labels[7].label[209] , \labels[7].label[208] , 
	\labels[7].label[207] , \labels[7].label[206] , 
	\labels[7].label[205] , \labels[7].label[204] , 
	\labels[7].label[203] , \labels[7].label[202] , 
	\labels[7].label[201] , \labels[7].label[200] , 
	\labels[7].label[199] , \labels[7].label[198] , 
	\labels[7].label[197] , \labels[7].label[196] , 
	\labels[7].label[195] , \labels[7].label[194] , 
	\labels[7].label[193] , \labels[7].label[192] , 
	\labels[7].label[191] , \labels[7].label[190] , 
	\labels[7].label[189] , \labels[7].label[188] , 
	\labels[7].label[187] , \labels[7].label[186] , 
	\labels[7].label[185] , \labels[7].label[184] , 
	\labels[7].label[183] , \labels[7].label[182] , 
	\labels[7].label[181] , \labels[7].label[180] , 
	\labels[7].label[179] , \labels[7].label[178] , 
	\labels[7].label[177] , \labels[7].label[176] , 
	\labels[7].label[175] , \labels[7].label[174] , 
	\labels[7].label[173] , \labels[7].label[172] , 
	\labels[7].label[171] , \labels[7].label[170] , 
	\labels[7].label[169] , \labels[7].label[168] , 
	\labels[7].label[167] , \labels[7].label[166] , 
	\labels[7].label[165] , \labels[7].label[164] , 
	\labels[7].label[163] , \labels[7].label[162] , 
	\labels[7].label[161] , \labels[7].label[160] , 
	\labels[7].label[159] , \labels[7].label[158] , 
	\labels[7].label[157] , \labels[7].label[156] , 
	\labels[7].label[155] , \labels[7].label[154] , 
	\labels[7].label[153] , \labels[7].label[152] , 
	\labels[7].label[151] , \labels[7].label[150] , 
	\labels[7].label[149] , \labels[7].label[148] , 
	\labels[7].label[147] , \labels[7].label[146] , 
	\labels[7].label[145] , \labels[7].label[144] , 
	\labels[7].label[143] , \labels[7].label[142] , 
	\labels[7].label[141] , \labels[7].label[140] , 
	\labels[7].label[139] , \labels[7].label[138] , 
	\labels[7].label[137] , \labels[7].label[136] , 
	\labels[7].label[135] , \labels[7].label[134] , 
	\labels[7].label[133] , \labels[7].label[132] , 
	\labels[7].label[131] , \labels[7].label[130] , 
	\labels[7].label[129] , \labels[7].label[128] , 
	\labels[7].label[127] , \labels[7].label[126] , 
	\labels[7].label[125] , \labels[7].label[124] , 
	\labels[7].label[123] , \labels[7].label[122] , 
	\labels[7].label[121] , \labels[7].label[120] , 
	\labels[7].label[119] , \labels[7].label[118] , 
	\labels[7].label[117] , \labels[7].label[116] , 
	\labels[7].label[115] , \labels[7].label[114] , 
	\labels[7].label[113] , \labels[7].label[112] , 
	\labels[7].label[111] , \labels[7].label[110] , 
	\labels[7].label[109] , \labels[7].label[108] , 
	\labels[7].label[107] , \labels[7].label[106] , 
	\labels[7].label[105] , \labels[7].label[104] , 
	\labels[7].label[103] , \labels[7].label[102] , 
	\labels[7].label[101] , \labels[7].label[100] , 
	\labels[7].label[99] , \labels[7].label[98] , \labels[7].label[97] , 
	\labels[7].label[96] , \labels[7].label[95] , \labels[7].label[94] , 
	\labels[7].label[93] , \labels[7].label[92] , \labels[7].label[91] , 
	\labels[7].label[90] , \labels[7].label[89] , \labels[7].label[88] , 
	\labels[7].label[87] , \labels[7].label[86] , \labels[7].label[85] , 
	\labels[7].label[84] , \labels[7].label[83] , \labels[7].label[82] , 
	\labels[7].label[81] , \labels[7].label[80] , \labels[7].label[79] , 
	\labels[7].label[78] , \labels[7].label[77] , \labels[7].label[76] , 
	\labels[7].label[75] , \labels[7].label[74] , \labels[7].label[73] , 
	\labels[7].label[72] , \labels[7].label[71] , \labels[7].label[70] , 
	\labels[7].label[69] , \labels[7].label[68] , \labels[7].label[67] , 
	\labels[7].label[66] , \labels[7].label[65] , \labels[7].label[64] , 
	\labels[7].label[63] , \labels[7].label[62] , \labels[7].label[61] , 
	\labels[7].label[60] , \labels[7].label[59] , \labels[7].label[58] , 
	\labels[7].label[57] , \labels[7].label[56] , \labels[7].label[55] , 
	\labels[7].label[54] , \labels[7].label[53] , \labels[7].label[52] , 
	\labels[7].label[51] , \labels[7].label[50] , \labels[7].label[49] , 
	\labels[7].label[48] , \labels[7].label[47] , \labels[7].label[46] , 
	\labels[7].label[45] , \labels[7].label[44] , \labels[7].label[43] , 
	\labels[7].label[42] , \labels[7].label[41] , \labels[7].label[40] , 
	\labels[7].label[39] , \labels[7].label[38] , \labels[7].label[37] , 
	\labels[7].label[36] , \labels[7].label[35] , \labels[7].label[34] , 
	\labels[7].label[33] , \labels[7].label[32] , \labels[7].label[31] , 
	\labels[7].label[30] , \labels[7].label[29] , \labels[7].label[28] , 
	\labels[7].label[27] , \labels[7].label[26] , \labels[7].label[25] , 
	\labels[7].label[24] , \labels[7].label[23] , \labels[7].label[22] , 
	\labels[7].label[21] , \labels[7].label[20] , \labels[7].label[19] , 
	\labels[7].label[18] , \labels[7].label[17] , \labels[7].label[16] , 
	\labels[7].label[15] , \labels[7].label[14] , \labels[7].label[13] , 
	\labels[7].label[12] , \labels[7].label[11] , \labels[7].label[10] , 
	\labels[7].label[9] , \labels[7].label[8] , \labels[7].label[7] , 
	\labels[7].label[6] , \labels[7].label[5] , \labels[7].label[4] , 
	\labels[7].label[3] , \labels[7].label[2] , \labels[7].label[1] , 
	\labels[7].label[0] , \labels[7].delimiter_valid[0] , 
	\labels[7].delimiter[7] , \labels[7].delimiter[6] , 
	\labels[7].delimiter[5] , \labels[7].delimiter[4] , 
	\labels[7].delimiter[3] , \labels[7].delimiter[2] , 
	\labels[7].delimiter[1] , \labels[7].delimiter[0] , 
	\labels[6].guid_size[0] , \labels[6].label_size[5] , 
	\labels[6].label_size[4] , \labels[6].label_size[3] , 
	\labels[6].label_size[2] , \labels[6].label_size[1] , 
	\labels[6].label_size[0] , \labels[6].label[255] , 
	\labels[6].label[254] , \labels[6].label[253] , 
	\labels[6].label[252] , \labels[6].label[251] , 
	\labels[6].label[250] , \labels[6].label[249] , 
	\labels[6].label[248] , \labels[6].label[247] , 
	\labels[6].label[246] , \labels[6].label[245] , 
	\labels[6].label[244] , \labels[6].label[243] , 
	\labels[6].label[242] , \labels[6].label[241] , 
	\labels[6].label[240] , \labels[6].label[239] , 
	\labels[6].label[238] , \labels[6].label[237] , 
	\labels[6].label[236] , \labels[6].label[235] , 
	\labels[6].label[234] , \labels[6].label[233] , 
	\labels[6].label[232] , \labels[6].label[231] , 
	\labels[6].label[230] , \labels[6].label[229] , 
	\labels[6].label[228] , \labels[6].label[227] , 
	\labels[6].label[226] , \labels[6].label[225] , 
	\labels[6].label[224] , \labels[6].label[223] , 
	\labels[6].label[222] , \labels[6].label[221] , 
	\labels[6].label[220] , \labels[6].label[219] , 
	\labels[6].label[218] , \labels[6].label[217] , 
	\labels[6].label[216] , \labels[6].label[215] , 
	\labels[6].label[214] , \labels[6].label[213] , 
	\labels[6].label[212] , \labels[6].label[211] , 
	\labels[6].label[210] , \labels[6].label[209] , 
	\labels[6].label[208] , \labels[6].label[207] , 
	\labels[6].label[206] , \labels[6].label[205] , 
	\labels[6].label[204] , \labels[6].label[203] , 
	\labels[6].label[202] , \labels[6].label[201] , 
	\labels[6].label[200] , \labels[6].label[199] , 
	\labels[6].label[198] , \labels[6].label[197] , 
	\labels[6].label[196] , \labels[6].label[195] , 
	\labels[6].label[194] , \labels[6].label[193] , 
	\labels[6].label[192] , \labels[6].label[191] , 
	\labels[6].label[190] , \labels[6].label[189] , 
	\labels[6].label[188] , \labels[6].label[187] , 
	\labels[6].label[186] , \labels[6].label[185] , 
	\labels[6].label[184] , \labels[6].label[183] , 
	\labels[6].label[182] , \labels[6].label[181] , 
	\labels[6].label[180] , \labels[6].label[179] , 
	\labels[6].label[178] , \labels[6].label[177] , 
	\labels[6].label[176] , \labels[6].label[175] , 
	\labels[6].label[174] , \labels[6].label[173] , 
	\labels[6].label[172] , \labels[6].label[171] , 
	\labels[6].label[170] , \labels[6].label[169] , 
	\labels[6].label[168] , \labels[6].label[167] , 
	\labels[6].label[166] , \labels[6].label[165] , 
	\labels[6].label[164] , \labels[6].label[163] , 
	\labels[6].label[162] , \labels[6].label[161] , 
	\labels[6].label[160] , \labels[6].label[159] , 
	\labels[6].label[158] , \labels[6].label[157] , 
	\labels[6].label[156] , \labels[6].label[155] , 
	\labels[6].label[154] , \labels[6].label[153] , 
	\labels[6].label[152] , \labels[6].label[151] , 
	\labels[6].label[150] , \labels[6].label[149] , 
	\labels[6].label[148] , \labels[6].label[147] , 
	\labels[6].label[146] , \labels[6].label[145] , 
	\labels[6].label[144] , \labels[6].label[143] , 
	\labels[6].label[142] , \labels[6].label[141] , 
	\labels[6].label[140] , \labels[6].label[139] , 
	\labels[6].label[138] , \labels[6].label[137] , 
	\labels[6].label[136] , \labels[6].label[135] , 
	\labels[6].label[134] , \labels[6].label[133] , 
	\labels[6].label[132] , \labels[6].label[131] , 
	\labels[6].label[130] , \labels[6].label[129] , 
	\labels[6].label[128] , \labels[6].label[127] , 
	\labels[6].label[126] , \labels[6].label[125] , 
	\labels[6].label[124] , \labels[6].label[123] , 
	\labels[6].label[122] , \labels[6].label[121] , 
	\labels[6].label[120] , \labels[6].label[119] , 
	\labels[6].label[118] , \labels[6].label[117] , 
	\labels[6].label[116] , \labels[6].label[115] , 
	\labels[6].label[114] , \labels[6].label[113] , 
	\labels[6].label[112] , \labels[6].label[111] , 
	\labels[6].label[110] , \labels[6].label[109] , 
	\labels[6].label[108] , \labels[6].label[107] , 
	\labels[6].label[106] , \labels[6].label[105] , 
	\labels[6].label[104] , \labels[6].label[103] , 
	\labels[6].label[102] , \labels[6].label[101] , 
	\labels[6].label[100] , \labels[6].label[99] , \labels[6].label[98] , 
	\labels[6].label[97] , \labels[6].label[96] , \labels[6].label[95] , 
	\labels[6].label[94] , \labels[6].label[93] , \labels[6].label[92] , 
	\labels[6].label[91] , \labels[6].label[90] , \labels[6].label[89] , 
	\labels[6].label[88] , \labels[6].label[87] , \labels[6].label[86] , 
	\labels[6].label[85] , \labels[6].label[84] , \labels[6].label[83] , 
	\labels[6].label[82] , \labels[6].label[81] , \labels[6].label[80] , 
	\labels[6].label[79] , \labels[6].label[78] , \labels[6].label[77] , 
	\labels[6].label[76] , \labels[6].label[75] , \labels[6].label[74] , 
	\labels[6].label[73] , \labels[6].label[72] , \labels[6].label[71] , 
	\labels[6].label[70] , \labels[6].label[69] , \labels[6].label[68] , 
	\labels[6].label[67] , \labels[6].label[66] , \labels[6].label[65] , 
	\labels[6].label[64] , \labels[6].label[63] , \labels[6].label[62] , 
	\labels[6].label[61] , \labels[6].label[60] , \labels[6].label[59] , 
	\labels[6].label[58] , \labels[6].label[57] , \labels[6].label[56] , 
	\labels[6].label[55] , \labels[6].label[54] , \labels[6].label[53] , 
	\labels[6].label[52] , \labels[6].label[51] , \labels[6].label[50] , 
	\labels[6].label[49] , \labels[6].label[48] , \labels[6].label[47] , 
	\labels[6].label[46] , \labels[6].label[45] , \labels[6].label[44] , 
	\labels[6].label[43] , \labels[6].label[42] , \labels[6].label[41] , 
	\labels[6].label[40] , \labels[6].label[39] , \labels[6].label[38] , 
	\labels[6].label[37] , \labels[6].label[36] , \labels[6].label[35] , 
	\labels[6].label[34] , \labels[6].label[33] , \labels[6].label[32] , 
	\labels[6].label[31] , \labels[6].label[30] , \labels[6].label[29] , 
	\labels[6].label[28] , \labels[6].label[27] , \labels[6].label[26] , 
	\labels[6].label[25] , \labels[6].label[24] , \labels[6].label[23] , 
	\labels[6].label[22] , \labels[6].label[21] , \labels[6].label[20] , 
	\labels[6].label[19] , \labels[6].label[18] , \labels[6].label[17] , 
	\labels[6].label[16] , \labels[6].label[15] , \labels[6].label[14] , 
	\labels[6].label[13] , \labels[6].label[12] , \labels[6].label[11] , 
	\labels[6].label[10] , \labels[6].label[9] , \labels[6].label[8] , 
	\labels[6].label[7] , \labels[6].label[6] , \labels[6].label[5] , 
	\labels[6].label[4] , \labels[6].label[3] , \labels[6].label[2] , 
	\labels[6].label[1] , \labels[6].label[0] , 
	\labels[6].delimiter_valid[0] , \labels[6].delimiter[7] , 
	\labels[6].delimiter[6] , \labels[6].delimiter[5] , 
	\labels[6].delimiter[4] , \labels[6].delimiter[3] , 
	\labels[6].delimiter[2] , \labels[6].delimiter[1] , 
	\labels[6].delimiter[0] , \labels[5].guid_size[0] , 
	\labels[5].label_size[5] , \labels[5].label_size[4] , 
	\labels[5].label_size[3] , \labels[5].label_size[2] , 
	\labels[5].label_size[1] , \labels[5].label_size[0] , 
	\labels[5].label[255] , \labels[5].label[254] , 
	\labels[5].label[253] , \labels[5].label[252] , 
	\labels[5].label[251] , \labels[5].label[250] , 
	\labels[5].label[249] , \labels[5].label[248] , 
	\labels[5].label[247] , \labels[5].label[246] , 
	\labels[5].label[245] , \labels[5].label[244] , 
	\labels[5].label[243] , \labels[5].label[242] , 
	\labels[5].label[241] , \labels[5].label[240] , 
	\labels[5].label[239] , \labels[5].label[238] , 
	\labels[5].label[237] , \labels[5].label[236] , 
	\labels[5].label[235] , \labels[5].label[234] , 
	\labels[5].label[233] , \labels[5].label[232] , 
	\labels[5].label[231] , \labels[5].label[230] , 
	\labels[5].label[229] , \labels[5].label[228] , 
	\labels[5].label[227] , \labels[5].label[226] , 
	\labels[5].label[225] , \labels[5].label[224] , 
	\labels[5].label[223] , \labels[5].label[222] , 
	\labels[5].label[221] , \labels[5].label[220] , 
	\labels[5].label[219] , \labels[5].label[218] , 
	\labels[5].label[217] , \labels[5].label[216] , 
	\labels[5].label[215] , \labels[5].label[214] , 
	\labels[5].label[213] , \labels[5].label[212] , 
	\labels[5].label[211] , \labels[5].label[210] , 
	\labels[5].label[209] , \labels[5].label[208] , 
	\labels[5].label[207] , \labels[5].label[206] , 
	\labels[5].label[205] , \labels[5].label[204] , 
	\labels[5].label[203] , \labels[5].label[202] , 
	\labels[5].label[201] , \labels[5].label[200] , 
	\labels[5].label[199] , \labels[5].label[198] , 
	\labels[5].label[197] , \labels[5].label[196] , 
	\labels[5].label[195] , \labels[5].label[194] , 
	\labels[5].label[193] , \labels[5].label[192] , 
	\labels[5].label[191] , \labels[5].label[190] , 
	\labels[5].label[189] , \labels[5].label[188] , 
	\labels[5].label[187] , \labels[5].label[186] , 
	\labels[5].label[185] , \labels[5].label[184] , 
	\labels[5].label[183] , \labels[5].label[182] , 
	\labels[5].label[181] , \labels[5].label[180] , 
	\labels[5].label[179] , \labels[5].label[178] , 
	\labels[5].label[177] , \labels[5].label[176] , 
	\labels[5].label[175] , \labels[5].label[174] , 
	\labels[5].label[173] , \labels[5].label[172] , 
	\labels[5].label[171] , \labels[5].label[170] , 
	\labels[5].label[169] , \labels[5].label[168] , 
	\labels[5].label[167] , \labels[5].label[166] , 
	\labels[5].label[165] , \labels[5].label[164] , 
	\labels[5].label[163] , \labels[5].label[162] , 
	\labels[5].label[161] , \labels[5].label[160] , 
	\labels[5].label[159] , \labels[5].label[158] , 
	\labels[5].label[157] , \labels[5].label[156] , 
	\labels[5].label[155] , \labels[5].label[154] , 
	\labels[5].label[153] , \labels[5].label[152] , 
	\labels[5].label[151] , \labels[5].label[150] , 
	\labels[5].label[149] , \labels[5].label[148] , 
	\labels[5].label[147] , \labels[5].label[146] , 
	\labels[5].label[145] , \labels[5].label[144] , 
	\labels[5].label[143] , \labels[5].label[142] , 
	\labels[5].label[141] , \labels[5].label[140] , 
	\labels[5].label[139] , \labels[5].label[138] , 
	\labels[5].label[137] , \labels[5].label[136] , 
	\labels[5].label[135] , \labels[5].label[134] , 
	\labels[5].label[133] , \labels[5].label[132] , 
	\labels[5].label[131] , \labels[5].label[130] , 
	\labels[5].label[129] , \labels[5].label[128] , 
	\labels[5].label[127] , \labels[5].label[126] , 
	\labels[5].label[125] , \labels[5].label[124] , 
	\labels[5].label[123] , \labels[5].label[122] , 
	\labels[5].label[121] , \labels[5].label[120] , 
	\labels[5].label[119] , \labels[5].label[118] , 
	\labels[5].label[117] , \labels[5].label[116] , 
	\labels[5].label[115] , \labels[5].label[114] , 
	\labels[5].label[113] , \labels[5].label[112] , 
	\labels[5].label[111] , \labels[5].label[110] , 
	\labels[5].label[109] , \labels[5].label[108] , 
	\labels[5].label[107] , \labels[5].label[106] , 
	\labels[5].label[105] , \labels[5].label[104] , 
	\labels[5].label[103] , \labels[5].label[102] , 
	\labels[5].label[101] , \labels[5].label[100] , 
	\labels[5].label[99] , \labels[5].label[98] , \labels[5].label[97] , 
	\labels[5].label[96] , \labels[5].label[95] , \labels[5].label[94] , 
	\labels[5].label[93] , \labels[5].label[92] , \labels[5].label[91] , 
	\labels[5].label[90] , \labels[5].label[89] , \labels[5].label[88] , 
	\labels[5].label[87] , \labels[5].label[86] , \labels[5].label[85] , 
	\labels[5].label[84] , \labels[5].label[83] , \labels[5].label[82] , 
	\labels[5].label[81] , \labels[5].label[80] , \labels[5].label[79] , 
	\labels[5].label[78] , \labels[5].label[77] , \labels[5].label[76] , 
	\labels[5].label[75] , \labels[5].label[74] , \labels[5].label[73] , 
	\labels[5].label[72] , \labels[5].label[71] , \labels[5].label[70] , 
	\labels[5].label[69] , \labels[5].label[68] , \labels[5].label[67] , 
	\labels[5].label[66] , \labels[5].label[65] , \labels[5].label[64] , 
	\labels[5].label[63] , \labels[5].label[62] , \labels[5].label[61] , 
	\labels[5].label[60] , \labels[5].label[59] , \labels[5].label[58] , 
	\labels[5].label[57] , \labels[5].label[56] , \labels[5].label[55] , 
	\labels[5].label[54] , \labels[5].label[53] , \labels[5].label[52] , 
	\labels[5].label[51] , \labels[5].label[50] , \labels[5].label[49] , 
	\labels[5].label[48] , \labels[5].label[47] , \labels[5].label[46] , 
	\labels[5].label[45] , \labels[5].label[44] , \labels[5].label[43] , 
	\labels[5].label[42] , \labels[5].label[41] , \labels[5].label[40] , 
	\labels[5].label[39] , \labels[5].label[38] , \labels[5].label[37] , 
	\labels[5].label[36] , \labels[5].label[35] , \labels[5].label[34] , 
	\labels[5].label[33] , \labels[5].label[32] , \labels[5].label[31] , 
	\labels[5].label[30] , \labels[5].label[29] , \labels[5].label[28] , 
	\labels[5].label[27] , \labels[5].label[26] , \labels[5].label[25] , 
	\labels[5].label[24] , \labels[5].label[23] , \labels[5].label[22] , 
	\labels[5].label[21] , \labels[5].label[20] , \labels[5].label[19] , 
	\labels[5].label[18] , \labels[5].label[17] , \labels[5].label[16] , 
	\labels[5].label[15] , \labels[5].label[14] , \labels[5].label[13] , 
	\labels[5].label[12] , \labels[5].label[11] , \labels[5].label[10] , 
	\labels[5].label[9] , \labels[5].label[8] , \labels[5].label[7] , 
	\labels[5].label[6] , \labels[5].label[5] , \labels[5].label[4] , 
	\labels[5].label[3] , \labels[5].label[2] , \labels[5].label[1] , 
	\labels[5].label[0] , \labels[5].delimiter_valid[0] , 
	\labels[5].delimiter[7] , \labels[5].delimiter[6] , 
	\labels[5].delimiter[5] , \labels[5].delimiter[4] , 
	\labels[5].delimiter[3] , \labels[5].delimiter[2] , 
	\labels[5].delimiter[1] , \labels[5].delimiter[0] , 
	\labels[4].guid_size[0] , \labels[4].label_size[5] , 
	\labels[4].label_size[4] , \labels[4].label_size[3] , 
	\labels[4].label_size[2] , \labels[4].label_size[1] , 
	\labels[4].label_size[0] , \labels[4].label[255] , 
	\labels[4].label[254] , \labels[4].label[253] , 
	\labels[4].label[252] , \labels[4].label[251] , 
	\labels[4].label[250] , \labels[4].label[249] , 
	\labels[4].label[248] , \labels[4].label[247] , 
	\labels[4].label[246] , \labels[4].label[245] , 
	\labels[4].label[244] , \labels[4].label[243] , 
	\labels[4].label[242] , \labels[4].label[241] , 
	\labels[4].label[240] , \labels[4].label[239] , 
	\labels[4].label[238] , \labels[4].label[237] , 
	\labels[4].label[236] , \labels[4].label[235] , 
	\labels[4].label[234] , \labels[4].label[233] , 
	\labels[4].label[232] , \labels[4].label[231] , 
	\labels[4].label[230] , \labels[4].label[229] , 
	\labels[4].label[228] , \labels[4].label[227] , 
	\labels[4].label[226] , \labels[4].label[225] , 
	\labels[4].label[224] , \labels[4].label[223] , 
	\labels[4].label[222] , \labels[4].label[221] , 
	\labels[4].label[220] , \labels[4].label[219] , 
	\labels[4].label[218] , \labels[4].label[217] , 
	\labels[4].label[216] , \labels[4].label[215] , 
	\labels[4].label[214] , \labels[4].label[213] , 
	\labels[4].label[212] , \labels[4].label[211] , 
	\labels[4].label[210] , \labels[4].label[209] , 
	\labels[4].label[208] , \labels[4].label[207] , 
	\labels[4].label[206] , \labels[4].label[205] , 
	\labels[4].label[204] , \labels[4].label[203] , 
	\labels[4].label[202] , \labels[4].label[201] , 
	\labels[4].label[200] , \labels[4].label[199] , 
	\labels[4].label[198] , \labels[4].label[197] , 
	\labels[4].label[196] , \labels[4].label[195] , 
	\labels[4].label[194] , \labels[4].label[193] , 
	\labels[4].label[192] , \labels[4].label[191] , 
	\labels[4].label[190] , \labels[4].label[189] , 
	\labels[4].label[188] , \labels[4].label[187] , 
	\labels[4].label[186] , \labels[4].label[185] , 
	\labels[4].label[184] , \labels[4].label[183] , 
	\labels[4].label[182] , \labels[4].label[181] , 
	\labels[4].label[180] , \labels[4].label[179] , 
	\labels[4].label[178] , \labels[4].label[177] , 
	\labels[4].label[176] , \labels[4].label[175] , 
	\labels[4].label[174] , \labels[4].label[173] , 
	\labels[4].label[172] , \labels[4].label[171] , 
	\labels[4].label[170] , \labels[4].label[169] , 
	\labels[4].label[168] , \labels[4].label[167] , 
	\labels[4].label[166] , \labels[4].label[165] , 
	\labels[4].label[164] , \labels[4].label[163] , 
	\labels[4].label[162] , \labels[4].label[161] , 
	\labels[4].label[160] , \labels[4].label[159] , 
	\labels[4].label[158] , \labels[4].label[157] , 
	\labels[4].label[156] , \labels[4].label[155] , 
	\labels[4].label[154] , \labels[4].label[153] , 
	\labels[4].label[152] , \labels[4].label[151] , 
	\labels[4].label[150] , \labels[4].label[149] , 
	\labels[4].label[148] , \labels[4].label[147] , 
	\labels[4].label[146] , \labels[4].label[145] , 
	\labels[4].label[144] , \labels[4].label[143] , 
	\labels[4].label[142] , \labels[4].label[141] , 
	\labels[4].label[140] , \labels[4].label[139] , 
	\labels[4].label[138] , \labels[4].label[137] , 
	\labels[4].label[136] , \labels[4].label[135] , 
	\labels[4].label[134] , \labels[4].label[133] , 
	\labels[4].label[132] , \labels[4].label[131] , 
	\labels[4].label[130] , \labels[4].label[129] , 
	\labels[4].label[128] , \labels[4].label[127] , 
	\labels[4].label[126] , \labels[4].label[125] , 
	\labels[4].label[124] , \labels[4].label[123] , 
	\labels[4].label[122] , \labels[4].label[121] , 
	\labels[4].label[120] , \labels[4].label[119] , 
	\labels[4].label[118] , \labels[4].label[117] , 
	\labels[4].label[116] , \labels[4].label[115] , 
	\labels[4].label[114] , \labels[4].label[113] , 
	\labels[4].label[112] , \labels[4].label[111] , 
	\labels[4].label[110] , \labels[4].label[109] , 
	\labels[4].label[108] , \labels[4].label[107] , 
	\labels[4].label[106] , \labels[4].label[105] , 
	\labels[4].label[104] , \labels[4].label[103] , 
	\labels[4].label[102] , \labels[4].label[101] , 
	\labels[4].label[100] , \labels[4].label[99] , \labels[4].label[98] , 
	\labels[4].label[97] , \labels[4].label[96] , \labels[4].label[95] , 
	\labels[4].label[94] , \labels[4].label[93] , \labels[4].label[92] , 
	\labels[4].label[91] , \labels[4].label[90] , \labels[4].label[89] , 
	\labels[4].label[88] , \labels[4].label[87] , \labels[4].label[86] , 
	\labels[4].label[85] , \labels[4].label[84] , \labels[4].label[83] , 
	\labels[4].label[82] , \labels[4].label[81] , \labels[4].label[80] , 
	\labels[4].label[79] , \labels[4].label[78] , \labels[4].label[77] , 
	\labels[4].label[76] , \labels[4].label[75] , \labels[4].label[74] , 
	\labels[4].label[73] , \labels[4].label[72] , \labels[4].label[71] , 
	\labels[4].label[70] , \labels[4].label[69] , \labels[4].label[68] , 
	\labels[4].label[67] , \labels[4].label[66] , \labels[4].label[65] , 
	\labels[4].label[64] , \labels[4].label[63] , \labels[4].label[62] , 
	\labels[4].label[61] , \labels[4].label[60] , \labels[4].label[59] , 
	\labels[4].label[58] , \labels[4].label[57] , \labels[4].label[56] , 
	\labels[4].label[55] , \labels[4].label[54] , \labels[4].label[53] , 
	\labels[4].label[52] , \labels[4].label[51] , \labels[4].label[50] , 
	\labels[4].label[49] , \labels[4].label[48] , \labels[4].label[47] , 
	\labels[4].label[46] , \labels[4].label[45] , \labels[4].label[44] , 
	\labels[4].label[43] , \labels[4].label[42] , \labels[4].label[41] , 
	\labels[4].label[40] , \labels[4].label[39] , \labels[4].label[38] , 
	\labels[4].label[37] , \labels[4].label[36] , \labels[4].label[35] , 
	\labels[4].label[34] , \labels[4].label[33] , \labels[4].label[32] , 
	\labels[4].label[31] , \labels[4].label[30] , \labels[4].label[29] , 
	\labels[4].label[28] , \labels[4].label[27] , \labels[4].label[26] , 
	\labels[4].label[25] , \labels[4].label[24] , \labels[4].label[23] , 
	\labels[4].label[22] , \labels[4].label[21] , \labels[4].label[20] , 
	\labels[4].label[19] , \labels[4].label[18] , \labels[4].label[17] , 
	\labels[4].label[16] , \labels[4].label[15] , \labels[4].label[14] , 
	\labels[4].label[13] , \labels[4].label[12] , \labels[4].label[11] , 
	\labels[4].label[10] , \labels[4].label[9] , \labels[4].label[8] , 
	\labels[4].label[7] , \labels[4].label[6] , \labels[4].label[5] , 
	\labels[4].label[4] , \labels[4].label[3] , \labels[4].label[2] , 
	\labels[4].label[1] , \labels[4].label[0] , 
	\labels[4].delimiter_valid[0] , \labels[4].delimiter[7] , 
	\labels[4].delimiter[6] , \labels[4].delimiter[5] , 
	\labels[4].delimiter[4] , \labels[4].delimiter[3] , 
	\labels[4].delimiter[2] , \labels[4].delimiter[1] , 
	\labels[4].delimiter[0] , \labels[3].guid_size[0] , 
	\labels[3].label_size[5] , \labels[3].label_size[4] , 
	\labels[3].label_size[3] , \labels[3].label_size[2] , 
	\labels[3].label_size[1] , \labels[3].label_size[0] , 
	\labels[3].label[255] , \labels[3].label[254] , 
	\labels[3].label[253] , \labels[3].label[252] , 
	\labels[3].label[251] , \labels[3].label[250] , 
	\labels[3].label[249] , \labels[3].label[248] , 
	\labels[3].label[247] , \labels[3].label[246] , 
	\labels[3].label[245] , \labels[3].label[244] , 
	\labels[3].label[243] , \labels[3].label[242] , 
	\labels[3].label[241] , \labels[3].label[240] , 
	\labels[3].label[239] , \labels[3].label[238] , 
	\labels[3].label[237] , \labels[3].label[236] , 
	\labels[3].label[235] , \labels[3].label[234] , 
	\labels[3].label[233] , \labels[3].label[232] , 
	\labels[3].label[231] , \labels[3].label[230] , 
	\labels[3].label[229] , \labels[3].label[228] , 
	\labels[3].label[227] , \labels[3].label[226] , 
	\labels[3].label[225] , \labels[3].label[224] , 
	\labels[3].label[223] , \labels[3].label[222] , 
	\labels[3].label[221] , \labels[3].label[220] , 
	\labels[3].label[219] , \labels[3].label[218] , 
	\labels[3].label[217] , \labels[3].label[216] , 
	\labels[3].label[215] , \labels[3].label[214] , 
	\labels[3].label[213] , \labels[3].label[212] , 
	\labels[3].label[211] , \labels[3].label[210] , 
	\labels[3].label[209] , \labels[3].label[208] , 
	\labels[3].label[207] , \labels[3].label[206] , 
	\labels[3].label[205] , \labels[3].label[204] , 
	\labels[3].label[203] , \labels[3].label[202] , 
	\labels[3].label[201] , \labels[3].label[200] , 
	\labels[3].label[199] , \labels[3].label[198] , 
	\labels[3].label[197] , \labels[3].label[196] , 
	\labels[3].label[195] , \labels[3].label[194] , 
	\labels[3].label[193] , \labels[3].label[192] , 
	\labels[3].label[191] , \labels[3].label[190] , 
	\labels[3].label[189] , \labels[3].label[188] , 
	\labels[3].label[187] , \labels[3].label[186] , 
	\labels[3].label[185] , \labels[3].label[184] , 
	\labels[3].label[183] , \labels[3].label[182] , 
	\labels[3].label[181] , \labels[3].label[180] , 
	\labels[3].label[179] , \labels[3].label[178] , 
	\labels[3].label[177] , \labels[3].label[176] , 
	\labels[3].label[175] , \labels[3].label[174] , 
	\labels[3].label[173] , \labels[3].label[172] , 
	\labels[3].label[171] , \labels[3].label[170] , 
	\labels[3].label[169] , \labels[3].label[168] , 
	\labels[3].label[167] , \labels[3].label[166] , 
	\labels[3].label[165] , \labels[3].label[164] , 
	\labels[3].label[163] , \labels[3].label[162] , 
	\labels[3].label[161] , \labels[3].label[160] , 
	\labels[3].label[159] , \labels[3].label[158] , 
	\labels[3].label[157] , \labels[3].label[156] , 
	\labels[3].label[155] , \labels[3].label[154] , 
	\labels[3].label[153] , \labels[3].label[152] , 
	\labels[3].label[151] , \labels[3].label[150] , 
	\labels[3].label[149] , \labels[3].label[148] , 
	\labels[3].label[147] , \labels[3].label[146] , 
	\labels[3].label[145] , \labels[3].label[144] , 
	\labels[3].label[143] , \labels[3].label[142] , 
	\labels[3].label[141] , \labels[3].label[140] , 
	\labels[3].label[139] , \labels[3].label[138] , 
	\labels[3].label[137] , \labels[3].label[136] , 
	\labels[3].label[135] , \labels[3].label[134] , 
	\labels[3].label[133] , \labels[3].label[132] , 
	\labels[3].label[131] , \labels[3].label[130] , 
	\labels[3].label[129] , \labels[3].label[128] , 
	\labels[3].label[127] , \labels[3].label[126] , 
	\labels[3].label[125] , \labels[3].label[124] , 
	\labels[3].label[123] , \labels[3].label[122] , 
	\labels[3].label[121] , \labels[3].label[120] , 
	\labels[3].label[119] , \labels[3].label[118] , 
	\labels[3].label[117] , \labels[3].label[116] , 
	\labels[3].label[115] , \labels[3].label[114] , 
	\labels[3].label[113] , \labels[3].label[112] , 
	\labels[3].label[111] , \labels[3].label[110] , 
	\labels[3].label[109] , \labels[3].label[108] , 
	\labels[3].label[107] , \labels[3].label[106] , 
	\labels[3].label[105] , \labels[3].label[104] , 
	\labels[3].label[103] , \labels[3].label[102] , 
	\labels[3].label[101] , \labels[3].label[100] , 
	\labels[3].label[99] , \labels[3].label[98] , \labels[3].label[97] , 
	\labels[3].label[96] , \labels[3].label[95] , \labels[3].label[94] , 
	\labels[3].label[93] , \labels[3].label[92] , \labels[3].label[91] , 
	\labels[3].label[90] , \labels[3].label[89] , \labels[3].label[88] , 
	\labels[3].label[87] , \labels[3].label[86] , \labels[3].label[85] , 
	\labels[3].label[84] , \labels[3].label[83] , \labels[3].label[82] , 
	\labels[3].label[81] , \labels[3].label[80] , \labels[3].label[79] , 
	\labels[3].label[78] , \labels[3].label[77] , \labels[3].label[76] , 
	\labels[3].label[75] , \labels[3].label[74] , \labels[3].label[73] , 
	\labels[3].label[72] , \labels[3].label[71] , \labels[3].label[70] , 
	\labels[3].label[69] , \labels[3].label[68] , \labels[3].label[67] , 
	\labels[3].label[66] , \labels[3].label[65] , \labels[3].label[64] , 
	\labels[3].label[63] , \labels[3].label[62] , \labels[3].label[61] , 
	\labels[3].label[60] , \labels[3].label[59] , \labels[3].label[58] , 
	\labels[3].label[57] , \labels[3].label[56] , \labels[3].label[55] , 
	\labels[3].label[54] , \labels[3].label[53] , \labels[3].label[52] , 
	\labels[3].label[51] , \labels[3].label[50] , \labels[3].label[49] , 
	\labels[3].label[48] , \labels[3].label[47] , \labels[3].label[46] , 
	\labels[3].label[45] , \labels[3].label[44] , \labels[3].label[43] , 
	\labels[3].label[42] , \labels[3].label[41] , \labels[3].label[40] , 
	\labels[3].label[39] , \labels[3].label[38] , \labels[3].label[37] , 
	\labels[3].label[36] , \labels[3].label[35] , \labels[3].label[34] , 
	\labels[3].label[33] , \labels[3].label[32] , \labels[3].label[31] , 
	\labels[3].label[30] , \labels[3].label[29] , \labels[3].label[28] , 
	\labels[3].label[27] , \labels[3].label[26] , \labels[3].label[25] , 
	\labels[3].label[24] , \labels[3].label[23] , \labels[3].label[22] , 
	\labels[3].label[21] , \labels[3].label[20] , \labels[3].label[19] , 
	\labels[3].label[18] , \labels[3].label[17] , \labels[3].label[16] , 
	\labels[3].label[15] , \labels[3].label[14] , \labels[3].label[13] , 
	\labels[3].label[12] , \labels[3].label[11] , \labels[3].label[10] , 
	\labels[3].label[9] , \labels[3].label[8] , \labels[3].label[7] , 
	\labels[3].label[6] , \labels[3].label[5] , \labels[3].label[4] , 
	\labels[3].label[3] , \labels[3].label[2] , \labels[3].label[1] , 
	\labels[3].label[0] , \labels[3].delimiter_valid[0] , 
	\labels[3].delimiter[7] , \labels[3].delimiter[6] , 
	\labels[3].delimiter[5] , \labels[3].delimiter[4] , 
	\labels[3].delimiter[3] , \labels[3].delimiter[2] , 
	\labels[3].delimiter[1] , \labels[3].delimiter[0] , 
	\labels[2].guid_size[0] , \labels[2].label_size[5] , 
	\labels[2].label_size[4] , \labels[2].label_size[3] , 
	\labels[2].label_size[2] , \labels[2].label_size[1] , 
	\labels[2].label_size[0] , \labels[2].label[255] , 
	\labels[2].label[254] , \labels[2].label[253] , 
	\labels[2].label[252] , \labels[2].label[251] , 
	\labels[2].label[250] , \labels[2].label[249] , 
	\labels[2].label[248] , \labels[2].label[247] , 
	\labels[2].label[246] , \labels[2].label[245] , 
	\labels[2].label[244] , \labels[2].label[243] , 
	\labels[2].label[242] , \labels[2].label[241] , 
	\labels[2].label[240] , \labels[2].label[239] , 
	\labels[2].label[238] , \labels[2].label[237] , 
	\labels[2].label[236] , \labels[2].label[235] , 
	\labels[2].label[234] , \labels[2].label[233] , 
	\labels[2].label[232] , \labels[2].label[231] , 
	\labels[2].label[230] , \labels[2].label[229] , 
	\labels[2].label[228] , \labels[2].label[227] , 
	\labels[2].label[226] , \labels[2].label[225] , 
	\labels[2].label[224] , \labels[2].label[223] , 
	\labels[2].label[222] , \labels[2].label[221] , 
	\labels[2].label[220] , \labels[2].label[219] , 
	\labels[2].label[218] , \labels[2].label[217] , 
	\labels[2].label[216] , \labels[2].label[215] , 
	\labels[2].label[214] , \labels[2].label[213] , 
	\labels[2].label[212] , \labels[2].label[211] , 
	\labels[2].label[210] , \labels[2].label[209] , 
	\labels[2].label[208] , \labels[2].label[207] , 
	\labels[2].label[206] , \labels[2].label[205] , 
	\labels[2].label[204] , \labels[2].label[203] , 
	\labels[2].label[202] , \labels[2].label[201] , 
	\labels[2].label[200] , \labels[2].label[199] , 
	\labels[2].label[198] , \labels[2].label[197] , 
	\labels[2].label[196] , \labels[2].label[195] , 
	\labels[2].label[194] , \labels[2].label[193] , 
	\labels[2].label[192] , \labels[2].label[191] , 
	\labels[2].label[190] , \labels[2].label[189] , 
	\labels[2].label[188] , \labels[2].label[187] , 
	\labels[2].label[186] , \labels[2].label[185] , 
	\labels[2].label[184] , \labels[2].label[183] , 
	\labels[2].label[182] , \labels[2].label[181] , 
	\labels[2].label[180] , \labels[2].label[179] , 
	\labels[2].label[178] , \labels[2].label[177] , 
	\labels[2].label[176] , \labels[2].label[175] , 
	\labels[2].label[174] , \labels[2].label[173] , 
	\labels[2].label[172] , \labels[2].label[171] , 
	\labels[2].label[170] , \labels[2].label[169] , 
	\labels[2].label[168] , \labels[2].label[167] , 
	\labels[2].label[166] , \labels[2].label[165] , 
	\labels[2].label[164] , \labels[2].label[163] , 
	\labels[2].label[162] , \labels[2].label[161] , 
	\labels[2].label[160] , \labels[2].label[159] , 
	\labels[2].label[158] , \labels[2].label[157] , 
	\labels[2].label[156] , \labels[2].label[155] , 
	\labels[2].label[154] , \labels[2].label[153] , 
	\labels[2].label[152] , \labels[2].label[151] , 
	\labels[2].label[150] , \labels[2].label[149] , 
	\labels[2].label[148] , \labels[2].label[147] , 
	\labels[2].label[146] , \labels[2].label[145] , 
	\labels[2].label[144] , \labels[2].label[143] , 
	\labels[2].label[142] , \labels[2].label[141] , 
	\labels[2].label[140] , \labels[2].label[139] , 
	\labels[2].label[138] , \labels[2].label[137] , 
	\labels[2].label[136] , \labels[2].label[135] , 
	\labels[2].label[134] , \labels[2].label[133] , 
	\labels[2].label[132] , \labels[2].label[131] , 
	\labels[2].label[130] , \labels[2].label[129] , 
	\labels[2].label[128] , \labels[2].label[127] , 
	\labels[2].label[126] , \labels[2].label[125] , 
	\labels[2].label[124] , \labels[2].label[123] , 
	\labels[2].label[122] , \labels[2].label[121] , 
	\labels[2].label[120] , \labels[2].label[119] , 
	\labels[2].label[118] , \labels[2].label[117] , 
	\labels[2].label[116] , \labels[2].label[115] , 
	\labels[2].label[114] , \labels[2].label[113] , 
	\labels[2].label[112] , \labels[2].label[111] , 
	\labels[2].label[110] , \labels[2].label[109] , 
	\labels[2].label[108] , \labels[2].label[107] , 
	\labels[2].label[106] , \labels[2].label[105] , 
	\labels[2].label[104] , \labels[2].label[103] , 
	\labels[2].label[102] , \labels[2].label[101] , 
	\labels[2].label[100] , \labels[2].label[99] , \labels[2].label[98] , 
	\labels[2].label[97] , \labels[2].label[96] , \labels[2].label[95] , 
	\labels[2].label[94] , \labels[2].label[93] , \labels[2].label[92] , 
	\labels[2].label[91] , \labels[2].label[90] , \labels[2].label[89] , 
	\labels[2].label[88] , \labels[2].label[87] , \labels[2].label[86] , 
	\labels[2].label[85] , \labels[2].label[84] , \labels[2].label[83] , 
	\labels[2].label[82] , \labels[2].label[81] , \labels[2].label[80] , 
	\labels[2].label[79] , \labels[2].label[78] , \labels[2].label[77] , 
	\labels[2].label[76] , \labels[2].label[75] , \labels[2].label[74] , 
	\labels[2].label[73] , \labels[2].label[72] , \labels[2].label[71] , 
	\labels[2].label[70] , \labels[2].label[69] , \labels[2].label[68] , 
	\labels[2].label[67] , \labels[2].label[66] , \labels[2].label[65] , 
	\labels[2].label[64] , \labels[2].label[63] , \labels[2].label[62] , 
	\labels[2].label[61] , \labels[2].label[60] , \labels[2].label[59] , 
	\labels[2].label[58] , \labels[2].label[57] , \labels[2].label[56] , 
	\labels[2].label[55] , \labels[2].label[54] , \labels[2].label[53] , 
	\labels[2].label[52] , \labels[2].label[51] , \labels[2].label[50] , 
	\labels[2].label[49] , \labels[2].label[48] , \labels[2].label[47] , 
	\labels[2].label[46] , \labels[2].label[45] , \labels[2].label[44] , 
	\labels[2].label[43] , \labels[2].label[42] , \labels[2].label[41] , 
	\labels[2].label[40] , \labels[2].label[39] , \labels[2].label[38] , 
	\labels[2].label[37] , \labels[2].label[36] , \labels[2].label[35] , 
	\labels[2].label[34] , \labels[2].label[33] , \labels[2].label[32] , 
	\labels[2].label[31] , \labels[2].label[30] , \labels[2].label[29] , 
	\labels[2].label[28] , \labels[2].label[27] , \labels[2].label[26] , 
	\labels[2].label[25] , \labels[2].label[24] , \labels[2].label[23] , 
	\labels[2].label[22] , \labels[2].label[21] , \labels[2].label[20] , 
	\labels[2].label[19] , \labels[2].label[18] , \labels[2].label[17] , 
	\labels[2].label[16] , \labels[2].label[15] , \labels[2].label[14] , 
	\labels[2].label[13] , \labels[2].label[12] , \labels[2].label[11] , 
	\labels[2].label[10] , \labels[2].label[9] , \labels[2].label[8] , 
	\labels[2].label[7] , \labels[2].label[6] , \labels[2].label[5] , 
	\labels[2].label[4] , \labels[2].label[3] , \labels[2].label[2] , 
	\labels[2].label[1] , \labels[2].label[0] , 
	\labels[2].delimiter_valid[0] , \labels[2].delimiter[7] , 
	\labels[2].delimiter[6] , \labels[2].delimiter[5] , 
	\labels[2].delimiter[4] , \labels[2].delimiter[3] , 
	\labels[2].delimiter[2] , \labels[2].delimiter[1] , 
	\labels[2].delimiter[0] , \labels[1].guid_size[0] , 
	\labels[1].label_size[5] , \labels[1].label_size[4] , 
	\labels[1].label_size[3] , \labels[1].label_size[2] , 
	\labels[1].label_size[1] , \labels[1].label_size[0] , 
	\labels[1].label[255] , \labels[1].label[254] , 
	\labels[1].label[253] , \labels[1].label[252] , 
	\labels[1].label[251] , \labels[1].label[250] , 
	\labels[1].label[249] , \labels[1].label[248] , 
	\labels[1].label[247] , \labels[1].label[246] , 
	\labels[1].label[245] , \labels[1].label[244] , 
	\labels[1].label[243] , \labels[1].label[242] , 
	\labels[1].label[241] , \labels[1].label[240] , 
	\labels[1].label[239] , \labels[1].label[238] , 
	\labels[1].label[237] , \labels[1].label[236] , 
	\labels[1].label[235] , \labels[1].label[234] , 
	\labels[1].label[233] , \labels[1].label[232] , 
	\labels[1].label[231] , \labels[1].label[230] , 
	\labels[1].label[229] , \labels[1].label[228] , 
	\labels[1].label[227] , \labels[1].label[226] , 
	\labels[1].label[225] , \labels[1].label[224] , 
	\labels[1].label[223] , \labels[1].label[222] , 
	\labels[1].label[221] , \labels[1].label[220] , 
	\labels[1].label[219] , \labels[1].label[218] , 
	\labels[1].label[217] , \labels[1].label[216] , 
	\labels[1].label[215] , \labels[1].label[214] , 
	\labels[1].label[213] , \labels[1].label[212] , 
	\labels[1].label[211] , \labels[1].label[210] , 
	\labels[1].label[209] , \labels[1].label[208] , 
	\labels[1].label[207] , \labels[1].label[206] , 
	\labels[1].label[205] , \labels[1].label[204] , 
	\labels[1].label[203] , \labels[1].label[202] , 
	\labels[1].label[201] , \labels[1].label[200] , 
	\labels[1].label[199] , \labels[1].label[198] , 
	\labels[1].label[197] , \labels[1].label[196] , 
	\labels[1].label[195] , \labels[1].label[194] , 
	\labels[1].label[193] , \labels[1].label[192] , 
	\labels[1].label[191] , \labels[1].label[190] , 
	\labels[1].label[189] , \labels[1].label[188] , 
	\labels[1].label[187] , \labels[1].label[186] , 
	\labels[1].label[185] , \labels[1].label[184] , 
	\labels[1].label[183] , \labels[1].label[182] , 
	\labels[1].label[181] , \labels[1].label[180] , 
	\labels[1].label[179] , \labels[1].label[178] , 
	\labels[1].label[177] , \labels[1].label[176] , 
	\labels[1].label[175] , \labels[1].label[174] , 
	\labels[1].label[173] , \labels[1].label[172] , 
	\labels[1].label[171] , \labels[1].label[170] , 
	\labels[1].label[169] , \labels[1].label[168] , 
	\labels[1].label[167] , \labels[1].label[166] , 
	\labels[1].label[165] , \labels[1].label[164] , 
	\labels[1].label[163] , \labels[1].label[162] , 
	\labels[1].label[161] , \labels[1].label[160] , 
	\labels[1].label[159] , \labels[1].label[158] , 
	\labels[1].label[157] , \labels[1].label[156] , 
	\labels[1].label[155] , \labels[1].label[154] , 
	\labels[1].label[153] , \labels[1].label[152] , 
	\labels[1].label[151] , \labels[1].label[150] , 
	\labels[1].label[149] , \labels[1].label[148] , 
	\labels[1].label[147] , \labels[1].label[146] , 
	\labels[1].label[145] , \labels[1].label[144] , 
	\labels[1].label[143] , \labels[1].label[142] , 
	\labels[1].label[141] , \labels[1].label[140] , 
	\labels[1].label[139] , \labels[1].label[138] , 
	\labels[1].label[137] , \labels[1].label[136] , 
	\labels[1].label[135] , \labels[1].label[134] , 
	\labels[1].label[133] , \labels[1].label[132] , 
	\labels[1].label[131] , \labels[1].label[130] , 
	\labels[1].label[129] , \labels[1].label[128] , 
	\labels[1].label[127] , \labels[1].label[126] , 
	\labels[1].label[125] , \labels[1].label[124] , 
	\labels[1].label[123] , \labels[1].label[122] , 
	\labels[1].label[121] , \labels[1].label[120] , 
	\labels[1].label[119] , \labels[1].label[118] , 
	\labels[1].label[117] , \labels[1].label[116] , 
	\labels[1].label[115] , \labels[1].label[114] , 
	\labels[1].label[113] , \labels[1].label[112] , 
	\labels[1].label[111] , \labels[1].label[110] , 
	\labels[1].label[109] , \labels[1].label[108] , 
	\labels[1].label[107] , \labels[1].label[106] , 
	\labels[1].label[105] , \labels[1].label[104] , 
	\labels[1].label[103] , \labels[1].label[102] , 
	\labels[1].label[101] , \labels[1].label[100] , 
	\labels[1].label[99] , \labels[1].label[98] , \labels[1].label[97] , 
	\labels[1].label[96] , \labels[1].label[95] , \labels[1].label[94] , 
	\labels[1].label[93] , \labels[1].label[92] , \labels[1].label[91] , 
	\labels[1].label[90] , \labels[1].label[89] , \labels[1].label[88] , 
	\labels[1].label[87] , \labels[1].label[86] , \labels[1].label[85] , 
	\labels[1].label[84] , \labels[1].label[83] , \labels[1].label[82] , 
	\labels[1].label[81] , \labels[1].label[80] , \labels[1].label[79] , 
	\labels[1].label[78] , \labels[1].label[77] , \labels[1].label[76] , 
	\labels[1].label[75] , \labels[1].label[74] , \labels[1].label[73] , 
	\labels[1].label[72] , \labels[1].label[71] , \labels[1].label[70] , 
	\labels[1].label[69] , \labels[1].label[68] , \labels[1].label[67] , 
	\labels[1].label[66] , \labels[1].label[65] , \labels[1].label[64] , 
	\labels[1].label[63] , \labels[1].label[62] , \labels[1].label[61] , 
	\labels[1].label[60] , \labels[1].label[59] , \labels[1].label[58] , 
	\labels[1].label[57] , \labels[1].label[56] , \labels[1].label[55] , 
	\labels[1].label[54] , \labels[1].label[53] , \labels[1].label[52] , 
	\labels[1].label[51] , \labels[1].label[50] , \labels[1].label[49] , 
	\labels[1].label[48] , \labels[1].label[47] , \labels[1].label[46] , 
	\labels[1].label[45] , \labels[1].label[44] , \labels[1].label[43] , 
	\labels[1].label[42] , \labels[1].label[41] , \labels[1].label[40] , 
	\labels[1].label[39] , \labels[1].label[38] , \labels[1].label[37] , 
	\labels[1].label[36] , \labels[1].label[35] , \labels[1].label[34] , 
	\labels[1].label[33] , \labels[1].label[32] , \labels[1].label[31] , 
	\labels[1].label[30] , \labels[1].label[29] , \labels[1].label[28] , 
	\labels[1].label[27] , \labels[1].label[26] , \labels[1].label[25] , 
	\labels[1].label[24] , \labels[1].label[23] , \labels[1].label[22] , 
	\labels[1].label[21] , \labels[1].label[20] , \labels[1].label[19] , 
	\labels[1].label[18] , \labels[1].label[17] , \labels[1].label[16] , 
	\labels[1].label[15] , \labels[1].label[14] , \labels[1].label[13] , 
	\labels[1].label[12] , \labels[1].label[11] , \labels[1].label[10] , 
	\labels[1].label[9] , \labels[1].label[8] , \labels[1].label[7] , 
	\labels[1].label[6] , \labels[1].label[5] , \labels[1].label[4] , 
	\labels[1].label[3] , \labels[1].label[2] , \labels[1].label[1] , 
	\labels[1].label[0] , \labels[1].delimiter_valid[0] , 
	\labels[1].delimiter[7] , \labels[1].delimiter[6] , 
	\labels[1].delimiter[5] , \labels[1].delimiter[4] , 
	\labels[1].delimiter[3] , \labels[1].delimiter[2] , 
	\labels[1].delimiter[1] , \labels[1].delimiter[0] , 
	\labels[0].guid_size[0] , \labels[0].label_size[5] , 
	\labels[0].label_size[4] , \labels[0].label_size[3] , 
	\labels[0].label_size[2] , \labels[0].label_size[1] , 
	\labels[0].label_size[0] , \labels[0].label[255] , 
	\labels[0].label[254] , \labels[0].label[253] , 
	\labels[0].label[252] , \labels[0].label[251] , 
	\labels[0].label[250] , \labels[0].label[249] , 
	\labels[0].label[248] , \labels[0].label[247] , 
	\labels[0].label[246] , \labels[0].label[245] , 
	\labels[0].label[244] , \labels[0].label[243] , 
	\labels[0].label[242] , \labels[0].label[241] , 
	\labels[0].label[240] , \labels[0].label[239] , 
	\labels[0].label[238] , \labels[0].label[237] , 
	\labels[0].label[236] , \labels[0].label[235] , 
	\labels[0].label[234] , \labels[0].label[233] , 
	\labels[0].label[232] , \labels[0].label[231] , 
	\labels[0].label[230] , \labels[0].label[229] , 
	\labels[0].label[228] , \labels[0].label[227] , 
	\labels[0].label[226] , \labels[0].label[225] , 
	\labels[0].label[224] , \labels[0].label[223] , 
	\labels[0].label[222] , \labels[0].label[221] , 
	\labels[0].label[220] , \labels[0].label[219] , 
	\labels[0].label[218] , \labels[0].label[217] , 
	\labels[0].label[216] , \labels[0].label[215] , 
	\labels[0].label[214] , \labels[0].label[213] , 
	\labels[0].label[212] , \labels[0].label[211] , 
	\labels[0].label[210] , \labels[0].label[209] , 
	\labels[0].label[208] , \labels[0].label[207] , 
	\labels[0].label[206] , \labels[0].label[205] , 
	\labels[0].label[204] , \labels[0].label[203] , 
	\labels[0].label[202] , \labels[0].label[201] , 
	\labels[0].label[200] , \labels[0].label[199] , 
	\labels[0].label[198] , \labels[0].label[197] , 
	\labels[0].label[196] , \labels[0].label[195] , 
	\labels[0].label[194] , \labels[0].label[193] , 
	\labels[0].label[192] , \labels[0].label[191] , 
	\labels[0].label[190] , \labels[0].label[189] , 
	\labels[0].label[188] , \labels[0].label[187] , 
	\labels[0].label[186] , \labels[0].label[185] , 
	\labels[0].label[184] , \labels[0].label[183] , 
	\labels[0].label[182] , \labels[0].label[181] , 
	\labels[0].label[180] , \labels[0].label[179] , 
	\labels[0].label[178] , \labels[0].label[177] , 
	\labels[0].label[176] , \labels[0].label[175] , 
	\labels[0].label[174] , \labels[0].label[173] , 
	\labels[0].label[172] , \labels[0].label[171] , 
	\labels[0].label[170] , \labels[0].label[169] , 
	\labels[0].label[168] , \labels[0].label[167] , 
	\labels[0].label[166] , \labels[0].label[165] , 
	\labels[0].label[164] , \labels[0].label[163] , 
	\labels[0].label[162] , \labels[0].label[161] , 
	\labels[0].label[160] , \labels[0].label[159] , 
	\labels[0].label[158] , \labels[0].label[157] , 
	\labels[0].label[156] , \labels[0].label[155] , 
	\labels[0].label[154] , \labels[0].label[153] , 
	\labels[0].label[152] , \labels[0].label[151] , 
	\labels[0].label[150] , \labels[0].label[149] , 
	\labels[0].label[148] , \labels[0].label[147] , 
	\labels[0].label[146] , \labels[0].label[145] , 
	\labels[0].label[144] , \labels[0].label[143] , 
	\labels[0].label[142] , \labels[0].label[141] , 
	\labels[0].label[140] , \labels[0].label[139] , 
	\labels[0].label[138] , \labels[0].label[137] , 
	\labels[0].label[136] , \labels[0].label[135] , 
	\labels[0].label[134] , \labels[0].label[133] , 
	\labels[0].label[132] , \labels[0].label[131] , 
	\labels[0].label[130] , \labels[0].label[129] , 
	\labels[0].label[128] , \labels[0].label[127] , 
	\labels[0].label[126] , \labels[0].label[125] , 
	\labels[0].label[124] , \labels[0].label[123] , 
	\labels[0].label[122] , \labels[0].label[121] , 
	\labels[0].label[120] , \labels[0].label[119] , 
	\labels[0].label[118] , \labels[0].label[117] , 
	\labels[0].label[116] , \labels[0].label[115] , 
	\labels[0].label[114] , \labels[0].label[113] , 
	\labels[0].label[112] , \labels[0].label[111] , 
	\labels[0].label[110] , \labels[0].label[109] , 
	\labels[0].label[108] , \labels[0].label[107] , 
	\labels[0].label[106] , \labels[0].label[105] , 
	\labels[0].label[104] , \labels[0].label[103] , 
	\labels[0].label[102] , \labels[0].label[101] , 
	\labels[0].label[100] , \labels[0].label[99] , \labels[0].label[98] , 
	\labels[0].label[97] , \labels[0].label[96] , \labels[0].label[95] , 
	\labels[0].label[94] , \labels[0].label[93] , \labels[0].label[92] , 
	\labels[0].label[91] , \labels[0].label[90] , \labels[0].label[89] , 
	\labels[0].label[88] , \labels[0].label[87] , \labels[0].label[86] , 
	\labels[0].label[85] , \labels[0].label[84] , \labels[0].label[83] , 
	\labels[0].label[82] , \labels[0].label[81] , \labels[0].label[80] , 
	\labels[0].label[79] , \labels[0].label[78] , \labels[0].label[77] , 
	\labels[0].label[76] , \labels[0].label[75] , \labels[0].label[74] , 
	\labels[0].label[73] , \labels[0].label[72] , \labels[0].label[71] , 
	\labels[0].label[70] , \labels[0].label[69] , \labels[0].label[68] , 
	\labels[0].label[67] , \labels[0].label[66] , \labels[0].label[65] , 
	\labels[0].label[64] , \labels[0].label[63] , \labels[0].label[62] , 
	\labels[0].label[61] , \labels[0].label[60] , \labels[0].label[59] , 
	\labels[0].label[58] , \labels[0].label[57] , \labels[0].label[56] , 
	\labels[0].label[55] , \labels[0].label[54] , \labels[0].label[53] , 
	\labels[0].label[52] , \labels[0].label[51] , \labels[0].label[50] , 
	\labels[0].label[49] , \labels[0].label[48] , \labels[0].label[47] , 
	\labels[0].label[46] , \labels[0].label[45] , \labels[0].label[44] , 
	\labels[0].label[43] , \labels[0].label[42] , \labels[0].label[41] , 
	\labels[0].label[40] , \labels[0].label[39] , \labels[0].label[38] , 
	\labels[0].label[37] , \labels[0].label[36] , \labels[0].label[35] , 
	\labels[0].label[34] , \labels[0].label[33] , \labels[0].label[32] , 
	\labels[0].label[31] , \labels[0].label[30] , \labels[0].label[29] , 
	\labels[0].label[28] , \labels[0].label[27] , \labels[0].label[26] , 
	\labels[0].label[25] , \labels[0].label[24] , \labels[0].label[23] , 
	\labels[0].label[22] , \labels[0].label[21] , \labels[0].label[20] , 
	\labels[0].label[19] , \labels[0].label[18] , \labels[0].label[17] , 
	\labels[0].label[16] , \labels[0].label[15] , \labels[0].label[14] , 
	\labels[0].label[13] , \labels[0].label[12] , \labels[0].label[11] , 
	\labels[0].label[10] , \labels[0].label[9] , \labels[0].label[8] , 
	\labels[0].label[7] , \labels[0].label[6] , \labels[0].label[5] , 
	\labels[0].label[4] , \labels[0].label[3] , \labels[0].label[2] , 
	\labels[0].label[1] , \labels[0].label[0] , 
	\labels[0].delimiter_valid[0] , \labels[0].delimiter[7] , 
	\labels[0].delimiter[6] , \labels[0].delimiter[5] , 
	\labels[0].delimiter[4] , \labels[0].delimiter[3] , 
	\labels[0].delimiter[2] , \labels[0].delimiter[1] , 
	\labels[0].delimiter[0] } ), .kme_internal_out( {
	\kme_internal_out.sot [0], \kme_internal_out.eoi [0], 
	\kme_internal_out.eot [0], \kme_internal_out.id [3], 
	\kme_internal_out.id [2], \kme_internal_out.id [1], 
	\kme_internal_out.id [0], \kme_internal_out.tdata [63], 
	\kme_internal_out.tdata [62], \kme_internal_out.tdata [61], 
	\kme_internal_out.tdata [60], \kme_internal_out.tdata [59], 
	\kme_internal_out.tdata [58], \kme_internal_out.tdata [57], 
	\kme_internal_out.tdata [56], \kme_internal_out.tdata [55], 
	\kme_internal_out.tdata [54], \kme_internal_out.tdata [53], 
	\kme_internal_out.tdata [52], \kme_internal_out.tdata [51], 
	\kme_internal_out.tdata [50], \kme_internal_out.tdata [49], 
	\kme_internal_out.tdata [48], \kme_internal_out.tdata [47], 
	\kme_internal_out.tdata [46], \kme_internal_out.tdata [45], 
	\kme_internal_out.tdata [44], \kme_internal_out.tdata [43], 
	\kme_internal_out.tdata [42], \kme_internal_out.tdata [41], 
	\kme_internal_out.tdata [40], \kme_internal_out.tdata [39], 
	\kme_internal_out.tdata [38], \kme_internal_out.tdata [37], 
	\kme_internal_out.tdata [36], \kme_internal_out.tdata [35], 
	\kme_internal_out.tdata [34], \kme_internal_out.tdata [33], 
	\kme_internal_out.tdata [32], \kme_internal_out.tdata [31], 
	\kme_internal_out.tdata [30], \kme_internal_out.tdata [29], 
	\kme_internal_out.tdata [28], \kme_internal_out.tdata [27], 
	\kme_internal_out.tdata [26], \kme_internal_out.tdata [25], 
	\kme_internal_out.tdata [24], \kme_internal_out.tdata [23], 
	\kme_internal_out.tdata [22], \kme_internal_out.tdata [21], 
	\kme_internal_out.tdata [20], \kme_internal_out.tdata [19], 
	\kme_internal_out.tdata [18], \kme_internal_out.tdata [17], 
	\kme_internal_out.tdata [16], \kme_internal_out.tdata [15], 
	\kme_internal_out.tdata [14], \kme_internal_out.tdata [13], 
	\kme_internal_out.tdata [12], \kme_internal_out.tdata [11], 
	\kme_internal_out.tdata [10], \kme_internal_out.tdata [9], 
	\kme_internal_out.tdata [8], \kme_internal_out.tdata [7], 
	\kme_internal_out.tdata [6], \kme_internal_out.tdata [5], 
	\kme_internal_out.tdata [4], \kme_internal_out.tdata [3], 
	\kme_internal_out.tdata [2], \kme_internal_out.tdata [1], 
	\kme_internal_out.tdata [0]} ), kme_internal_out_valid, 
	key_tlv_ob_full, key_tlv_ob_afull, .kop_fifo_override( {
	\kop_fifo_override.r.part0 [6], \kop_fifo_override.r.part0 [5], 
	\kop_fifo_override.r.part0 [4], \kop_fifo_override.r.part0 [3], 
	\kop_fifo_override.r.part0 [2], \kop_fifo_override.r.part0 [1], 
	\kop_fifo_override.r.part0 [0]} ), kdf_test_key_size, 
	kdf_test_mode_en);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output kme_internal_out_ack;
output key_tlv_ob_wr;
output \key_tlv_ob_tlv.insert ;
output [12:0] \key_tlv_ob_tlv.ordern ;
output [7:0] \key_tlv_ob_tlv.typen ;
output \key_tlv_ob_tlv.sot ;
output \key_tlv_ob_tlv.eot ;
output \key_tlv_ob_tlv.tlast ;
output [0:0] \key_tlv_ob_tlv.tid ;
output [7:0] \key_tlv_ob_tlv.tstrb ;
output [7:0] \key_tlv_ob_tlv.tuser ;
output [63:0] \key_tlv_ob_tlv.tdata ;
wire [105:0] key_tlv_ob_tlv;
output set_gcm_tag_fail_int;
input clk;
input rst_n;
input scan_en;
input scan_mode;
input scan_rst_n;
input \labels[7].guid_size[0] ,\labels[7].label_size[5] 
	,\labels[7].label_size[4] ,\labels[7].label_size[3] 
	,\labels[7].label_size[2] ,\labels[7].label_size[1] 
	,\labels[7].label_size[0] ,\labels[7].label[255] 
	,\labels[7].label[254] ,\labels[7].label[253] ,\labels[7].label[252] 
	,\labels[7].label[251] ,\labels[7].label[250] ,\labels[7].label[249] 
	,\labels[7].label[248] ,\labels[7].label[247] ,\labels[7].label[246] 
	,\labels[7].label[245] ,\labels[7].label[244] ,\labels[7].label[243] 
	,\labels[7].label[242] ,\labels[7].label[241] ,\labels[7].label[240] 
	,\labels[7].label[239] ,\labels[7].label[238] ,\labels[7].label[237] 
	,\labels[7].label[236] ,\labels[7].label[235] ,\labels[7].label[234] 
	,\labels[7].label[233] ,\labels[7].label[232] ,\labels[7].label[231] 
	,\labels[7].label[230] ,\labels[7].label[229] ,\labels[7].label[228] 
	,\labels[7].label[227] ,\labels[7].label[226] ,\labels[7].label[225] 
	,\labels[7].label[224] ,\labels[7].label[223] ,\labels[7].label[222] 
	,\labels[7].label[221] ,\labels[7].label[220] ,\labels[7].label[219] 
	,\labels[7].label[218] ,\labels[7].label[217] ,\labels[7].label[216] 
	,\labels[7].label[215] ,\labels[7].label[214] ,\labels[7].label[213] 
	,\labels[7].label[212] ,\labels[7].label[211] ,\labels[7].label[210] 
	,\labels[7].label[209] ,\labels[7].label[208] ,\labels[7].label[207] 
	,\labels[7].label[206] ,\labels[7].label[205] ,\labels[7].label[204] 
	,\labels[7].label[203] ,\labels[7].label[202] ,\labels[7].label[201] 
	,\labels[7].label[200] ,\labels[7].label[199] ,\labels[7].label[198] 
	,\labels[7].label[197] ,\labels[7].label[196] ,\labels[7].label[195] 
	,\labels[7].label[194] ,\labels[7].label[193] ,\labels[7].label[192] 
	,\labels[7].label[191] ,\labels[7].label[190] ,\labels[7].label[189] 
	,\labels[7].label[188] ,\labels[7].label[187] ,\labels[7].label[186] 
	,\labels[7].label[185] ,\labels[7].label[184] ,\labels[7].label[183] 
	,\labels[7].label[182] ,\labels[7].label[181] ,\labels[7].label[180] 
	,\labels[7].label[179] ,\labels[7].label[178] ,\labels[7].label[177] 
	,\labels[7].label[176] ,\labels[7].label[175] ,\labels[7].label[174] 
	,\labels[7].label[173] ,\labels[7].label[172] ,\labels[7].label[171] 
	,\labels[7].label[170] ,\labels[7].label[169] ,\labels[7].label[168] 
	,\labels[7].label[167] ,\labels[7].label[166] ,\labels[7].label[165] 
	,\labels[7].label[164] ,\labels[7].label[163] ,\labels[7].label[162] 
	,\labels[7].label[161] ,\labels[7].label[160] ,\labels[7].label[159] 
	,\labels[7].label[158] ,\labels[7].label[157] ,\labels[7].label[156] 
	,\labels[7].label[155] ,\labels[7].label[154] ,\labels[7].label[153] 
	,\labels[7].label[152] ,\labels[7].label[151] ,\labels[7].label[150] 
	,\labels[7].label[149] ,\labels[7].label[148] ,\labels[7].label[147] 
	,\labels[7].label[146] ,\labels[7].label[145] ,\labels[7].label[144] 
	,\labels[7].label[143] ,\labels[7].label[142] ,\labels[7].label[141] 
	,\labels[7].label[140] ,\labels[7].label[139] ,\labels[7].label[138] 
	,\labels[7].label[137] ,\labels[7].label[136] ,\labels[7].label[135] 
	,\labels[7].label[134] ,\labels[7].label[133] ,\labels[7].label[132] 
	,\labels[7].label[131] ,\labels[7].label[130] ,\labels[7].label[129] 
	,\labels[7].label[128] ,\labels[7].label[127] ,\labels[7].label[126] 
	,\labels[7].label[125] ,\labels[7].label[124] ,\labels[7].label[123] 
	,\labels[7].label[122] ,\labels[7].label[121] ,\labels[7].label[120] 
	,\labels[7].label[119] ,\labels[7].label[118] ,\labels[7].label[117] 
	,\labels[7].label[116] ,\labels[7].label[115] ,\labels[7].label[114] 
	,\labels[7].label[113] ,\labels[7].label[112] ,\labels[7].label[111] 
	,\labels[7].label[110] ,\labels[7].label[109] ,\labels[7].label[108] 
	,\labels[7].label[107] ,\labels[7].label[106] ,\labels[7].label[105] 
	,\labels[7].label[104] ,\labels[7].label[103] ,\labels[7].label[102] 
	,\labels[7].label[101] ,\labels[7].label[100] ,\labels[7].label[99] 
	,\labels[7].label[98] ,\labels[7].label[97] ,\labels[7].label[96] 
	,\labels[7].label[95] ,\labels[7].label[94] ,\labels[7].label[93] 
	,\labels[7].label[92] ,\labels[7].label[91] ,\labels[7].label[90] 
	,\labels[7].label[89] ,\labels[7].label[88] ,\labels[7].label[87] 
	,\labels[7].label[86] ,\labels[7].label[85] ,\labels[7].label[84] 
	,\labels[7].label[83] ,\labels[7].label[82] ,\labels[7].label[81] 
	,\labels[7].label[80] ,\labels[7].label[79] ,\labels[7].label[78] 
	,\labels[7].label[77] ,\labels[7].label[76] ,\labels[7].label[75] 
	,\labels[7].label[74] ,\labels[7].label[73] ,\labels[7].label[72] 
	,\labels[7].label[71] ,\labels[7].label[70] ,\labels[7].label[69] 
	,\labels[7].label[68] ,\labels[7].label[67] ,\labels[7].label[66] 
	,\labels[7].label[65] ,\labels[7].label[64] ,\labels[7].label[63] 
	,\labels[7].label[62] ,\labels[7].label[61] ,\labels[7].label[60] 
	,\labels[7].label[59] ,\labels[7].label[58] ,\labels[7].label[57] 
	,\labels[7].label[56] ,\labels[7].label[55] ,\labels[7].label[54] 
	,\labels[7].label[53] ,\labels[7].label[52] ,\labels[7].label[51] 
	,\labels[7].label[50] ,\labels[7].label[49] ,\labels[7].label[48] 
	,\labels[7].label[47] ,\labels[7].label[46] ,\labels[7].label[45] 
	,\labels[7].label[44] ,\labels[7].label[43] ,\labels[7].label[42] 
	,\labels[7].label[41] ,\labels[7].label[40] ,\labels[7].label[39] 
	,\labels[7].label[38] ,\labels[7].label[37] ,\labels[7].label[36] 
	,\labels[7].label[35] ,\labels[7].label[34] ,\labels[7].label[33] 
	,\labels[7].label[32] ,\labels[7].label[31] ,\labels[7].label[30] 
	,\labels[7].label[29] ,\labels[7].label[28] ,\labels[7].label[27] 
	,\labels[7].label[26] ,\labels[7].label[25] ,\labels[7].label[24] 
	,\labels[7].label[23] ,\labels[7].label[22] ,\labels[7].label[21] 
	,\labels[7].label[20] ,\labels[7].label[19] ,\labels[7].label[18] 
	,\labels[7].label[17] ,\labels[7].label[16] ,\labels[7].label[15] 
	,\labels[7].label[14] ,\labels[7].label[13] ,\labels[7].label[12] 
	,\labels[7].label[11] ,\labels[7].label[10] ,\labels[7].label[9] 
	,\labels[7].label[8] ,\labels[7].label[7] ,\labels[7].label[6] 
	,\labels[7].label[5] ,\labels[7].label[4] ,\labels[7].label[3] 
	,\labels[7].label[2] ,\labels[7].label[1] ,\labels[7].label[0] 
	,\labels[7].delimiter_valid[0] ,\labels[7].delimiter[7] 
	,\labels[7].delimiter[6] ,\labels[7].delimiter[5] 
	,\labels[7].delimiter[4] ,\labels[7].delimiter[3] 
	,\labels[7].delimiter[2] ,\labels[7].delimiter[1] 
	,\labels[7].delimiter[0] ,\labels[6].guid_size[0] 
	,\labels[6].label_size[5] ,\labels[6].label_size[4] 
	,\labels[6].label_size[3] ,\labels[6].label_size[2] 
	,\labels[6].label_size[1] ,\labels[6].label_size[0] 
	,\labels[6].label[255] ,\labels[6].label[254] ,\labels[6].label[253] 
	,\labels[6].label[252] ,\labels[6].label[251] ,\labels[6].label[250] 
	,\labels[6].label[249] ,\labels[6].label[248] ,\labels[6].label[247] 
	,\labels[6].label[246] ,\labels[6].label[245] ,\labels[6].label[244] 
	,\labels[6].label[243] ,\labels[6].label[242] ,\labels[6].label[241] 
	,\labels[6].label[240] ,\labels[6].label[239] ,\labels[6].label[238] 
	,\labels[6].label[237] ,\labels[6].label[236] ,\labels[6].label[235] 
	,\labels[6].label[234] ,\labels[6].label[233] ,\labels[6].label[232] 
	,\labels[6].label[231] ,\labels[6].label[230] ,\labels[6].label[229] 
	,\labels[6].label[228] ,\labels[6].label[227] ,\labels[6].label[226] 
	,\labels[6].label[225] ,\labels[6].label[224] ,\labels[6].label[223] 
	,\labels[6].label[222] ,\labels[6].label[221] ,\labels[6].label[220] 
	,\labels[6].label[219] ,\labels[6].label[218] ,\labels[6].label[217] 
	,\labels[6].label[216] ,\labels[6].label[215] ,\labels[6].label[214] 
	,\labels[6].label[213] ,\labels[6].label[212] ,\labels[6].label[211] 
	,\labels[6].label[210] ,\labels[6].label[209] ,\labels[6].label[208] 
	,\labels[6].label[207] ,\labels[6].label[206] ,\labels[6].label[205] 
	,\labels[6].label[204] ,\labels[6].label[203] ,\labels[6].label[202] 
	,\labels[6].label[201] ,\labels[6].label[200] ,\labels[6].label[199] 
	,\labels[6].label[198] ,\labels[6].label[197] ,\labels[6].label[196] 
	,\labels[6].label[195] ,\labels[6].label[194] ,\labels[6].label[193] 
	,\labels[6].label[192] ,\labels[6].label[191] ,\labels[6].label[190] 
	,\labels[6].label[189] ,\labels[6].label[188] ,\labels[6].label[187] 
	,\labels[6].label[186] ,\labels[6].label[185] ,\labels[6].label[184] 
	,\labels[6].label[183] ,\labels[6].label[182] ,\labels[6].label[181] 
	,\labels[6].label[180] ,\labels[6].label[179] ,\labels[6].label[178] 
	,\labels[6].label[177] ,\labels[6].label[176] ,\labels[6].label[175] 
	,\labels[6].label[174] ,\labels[6].label[173] ,\labels[6].label[172] 
	,\labels[6].label[171] ,\labels[6].label[170] ,\labels[6].label[169] 
	,\labels[6].label[168] ,\labels[6].label[167] ,\labels[6].label[166] 
	,\labels[6].label[165] ,\labels[6].label[164] ,\labels[6].label[163] 
	,\labels[6].label[162] ,\labels[6].label[161] ,\labels[6].label[160] 
	,\labels[6].label[159] ,\labels[6].label[158] ,\labels[6].label[157] 
	,\labels[6].label[156] ,\labels[6].label[155] ,\labels[6].label[154] 
	,\labels[6].label[153] ,\labels[6].label[152] ,\labels[6].label[151] 
	,\labels[6].label[150] ,\labels[6].label[149] ,\labels[6].label[148] 
	,\labels[6].label[147] ,\labels[6].label[146] ,\labels[6].label[145] 
	,\labels[6].label[144] ,\labels[6].label[143] ,\labels[6].label[142] 
	,\labels[6].label[141] ,\labels[6].label[140] ,\labels[6].label[139] 
	,\labels[6].label[138] ,\labels[6].label[137] ,\labels[6].label[136] 
	,\labels[6].label[135] ,\labels[6].label[134] ,\labels[6].label[133] 
	,\labels[6].label[132] ,\labels[6].label[131] ,\labels[6].label[130] 
	,\labels[6].label[129] ,\labels[6].label[128] ,\labels[6].label[127] 
	,\labels[6].label[126] ,\labels[6].label[125] ,\labels[6].label[124] 
	,\labels[6].label[123] ,\labels[6].label[122] ,\labels[6].label[121] 
	,\labels[6].label[120] ,\labels[6].label[119] ,\labels[6].label[118] 
	,\labels[6].label[117] ,\labels[6].label[116] ,\labels[6].label[115] 
	,\labels[6].label[114] ,\labels[6].label[113] ,\labels[6].label[112] 
	,\labels[6].label[111] ,\labels[6].label[110] ,\labels[6].label[109] 
	,\labels[6].label[108] ,\labels[6].label[107] ,\labels[6].label[106] 
	,\labels[6].label[105] ,\labels[6].label[104] ,\labels[6].label[103] 
	,\labels[6].label[102] ,\labels[6].label[101] ,\labels[6].label[100] 
	,\labels[6].label[99] ,\labels[6].label[98] ,\labels[6].label[97] 
	,\labels[6].label[96] ,\labels[6].label[95] ,\labels[6].label[94] 
	,\labels[6].label[93] ,\labels[6].label[92] ,\labels[6].label[91] 
	,\labels[6].label[90] ,\labels[6].label[89] ,\labels[6].label[88] 
	,\labels[6].label[87] ,\labels[6].label[86] ,\labels[6].label[85] 
	,\labels[6].label[84] ,\labels[6].label[83] ,\labels[6].label[82] 
	,\labels[6].label[81] ,\labels[6].label[80] ,\labels[6].label[79] 
	,\labels[6].label[78] ,\labels[6].label[77] ,\labels[6].label[76] 
	,\labels[6].label[75] ,\labels[6].label[74] ,\labels[6].label[73] 
	,\labels[6].label[72] ,\labels[6].label[71] ,\labels[6].label[70] 
	,\labels[6].label[69] ,\labels[6].label[68] ,\labels[6].label[67] 
	,\labels[6].label[66] ,\labels[6].label[65] ,\labels[6].label[64] 
	,\labels[6].label[63] ,\labels[6].label[62] ,\labels[6].label[61] 
	,\labels[6].label[60] ,\labels[6].label[59] ,\labels[6].label[58] 
	,\labels[6].label[57] ,\labels[6].label[56] ,\labels[6].label[55] 
	,\labels[6].label[54] ,\labels[6].label[53] ,\labels[6].label[52] 
	,\labels[6].label[51] ,\labels[6].label[50] ,\labels[6].label[49] 
	,\labels[6].label[48] ,\labels[6].label[47] ,\labels[6].label[46] 
	,\labels[6].label[45] ,\labels[6].label[44] ,\labels[6].label[43] 
	,\labels[6].label[42] ,\labels[6].label[41] ,\labels[6].label[40] 
	,\labels[6].label[39] ,\labels[6].label[38] ,\labels[6].label[37] 
	,\labels[6].label[36] ,\labels[6].label[35] ,\labels[6].label[34] 
	,\labels[6].label[33] ,\labels[6].label[32] ,\labels[6].label[31] 
	,\labels[6].label[30] ,\labels[6].label[29] ,\labels[6].label[28] 
	,\labels[6].label[27] ,\labels[6].label[26] ,\labels[6].label[25] 
	,\labels[6].label[24] ,\labels[6].label[23] ,\labels[6].label[22] 
	,\labels[6].label[21] ,\labels[6].label[20] ,\labels[6].label[19] 
	,\labels[6].label[18] ,\labels[6].label[17] ,\labels[6].label[16] 
	,\labels[6].label[15] ,\labels[6].label[14] ,\labels[6].label[13] 
	,\labels[6].label[12] ,\labels[6].label[11] ,\labels[6].label[10] 
	,\labels[6].label[9] ,\labels[6].label[8] ,\labels[6].label[7] 
	,\labels[6].label[6] ,\labels[6].label[5] ,\labels[6].label[4] 
	,\labels[6].label[3] ,\labels[6].label[2] ,\labels[6].label[1] 
	,\labels[6].label[0] ,\labels[6].delimiter_valid[0] 
	,\labels[6].delimiter[7] ,\labels[6].delimiter[6] 
	,\labels[6].delimiter[5] ,\labels[6].delimiter[4] 
	,\labels[6].delimiter[3] ,\labels[6].delimiter[2] 
	,\labels[6].delimiter[1] ,\labels[6].delimiter[0] 
	,\labels[5].guid_size[0] ,\labels[5].label_size[5] 
	,\labels[5].label_size[4] ,\labels[5].label_size[3] 
	,\labels[5].label_size[2] ,\labels[5].label_size[1] 
	,\labels[5].label_size[0] ,\labels[5].label[255] 
	,\labels[5].label[254] ,\labels[5].label[253] ,\labels[5].label[252] 
	,\labels[5].label[251] ,\labels[5].label[250] ,\labels[5].label[249] 
	,\labels[5].label[248] ,\labels[5].label[247] ,\labels[5].label[246] 
	,\labels[5].label[245] ,\labels[5].label[244] ,\labels[5].label[243] 
	,\labels[5].label[242] ,\labels[5].label[241] ,\labels[5].label[240] 
	,\labels[5].label[239] ,\labels[5].label[238] ,\labels[5].label[237] 
	,\labels[5].label[236] ,\labels[5].label[235] ,\labels[5].label[234] 
	,\labels[5].label[233] ,\labels[5].label[232] ,\labels[5].label[231] 
	,\labels[5].label[230] ,\labels[5].label[229] ,\labels[5].label[228] 
	,\labels[5].label[227] ,\labels[5].label[226] ,\labels[5].label[225] 
	,\labels[5].label[224] ,\labels[5].label[223] ,\labels[5].label[222] 
	,\labels[5].label[221] ,\labels[5].label[220] ,\labels[5].label[219] 
	,\labels[5].label[218] ,\labels[5].label[217] ,\labels[5].label[216] 
	,\labels[5].label[215] ,\labels[5].label[214] ,\labels[5].label[213] 
	,\labels[5].label[212] ,\labels[5].label[211] ,\labels[5].label[210] 
	,\labels[5].label[209] ,\labels[5].label[208] ,\labels[5].label[207] 
	,\labels[5].label[206] ,\labels[5].label[205] ,\labels[5].label[204] 
	,\labels[5].label[203] ,\labels[5].label[202] ,\labels[5].label[201] 
	,\labels[5].label[200] ,\labels[5].label[199] ,\labels[5].label[198] 
	,\labels[5].label[197] ,\labels[5].label[196] ,\labels[5].label[195] 
	,\labels[5].label[194] ,\labels[5].label[193] ,\labels[5].label[192] 
	,\labels[5].label[191] ,\labels[5].label[190] ,\labels[5].label[189] 
	,\labels[5].label[188] ,\labels[5].label[187] ,\labels[5].label[186] 
	,\labels[5].label[185] ,\labels[5].label[184] ,\labels[5].label[183] 
	,\labels[5].label[182] ,\labels[5].label[181] ,\labels[5].label[180] 
	,\labels[5].label[179] ,\labels[5].label[178] ,\labels[5].label[177] 
	,\labels[5].label[176] ,\labels[5].label[175] ,\labels[5].label[174] 
	,\labels[5].label[173] ,\labels[5].label[172] ,\labels[5].label[171] 
	,\labels[5].label[170] ,\labels[5].label[169] ,\labels[5].label[168] 
	,\labels[5].label[167] ,\labels[5].label[166] ,\labels[5].label[165] 
	,\labels[5].label[164] ,\labels[5].label[163] ,\labels[5].label[162] 
	,\labels[5].label[161] ,\labels[5].label[160] ,\labels[5].label[159] 
	,\labels[5].label[158] ,\labels[5].label[157] ,\labels[5].label[156] 
	,\labels[5].label[155] ,\labels[5].label[154] ,\labels[5].label[153] 
	,\labels[5].label[152] ,\labels[5].label[151] ,\labels[5].label[150] 
	,\labels[5].label[149] ,\labels[5].label[148] ,\labels[5].label[147] 
	,\labels[5].label[146] ,\labels[5].label[145] ,\labels[5].label[144] 
	,\labels[5].label[143] ,\labels[5].label[142] ,\labels[5].label[141] 
	,\labels[5].label[140] ,\labels[5].label[139] ,\labels[5].label[138] 
	,\labels[5].label[137] ,\labels[5].label[136] ,\labels[5].label[135] 
	,\labels[5].label[134] ,\labels[5].label[133] ,\labels[5].label[132] 
	,\labels[5].label[131] ,\labels[5].label[130] ,\labels[5].label[129] 
	,\labels[5].label[128] ,\labels[5].label[127] ,\labels[5].label[126] 
	,\labels[5].label[125] ,\labels[5].label[124] ,\labels[5].label[123] 
	,\labels[5].label[122] ,\labels[5].label[121] ,\labels[5].label[120] 
	,\labels[5].label[119] ,\labels[5].label[118] ,\labels[5].label[117] 
	,\labels[5].label[116] ,\labels[5].label[115] ,\labels[5].label[114] 
	,\labels[5].label[113] ,\labels[5].label[112] ,\labels[5].label[111] 
	,\labels[5].label[110] ,\labels[5].label[109] ,\labels[5].label[108] 
	,\labels[5].label[107] ,\labels[5].label[106] ,\labels[5].label[105] 
	,\labels[5].label[104] ,\labels[5].label[103] ,\labels[5].label[102] 
	,\labels[5].label[101] ,\labels[5].label[100] ,\labels[5].label[99] 
	,\labels[5].label[98] ,\labels[5].label[97] ,\labels[5].label[96] 
	,\labels[5].label[95] ,\labels[5].label[94] ,\labels[5].label[93] 
	,\labels[5].label[92] ,\labels[5].label[91] ,\labels[5].label[90] 
	,\labels[5].label[89] ,\labels[5].label[88] ,\labels[5].label[87] 
	,\labels[5].label[86] ,\labels[5].label[85] ,\labels[5].label[84] 
	,\labels[5].label[83] ,\labels[5].label[82] ,\labels[5].label[81] 
	,\labels[5].label[80] ,\labels[5].label[79] ,\labels[5].label[78] 
	,\labels[5].label[77] ,\labels[5].label[76] ,\labels[5].label[75] 
	,\labels[5].label[74] ,\labels[5].label[73] ,\labels[5].label[72] 
	,\labels[5].label[71] ,\labels[5].label[70] ,\labels[5].label[69] 
	,\labels[5].label[68] ,\labels[5].label[67] ,\labels[5].label[66] 
	,\labels[5].label[65] ,\labels[5].label[64] ,\labels[5].label[63] 
	,\labels[5].label[62] ,\labels[5].label[61] ,\labels[5].label[60] 
	,\labels[5].label[59] ,\labels[5].label[58] ,\labels[5].label[57] 
	,\labels[5].label[56] ,\labels[5].label[55] ,\labels[5].label[54] 
	,\labels[5].label[53] ,\labels[5].label[52] ,\labels[5].label[51] 
	,\labels[5].label[50] ,\labels[5].label[49] ,\labels[5].label[48] 
	,\labels[5].label[47] ,\labels[5].label[46] ,\labels[5].label[45] 
	,\labels[5].label[44] ,\labels[5].label[43] ,\labels[5].label[42] 
	,\labels[5].label[41] ,\labels[5].label[40] ,\labels[5].label[39] 
	,\labels[5].label[38] ,\labels[5].label[37] ,\labels[5].label[36] 
	,\labels[5].label[35] ,\labels[5].label[34] ,\labels[5].label[33] 
	,\labels[5].label[32] ,\labels[5].label[31] ,\labels[5].label[30] 
	,\labels[5].label[29] ,\labels[5].label[28] ,\labels[5].label[27] 
	,\labels[5].label[26] ,\labels[5].label[25] ,\labels[5].label[24] 
	,\labels[5].label[23] ,\labels[5].label[22] ,\labels[5].label[21] 
	,\labels[5].label[20] ,\labels[5].label[19] ,\labels[5].label[18] 
	,\labels[5].label[17] ,\labels[5].label[16] ,\labels[5].label[15] 
	,\labels[5].label[14] ,\labels[5].label[13] ,\labels[5].label[12] 
	,\labels[5].label[11] ,\labels[5].label[10] ,\labels[5].label[9] 
	,\labels[5].label[8] ,\labels[5].label[7] ,\labels[5].label[6] 
	,\labels[5].label[5] ,\labels[5].label[4] ,\labels[5].label[3] 
	,\labels[5].label[2] ,\labels[5].label[1] ,\labels[5].label[0] 
	,\labels[5].delimiter_valid[0] ,\labels[5].delimiter[7] 
	,\labels[5].delimiter[6] ,\labels[5].delimiter[5] 
	,\labels[5].delimiter[4] ,\labels[5].delimiter[3] 
	,\labels[5].delimiter[2] ,\labels[5].delimiter[1] 
	,\labels[5].delimiter[0] ,\labels[4].guid_size[0] 
	,\labels[4].label_size[5] ,\labels[4].label_size[4] 
	,\labels[4].label_size[3] ,\labels[4].label_size[2] 
	,\labels[4].label_size[1] ,\labels[4].label_size[0] 
	,\labels[4].label[255] ,\labels[4].label[254] ,\labels[4].label[253] 
	,\labels[4].label[252] ,\labels[4].label[251] ,\labels[4].label[250] 
	,\labels[4].label[249] ,\labels[4].label[248] ,\labels[4].label[247] 
	,\labels[4].label[246] ,\labels[4].label[245] ,\labels[4].label[244] 
	,\labels[4].label[243] ,\labels[4].label[242] ,\labels[4].label[241] 
	,\labels[4].label[240] ,\labels[4].label[239] ,\labels[4].label[238] 
	,\labels[4].label[237] ,\labels[4].label[236] ,\labels[4].label[235] 
	,\labels[4].label[234] ,\labels[4].label[233] ,\labels[4].label[232] 
	,\labels[4].label[231] ,\labels[4].label[230] ,\labels[4].label[229] 
	,\labels[4].label[228] ,\labels[4].label[227] ,\labels[4].label[226] 
	,\labels[4].label[225] ,\labels[4].label[224] ,\labels[4].label[223] 
	,\labels[4].label[222] ,\labels[4].label[221] ,\labels[4].label[220] 
	,\labels[4].label[219] ,\labels[4].label[218] ,\labels[4].label[217] 
	,\labels[4].label[216] ,\labels[4].label[215] ,\labels[4].label[214] 
	,\labels[4].label[213] ,\labels[4].label[212] ,\labels[4].label[211] 
	,\labels[4].label[210] ,\labels[4].label[209] ,\labels[4].label[208] 
	,\labels[4].label[207] ,\labels[4].label[206] ,\labels[4].label[205] 
	,\labels[4].label[204] ,\labels[4].label[203] ,\labels[4].label[202] 
	,\labels[4].label[201] ,\labels[4].label[200] ,\labels[4].label[199] 
	,\labels[4].label[198] ,\labels[4].label[197] ,\labels[4].label[196] 
	,\labels[4].label[195] ,\labels[4].label[194] ,\labels[4].label[193] 
	,\labels[4].label[192] ,\labels[4].label[191] ,\labels[4].label[190] 
	,\labels[4].label[189] ,\labels[4].label[188] ,\labels[4].label[187] 
	,\labels[4].label[186] ,\labels[4].label[185] ,\labels[4].label[184] 
	,\labels[4].label[183] ,\labels[4].label[182] ,\labels[4].label[181] 
	,\labels[4].label[180] ,\labels[4].label[179] ,\labels[4].label[178] 
	,\labels[4].label[177] ,\labels[4].label[176] ,\labels[4].label[175] 
	,\labels[4].label[174] ,\labels[4].label[173] ,\labels[4].label[172] 
	,\labels[4].label[171] ,\labels[4].label[170] ,\labels[4].label[169] 
	,\labels[4].label[168] ,\labels[4].label[167] ,\labels[4].label[166] 
	,\labels[4].label[165] ,\labels[4].label[164] ,\labels[4].label[163] 
	,\labels[4].label[162] ,\labels[4].label[161] ,\labels[4].label[160] 
	,\labels[4].label[159] ,\labels[4].label[158] ,\labels[4].label[157] 
	,\labels[4].label[156] ,\labels[4].label[155] ,\labels[4].label[154] 
	,\labels[4].label[153] ,\labels[4].label[152] ,\labels[4].label[151] 
	,\labels[4].label[150] ,\labels[4].label[149] ,\labels[4].label[148] 
	,\labels[4].label[147] ,\labels[4].label[146] ,\labels[4].label[145] 
	,\labels[4].label[144] ,\labels[4].label[143] ,\labels[4].label[142] 
	,\labels[4].label[141] ,\labels[4].label[140] ,\labels[4].label[139] 
	,\labels[4].label[138] ,\labels[4].label[137] ,\labels[4].label[136] 
	,\labels[4].label[135] ,\labels[4].label[134] ,\labels[4].label[133] 
	,\labels[4].label[132] ,\labels[4].label[131] ,\labels[4].label[130] 
	,\labels[4].label[129] ,\labels[4].label[128] ,\labels[4].label[127] 
	,\labels[4].label[126] ,\labels[4].label[125] ,\labels[4].label[124] 
	,\labels[4].label[123] ,\labels[4].label[122] ,\labels[4].label[121] 
	,\labels[4].label[120] ,\labels[4].label[119] ,\labels[4].label[118] 
	,\labels[4].label[117] ,\labels[4].label[116] ,\labels[4].label[115] 
	,\labels[4].label[114] ,\labels[4].label[113] ,\labels[4].label[112] 
	,\labels[4].label[111] ,\labels[4].label[110] ,\labels[4].label[109] 
	,\labels[4].label[108] ,\labels[4].label[107] ,\labels[4].label[106] 
	,\labels[4].label[105] ,\labels[4].label[104] ,\labels[4].label[103] 
	,\labels[4].label[102] ,\labels[4].label[101] ,\labels[4].label[100] 
	,\labels[4].label[99] ,\labels[4].label[98] ,\labels[4].label[97] 
	,\labels[4].label[96] ,\labels[4].label[95] ,\labels[4].label[94] 
	,\labels[4].label[93] ,\labels[4].label[92] ,\labels[4].label[91] 
	,\labels[4].label[90] ,\labels[4].label[89] ,\labels[4].label[88] 
	,\labels[4].label[87] ,\labels[4].label[86] ,\labels[4].label[85] 
	,\labels[4].label[84] ,\labels[4].label[83] ,\labels[4].label[82] 
	,\labels[4].label[81] ,\labels[4].label[80] ,\labels[4].label[79] 
	,\labels[4].label[78] ,\labels[4].label[77] ,\labels[4].label[76] 
	,\labels[4].label[75] ,\labels[4].label[74] ,\labels[4].label[73] 
	,\labels[4].label[72] ,\labels[4].label[71] ,\labels[4].label[70] 
	,\labels[4].label[69] ,\labels[4].label[68] ,\labels[4].label[67] 
	,\labels[4].label[66] ,\labels[4].label[65] ,\labels[4].label[64] 
	,\labels[4].label[63] ,\labels[4].label[62] ,\labels[4].label[61] 
	,\labels[4].label[60] ,\labels[4].label[59] ,\labels[4].label[58] 
	,\labels[4].label[57] ,\labels[4].label[56] ,\labels[4].label[55] 
	,\labels[4].label[54] ,\labels[4].label[53] ,\labels[4].label[52] 
	,\labels[4].label[51] ,\labels[4].label[50] ,\labels[4].label[49] 
	,\labels[4].label[48] ,\labels[4].label[47] ,\labels[4].label[46] 
	,\labels[4].label[45] ,\labels[4].label[44] ,\labels[4].label[43] 
	,\labels[4].label[42] ,\labels[4].label[41] ,\labels[4].label[40] 
	,\labels[4].label[39] ,\labels[4].label[38] ,\labels[4].label[37] 
	,\labels[4].label[36] ,\labels[4].label[35] ,\labels[4].label[34] 
	,\labels[4].label[33] ,\labels[4].label[32] ,\labels[4].label[31] 
	,\labels[4].label[30] ,\labels[4].label[29] ,\labels[4].label[28] 
	,\labels[4].label[27] ,\labels[4].label[26] ,\labels[4].label[25] 
	,\labels[4].label[24] ,\labels[4].label[23] ,\labels[4].label[22] 
	,\labels[4].label[21] ,\labels[4].label[20] ,\labels[4].label[19] 
	,\labels[4].label[18] ,\labels[4].label[17] ,\labels[4].label[16] 
	,\labels[4].label[15] ,\labels[4].label[14] ,\labels[4].label[13] 
	,\labels[4].label[12] ,\labels[4].label[11] ,\labels[4].label[10] 
	,\labels[4].label[9] ,\labels[4].label[8] ,\labels[4].label[7] 
	,\labels[4].label[6] ,\labels[4].label[5] ,\labels[4].label[4] 
	,\labels[4].label[3] ,\labels[4].label[2] ,\labels[4].label[1] 
	,\labels[4].label[0] ,\labels[4].delimiter_valid[0] 
	,\labels[4].delimiter[7] ,\labels[4].delimiter[6] 
	,\labels[4].delimiter[5] ,\labels[4].delimiter[4] 
	,\labels[4].delimiter[3] ,\labels[4].delimiter[2] 
	,\labels[4].delimiter[1] ,\labels[4].delimiter[0] 
	,\labels[3].guid_size[0] ,\labels[3].label_size[5] 
	,\labels[3].label_size[4] ,\labels[3].label_size[3] 
	,\labels[3].label_size[2] ,\labels[3].label_size[1] 
	,\labels[3].label_size[0] ,\labels[3].label[255] 
	,\labels[3].label[254] ,\labels[3].label[253] ,\labels[3].label[252] 
	,\labels[3].label[251] ,\labels[3].label[250] ,\labels[3].label[249] 
	,\labels[3].label[248] ,\labels[3].label[247] ,\labels[3].label[246] 
	,\labels[3].label[245] ,\labels[3].label[244] ,\labels[3].label[243] 
	,\labels[3].label[242] ,\labels[3].label[241] ,\labels[3].label[240] 
	,\labels[3].label[239] ,\labels[3].label[238] ,\labels[3].label[237] 
	,\labels[3].label[236] ,\labels[3].label[235] ,\labels[3].label[234] 
	,\labels[3].label[233] ,\labels[3].label[232] ,\labels[3].label[231] 
	,\labels[3].label[230] ,\labels[3].label[229] ,\labels[3].label[228] 
	,\labels[3].label[227] ,\labels[3].label[226] ,\labels[3].label[225] 
	,\labels[3].label[224] ,\labels[3].label[223] ,\labels[3].label[222] 
	,\labels[3].label[221] ,\labels[3].label[220] ,\labels[3].label[219] 
	,\labels[3].label[218] ,\labels[3].label[217] ,\labels[3].label[216] 
	,\labels[3].label[215] ,\labels[3].label[214] ,\labels[3].label[213] 
	,\labels[3].label[212] ,\labels[3].label[211] ,\labels[3].label[210] 
	,\labels[3].label[209] ,\labels[3].label[208] ,\labels[3].label[207] 
	,\labels[3].label[206] ,\labels[3].label[205] ,\labels[3].label[204] 
	,\labels[3].label[203] ,\labels[3].label[202] ,\labels[3].label[201] 
	,\labels[3].label[200] ,\labels[3].label[199] ,\labels[3].label[198] 
	,\labels[3].label[197] ,\labels[3].label[196] ,\labels[3].label[195] 
	,\labels[3].label[194] ,\labels[3].label[193] ,\labels[3].label[192] 
	,\labels[3].label[191] ,\labels[3].label[190] ,\labels[3].label[189] 
	,\labels[3].label[188] ,\labels[3].label[187] ,\labels[3].label[186] 
	,\labels[3].label[185] ,\labels[3].label[184] ,\labels[3].label[183] 
	,\labels[3].label[182] ,\labels[3].label[181] ,\labels[3].label[180] 
	,\labels[3].label[179] ,\labels[3].label[178] ,\labels[3].label[177] 
	,\labels[3].label[176] ,\labels[3].label[175] ,\labels[3].label[174] 
	,\labels[3].label[173] ,\labels[3].label[172] ,\labels[3].label[171] 
	,\labels[3].label[170] ,\labels[3].label[169] ,\labels[3].label[168] 
	,\labels[3].label[167] ,\labels[3].label[166] ,\labels[3].label[165] 
	,\labels[3].label[164] ,\labels[3].label[163] ,\labels[3].label[162] 
	,\labels[3].label[161] ,\labels[3].label[160] ,\labels[3].label[159] 
	,\labels[3].label[158] ,\labels[3].label[157] ,\labels[3].label[156] 
	,\labels[3].label[155] ,\labels[3].label[154] ,\labels[3].label[153] 
	,\labels[3].label[152] ,\labels[3].label[151] ,\labels[3].label[150] 
	,\labels[3].label[149] ,\labels[3].label[148] ,\labels[3].label[147] 
	,\labels[3].label[146] ,\labels[3].label[145] ,\labels[3].label[144] 
	,\labels[3].label[143] ,\labels[3].label[142] ,\labels[3].label[141] 
	,\labels[3].label[140] ,\labels[3].label[139] ,\labels[3].label[138] 
	,\labels[3].label[137] ,\labels[3].label[136] ,\labels[3].label[135] 
	,\labels[3].label[134] ,\labels[3].label[133] ,\labels[3].label[132] 
	,\labels[3].label[131] ,\labels[3].label[130] ,\labels[3].label[129] 
	,\labels[3].label[128] ,\labels[3].label[127] ,\labels[3].label[126] 
	,\labels[3].label[125] ,\labels[3].label[124] ,\labels[3].label[123] 
	,\labels[3].label[122] ,\labels[3].label[121] ,\labels[3].label[120] 
	,\labels[3].label[119] ,\labels[3].label[118] ,\labels[3].label[117] 
	,\labels[3].label[116] ,\labels[3].label[115] ,\labels[3].label[114] 
	,\labels[3].label[113] ,\labels[3].label[112] ,\labels[3].label[111] 
	,\labels[3].label[110] ,\labels[3].label[109] ,\labels[3].label[108] 
	,\labels[3].label[107] ,\labels[3].label[106] ,\labels[3].label[105] 
	,\labels[3].label[104] ,\labels[3].label[103] ,\labels[3].label[102] 
	,\labels[3].label[101] ,\labels[3].label[100] ,\labels[3].label[99] 
	,\labels[3].label[98] ,\labels[3].label[97] ,\labels[3].label[96] 
	,\labels[3].label[95] ,\labels[3].label[94] ,\labels[3].label[93] 
	,\labels[3].label[92] ,\labels[3].label[91] ,\labels[3].label[90] 
	,\labels[3].label[89] ,\labels[3].label[88] ,\labels[3].label[87] 
	,\labels[3].label[86] ,\labels[3].label[85] ,\labels[3].label[84] 
	,\labels[3].label[83] ,\labels[3].label[82] ,\labels[3].label[81] 
	,\labels[3].label[80] ,\labels[3].label[79] ,\labels[3].label[78] 
	,\labels[3].label[77] ,\labels[3].label[76] ,\labels[3].label[75] 
	,\labels[3].label[74] ,\labels[3].label[73] ,\labels[3].label[72] 
	,\labels[3].label[71] ,\labels[3].label[70] ,\labels[3].label[69] 
	,\labels[3].label[68] ,\labels[3].label[67] ,\labels[3].label[66] 
	,\labels[3].label[65] ,\labels[3].label[64] ,\labels[3].label[63] 
	,\labels[3].label[62] ,\labels[3].label[61] ,\labels[3].label[60] 
	,\labels[3].label[59] ,\labels[3].label[58] ,\labels[3].label[57] 
	,\labels[3].label[56] ,\labels[3].label[55] ,\labels[3].label[54] 
	,\labels[3].label[53] ,\labels[3].label[52] ,\labels[3].label[51] 
	,\labels[3].label[50] ,\labels[3].label[49] ,\labels[3].label[48] 
	,\labels[3].label[47] ,\labels[3].label[46] ,\labels[3].label[45] 
	,\labels[3].label[44] ,\labels[3].label[43] ,\labels[3].label[42] 
	,\labels[3].label[41] ,\labels[3].label[40] ,\labels[3].label[39] 
	,\labels[3].label[38] ,\labels[3].label[37] ,\labels[3].label[36] 
	,\labels[3].label[35] ,\labels[3].label[34] ,\labels[3].label[33] 
	,\labels[3].label[32] ,\labels[3].label[31] ,\labels[3].label[30] 
	,\labels[3].label[29] ,\labels[3].label[28] ,\labels[3].label[27] 
	,\labels[3].label[26] ,\labels[3].label[25] ,\labels[3].label[24] 
	,\labels[3].label[23] ,\labels[3].label[22] ,\labels[3].label[21] 
	,\labels[3].label[20] ,\labels[3].label[19] ,\labels[3].label[18] 
	,\labels[3].label[17] ,\labels[3].label[16] ,\labels[3].label[15] 
	,\labels[3].label[14] ,\labels[3].label[13] ,\labels[3].label[12] 
	,\labels[3].label[11] ,\labels[3].label[10] ,\labels[3].label[9] 
	,\labels[3].label[8] ,\labels[3].label[7] ,\labels[3].label[6] 
	,\labels[3].label[5] ,\labels[3].label[4] ,\labels[3].label[3] 
	,\labels[3].label[2] ,\labels[3].label[1] ,\labels[3].label[0] 
	,\labels[3].delimiter_valid[0] ,\labels[3].delimiter[7] 
	,\labels[3].delimiter[6] ,\labels[3].delimiter[5] 
	,\labels[3].delimiter[4] ,\labels[3].delimiter[3] 
	,\labels[3].delimiter[2] ,\labels[3].delimiter[1] 
	,\labels[3].delimiter[0] ,\labels[2].guid_size[0] 
	,\labels[2].label_size[5] ,\labels[2].label_size[4] 
	,\labels[2].label_size[3] ,\labels[2].label_size[2] 
	,\labels[2].label_size[1] ,\labels[2].label_size[0] 
	,\labels[2].label[255] ,\labels[2].label[254] ,\labels[2].label[253] 
	,\labels[2].label[252] ,\labels[2].label[251] ,\labels[2].label[250] 
	,\labels[2].label[249] ,\labels[2].label[248] ,\labels[2].label[247] 
	,\labels[2].label[246] ,\labels[2].label[245] ,\labels[2].label[244] 
	,\labels[2].label[243] ,\labels[2].label[242] ,\labels[2].label[241] 
	,\labels[2].label[240] ,\labels[2].label[239] ,\labels[2].label[238] 
	,\labels[2].label[237] ,\labels[2].label[236] ,\labels[2].label[235] 
	,\labels[2].label[234] ,\labels[2].label[233] ,\labels[2].label[232] 
	,\labels[2].label[231] ,\labels[2].label[230] ,\labels[2].label[229] 
	,\labels[2].label[228] ,\labels[2].label[227] ,\labels[2].label[226] 
	,\labels[2].label[225] ,\labels[2].label[224] ,\labels[2].label[223] 
	,\labels[2].label[222] ,\labels[2].label[221] ,\labels[2].label[220] 
	,\labels[2].label[219] ,\labels[2].label[218] ,\labels[2].label[217] 
	,\labels[2].label[216] ,\labels[2].label[215] ,\labels[2].label[214] 
	,\labels[2].label[213] ,\labels[2].label[212] ,\labels[2].label[211] 
	,\labels[2].label[210] ,\labels[2].label[209] ,\labels[2].label[208] 
	,\labels[2].label[207] ,\labels[2].label[206] ,\labels[2].label[205] 
	,\labels[2].label[204] ,\labels[2].label[203] ,\labels[2].label[202] 
	,\labels[2].label[201] ,\labels[2].label[200] ,\labels[2].label[199] 
	,\labels[2].label[198] ,\labels[2].label[197] ,\labels[2].label[196] 
	,\labels[2].label[195] ,\labels[2].label[194] ,\labels[2].label[193] 
	,\labels[2].label[192] ,\labels[2].label[191] ,\labels[2].label[190] 
	,\labels[2].label[189] ,\labels[2].label[188] ,\labels[2].label[187] 
	,\labels[2].label[186] ,\labels[2].label[185] ,\labels[2].label[184] 
	,\labels[2].label[183] ,\labels[2].label[182] ,\labels[2].label[181] 
	,\labels[2].label[180] ,\labels[2].label[179] ,\labels[2].label[178] 
	,\labels[2].label[177] ,\labels[2].label[176] ,\labels[2].label[175] 
	,\labels[2].label[174] ,\labels[2].label[173] ,\labels[2].label[172] 
	,\labels[2].label[171] ,\labels[2].label[170] ,\labels[2].label[169] 
	,\labels[2].label[168] ,\labels[2].label[167] ,\labels[2].label[166] 
	,\labels[2].label[165] ,\labels[2].label[164] ,\labels[2].label[163] 
	,\labels[2].label[162] ,\labels[2].label[161] ,\labels[2].label[160] 
	,\labels[2].label[159] ,\labels[2].label[158] ,\labels[2].label[157] 
	,\labels[2].label[156] ,\labels[2].label[155] ,\labels[2].label[154] 
	,\labels[2].label[153] ,\labels[2].label[152] ,\labels[2].label[151] 
	,\labels[2].label[150] ,\labels[2].label[149] ,\labels[2].label[148] 
	,\labels[2].label[147] ,\labels[2].label[146] ,\labels[2].label[145] 
	,\labels[2].label[144] ,\labels[2].label[143] ,\labels[2].label[142] 
	,\labels[2].label[141] ,\labels[2].label[140] ,\labels[2].label[139] 
	,\labels[2].label[138] ,\labels[2].label[137] ,\labels[2].label[136] 
	,\labels[2].label[135] ,\labels[2].label[134] ,\labels[2].label[133] 
	,\labels[2].label[132] ,\labels[2].label[131] ,\labels[2].label[130] 
	,\labels[2].label[129] ,\labels[2].label[128] ,\labels[2].label[127] 
	,\labels[2].label[126] ,\labels[2].label[125] ,\labels[2].label[124] 
	,\labels[2].label[123] ,\labels[2].label[122] ,\labels[2].label[121] 
	,\labels[2].label[120] ,\labels[2].label[119] ,\labels[2].label[118] 
	,\labels[2].label[117] ,\labels[2].label[116] ,\labels[2].label[115] 
	,\labels[2].label[114] ,\labels[2].label[113] ,\labels[2].label[112] 
	,\labels[2].label[111] ,\labels[2].label[110] ,\labels[2].label[109] 
	,\labels[2].label[108] ,\labels[2].label[107] ,\labels[2].label[106] 
	,\labels[2].label[105] ,\labels[2].label[104] ,\labels[2].label[103] 
	,\labels[2].label[102] ,\labels[2].label[101] ,\labels[2].label[100] 
	,\labels[2].label[99] ,\labels[2].label[98] ,\labels[2].label[97] 
	,\labels[2].label[96] ,\labels[2].label[95] ,\labels[2].label[94] 
	,\labels[2].label[93] ,\labels[2].label[92] ,\labels[2].label[91] 
	,\labels[2].label[90] ,\labels[2].label[89] ,\labels[2].label[88] 
	,\labels[2].label[87] ,\labels[2].label[86] ,\labels[2].label[85] 
	,\labels[2].label[84] ,\labels[2].label[83] ,\labels[2].label[82] 
	,\labels[2].label[81] ,\labels[2].label[80] ,\labels[2].label[79] 
	,\labels[2].label[78] ,\labels[2].label[77] ,\labels[2].label[76] 
	,\labels[2].label[75] ,\labels[2].label[74] ,\labels[2].label[73] 
	,\labels[2].label[72] ,\labels[2].label[71] ,\labels[2].label[70] 
	,\labels[2].label[69] ,\labels[2].label[68] ,\labels[2].label[67] 
	,\labels[2].label[66] ,\labels[2].label[65] ,\labels[2].label[64] 
	,\labels[2].label[63] ,\labels[2].label[62] ,\labels[2].label[61] 
	,\labels[2].label[60] ,\labels[2].label[59] ,\labels[2].label[58] 
	,\labels[2].label[57] ,\labels[2].label[56] ,\labels[2].label[55] 
	,\labels[2].label[54] ,\labels[2].label[53] ,\labels[2].label[52] 
	,\labels[2].label[51] ,\labels[2].label[50] ,\labels[2].label[49] 
	,\labels[2].label[48] ,\labels[2].label[47] ,\labels[2].label[46] 
	,\labels[2].label[45] ,\labels[2].label[44] ,\labels[2].label[43] 
	,\labels[2].label[42] ,\labels[2].label[41] ,\labels[2].label[40] 
	,\labels[2].label[39] ,\labels[2].label[38] ,\labels[2].label[37] 
	,\labels[2].label[36] ,\labels[2].label[35] ,\labels[2].label[34] 
	,\labels[2].label[33] ,\labels[2].label[32] ,\labels[2].label[31] 
	,\labels[2].label[30] ,\labels[2].label[29] ,\labels[2].label[28] 
	,\labels[2].label[27] ,\labels[2].label[26] ,\labels[2].label[25] 
	,\labels[2].label[24] ,\labels[2].label[23] ,\labels[2].label[22] 
	,\labels[2].label[21] ,\labels[2].label[20] ,\labels[2].label[19] 
	,\labels[2].label[18] ,\labels[2].label[17] ,\labels[2].label[16] 
	,\labels[2].label[15] ,\labels[2].label[14] ,\labels[2].label[13] 
	,\labels[2].label[12] ,\labels[2].label[11] ,\labels[2].label[10] 
	,\labels[2].label[9] ,\labels[2].label[8] ,\labels[2].label[7] 
	,\labels[2].label[6] ,\labels[2].label[5] ,\labels[2].label[4] 
	,\labels[2].label[3] ,\labels[2].label[2] ,\labels[2].label[1] 
	,\labels[2].label[0] ,\labels[2].delimiter_valid[0] 
	,\labels[2].delimiter[7] ,\labels[2].delimiter[6] 
	,\labels[2].delimiter[5] ,\labels[2].delimiter[4] 
	,\labels[2].delimiter[3] ,\labels[2].delimiter[2] 
	,\labels[2].delimiter[1] ,\labels[2].delimiter[0] 
	,\labels[1].guid_size[0] ,\labels[1].label_size[5] 
	,\labels[1].label_size[4] ,\labels[1].label_size[3] 
	,\labels[1].label_size[2] ,\labels[1].label_size[1] 
	,\labels[1].label_size[0] ,\labels[1].label[255] 
	,\labels[1].label[254] ,\labels[1].label[253] ,\labels[1].label[252] 
	,\labels[1].label[251] ,\labels[1].label[250] ,\labels[1].label[249] 
	,\labels[1].label[248] ,\labels[1].label[247] ,\labels[1].label[246] 
	,\labels[1].label[245] ,\labels[1].label[244] ,\labels[1].label[243] 
	,\labels[1].label[242] ,\labels[1].label[241] ,\labels[1].label[240] 
	,\labels[1].label[239] ,\labels[1].label[238] ,\labels[1].label[237] 
	,\labels[1].label[236] ,\labels[1].label[235] ,\labels[1].label[234] 
	,\labels[1].label[233] ,\labels[1].label[232] ,\labels[1].label[231] 
	,\labels[1].label[230] ,\labels[1].label[229] ,\labels[1].label[228] 
	,\labels[1].label[227] ,\labels[1].label[226] ,\labels[1].label[225] 
	,\labels[1].label[224] ,\labels[1].label[223] ,\labels[1].label[222] 
	,\labels[1].label[221] ,\labels[1].label[220] ,\labels[1].label[219] 
	,\labels[1].label[218] ,\labels[1].label[217] ,\labels[1].label[216] 
	,\labels[1].label[215] ,\labels[1].label[214] ,\labels[1].label[213] 
	,\labels[1].label[212] ,\labels[1].label[211] ,\labels[1].label[210] 
	,\labels[1].label[209] ,\labels[1].label[208] ,\labels[1].label[207] 
	,\labels[1].label[206] ,\labels[1].label[205] ,\labels[1].label[204] 
	,\labels[1].label[203] ,\labels[1].label[202] ,\labels[1].label[201] 
	,\labels[1].label[200] ,\labels[1].label[199] ,\labels[1].label[198] 
	,\labels[1].label[197] ,\labels[1].label[196] ,\labels[1].label[195] 
	,\labels[1].label[194] ,\labels[1].label[193] ,\labels[1].label[192] 
	,\labels[1].label[191] ,\labels[1].label[190] ,\labels[1].label[189] 
	,\labels[1].label[188] ,\labels[1].label[187] ,\labels[1].label[186] 
	,\labels[1].label[185] ,\labels[1].label[184] ,\labels[1].label[183] 
	,\labels[1].label[182] ,\labels[1].label[181] ,\labels[1].label[180] 
	,\labels[1].label[179] ,\labels[1].label[178] ,\labels[1].label[177] 
	,\labels[1].label[176] ,\labels[1].label[175] ,\labels[1].label[174] 
	,\labels[1].label[173] ,\labels[1].label[172] ,\labels[1].label[171] 
	,\labels[1].label[170] ,\labels[1].label[169] ,\labels[1].label[168] 
	,\labels[1].label[167] ,\labels[1].label[166] ,\labels[1].label[165] 
	,\labels[1].label[164] ,\labels[1].label[163] ,\labels[1].label[162] 
	,\labels[1].label[161] ,\labels[1].label[160] ,\labels[1].label[159] 
	,\labels[1].label[158] ,\labels[1].label[157] ,\labels[1].label[156] 
	,\labels[1].label[155] ,\labels[1].label[154] ,\labels[1].label[153] 
	,\labels[1].label[152] ,\labels[1].label[151] ,\labels[1].label[150] 
	,\labels[1].label[149] ,\labels[1].label[148] ,\labels[1].label[147] 
	,\labels[1].label[146] ,\labels[1].label[145] ,\labels[1].label[144] 
	,\labels[1].label[143] ,\labels[1].label[142] ,\labels[1].label[141] 
	,\labels[1].label[140] ,\labels[1].label[139] ,\labels[1].label[138] 
	,\labels[1].label[137] ,\labels[1].label[136] ,\labels[1].label[135] 
	,\labels[1].label[134] ,\labels[1].label[133] ,\labels[1].label[132] 
	,\labels[1].label[131] ,\labels[1].label[130] ,\labels[1].label[129] 
	,\labels[1].label[128] ,\labels[1].label[127] ,\labels[1].label[126] 
	,\labels[1].label[125] ,\labels[1].label[124] ,\labels[1].label[123] 
	,\labels[1].label[122] ,\labels[1].label[121] ,\labels[1].label[120] 
	,\labels[1].label[119] ,\labels[1].label[118] ,\labels[1].label[117] 
	,\labels[1].label[116] ,\labels[1].label[115] ,\labels[1].label[114] 
	,\labels[1].label[113] ,\labels[1].label[112] ,\labels[1].label[111] 
	,\labels[1].label[110] ,\labels[1].label[109] ,\labels[1].label[108] 
	,\labels[1].label[107] ,\labels[1].label[106] ,\labels[1].label[105] 
	,\labels[1].label[104] ,\labels[1].label[103] ,\labels[1].label[102] 
	,\labels[1].label[101] ,\labels[1].label[100] ,\labels[1].label[99] 
	,\labels[1].label[98] ,\labels[1].label[97] ,\labels[1].label[96] 
	,\labels[1].label[95] ,\labels[1].label[94] ,\labels[1].label[93] 
	,\labels[1].label[92] ,\labels[1].label[91] ,\labels[1].label[90] 
	,\labels[1].label[89] ,\labels[1].label[88] ,\labels[1].label[87] 
	,\labels[1].label[86] ,\labels[1].label[85] ,\labels[1].label[84] 
	,\labels[1].label[83] ,\labels[1].label[82] ,\labels[1].label[81] 
	,\labels[1].label[80] ,\labels[1].label[79] ,\labels[1].label[78] 
	,\labels[1].label[77] ,\labels[1].label[76] ,\labels[1].label[75] 
	,\labels[1].label[74] ,\labels[1].label[73] ,\labels[1].label[72] 
	,\labels[1].label[71] ,\labels[1].label[70] ,\labels[1].label[69] 
	,\labels[1].label[68] ,\labels[1].label[67] ,\labels[1].label[66] 
	,\labels[1].label[65] ,\labels[1].label[64] ,\labels[1].label[63] 
	,\labels[1].label[62] ,\labels[1].label[61] ,\labels[1].label[60] 
	,\labels[1].label[59] ,\labels[1].label[58] ,\labels[1].label[57] 
	,\labels[1].label[56] ,\labels[1].label[55] ,\labels[1].label[54] 
	,\labels[1].label[53] ,\labels[1].label[52] ,\labels[1].label[51] 
	,\labels[1].label[50] ,\labels[1].label[49] ,\labels[1].label[48] 
	,\labels[1].label[47] ,\labels[1].label[46] ,\labels[1].label[45] 
	,\labels[1].label[44] ,\labels[1].label[43] ,\labels[1].label[42] 
	,\labels[1].label[41] ,\labels[1].label[40] ,\labels[1].label[39] 
	,\labels[1].label[38] ,\labels[1].label[37] ,\labels[1].label[36] 
	,\labels[1].label[35] ,\labels[1].label[34] ,\labels[1].label[33] 
	,\labels[1].label[32] ,\labels[1].label[31] ,\labels[1].label[30] 
	,\labels[1].label[29] ,\labels[1].label[28] ,\labels[1].label[27] 
	,\labels[1].label[26] ,\labels[1].label[25] ,\labels[1].label[24] 
	,\labels[1].label[23] ,\labels[1].label[22] ,\labels[1].label[21] 
	,\labels[1].label[20] ,\labels[1].label[19] ,\labels[1].label[18] 
	,\labels[1].label[17] ,\labels[1].label[16] ,\labels[1].label[15] 
	,\labels[1].label[14] ,\labels[1].label[13] ,\labels[1].label[12] 
	,\labels[1].label[11] ,\labels[1].label[10] ,\labels[1].label[9] 
	,\labels[1].label[8] ,\labels[1].label[7] ,\labels[1].label[6] 
	,\labels[1].label[5] ,\labels[1].label[4] ,\labels[1].label[3] 
	,\labels[1].label[2] ,\labels[1].label[1] ,\labels[1].label[0] 
	,\labels[1].delimiter_valid[0] ,\labels[1].delimiter[7] 
	,\labels[1].delimiter[6] ,\labels[1].delimiter[5] 
	,\labels[1].delimiter[4] ,\labels[1].delimiter[3] 
	,\labels[1].delimiter[2] ,\labels[1].delimiter[1] 
	,\labels[1].delimiter[0] ,\labels[0].guid_size[0] 
	,\labels[0].label_size[5] ,\labels[0].label_size[4] 
	,\labels[0].label_size[3] ,\labels[0].label_size[2] 
	,\labels[0].label_size[1] ,\labels[0].label_size[0] 
	,\labels[0].label[255] ,\labels[0].label[254] ,\labels[0].label[253] 
	,\labels[0].label[252] ,\labels[0].label[251] ,\labels[0].label[250] 
	,\labels[0].label[249] ,\labels[0].label[248] ,\labels[0].label[247] 
	,\labels[0].label[246] ,\labels[0].label[245] ,\labels[0].label[244] 
	,\labels[0].label[243] ,\labels[0].label[242] ,\labels[0].label[241] 
	,\labels[0].label[240] ,\labels[0].label[239] ,\labels[0].label[238] 
	,\labels[0].label[237] ,\labels[0].label[236] ,\labels[0].label[235] 
	,\labels[0].label[234] ,\labels[0].label[233] ,\labels[0].label[232] 
	,\labels[0].label[231] ,\labels[0].label[230] ,\labels[0].label[229] 
	,\labels[0].label[228] ,\labels[0].label[227] ,\labels[0].label[226] 
	,\labels[0].label[225] ,\labels[0].label[224] ,\labels[0].label[223] 
	,\labels[0].label[222] ,\labels[0].label[221] ,\labels[0].label[220] 
	,\labels[0].label[219] ,\labels[0].label[218] ,\labels[0].label[217] 
	,\labels[0].label[216] ,\labels[0].label[215] ,\labels[0].label[214] 
	,\labels[0].label[213] ,\labels[0].label[212] ,\labels[0].label[211] 
	,\labels[0].label[210] ,\labels[0].label[209] ,\labels[0].label[208] 
	,\labels[0].label[207] ,\labels[0].label[206] ,\labels[0].label[205] 
	,\labels[0].label[204] ,\labels[0].label[203] ,\labels[0].label[202] 
	,\labels[0].label[201] ,\labels[0].label[200] ,\labels[0].label[199] 
	,\labels[0].label[198] ,\labels[0].label[197] ,\labels[0].label[196] 
	,\labels[0].label[195] ,\labels[0].label[194] ,\labels[0].label[193] 
	,\labels[0].label[192] ,\labels[0].label[191] ,\labels[0].label[190] 
	,\labels[0].label[189] ,\labels[0].label[188] ,\labels[0].label[187] 
	,\labels[0].label[186] ,\labels[0].label[185] ,\labels[0].label[184] 
	,\labels[0].label[183] ,\labels[0].label[182] ,\labels[0].label[181] 
	,\labels[0].label[180] ,\labels[0].label[179] ,\labels[0].label[178] 
	,\labels[0].label[177] ,\labels[0].label[176] ,\labels[0].label[175] 
	,\labels[0].label[174] ,\labels[0].label[173] ,\labels[0].label[172] 
	,\labels[0].label[171] ,\labels[0].label[170] ,\labels[0].label[169] 
	,\labels[0].label[168] ,\labels[0].label[167] ,\labels[0].label[166] 
	,\labels[0].label[165] ,\labels[0].label[164] ,\labels[0].label[163] 
	,\labels[0].label[162] ,\labels[0].label[161] ,\labels[0].label[160] 
	,\labels[0].label[159] ,\labels[0].label[158] ,\labels[0].label[157] 
	,\labels[0].label[156] ,\labels[0].label[155] ,\labels[0].label[154] 
	,\labels[0].label[153] ,\labels[0].label[152] ,\labels[0].label[151] 
	,\labels[0].label[150] ,\labels[0].label[149] ,\labels[0].label[148] 
	,\labels[0].label[147] ,\labels[0].label[146] ,\labels[0].label[145] 
	,\labels[0].label[144] ,\labels[0].label[143] ,\labels[0].label[142] 
	,\labels[0].label[141] ,\labels[0].label[140] ,\labels[0].label[139] 
	,\labels[0].label[138] ,\labels[0].label[137] ,\labels[0].label[136] 
	,\labels[0].label[135] ,\labels[0].label[134] ,\labels[0].label[133] 
	,\labels[0].label[132] ,\labels[0].label[131] ,\labels[0].label[130] 
	,\labels[0].label[129] ,\labels[0].label[128] ,\labels[0].label[127] 
	,\labels[0].label[126] ,\labels[0].label[125] ,\labels[0].label[124] 
	,\labels[0].label[123] ,\labels[0].label[122] ,\labels[0].label[121] 
	,\labels[0].label[120] ,\labels[0].label[119] ,\labels[0].label[118] 
	,\labels[0].label[117] ,\labels[0].label[116] ,\labels[0].label[115] 
	,\labels[0].label[114] ,\labels[0].label[113] ,\labels[0].label[112] 
	,\labels[0].label[111] ,\labels[0].label[110] ,\labels[0].label[109] 
	,\labels[0].label[108] ,\labels[0].label[107] ,\labels[0].label[106] 
	,\labels[0].label[105] ,\labels[0].label[104] ,\labels[0].label[103] 
	,\labels[0].label[102] ,\labels[0].label[101] ,\labels[0].label[100] 
	,\labels[0].label[99] ,\labels[0].label[98] ,\labels[0].label[97] 
	,\labels[0].label[96] ,\labels[0].label[95] ,\labels[0].label[94] 
	,\labels[0].label[93] ,\labels[0].label[92] ,\labels[0].label[91] 
	,\labels[0].label[90] ,\labels[0].label[89] ,\labels[0].label[88] 
	,\labels[0].label[87] ,\labels[0].label[86] ,\labels[0].label[85] 
	,\labels[0].label[84] ,\labels[0].label[83] ,\labels[0].label[82] 
	,\labels[0].label[81] ,\labels[0].label[80] ,\labels[0].label[79] 
	,\labels[0].label[78] ,\labels[0].label[77] ,\labels[0].label[76] 
	,\labels[0].label[75] ,\labels[0].label[74] ,\labels[0].label[73] 
	,\labels[0].label[72] ,\labels[0].label[71] ,\labels[0].label[70] 
	,\labels[0].label[69] ,\labels[0].label[68] ,\labels[0].label[67] 
	,\labels[0].label[66] ,\labels[0].label[65] ,\labels[0].label[64] 
	,\labels[0].label[63] ,\labels[0].label[62] ,\labels[0].label[61] 
	,\labels[0].label[60] ,\labels[0].label[59] ,\labels[0].label[58] 
	,\labels[0].label[57] ,\labels[0].label[56] ,\labels[0].label[55] 
	,\labels[0].label[54] ,\labels[0].label[53] ,\labels[0].label[52] 
	,\labels[0].label[51] ,\labels[0].label[50] ,\labels[0].label[49] 
	,\labels[0].label[48] ,\labels[0].label[47] ,\labels[0].label[46] 
	,\labels[0].label[45] ,\labels[0].label[44] ,\labels[0].label[43] 
	,\labels[0].label[42] ,\labels[0].label[41] ,\labels[0].label[40] 
	,\labels[0].label[39] ,\labels[0].label[38] ,\labels[0].label[37] 
	,\labels[0].label[36] ,\labels[0].label[35] ,\labels[0].label[34] 
	,\labels[0].label[33] ,\labels[0].label[32] ,\labels[0].label[31] 
	,\labels[0].label[30] ,\labels[0].label[29] ,\labels[0].label[28] 
	,\labels[0].label[27] ,\labels[0].label[26] ,\labels[0].label[25] 
	,\labels[0].label[24] ,\labels[0].label[23] ,\labels[0].label[22] 
	,\labels[0].label[21] ,\labels[0].label[20] ,\labels[0].label[19] 
	,\labels[0].label[18] ,\labels[0].label[17] ,\labels[0].label[16] 
	,\labels[0].label[15] ,\labels[0].label[14] ,\labels[0].label[13] 
	,\labels[0].label[12] ,\labels[0].label[11] ,\labels[0].label[10] 
	,\labels[0].label[9] ,\labels[0].label[8] ,\labels[0].label[7] 
	,\labels[0].label[6] ,\labels[0].label[5] ,\labels[0].label[4] 
	,\labels[0].label[3] ,\labels[0].label[2] ,\labels[0].label[1] 
	,\labels[0].label[0] ,\labels[0].delimiter_valid[0] 
	,\labels[0].delimiter[7] ,\labels[0].delimiter[6] 
	,\labels[0].delimiter[5] ,\labels[0].delimiter[4] 
	,\labels[0].delimiter[3] ,\labels[0].delimiter[2] 
	,\labels[0].delimiter[1] ,\labels[0].delimiter[0] ;
input [0:0] \kme_internal_out.sot ;
input [0:0] \kme_internal_out.eoi ;
input [0:0] \kme_internal_out.eot ;
input [3:0] \kme_internal_out.id ;
input [63:0] \kme_internal_out.tdata ;
wire [70:0] kme_internal_out;
input kme_internal_out_valid;
input key_tlv_ob_full;
input key_tlv_ob_afull;
input [6:0] \kop_fifo_override.r.part0 ;
wire \kop_fifo_override.f.gcm_status_data_fifo ;
wire \kop_fifo_override.f.tlv_sb_data_fifo ;
wire \kop_fifo_override.f.kdf_cmd_fifo ;
wire \kop_fifo_override.f.kdfstream_cmd_fifo ;
wire \kop_fifo_override.f.keyfilter_cmd_fifo ;
wire \kop_fifo_override.f.gcm_tag_data_fifo ;
wire \kop_fifo_override.f.gcm_cmd_fifo ;
wire [6:0] kop_fifo_override;
input [31:0] kdf_test_key_size;
input kdf_test_mode_en;
wire [610:0] cmdfifo_gcm_cmd;
wire cmdfifo_gcm_valid;
wire [3:0] cmdfifo_kdf_cmd;
wire cmdfifo_kdf_valid;
wire [262:0] cmdfifo_kdfstream_cmd;
wire cmdfifo_kdfstream_valid;
wire [0:0] cmdfifo_keyfilter_cmd;
wire cmdfifo_keyfilter_valid;
wire gcm_cmd_in_stall;
wire gcm_cmd_in_valid;
wire gcm_cmdfifo_ack;
wire [127:0] gcm_kdf_data;
wire gcm_kdf_eof;
wire gcm_kdf_valid;
wire gcm_status_data_in_stall;
wire gcm_status_data_in_valid;
wire [0:0] gcm_status_data_out;
wire gcm_status_data_out_ack;
wire gcm_status_data_out_valid;
wire [95:0] gcm_tag_data_in;
wire gcm_tag_data_in_stall;
wire gcm_tag_data_in_valid;
wire [95:0] gcm_tag_data_out;
wire gcm_tag_data_out_ack;
wire gcm_tag_data_out_valid;
wire gcm_upsizer_stall;
wire [63:0] inspector_upsizer_data;
wire inspector_upsizer_eof;
wire inspector_upsizer_valid;
wire kdf_cmd_in_stall;
wire kdf_cmd_in_valid;
wire kdf_cmdfifo_ack;
wire kdf_gcm_stall;
wire [63:0] kdf_keybuilder_data;
wire kdf_keybuilder_valid;
wire kdfstream_cmd_in_stall;
wire kdfstream_cmd_in_valid;
wire kdfstream_cmdfifo_ack;
wire keybuilder_kdf_stall;
wire keyfilter_cmd_in_stall;
wire keyfilter_cmd_in_valid;
wire keyfilter_cmdfifo_ack;
wire [63:0] tlv_sb_data_in;
wire tlv_sb_data_in_stall;
wire tlv_sb_data_in_valid;
wire [63:0] tlv_sb_data_out;
wire tlv_sb_data_out_ack;
wire tlv_sb_data_out_valid;
wire [127:0] upsizer_gcm_data;
wire upsizer_gcm_eof;
wire upsizer_gcm_valid;
wire upsizer_inspector_stall;
wire [0:105] _zy_simnet_key_tlv_ob_tlv_0_w$;
wire [0:610] _zy_simnet_gcm_cmd_in_1_w$;
wire _zy_simnet_keyfilter_cmd_in_2_w$;
wire [0:262] _zy_simnet_kdfstream_cmd_in_3_w$;
wire [0:3] _zy_simnet_kdf_cmd_in_4_w$;
wire _zy_simnet_gcm_status_data_in_5_w$;
wire [0:105] _zy_simnet_key_tlv_ob_tlv_6_w$;
wire _zy_simnet_dio_7;
wire _zy_simnet_dio_8;
wire [0:610] _zy_simnet_gcm_cmd_in_9_w$;
wire _zy_simnet_dio_10;
wire _zy_simnet_dio_11;
wire _zy_simnet_keyfilter_cmd_in_12_w$;
wire _zy_simnet_dio_13;
wire _zy_simnet_dio_14;
wire [0:3] _zy_simnet_kdf_cmd_in_15_w$;
wire _zy_simnet_dio_16;
wire _zy_simnet_dio_17;
wire [0:262] _zy_simnet_kdfstream_cmd_in_18_w$;
wire _zy_simnet_dio_19;
wire _zy_simnet_dio_20;
wire _zy_simnet_dio_21;
wire _zy_simnet_dio_22;
wire _zy_simnet_dio_23;
wire _zy_simnet_dio_24;
wire _zy_simnet_gcm_status_data_in_25_w$;
wire [610:0] gcm_cmd_in;
wire [0:0] gcm_status_data_in;
wire [3:0] kdf_cmd_in;
wire [262:0] kdfstream_cmd_in;
wire [0:0] keyfilter_cmd_in;
wire [255:0] \gcm_cmd_in.key0 ;
wire [255:0] \gcm_cmd_in.key1 ;
wire [95:0] \gcm_cmd_in.iv ;
wire [2:0] \gcm_cmd_in.op ;
wire [0:0] \gcm_status_data_in.tag_mismatch ;
wire [0:0] \kdf_cmd_in.kdf_dek_iter ;
wire [0:0] \kdf_cmd_in.combo_mode ;
wire [0:0] \kdf_cmd_in.dek_key_op ;
wire [0:0] \kdf_cmd_in.dak_key_op ;
wire [0:0] \kdfstream_cmd_in.combo_mode ;
wire [0:0] \kdfstream_cmd_in.skip ;
wire [255:0] \kdfstream_cmd_in.guid ;
wire [2:0] \kdfstream_cmd_in.label_index ;
wire [1:0] \kdfstream_cmd_in.num_iter ;
wire [0:0] \keyfilter_cmd_in.combo_mode ;
tran (key_tlv_ob_tlv[105], \key_tlv_ob_tlv.insert );
tran (key_tlv_ob_tlv[104], \key_tlv_ob_tlv.ordern [12]);
tran (key_tlv_ob_tlv[103], \key_tlv_ob_tlv.ordern [11]);
tran (key_tlv_ob_tlv[102], \key_tlv_ob_tlv.ordern [10]);
tran (key_tlv_ob_tlv[101], \key_tlv_ob_tlv.ordern [9]);
tran (key_tlv_ob_tlv[100], \key_tlv_ob_tlv.ordern [8]);
tran (key_tlv_ob_tlv[99], \key_tlv_ob_tlv.ordern [7]);
tran (key_tlv_ob_tlv[98], \key_tlv_ob_tlv.ordern [6]);
tran (key_tlv_ob_tlv[97], \key_tlv_ob_tlv.ordern [5]);
tran (key_tlv_ob_tlv[96], \key_tlv_ob_tlv.ordern [4]);
tran (key_tlv_ob_tlv[95], \key_tlv_ob_tlv.ordern [3]);
tran (key_tlv_ob_tlv[94], \key_tlv_ob_tlv.ordern [2]);
tran (key_tlv_ob_tlv[93], \key_tlv_ob_tlv.ordern [1]);
tran (key_tlv_ob_tlv[92], \key_tlv_ob_tlv.ordern [0]);
tran (key_tlv_ob_tlv[91], \key_tlv_ob_tlv.typen [7]);
tran (key_tlv_ob_tlv[90], \key_tlv_ob_tlv.typen [6]);
tran (key_tlv_ob_tlv[89], \key_tlv_ob_tlv.typen [5]);
tran (key_tlv_ob_tlv[88], \key_tlv_ob_tlv.typen [4]);
tran (key_tlv_ob_tlv[87], \key_tlv_ob_tlv.typen [3]);
tran (key_tlv_ob_tlv[86], \key_tlv_ob_tlv.typen [2]);
tran (key_tlv_ob_tlv[85], \key_tlv_ob_tlv.typen [1]);
tran (key_tlv_ob_tlv[84], \key_tlv_ob_tlv.typen [0]);
tran (key_tlv_ob_tlv[83], \key_tlv_ob_tlv.sot );
tran (key_tlv_ob_tlv[82], \key_tlv_ob_tlv.eot );
tran (key_tlv_ob_tlv[81], \key_tlv_ob_tlv.tlast );
tran (key_tlv_ob_tlv[80], \key_tlv_ob_tlv.tid [0]);
tran (key_tlv_ob_tlv[79], \key_tlv_ob_tlv.tstrb [7]);
tran (key_tlv_ob_tlv[78], \key_tlv_ob_tlv.tstrb [6]);
tran (key_tlv_ob_tlv[77], \key_tlv_ob_tlv.tstrb [5]);
tran (key_tlv_ob_tlv[76], \key_tlv_ob_tlv.tstrb [4]);
tran (key_tlv_ob_tlv[75], \key_tlv_ob_tlv.tstrb [3]);
tran (key_tlv_ob_tlv[74], \key_tlv_ob_tlv.tstrb [2]);
tran (key_tlv_ob_tlv[73], \key_tlv_ob_tlv.tstrb [1]);
tran (key_tlv_ob_tlv[72], \key_tlv_ob_tlv.tstrb [0]);
tran (key_tlv_ob_tlv[71], \key_tlv_ob_tlv.tuser [7]);
tran (key_tlv_ob_tlv[70], \key_tlv_ob_tlv.tuser [6]);
tran (key_tlv_ob_tlv[69], \key_tlv_ob_tlv.tuser [5]);
tran (key_tlv_ob_tlv[68], \key_tlv_ob_tlv.tuser [4]);
tran (key_tlv_ob_tlv[67], \key_tlv_ob_tlv.tuser [3]);
tran (key_tlv_ob_tlv[66], \key_tlv_ob_tlv.tuser [2]);
tran (key_tlv_ob_tlv[65], \key_tlv_ob_tlv.tuser [1]);
tran (key_tlv_ob_tlv[64], \key_tlv_ob_tlv.tuser [0]);
tran (key_tlv_ob_tlv[63], \key_tlv_ob_tlv.tdata [63]);
tran (key_tlv_ob_tlv[62], \key_tlv_ob_tlv.tdata [62]);
tran (key_tlv_ob_tlv[61], \key_tlv_ob_tlv.tdata [61]);
tran (key_tlv_ob_tlv[60], \key_tlv_ob_tlv.tdata [60]);
tran (key_tlv_ob_tlv[59], \key_tlv_ob_tlv.tdata [59]);
tran (key_tlv_ob_tlv[58], \key_tlv_ob_tlv.tdata [58]);
tran (key_tlv_ob_tlv[57], \key_tlv_ob_tlv.tdata [57]);
tran (key_tlv_ob_tlv[56], \key_tlv_ob_tlv.tdata [56]);
tran (key_tlv_ob_tlv[55], \key_tlv_ob_tlv.tdata [55]);
tran (key_tlv_ob_tlv[54], \key_tlv_ob_tlv.tdata [54]);
tran (key_tlv_ob_tlv[53], \key_tlv_ob_tlv.tdata [53]);
tran (key_tlv_ob_tlv[52], \key_tlv_ob_tlv.tdata [52]);
tran (key_tlv_ob_tlv[51], \key_tlv_ob_tlv.tdata [51]);
tran (key_tlv_ob_tlv[50], \key_tlv_ob_tlv.tdata [50]);
tran (key_tlv_ob_tlv[49], \key_tlv_ob_tlv.tdata [49]);
tran (key_tlv_ob_tlv[48], \key_tlv_ob_tlv.tdata [48]);
tran (key_tlv_ob_tlv[47], \key_tlv_ob_tlv.tdata [47]);
tran (key_tlv_ob_tlv[46], \key_tlv_ob_tlv.tdata [46]);
tran (key_tlv_ob_tlv[45], \key_tlv_ob_tlv.tdata [45]);
tran (key_tlv_ob_tlv[44], \key_tlv_ob_tlv.tdata [44]);
tran (key_tlv_ob_tlv[43], \key_tlv_ob_tlv.tdata [43]);
tran (key_tlv_ob_tlv[42], \key_tlv_ob_tlv.tdata [42]);
tran (key_tlv_ob_tlv[41], \key_tlv_ob_tlv.tdata [41]);
tran (key_tlv_ob_tlv[40], \key_tlv_ob_tlv.tdata [40]);
tran (key_tlv_ob_tlv[39], \key_tlv_ob_tlv.tdata [39]);
tran (key_tlv_ob_tlv[38], \key_tlv_ob_tlv.tdata [38]);
tran (key_tlv_ob_tlv[37], \key_tlv_ob_tlv.tdata [37]);
tran (key_tlv_ob_tlv[36], \key_tlv_ob_tlv.tdata [36]);
tran (key_tlv_ob_tlv[35], \key_tlv_ob_tlv.tdata [35]);
tran (key_tlv_ob_tlv[34], \key_tlv_ob_tlv.tdata [34]);
tran (key_tlv_ob_tlv[33], \key_tlv_ob_tlv.tdata [33]);
tran (key_tlv_ob_tlv[32], \key_tlv_ob_tlv.tdata [32]);
tran (key_tlv_ob_tlv[31], \key_tlv_ob_tlv.tdata [31]);
tran (key_tlv_ob_tlv[30], \key_tlv_ob_tlv.tdata [30]);
tran (key_tlv_ob_tlv[29], \key_tlv_ob_tlv.tdata [29]);
tran (key_tlv_ob_tlv[28], \key_tlv_ob_tlv.tdata [28]);
tran (key_tlv_ob_tlv[27], \key_tlv_ob_tlv.tdata [27]);
tran (key_tlv_ob_tlv[26], \key_tlv_ob_tlv.tdata [26]);
tran (key_tlv_ob_tlv[25], \key_tlv_ob_tlv.tdata [25]);
tran (key_tlv_ob_tlv[24], \key_tlv_ob_tlv.tdata [24]);
tran (key_tlv_ob_tlv[23], \key_tlv_ob_tlv.tdata [23]);
tran (key_tlv_ob_tlv[22], \key_tlv_ob_tlv.tdata [22]);
tran (key_tlv_ob_tlv[21], \key_tlv_ob_tlv.tdata [21]);
tran (key_tlv_ob_tlv[20], \key_tlv_ob_tlv.tdata [20]);
tran (key_tlv_ob_tlv[19], \key_tlv_ob_tlv.tdata [19]);
tran (key_tlv_ob_tlv[18], \key_tlv_ob_tlv.tdata [18]);
tran (key_tlv_ob_tlv[17], \key_tlv_ob_tlv.tdata [17]);
tran (key_tlv_ob_tlv[16], \key_tlv_ob_tlv.tdata [16]);
tran (key_tlv_ob_tlv[15], \key_tlv_ob_tlv.tdata [15]);
tran (key_tlv_ob_tlv[14], \key_tlv_ob_tlv.tdata [14]);
tran (key_tlv_ob_tlv[13], \key_tlv_ob_tlv.tdata [13]);
tran (key_tlv_ob_tlv[12], \key_tlv_ob_tlv.tdata [12]);
tran (key_tlv_ob_tlv[11], \key_tlv_ob_tlv.tdata [11]);
tran (key_tlv_ob_tlv[10], \key_tlv_ob_tlv.tdata [10]);
tran (key_tlv_ob_tlv[9], \key_tlv_ob_tlv.tdata [9]);
tran (key_tlv_ob_tlv[8], \key_tlv_ob_tlv.tdata [8]);
tran (key_tlv_ob_tlv[7], \key_tlv_ob_tlv.tdata [7]);
tran (key_tlv_ob_tlv[6], \key_tlv_ob_tlv.tdata [6]);
tran (key_tlv_ob_tlv[5], \key_tlv_ob_tlv.tdata [5]);
tran (key_tlv_ob_tlv[4], \key_tlv_ob_tlv.tdata [4]);
tran (key_tlv_ob_tlv[3], \key_tlv_ob_tlv.tdata [3]);
tran (key_tlv_ob_tlv[2], \key_tlv_ob_tlv.tdata [2]);
tran (key_tlv_ob_tlv[1], \key_tlv_ob_tlv.tdata [1]);
tran (key_tlv_ob_tlv[0], \key_tlv_ob_tlv.tdata [0]);
tran (\labels[0][0] , \labels[0].delimiter[0] );
tran (\labels[0][1] , \labels[0].delimiter[1] );
tran (\labels[0][2] , \labels[0].delimiter[2] );
tran (\labels[0][3] , \labels[0].delimiter[3] );
tran (\labels[0][4] , \labels[0].delimiter[4] );
tran (\labels[0][5] , \labels[0].delimiter[5] );
tran (\labels[0][6] , \labels[0].delimiter[6] );
tran (\labels[0][7] , \labels[0].delimiter[7] );
tran (\labels[0][8] , \labels[0].delimiter_valid[0] );
tran (\labels[0][9] , \labels[0].label[0] );
tran (\labels[0][10] , \labels[0].label[1] );
tran (\labels[0][11] , \labels[0].label[2] );
tran (\labels[0][12] , \labels[0].label[3] );
tran (\labels[0][13] , \labels[0].label[4] );
tran (\labels[0][14] , \labels[0].label[5] );
tran (\labels[0][15] , \labels[0].label[6] );
tran (\labels[0][16] , \labels[0].label[7] );
tran (\labels[0][17] , \labels[0].label[8] );
tran (\labels[0][18] , \labels[0].label[9] );
tran (\labels[0][19] , \labels[0].label[10] );
tran (\labels[0][20] , \labels[0].label[11] );
tran (\labels[0][21] , \labels[0].label[12] );
tran (\labels[0][22] , \labels[0].label[13] );
tran (\labels[0][23] , \labels[0].label[14] );
tran (\labels[0][24] , \labels[0].label[15] );
tran (\labels[0][25] , \labels[0].label[16] );
tran (\labels[0][26] , \labels[0].label[17] );
tran (\labels[0][27] , \labels[0].label[18] );
tran (\labels[0][28] , \labels[0].label[19] );
tran (\labels[0][29] , \labels[0].label[20] );
tran (\labels[0][30] , \labels[0].label[21] );
tran (\labels[0][31] , \labels[0].label[22] );
tran (\labels[0][32] , \labels[0].label[23] );
tran (\labels[0][33] , \labels[0].label[24] );
tran (\labels[0][34] , \labels[0].label[25] );
tran (\labels[0][35] , \labels[0].label[26] );
tran (\labels[0][36] , \labels[0].label[27] );
tran (\labels[0][37] , \labels[0].label[28] );
tran (\labels[0][38] , \labels[0].label[29] );
tran (\labels[0][39] , \labels[0].label[30] );
tran (\labels[0][40] , \labels[0].label[31] );
tran (\labels[0][41] , \labels[0].label[32] );
tran (\labels[0][42] , \labels[0].label[33] );
tran (\labels[0][43] , \labels[0].label[34] );
tran (\labels[0][44] , \labels[0].label[35] );
tran (\labels[0][45] , \labels[0].label[36] );
tran (\labels[0][46] , \labels[0].label[37] );
tran (\labels[0][47] , \labels[0].label[38] );
tran (\labels[0][48] , \labels[0].label[39] );
tran (\labels[0][49] , \labels[0].label[40] );
tran (\labels[0][50] , \labels[0].label[41] );
tran (\labels[0][51] , \labels[0].label[42] );
tran (\labels[0][52] , \labels[0].label[43] );
tran (\labels[0][53] , \labels[0].label[44] );
tran (\labels[0][54] , \labels[0].label[45] );
tran (\labels[0][55] , \labels[0].label[46] );
tran (\labels[0][56] , \labels[0].label[47] );
tran (\labels[0][57] , \labels[0].label[48] );
tran (\labels[0][58] , \labels[0].label[49] );
tran (\labels[0][59] , \labels[0].label[50] );
tran (\labels[0][60] , \labels[0].label[51] );
tran (\labels[0][61] , \labels[0].label[52] );
tran (\labels[0][62] , \labels[0].label[53] );
tran (\labels[0][63] , \labels[0].label[54] );
tran (\labels[0][64] , \labels[0].label[55] );
tran (\labels[0][65] , \labels[0].label[56] );
tran (\labels[0][66] , \labels[0].label[57] );
tran (\labels[0][67] , \labels[0].label[58] );
tran (\labels[0][68] , \labels[0].label[59] );
tran (\labels[0][69] , \labels[0].label[60] );
tran (\labels[0][70] , \labels[0].label[61] );
tran (\labels[0][71] , \labels[0].label[62] );
tran (\labels[0][72] , \labels[0].label[63] );
tran (\labels[0][73] , \labels[0].label[64] );
tran (\labels[0][74] , \labels[0].label[65] );
tran (\labels[0][75] , \labels[0].label[66] );
tran (\labels[0][76] , \labels[0].label[67] );
tran (\labels[0][77] , \labels[0].label[68] );
tran (\labels[0][78] , \labels[0].label[69] );
tran (\labels[0][79] , \labels[0].label[70] );
tran (\labels[0][80] , \labels[0].label[71] );
tran (\labels[0][81] , \labels[0].label[72] );
tran (\labels[0][82] , \labels[0].label[73] );
tran (\labels[0][83] , \labels[0].label[74] );
tran (\labels[0][84] , \labels[0].label[75] );
tran (\labels[0][85] , \labels[0].label[76] );
tran (\labels[0][86] , \labels[0].label[77] );
tran (\labels[0][87] , \labels[0].label[78] );
tran (\labels[0][88] , \labels[0].label[79] );
tran (\labels[0][89] , \labels[0].label[80] );
tran (\labels[0][90] , \labels[0].label[81] );
tran (\labels[0][91] , \labels[0].label[82] );
tran (\labels[0][92] , \labels[0].label[83] );
tran (\labels[0][93] , \labels[0].label[84] );
tran (\labels[0][94] , \labels[0].label[85] );
tran (\labels[0][95] , \labels[0].label[86] );
tran (\labels[0][96] , \labels[0].label[87] );
tran (\labels[0][97] , \labels[0].label[88] );
tran (\labels[0][98] , \labels[0].label[89] );
tran (\labels[0][99] , \labels[0].label[90] );
tran (\labels[0][100] , \labels[0].label[91] );
tran (\labels[0][101] , \labels[0].label[92] );
tran (\labels[0][102] , \labels[0].label[93] );
tran (\labels[0][103] , \labels[0].label[94] );
tran (\labels[0][104] , \labels[0].label[95] );
tran (\labels[0][105] , \labels[0].label[96] );
tran (\labels[0][106] , \labels[0].label[97] );
tran (\labels[0][107] , \labels[0].label[98] );
tran (\labels[0][108] , \labels[0].label[99] );
tran (\labels[0][109] , \labels[0].label[100] );
tran (\labels[0][110] , \labels[0].label[101] );
tran (\labels[0][111] , \labels[0].label[102] );
tran (\labels[0][112] , \labels[0].label[103] );
tran (\labels[0][113] , \labels[0].label[104] );
tran (\labels[0][114] , \labels[0].label[105] );
tran (\labels[0][115] , \labels[0].label[106] );
tran (\labels[0][116] , \labels[0].label[107] );
tran (\labels[0][117] , \labels[0].label[108] );
tran (\labels[0][118] , \labels[0].label[109] );
tran (\labels[0][119] , \labels[0].label[110] );
tran (\labels[0][120] , \labels[0].label[111] );
tran (\labels[0][121] , \labels[0].label[112] );
tran (\labels[0][122] , \labels[0].label[113] );
tran (\labels[0][123] , \labels[0].label[114] );
tran (\labels[0][124] , \labels[0].label[115] );
tran (\labels[0][125] , \labels[0].label[116] );
tran (\labels[0][126] , \labels[0].label[117] );
tran (\labels[0][127] , \labels[0].label[118] );
tran (\labels[0][128] , \labels[0].label[119] );
tran (\labels[0][129] , \labels[0].label[120] );
tran (\labels[0][130] , \labels[0].label[121] );
tran (\labels[0][131] , \labels[0].label[122] );
tran (\labels[0][132] , \labels[0].label[123] );
tran (\labels[0][133] , \labels[0].label[124] );
tran (\labels[0][134] , \labels[0].label[125] );
tran (\labels[0][135] , \labels[0].label[126] );
tran (\labels[0][136] , \labels[0].label[127] );
tran (\labels[0][137] , \labels[0].label[128] );
tran (\labels[0][138] , \labels[0].label[129] );
tran (\labels[0][139] , \labels[0].label[130] );
tran (\labels[0][140] , \labels[0].label[131] );
tran (\labels[0][141] , \labels[0].label[132] );
tran (\labels[0][142] , \labels[0].label[133] );
tran (\labels[0][143] , \labels[0].label[134] );
tran (\labels[0][144] , \labels[0].label[135] );
tran (\labels[0][145] , \labels[0].label[136] );
tran (\labels[0][146] , \labels[0].label[137] );
tran (\labels[0][147] , \labels[0].label[138] );
tran (\labels[0][148] , \labels[0].label[139] );
tran (\labels[0][149] , \labels[0].label[140] );
tran (\labels[0][150] , \labels[0].label[141] );
tran (\labels[0][151] , \labels[0].label[142] );
tran (\labels[0][152] , \labels[0].label[143] );
tran (\labels[0][153] , \labels[0].label[144] );
tran (\labels[0][154] , \labels[0].label[145] );
tran (\labels[0][155] , \labels[0].label[146] );
tran (\labels[0][156] , \labels[0].label[147] );
tran (\labels[0][157] , \labels[0].label[148] );
tran (\labels[0][158] , \labels[0].label[149] );
tran (\labels[0][159] , \labels[0].label[150] );
tran (\labels[0][160] , \labels[0].label[151] );
tran (\labels[0][161] , \labels[0].label[152] );
tran (\labels[0][162] , \labels[0].label[153] );
tran (\labels[0][163] , \labels[0].label[154] );
tran (\labels[0][164] , \labels[0].label[155] );
tran (\labels[0][165] , \labels[0].label[156] );
tran (\labels[0][166] , \labels[0].label[157] );
tran (\labels[0][167] , \labels[0].label[158] );
tran (\labels[0][168] , \labels[0].label[159] );
tran (\labels[0][169] , \labels[0].label[160] );
tran (\labels[0][170] , \labels[0].label[161] );
tran (\labels[0][171] , \labels[0].label[162] );
tran (\labels[0][172] , \labels[0].label[163] );
tran (\labels[0][173] , \labels[0].label[164] );
tran (\labels[0][174] , \labels[0].label[165] );
tran (\labels[0][175] , \labels[0].label[166] );
tran (\labels[0][176] , \labels[0].label[167] );
tran (\labels[0][177] , \labels[0].label[168] );
tran (\labels[0][178] , \labels[0].label[169] );
tran (\labels[0][179] , \labels[0].label[170] );
tran (\labels[0][180] , \labels[0].label[171] );
tran (\labels[0][181] , \labels[0].label[172] );
tran (\labels[0][182] , \labels[0].label[173] );
tran (\labels[0][183] , \labels[0].label[174] );
tran (\labels[0][184] , \labels[0].label[175] );
tran (\labels[0][185] , \labels[0].label[176] );
tran (\labels[0][186] , \labels[0].label[177] );
tran (\labels[0][187] , \labels[0].label[178] );
tran (\labels[0][188] , \labels[0].label[179] );
tran (\labels[0][189] , \labels[0].label[180] );
tran (\labels[0][190] , \labels[0].label[181] );
tran (\labels[0][191] , \labels[0].label[182] );
tran (\labels[0][192] , \labels[0].label[183] );
tran (\labels[0][193] , \labels[0].label[184] );
tran (\labels[0][194] , \labels[0].label[185] );
tran (\labels[0][195] , \labels[0].label[186] );
tran (\labels[0][196] , \labels[0].label[187] );
tran (\labels[0][197] , \labels[0].label[188] );
tran (\labels[0][198] , \labels[0].label[189] );
tran (\labels[0][199] , \labels[0].label[190] );
tran (\labels[0][200] , \labels[0].label[191] );
tran (\labels[0][201] , \labels[0].label[192] );
tran (\labels[0][202] , \labels[0].label[193] );
tran (\labels[0][203] , \labels[0].label[194] );
tran (\labels[0][204] , \labels[0].label[195] );
tran (\labels[0][205] , \labels[0].label[196] );
tran (\labels[0][206] , \labels[0].label[197] );
tran (\labels[0][207] , \labels[0].label[198] );
tran (\labels[0][208] , \labels[0].label[199] );
tran (\labels[0][209] , \labels[0].label[200] );
tran (\labels[0][210] , \labels[0].label[201] );
tran (\labels[0][211] , \labels[0].label[202] );
tran (\labels[0][212] , \labels[0].label[203] );
tran (\labels[0][213] , \labels[0].label[204] );
tran (\labels[0][214] , \labels[0].label[205] );
tran (\labels[0][215] , \labels[0].label[206] );
tran (\labels[0][216] , \labels[0].label[207] );
tran (\labels[0][217] , \labels[0].label[208] );
tran (\labels[0][218] , \labels[0].label[209] );
tran (\labels[0][219] , \labels[0].label[210] );
tran (\labels[0][220] , \labels[0].label[211] );
tran (\labels[0][221] , \labels[0].label[212] );
tran (\labels[0][222] , \labels[0].label[213] );
tran (\labels[0][223] , \labels[0].label[214] );
tran (\labels[0][224] , \labels[0].label[215] );
tran (\labels[0][225] , \labels[0].label[216] );
tran (\labels[0][226] , \labels[0].label[217] );
tran (\labels[0][227] , \labels[0].label[218] );
tran (\labels[0][228] , \labels[0].label[219] );
tran (\labels[0][229] , \labels[0].label[220] );
tran (\labels[0][230] , \labels[0].label[221] );
tran (\labels[0][231] , \labels[0].label[222] );
tran (\labels[0][232] , \labels[0].label[223] );
tran (\labels[0][233] , \labels[0].label[224] );
tran (\labels[0][234] , \labels[0].label[225] );
tran (\labels[0][235] , \labels[0].label[226] );
tran (\labels[0][236] , \labels[0].label[227] );
tran (\labels[0][237] , \labels[0].label[228] );
tran (\labels[0][238] , \labels[0].label[229] );
tran (\labels[0][239] , \labels[0].label[230] );
tran (\labels[0][240] , \labels[0].label[231] );
tran (\labels[0][241] , \labels[0].label[232] );
tran (\labels[0][242] , \labels[0].label[233] );
tran (\labels[0][243] , \labels[0].label[234] );
tran (\labels[0][244] , \labels[0].label[235] );
tran (\labels[0][245] , \labels[0].label[236] );
tran (\labels[0][246] , \labels[0].label[237] );
tran (\labels[0][247] , \labels[0].label[238] );
tran (\labels[0][248] , \labels[0].label[239] );
tran (\labels[0][249] , \labels[0].label[240] );
tran (\labels[0][250] , \labels[0].label[241] );
tran (\labels[0][251] , \labels[0].label[242] );
tran (\labels[0][252] , \labels[0].label[243] );
tran (\labels[0][253] , \labels[0].label[244] );
tran (\labels[0][254] , \labels[0].label[245] );
tran (\labels[0][255] , \labels[0].label[246] );
tran (\labels[0][256] , \labels[0].label[247] );
tran (\labels[0][257] , \labels[0].label[248] );
tran (\labels[0][258] , \labels[0].label[249] );
tran (\labels[0][259] , \labels[0].label[250] );
tran (\labels[0][260] , \labels[0].label[251] );
tran (\labels[0][261] , \labels[0].label[252] );
tran (\labels[0][262] , \labels[0].label[253] );
tran (\labels[0][263] , \labels[0].label[254] );
tran (\labels[0][264] , \labels[0].label[255] );
tran (\labels[0][265] , \labels[0].label_size[0] );
tran (\labels[0][266] , \labels[0].label_size[1] );
tran (\labels[0][267] , \labels[0].label_size[2] );
tran (\labels[0][268] , \labels[0].label_size[3] );
tran (\labels[0][269] , \labels[0].label_size[4] );
tran (\labels[0][270] , \labels[0].label_size[5] );
tran (\labels[0][271] , \labels[0].guid_size[0] );
tran (\labels[1][0] , \labels[1].delimiter[0] );
tran (\labels[1][1] , \labels[1].delimiter[1] );
tran (\labels[1][2] , \labels[1].delimiter[2] );
tran (\labels[1][3] , \labels[1].delimiter[3] );
tran (\labels[1][4] , \labels[1].delimiter[4] );
tran (\labels[1][5] , \labels[1].delimiter[5] );
tran (\labels[1][6] , \labels[1].delimiter[6] );
tran (\labels[1][7] , \labels[1].delimiter[7] );
tran (\labels[1][8] , \labels[1].delimiter_valid[0] );
tran (\labels[1][9] , \labels[1].label[0] );
tran (\labels[1][10] , \labels[1].label[1] );
tran (\labels[1][11] , \labels[1].label[2] );
tran (\labels[1][12] , \labels[1].label[3] );
tran (\labels[1][13] , \labels[1].label[4] );
tran (\labels[1][14] , \labels[1].label[5] );
tran (\labels[1][15] , \labels[1].label[6] );
tran (\labels[1][16] , \labels[1].label[7] );
tran (\labels[1][17] , \labels[1].label[8] );
tran (\labels[1][18] , \labels[1].label[9] );
tran (\labels[1][19] , \labels[1].label[10] );
tran (\labels[1][20] , \labels[1].label[11] );
tran (\labels[1][21] , \labels[1].label[12] );
tran (\labels[1][22] , \labels[1].label[13] );
tran (\labels[1][23] , \labels[1].label[14] );
tran (\labels[1][24] , \labels[1].label[15] );
tran (\labels[1][25] , \labels[1].label[16] );
tran (\labels[1][26] , \labels[1].label[17] );
tran (\labels[1][27] , \labels[1].label[18] );
tran (\labels[1][28] , \labels[1].label[19] );
tran (\labels[1][29] , \labels[1].label[20] );
tran (\labels[1][30] , \labels[1].label[21] );
tran (\labels[1][31] , \labels[1].label[22] );
tran (\labels[1][32] , \labels[1].label[23] );
tran (\labels[1][33] , \labels[1].label[24] );
tran (\labels[1][34] , \labels[1].label[25] );
tran (\labels[1][35] , \labels[1].label[26] );
tran (\labels[1][36] , \labels[1].label[27] );
tran (\labels[1][37] , \labels[1].label[28] );
tran (\labels[1][38] , \labels[1].label[29] );
tran (\labels[1][39] , \labels[1].label[30] );
tran (\labels[1][40] , \labels[1].label[31] );
tran (\labels[1][41] , \labels[1].label[32] );
tran (\labels[1][42] , \labels[1].label[33] );
tran (\labels[1][43] , \labels[1].label[34] );
tran (\labels[1][44] , \labels[1].label[35] );
tran (\labels[1][45] , \labels[1].label[36] );
tran (\labels[1][46] , \labels[1].label[37] );
tran (\labels[1][47] , \labels[1].label[38] );
tran (\labels[1][48] , \labels[1].label[39] );
tran (\labels[1][49] , \labels[1].label[40] );
tran (\labels[1][50] , \labels[1].label[41] );
tran (\labels[1][51] , \labels[1].label[42] );
tran (\labels[1][52] , \labels[1].label[43] );
tran (\labels[1][53] , \labels[1].label[44] );
tran (\labels[1][54] , \labels[1].label[45] );
tran (\labels[1][55] , \labels[1].label[46] );
tran (\labels[1][56] , \labels[1].label[47] );
tran (\labels[1][57] , \labels[1].label[48] );
tran (\labels[1][58] , \labels[1].label[49] );
tran (\labels[1][59] , \labels[1].label[50] );
tran (\labels[1][60] , \labels[1].label[51] );
tran (\labels[1][61] , \labels[1].label[52] );
tran (\labels[1][62] , \labels[1].label[53] );
tran (\labels[1][63] , \labels[1].label[54] );
tran (\labels[1][64] , \labels[1].label[55] );
tran (\labels[1][65] , \labels[1].label[56] );
tran (\labels[1][66] , \labels[1].label[57] );
tran (\labels[1][67] , \labels[1].label[58] );
tran (\labels[1][68] , \labels[1].label[59] );
tran (\labels[1][69] , \labels[1].label[60] );
tran (\labels[1][70] , \labels[1].label[61] );
tran (\labels[1][71] , \labels[1].label[62] );
tran (\labels[1][72] , \labels[1].label[63] );
tran (\labels[1][73] , \labels[1].label[64] );
tran (\labels[1][74] , \labels[1].label[65] );
tran (\labels[1][75] , \labels[1].label[66] );
tran (\labels[1][76] , \labels[1].label[67] );
tran (\labels[1][77] , \labels[1].label[68] );
tran (\labels[1][78] , \labels[1].label[69] );
tran (\labels[1][79] , \labels[1].label[70] );
tran (\labels[1][80] , \labels[1].label[71] );
tran (\labels[1][81] , \labels[1].label[72] );
tran (\labels[1][82] , \labels[1].label[73] );
tran (\labels[1][83] , \labels[1].label[74] );
tran (\labels[1][84] , \labels[1].label[75] );
tran (\labels[1][85] , \labels[1].label[76] );
tran (\labels[1][86] , \labels[1].label[77] );
tran (\labels[1][87] , \labels[1].label[78] );
tran (\labels[1][88] , \labels[1].label[79] );
tran (\labels[1][89] , \labels[1].label[80] );
tran (\labels[1][90] , \labels[1].label[81] );
tran (\labels[1][91] , \labels[1].label[82] );
tran (\labels[1][92] , \labels[1].label[83] );
tran (\labels[1][93] , \labels[1].label[84] );
tran (\labels[1][94] , \labels[1].label[85] );
tran (\labels[1][95] , \labels[1].label[86] );
tran (\labels[1][96] , \labels[1].label[87] );
tran (\labels[1][97] , \labels[1].label[88] );
tran (\labels[1][98] , \labels[1].label[89] );
tran (\labels[1][99] , \labels[1].label[90] );
tran (\labels[1][100] , \labels[1].label[91] );
tran (\labels[1][101] , \labels[1].label[92] );
tran (\labels[1][102] , \labels[1].label[93] );
tran (\labels[1][103] , \labels[1].label[94] );
tran (\labels[1][104] , \labels[1].label[95] );
tran (\labels[1][105] , \labels[1].label[96] );
tran (\labels[1][106] , \labels[1].label[97] );
tran (\labels[1][107] , \labels[1].label[98] );
tran (\labels[1][108] , \labels[1].label[99] );
tran (\labels[1][109] , \labels[1].label[100] );
tran (\labels[1][110] , \labels[1].label[101] );
tran (\labels[1][111] , \labels[1].label[102] );
tran (\labels[1][112] , \labels[1].label[103] );
tran (\labels[1][113] , \labels[1].label[104] );
tran (\labels[1][114] , \labels[1].label[105] );
tran (\labels[1][115] , \labels[1].label[106] );
tran (\labels[1][116] , \labels[1].label[107] );
tran (\labels[1][117] , \labels[1].label[108] );
tran (\labels[1][118] , \labels[1].label[109] );
tran (\labels[1][119] , \labels[1].label[110] );
tran (\labels[1][120] , \labels[1].label[111] );
tran (\labels[1][121] , \labels[1].label[112] );
tran (\labels[1][122] , \labels[1].label[113] );
tran (\labels[1][123] , \labels[1].label[114] );
tran (\labels[1][124] , \labels[1].label[115] );
tran (\labels[1][125] , \labels[1].label[116] );
tran (\labels[1][126] , \labels[1].label[117] );
tran (\labels[1][127] , \labels[1].label[118] );
tran (\labels[1][128] , \labels[1].label[119] );
tran (\labels[1][129] , \labels[1].label[120] );
tran (\labels[1][130] , \labels[1].label[121] );
tran (\labels[1][131] , \labels[1].label[122] );
tran (\labels[1][132] , \labels[1].label[123] );
tran (\labels[1][133] , \labels[1].label[124] );
tran (\labels[1][134] , \labels[1].label[125] );
tran (\labels[1][135] , \labels[1].label[126] );
tran (\labels[1][136] , \labels[1].label[127] );
tran (\labels[1][137] , \labels[1].label[128] );
tran (\labels[1][138] , \labels[1].label[129] );
tran (\labels[1][139] , \labels[1].label[130] );
tran (\labels[1][140] , \labels[1].label[131] );
tran (\labels[1][141] , \labels[1].label[132] );
tran (\labels[1][142] , \labels[1].label[133] );
tran (\labels[1][143] , \labels[1].label[134] );
tran (\labels[1][144] , \labels[1].label[135] );
tran (\labels[1][145] , \labels[1].label[136] );
tran (\labels[1][146] , \labels[1].label[137] );
tran (\labels[1][147] , \labels[1].label[138] );
tran (\labels[1][148] , \labels[1].label[139] );
tran (\labels[1][149] , \labels[1].label[140] );
tran (\labels[1][150] , \labels[1].label[141] );
tran (\labels[1][151] , \labels[1].label[142] );
tran (\labels[1][152] , \labels[1].label[143] );
tran (\labels[1][153] , \labels[1].label[144] );
tran (\labels[1][154] , \labels[1].label[145] );
tran (\labels[1][155] , \labels[1].label[146] );
tran (\labels[1][156] , \labels[1].label[147] );
tran (\labels[1][157] , \labels[1].label[148] );
tran (\labels[1][158] , \labels[1].label[149] );
tran (\labels[1][159] , \labels[1].label[150] );
tran (\labels[1][160] , \labels[1].label[151] );
tran (\labels[1][161] , \labels[1].label[152] );
tran (\labels[1][162] , \labels[1].label[153] );
tran (\labels[1][163] , \labels[1].label[154] );
tran (\labels[1][164] , \labels[1].label[155] );
tran (\labels[1][165] , \labels[1].label[156] );
tran (\labels[1][166] , \labels[1].label[157] );
tran (\labels[1][167] , \labels[1].label[158] );
tran (\labels[1][168] , \labels[1].label[159] );
tran (\labels[1][169] , \labels[1].label[160] );
tran (\labels[1][170] , \labels[1].label[161] );
tran (\labels[1][171] , \labels[1].label[162] );
tran (\labels[1][172] , \labels[1].label[163] );
tran (\labels[1][173] , \labels[1].label[164] );
tran (\labels[1][174] , \labels[1].label[165] );
tran (\labels[1][175] , \labels[1].label[166] );
tran (\labels[1][176] , \labels[1].label[167] );
tran (\labels[1][177] , \labels[1].label[168] );
tran (\labels[1][178] , \labels[1].label[169] );
tran (\labels[1][179] , \labels[1].label[170] );
tran (\labels[1][180] , \labels[1].label[171] );
tran (\labels[1][181] , \labels[1].label[172] );
tran (\labels[1][182] , \labels[1].label[173] );
tran (\labels[1][183] , \labels[1].label[174] );
tran (\labels[1][184] , \labels[1].label[175] );
tran (\labels[1][185] , \labels[1].label[176] );
tran (\labels[1][186] , \labels[1].label[177] );
tran (\labels[1][187] , \labels[1].label[178] );
tran (\labels[1][188] , \labels[1].label[179] );
tran (\labels[1][189] , \labels[1].label[180] );
tran (\labels[1][190] , \labels[1].label[181] );
tran (\labels[1][191] , \labels[1].label[182] );
tran (\labels[1][192] , \labels[1].label[183] );
tran (\labels[1][193] , \labels[1].label[184] );
tran (\labels[1][194] , \labels[1].label[185] );
tran (\labels[1][195] , \labels[1].label[186] );
tran (\labels[1][196] , \labels[1].label[187] );
tran (\labels[1][197] , \labels[1].label[188] );
tran (\labels[1][198] , \labels[1].label[189] );
tran (\labels[1][199] , \labels[1].label[190] );
tran (\labels[1][200] , \labels[1].label[191] );
tran (\labels[1][201] , \labels[1].label[192] );
tran (\labels[1][202] , \labels[1].label[193] );
tran (\labels[1][203] , \labels[1].label[194] );
tran (\labels[1][204] , \labels[1].label[195] );
tran (\labels[1][205] , \labels[1].label[196] );
tran (\labels[1][206] , \labels[1].label[197] );
tran (\labels[1][207] , \labels[1].label[198] );
tran (\labels[1][208] , \labels[1].label[199] );
tran (\labels[1][209] , \labels[1].label[200] );
tran (\labels[1][210] , \labels[1].label[201] );
tran (\labels[1][211] , \labels[1].label[202] );
tran (\labels[1][212] , \labels[1].label[203] );
tran (\labels[1][213] , \labels[1].label[204] );
tran (\labels[1][214] , \labels[1].label[205] );
tran (\labels[1][215] , \labels[1].label[206] );
tran (\labels[1][216] , \labels[1].label[207] );
tran (\labels[1][217] , \labels[1].label[208] );
tran (\labels[1][218] , \labels[1].label[209] );
tran (\labels[1][219] , \labels[1].label[210] );
tran (\labels[1][220] , \labels[1].label[211] );
tran (\labels[1][221] , \labels[1].label[212] );
tran (\labels[1][222] , \labels[1].label[213] );
tran (\labels[1][223] , \labels[1].label[214] );
tran (\labels[1][224] , \labels[1].label[215] );
tran (\labels[1][225] , \labels[1].label[216] );
tran (\labels[1][226] , \labels[1].label[217] );
tran (\labels[1][227] , \labels[1].label[218] );
tran (\labels[1][228] , \labels[1].label[219] );
tran (\labels[1][229] , \labels[1].label[220] );
tran (\labels[1][230] , \labels[1].label[221] );
tran (\labels[1][231] , \labels[1].label[222] );
tran (\labels[1][232] , \labels[1].label[223] );
tran (\labels[1][233] , \labels[1].label[224] );
tran (\labels[1][234] , \labels[1].label[225] );
tran (\labels[1][235] , \labels[1].label[226] );
tran (\labels[1][236] , \labels[1].label[227] );
tran (\labels[1][237] , \labels[1].label[228] );
tran (\labels[1][238] , \labels[1].label[229] );
tran (\labels[1][239] , \labels[1].label[230] );
tran (\labels[1][240] , \labels[1].label[231] );
tran (\labels[1][241] , \labels[1].label[232] );
tran (\labels[1][242] , \labels[1].label[233] );
tran (\labels[1][243] , \labels[1].label[234] );
tran (\labels[1][244] , \labels[1].label[235] );
tran (\labels[1][245] , \labels[1].label[236] );
tran (\labels[1][246] , \labels[1].label[237] );
tran (\labels[1][247] , \labels[1].label[238] );
tran (\labels[1][248] , \labels[1].label[239] );
tran (\labels[1][249] , \labels[1].label[240] );
tran (\labels[1][250] , \labels[1].label[241] );
tran (\labels[1][251] , \labels[1].label[242] );
tran (\labels[1][252] , \labels[1].label[243] );
tran (\labels[1][253] , \labels[1].label[244] );
tran (\labels[1][254] , \labels[1].label[245] );
tran (\labels[1][255] , \labels[1].label[246] );
tran (\labels[1][256] , \labels[1].label[247] );
tran (\labels[1][257] , \labels[1].label[248] );
tran (\labels[1][258] , \labels[1].label[249] );
tran (\labels[1][259] , \labels[1].label[250] );
tran (\labels[1][260] , \labels[1].label[251] );
tran (\labels[1][261] , \labels[1].label[252] );
tran (\labels[1][262] , \labels[1].label[253] );
tran (\labels[1][263] , \labels[1].label[254] );
tran (\labels[1][264] , \labels[1].label[255] );
tran (\labels[1][265] , \labels[1].label_size[0] );
tran (\labels[1][266] , \labels[1].label_size[1] );
tran (\labels[1][267] , \labels[1].label_size[2] );
tran (\labels[1][268] , \labels[1].label_size[3] );
tran (\labels[1][269] , \labels[1].label_size[4] );
tran (\labels[1][270] , \labels[1].label_size[5] );
tran (\labels[1][271] , \labels[1].guid_size[0] );
tran (\labels[2][0] , \labels[2].delimiter[0] );
tran (\labels[2][1] , \labels[2].delimiter[1] );
tran (\labels[2][2] , \labels[2].delimiter[2] );
tran (\labels[2][3] , \labels[2].delimiter[3] );
tran (\labels[2][4] , \labels[2].delimiter[4] );
tran (\labels[2][5] , \labels[2].delimiter[5] );
tran (\labels[2][6] , \labels[2].delimiter[6] );
tran (\labels[2][7] , \labels[2].delimiter[7] );
tran (\labels[2][8] , \labels[2].delimiter_valid[0] );
tran (\labels[2][9] , \labels[2].label[0] );
tran (\labels[2][10] , \labels[2].label[1] );
tran (\labels[2][11] , \labels[2].label[2] );
tran (\labels[2][12] , \labels[2].label[3] );
tran (\labels[2][13] , \labels[2].label[4] );
tran (\labels[2][14] , \labels[2].label[5] );
tran (\labels[2][15] , \labels[2].label[6] );
tran (\labels[2][16] , \labels[2].label[7] );
tran (\labels[2][17] , \labels[2].label[8] );
tran (\labels[2][18] , \labels[2].label[9] );
tran (\labels[2][19] , \labels[2].label[10] );
tran (\labels[2][20] , \labels[2].label[11] );
tran (\labels[2][21] , \labels[2].label[12] );
tran (\labels[2][22] , \labels[2].label[13] );
tran (\labels[2][23] , \labels[2].label[14] );
tran (\labels[2][24] , \labels[2].label[15] );
tran (\labels[2][25] , \labels[2].label[16] );
tran (\labels[2][26] , \labels[2].label[17] );
tran (\labels[2][27] , \labels[2].label[18] );
tran (\labels[2][28] , \labels[2].label[19] );
tran (\labels[2][29] , \labels[2].label[20] );
tran (\labels[2][30] , \labels[2].label[21] );
tran (\labels[2][31] , \labels[2].label[22] );
tran (\labels[2][32] , \labels[2].label[23] );
tran (\labels[2][33] , \labels[2].label[24] );
tran (\labels[2][34] , \labels[2].label[25] );
tran (\labels[2][35] , \labels[2].label[26] );
tran (\labels[2][36] , \labels[2].label[27] );
tran (\labels[2][37] , \labels[2].label[28] );
tran (\labels[2][38] , \labels[2].label[29] );
tran (\labels[2][39] , \labels[2].label[30] );
tran (\labels[2][40] , \labels[2].label[31] );
tran (\labels[2][41] , \labels[2].label[32] );
tran (\labels[2][42] , \labels[2].label[33] );
tran (\labels[2][43] , \labels[2].label[34] );
tran (\labels[2][44] , \labels[2].label[35] );
tran (\labels[2][45] , \labels[2].label[36] );
tran (\labels[2][46] , \labels[2].label[37] );
tran (\labels[2][47] , \labels[2].label[38] );
tran (\labels[2][48] , \labels[2].label[39] );
tran (\labels[2][49] , \labels[2].label[40] );
tran (\labels[2][50] , \labels[2].label[41] );
tran (\labels[2][51] , \labels[2].label[42] );
tran (\labels[2][52] , \labels[2].label[43] );
tran (\labels[2][53] , \labels[2].label[44] );
tran (\labels[2][54] , \labels[2].label[45] );
tran (\labels[2][55] , \labels[2].label[46] );
tran (\labels[2][56] , \labels[2].label[47] );
tran (\labels[2][57] , \labels[2].label[48] );
tran (\labels[2][58] , \labels[2].label[49] );
tran (\labels[2][59] , \labels[2].label[50] );
tran (\labels[2][60] , \labels[2].label[51] );
tran (\labels[2][61] , \labels[2].label[52] );
tran (\labels[2][62] , \labels[2].label[53] );
tran (\labels[2][63] , \labels[2].label[54] );
tran (\labels[2][64] , \labels[2].label[55] );
tran (\labels[2][65] , \labels[2].label[56] );
tran (\labels[2][66] , \labels[2].label[57] );
tran (\labels[2][67] , \labels[2].label[58] );
tran (\labels[2][68] , \labels[2].label[59] );
tran (\labels[2][69] , \labels[2].label[60] );
tran (\labels[2][70] , \labels[2].label[61] );
tran (\labels[2][71] , \labels[2].label[62] );
tran (\labels[2][72] , \labels[2].label[63] );
tran (\labels[2][73] , \labels[2].label[64] );
tran (\labels[2][74] , \labels[2].label[65] );
tran (\labels[2][75] , \labels[2].label[66] );
tran (\labels[2][76] , \labels[2].label[67] );
tran (\labels[2][77] , \labels[2].label[68] );
tran (\labels[2][78] , \labels[2].label[69] );
tran (\labels[2][79] , \labels[2].label[70] );
tran (\labels[2][80] , \labels[2].label[71] );
tran (\labels[2][81] , \labels[2].label[72] );
tran (\labels[2][82] , \labels[2].label[73] );
tran (\labels[2][83] , \labels[2].label[74] );
tran (\labels[2][84] , \labels[2].label[75] );
tran (\labels[2][85] , \labels[2].label[76] );
tran (\labels[2][86] , \labels[2].label[77] );
tran (\labels[2][87] , \labels[2].label[78] );
tran (\labels[2][88] , \labels[2].label[79] );
tran (\labels[2][89] , \labels[2].label[80] );
tran (\labels[2][90] , \labels[2].label[81] );
tran (\labels[2][91] , \labels[2].label[82] );
tran (\labels[2][92] , \labels[2].label[83] );
tran (\labels[2][93] , \labels[2].label[84] );
tran (\labels[2][94] , \labels[2].label[85] );
tran (\labels[2][95] , \labels[2].label[86] );
tran (\labels[2][96] , \labels[2].label[87] );
tran (\labels[2][97] , \labels[2].label[88] );
tran (\labels[2][98] , \labels[2].label[89] );
tran (\labels[2][99] , \labels[2].label[90] );
tran (\labels[2][100] , \labels[2].label[91] );
tran (\labels[2][101] , \labels[2].label[92] );
tran (\labels[2][102] , \labels[2].label[93] );
tran (\labels[2][103] , \labels[2].label[94] );
tran (\labels[2][104] , \labels[2].label[95] );
tran (\labels[2][105] , \labels[2].label[96] );
tran (\labels[2][106] , \labels[2].label[97] );
tran (\labels[2][107] , \labels[2].label[98] );
tran (\labels[2][108] , \labels[2].label[99] );
tran (\labels[2][109] , \labels[2].label[100] );
tran (\labels[2][110] , \labels[2].label[101] );
tran (\labels[2][111] , \labels[2].label[102] );
tran (\labels[2][112] , \labels[2].label[103] );
tran (\labels[2][113] , \labels[2].label[104] );
tran (\labels[2][114] , \labels[2].label[105] );
tran (\labels[2][115] , \labels[2].label[106] );
tran (\labels[2][116] , \labels[2].label[107] );
tran (\labels[2][117] , \labels[2].label[108] );
tran (\labels[2][118] , \labels[2].label[109] );
tran (\labels[2][119] , \labels[2].label[110] );
tran (\labels[2][120] , \labels[2].label[111] );
tran (\labels[2][121] , \labels[2].label[112] );
tran (\labels[2][122] , \labels[2].label[113] );
tran (\labels[2][123] , \labels[2].label[114] );
tran (\labels[2][124] , \labels[2].label[115] );
tran (\labels[2][125] , \labels[2].label[116] );
tran (\labels[2][126] , \labels[2].label[117] );
tran (\labels[2][127] , \labels[2].label[118] );
tran (\labels[2][128] , \labels[2].label[119] );
tran (\labels[2][129] , \labels[2].label[120] );
tran (\labels[2][130] , \labels[2].label[121] );
tran (\labels[2][131] , \labels[2].label[122] );
tran (\labels[2][132] , \labels[2].label[123] );
tran (\labels[2][133] , \labels[2].label[124] );
tran (\labels[2][134] , \labels[2].label[125] );
tran (\labels[2][135] , \labels[2].label[126] );
tran (\labels[2][136] , \labels[2].label[127] );
tran (\labels[2][137] , \labels[2].label[128] );
tran (\labels[2][138] , \labels[2].label[129] );
tran (\labels[2][139] , \labels[2].label[130] );
tran (\labels[2][140] , \labels[2].label[131] );
tran (\labels[2][141] , \labels[2].label[132] );
tran (\labels[2][142] , \labels[2].label[133] );
tran (\labels[2][143] , \labels[2].label[134] );
tran (\labels[2][144] , \labels[2].label[135] );
tran (\labels[2][145] , \labels[2].label[136] );
tran (\labels[2][146] , \labels[2].label[137] );
tran (\labels[2][147] , \labels[2].label[138] );
tran (\labels[2][148] , \labels[2].label[139] );
tran (\labels[2][149] , \labels[2].label[140] );
tran (\labels[2][150] , \labels[2].label[141] );
tran (\labels[2][151] , \labels[2].label[142] );
tran (\labels[2][152] , \labels[2].label[143] );
tran (\labels[2][153] , \labels[2].label[144] );
tran (\labels[2][154] , \labels[2].label[145] );
tran (\labels[2][155] , \labels[2].label[146] );
tran (\labels[2][156] , \labels[2].label[147] );
tran (\labels[2][157] , \labels[2].label[148] );
tran (\labels[2][158] , \labels[2].label[149] );
tran (\labels[2][159] , \labels[2].label[150] );
tran (\labels[2][160] , \labels[2].label[151] );
tran (\labels[2][161] , \labels[2].label[152] );
tran (\labels[2][162] , \labels[2].label[153] );
tran (\labels[2][163] , \labels[2].label[154] );
tran (\labels[2][164] , \labels[2].label[155] );
tran (\labels[2][165] , \labels[2].label[156] );
tran (\labels[2][166] , \labels[2].label[157] );
tran (\labels[2][167] , \labels[2].label[158] );
tran (\labels[2][168] , \labels[2].label[159] );
tran (\labels[2][169] , \labels[2].label[160] );
tran (\labels[2][170] , \labels[2].label[161] );
tran (\labels[2][171] , \labels[2].label[162] );
tran (\labels[2][172] , \labels[2].label[163] );
tran (\labels[2][173] , \labels[2].label[164] );
tran (\labels[2][174] , \labels[2].label[165] );
tran (\labels[2][175] , \labels[2].label[166] );
tran (\labels[2][176] , \labels[2].label[167] );
tran (\labels[2][177] , \labels[2].label[168] );
tran (\labels[2][178] , \labels[2].label[169] );
tran (\labels[2][179] , \labels[2].label[170] );
tran (\labels[2][180] , \labels[2].label[171] );
tran (\labels[2][181] , \labels[2].label[172] );
tran (\labels[2][182] , \labels[2].label[173] );
tran (\labels[2][183] , \labels[2].label[174] );
tran (\labels[2][184] , \labels[2].label[175] );
tran (\labels[2][185] , \labels[2].label[176] );
tran (\labels[2][186] , \labels[2].label[177] );
tran (\labels[2][187] , \labels[2].label[178] );
tran (\labels[2][188] , \labels[2].label[179] );
tran (\labels[2][189] , \labels[2].label[180] );
tran (\labels[2][190] , \labels[2].label[181] );
tran (\labels[2][191] , \labels[2].label[182] );
tran (\labels[2][192] , \labels[2].label[183] );
tran (\labels[2][193] , \labels[2].label[184] );
tran (\labels[2][194] , \labels[2].label[185] );
tran (\labels[2][195] , \labels[2].label[186] );
tran (\labels[2][196] , \labels[2].label[187] );
tran (\labels[2][197] , \labels[2].label[188] );
tran (\labels[2][198] , \labels[2].label[189] );
tran (\labels[2][199] , \labels[2].label[190] );
tran (\labels[2][200] , \labels[2].label[191] );
tran (\labels[2][201] , \labels[2].label[192] );
tran (\labels[2][202] , \labels[2].label[193] );
tran (\labels[2][203] , \labels[2].label[194] );
tran (\labels[2][204] , \labels[2].label[195] );
tran (\labels[2][205] , \labels[2].label[196] );
tran (\labels[2][206] , \labels[2].label[197] );
tran (\labels[2][207] , \labels[2].label[198] );
tran (\labels[2][208] , \labels[2].label[199] );
tran (\labels[2][209] , \labels[2].label[200] );
tran (\labels[2][210] , \labels[2].label[201] );
tran (\labels[2][211] , \labels[2].label[202] );
tran (\labels[2][212] , \labels[2].label[203] );
tran (\labels[2][213] , \labels[2].label[204] );
tran (\labels[2][214] , \labels[2].label[205] );
tran (\labels[2][215] , \labels[2].label[206] );
tran (\labels[2][216] , \labels[2].label[207] );
tran (\labels[2][217] , \labels[2].label[208] );
tran (\labels[2][218] , \labels[2].label[209] );
tran (\labels[2][219] , \labels[2].label[210] );
tran (\labels[2][220] , \labels[2].label[211] );
tran (\labels[2][221] , \labels[2].label[212] );
tran (\labels[2][222] , \labels[2].label[213] );
tran (\labels[2][223] , \labels[2].label[214] );
tran (\labels[2][224] , \labels[2].label[215] );
tran (\labels[2][225] , \labels[2].label[216] );
tran (\labels[2][226] , \labels[2].label[217] );
tran (\labels[2][227] , \labels[2].label[218] );
tran (\labels[2][228] , \labels[2].label[219] );
tran (\labels[2][229] , \labels[2].label[220] );
tran (\labels[2][230] , \labels[2].label[221] );
tran (\labels[2][231] , \labels[2].label[222] );
tran (\labels[2][232] , \labels[2].label[223] );
tran (\labels[2][233] , \labels[2].label[224] );
tran (\labels[2][234] , \labels[2].label[225] );
tran (\labels[2][235] , \labels[2].label[226] );
tran (\labels[2][236] , \labels[2].label[227] );
tran (\labels[2][237] , \labels[2].label[228] );
tran (\labels[2][238] , \labels[2].label[229] );
tran (\labels[2][239] , \labels[2].label[230] );
tran (\labels[2][240] , \labels[2].label[231] );
tran (\labels[2][241] , \labels[2].label[232] );
tran (\labels[2][242] , \labels[2].label[233] );
tran (\labels[2][243] , \labels[2].label[234] );
tran (\labels[2][244] , \labels[2].label[235] );
tran (\labels[2][245] , \labels[2].label[236] );
tran (\labels[2][246] , \labels[2].label[237] );
tran (\labels[2][247] , \labels[2].label[238] );
tran (\labels[2][248] , \labels[2].label[239] );
tran (\labels[2][249] , \labels[2].label[240] );
tran (\labels[2][250] , \labels[2].label[241] );
tran (\labels[2][251] , \labels[2].label[242] );
tran (\labels[2][252] , \labels[2].label[243] );
tran (\labels[2][253] , \labels[2].label[244] );
tran (\labels[2][254] , \labels[2].label[245] );
tran (\labels[2][255] , \labels[2].label[246] );
tran (\labels[2][256] , \labels[2].label[247] );
tran (\labels[2][257] , \labels[2].label[248] );
tran (\labels[2][258] , \labels[2].label[249] );
tran (\labels[2][259] , \labels[2].label[250] );
tran (\labels[2][260] , \labels[2].label[251] );
tran (\labels[2][261] , \labels[2].label[252] );
tran (\labels[2][262] , \labels[2].label[253] );
tran (\labels[2][263] , \labels[2].label[254] );
tran (\labels[2][264] , \labels[2].label[255] );
tran (\labels[2][265] , \labels[2].label_size[0] );
tran (\labels[2][266] , \labels[2].label_size[1] );
tran (\labels[2][267] , \labels[2].label_size[2] );
tran (\labels[2][268] , \labels[2].label_size[3] );
tran (\labels[2][269] , \labels[2].label_size[4] );
tran (\labels[2][270] , \labels[2].label_size[5] );
tran (\labels[2][271] , \labels[2].guid_size[0] );
tran (\labels[3][0] , \labels[3].delimiter[0] );
tran (\labels[3][1] , \labels[3].delimiter[1] );
tran (\labels[3][2] , \labels[3].delimiter[2] );
tran (\labels[3][3] , \labels[3].delimiter[3] );
tran (\labels[3][4] , \labels[3].delimiter[4] );
tran (\labels[3][5] , \labels[3].delimiter[5] );
tran (\labels[3][6] , \labels[3].delimiter[6] );
tran (\labels[3][7] , \labels[3].delimiter[7] );
tran (\labels[3][8] , \labels[3].delimiter_valid[0] );
tran (\labels[3][9] , \labels[3].label[0] );
tran (\labels[3][10] , \labels[3].label[1] );
tran (\labels[3][11] , \labels[3].label[2] );
tran (\labels[3][12] , \labels[3].label[3] );
tran (\labels[3][13] , \labels[3].label[4] );
tran (\labels[3][14] , \labels[3].label[5] );
tran (\labels[3][15] , \labels[3].label[6] );
tran (\labels[3][16] , \labels[3].label[7] );
tran (\labels[3][17] , \labels[3].label[8] );
tran (\labels[3][18] , \labels[3].label[9] );
tran (\labels[3][19] , \labels[3].label[10] );
tran (\labels[3][20] , \labels[3].label[11] );
tran (\labels[3][21] , \labels[3].label[12] );
tran (\labels[3][22] , \labels[3].label[13] );
tran (\labels[3][23] , \labels[3].label[14] );
tran (\labels[3][24] , \labels[3].label[15] );
tran (\labels[3][25] , \labels[3].label[16] );
tran (\labels[3][26] , \labels[3].label[17] );
tran (\labels[3][27] , \labels[3].label[18] );
tran (\labels[3][28] , \labels[3].label[19] );
tran (\labels[3][29] , \labels[3].label[20] );
tran (\labels[3][30] , \labels[3].label[21] );
tran (\labels[3][31] , \labels[3].label[22] );
tran (\labels[3][32] , \labels[3].label[23] );
tran (\labels[3][33] , \labels[3].label[24] );
tran (\labels[3][34] , \labels[3].label[25] );
tran (\labels[3][35] , \labels[3].label[26] );
tran (\labels[3][36] , \labels[3].label[27] );
tran (\labels[3][37] , \labels[3].label[28] );
tran (\labels[3][38] , \labels[3].label[29] );
tran (\labels[3][39] , \labels[3].label[30] );
tran (\labels[3][40] , \labels[3].label[31] );
tran (\labels[3][41] , \labels[3].label[32] );
tran (\labels[3][42] , \labels[3].label[33] );
tran (\labels[3][43] , \labels[3].label[34] );
tran (\labels[3][44] , \labels[3].label[35] );
tran (\labels[3][45] , \labels[3].label[36] );
tran (\labels[3][46] , \labels[3].label[37] );
tran (\labels[3][47] , \labels[3].label[38] );
tran (\labels[3][48] , \labels[3].label[39] );
tran (\labels[3][49] , \labels[3].label[40] );
tran (\labels[3][50] , \labels[3].label[41] );
tran (\labels[3][51] , \labels[3].label[42] );
tran (\labels[3][52] , \labels[3].label[43] );
tran (\labels[3][53] , \labels[3].label[44] );
tran (\labels[3][54] , \labels[3].label[45] );
tran (\labels[3][55] , \labels[3].label[46] );
tran (\labels[3][56] , \labels[3].label[47] );
tran (\labels[3][57] , \labels[3].label[48] );
tran (\labels[3][58] , \labels[3].label[49] );
tran (\labels[3][59] , \labels[3].label[50] );
tran (\labels[3][60] , \labels[3].label[51] );
tran (\labels[3][61] , \labels[3].label[52] );
tran (\labels[3][62] , \labels[3].label[53] );
tran (\labels[3][63] , \labels[3].label[54] );
tran (\labels[3][64] , \labels[3].label[55] );
tran (\labels[3][65] , \labels[3].label[56] );
tran (\labels[3][66] , \labels[3].label[57] );
tran (\labels[3][67] , \labels[3].label[58] );
tran (\labels[3][68] , \labels[3].label[59] );
tran (\labels[3][69] , \labels[3].label[60] );
tran (\labels[3][70] , \labels[3].label[61] );
tran (\labels[3][71] , \labels[3].label[62] );
tran (\labels[3][72] , \labels[3].label[63] );
tran (\labels[3][73] , \labels[3].label[64] );
tran (\labels[3][74] , \labels[3].label[65] );
tran (\labels[3][75] , \labels[3].label[66] );
tran (\labels[3][76] , \labels[3].label[67] );
tran (\labels[3][77] , \labels[3].label[68] );
tran (\labels[3][78] , \labels[3].label[69] );
tran (\labels[3][79] , \labels[3].label[70] );
tran (\labels[3][80] , \labels[3].label[71] );
tran (\labels[3][81] , \labels[3].label[72] );
tran (\labels[3][82] , \labels[3].label[73] );
tran (\labels[3][83] , \labels[3].label[74] );
tran (\labels[3][84] , \labels[3].label[75] );
tran (\labels[3][85] , \labels[3].label[76] );
tran (\labels[3][86] , \labels[3].label[77] );
tran (\labels[3][87] , \labels[3].label[78] );
tran (\labels[3][88] , \labels[3].label[79] );
tran (\labels[3][89] , \labels[3].label[80] );
tran (\labels[3][90] , \labels[3].label[81] );
tran (\labels[3][91] , \labels[3].label[82] );
tran (\labels[3][92] , \labels[3].label[83] );
tran (\labels[3][93] , \labels[3].label[84] );
tran (\labels[3][94] , \labels[3].label[85] );
tran (\labels[3][95] , \labels[3].label[86] );
tran (\labels[3][96] , \labels[3].label[87] );
tran (\labels[3][97] , \labels[3].label[88] );
tran (\labels[3][98] , \labels[3].label[89] );
tran (\labels[3][99] , \labels[3].label[90] );
tran (\labels[3][100] , \labels[3].label[91] );
tran (\labels[3][101] , \labels[3].label[92] );
tran (\labels[3][102] , \labels[3].label[93] );
tran (\labels[3][103] , \labels[3].label[94] );
tran (\labels[3][104] , \labels[3].label[95] );
tran (\labels[3][105] , \labels[3].label[96] );
tran (\labels[3][106] , \labels[3].label[97] );
tran (\labels[3][107] , \labels[3].label[98] );
tran (\labels[3][108] , \labels[3].label[99] );
tran (\labels[3][109] , \labels[3].label[100] );
tran (\labels[3][110] , \labels[3].label[101] );
tran (\labels[3][111] , \labels[3].label[102] );
tran (\labels[3][112] , \labels[3].label[103] );
tran (\labels[3][113] , \labels[3].label[104] );
tran (\labels[3][114] , \labels[3].label[105] );
tran (\labels[3][115] , \labels[3].label[106] );
tran (\labels[3][116] , \labels[3].label[107] );
tran (\labels[3][117] , \labels[3].label[108] );
tran (\labels[3][118] , \labels[3].label[109] );
tran (\labels[3][119] , \labels[3].label[110] );
tran (\labels[3][120] , \labels[3].label[111] );
tran (\labels[3][121] , \labels[3].label[112] );
tran (\labels[3][122] , \labels[3].label[113] );
tran (\labels[3][123] , \labels[3].label[114] );
tran (\labels[3][124] , \labels[3].label[115] );
tran (\labels[3][125] , \labels[3].label[116] );
tran (\labels[3][126] , \labels[3].label[117] );
tran (\labels[3][127] , \labels[3].label[118] );
tran (\labels[3][128] , \labels[3].label[119] );
tran (\labels[3][129] , \labels[3].label[120] );
tran (\labels[3][130] , \labels[3].label[121] );
tran (\labels[3][131] , \labels[3].label[122] );
tran (\labels[3][132] , \labels[3].label[123] );
tran (\labels[3][133] , \labels[3].label[124] );
tran (\labels[3][134] , \labels[3].label[125] );
tran (\labels[3][135] , \labels[3].label[126] );
tran (\labels[3][136] , \labels[3].label[127] );
tran (\labels[3][137] , \labels[3].label[128] );
tran (\labels[3][138] , \labels[3].label[129] );
tran (\labels[3][139] , \labels[3].label[130] );
tran (\labels[3][140] , \labels[3].label[131] );
tran (\labels[3][141] , \labels[3].label[132] );
tran (\labels[3][142] , \labels[3].label[133] );
tran (\labels[3][143] , \labels[3].label[134] );
tran (\labels[3][144] , \labels[3].label[135] );
tran (\labels[3][145] , \labels[3].label[136] );
tran (\labels[3][146] , \labels[3].label[137] );
tran (\labels[3][147] , \labels[3].label[138] );
tran (\labels[3][148] , \labels[3].label[139] );
tran (\labels[3][149] , \labels[3].label[140] );
tran (\labels[3][150] , \labels[3].label[141] );
tran (\labels[3][151] , \labels[3].label[142] );
tran (\labels[3][152] , \labels[3].label[143] );
tran (\labels[3][153] , \labels[3].label[144] );
tran (\labels[3][154] , \labels[3].label[145] );
tran (\labels[3][155] , \labels[3].label[146] );
tran (\labels[3][156] , \labels[3].label[147] );
tran (\labels[3][157] , \labels[3].label[148] );
tran (\labels[3][158] , \labels[3].label[149] );
tran (\labels[3][159] , \labels[3].label[150] );
tran (\labels[3][160] , \labels[3].label[151] );
tran (\labels[3][161] , \labels[3].label[152] );
tran (\labels[3][162] , \labels[3].label[153] );
tran (\labels[3][163] , \labels[3].label[154] );
tran (\labels[3][164] , \labels[3].label[155] );
tran (\labels[3][165] , \labels[3].label[156] );
tran (\labels[3][166] , \labels[3].label[157] );
tran (\labels[3][167] , \labels[3].label[158] );
tran (\labels[3][168] , \labels[3].label[159] );
tran (\labels[3][169] , \labels[3].label[160] );
tran (\labels[3][170] , \labels[3].label[161] );
tran (\labels[3][171] , \labels[3].label[162] );
tran (\labels[3][172] , \labels[3].label[163] );
tran (\labels[3][173] , \labels[3].label[164] );
tran (\labels[3][174] , \labels[3].label[165] );
tran (\labels[3][175] , \labels[3].label[166] );
tran (\labels[3][176] , \labels[3].label[167] );
tran (\labels[3][177] , \labels[3].label[168] );
tran (\labels[3][178] , \labels[3].label[169] );
tran (\labels[3][179] , \labels[3].label[170] );
tran (\labels[3][180] , \labels[3].label[171] );
tran (\labels[3][181] , \labels[3].label[172] );
tran (\labels[3][182] , \labels[3].label[173] );
tran (\labels[3][183] , \labels[3].label[174] );
tran (\labels[3][184] , \labels[3].label[175] );
tran (\labels[3][185] , \labels[3].label[176] );
tran (\labels[3][186] , \labels[3].label[177] );
tran (\labels[3][187] , \labels[3].label[178] );
tran (\labels[3][188] , \labels[3].label[179] );
tran (\labels[3][189] , \labels[3].label[180] );
tran (\labels[3][190] , \labels[3].label[181] );
tran (\labels[3][191] , \labels[3].label[182] );
tran (\labels[3][192] , \labels[3].label[183] );
tran (\labels[3][193] , \labels[3].label[184] );
tran (\labels[3][194] , \labels[3].label[185] );
tran (\labels[3][195] , \labels[3].label[186] );
tran (\labels[3][196] , \labels[3].label[187] );
tran (\labels[3][197] , \labels[3].label[188] );
tran (\labels[3][198] , \labels[3].label[189] );
tran (\labels[3][199] , \labels[3].label[190] );
tran (\labels[3][200] , \labels[3].label[191] );
tran (\labels[3][201] , \labels[3].label[192] );
tran (\labels[3][202] , \labels[3].label[193] );
tran (\labels[3][203] , \labels[3].label[194] );
tran (\labels[3][204] , \labels[3].label[195] );
tran (\labels[3][205] , \labels[3].label[196] );
tran (\labels[3][206] , \labels[3].label[197] );
tran (\labels[3][207] , \labels[3].label[198] );
tran (\labels[3][208] , \labels[3].label[199] );
tran (\labels[3][209] , \labels[3].label[200] );
tran (\labels[3][210] , \labels[3].label[201] );
tran (\labels[3][211] , \labels[3].label[202] );
tran (\labels[3][212] , \labels[3].label[203] );
tran (\labels[3][213] , \labels[3].label[204] );
tran (\labels[3][214] , \labels[3].label[205] );
tran (\labels[3][215] , \labels[3].label[206] );
tran (\labels[3][216] , \labels[3].label[207] );
tran (\labels[3][217] , \labels[3].label[208] );
tran (\labels[3][218] , \labels[3].label[209] );
tran (\labels[3][219] , \labels[3].label[210] );
tran (\labels[3][220] , \labels[3].label[211] );
tran (\labels[3][221] , \labels[3].label[212] );
tran (\labels[3][222] , \labels[3].label[213] );
tran (\labels[3][223] , \labels[3].label[214] );
tran (\labels[3][224] , \labels[3].label[215] );
tran (\labels[3][225] , \labels[3].label[216] );
tran (\labels[3][226] , \labels[3].label[217] );
tran (\labels[3][227] , \labels[3].label[218] );
tran (\labels[3][228] , \labels[3].label[219] );
tran (\labels[3][229] , \labels[3].label[220] );
tran (\labels[3][230] , \labels[3].label[221] );
tran (\labels[3][231] , \labels[3].label[222] );
tran (\labels[3][232] , \labels[3].label[223] );
tran (\labels[3][233] , \labels[3].label[224] );
tran (\labels[3][234] , \labels[3].label[225] );
tran (\labels[3][235] , \labels[3].label[226] );
tran (\labels[3][236] , \labels[3].label[227] );
tran (\labels[3][237] , \labels[3].label[228] );
tran (\labels[3][238] , \labels[3].label[229] );
tran (\labels[3][239] , \labels[3].label[230] );
tran (\labels[3][240] , \labels[3].label[231] );
tran (\labels[3][241] , \labels[3].label[232] );
tran (\labels[3][242] , \labels[3].label[233] );
tran (\labels[3][243] , \labels[3].label[234] );
tran (\labels[3][244] , \labels[3].label[235] );
tran (\labels[3][245] , \labels[3].label[236] );
tran (\labels[3][246] , \labels[3].label[237] );
tran (\labels[3][247] , \labels[3].label[238] );
tran (\labels[3][248] , \labels[3].label[239] );
tran (\labels[3][249] , \labels[3].label[240] );
tran (\labels[3][250] , \labels[3].label[241] );
tran (\labels[3][251] , \labels[3].label[242] );
tran (\labels[3][252] , \labels[3].label[243] );
tran (\labels[3][253] , \labels[3].label[244] );
tran (\labels[3][254] , \labels[3].label[245] );
tran (\labels[3][255] , \labels[3].label[246] );
tran (\labels[3][256] , \labels[3].label[247] );
tran (\labels[3][257] , \labels[3].label[248] );
tran (\labels[3][258] , \labels[3].label[249] );
tran (\labels[3][259] , \labels[3].label[250] );
tran (\labels[3][260] , \labels[3].label[251] );
tran (\labels[3][261] , \labels[3].label[252] );
tran (\labels[3][262] , \labels[3].label[253] );
tran (\labels[3][263] , \labels[3].label[254] );
tran (\labels[3][264] , \labels[3].label[255] );
tran (\labels[3][265] , \labels[3].label_size[0] );
tran (\labels[3][266] , \labels[3].label_size[1] );
tran (\labels[3][267] , \labels[3].label_size[2] );
tran (\labels[3][268] , \labels[3].label_size[3] );
tran (\labels[3][269] , \labels[3].label_size[4] );
tran (\labels[3][270] , \labels[3].label_size[5] );
tran (\labels[3][271] , \labels[3].guid_size[0] );
tran (\labels[4][0] , \labels[4].delimiter[0] );
tran (\labels[4][1] , \labels[4].delimiter[1] );
tran (\labels[4][2] , \labels[4].delimiter[2] );
tran (\labels[4][3] , \labels[4].delimiter[3] );
tran (\labels[4][4] , \labels[4].delimiter[4] );
tran (\labels[4][5] , \labels[4].delimiter[5] );
tran (\labels[4][6] , \labels[4].delimiter[6] );
tran (\labels[4][7] , \labels[4].delimiter[7] );
tran (\labels[4][8] , \labels[4].delimiter_valid[0] );
tran (\labels[4][9] , \labels[4].label[0] );
tran (\labels[4][10] , \labels[4].label[1] );
tran (\labels[4][11] , \labels[4].label[2] );
tran (\labels[4][12] , \labels[4].label[3] );
tran (\labels[4][13] , \labels[4].label[4] );
tran (\labels[4][14] , \labels[4].label[5] );
tran (\labels[4][15] , \labels[4].label[6] );
tran (\labels[4][16] , \labels[4].label[7] );
tran (\labels[4][17] , \labels[4].label[8] );
tran (\labels[4][18] , \labels[4].label[9] );
tran (\labels[4][19] , \labels[4].label[10] );
tran (\labels[4][20] , \labels[4].label[11] );
tran (\labels[4][21] , \labels[4].label[12] );
tran (\labels[4][22] , \labels[4].label[13] );
tran (\labels[4][23] , \labels[4].label[14] );
tran (\labels[4][24] , \labels[4].label[15] );
tran (\labels[4][25] , \labels[4].label[16] );
tran (\labels[4][26] , \labels[4].label[17] );
tran (\labels[4][27] , \labels[4].label[18] );
tran (\labels[4][28] , \labels[4].label[19] );
tran (\labels[4][29] , \labels[4].label[20] );
tran (\labels[4][30] , \labels[4].label[21] );
tran (\labels[4][31] , \labels[4].label[22] );
tran (\labels[4][32] , \labels[4].label[23] );
tran (\labels[4][33] , \labels[4].label[24] );
tran (\labels[4][34] , \labels[4].label[25] );
tran (\labels[4][35] , \labels[4].label[26] );
tran (\labels[4][36] , \labels[4].label[27] );
tran (\labels[4][37] , \labels[4].label[28] );
tran (\labels[4][38] , \labels[4].label[29] );
tran (\labels[4][39] , \labels[4].label[30] );
tran (\labels[4][40] , \labels[4].label[31] );
tran (\labels[4][41] , \labels[4].label[32] );
tran (\labels[4][42] , \labels[4].label[33] );
tran (\labels[4][43] , \labels[4].label[34] );
tran (\labels[4][44] , \labels[4].label[35] );
tran (\labels[4][45] , \labels[4].label[36] );
tran (\labels[4][46] , \labels[4].label[37] );
tran (\labels[4][47] , \labels[4].label[38] );
tran (\labels[4][48] , \labels[4].label[39] );
tran (\labels[4][49] , \labels[4].label[40] );
tran (\labels[4][50] , \labels[4].label[41] );
tran (\labels[4][51] , \labels[4].label[42] );
tran (\labels[4][52] , \labels[4].label[43] );
tran (\labels[4][53] , \labels[4].label[44] );
tran (\labels[4][54] , \labels[4].label[45] );
tran (\labels[4][55] , \labels[4].label[46] );
tran (\labels[4][56] , \labels[4].label[47] );
tran (\labels[4][57] , \labels[4].label[48] );
tran (\labels[4][58] , \labels[4].label[49] );
tran (\labels[4][59] , \labels[4].label[50] );
tran (\labels[4][60] , \labels[4].label[51] );
tran (\labels[4][61] , \labels[4].label[52] );
tran (\labels[4][62] , \labels[4].label[53] );
tran (\labels[4][63] , \labels[4].label[54] );
tran (\labels[4][64] , \labels[4].label[55] );
tran (\labels[4][65] , \labels[4].label[56] );
tran (\labels[4][66] , \labels[4].label[57] );
tran (\labels[4][67] , \labels[4].label[58] );
tran (\labels[4][68] , \labels[4].label[59] );
tran (\labels[4][69] , \labels[4].label[60] );
tran (\labels[4][70] , \labels[4].label[61] );
tran (\labels[4][71] , \labels[4].label[62] );
tran (\labels[4][72] , \labels[4].label[63] );
tran (\labels[4][73] , \labels[4].label[64] );
tran (\labels[4][74] , \labels[4].label[65] );
tran (\labels[4][75] , \labels[4].label[66] );
tran (\labels[4][76] , \labels[4].label[67] );
tran (\labels[4][77] , \labels[4].label[68] );
tran (\labels[4][78] , \labels[4].label[69] );
tran (\labels[4][79] , \labels[4].label[70] );
tran (\labels[4][80] , \labels[4].label[71] );
tran (\labels[4][81] , \labels[4].label[72] );
tran (\labels[4][82] , \labels[4].label[73] );
tran (\labels[4][83] , \labels[4].label[74] );
tran (\labels[4][84] , \labels[4].label[75] );
tran (\labels[4][85] , \labels[4].label[76] );
tran (\labels[4][86] , \labels[4].label[77] );
tran (\labels[4][87] , \labels[4].label[78] );
tran (\labels[4][88] , \labels[4].label[79] );
tran (\labels[4][89] , \labels[4].label[80] );
tran (\labels[4][90] , \labels[4].label[81] );
tran (\labels[4][91] , \labels[4].label[82] );
tran (\labels[4][92] , \labels[4].label[83] );
tran (\labels[4][93] , \labels[4].label[84] );
tran (\labels[4][94] , \labels[4].label[85] );
tran (\labels[4][95] , \labels[4].label[86] );
tran (\labels[4][96] , \labels[4].label[87] );
tran (\labels[4][97] , \labels[4].label[88] );
tran (\labels[4][98] , \labels[4].label[89] );
tran (\labels[4][99] , \labels[4].label[90] );
tran (\labels[4][100] , \labels[4].label[91] );
tran (\labels[4][101] , \labels[4].label[92] );
tran (\labels[4][102] , \labels[4].label[93] );
tran (\labels[4][103] , \labels[4].label[94] );
tran (\labels[4][104] , \labels[4].label[95] );
tran (\labels[4][105] , \labels[4].label[96] );
tran (\labels[4][106] , \labels[4].label[97] );
tran (\labels[4][107] , \labels[4].label[98] );
tran (\labels[4][108] , \labels[4].label[99] );
tran (\labels[4][109] , \labels[4].label[100] );
tran (\labels[4][110] , \labels[4].label[101] );
tran (\labels[4][111] , \labels[4].label[102] );
tran (\labels[4][112] , \labels[4].label[103] );
tran (\labels[4][113] , \labels[4].label[104] );
tran (\labels[4][114] , \labels[4].label[105] );
tran (\labels[4][115] , \labels[4].label[106] );
tran (\labels[4][116] , \labels[4].label[107] );
tran (\labels[4][117] , \labels[4].label[108] );
tran (\labels[4][118] , \labels[4].label[109] );
tran (\labels[4][119] , \labels[4].label[110] );
tran (\labels[4][120] , \labels[4].label[111] );
tran (\labels[4][121] , \labels[4].label[112] );
tran (\labels[4][122] , \labels[4].label[113] );
tran (\labels[4][123] , \labels[4].label[114] );
tran (\labels[4][124] , \labels[4].label[115] );
tran (\labels[4][125] , \labels[4].label[116] );
tran (\labels[4][126] , \labels[4].label[117] );
tran (\labels[4][127] , \labels[4].label[118] );
tran (\labels[4][128] , \labels[4].label[119] );
tran (\labels[4][129] , \labels[4].label[120] );
tran (\labels[4][130] , \labels[4].label[121] );
tran (\labels[4][131] , \labels[4].label[122] );
tran (\labels[4][132] , \labels[4].label[123] );
tran (\labels[4][133] , \labels[4].label[124] );
tran (\labels[4][134] , \labels[4].label[125] );
tran (\labels[4][135] , \labels[4].label[126] );
tran (\labels[4][136] , \labels[4].label[127] );
tran (\labels[4][137] , \labels[4].label[128] );
tran (\labels[4][138] , \labels[4].label[129] );
tran (\labels[4][139] , \labels[4].label[130] );
tran (\labels[4][140] , \labels[4].label[131] );
tran (\labels[4][141] , \labels[4].label[132] );
tran (\labels[4][142] , \labels[4].label[133] );
tran (\labels[4][143] , \labels[4].label[134] );
tran (\labels[4][144] , \labels[4].label[135] );
tran (\labels[4][145] , \labels[4].label[136] );
tran (\labels[4][146] , \labels[4].label[137] );
tran (\labels[4][147] , \labels[4].label[138] );
tran (\labels[4][148] , \labels[4].label[139] );
tran (\labels[4][149] , \labels[4].label[140] );
tran (\labels[4][150] , \labels[4].label[141] );
tran (\labels[4][151] , \labels[4].label[142] );
tran (\labels[4][152] , \labels[4].label[143] );
tran (\labels[4][153] , \labels[4].label[144] );
tran (\labels[4][154] , \labels[4].label[145] );
tran (\labels[4][155] , \labels[4].label[146] );
tran (\labels[4][156] , \labels[4].label[147] );
tran (\labels[4][157] , \labels[4].label[148] );
tran (\labels[4][158] , \labels[4].label[149] );
tran (\labels[4][159] , \labels[4].label[150] );
tran (\labels[4][160] , \labels[4].label[151] );
tran (\labels[4][161] , \labels[4].label[152] );
tran (\labels[4][162] , \labels[4].label[153] );
tran (\labels[4][163] , \labels[4].label[154] );
tran (\labels[4][164] , \labels[4].label[155] );
tran (\labels[4][165] , \labels[4].label[156] );
tran (\labels[4][166] , \labels[4].label[157] );
tran (\labels[4][167] , \labels[4].label[158] );
tran (\labels[4][168] , \labels[4].label[159] );
tran (\labels[4][169] , \labels[4].label[160] );
tran (\labels[4][170] , \labels[4].label[161] );
tran (\labels[4][171] , \labels[4].label[162] );
tran (\labels[4][172] , \labels[4].label[163] );
tran (\labels[4][173] , \labels[4].label[164] );
tran (\labels[4][174] , \labels[4].label[165] );
tran (\labels[4][175] , \labels[4].label[166] );
tran (\labels[4][176] , \labels[4].label[167] );
tran (\labels[4][177] , \labels[4].label[168] );
tran (\labels[4][178] , \labels[4].label[169] );
tran (\labels[4][179] , \labels[4].label[170] );
tran (\labels[4][180] , \labels[4].label[171] );
tran (\labels[4][181] , \labels[4].label[172] );
tran (\labels[4][182] , \labels[4].label[173] );
tran (\labels[4][183] , \labels[4].label[174] );
tran (\labels[4][184] , \labels[4].label[175] );
tran (\labels[4][185] , \labels[4].label[176] );
tran (\labels[4][186] , \labels[4].label[177] );
tran (\labels[4][187] , \labels[4].label[178] );
tran (\labels[4][188] , \labels[4].label[179] );
tran (\labels[4][189] , \labels[4].label[180] );
tran (\labels[4][190] , \labels[4].label[181] );
tran (\labels[4][191] , \labels[4].label[182] );
tran (\labels[4][192] , \labels[4].label[183] );
tran (\labels[4][193] , \labels[4].label[184] );
tran (\labels[4][194] , \labels[4].label[185] );
tran (\labels[4][195] , \labels[4].label[186] );
tran (\labels[4][196] , \labels[4].label[187] );
tran (\labels[4][197] , \labels[4].label[188] );
tran (\labels[4][198] , \labels[4].label[189] );
tran (\labels[4][199] , \labels[4].label[190] );
tran (\labels[4][200] , \labels[4].label[191] );
tran (\labels[4][201] , \labels[4].label[192] );
tran (\labels[4][202] , \labels[4].label[193] );
tran (\labels[4][203] , \labels[4].label[194] );
tran (\labels[4][204] , \labels[4].label[195] );
tran (\labels[4][205] , \labels[4].label[196] );
tran (\labels[4][206] , \labels[4].label[197] );
tran (\labels[4][207] , \labels[4].label[198] );
tran (\labels[4][208] , \labels[4].label[199] );
tran (\labels[4][209] , \labels[4].label[200] );
tran (\labels[4][210] , \labels[4].label[201] );
tran (\labels[4][211] , \labels[4].label[202] );
tran (\labels[4][212] , \labels[4].label[203] );
tran (\labels[4][213] , \labels[4].label[204] );
tran (\labels[4][214] , \labels[4].label[205] );
tran (\labels[4][215] , \labels[4].label[206] );
tran (\labels[4][216] , \labels[4].label[207] );
tran (\labels[4][217] , \labels[4].label[208] );
tran (\labels[4][218] , \labels[4].label[209] );
tran (\labels[4][219] , \labels[4].label[210] );
tran (\labels[4][220] , \labels[4].label[211] );
tran (\labels[4][221] , \labels[4].label[212] );
tran (\labels[4][222] , \labels[4].label[213] );
tran (\labels[4][223] , \labels[4].label[214] );
tran (\labels[4][224] , \labels[4].label[215] );
tran (\labels[4][225] , \labels[4].label[216] );
tran (\labels[4][226] , \labels[4].label[217] );
tran (\labels[4][227] , \labels[4].label[218] );
tran (\labels[4][228] , \labels[4].label[219] );
tran (\labels[4][229] , \labels[4].label[220] );
tran (\labels[4][230] , \labels[4].label[221] );
tran (\labels[4][231] , \labels[4].label[222] );
tran (\labels[4][232] , \labels[4].label[223] );
tran (\labels[4][233] , \labels[4].label[224] );
tran (\labels[4][234] , \labels[4].label[225] );
tran (\labels[4][235] , \labels[4].label[226] );
tran (\labels[4][236] , \labels[4].label[227] );
tran (\labels[4][237] , \labels[4].label[228] );
tran (\labels[4][238] , \labels[4].label[229] );
tran (\labels[4][239] , \labels[4].label[230] );
tran (\labels[4][240] , \labels[4].label[231] );
tran (\labels[4][241] , \labels[4].label[232] );
tran (\labels[4][242] , \labels[4].label[233] );
tran (\labels[4][243] , \labels[4].label[234] );
tran (\labels[4][244] , \labels[4].label[235] );
tran (\labels[4][245] , \labels[4].label[236] );
tran (\labels[4][246] , \labels[4].label[237] );
tran (\labels[4][247] , \labels[4].label[238] );
tran (\labels[4][248] , \labels[4].label[239] );
tran (\labels[4][249] , \labels[4].label[240] );
tran (\labels[4][250] , \labels[4].label[241] );
tran (\labels[4][251] , \labels[4].label[242] );
tran (\labels[4][252] , \labels[4].label[243] );
tran (\labels[4][253] , \labels[4].label[244] );
tran (\labels[4][254] , \labels[4].label[245] );
tran (\labels[4][255] , \labels[4].label[246] );
tran (\labels[4][256] , \labels[4].label[247] );
tran (\labels[4][257] , \labels[4].label[248] );
tran (\labels[4][258] , \labels[4].label[249] );
tran (\labels[4][259] , \labels[4].label[250] );
tran (\labels[4][260] , \labels[4].label[251] );
tran (\labels[4][261] , \labels[4].label[252] );
tran (\labels[4][262] , \labels[4].label[253] );
tran (\labels[4][263] , \labels[4].label[254] );
tran (\labels[4][264] , \labels[4].label[255] );
tran (\labels[4][265] , \labels[4].label_size[0] );
tran (\labels[4][266] , \labels[4].label_size[1] );
tran (\labels[4][267] , \labels[4].label_size[2] );
tran (\labels[4][268] , \labels[4].label_size[3] );
tran (\labels[4][269] , \labels[4].label_size[4] );
tran (\labels[4][270] , \labels[4].label_size[5] );
tran (\labels[4][271] , \labels[4].guid_size[0] );
tran (\labels[5][0] , \labels[5].delimiter[0] );
tran (\labels[5][1] , \labels[5].delimiter[1] );
tran (\labels[5][2] , \labels[5].delimiter[2] );
tran (\labels[5][3] , \labels[5].delimiter[3] );
tran (\labels[5][4] , \labels[5].delimiter[4] );
tran (\labels[5][5] , \labels[5].delimiter[5] );
tran (\labels[5][6] , \labels[5].delimiter[6] );
tran (\labels[5][7] , \labels[5].delimiter[7] );
tran (\labels[5][8] , \labels[5].delimiter_valid[0] );
tran (\labels[5][9] , \labels[5].label[0] );
tran (\labels[5][10] , \labels[5].label[1] );
tran (\labels[5][11] , \labels[5].label[2] );
tran (\labels[5][12] , \labels[5].label[3] );
tran (\labels[5][13] , \labels[5].label[4] );
tran (\labels[5][14] , \labels[5].label[5] );
tran (\labels[5][15] , \labels[5].label[6] );
tran (\labels[5][16] , \labels[5].label[7] );
tran (\labels[5][17] , \labels[5].label[8] );
tran (\labels[5][18] , \labels[5].label[9] );
tran (\labels[5][19] , \labels[5].label[10] );
tran (\labels[5][20] , \labels[5].label[11] );
tran (\labels[5][21] , \labels[5].label[12] );
tran (\labels[5][22] , \labels[5].label[13] );
tran (\labels[5][23] , \labels[5].label[14] );
tran (\labels[5][24] , \labels[5].label[15] );
tran (\labels[5][25] , \labels[5].label[16] );
tran (\labels[5][26] , \labels[5].label[17] );
tran (\labels[5][27] , \labels[5].label[18] );
tran (\labels[5][28] , \labels[5].label[19] );
tran (\labels[5][29] , \labels[5].label[20] );
tran (\labels[5][30] , \labels[5].label[21] );
tran (\labels[5][31] , \labels[5].label[22] );
tran (\labels[5][32] , \labels[5].label[23] );
tran (\labels[5][33] , \labels[5].label[24] );
tran (\labels[5][34] , \labels[5].label[25] );
tran (\labels[5][35] , \labels[5].label[26] );
tran (\labels[5][36] , \labels[5].label[27] );
tran (\labels[5][37] , \labels[5].label[28] );
tran (\labels[5][38] , \labels[5].label[29] );
tran (\labels[5][39] , \labels[5].label[30] );
tran (\labels[5][40] , \labels[5].label[31] );
tran (\labels[5][41] , \labels[5].label[32] );
tran (\labels[5][42] , \labels[5].label[33] );
tran (\labels[5][43] , \labels[5].label[34] );
tran (\labels[5][44] , \labels[5].label[35] );
tran (\labels[5][45] , \labels[5].label[36] );
tran (\labels[5][46] , \labels[5].label[37] );
tran (\labels[5][47] , \labels[5].label[38] );
tran (\labels[5][48] , \labels[5].label[39] );
tran (\labels[5][49] , \labels[5].label[40] );
tran (\labels[5][50] , \labels[5].label[41] );
tran (\labels[5][51] , \labels[5].label[42] );
tran (\labels[5][52] , \labels[5].label[43] );
tran (\labels[5][53] , \labels[5].label[44] );
tran (\labels[5][54] , \labels[5].label[45] );
tran (\labels[5][55] , \labels[5].label[46] );
tran (\labels[5][56] , \labels[5].label[47] );
tran (\labels[5][57] , \labels[5].label[48] );
tran (\labels[5][58] , \labels[5].label[49] );
tran (\labels[5][59] , \labels[5].label[50] );
tran (\labels[5][60] , \labels[5].label[51] );
tran (\labels[5][61] , \labels[5].label[52] );
tran (\labels[5][62] , \labels[5].label[53] );
tran (\labels[5][63] , \labels[5].label[54] );
tran (\labels[5][64] , \labels[5].label[55] );
tran (\labels[5][65] , \labels[5].label[56] );
tran (\labels[5][66] , \labels[5].label[57] );
tran (\labels[5][67] , \labels[5].label[58] );
tran (\labels[5][68] , \labels[5].label[59] );
tran (\labels[5][69] , \labels[5].label[60] );
tran (\labels[5][70] , \labels[5].label[61] );
tran (\labels[5][71] , \labels[5].label[62] );
tran (\labels[5][72] , \labels[5].label[63] );
tran (\labels[5][73] , \labels[5].label[64] );
tran (\labels[5][74] , \labels[5].label[65] );
tran (\labels[5][75] , \labels[5].label[66] );
tran (\labels[5][76] , \labels[5].label[67] );
tran (\labels[5][77] , \labels[5].label[68] );
tran (\labels[5][78] , \labels[5].label[69] );
tran (\labels[5][79] , \labels[5].label[70] );
tran (\labels[5][80] , \labels[5].label[71] );
tran (\labels[5][81] , \labels[5].label[72] );
tran (\labels[5][82] , \labels[5].label[73] );
tran (\labels[5][83] , \labels[5].label[74] );
tran (\labels[5][84] , \labels[5].label[75] );
tran (\labels[5][85] , \labels[5].label[76] );
tran (\labels[5][86] , \labels[5].label[77] );
tran (\labels[5][87] , \labels[5].label[78] );
tran (\labels[5][88] , \labels[5].label[79] );
tran (\labels[5][89] , \labels[5].label[80] );
tran (\labels[5][90] , \labels[5].label[81] );
tran (\labels[5][91] , \labels[5].label[82] );
tran (\labels[5][92] , \labels[5].label[83] );
tran (\labels[5][93] , \labels[5].label[84] );
tran (\labels[5][94] , \labels[5].label[85] );
tran (\labels[5][95] , \labels[5].label[86] );
tran (\labels[5][96] , \labels[5].label[87] );
tran (\labels[5][97] , \labels[5].label[88] );
tran (\labels[5][98] , \labels[5].label[89] );
tran (\labels[5][99] , \labels[5].label[90] );
tran (\labels[5][100] , \labels[5].label[91] );
tran (\labels[5][101] , \labels[5].label[92] );
tran (\labels[5][102] , \labels[5].label[93] );
tran (\labels[5][103] , \labels[5].label[94] );
tran (\labels[5][104] , \labels[5].label[95] );
tran (\labels[5][105] , \labels[5].label[96] );
tran (\labels[5][106] , \labels[5].label[97] );
tran (\labels[5][107] , \labels[5].label[98] );
tran (\labels[5][108] , \labels[5].label[99] );
tran (\labels[5][109] , \labels[5].label[100] );
tran (\labels[5][110] , \labels[5].label[101] );
tran (\labels[5][111] , \labels[5].label[102] );
tran (\labels[5][112] , \labels[5].label[103] );
tran (\labels[5][113] , \labels[5].label[104] );
tran (\labels[5][114] , \labels[5].label[105] );
tran (\labels[5][115] , \labels[5].label[106] );
tran (\labels[5][116] , \labels[5].label[107] );
tran (\labels[5][117] , \labels[5].label[108] );
tran (\labels[5][118] , \labels[5].label[109] );
tran (\labels[5][119] , \labels[5].label[110] );
tran (\labels[5][120] , \labels[5].label[111] );
tran (\labels[5][121] , \labels[5].label[112] );
tran (\labels[5][122] , \labels[5].label[113] );
tran (\labels[5][123] , \labels[5].label[114] );
tran (\labels[5][124] , \labels[5].label[115] );
tran (\labels[5][125] , \labels[5].label[116] );
tran (\labels[5][126] , \labels[5].label[117] );
tran (\labels[5][127] , \labels[5].label[118] );
tran (\labels[5][128] , \labels[5].label[119] );
tran (\labels[5][129] , \labels[5].label[120] );
tran (\labels[5][130] , \labels[5].label[121] );
tran (\labels[5][131] , \labels[5].label[122] );
tran (\labels[5][132] , \labels[5].label[123] );
tran (\labels[5][133] , \labels[5].label[124] );
tran (\labels[5][134] , \labels[5].label[125] );
tran (\labels[5][135] , \labels[5].label[126] );
tran (\labels[5][136] , \labels[5].label[127] );
tran (\labels[5][137] , \labels[5].label[128] );
tran (\labels[5][138] , \labels[5].label[129] );
tran (\labels[5][139] , \labels[5].label[130] );
tran (\labels[5][140] , \labels[5].label[131] );
tran (\labels[5][141] , \labels[5].label[132] );
tran (\labels[5][142] , \labels[5].label[133] );
tran (\labels[5][143] , \labels[5].label[134] );
tran (\labels[5][144] , \labels[5].label[135] );
tran (\labels[5][145] , \labels[5].label[136] );
tran (\labels[5][146] , \labels[5].label[137] );
tran (\labels[5][147] , \labels[5].label[138] );
tran (\labels[5][148] , \labels[5].label[139] );
tran (\labels[5][149] , \labels[5].label[140] );
tran (\labels[5][150] , \labels[5].label[141] );
tran (\labels[5][151] , \labels[5].label[142] );
tran (\labels[5][152] , \labels[5].label[143] );
tran (\labels[5][153] , \labels[5].label[144] );
tran (\labels[5][154] , \labels[5].label[145] );
tran (\labels[5][155] , \labels[5].label[146] );
tran (\labels[5][156] , \labels[5].label[147] );
tran (\labels[5][157] , \labels[5].label[148] );
tran (\labels[5][158] , \labels[5].label[149] );
tran (\labels[5][159] , \labels[5].label[150] );
tran (\labels[5][160] , \labels[5].label[151] );
tran (\labels[5][161] , \labels[5].label[152] );
tran (\labels[5][162] , \labels[5].label[153] );
tran (\labels[5][163] , \labels[5].label[154] );
tran (\labels[5][164] , \labels[5].label[155] );
tran (\labels[5][165] , \labels[5].label[156] );
tran (\labels[5][166] , \labels[5].label[157] );
tran (\labels[5][167] , \labels[5].label[158] );
tran (\labels[5][168] , \labels[5].label[159] );
tran (\labels[5][169] , \labels[5].label[160] );
tran (\labels[5][170] , \labels[5].label[161] );
tran (\labels[5][171] , \labels[5].label[162] );
tran (\labels[5][172] , \labels[5].label[163] );
tran (\labels[5][173] , \labels[5].label[164] );
tran (\labels[5][174] , \labels[5].label[165] );
tran (\labels[5][175] , \labels[5].label[166] );
tran (\labels[5][176] , \labels[5].label[167] );
tran (\labels[5][177] , \labels[5].label[168] );
tran (\labels[5][178] , \labels[5].label[169] );
tran (\labels[5][179] , \labels[5].label[170] );
tran (\labels[5][180] , \labels[5].label[171] );
tran (\labels[5][181] , \labels[5].label[172] );
tran (\labels[5][182] , \labels[5].label[173] );
tran (\labels[5][183] , \labels[5].label[174] );
tran (\labels[5][184] , \labels[5].label[175] );
tran (\labels[5][185] , \labels[5].label[176] );
tran (\labels[5][186] , \labels[5].label[177] );
tran (\labels[5][187] , \labels[5].label[178] );
tran (\labels[5][188] , \labels[5].label[179] );
tran (\labels[5][189] , \labels[5].label[180] );
tran (\labels[5][190] , \labels[5].label[181] );
tran (\labels[5][191] , \labels[5].label[182] );
tran (\labels[5][192] , \labels[5].label[183] );
tran (\labels[5][193] , \labels[5].label[184] );
tran (\labels[5][194] , \labels[5].label[185] );
tran (\labels[5][195] , \labels[5].label[186] );
tran (\labels[5][196] , \labels[5].label[187] );
tran (\labels[5][197] , \labels[5].label[188] );
tran (\labels[5][198] , \labels[5].label[189] );
tran (\labels[5][199] , \labels[5].label[190] );
tran (\labels[5][200] , \labels[5].label[191] );
tran (\labels[5][201] , \labels[5].label[192] );
tran (\labels[5][202] , \labels[5].label[193] );
tran (\labels[5][203] , \labels[5].label[194] );
tran (\labels[5][204] , \labels[5].label[195] );
tran (\labels[5][205] , \labels[5].label[196] );
tran (\labels[5][206] , \labels[5].label[197] );
tran (\labels[5][207] , \labels[5].label[198] );
tran (\labels[5][208] , \labels[5].label[199] );
tran (\labels[5][209] , \labels[5].label[200] );
tran (\labels[5][210] , \labels[5].label[201] );
tran (\labels[5][211] , \labels[5].label[202] );
tran (\labels[5][212] , \labels[5].label[203] );
tran (\labels[5][213] , \labels[5].label[204] );
tran (\labels[5][214] , \labels[5].label[205] );
tran (\labels[5][215] , \labels[5].label[206] );
tran (\labels[5][216] , \labels[5].label[207] );
tran (\labels[5][217] , \labels[5].label[208] );
tran (\labels[5][218] , \labels[5].label[209] );
tran (\labels[5][219] , \labels[5].label[210] );
tran (\labels[5][220] , \labels[5].label[211] );
tran (\labels[5][221] , \labels[5].label[212] );
tran (\labels[5][222] , \labels[5].label[213] );
tran (\labels[5][223] , \labels[5].label[214] );
tran (\labels[5][224] , \labels[5].label[215] );
tran (\labels[5][225] , \labels[5].label[216] );
tran (\labels[5][226] , \labels[5].label[217] );
tran (\labels[5][227] , \labels[5].label[218] );
tran (\labels[5][228] , \labels[5].label[219] );
tran (\labels[5][229] , \labels[5].label[220] );
tran (\labels[5][230] , \labels[5].label[221] );
tran (\labels[5][231] , \labels[5].label[222] );
tran (\labels[5][232] , \labels[5].label[223] );
tran (\labels[5][233] , \labels[5].label[224] );
tran (\labels[5][234] , \labels[5].label[225] );
tran (\labels[5][235] , \labels[5].label[226] );
tran (\labels[5][236] , \labels[5].label[227] );
tran (\labels[5][237] , \labels[5].label[228] );
tran (\labels[5][238] , \labels[5].label[229] );
tran (\labels[5][239] , \labels[5].label[230] );
tran (\labels[5][240] , \labels[5].label[231] );
tran (\labels[5][241] , \labels[5].label[232] );
tran (\labels[5][242] , \labels[5].label[233] );
tran (\labels[5][243] , \labels[5].label[234] );
tran (\labels[5][244] , \labels[5].label[235] );
tran (\labels[5][245] , \labels[5].label[236] );
tran (\labels[5][246] , \labels[5].label[237] );
tran (\labels[5][247] , \labels[5].label[238] );
tran (\labels[5][248] , \labels[5].label[239] );
tran (\labels[5][249] , \labels[5].label[240] );
tran (\labels[5][250] , \labels[5].label[241] );
tran (\labels[5][251] , \labels[5].label[242] );
tran (\labels[5][252] , \labels[5].label[243] );
tran (\labels[5][253] , \labels[5].label[244] );
tran (\labels[5][254] , \labels[5].label[245] );
tran (\labels[5][255] , \labels[5].label[246] );
tran (\labels[5][256] , \labels[5].label[247] );
tran (\labels[5][257] , \labels[5].label[248] );
tran (\labels[5][258] , \labels[5].label[249] );
tran (\labels[5][259] , \labels[5].label[250] );
tran (\labels[5][260] , \labels[5].label[251] );
tran (\labels[5][261] , \labels[5].label[252] );
tran (\labels[5][262] , \labels[5].label[253] );
tran (\labels[5][263] , \labels[5].label[254] );
tran (\labels[5][264] , \labels[5].label[255] );
tran (\labels[5][265] , \labels[5].label_size[0] );
tran (\labels[5][266] , \labels[5].label_size[1] );
tran (\labels[5][267] , \labels[5].label_size[2] );
tran (\labels[5][268] , \labels[5].label_size[3] );
tran (\labels[5][269] , \labels[5].label_size[4] );
tran (\labels[5][270] , \labels[5].label_size[5] );
tran (\labels[5][271] , \labels[5].guid_size[0] );
tran (\labels[6][0] , \labels[6].delimiter[0] );
tran (\labels[6][1] , \labels[6].delimiter[1] );
tran (\labels[6][2] , \labels[6].delimiter[2] );
tran (\labels[6][3] , \labels[6].delimiter[3] );
tran (\labels[6][4] , \labels[6].delimiter[4] );
tran (\labels[6][5] , \labels[6].delimiter[5] );
tran (\labels[6][6] , \labels[6].delimiter[6] );
tran (\labels[6][7] , \labels[6].delimiter[7] );
tran (\labels[6][8] , \labels[6].delimiter_valid[0] );
tran (\labels[6][9] , \labels[6].label[0] );
tran (\labels[6][10] , \labels[6].label[1] );
tran (\labels[6][11] , \labels[6].label[2] );
tran (\labels[6][12] , \labels[6].label[3] );
tran (\labels[6][13] , \labels[6].label[4] );
tran (\labels[6][14] , \labels[6].label[5] );
tran (\labels[6][15] , \labels[6].label[6] );
tran (\labels[6][16] , \labels[6].label[7] );
tran (\labels[6][17] , \labels[6].label[8] );
tran (\labels[6][18] , \labels[6].label[9] );
tran (\labels[6][19] , \labels[6].label[10] );
tran (\labels[6][20] , \labels[6].label[11] );
tran (\labels[6][21] , \labels[6].label[12] );
tran (\labels[6][22] , \labels[6].label[13] );
tran (\labels[6][23] , \labels[6].label[14] );
tran (\labels[6][24] , \labels[6].label[15] );
tran (\labels[6][25] , \labels[6].label[16] );
tran (\labels[6][26] , \labels[6].label[17] );
tran (\labels[6][27] , \labels[6].label[18] );
tran (\labels[6][28] , \labels[6].label[19] );
tran (\labels[6][29] , \labels[6].label[20] );
tran (\labels[6][30] , \labels[6].label[21] );
tran (\labels[6][31] , \labels[6].label[22] );
tran (\labels[6][32] , \labels[6].label[23] );
tran (\labels[6][33] , \labels[6].label[24] );
tran (\labels[6][34] , \labels[6].label[25] );
tran (\labels[6][35] , \labels[6].label[26] );
tran (\labels[6][36] , \labels[6].label[27] );
tran (\labels[6][37] , \labels[6].label[28] );
tran (\labels[6][38] , \labels[6].label[29] );
tran (\labels[6][39] , \labels[6].label[30] );
tran (\labels[6][40] , \labels[6].label[31] );
tran (\labels[6][41] , \labels[6].label[32] );
tran (\labels[6][42] , \labels[6].label[33] );
tran (\labels[6][43] , \labels[6].label[34] );
tran (\labels[6][44] , \labels[6].label[35] );
tran (\labels[6][45] , \labels[6].label[36] );
tran (\labels[6][46] , \labels[6].label[37] );
tran (\labels[6][47] , \labels[6].label[38] );
tran (\labels[6][48] , \labels[6].label[39] );
tran (\labels[6][49] , \labels[6].label[40] );
tran (\labels[6][50] , \labels[6].label[41] );
tran (\labels[6][51] , \labels[6].label[42] );
tran (\labels[6][52] , \labels[6].label[43] );
tran (\labels[6][53] , \labels[6].label[44] );
tran (\labels[6][54] , \labels[6].label[45] );
tran (\labels[6][55] , \labels[6].label[46] );
tran (\labels[6][56] , \labels[6].label[47] );
tran (\labels[6][57] , \labels[6].label[48] );
tran (\labels[6][58] , \labels[6].label[49] );
tran (\labels[6][59] , \labels[6].label[50] );
tran (\labels[6][60] , \labels[6].label[51] );
tran (\labels[6][61] , \labels[6].label[52] );
tran (\labels[6][62] , \labels[6].label[53] );
tran (\labels[6][63] , \labels[6].label[54] );
tran (\labels[6][64] , \labels[6].label[55] );
tran (\labels[6][65] , \labels[6].label[56] );
tran (\labels[6][66] , \labels[6].label[57] );
tran (\labels[6][67] , \labels[6].label[58] );
tran (\labels[6][68] , \labels[6].label[59] );
tran (\labels[6][69] , \labels[6].label[60] );
tran (\labels[6][70] , \labels[6].label[61] );
tran (\labels[6][71] , \labels[6].label[62] );
tran (\labels[6][72] , \labels[6].label[63] );
tran (\labels[6][73] , \labels[6].label[64] );
tran (\labels[6][74] , \labels[6].label[65] );
tran (\labels[6][75] , \labels[6].label[66] );
tran (\labels[6][76] , \labels[6].label[67] );
tran (\labels[6][77] , \labels[6].label[68] );
tran (\labels[6][78] , \labels[6].label[69] );
tran (\labels[6][79] , \labels[6].label[70] );
tran (\labels[6][80] , \labels[6].label[71] );
tran (\labels[6][81] , \labels[6].label[72] );
tran (\labels[6][82] , \labels[6].label[73] );
tran (\labels[6][83] , \labels[6].label[74] );
tran (\labels[6][84] , \labels[6].label[75] );
tran (\labels[6][85] , \labels[6].label[76] );
tran (\labels[6][86] , \labels[6].label[77] );
tran (\labels[6][87] , \labels[6].label[78] );
tran (\labels[6][88] , \labels[6].label[79] );
tran (\labels[6][89] , \labels[6].label[80] );
tran (\labels[6][90] , \labels[6].label[81] );
tran (\labels[6][91] , \labels[6].label[82] );
tran (\labels[6][92] , \labels[6].label[83] );
tran (\labels[6][93] , \labels[6].label[84] );
tran (\labels[6][94] , \labels[6].label[85] );
tran (\labels[6][95] , \labels[6].label[86] );
tran (\labels[6][96] , \labels[6].label[87] );
tran (\labels[6][97] , \labels[6].label[88] );
tran (\labels[6][98] , \labels[6].label[89] );
tran (\labels[6][99] , \labels[6].label[90] );
tran (\labels[6][100] , \labels[6].label[91] );
tran (\labels[6][101] , \labels[6].label[92] );
tran (\labels[6][102] , \labels[6].label[93] );
tran (\labels[6][103] , \labels[6].label[94] );
tran (\labels[6][104] , \labels[6].label[95] );
tran (\labels[6][105] , \labels[6].label[96] );
tran (\labels[6][106] , \labels[6].label[97] );
tran (\labels[6][107] , \labels[6].label[98] );
tran (\labels[6][108] , \labels[6].label[99] );
tran (\labels[6][109] , \labels[6].label[100] );
tran (\labels[6][110] , \labels[6].label[101] );
tran (\labels[6][111] , \labels[6].label[102] );
tran (\labels[6][112] , \labels[6].label[103] );
tran (\labels[6][113] , \labels[6].label[104] );
tran (\labels[6][114] , \labels[6].label[105] );
tran (\labels[6][115] , \labels[6].label[106] );
tran (\labels[6][116] , \labels[6].label[107] );
tran (\labels[6][117] , \labels[6].label[108] );
tran (\labels[6][118] , \labels[6].label[109] );
tran (\labels[6][119] , \labels[6].label[110] );
tran (\labels[6][120] , \labels[6].label[111] );
tran (\labels[6][121] , \labels[6].label[112] );
tran (\labels[6][122] , \labels[6].label[113] );
tran (\labels[6][123] , \labels[6].label[114] );
tran (\labels[6][124] , \labels[6].label[115] );
tran (\labels[6][125] , \labels[6].label[116] );
tran (\labels[6][126] , \labels[6].label[117] );
tran (\labels[6][127] , \labels[6].label[118] );
tran (\labels[6][128] , \labels[6].label[119] );
tran (\labels[6][129] , \labels[6].label[120] );
tran (\labels[6][130] , \labels[6].label[121] );
tran (\labels[6][131] , \labels[6].label[122] );
tran (\labels[6][132] , \labels[6].label[123] );
tran (\labels[6][133] , \labels[6].label[124] );
tran (\labels[6][134] , \labels[6].label[125] );
tran (\labels[6][135] , \labels[6].label[126] );
tran (\labels[6][136] , \labels[6].label[127] );
tran (\labels[6][137] , \labels[6].label[128] );
tran (\labels[6][138] , \labels[6].label[129] );
tran (\labels[6][139] , \labels[6].label[130] );
tran (\labels[6][140] , \labels[6].label[131] );
tran (\labels[6][141] , \labels[6].label[132] );
tran (\labels[6][142] , \labels[6].label[133] );
tran (\labels[6][143] , \labels[6].label[134] );
tran (\labels[6][144] , \labels[6].label[135] );
tran (\labels[6][145] , \labels[6].label[136] );
tran (\labels[6][146] , \labels[6].label[137] );
tran (\labels[6][147] , \labels[6].label[138] );
tran (\labels[6][148] , \labels[6].label[139] );
tran (\labels[6][149] , \labels[6].label[140] );
tran (\labels[6][150] , \labels[6].label[141] );
tran (\labels[6][151] , \labels[6].label[142] );
tran (\labels[6][152] , \labels[6].label[143] );
tran (\labels[6][153] , \labels[6].label[144] );
tran (\labels[6][154] , \labels[6].label[145] );
tran (\labels[6][155] , \labels[6].label[146] );
tran (\labels[6][156] , \labels[6].label[147] );
tran (\labels[6][157] , \labels[6].label[148] );
tran (\labels[6][158] , \labels[6].label[149] );
tran (\labels[6][159] , \labels[6].label[150] );
tran (\labels[6][160] , \labels[6].label[151] );
tran (\labels[6][161] , \labels[6].label[152] );
tran (\labels[6][162] , \labels[6].label[153] );
tran (\labels[6][163] , \labels[6].label[154] );
tran (\labels[6][164] , \labels[6].label[155] );
tran (\labels[6][165] , \labels[6].label[156] );
tran (\labels[6][166] , \labels[6].label[157] );
tran (\labels[6][167] , \labels[6].label[158] );
tran (\labels[6][168] , \labels[6].label[159] );
tran (\labels[6][169] , \labels[6].label[160] );
tran (\labels[6][170] , \labels[6].label[161] );
tran (\labels[6][171] , \labels[6].label[162] );
tran (\labels[6][172] , \labels[6].label[163] );
tran (\labels[6][173] , \labels[6].label[164] );
tran (\labels[6][174] , \labels[6].label[165] );
tran (\labels[6][175] , \labels[6].label[166] );
tran (\labels[6][176] , \labels[6].label[167] );
tran (\labels[6][177] , \labels[6].label[168] );
tran (\labels[6][178] , \labels[6].label[169] );
tran (\labels[6][179] , \labels[6].label[170] );
tran (\labels[6][180] , \labels[6].label[171] );
tran (\labels[6][181] , \labels[6].label[172] );
tran (\labels[6][182] , \labels[6].label[173] );
tran (\labels[6][183] , \labels[6].label[174] );
tran (\labels[6][184] , \labels[6].label[175] );
tran (\labels[6][185] , \labels[6].label[176] );
tran (\labels[6][186] , \labels[6].label[177] );
tran (\labels[6][187] , \labels[6].label[178] );
tran (\labels[6][188] , \labels[6].label[179] );
tran (\labels[6][189] , \labels[6].label[180] );
tran (\labels[6][190] , \labels[6].label[181] );
tran (\labels[6][191] , \labels[6].label[182] );
tran (\labels[6][192] , \labels[6].label[183] );
tran (\labels[6][193] , \labels[6].label[184] );
tran (\labels[6][194] , \labels[6].label[185] );
tran (\labels[6][195] , \labels[6].label[186] );
tran (\labels[6][196] , \labels[6].label[187] );
tran (\labels[6][197] , \labels[6].label[188] );
tran (\labels[6][198] , \labels[6].label[189] );
tran (\labels[6][199] , \labels[6].label[190] );
tran (\labels[6][200] , \labels[6].label[191] );
tran (\labels[6][201] , \labels[6].label[192] );
tran (\labels[6][202] , \labels[6].label[193] );
tran (\labels[6][203] , \labels[6].label[194] );
tran (\labels[6][204] , \labels[6].label[195] );
tran (\labels[6][205] , \labels[6].label[196] );
tran (\labels[6][206] , \labels[6].label[197] );
tran (\labels[6][207] , \labels[6].label[198] );
tran (\labels[6][208] , \labels[6].label[199] );
tran (\labels[6][209] , \labels[6].label[200] );
tran (\labels[6][210] , \labels[6].label[201] );
tran (\labels[6][211] , \labels[6].label[202] );
tran (\labels[6][212] , \labels[6].label[203] );
tran (\labels[6][213] , \labels[6].label[204] );
tran (\labels[6][214] , \labels[6].label[205] );
tran (\labels[6][215] , \labels[6].label[206] );
tran (\labels[6][216] , \labels[6].label[207] );
tran (\labels[6][217] , \labels[6].label[208] );
tran (\labels[6][218] , \labels[6].label[209] );
tran (\labels[6][219] , \labels[6].label[210] );
tran (\labels[6][220] , \labels[6].label[211] );
tran (\labels[6][221] , \labels[6].label[212] );
tran (\labels[6][222] , \labels[6].label[213] );
tran (\labels[6][223] , \labels[6].label[214] );
tran (\labels[6][224] , \labels[6].label[215] );
tran (\labels[6][225] , \labels[6].label[216] );
tran (\labels[6][226] , \labels[6].label[217] );
tran (\labels[6][227] , \labels[6].label[218] );
tran (\labels[6][228] , \labels[6].label[219] );
tran (\labels[6][229] , \labels[6].label[220] );
tran (\labels[6][230] , \labels[6].label[221] );
tran (\labels[6][231] , \labels[6].label[222] );
tran (\labels[6][232] , \labels[6].label[223] );
tran (\labels[6][233] , \labels[6].label[224] );
tran (\labels[6][234] , \labels[6].label[225] );
tran (\labels[6][235] , \labels[6].label[226] );
tran (\labels[6][236] , \labels[6].label[227] );
tran (\labels[6][237] , \labels[6].label[228] );
tran (\labels[6][238] , \labels[6].label[229] );
tran (\labels[6][239] , \labels[6].label[230] );
tran (\labels[6][240] , \labels[6].label[231] );
tran (\labels[6][241] , \labels[6].label[232] );
tran (\labels[6][242] , \labels[6].label[233] );
tran (\labels[6][243] , \labels[6].label[234] );
tran (\labels[6][244] , \labels[6].label[235] );
tran (\labels[6][245] , \labels[6].label[236] );
tran (\labels[6][246] , \labels[6].label[237] );
tran (\labels[6][247] , \labels[6].label[238] );
tran (\labels[6][248] , \labels[6].label[239] );
tran (\labels[6][249] , \labels[6].label[240] );
tran (\labels[6][250] , \labels[6].label[241] );
tran (\labels[6][251] , \labels[6].label[242] );
tran (\labels[6][252] , \labels[6].label[243] );
tran (\labels[6][253] , \labels[6].label[244] );
tran (\labels[6][254] , \labels[6].label[245] );
tran (\labels[6][255] , \labels[6].label[246] );
tran (\labels[6][256] , \labels[6].label[247] );
tran (\labels[6][257] , \labels[6].label[248] );
tran (\labels[6][258] , \labels[6].label[249] );
tran (\labels[6][259] , \labels[6].label[250] );
tran (\labels[6][260] , \labels[6].label[251] );
tran (\labels[6][261] , \labels[6].label[252] );
tran (\labels[6][262] , \labels[6].label[253] );
tran (\labels[6][263] , \labels[6].label[254] );
tran (\labels[6][264] , \labels[6].label[255] );
tran (\labels[6][265] , \labels[6].label_size[0] );
tran (\labels[6][266] , \labels[6].label_size[1] );
tran (\labels[6][267] , \labels[6].label_size[2] );
tran (\labels[6][268] , \labels[6].label_size[3] );
tran (\labels[6][269] , \labels[6].label_size[4] );
tran (\labels[6][270] , \labels[6].label_size[5] );
tran (\labels[6][271] , \labels[6].guid_size[0] );
tran (\labels[7][0] , \labels[7].delimiter[0] );
tran (\labels[7][1] , \labels[7].delimiter[1] );
tran (\labels[7][2] , \labels[7].delimiter[2] );
tran (\labels[7][3] , \labels[7].delimiter[3] );
tran (\labels[7][4] , \labels[7].delimiter[4] );
tran (\labels[7][5] , \labels[7].delimiter[5] );
tran (\labels[7][6] , \labels[7].delimiter[6] );
tran (\labels[7][7] , \labels[7].delimiter[7] );
tran (\labels[7][8] , \labels[7].delimiter_valid[0] );
tran (\labels[7][9] , \labels[7].label[0] );
tran (\labels[7][10] , \labels[7].label[1] );
tran (\labels[7][11] , \labels[7].label[2] );
tran (\labels[7][12] , \labels[7].label[3] );
tran (\labels[7][13] , \labels[7].label[4] );
tran (\labels[7][14] , \labels[7].label[5] );
tran (\labels[7][15] , \labels[7].label[6] );
tran (\labels[7][16] , \labels[7].label[7] );
tran (\labels[7][17] , \labels[7].label[8] );
tran (\labels[7][18] , \labels[7].label[9] );
tran (\labels[7][19] , \labels[7].label[10] );
tran (\labels[7][20] , \labels[7].label[11] );
tran (\labels[7][21] , \labels[7].label[12] );
tran (\labels[7][22] , \labels[7].label[13] );
tran (\labels[7][23] , \labels[7].label[14] );
tran (\labels[7][24] , \labels[7].label[15] );
tran (\labels[7][25] , \labels[7].label[16] );
tran (\labels[7][26] , \labels[7].label[17] );
tran (\labels[7][27] , \labels[7].label[18] );
tran (\labels[7][28] , \labels[7].label[19] );
tran (\labels[7][29] , \labels[7].label[20] );
tran (\labels[7][30] , \labels[7].label[21] );
tran (\labels[7][31] , \labels[7].label[22] );
tran (\labels[7][32] , \labels[7].label[23] );
tran (\labels[7][33] , \labels[7].label[24] );
tran (\labels[7][34] , \labels[7].label[25] );
tran (\labels[7][35] , \labels[7].label[26] );
tran (\labels[7][36] , \labels[7].label[27] );
tran (\labels[7][37] , \labels[7].label[28] );
tran (\labels[7][38] , \labels[7].label[29] );
tran (\labels[7][39] , \labels[7].label[30] );
tran (\labels[7][40] , \labels[7].label[31] );
tran (\labels[7][41] , \labels[7].label[32] );
tran (\labels[7][42] , \labels[7].label[33] );
tran (\labels[7][43] , \labels[7].label[34] );
tran (\labels[7][44] , \labels[7].label[35] );
tran (\labels[7][45] , \labels[7].label[36] );
tran (\labels[7][46] , \labels[7].label[37] );
tran (\labels[7][47] , \labels[7].label[38] );
tran (\labels[7][48] , \labels[7].label[39] );
tran (\labels[7][49] , \labels[7].label[40] );
tran (\labels[7][50] , \labels[7].label[41] );
tran (\labels[7][51] , \labels[7].label[42] );
tran (\labels[7][52] , \labels[7].label[43] );
tran (\labels[7][53] , \labels[7].label[44] );
tran (\labels[7][54] , \labels[7].label[45] );
tran (\labels[7][55] , \labels[7].label[46] );
tran (\labels[7][56] , \labels[7].label[47] );
tran (\labels[7][57] , \labels[7].label[48] );
tran (\labels[7][58] , \labels[7].label[49] );
tran (\labels[7][59] , \labels[7].label[50] );
tran (\labels[7][60] , \labels[7].label[51] );
tran (\labels[7][61] , \labels[7].label[52] );
tran (\labels[7][62] , \labels[7].label[53] );
tran (\labels[7][63] , \labels[7].label[54] );
tran (\labels[7][64] , \labels[7].label[55] );
tran (\labels[7][65] , \labels[7].label[56] );
tran (\labels[7][66] , \labels[7].label[57] );
tran (\labels[7][67] , \labels[7].label[58] );
tran (\labels[7][68] , \labels[7].label[59] );
tran (\labels[7][69] , \labels[7].label[60] );
tran (\labels[7][70] , \labels[7].label[61] );
tran (\labels[7][71] , \labels[7].label[62] );
tran (\labels[7][72] , \labels[7].label[63] );
tran (\labels[7][73] , \labels[7].label[64] );
tran (\labels[7][74] , \labels[7].label[65] );
tran (\labels[7][75] , \labels[7].label[66] );
tran (\labels[7][76] , \labels[7].label[67] );
tran (\labels[7][77] , \labels[7].label[68] );
tran (\labels[7][78] , \labels[7].label[69] );
tran (\labels[7][79] , \labels[7].label[70] );
tran (\labels[7][80] , \labels[7].label[71] );
tran (\labels[7][81] , \labels[7].label[72] );
tran (\labels[7][82] , \labels[7].label[73] );
tran (\labels[7][83] , \labels[7].label[74] );
tran (\labels[7][84] , \labels[7].label[75] );
tran (\labels[7][85] , \labels[7].label[76] );
tran (\labels[7][86] , \labels[7].label[77] );
tran (\labels[7][87] , \labels[7].label[78] );
tran (\labels[7][88] , \labels[7].label[79] );
tran (\labels[7][89] , \labels[7].label[80] );
tran (\labels[7][90] , \labels[7].label[81] );
tran (\labels[7][91] , \labels[7].label[82] );
tran (\labels[7][92] , \labels[7].label[83] );
tran (\labels[7][93] , \labels[7].label[84] );
tran (\labels[7][94] , \labels[7].label[85] );
tran (\labels[7][95] , \labels[7].label[86] );
tran (\labels[7][96] , \labels[7].label[87] );
tran (\labels[7][97] , \labels[7].label[88] );
tran (\labels[7][98] , \labels[7].label[89] );
tran (\labels[7][99] , \labels[7].label[90] );
tran (\labels[7][100] , \labels[7].label[91] );
tran (\labels[7][101] , \labels[7].label[92] );
tran (\labels[7][102] , \labels[7].label[93] );
tran (\labels[7][103] , \labels[7].label[94] );
tran (\labels[7][104] , \labels[7].label[95] );
tran (\labels[7][105] , \labels[7].label[96] );
tran (\labels[7][106] , \labels[7].label[97] );
tran (\labels[7][107] , \labels[7].label[98] );
tran (\labels[7][108] , \labels[7].label[99] );
tran (\labels[7][109] , \labels[7].label[100] );
tran (\labels[7][110] , \labels[7].label[101] );
tran (\labels[7][111] , \labels[7].label[102] );
tran (\labels[7][112] , \labels[7].label[103] );
tran (\labels[7][113] , \labels[7].label[104] );
tran (\labels[7][114] , \labels[7].label[105] );
tran (\labels[7][115] , \labels[7].label[106] );
tran (\labels[7][116] , \labels[7].label[107] );
tran (\labels[7][117] , \labels[7].label[108] );
tran (\labels[7][118] , \labels[7].label[109] );
tran (\labels[7][119] , \labels[7].label[110] );
tran (\labels[7][120] , \labels[7].label[111] );
tran (\labels[7][121] , \labels[7].label[112] );
tran (\labels[7][122] , \labels[7].label[113] );
tran (\labels[7][123] , \labels[7].label[114] );
tran (\labels[7][124] , \labels[7].label[115] );
tran (\labels[7][125] , \labels[7].label[116] );
tran (\labels[7][126] , \labels[7].label[117] );
tran (\labels[7][127] , \labels[7].label[118] );
tran (\labels[7][128] , \labels[7].label[119] );
tran (\labels[7][129] , \labels[7].label[120] );
tran (\labels[7][130] , \labels[7].label[121] );
tran (\labels[7][131] , \labels[7].label[122] );
tran (\labels[7][132] , \labels[7].label[123] );
tran (\labels[7][133] , \labels[7].label[124] );
tran (\labels[7][134] , \labels[7].label[125] );
tran (\labels[7][135] , \labels[7].label[126] );
tran (\labels[7][136] , \labels[7].label[127] );
tran (\labels[7][137] , \labels[7].label[128] );
tran (\labels[7][138] , \labels[7].label[129] );
tran (\labels[7][139] , \labels[7].label[130] );
tran (\labels[7][140] , \labels[7].label[131] );
tran (\labels[7][141] , \labels[7].label[132] );
tran (\labels[7][142] , \labels[7].label[133] );
tran (\labels[7][143] , \labels[7].label[134] );
tran (\labels[7][144] , \labels[7].label[135] );
tran (\labels[7][145] , \labels[7].label[136] );
tran (\labels[7][146] , \labels[7].label[137] );
tran (\labels[7][147] , \labels[7].label[138] );
tran (\labels[7][148] , \labels[7].label[139] );
tran (\labels[7][149] , \labels[7].label[140] );
tran (\labels[7][150] , \labels[7].label[141] );
tran (\labels[7][151] , \labels[7].label[142] );
tran (\labels[7][152] , \labels[7].label[143] );
tran (\labels[7][153] , \labels[7].label[144] );
tran (\labels[7][154] , \labels[7].label[145] );
tran (\labels[7][155] , \labels[7].label[146] );
tran (\labels[7][156] , \labels[7].label[147] );
tran (\labels[7][157] , \labels[7].label[148] );
tran (\labels[7][158] , \labels[7].label[149] );
tran (\labels[7][159] , \labels[7].label[150] );
tran (\labels[7][160] , \labels[7].label[151] );
tran (\labels[7][161] , \labels[7].label[152] );
tran (\labels[7][162] , \labels[7].label[153] );
tran (\labels[7][163] , \labels[7].label[154] );
tran (\labels[7][164] , \labels[7].label[155] );
tran (\labels[7][165] , \labels[7].label[156] );
tran (\labels[7][166] , \labels[7].label[157] );
tran (\labels[7][167] , \labels[7].label[158] );
tran (\labels[7][168] , \labels[7].label[159] );
tran (\labels[7][169] , \labels[7].label[160] );
tran (\labels[7][170] , \labels[7].label[161] );
tran (\labels[7][171] , \labels[7].label[162] );
tran (\labels[7][172] , \labels[7].label[163] );
tran (\labels[7][173] , \labels[7].label[164] );
tran (\labels[7][174] , \labels[7].label[165] );
tran (\labels[7][175] , \labels[7].label[166] );
tran (\labels[7][176] , \labels[7].label[167] );
tran (\labels[7][177] , \labels[7].label[168] );
tran (\labels[7][178] , \labels[7].label[169] );
tran (\labels[7][179] , \labels[7].label[170] );
tran (\labels[7][180] , \labels[7].label[171] );
tran (\labels[7][181] , \labels[7].label[172] );
tran (\labels[7][182] , \labels[7].label[173] );
tran (\labels[7][183] , \labels[7].label[174] );
tran (\labels[7][184] , \labels[7].label[175] );
tran (\labels[7][185] , \labels[7].label[176] );
tran (\labels[7][186] , \labels[7].label[177] );
tran (\labels[7][187] , \labels[7].label[178] );
tran (\labels[7][188] , \labels[7].label[179] );
tran (\labels[7][189] , \labels[7].label[180] );
tran (\labels[7][190] , \labels[7].label[181] );
tran (\labels[7][191] , \labels[7].label[182] );
tran (\labels[7][192] , \labels[7].label[183] );
tran (\labels[7][193] , \labels[7].label[184] );
tran (\labels[7][194] , \labels[7].label[185] );
tran (\labels[7][195] , \labels[7].label[186] );
tran (\labels[7][196] , \labels[7].label[187] );
tran (\labels[7][197] , \labels[7].label[188] );
tran (\labels[7][198] , \labels[7].label[189] );
tran (\labels[7][199] , \labels[7].label[190] );
tran (\labels[7][200] , \labels[7].label[191] );
tran (\labels[7][201] , \labels[7].label[192] );
tran (\labels[7][202] , \labels[7].label[193] );
tran (\labels[7][203] , \labels[7].label[194] );
tran (\labels[7][204] , \labels[7].label[195] );
tran (\labels[7][205] , \labels[7].label[196] );
tran (\labels[7][206] , \labels[7].label[197] );
tran (\labels[7][207] , \labels[7].label[198] );
tran (\labels[7][208] , \labels[7].label[199] );
tran (\labels[7][209] , \labels[7].label[200] );
tran (\labels[7][210] , \labels[7].label[201] );
tran (\labels[7][211] , \labels[7].label[202] );
tran (\labels[7][212] , \labels[7].label[203] );
tran (\labels[7][213] , \labels[7].label[204] );
tran (\labels[7][214] , \labels[7].label[205] );
tran (\labels[7][215] , \labels[7].label[206] );
tran (\labels[7][216] , \labels[7].label[207] );
tran (\labels[7][217] , \labels[7].label[208] );
tran (\labels[7][218] , \labels[7].label[209] );
tran (\labels[7][219] , \labels[7].label[210] );
tran (\labels[7][220] , \labels[7].label[211] );
tran (\labels[7][221] , \labels[7].label[212] );
tran (\labels[7][222] , \labels[7].label[213] );
tran (\labels[7][223] , \labels[7].label[214] );
tran (\labels[7][224] , \labels[7].label[215] );
tran (\labels[7][225] , \labels[7].label[216] );
tran (\labels[7][226] , \labels[7].label[217] );
tran (\labels[7][227] , \labels[7].label[218] );
tran (\labels[7][228] , \labels[7].label[219] );
tran (\labels[7][229] , \labels[7].label[220] );
tran (\labels[7][230] , \labels[7].label[221] );
tran (\labels[7][231] , \labels[7].label[222] );
tran (\labels[7][232] , \labels[7].label[223] );
tran (\labels[7][233] , \labels[7].label[224] );
tran (\labels[7][234] , \labels[7].label[225] );
tran (\labels[7][235] , \labels[7].label[226] );
tran (\labels[7][236] , \labels[7].label[227] );
tran (\labels[7][237] , \labels[7].label[228] );
tran (\labels[7][238] , \labels[7].label[229] );
tran (\labels[7][239] , \labels[7].label[230] );
tran (\labels[7][240] , \labels[7].label[231] );
tran (\labels[7][241] , \labels[7].label[232] );
tran (\labels[7][242] , \labels[7].label[233] );
tran (\labels[7][243] , \labels[7].label[234] );
tran (\labels[7][244] , \labels[7].label[235] );
tran (\labels[7][245] , \labels[7].label[236] );
tran (\labels[7][246] , \labels[7].label[237] );
tran (\labels[7][247] , \labels[7].label[238] );
tran (\labels[7][248] , \labels[7].label[239] );
tran (\labels[7][249] , \labels[7].label[240] );
tran (\labels[7][250] , \labels[7].label[241] );
tran (\labels[7][251] , \labels[7].label[242] );
tran (\labels[7][252] , \labels[7].label[243] );
tran (\labels[7][253] , \labels[7].label[244] );
tran (\labels[7][254] , \labels[7].label[245] );
tran (\labels[7][255] , \labels[7].label[246] );
tran (\labels[7][256] , \labels[7].label[247] );
tran (\labels[7][257] , \labels[7].label[248] );
tran (\labels[7][258] , \labels[7].label[249] );
tran (\labels[7][259] , \labels[7].label[250] );
tran (\labels[7][260] , \labels[7].label[251] );
tran (\labels[7][261] , \labels[7].label[252] );
tran (\labels[7][262] , \labels[7].label[253] );
tran (\labels[7][263] , \labels[7].label[254] );
tran (\labels[7][264] , \labels[7].label[255] );
tran (\labels[7][265] , \labels[7].label_size[0] );
tran (\labels[7][266] , \labels[7].label_size[1] );
tran (\labels[7][267] , \labels[7].label_size[2] );
tran (\labels[7][268] , \labels[7].label_size[3] );
tran (\labels[7][269] , \labels[7].label_size[4] );
tran (\labels[7][270] , \labels[7].label_size[5] );
tran (\labels[7][271] , \labels[7].guid_size[0] );
tran (kme_internal_out[70], \kme_internal_out.sot [0]);
tran (kme_internal_out[69], \kme_internal_out.eoi [0]);
tran (kme_internal_out[68], \kme_internal_out.eot [0]);
tran (kme_internal_out[67], \kme_internal_out.id [3]);
tran (kme_internal_out[66], \kme_internal_out.id [2]);
tran (kme_internal_out[65], \kme_internal_out.id [1]);
tran (kme_internal_out[64], \kme_internal_out.id [0]);
tran (kme_internal_out[63], \kme_internal_out.tdata [63]);
tran (kme_internal_out[62], \kme_internal_out.tdata [62]);
tran (kme_internal_out[61], \kme_internal_out.tdata [61]);
tran (kme_internal_out[60], \kme_internal_out.tdata [60]);
tran (kme_internal_out[59], \kme_internal_out.tdata [59]);
tran (kme_internal_out[58], \kme_internal_out.tdata [58]);
tran (kme_internal_out[57], \kme_internal_out.tdata [57]);
tran (kme_internal_out[56], \kme_internal_out.tdata [56]);
tran (kme_internal_out[55], \kme_internal_out.tdata [55]);
tran (kme_internal_out[54], \kme_internal_out.tdata [54]);
tran (kme_internal_out[53], \kme_internal_out.tdata [53]);
tran (kme_internal_out[52], \kme_internal_out.tdata [52]);
tran (kme_internal_out[51], \kme_internal_out.tdata [51]);
tran (kme_internal_out[50], \kme_internal_out.tdata [50]);
tran (kme_internal_out[49], \kme_internal_out.tdata [49]);
tran (kme_internal_out[48], \kme_internal_out.tdata [48]);
tran (kme_internal_out[47], \kme_internal_out.tdata [47]);
tran (kme_internal_out[46], \kme_internal_out.tdata [46]);
tran (kme_internal_out[45], \kme_internal_out.tdata [45]);
tran (kme_internal_out[44], \kme_internal_out.tdata [44]);
tran (kme_internal_out[43], \kme_internal_out.tdata [43]);
tran (kme_internal_out[42], \kme_internal_out.tdata [42]);
tran (kme_internal_out[41], \kme_internal_out.tdata [41]);
tran (kme_internal_out[40], \kme_internal_out.tdata [40]);
tran (kme_internal_out[39], \kme_internal_out.tdata [39]);
tran (kme_internal_out[38], \kme_internal_out.tdata [38]);
tran (kme_internal_out[37], \kme_internal_out.tdata [37]);
tran (kme_internal_out[36], \kme_internal_out.tdata [36]);
tran (kme_internal_out[35], \kme_internal_out.tdata [35]);
tran (kme_internal_out[34], \kme_internal_out.tdata [34]);
tran (kme_internal_out[33], \kme_internal_out.tdata [33]);
tran (kme_internal_out[32], \kme_internal_out.tdata [32]);
tran (kme_internal_out[31], \kme_internal_out.tdata [31]);
tran (kme_internal_out[30], \kme_internal_out.tdata [30]);
tran (kme_internal_out[29], \kme_internal_out.tdata [29]);
tran (kme_internal_out[28], \kme_internal_out.tdata [28]);
tran (kme_internal_out[27], \kme_internal_out.tdata [27]);
tran (kme_internal_out[26], \kme_internal_out.tdata [26]);
tran (kme_internal_out[25], \kme_internal_out.tdata [25]);
tran (kme_internal_out[24], \kme_internal_out.tdata [24]);
tran (kme_internal_out[23], \kme_internal_out.tdata [23]);
tran (kme_internal_out[22], \kme_internal_out.tdata [22]);
tran (kme_internal_out[21], \kme_internal_out.tdata [21]);
tran (kme_internal_out[20], \kme_internal_out.tdata [20]);
tran (kme_internal_out[19], \kme_internal_out.tdata [19]);
tran (kme_internal_out[18], \kme_internal_out.tdata [18]);
tran (kme_internal_out[17], \kme_internal_out.tdata [17]);
tran (kme_internal_out[16], \kme_internal_out.tdata [16]);
tran (kme_internal_out[15], \kme_internal_out.tdata [15]);
tran (kme_internal_out[14], \kme_internal_out.tdata [14]);
tran (kme_internal_out[13], \kme_internal_out.tdata [13]);
tran (kme_internal_out[12], \kme_internal_out.tdata [12]);
tran (kme_internal_out[11], \kme_internal_out.tdata [11]);
tran (kme_internal_out[10], \kme_internal_out.tdata [10]);
tran (kme_internal_out[9], \kme_internal_out.tdata [9]);
tran (kme_internal_out[8], \kme_internal_out.tdata [8]);
tran (kme_internal_out[7], \kme_internal_out.tdata [7]);
tran (kme_internal_out[6], \kme_internal_out.tdata [6]);
tran (kme_internal_out[5], \kme_internal_out.tdata [5]);
tran (kme_internal_out[4], \kme_internal_out.tdata [4]);
tran (kme_internal_out[3], \kme_internal_out.tdata [3]);
tran (kme_internal_out[2], \kme_internal_out.tdata [2]);
tran (kme_internal_out[1], \kme_internal_out.tdata [1]);
tran (kme_internal_out[0], \kme_internal_out.tdata [0]);
tran (kop_fifo_override[6], \kop_fifo_override.r.part0 [6]);
tran (kop_fifo_override[6], \kop_fifo_override.f.gcm_status_data_fifo );
tran (kop_fifo_override[5], \kop_fifo_override.r.part0 [5]);
tran (kop_fifo_override[5], \kop_fifo_override.f.tlv_sb_data_fifo );
tran (kop_fifo_override[4], \kop_fifo_override.r.part0 [4]);
tran (kop_fifo_override[4], \kop_fifo_override.f.kdf_cmd_fifo );
tran (kop_fifo_override[3], \kop_fifo_override.r.part0 [3]);
tran (kop_fifo_override[3], \kop_fifo_override.f.kdfstream_cmd_fifo );
tran (kop_fifo_override[2], \kop_fifo_override.r.part0 [2]);
tran (kop_fifo_override[2], \kop_fifo_override.f.keyfilter_cmd_fifo );
tran (kop_fifo_override[1], \kop_fifo_override.r.part0 [1]);
tran (kop_fifo_override[1], \kop_fifo_override.f.gcm_tag_data_fifo );
tran (kop_fifo_override[0], \kop_fifo_override.r.part0 [0]);
tran (kop_fifo_override[0], \kop_fifo_override.f.gcm_cmd_fifo );
tran (gcm_cmd_in[610], \gcm_cmd_in.key0 [255]);
tran (gcm_cmd_in[609], \gcm_cmd_in.key0 [254]);
tran (gcm_cmd_in[608], \gcm_cmd_in.key0 [253]);
tran (gcm_cmd_in[607], \gcm_cmd_in.key0 [252]);
tran (gcm_cmd_in[606], \gcm_cmd_in.key0 [251]);
tran (gcm_cmd_in[605], \gcm_cmd_in.key0 [250]);
tran (gcm_cmd_in[604], \gcm_cmd_in.key0 [249]);
tran (gcm_cmd_in[603], \gcm_cmd_in.key0 [248]);
tran (gcm_cmd_in[602], \gcm_cmd_in.key0 [247]);
tran (gcm_cmd_in[601], \gcm_cmd_in.key0 [246]);
tran (gcm_cmd_in[600], \gcm_cmd_in.key0 [245]);
tran (gcm_cmd_in[599], \gcm_cmd_in.key0 [244]);
tran (gcm_cmd_in[598], \gcm_cmd_in.key0 [243]);
tran (gcm_cmd_in[597], \gcm_cmd_in.key0 [242]);
tran (gcm_cmd_in[596], \gcm_cmd_in.key0 [241]);
tran (gcm_cmd_in[595], \gcm_cmd_in.key0 [240]);
tran (gcm_cmd_in[594], \gcm_cmd_in.key0 [239]);
tran (gcm_cmd_in[593], \gcm_cmd_in.key0 [238]);
tran (gcm_cmd_in[592], \gcm_cmd_in.key0 [237]);
tran (gcm_cmd_in[591], \gcm_cmd_in.key0 [236]);
tran (gcm_cmd_in[590], \gcm_cmd_in.key0 [235]);
tran (gcm_cmd_in[589], \gcm_cmd_in.key0 [234]);
tran (gcm_cmd_in[588], \gcm_cmd_in.key0 [233]);
tran (gcm_cmd_in[587], \gcm_cmd_in.key0 [232]);
tran (gcm_cmd_in[586], \gcm_cmd_in.key0 [231]);
tran (gcm_cmd_in[585], \gcm_cmd_in.key0 [230]);
tran (gcm_cmd_in[584], \gcm_cmd_in.key0 [229]);
tran (gcm_cmd_in[583], \gcm_cmd_in.key0 [228]);
tran (gcm_cmd_in[582], \gcm_cmd_in.key0 [227]);
tran (gcm_cmd_in[581], \gcm_cmd_in.key0 [226]);
tran (gcm_cmd_in[580], \gcm_cmd_in.key0 [225]);
tran (gcm_cmd_in[579], \gcm_cmd_in.key0 [224]);
tran (gcm_cmd_in[578], \gcm_cmd_in.key0 [223]);
tran (gcm_cmd_in[577], \gcm_cmd_in.key0 [222]);
tran (gcm_cmd_in[576], \gcm_cmd_in.key0 [221]);
tran (gcm_cmd_in[575], \gcm_cmd_in.key0 [220]);
tran (gcm_cmd_in[574], \gcm_cmd_in.key0 [219]);
tran (gcm_cmd_in[573], \gcm_cmd_in.key0 [218]);
tran (gcm_cmd_in[572], \gcm_cmd_in.key0 [217]);
tran (gcm_cmd_in[571], \gcm_cmd_in.key0 [216]);
tran (gcm_cmd_in[570], \gcm_cmd_in.key0 [215]);
tran (gcm_cmd_in[569], \gcm_cmd_in.key0 [214]);
tran (gcm_cmd_in[568], \gcm_cmd_in.key0 [213]);
tran (gcm_cmd_in[567], \gcm_cmd_in.key0 [212]);
tran (gcm_cmd_in[566], \gcm_cmd_in.key0 [211]);
tran (gcm_cmd_in[565], \gcm_cmd_in.key0 [210]);
tran (gcm_cmd_in[564], \gcm_cmd_in.key0 [209]);
tran (gcm_cmd_in[563], \gcm_cmd_in.key0 [208]);
tran (gcm_cmd_in[562], \gcm_cmd_in.key0 [207]);
tran (gcm_cmd_in[561], \gcm_cmd_in.key0 [206]);
tran (gcm_cmd_in[560], \gcm_cmd_in.key0 [205]);
tran (gcm_cmd_in[559], \gcm_cmd_in.key0 [204]);
tran (gcm_cmd_in[558], \gcm_cmd_in.key0 [203]);
tran (gcm_cmd_in[557], \gcm_cmd_in.key0 [202]);
tran (gcm_cmd_in[556], \gcm_cmd_in.key0 [201]);
tran (gcm_cmd_in[555], \gcm_cmd_in.key0 [200]);
tran (gcm_cmd_in[554], \gcm_cmd_in.key0 [199]);
tran (gcm_cmd_in[553], \gcm_cmd_in.key0 [198]);
tran (gcm_cmd_in[552], \gcm_cmd_in.key0 [197]);
tran (gcm_cmd_in[551], \gcm_cmd_in.key0 [196]);
tran (gcm_cmd_in[550], \gcm_cmd_in.key0 [195]);
tran (gcm_cmd_in[549], \gcm_cmd_in.key0 [194]);
tran (gcm_cmd_in[548], \gcm_cmd_in.key0 [193]);
tran (gcm_cmd_in[547], \gcm_cmd_in.key0 [192]);
tran (gcm_cmd_in[546], \gcm_cmd_in.key0 [191]);
tran (gcm_cmd_in[545], \gcm_cmd_in.key0 [190]);
tran (gcm_cmd_in[544], \gcm_cmd_in.key0 [189]);
tran (gcm_cmd_in[543], \gcm_cmd_in.key0 [188]);
tran (gcm_cmd_in[542], \gcm_cmd_in.key0 [187]);
tran (gcm_cmd_in[541], \gcm_cmd_in.key0 [186]);
tran (gcm_cmd_in[540], \gcm_cmd_in.key0 [185]);
tran (gcm_cmd_in[539], \gcm_cmd_in.key0 [184]);
tran (gcm_cmd_in[538], \gcm_cmd_in.key0 [183]);
tran (gcm_cmd_in[537], \gcm_cmd_in.key0 [182]);
tran (gcm_cmd_in[536], \gcm_cmd_in.key0 [181]);
tran (gcm_cmd_in[535], \gcm_cmd_in.key0 [180]);
tran (gcm_cmd_in[534], \gcm_cmd_in.key0 [179]);
tran (gcm_cmd_in[533], \gcm_cmd_in.key0 [178]);
tran (gcm_cmd_in[532], \gcm_cmd_in.key0 [177]);
tran (gcm_cmd_in[531], \gcm_cmd_in.key0 [176]);
tran (gcm_cmd_in[530], \gcm_cmd_in.key0 [175]);
tran (gcm_cmd_in[529], \gcm_cmd_in.key0 [174]);
tran (gcm_cmd_in[528], \gcm_cmd_in.key0 [173]);
tran (gcm_cmd_in[527], \gcm_cmd_in.key0 [172]);
tran (gcm_cmd_in[526], \gcm_cmd_in.key0 [171]);
tran (gcm_cmd_in[525], \gcm_cmd_in.key0 [170]);
tran (gcm_cmd_in[524], \gcm_cmd_in.key0 [169]);
tran (gcm_cmd_in[523], \gcm_cmd_in.key0 [168]);
tran (gcm_cmd_in[522], \gcm_cmd_in.key0 [167]);
tran (gcm_cmd_in[521], \gcm_cmd_in.key0 [166]);
tran (gcm_cmd_in[520], \gcm_cmd_in.key0 [165]);
tran (gcm_cmd_in[519], \gcm_cmd_in.key0 [164]);
tran (gcm_cmd_in[518], \gcm_cmd_in.key0 [163]);
tran (gcm_cmd_in[517], \gcm_cmd_in.key0 [162]);
tran (gcm_cmd_in[516], \gcm_cmd_in.key0 [161]);
tran (gcm_cmd_in[515], \gcm_cmd_in.key0 [160]);
tran (gcm_cmd_in[514], \gcm_cmd_in.key0 [159]);
tran (gcm_cmd_in[513], \gcm_cmd_in.key0 [158]);
tran (gcm_cmd_in[512], \gcm_cmd_in.key0 [157]);
tran (gcm_cmd_in[511], \gcm_cmd_in.key0 [156]);
tran (gcm_cmd_in[510], \gcm_cmd_in.key0 [155]);
tran (gcm_cmd_in[509], \gcm_cmd_in.key0 [154]);
tran (gcm_cmd_in[508], \gcm_cmd_in.key0 [153]);
tran (gcm_cmd_in[507], \gcm_cmd_in.key0 [152]);
tran (gcm_cmd_in[506], \gcm_cmd_in.key0 [151]);
tran (gcm_cmd_in[505], \gcm_cmd_in.key0 [150]);
tran (gcm_cmd_in[504], \gcm_cmd_in.key0 [149]);
tran (gcm_cmd_in[503], \gcm_cmd_in.key0 [148]);
tran (gcm_cmd_in[502], \gcm_cmd_in.key0 [147]);
tran (gcm_cmd_in[501], \gcm_cmd_in.key0 [146]);
tran (gcm_cmd_in[500], \gcm_cmd_in.key0 [145]);
tran (gcm_cmd_in[499], \gcm_cmd_in.key0 [144]);
tran (gcm_cmd_in[498], \gcm_cmd_in.key0 [143]);
tran (gcm_cmd_in[497], \gcm_cmd_in.key0 [142]);
tran (gcm_cmd_in[496], \gcm_cmd_in.key0 [141]);
tran (gcm_cmd_in[495], \gcm_cmd_in.key0 [140]);
tran (gcm_cmd_in[494], \gcm_cmd_in.key0 [139]);
tran (gcm_cmd_in[493], \gcm_cmd_in.key0 [138]);
tran (gcm_cmd_in[492], \gcm_cmd_in.key0 [137]);
tran (gcm_cmd_in[491], \gcm_cmd_in.key0 [136]);
tran (gcm_cmd_in[490], \gcm_cmd_in.key0 [135]);
tran (gcm_cmd_in[489], \gcm_cmd_in.key0 [134]);
tran (gcm_cmd_in[488], \gcm_cmd_in.key0 [133]);
tran (gcm_cmd_in[487], \gcm_cmd_in.key0 [132]);
tran (gcm_cmd_in[486], \gcm_cmd_in.key0 [131]);
tran (gcm_cmd_in[485], \gcm_cmd_in.key0 [130]);
tran (gcm_cmd_in[484], \gcm_cmd_in.key0 [129]);
tran (gcm_cmd_in[483], \gcm_cmd_in.key0 [128]);
tran (gcm_cmd_in[482], \gcm_cmd_in.key0 [127]);
tran (gcm_cmd_in[481], \gcm_cmd_in.key0 [126]);
tran (gcm_cmd_in[480], \gcm_cmd_in.key0 [125]);
tran (gcm_cmd_in[479], \gcm_cmd_in.key0 [124]);
tran (gcm_cmd_in[478], \gcm_cmd_in.key0 [123]);
tran (gcm_cmd_in[477], \gcm_cmd_in.key0 [122]);
tran (gcm_cmd_in[476], \gcm_cmd_in.key0 [121]);
tran (gcm_cmd_in[475], \gcm_cmd_in.key0 [120]);
tran (gcm_cmd_in[474], \gcm_cmd_in.key0 [119]);
tran (gcm_cmd_in[473], \gcm_cmd_in.key0 [118]);
tran (gcm_cmd_in[472], \gcm_cmd_in.key0 [117]);
tran (gcm_cmd_in[471], \gcm_cmd_in.key0 [116]);
tran (gcm_cmd_in[470], \gcm_cmd_in.key0 [115]);
tran (gcm_cmd_in[469], \gcm_cmd_in.key0 [114]);
tran (gcm_cmd_in[468], \gcm_cmd_in.key0 [113]);
tran (gcm_cmd_in[467], \gcm_cmd_in.key0 [112]);
tran (gcm_cmd_in[466], \gcm_cmd_in.key0 [111]);
tran (gcm_cmd_in[465], \gcm_cmd_in.key0 [110]);
tran (gcm_cmd_in[464], \gcm_cmd_in.key0 [109]);
tran (gcm_cmd_in[463], \gcm_cmd_in.key0 [108]);
tran (gcm_cmd_in[462], \gcm_cmd_in.key0 [107]);
tran (gcm_cmd_in[461], \gcm_cmd_in.key0 [106]);
tran (gcm_cmd_in[460], \gcm_cmd_in.key0 [105]);
tran (gcm_cmd_in[459], \gcm_cmd_in.key0 [104]);
tran (gcm_cmd_in[458], \gcm_cmd_in.key0 [103]);
tran (gcm_cmd_in[457], \gcm_cmd_in.key0 [102]);
tran (gcm_cmd_in[456], \gcm_cmd_in.key0 [101]);
tran (gcm_cmd_in[455], \gcm_cmd_in.key0 [100]);
tran (gcm_cmd_in[454], \gcm_cmd_in.key0 [99]);
tran (gcm_cmd_in[453], \gcm_cmd_in.key0 [98]);
tran (gcm_cmd_in[452], \gcm_cmd_in.key0 [97]);
tran (gcm_cmd_in[451], \gcm_cmd_in.key0 [96]);
tran (gcm_cmd_in[450], \gcm_cmd_in.key0 [95]);
tran (gcm_cmd_in[449], \gcm_cmd_in.key0 [94]);
tran (gcm_cmd_in[448], \gcm_cmd_in.key0 [93]);
tran (gcm_cmd_in[447], \gcm_cmd_in.key0 [92]);
tran (gcm_cmd_in[446], \gcm_cmd_in.key0 [91]);
tran (gcm_cmd_in[445], \gcm_cmd_in.key0 [90]);
tran (gcm_cmd_in[444], \gcm_cmd_in.key0 [89]);
tran (gcm_cmd_in[443], \gcm_cmd_in.key0 [88]);
tran (gcm_cmd_in[442], \gcm_cmd_in.key0 [87]);
tran (gcm_cmd_in[441], \gcm_cmd_in.key0 [86]);
tran (gcm_cmd_in[440], \gcm_cmd_in.key0 [85]);
tran (gcm_cmd_in[439], \gcm_cmd_in.key0 [84]);
tran (gcm_cmd_in[438], \gcm_cmd_in.key0 [83]);
tran (gcm_cmd_in[437], \gcm_cmd_in.key0 [82]);
tran (gcm_cmd_in[436], \gcm_cmd_in.key0 [81]);
tran (gcm_cmd_in[435], \gcm_cmd_in.key0 [80]);
tran (gcm_cmd_in[434], \gcm_cmd_in.key0 [79]);
tran (gcm_cmd_in[433], \gcm_cmd_in.key0 [78]);
tran (gcm_cmd_in[432], \gcm_cmd_in.key0 [77]);
tran (gcm_cmd_in[431], \gcm_cmd_in.key0 [76]);
tran (gcm_cmd_in[430], \gcm_cmd_in.key0 [75]);
tran (gcm_cmd_in[429], \gcm_cmd_in.key0 [74]);
tran (gcm_cmd_in[428], \gcm_cmd_in.key0 [73]);
tran (gcm_cmd_in[427], \gcm_cmd_in.key0 [72]);
tran (gcm_cmd_in[426], \gcm_cmd_in.key0 [71]);
tran (gcm_cmd_in[425], \gcm_cmd_in.key0 [70]);
tran (gcm_cmd_in[424], \gcm_cmd_in.key0 [69]);
tran (gcm_cmd_in[423], \gcm_cmd_in.key0 [68]);
tran (gcm_cmd_in[422], \gcm_cmd_in.key0 [67]);
tran (gcm_cmd_in[421], \gcm_cmd_in.key0 [66]);
tran (gcm_cmd_in[420], \gcm_cmd_in.key0 [65]);
tran (gcm_cmd_in[419], \gcm_cmd_in.key0 [64]);
tran (gcm_cmd_in[418], \gcm_cmd_in.key0 [63]);
tran (gcm_cmd_in[417], \gcm_cmd_in.key0 [62]);
tran (gcm_cmd_in[416], \gcm_cmd_in.key0 [61]);
tran (gcm_cmd_in[415], \gcm_cmd_in.key0 [60]);
tran (gcm_cmd_in[414], \gcm_cmd_in.key0 [59]);
tran (gcm_cmd_in[413], \gcm_cmd_in.key0 [58]);
tran (gcm_cmd_in[412], \gcm_cmd_in.key0 [57]);
tran (gcm_cmd_in[411], \gcm_cmd_in.key0 [56]);
tran (gcm_cmd_in[410], \gcm_cmd_in.key0 [55]);
tran (gcm_cmd_in[409], \gcm_cmd_in.key0 [54]);
tran (gcm_cmd_in[408], \gcm_cmd_in.key0 [53]);
tran (gcm_cmd_in[407], \gcm_cmd_in.key0 [52]);
tran (gcm_cmd_in[406], \gcm_cmd_in.key0 [51]);
tran (gcm_cmd_in[405], \gcm_cmd_in.key0 [50]);
tran (gcm_cmd_in[404], \gcm_cmd_in.key0 [49]);
tran (gcm_cmd_in[403], \gcm_cmd_in.key0 [48]);
tran (gcm_cmd_in[402], \gcm_cmd_in.key0 [47]);
tran (gcm_cmd_in[401], \gcm_cmd_in.key0 [46]);
tran (gcm_cmd_in[400], \gcm_cmd_in.key0 [45]);
tran (gcm_cmd_in[399], \gcm_cmd_in.key0 [44]);
tran (gcm_cmd_in[398], \gcm_cmd_in.key0 [43]);
tran (gcm_cmd_in[397], \gcm_cmd_in.key0 [42]);
tran (gcm_cmd_in[396], \gcm_cmd_in.key0 [41]);
tran (gcm_cmd_in[395], \gcm_cmd_in.key0 [40]);
tran (gcm_cmd_in[394], \gcm_cmd_in.key0 [39]);
tran (gcm_cmd_in[393], \gcm_cmd_in.key0 [38]);
tran (gcm_cmd_in[392], \gcm_cmd_in.key0 [37]);
tran (gcm_cmd_in[391], \gcm_cmd_in.key0 [36]);
tran (gcm_cmd_in[390], \gcm_cmd_in.key0 [35]);
tran (gcm_cmd_in[389], \gcm_cmd_in.key0 [34]);
tran (gcm_cmd_in[388], \gcm_cmd_in.key0 [33]);
tran (gcm_cmd_in[387], \gcm_cmd_in.key0 [32]);
tran (gcm_cmd_in[386], \gcm_cmd_in.key0 [31]);
tran (gcm_cmd_in[385], \gcm_cmd_in.key0 [30]);
tran (gcm_cmd_in[384], \gcm_cmd_in.key0 [29]);
tran (gcm_cmd_in[383], \gcm_cmd_in.key0 [28]);
tran (gcm_cmd_in[382], \gcm_cmd_in.key0 [27]);
tran (gcm_cmd_in[381], \gcm_cmd_in.key0 [26]);
tran (gcm_cmd_in[380], \gcm_cmd_in.key0 [25]);
tran (gcm_cmd_in[379], \gcm_cmd_in.key0 [24]);
tran (gcm_cmd_in[378], \gcm_cmd_in.key0 [23]);
tran (gcm_cmd_in[377], \gcm_cmd_in.key0 [22]);
tran (gcm_cmd_in[376], \gcm_cmd_in.key0 [21]);
tran (gcm_cmd_in[375], \gcm_cmd_in.key0 [20]);
tran (gcm_cmd_in[374], \gcm_cmd_in.key0 [19]);
tran (gcm_cmd_in[373], \gcm_cmd_in.key0 [18]);
tran (gcm_cmd_in[372], \gcm_cmd_in.key0 [17]);
tran (gcm_cmd_in[371], \gcm_cmd_in.key0 [16]);
tran (gcm_cmd_in[370], \gcm_cmd_in.key0 [15]);
tran (gcm_cmd_in[369], \gcm_cmd_in.key0 [14]);
tran (gcm_cmd_in[368], \gcm_cmd_in.key0 [13]);
tran (gcm_cmd_in[367], \gcm_cmd_in.key0 [12]);
tran (gcm_cmd_in[366], \gcm_cmd_in.key0 [11]);
tran (gcm_cmd_in[365], \gcm_cmd_in.key0 [10]);
tran (gcm_cmd_in[364], \gcm_cmd_in.key0 [9]);
tran (gcm_cmd_in[363], \gcm_cmd_in.key0 [8]);
tran (gcm_cmd_in[362], \gcm_cmd_in.key0 [7]);
tran (gcm_cmd_in[361], \gcm_cmd_in.key0 [6]);
tran (gcm_cmd_in[360], \gcm_cmd_in.key0 [5]);
tran (gcm_cmd_in[359], \gcm_cmd_in.key0 [4]);
tran (gcm_cmd_in[358], \gcm_cmd_in.key0 [3]);
tran (gcm_cmd_in[357], \gcm_cmd_in.key0 [2]);
tran (gcm_cmd_in[356], \gcm_cmd_in.key0 [1]);
tran (gcm_cmd_in[355], \gcm_cmd_in.key0 [0]);
tran (gcm_cmd_in[354], \gcm_cmd_in.key1 [255]);
tran (gcm_cmd_in[353], \gcm_cmd_in.key1 [254]);
tran (gcm_cmd_in[352], \gcm_cmd_in.key1 [253]);
tran (gcm_cmd_in[351], \gcm_cmd_in.key1 [252]);
tran (gcm_cmd_in[350], \gcm_cmd_in.key1 [251]);
tran (gcm_cmd_in[349], \gcm_cmd_in.key1 [250]);
tran (gcm_cmd_in[348], \gcm_cmd_in.key1 [249]);
tran (gcm_cmd_in[347], \gcm_cmd_in.key1 [248]);
tran (gcm_cmd_in[346], \gcm_cmd_in.key1 [247]);
tran (gcm_cmd_in[345], \gcm_cmd_in.key1 [246]);
tran (gcm_cmd_in[344], \gcm_cmd_in.key1 [245]);
tran (gcm_cmd_in[343], \gcm_cmd_in.key1 [244]);
tran (gcm_cmd_in[342], \gcm_cmd_in.key1 [243]);
tran (gcm_cmd_in[341], \gcm_cmd_in.key1 [242]);
tran (gcm_cmd_in[340], \gcm_cmd_in.key1 [241]);
tran (gcm_cmd_in[339], \gcm_cmd_in.key1 [240]);
tran (gcm_cmd_in[338], \gcm_cmd_in.key1 [239]);
tran (gcm_cmd_in[337], \gcm_cmd_in.key1 [238]);
tran (gcm_cmd_in[336], \gcm_cmd_in.key1 [237]);
tran (gcm_cmd_in[335], \gcm_cmd_in.key1 [236]);
tran (gcm_cmd_in[334], \gcm_cmd_in.key1 [235]);
tran (gcm_cmd_in[333], \gcm_cmd_in.key1 [234]);
tran (gcm_cmd_in[332], \gcm_cmd_in.key1 [233]);
tran (gcm_cmd_in[331], \gcm_cmd_in.key1 [232]);
tran (gcm_cmd_in[330], \gcm_cmd_in.key1 [231]);
tran (gcm_cmd_in[329], \gcm_cmd_in.key1 [230]);
tran (gcm_cmd_in[328], \gcm_cmd_in.key1 [229]);
tran (gcm_cmd_in[327], \gcm_cmd_in.key1 [228]);
tran (gcm_cmd_in[326], \gcm_cmd_in.key1 [227]);
tran (gcm_cmd_in[325], \gcm_cmd_in.key1 [226]);
tran (gcm_cmd_in[324], \gcm_cmd_in.key1 [225]);
tran (gcm_cmd_in[323], \gcm_cmd_in.key1 [224]);
tran (gcm_cmd_in[322], \gcm_cmd_in.key1 [223]);
tran (gcm_cmd_in[321], \gcm_cmd_in.key1 [222]);
tran (gcm_cmd_in[320], \gcm_cmd_in.key1 [221]);
tran (gcm_cmd_in[319], \gcm_cmd_in.key1 [220]);
tran (gcm_cmd_in[318], \gcm_cmd_in.key1 [219]);
tran (gcm_cmd_in[317], \gcm_cmd_in.key1 [218]);
tran (gcm_cmd_in[316], \gcm_cmd_in.key1 [217]);
tran (gcm_cmd_in[315], \gcm_cmd_in.key1 [216]);
tran (gcm_cmd_in[314], \gcm_cmd_in.key1 [215]);
tran (gcm_cmd_in[313], \gcm_cmd_in.key1 [214]);
tran (gcm_cmd_in[312], \gcm_cmd_in.key1 [213]);
tran (gcm_cmd_in[311], \gcm_cmd_in.key1 [212]);
tran (gcm_cmd_in[310], \gcm_cmd_in.key1 [211]);
tran (gcm_cmd_in[309], \gcm_cmd_in.key1 [210]);
tran (gcm_cmd_in[308], \gcm_cmd_in.key1 [209]);
tran (gcm_cmd_in[307], \gcm_cmd_in.key1 [208]);
tran (gcm_cmd_in[306], \gcm_cmd_in.key1 [207]);
tran (gcm_cmd_in[305], \gcm_cmd_in.key1 [206]);
tran (gcm_cmd_in[304], \gcm_cmd_in.key1 [205]);
tran (gcm_cmd_in[303], \gcm_cmd_in.key1 [204]);
tran (gcm_cmd_in[302], \gcm_cmd_in.key1 [203]);
tran (gcm_cmd_in[301], \gcm_cmd_in.key1 [202]);
tran (gcm_cmd_in[300], \gcm_cmd_in.key1 [201]);
tran (gcm_cmd_in[299], \gcm_cmd_in.key1 [200]);
tran (gcm_cmd_in[298], \gcm_cmd_in.key1 [199]);
tran (gcm_cmd_in[297], \gcm_cmd_in.key1 [198]);
tran (gcm_cmd_in[296], \gcm_cmd_in.key1 [197]);
tran (gcm_cmd_in[295], \gcm_cmd_in.key1 [196]);
tran (gcm_cmd_in[294], \gcm_cmd_in.key1 [195]);
tran (gcm_cmd_in[293], \gcm_cmd_in.key1 [194]);
tran (gcm_cmd_in[292], \gcm_cmd_in.key1 [193]);
tran (gcm_cmd_in[291], \gcm_cmd_in.key1 [192]);
tran (gcm_cmd_in[290], \gcm_cmd_in.key1 [191]);
tran (gcm_cmd_in[289], \gcm_cmd_in.key1 [190]);
tran (gcm_cmd_in[288], \gcm_cmd_in.key1 [189]);
tran (gcm_cmd_in[287], \gcm_cmd_in.key1 [188]);
tran (gcm_cmd_in[286], \gcm_cmd_in.key1 [187]);
tran (gcm_cmd_in[285], \gcm_cmd_in.key1 [186]);
tran (gcm_cmd_in[284], \gcm_cmd_in.key1 [185]);
tran (gcm_cmd_in[283], \gcm_cmd_in.key1 [184]);
tran (gcm_cmd_in[282], \gcm_cmd_in.key1 [183]);
tran (gcm_cmd_in[281], \gcm_cmd_in.key1 [182]);
tran (gcm_cmd_in[280], \gcm_cmd_in.key1 [181]);
tran (gcm_cmd_in[279], \gcm_cmd_in.key1 [180]);
tran (gcm_cmd_in[278], \gcm_cmd_in.key1 [179]);
tran (gcm_cmd_in[277], \gcm_cmd_in.key1 [178]);
tran (gcm_cmd_in[276], \gcm_cmd_in.key1 [177]);
tran (gcm_cmd_in[275], \gcm_cmd_in.key1 [176]);
tran (gcm_cmd_in[274], \gcm_cmd_in.key1 [175]);
tran (gcm_cmd_in[273], \gcm_cmd_in.key1 [174]);
tran (gcm_cmd_in[272], \gcm_cmd_in.key1 [173]);
tran (gcm_cmd_in[271], \gcm_cmd_in.key1 [172]);
tran (gcm_cmd_in[270], \gcm_cmd_in.key1 [171]);
tran (gcm_cmd_in[269], \gcm_cmd_in.key1 [170]);
tran (gcm_cmd_in[268], \gcm_cmd_in.key1 [169]);
tran (gcm_cmd_in[267], \gcm_cmd_in.key1 [168]);
tran (gcm_cmd_in[266], \gcm_cmd_in.key1 [167]);
tran (gcm_cmd_in[265], \gcm_cmd_in.key1 [166]);
tran (gcm_cmd_in[264], \gcm_cmd_in.key1 [165]);
tran (gcm_cmd_in[263], \gcm_cmd_in.key1 [164]);
tran (gcm_cmd_in[262], \gcm_cmd_in.key1 [163]);
tran (gcm_cmd_in[261], \gcm_cmd_in.key1 [162]);
tran (gcm_cmd_in[260], \gcm_cmd_in.key1 [161]);
tran (gcm_cmd_in[259], \gcm_cmd_in.key1 [160]);
tran (gcm_cmd_in[258], \gcm_cmd_in.key1 [159]);
tran (gcm_cmd_in[257], \gcm_cmd_in.key1 [158]);
tran (gcm_cmd_in[256], \gcm_cmd_in.key1 [157]);
tran (gcm_cmd_in[255], \gcm_cmd_in.key1 [156]);
tran (gcm_cmd_in[254], \gcm_cmd_in.key1 [155]);
tran (gcm_cmd_in[253], \gcm_cmd_in.key1 [154]);
tran (gcm_cmd_in[252], \gcm_cmd_in.key1 [153]);
tran (gcm_cmd_in[251], \gcm_cmd_in.key1 [152]);
tran (gcm_cmd_in[250], \gcm_cmd_in.key1 [151]);
tran (gcm_cmd_in[249], \gcm_cmd_in.key1 [150]);
tran (gcm_cmd_in[248], \gcm_cmd_in.key1 [149]);
tran (gcm_cmd_in[247], \gcm_cmd_in.key1 [148]);
tran (gcm_cmd_in[246], \gcm_cmd_in.key1 [147]);
tran (gcm_cmd_in[245], \gcm_cmd_in.key1 [146]);
tran (gcm_cmd_in[244], \gcm_cmd_in.key1 [145]);
tran (gcm_cmd_in[243], \gcm_cmd_in.key1 [144]);
tran (gcm_cmd_in[242], \gcm_cmd_in.key1 [143]);
tran (gcm_cmd_in[241], \gcm_cmd_in.key1 [142]);
tran (gcm_cmd_in[240], \gcm_cmd_in.key1 [141]);
tran (gcm_cmd_in[239], \gcm_cmd_in.key1 [140]);
tran (gcm_cmd_in[238], \gcm_cmd_in.key1 [139]);
tran (gcm_cmd_in[237], \gcm_cmd_in.key1 [138]);
tran (gcm_cmd_in[236], \gcm_cmd_in.key1 [137]);
tran (gcm_cmd_in[235], \gcm_cmd_in.key1 [136]);
tran (gcm_cmd_in[234], \gcm_cmd_in.key1 [135]);
tran (gcm_cmd_in[233], \gcm_cmd_in.key1 [134]);
tran (gcm_cmd_in[232], \gcm_cmd_in.key1 [133]);
tran (gcm_cmd_in[231], \gcm_cmd_in.key1 [132]);
tran (gcm_cmd_in[230], \gcm_cmd_in.key1 [131]);
tran (gcm_cmd_in[229], \gcm_cmd_in.key1 [130]);
tran (gcm_cmd_in[228], \gcm_cmd_in.key1 [129]);
tran (gcm_cmd_in[227], \gcm_cmd_in.key1 [128]);
tran (gcm_cmd_in[226], \gcm_cmd_in.key1 [127]);
tran (gcm_cmd_in[225], \gcm_cmd_in.key1 [126]);
tran (gcm_cmd_in[224], \gcm_cmd_in.key1 [125]);
tran (gcm_cmd_in[223], \gcm_cmd_in.key1 [124]);
tran (gcm_cmd_in[222], \gcm_cmd_in.key1 [123]);
tran (gcm_cmd_in[221], \gcm_cmd_in.key1 [122]);
tran (gcm_cmd_in[220], \gcm_cmd_in.key1 [121]);
tran (gcm_cmd_in[219], \gcm_cmd_in.key1 [120]);
tran (gcm_cmd_in[218], \gcm_cmd_in.key1 [119]);
tran (gcm_cmd_in[217], \gcm_cmd_in.key1 [118]);
tran (gcm_cmd_in[216], \gcm_cmd_in.key1 [117]);
tran (gcm_cmd_in[215], \gcm_cmd_in.key1 [116]);
tran (gcm_cmd_in[214], \gcm_cmd_in.key1 [115]);
tran (gcm_cmd_in[213], \gcm_cmd_in.key1 [114]);
tran (gcm_cmd_in[212], \gcm_cmd_in.key1 [113]);
tran (gcm_cmd_in[211], \gcm_cmd_in.key1 [112]);
tran (gcm_cmd_in[210], \gcm_cmd_in.key1 [111]);
tran (gcm_cmd_in[209], \gcm_cmd_in.key1 [110]);
tran (gcm_cmd_in[208], \gcm_cmd_in.key1 [109]);
tran (gcm_cmd_in[207], \gcm_cmd_in.key1 [108]);
tran (gcm_cmd_in[206], \gcm_cmd_in.key1 [107]);
tran (gcm_cmd_in[205], \gcm_cmd_in.key1 [106]);
tran (gcm_cmd_in[204], \gcm_cmd_in.key1 [105]);
tran (gcm_cmd_in[203], \gcm_cmd_in.key1 [104]);
tran (gcm_cmd_in[202], \gcm_cmd_in.key1 [103]);
tran (gcm_cmd_in[201], \gcm_cmd_in.key1 [102]);
tran (gcm_cmd_in[200], \gcm_cmd_in.key1 [101]);
tran (gcm_cmd_in[199], \gcm_cmd_in.key1 [100]);
tran (gcm_cmd_in[198], \gcm_cmd_in.key1 [99]);
tran (gcm_cmd_in[197], \gcm_cmd_in.key1 [98]);
tran (gcm_cmd_in[196], \gcm_cmd_in.key1 [97]);
tran (gcm_cmd_in[195], \gcm_cmd_in.key1 [96]);
tran (gcm_cmd_in[194], \gcm_cmd_in.key1 [95]);
tran (gcm_cmd_in[193], \gcm_cmd_in.key1 [94]);
tran (gcm_cmd_in[192], \gcm_cmd_in.key1 [93]);
tran (gcm_cmd_in[191], \gcm_cmd_in.key1 [92]);
tran (gcm_cmd_in[190], \gcm_cmd_in.key1 [91]);
tran (gcm_cmd_in[189], \gcm_cmd_in.key1 [90]);
tran (gcm_cmd_in[188], \gcm_cmd_in.key1 [89]);
tran (gcm_cmd_in[187], \gcm_cmd_in.key1 [88]);
tran (gcm_cmd_in[186], \gcm_cmd_in.key1 [87]);
tran (gcm_cmd_in[185], \gcm_cmd_in.key1 [86]);
tran (gcm_cmd_in[184], \gcm_cmd_in.key1 [85]);
tran (gcm_cmd_in[183], \gcm_cmd_in.key1 [84]);
tran (gcm_cmd_in[182], \gcm_cmd_in.key1 [83]);
tran (gcm_cmd_in[181], \gcm_cmd_in.key1 [82]);
tran (gcm_cmd_in[180], \gcm_cmd_in.key1 [81]);
tran (gcm_cmd_in[179], \gcm_cmd_in.key1 [80]);
tran (gcm_cmd_in[178], \gcm_cmd_in.key1 [79]);
tran (gcm_cmd_in[177], \gcm_cmd_in.key1 [78]);
tran (gcm_cmd_in[176], \gcm_cmd_in.key1 [77]);
tran (gcm_cmd_in[175], \gcm_cmd_in.key1 [76]);
tran (gcm_cmd_in[174], \gcm_cmd_in.key1 [75]);
tran (gcm_cmd_in[173], \gcm_cmd_in.key1 [74]);
tran (gcm_cmd_in[172], \gcm_cmd_in.key1 [73]);
tran (gcm_cmd_in[171], \gcm_cmd_in.key1 [72]);
tran (gcm_cmd_in[170], \gcm_cmd_in.key1 [71]);
tran (gcm_cmd_in[169], \gcm_cmd_in.key1 [70]);
tran (gcm_cmd_in[168], \gcm_cmd_in.key1 [69]);
tran (gcm_cmd_in[167], \gcm_cmd_in.key1 [68]);
tran (gcm_cmd_in[166], \gcm_cmd_in.key1 [67]);
tran (gcm_cmd_in[165], \gcm_cmd_in.key1 [66]);
tran (gcm_cmd_in[164], \gcm_cmd_in.key1 [65]);
tran (gcm_cmd_in[163], \gcm_cmd_in.key1 [64]);
tran (gcm_cmd_in[162], \gcm_cmd_in.key1 [63]);
tran (gcm_cmd_in[161], \gcm_cmd_in.key1 [62]);
tran (gcm_cmd_in[160], \gcm_cmd_in.key1 [61]);
tran (gcm_cmd_in[159], \gcm_cmd_in.key1 [60]);
tran (gcm_cmd_in[158], \gcm_cmd_in.key1 [59]);
tran (gcm_cmd_in[157], \gcm_cmd_in.key1 [58]);
tran (gcm_cmd_in[156], \gcm_cmd_in.key1 [57]);
tran (gcm_cmd_in[155], \gcm_cmd_in.key1 [56]);
tran (gcm_cmd_in[154], \gcm_cmd_in.key1 [55]);
tran (gcm_cmd_in[153], \gcm_cmd_in.key1 [54]);
tran (gcm_cmd_in[152], \gcm_cmd_in.key1 [53]);
tran (gcm_cmd_in[151], \gcm_cmd_in.key1 [52]);
tran (gcm_cmd_in[150], \gcm_cmd_in.key1 [51]);
tran (gcm_cmd_in[149], \gcm_cmd_in.key1 [50]);
tran (gcm_cmd_in[148], \gcm_cmd_in.key1 [49]);
tran (gcm_cmd_in[147], \gcm_cmd_in.key1 [48]);
tran (gcm_cmd_in[146], \gcm_cmd_in.key1 [47]);
tran (gcm_cmd_in[145], \gcm_cmd_in.key1 [46]);
tran (gcm_cmd_in[144], \gcm_cmd_in.key1 [45]);
tran (gcm_cmd_in[143], \gcm_cmd_in.key1 [44]);
tran (gcm_cmd_in[142], \gcm_cmd_in.key1 [43]);
tran (gcm_cmd_in[141], \gcm_cmd_in.key1 [42]);
tran (gcm_cmd_in[140], \gcm_cmd_in.key1 [41]);
tran (gcm_cmd_in[139], \gcm_cmd_in.key1 [40]);
tran (gcm_cmd_in[138], \gcm_cmd_in.key1 [39]);
tran (gcm_cmd_in[137], \gcm_cmd_in.key1 [38]);
tran (gcm_cmd_in[136], \gcm_cmd_in.key1 [37]);
tran (gcm_cmd_in[135], \gcm_cmd_in.key1 [36]);
tran (gcm_cmd_in[134], \gcm_cmd_in.key1 [35]);
tran (gcm_cmd_in[133], \gcm_cmd_in.key1 [34]);
tran (gcm_cmd_in[132], \gcm_cmd_in.key1 [33]);
tran (gcm_cmd_in[131], \gcm_cmd_in.key1 [32]);
tran (gcm_cmd_in[130], \gcm_cmd_in.key1 [31]);
tran (gcm_cmd_in[129], \gcm_cmd_in.key1 [30]);
tran (gcm_cmd_in[128], \gcm_cmd_in.key1 [29]);
tran (gcm_cmd_in[127], \gcm_cmd_in.key1 [28]);
tran (gcm_cmd_in[126], \gcm_cmd_in.key1 [27]);
tran (gcm_cmd_in[125], \gcm_cmd_in.key1 [26]);
tran (gcm_cmd_in[124], \gcm_cmd_in.key1 [25]);
tran (gcm_cmd_in[123], \gcm_cmd_in.key1 [24]);
tran (gcm_cmd_in[122], \gcm_cmd_in.key1 [23]);
tran (gcm_cmd_in[121], \gcm_cmd_in.key1 [22]);
tran (gcm_cmd_in[120], \gcm_cmd_in.key1 [21]);
tran (gcm_cmd_in[119], \gcm_cmd_in.key1 [20]);
tran (gcm_cmd_in[118], \gcm_cmd_in.key1 [19]);
tran (gcm_cmd_in[117], \gcm_cmd_in.key1 [18]);
tran (gcm_cmd_in[116], \gcm_cmd_in.key1 [17]);
tran (gcm_cmd_in[115], \gcm_cmd_in.key1 [16]);
tran (gcm_cmd_in[114], \gcm_cmd_in.key1 [15]);
tran (gcm_cmd_in[113], \gcm_cmd_in.key1 [14]);
tran (gcm_cmd_in[112], \gcm_cmd_in.key1 [13]);
tran (gcm_cmd_in[111], \gcm_cmd_in.key1 [12]);
tran (gcm_cmd_in[110], \gcm_cmd_in.key1 [11]);
tran (gcm_cmd_in[109], \gcm_cmd_in.key1 [10]);
tran (gcm_cmd_in[108], \gcm_cmd_in.key1 [9]);
tran (gcm_cmd_in[107], \gcm_cmd_in.key1 [8]);
tran (gcm_cmd_in[106], \gcm_cmd_in.key1 [7]);
tran (gcm_cmd_in[105], \gcm_cmd_in.key1 [6]);
tran (gcm_cmd_in[104], \gcm_cmd_in.key1 [5]);
tran (gcm_cmd_in[103], \gcm_cmd_in.key1 [4]);
tran (gcm_cmd_in[102], \gcm_cmd_in.key1 [3]);
tran (gcm_cmd_in[101], \gcm_cmd_in.key1 [2]);
tran (gcm_cmd_in[100], \gcm_cmd_in.key1 [1]);
tran (gcm_cmd_in[99], \gcm_cmd_in.key1 [0]);
tran (gcm_cmd_in[98], \gcm_cmd_in.iv [95]);
tran (gcm_cmd_in[97], \gcm_cmd_in.iv [94]);
tran (gcm_cmd_in[96], \gcm_cmd_in.iv [93]);
tran (gcm_cmd_in[95], \gcm_cmd_in.iv [92]);
tran (gcm_cmd_in[94], \gcm_cmd_in.iv [91]);
tran (gcm_cmd_in[93], \gcm_cmd_in.iv [90]);
tran (gcm_cmd_in[92], \gcm_cmd_in.iv [89]);
tran (gcm_cmd_in[91], \gcm_cmd_in.iv [88]);
tran (gcm_cmd_in[90], \gcm_cmd_in.iv [87]);
tran (gcm_cmd_in[89], \gcm_cmd_in.iv [86]);
tran (gcm_cmd_in[88], \gcm_cmd_in.iv [85]);
tran (gcm_cmd_in[87], \gcm_cmd_in.iv [84]);
tran (gcm_cmd_in[86], \gcm_cmd_in.iv [83]);
tran (gcm_cmd_in[85], \gcm_cmd_in.iv [82]);
tran (gcm_cmd_in[84], \gcm_cmd_in.iv [81]);
tran (gcm_cmd_in[83], \gcm_cmd_in.iv [80]);
tran (gcm_cmd_in[82], \gcm_cmd_in.iv [79]);
tran (gcm_cmd_in[81], \gcm_cmd_in.iv [78]);
tran (gcm_cmd_in[80], \gcm_cmd_in.iv [77]);
tran (gcm_cmd_in[79], \gcm_cmd_in.iv [76]);
tran (gcm_cmd_in[78], \gcm_cmd_in.iv [75]);
tran (gcm_cmd_in[77], \gcm_cmd_in.iv [74]);
tran (gcm_cmd_in[76], \gcm_cmd_in.iv [73]);
tran (gcm_cmd_in[75], \gcm_cmd_in.iv [72]);
tran (gcm_cmd_in[74], \gcm_cmd_in.iv [71]);
tran (gcm_cmd_in[73], \gcm_cmd_in.iv [70]);
tran (gcm_cmd_in[72], \gcm_cmd_in.iv [69]);
tran (gcm_cmd_in[71], \gcm_cmd_in.iv [68]);
tran (gcm_cmd_in[70], \gcm_cmd_in.iv [67]);
tran (gcm_cmd_in[69], \gcm_cmd_in.iv [66]);
tran (gcm_cmd_in[68], \gcm_cmd_in.iv [65]);
tran (gcm_cmd_in[67], \gcm_cmd_in.iv [64]);
tran (gcm_cmd_in[66], \gcm_cmd_in.iv [63]);
tran (gcm_cmd_in[65], \gcm_cmd_in.iv [62]);
tran (gcm_cmd_in[64], \gcm_cmd_in.iv [61]);
tran (gcm_cmd_in[63], \gcm_cmd_in.iv [60]);
tran (gcm_cmd_in[62], \gcm_cmd_in.iv [59]);
tran (gcm_cmd_in[61], \gcm_cmd_in.iv [58]);
tran (gcm_cmd_in[60], \gcm_cmd_in.iv [57]);
tran (gcm_cmd_in[59], \gcm_cmd_in.iv [56]);
tran (gcm_cmd_in[58], \gcm_cmd_in.iv [55]);
tran (gcm_cmd_in[57], \gcm_cmd_in.iv [54]);
tran (gcm_cmd_in[56], \gcm_cmd_in.iv [53]);
tran (gcm_cmd_in[55], \gcm_cmd_in.iv [52]);
tran (gcm_cmd_in[54], \gcm_cmd_in.iv [51]);
tran (gcm_cmd_in[53], \gcm_cmd_in.iv [50]);
tran (gcm_cmd_in[52], \gcm_cmd_in.iv [49]);
tran (gcm_cmd_in[51], \gcm_cmd_in.iv [48]);
tran (gcm_cmd_in[50], \gcm_cmd_in.iv [47]);
tran (gcm_cmd_in[49], \gcm_cmd_in.iv [46]);
tran (gcm_cmd_in[48], \gcm_cmd_in.iv [45]);
tran (gcm_cmd_in[47], \gcm_cmd_in.iv [44]);
tran (gcm_cmd_in[46], \gcm_cmd_in.iv [43]);
tran (gcm_cmd_in[45], \gcm_cmd_in.iv [42]);
tran (gcm_cmd_in[44], \gcm_cmd_in.iv [41]);
tran (gcm_cmd_in[43], \gcm_cmd_in.iv [40]);
tran (gcm_cmd_in[42], \gcm_cmd_in.iv [39]);
tran (gcm_cmd_in[41], \gcm_cmd_in.iv [38]);
tran (gcm_cmd_in[40], \gcm_cmd_in.iv [37]);
tran (gcm_cmd_in[39], \gcm_cmd_in.iv [36]);
tran (gcm_cmd_in[38], \gcm_cmd_in.iv [35]);
tran (gcm_cmd_in[37], \gcm_cmd_in.iv [34]);
tran (gcm_cmd_in[36], \gcm_cmd_in.iv [33]);
tran (gcm_cmd_in[35], \gcm_cmd_in.iv [32]);
tran (gcm_cmd_in[34], \gcm_cmd_in.iv [31]);
tran (gcm_cmd_in[33], \gcm_cmd_in.iv [30]);
tran (gcm_cmd_in[32], \gcm_cmd_in.iv [29]);
tran (gcm_cmd_in[31], \gcm_cmd_in.iv [28]);
tran (gcm_cmd_in[30], \gcm_cmd_in.iv [27]);
tran (gcm_cmd_in[29], \gcm_cmd_in.iv [26]);
tran (gcm_cmd_in[28], \gcm_cmd_in.iv [25]);
tran (gcm_cmd_in[27], \gcm_cmd_in.iv [24]);
tran (gcm_cmd_in[26], \gcm_cmd_in.iv [23]);
tran (gcm_cmd_in[25], \gcm_cmd_in.iv [22]);
tran (gcm_cmd_in[24], \gcm_cmd_in.iv [21]);
tran (gcm_cmd_in[23], \gcm_cmd_in.iv [20]);
tran (gcm_cmd_in[22], \gcm_cmd_in.iv [19]);
tran (gcm_cmd_in[21], \gcm_cmd_in.iv [18]);
tran (gcm_cmd_in[20], \gcm_cmd_in.iv [17]);
tran (gcm_cmd_in[19], \gcm_cmd_in.iv [16]);
tran (gcm_cmd_in[18], \gcm_cmd_in.iv [15]);
tran (gcm_cmd_in[17], \gcm_cmd_in.iv [14]);
tran (gcm_cmd_in[16], \gcm_cmd_in.iv [13]);
tran (gcm_cmd_in[15], \gcm_cmd_in.iv [12]);
tran (gcm_cmd_in[14], \gcm_cmd_in.iv [11]);
tran (gcm_cmd_in[13], \gcm_cmd_in.iv [10]);
tran (gcm_cmd_in[12], \gcm_cmd_in.iv [9]);
tran (gcm_cmd_in[11], \gcm_cmd_in.iv [8]);
tran (gcm_cmd_in[10], \gcm_cmd_in.iv [7]);
tran (gcm_cmd_in[9], \gcm_cmd_in.iv [6]);
tran (gcm_cmd_in[8], \gcm_cmd_in.iv [5]);
tran (gcm_cmd_in[7], \gcm_cmd_in.iv [4]);
tran (gcm_cmd_in[6], \gcm_cmd_in.iv [3]);
tran (gcm_cmd_in[5], \gcm_cmd_in.iv [2]);
tran (gcm_cmd_in[4], \gcm_cmd_in.iv [1]);
tran (gcm_cmd_in[3], \gcm_cmd_in.iv [0]);
tran (gcm_cmd_in[2], \gcm_cmd_in.op [2]);
tran (gcm_cmd_in[1], \gcm_cmd_in.op [1]);
tran (gcm_cmd_in[0], \gcm_cmd_in.op [0]);
tran (keyfilter_cmd_in[0], \keyfilter_cmd_in.combo_mode [0]);
tran (kdfstream_cmd_in[262], \kdfstream_cmd_in.combo_mode [0]);
tran (kdfstream_cmd_in[261], \kdfstream_cmd_in.skip [0]);
tran (kdfstream_cmd_in[260], \kdfstream_cmd_in.guid [255]);
tran (kdfstream_cmd_in[259], \kdfstream_cmd_in.guid [254]);
tran (kdfstream_cmd_in[258], \kdfstream_cmd_in.guid [253]);
tran (kdfstream_cmd_in[257], \kdfstream_cmd_in.guid [252]);
tran (kdfstream_cmd_in[256], \kdfstream_cmd_in.guid [251]);
tran (kdfstream_cmd_in[255], \kdfstream_cmd_in.guid [250]);
tran (kdfstream_cmd_in[254], \kdfstream_cmd_in.guid [249]);
tran (kdfstream_cmd_in[253], \kdfstream_cmd_in.guid [248]);
tran (kdfstream_cmd_in[252], \kdfstream_cmd_in.guid [247]);
tran (kdfstream_cmd_in[251], \kdfstream_cmd_in.guid [246]);
tran (kdfstream_cmd_in[250], \kdfstream_cmd_in.guid [245]);
tran (kdfstream_cmd_in[249], \kdfstream_cmd_in.guid [244]);
tran (kdfstream_cmd_in[248], \kdfstream_cmd_in.guid [243]);
tran (kdfstream_cmd_in[247], \kdfstream_cmd_in.guid [242]);
tran (kdfstream_cmd_in[246], \kdfstream_cmd_in.guid [241]);
tran (kdfstream_cmd_in[245], \kdfstream_cmd_in.guid [240]);
tran (kdfstream_cmd_in[244], \kdfstream_cmd_in.guid [239]);
tran (kdfstream_cmd_in[243], \kdfstream_cmd_in.guid [238]);
tran (kdfstream_cmd_in[242], \kdfstream_cmd_in.guid [237]);
tran (kdfstream_cmd_in[241], \kdfstream_cmd_in.guid [236]);
tran (kdfstream_cmd_in[240], \kdfstream_cmd_in.guid [235]);
tran (kdfstream_cmd_in[239], \kdfstream_cmd_in.guid [234]);
tran (kdfstream_cmd_in[238], \kdfstream_cmd_in.guid [233]);
tran (kdfstream_cmd_in[237], \kdfstream_cmd_in.guid [232]);
tran (kdfstream_cmd_in[236], \kdfstream_cmd_in.guid [231]);
tran (kdfstream_cmd_in[235], \kdfstream_cmd_in.guid [230]);
tran (kdfstream_cmd_in[234], \kdfstream_cmd_in.guid [229]);
tran (kdfstream_cmd_in[233], \kdfstream_cmd_in.guid [228]);
tran (kdfstream_cmd_in[232], \kdfstream_cmd_in.guid [227]);
tran (kdfstream_cmd_in[231], \kdfstream_cmd_in.guid [226]);
tran (kdfstream_cmd_in[230], \kdfstream_cmd_in.guid [225]);
tran (kdfstream_cmd_in[229], \kdfstream_cmd_in.guid [224]);
tran (kdfstream_cmd_in[228], \kdfstream_cmd_in.guid [223]);
tran (kdfstream_cmd_in[227], \kdfstream_cmd_in.guid [222]);
tran (kdfstream_cmd_in[226], \kdfstream_cmd_in.guid [221]);
tran (kdfstream_cmd_in[225], \kdfstream_cmd_in.guid [220]);
tran (kdfstream_cmd_in[224], \kdfstream_cmd_in.guid [219]);
tran (kdfstream_cmd_in[223], \kdfstream_cmd_in.guid [218]);
tran (kdfstream_cmd_in[222], \kdfstream_cmd_in.guid [217]);
tran (kdfstream_cmd_in[221], \kdfstream_cmd_in.guid [216]);
tran (kdfstream_cmd_in[220], \kdfstream_cmd_in.guid [215]);
tran (kdfstream_cmd_in[219], \kdfstream_cmd_in.guid [214]);
tran (kdfstream_cmd_in[218], \kdfstream_cmd_in.guid [213]);
tran (kdfstream_cmd_in[217], \kdfstream_cmd_in.guid [212]);
tran (kdfstream_cmd_in[216], \kdfstream_cmd_in.guid [211]);
tran (kdfstream_cmd_in[215], \kdfstream_cmd_in.guid [210]);
tran (kdfstream_cmd_in[214], \kdfstream_cmd_in.guid [209]);
tran (kdfstream_cmd_in[213], \kdfstream_cmd_in.guid [208]);
tran (kdfstream_cmd_in[212], \kdfstream_cmd_in.guid [207]);
tran (kdfstream_cmd_in[211], \kdfstream_cmd_in.guid [206]);
tran (kdfstream_cmd_in[210], \kdfstream_cmd_in.guid [205]);
tran (kdfstream_cmd_in[209], \kdfstream_cmd_in.guid [204]);
tran (kdfstream_cmd_in[208], \kdfstream_cmd_in.guid [203]);
tran (kdfstream_cmd_in[207], \kdfstream_cmd_in.guid [202]);
tran (kdfstream_cmd_in[206], \kdfstream_cmd_in.guid [201]);
tran (kdfstream_cmd_in[205], \kdfstream_cmd_in.guid [200]);
tran (kdfstream_cmd_in[204], \kdfstream_cmd_in.guid [199]);
tran (kdfstream_cmd_in[203], \kdfstream_cmd_in.guid [198]);
tran (kdfstream_cmd_in[202], \kdfstream_cmd_in.guid [197]);
tran (kdfstream_cmd_in[201], \kdfstream_cmd_in.guid [196]);
tran (kdfstream_cmd_in[200], \kdfstream_cmd_in.guid [195]);
tran (kdfstream_cmd_in[199], \kdfstream_cmd_in.guid [194]);
tran (kdfstream_cmd_in[198], \kdfstream_cmd_in.guid [193]);
tran (kdfstream_cmd_in[197], \kdfstream_cmd_in.guid [192]);
tran (kdfstream_cmd_in[196], \kdfstream_cmd_in.guid [191]);
tran (kdfstream_cmd_in[195], \kdfstream_cmd_in.guid [190]);
tran (kdfstream_cmd_in[194], \kdfstream_cmd_in.guid [189]);
tran (kdfstream_cmd_in[193], \kdfstream_cmd_in.guid [188]);
tran (kdfstream_cmd_in[192], \kdfstream_cmd_in.guid [187]);
tran (kdfstream_cmd_in[191], \kdfstream_cmd_in.guid [186]);
tran (kdfstream_cmd_in[190], \kdfstream_cmd_in.guid [185]);
tran (kdfstream_cmd_in[189], \kdfstream_cmd_in.guid [184]);
tran (kdfstream_cmd_in[188], \kdfstream_cmd_in.guid [183]);
tran (kdfstream_cmd_in[187], \kdfstream_cmd_in.guid [182]);
tran (kdfstream_cmd_in[186], \kdfstream_cmd_in.guid [181]);
tran (kdfstream_cmd_in[185], \kdfstream_cmd_in.guid [180]);
tran (kdfstream_cmd_in[184], \kdfstream_cmd_in.guid [179]);
tran (kdfstream_cmd_in[183], \kdfstream_cmd_in.guid [178]);
tran (kdfstream_cmd_in[182], \kdfstream_cmd_in.guid [177]);
tran (kdfstream_cmd_in[181], \kdfstream_cmd_in.guid [176]);
tran (kdfstream_cmd_in[180], \kdfstream_cmd_in.guid [175]);
tran (kdfstream_cmd_in[179], \kdfstream_cmd_in.guid [174]);
tran (kdfstream_cmd_in[178], \kdfstream_cmd_in.guid [173]);
tran (kdfstream_cmd_in[177], \kdfstream_cmd_in.guid [172]);
tran (kdfstream_cmd_in[176], \kdfstream_cmd_in.guid [171]);
tran (kdfstream_cmd_in[175], \kdfstream_cmd_in.guid [170]);
tran (kdfstream_cmd_in[174], \kdfstream_cmd_in.guid [169]);
tran (kdfstream_cmd_in[173], \kdfstream_cmd_in.guid [168]);
tran (kdfstream_cmd_in[172], \kdfstream_cmd_in.guid [167]);
tran (kdfstream_cmd_in[171], \kdfstream_cmd_in.guid [166]);
tran (kdfstream_cmd_in[170], \kdfstream_cmd_in.guid [165]);
tran (kdfstream_cmd_in[169], \kdfstream_cmd_in.guid [164]);
tran (kdfstream_cmd_in[168], \kdfstream_cmd_in.guid [163]);
tran (kdfstream_cmd_in[167], \kdfstream_cmd_in.guid [162]);
tran (kdfstream_cmd_in[166], \kdfstream_cmd_in.guid [161]);
tran (kdfstream_cmd_in[165], \kdfstream_cmd_in.guid [160]);
tran (kdfstream_cmd_in[164], \kdfstream_cmd_in.guid [159]);
tran (kdfstream_cmd_in[163], \kdfstream_cmd_in.guid [158]);
tran (kdfstream_cmd_in[162], \kdfstream_cmd_in.guid [157]);
tran (kdfstream_cmd_in[161], \kdfstream_cmd_in.guid [156]);
tran (kdfstream_cmd_in[160], \kdfstream_cmd_in.guid [155]);
tran (kdfstream_cmd_in[159], \kdfstream_cmd_in.guid [154]);
tran (kdfstream_cmd_in[158], \kdfstream_cmd_in.guid [153]);
tran (kdfstream_cmd_in[157], \kdfstream_cmd_in.guid [152]);
tran (kdfstream_cmd_in[156], \kdfstream_cmd_in.guid [151]);
tran (kdfstream_cmd_in[155], \kdfstream_cmd_in.guid [150]);
tran (kdfstream_cmd_in[154], \kdfstream_cmd_in.guid [149]);
tran (kdfstream_cmd_in[153], \kdfstream_cmd_in.guid [148]);
tran (kdfstream_cmd_in[152], \kdfstream_cmd_in.guid [147]);
tran (kdfstream_cmd_in[151], \kdfstream_cmd_in.guid [146]);
tran (kdfstream_cmd_in[150], \kdfstream_cmd_in.guid [145]);
tran (kdfstream_cmd_in[149], \kdfstream_cmd_in.guid [144]);
tran (kdfstream_cmd_in[148], \kdfstream_cmd_in.guid [143]);
tran (kdfstream_cmd_in[147], \kdfstream_cmd_in.guid [142]);
tran (kdfstream_cmd_in[146], \kdfstream_cmd_in.guid [141]);
tran (kdfstream_cmd_in[145], \kdfstream_cmd_in.guid [140]);
tran (kdfstream_cmd_in[144], \kdfstream_cmd_in.guid [139]);
tran (kdfstream_cmd_in[143], \kdfstream_cmd_in.guid [138]);
tran (kdfstream_cmd_in[142], \kdfstream_cmd_in.guid [137]);
tran (kdfstream_cmd_in[141], \kdfstream_cmd_in.guid [136]);
tran (kdfstream_cmd_in[140], \kdfstream_cmd_in.guid [135]);
tran (kdfstream_cmd_in[139], \kdfstream_cmd_in.guid [134]);
tran (kdfstream_cmd_in[138], \kdfstream_cmd_in.guid [133]);
tran (kdfstream_cmd_in[137], \kdfstream_cmd_in.guid [132]);
tran (kdfstream_cmd_in[136], \kdfstream_cmd_in.guid [131]);
tran (kdfstream_cmd_in[135], \kdfstream_cmd_in.guid [130]);
tran (kdfstream_cmd_in[134], \kdfstream_cmd_in.guid [129]);
tran (kdfstream_cmd_in[133], \kdfstream_cmd_in.guid [128]);
tran (kdfstream_cmd_in[132], \kdfstream_cmd_in.guid [127]);
tran (kdfstream_cmd_in[131], \kdfstream_cmd_in.guid [126]);
tran (kdfstream_cmd_in[130], \kdfstream_cmd_in.guid [125]);
tran (kdfstream_cmd_in[129], \kdfstream_cmd_in.guid [124]);
tran (kdfstream_cmd_in[128], \kdfstream_cmd_in.guid [123]);
tran (kdfstream_cmd_in[127], \kdfstream_cmd_in.guid [122]);
tran (kdfstream_cmd_in[126], \kdfstream_cmd_in.guid [121]);
tran (kdfstream_cmd_in[125], \kdfstream_cmd_in.guid [120]);
tran (kdfstream_cmd_in[124], \kdfstream_cmd_in.guid [119]);
tran (kdfstream_cmd_in[123], \kdfstream_cmd_in.guid [118]);
tran (kdfstream_cmd_in[122], \kdfstream_cmd_in.guid [117]);
tran (kdfstream_cmd_in[121], \kdfstream_cmd_in.guid [116]);
tran (kdfstream_cmd_in[120], \kdfstream_cmd_in.guid [115]);
tran (kdfstream_cmd_in[119], \kdfstream_cmd_in.guid [114]);
tran (kdfstream_cmd_in[118], \kdfstream_cmd_in.guid [113]);
tran (kdfstream_cmd_in[117], \kdfstream_cmd_in.guid [112]);
tran (kdfstream_cmd_in[116], \kdfstream_cmd_in.guid [111]);
tran (kdfstream_cmd_in[115], \kdfstream_cmd_in.guid [110]);
tran (kdfstream_cmd_in[114], \kdfstream_cmd_in.guid [109]);
tran (kdfstream_cmd_in[113], \kdfstream_cmd_in.guid [108]);
tran (kdfstream_cmd_in[112], \kdfstream_cmd_in.guid [107]);
tran (kdfstream_cmd_in[111], \kdfstream_cmd_in.guid [106]);
tran (kdfstream_cmd_in[110], \kdfstream_cmd_in.guid [105]);
tran (kdfstream_cmd_in[109], \kdfstream_cmd_in.guid [104]);
tran (kdfstream_cmd_in[108], \kdfstream_cmd_in.guid [103]);
tran (kdfstream_cmd_in[107], \kdfstream_cmd_in.guid [102]);
tran (kdfstream_cmd_in[106], \kdfstream_cmd_in.guid [101]);
tran (kdfstream_cmd_in[105], \kdfstream_cmd_in.guid [100]);
tran (kdfstream_cmd_in[104], \kdfstream_cmd_in.guid [99]);
tran (kdfstream_cmd_in[103], \kdfstream_cmd_in.guid [98]);
tran (kdfstream_cmd_in[102], \kdfstream_cmd_in.guid [97]);
tran (kdfstream_cmd_in[101], \kdfstream_cmd_in.guid [96]);
tran (kdfstream_cmd_in[100], \kdfstream_cmd_in.guid [95]);
tran (kdfstream_cmd_in[99], \kdfstream_cmd_in.guid [94]);
tran (kdfstream_cmd_in[98], \kdfstream_cmd_in.guid [93]);
tran (kdfstream_cmd_in[97], \kdfstream_cmd_in.guid [92]);
tran (kdfstream_cmd_in[96], \kdfstream_cmd_in.guid [91]);
tran (kdfstream_cmd_in[95], \kdfstream_cmd_in.guid [90]);
tran (kdfstream_cmd_in[94], \kdfstream_cmd_in.guid [89]);
tran (kdfstream_cmd_in[93], \kdfstream_cmd_in.guid [88]);
tran (kdfstream_cmd_in[92], \kdfstream_cmd_in.guid [87]);
tran (kdfstream_cmd_in[91], \kdfstream_cmd_in.guid [86]);
tran (kdfstream_cmd_in[90], \kdfstream_cmd_in.guid [85]);
tran (kdfstream_cmd_in[89], \kdfstream_cmd_in.guid [84]);
tran (kdfstream_cmd_in[88], \kdfstream_cmd_in.guid [83]);
tran (kdfstream_cmd_in[87], \kdfstream_cmd_in.guid [82]);
tran (kdfstream_cmd_in[86], \kdfstream_cmd_in.guid [81]);
tran (kdfstream_cmd_in[85], \kdfstream_cmd_in.guid [80]);
tran (kdfstream_cmd_in[84], \kdfstream_cmd_in.guid [79]);
tran (kdfstream_cmd_in[83], \kdfstream_cmd_in.guid [78]);
tran (kdfstream_cmd_in[82], \kdfstream_cmd_in.guid [77]);
tran (kdfstream_cmd_in[81], \kdfstream_cmd_in.guid [76]);
tran (kdfstream_cmd_in[80], \kdfstream_cmd_in.guid [75]);
tran (kdfstream_cmd_in[79], \kdfstream_cmd_in.guid [74]);
tran (kdfstream_cmd_in[78], \kdfstream_cmd_in.guid [73]);
tran (kdfstream_cmd_in[77], \kdfstream_cmd_in.guid [72]);
tran (kdfstream_cmd_in[76], \kdfstream_cmd_in.guid [71]);
tran (kdfstream_cmd_in[75], \kdfstream_cmd_in.guid [70]);
tran (kdfstream_cmd_in[74], \kdfstream_cmd_in.guid [69]);
tran (kdfstream_cmd_in[73], \kdfstream_cmd_in.guid [68]);
tran (kdfstream_cmd_in[72], \kdfstream_cmd_in.guid [67]);
tran (kdfstream_cmd_in[71], \kdfstream_cmd_in.guid [66]);
tran (kdfstream_cmd_in[70], \kdfstream_cmd_in.guid [65]);
tran (kdfstream_cmd_in[69], \kdfstream_cmd_in.guid [64]);
tran (kdfstream_cmd_in[68], \kdfstream_cmd_in.guid [63]);
tran (kdfstream_cmd_in[67], \kdfstream_cmd_in.guid [62]);
tran (kdfstream_cmd_in[66], \kdfstream_cmd_in.guid [61]);
tran (kdfstream_cmd_in[65], \kdfstream_cmd_in.guid [60]);
tran (kdfstream_cmd_in[64], \kdfstream_cmd_in.guid [59]);
tran (kdfstream_cmd_in[63], \kdfstream_cmd_in.guid [58]);
tran (kdfstream_cmd_in[62], \kdfstream_cmd_in.guid [57]);
tran (kdfstream_cmd_in[61], \kdfstream_cmd_in.guid [56]);
tran (kdfstream_cmd_in[60], \kdfstream_cmd_in.guid [55]);
tran (kdfstream_cmd_in[59], \kdfstream_cmd_in.guid [54]);
tran (kdfstream_cmd_in[58], \kdfstream_cmd_in.guid [53]);
tran (kdfstream_cmd_in[57], \kdfstream_cmd_in.guid [52]);
tran (kdfstream_cmd_in[56], \kdfstream_cmd_in.guid [51]);
tran (kdfstream_cmd_in[55], \kdfstream_cmd_in.guid [50]);
tran (kdfstream_cmd_in[54], \kdfstream_cmd_in.guid [49]);
tran (kdfstream_cmd_in[53], \kdfstream_cmd_in.guid [48]);
tran (kdfstream_cmd_in[52], \kdfstream_cmd_in.guid [47]);
tran (kdfstream_cmd_in[51], \kdfstream_cmd_in.guid [46]);
tran (kdfstream_cmd_in[50], \kdfstream_cmd_in.guid [45]);
tran (kdfstream_cmd_in[49], \kdfstream_cmd_in.guid [44]);
tran (kdfstream_cmd_in[48], \kdfstream_cmd_in.guid [43]);
tran (kdfstream_cmd_in[47], \kdfstream_cmd_in.guid [42]);
tran (kdfstream_cmd_in[46], \kdfstream_cmd_in.guid [41]);
tran (kdfstream_cmd_in[45], \kdfstream_cmd_in.guid [40]);
tran (kdfstream_cmd_in[44], \kdfstream_cmd_in.guid [39]);
tran (kdfstream_cmd_in[43], \kdfstream_cmd_in.guid [38]);
tran (kdfstream_cmd_in[42], \kdfstream_cmd_in.guid [37]);
tran (kdfstream_cmd_in[41], \kdfstream_cmd_in.guid [36]);
tran (kdfstream_cmd_in[40], \kdfstream_cmd_in.guid [35]);
tran (kdfstream_cmd_in[39], \kdfstream_cmd_in.guid [34]);
tran (kdfstream_cmd_in[38], \kdfstream_cmd_in.guid [33]);
tran (kdfstream_cmd_in[37], \kdfstream_cmd_in.guid [32]);
tran (kdfstream_cmd_in[36], \kdfstream_cmd_in.guid [31]);
tran (kdfstream_cmd_in[35], \kdfstream_cmd_in.guid [30]);
tran (kdfstream_cmd_in[34], \kdfstream_cmd_in.guid [29]);
tran (kdfstream_cmd_in[33], \kdfstream_cmd_in.guid [28]);
tran (kdfstream_cmd_in[32], \kdfstream_cmd_in.guid [27]);
tran (kdfstream_cmd_in[31], \kdfstream_cmd_in.guid [26]);
tran (kdfstream_cmd_in[30], \kdfstream_cmd_in.guid [25]);
tran (kdfstream_cmd_in[29], \kdfstream_cmd_in.guid [24]);
tran (kdfstream_cmd_in[28], \kdfstream_cmd_in.guid [23]);
tran (kdfstream_cmd_in[27], \kdfstream_cmd_in.guid [22]);
tran (kdfstream_cmd_in[26], \kdfstream_cmd_in.guid [21]);
tran (kdfstream_cmd_in[25], \kdfstream_cmd_in.guid [20]);
tran (kdfstream_cmd_in[24], \kdfstream_cmd_in.guid [19]);
tran (kdfstream_cmd_in[23], \kdfstream_cmd_in.guid [18]);
tran (kdfstream_cmd_in[22], \kdfstream_cmd_in.guid [17]);
tran (kdfstream_cmd_in[21], \kdfstream_cmd_in.guid [16]);
tran (kdfstream_cmd_in[20], \kdfstream_cmd_in.guid [15]);
tran (kdfstream_cmd_in[19], \kdfstream_cmd_in.guid [14]);
tran (kdfstream_cmd_in[18], \kdfstream_cmd_in.guid [13]);
tran (kdfstream_cmd_in[17], \kdfstream_cmd_in.guid [12]);
tran (kdfstream_cmd_in[16], \kdfstream_cmd_in.guid [11]);
tran (kdfstream_cmd_in[15], \kdfstream_cmd_in.guid [10]);
tran (kdfstream_cmd_in[14], \kdfstream_cmd_in.guid [9]);
tran (kdfstream_cmd_in[13], \kdfstream_cmd_in.guid [8]);
tran (kdfstream_cmd_in[12], \kdfstream_cmd_in.guid [7]);
tran (kdfstream_cmd_in[11], \kdfstream_cmd_in.guid [6]);
tran (kdfstream_cmd_in[10], \kdfstream_cmd_in.guid [5]);
tran (kdfstream_cmd_in[9], \kdfstream_cmd_in.guid [4]);
tran (kdfstream_cmd_in[8], \kdfstream_cmd_in.guid [3]);
tran (kdfstream_cmd_in[7], \kdfstream_cmd_in.guid [2]);
tran (kdfstream_cmd_in[6], \kdfstream_cmd_in.guid [1]);
tran (kdfstream_cmd_in[5], \kdfstream_cmd_in.guid [0]);
tran (kdfstream_cmd_in[4], \kdfstream_cmd_in.label_index [2]);
tran (kdfstream_cmd_in[3], \kdfstream_cmd_in.label_index [1]);
tran (kdfstream_cmd_in[2], \kdfstream_cmd_in.label_index [0]);
tran (kdfstream_cmd_in[1], \kdfstream_cmd_in.num_iter [1]);
tran (kdfstream_cmd_in[0], \kdfstream_cmd_in.num_iter [0]);
tran (kdf_cmd_in[3], \kdf_cmd_in.kdf_dek_iter [0]);
tran (kdf_cmd_in[2], \kdf_cmd_in.combo_mode [0]);
tran (kdf_cmd_in[1], \kdf_cmd_in.dek_key_op [0]);
tran (kdf_cmd_in[0], \kdf_cmd_in.dak_key_op [0]);
tran (gcm_status_data_in[0], \gcm_status_data_in.tag_mismatch [0]);
ixc_assign_106 _zz_strnp_0 ( _zy_simnet_key_tlv_ob_tlv_0_w$[0:105], 
	key_tlv_ob_tlv[105:0]);
ixc_assign_611 _zz_strnp_1 ( gcm_cmd_in[610:0], 
	_zy_simnet_gcm_cmd_in_1_w$[0:610]);
ixc_assign _zz_strnp_2 ( keyfilter_cmd_in[0], 
	_zy_simnet_keyfilter_cmd_in_2_w$);
ixc_assign_263 _zz_strnp_3 ( kdfstream_cmd_in[262:0], 
	_zy_simnet_kdfstream_cmd_in_3_w$[0:262]);
ixc_assign_4 _zz_strnp_4 ( kdf_cmd_in[3:0], _zy_simnet_kdf_cmd_in_4_w$[0:3]);
ixc_assign _zz_strnp_5 ( gcm_status_data_in[0], 
	_zy_simnet_gcm_status_data_in_5_w$);
ixc_assign_106 _zz_strnp_6 ( key_tlv_ob_tlv[105:0], 
	_zy_simnet_key_tlv_ob_tlv_6_w$[0:105]);
ixc_assign_611 _zz_strnp_7 ( _zy_simnet_gcm_cmd_in_9_w$[0:610], 
	gcm_cmd_in[610:0]);
ixc_assign _zz_strnp_8 ( _zy_simnet_keyfilter_cmd_in_12_w$, 
	keyfilter_cmd_in[0]);
ixc_assign_4 _zz_strnp_9 ( _zy_simnet_kdf_cmd_in_15_w$[0:3], kdf_cmd_in[3:0]);
ixc_assign_263 _zz_strnp_10 ( _zy_simnet_kdfstream_cmd_in_18_w$[0:262], 
	kdfstream_cmd_in[262:0]);
ixc_assign _zz_strnp_11 ( _zy_simnet_gcm_status_data_in_25_w$, 
	gcm_status_data_in[0]);
cr_kme_kop_tlv_inspector_xcm69 tlv_inspector ( .kme_internal_out_ack( 
	kme_internal_out_ack), .gcm_cmd_in( _zy_simnet_gcm_cmd_in_1_w$[0:610]), 
	.gcm_cmd_in_valid( gcm_cmd_in_valid), .gcm_tag_data_in( 
	gcm_tag_data_in[95:0]), .gcm_tag_data_in_valid( 
	gcm_tag_data_in_valid), .inspector_upsizer_valid( 
	inspector_upsizer_valid), .inspector_upsizer_eof( 
	inspector_upsizer_eof), .inspector_upsizer_data( 
	inspector_upsizer_data[63:0]), .keyfilter_cmd_in( 
	_zy_simnet_keyfilter_cmd_in_2_w$), .keyfilter_cmd_in_valid( 
	keyfilter_cmd_in_valid), .kdfstream_cmd_in( 
	_zy_simnet_kdfstream_cmd_in_3_w$[0:262]), .kdfstream_cmd_in_valid( 
	kdfstream_cmd_in_valid), .kdf_cmd_in( 
	_zy_simnet_kdf_cmd_in_4_w$[0:3]), .kdf_cmd_in_valid( kdf_cmd_in_valid), 
	.tlv_sb_data_in( tlv_sb_data_in[63:0]), .tlv_sb_data_in_valid( 
	tlv_sb_data_in_valid), .clk( clk), .rst_n( rst_n), .labels( { 
	\labels[7][271] , \labels[7][270] , \labels[7][269] , 
	\labels[7][268] , \labels[7][267] , \labels[7][266] , 
	\labels[7][265] , \labels[7][264] , \labels[7][263] , 
	\labels[7][262] , \labels[7][261] , \labels[7][260] , 
	\labels[7][259] , \labels[7][258] , \labels[7][257] , 
	\labels[7][256] , \labels[7][255] , \labels[7][254] , 
	\labels[7][253] , \labels[7][252] , \labels[7][251] , 
	\labels[7][250] , \labels[7][249] , \labels[7][248] , 
	\labels[7][247] , \labels[7][246] , \labels[7][245] , 
	\labels[7][244] , \labels[7][243] , \labels[7][242] , 
	\labels[7][241] , \labels[7][240] , \labels[7][239] , 
	\labels[7][238] , \labels[7][237] , \labels[7][236] , 
	\labels[7][235] , \labels[7][234] , \labels[7][233] , 
	\labels[7][232] , \labels[7][231] , \labels[7][230] , 
	\labels[7][229] , \labels[7][228] , \labels[7][227] , 
	\labels[7][226] , \labels[7][225] , \labels[7][224] , 
	\labels[7][223] , \labels[7][222] , \labels[7][221] , 
	\labels[7][220] , \labels[7][219] , \labels[7][218] , 
	\labels[7][217] , \labels[7][216] , \labels[7][215] , 
	\labels[7][214] , \labels[7][213] , \labels[7][212] , 
	\labels[7][211] , \labels[7][210] , \labels[7][209] , 
	\labels[7][208] , \labels[7][207] , \labels[7][206] , 
	\labels[7][205] , \labels[7][204] , \labels[7][203] , 
	\labels[7][202] , \labels[7][201] , \labels[7][200] , 
	\labels[7][199] , \labels[7][198] , \labels[7][197] , 
	\labels[7][196] , \labels[7][195] , \labels[7][194] , 
	\labels[7][193] , \labels[7][192] , \labels[7][191] , 
	\labels[7][190] , \labels[7][189] , \labels[7][188] , 
	\labels[7][187] , \labels[7][186] , \labels[7][185] , 
	\labels[7][184] , \labels[7][183] , \labels[7][182] , 
	\labels[7][181] , \labels[7][180] , \labels[7][179] , 
	\labels[7][178] , \labels[7][177] , \labels[7][176] , 
	\labels[7][175] , \labels[7][174] , \labels[7][173] , 
	\labels[7][172] , \labels[7][171] , \labels[7][170] , 
	\labels[7][169] , \labels[7][168] , \labels[7][167] , 
	\labels[7][166] , \labels[7][165] , \labels[7][164] , 
	\labels[7][163] , \labels[7][162] , \labels[7][161] , 
	\labels[7][160] , \labels[7][159] , \labels[7][158] , 
	\labels[7][157] , \labels[7][156] , \labels[7][155] , 
	\labels[7][154] , \labels[7][153] , \labels[7][152] , 
	\labels[7][151] , \labels[7][150] , \labels[7][149] , 
	\labels[7][148] , \labels[7][147] , \labels[7][146] , 
	\labels[7][145] , \labels[7][144] , \labels[7][143] , 
	\labels[7][142] , \labels[7][141] , \labels[7][140] , 
	\labels[7][139] , \labels[7][138] , \labels[7][137] , 
	\labels[7][136] , \labels[7][135] , \labels[7][134] , 
	\labels[7][133] , \labels[7][132] , \labels[7][131] , 
	\labels[7][130] , \labels[7][129] , \labels[7][128] , 
	\labels[7][127] , \labels[7][126] , \labels[7][125] , 
	\labels[7][124] , \labels[7][123] , \labels[7][122] , 
	\labels[7][121] , \labels[7][120] , \labels[7][119] , 
	\labels[7][118] , \labels[7][117] , \labels[7][116] , 
	\labels[7][115] , \labels[7][114] , \labels[7][113] , 
	\labels[7][112] , \labels[7][111] , \labels[7][110] , 
	\labels[7][109] , \labels[7][108] , \labels[7][107] , 
	\labels[7][106] , \labels[7][105] , \labels[7][104] , 
	\labels[7][103] , \labels[7][102] , \labels[7][101] , 
	\labels[7][100] , \labels[7][99] , \labels[7][98] , \labels[7][97] , 
	\labels[7][96] , \labels[7][95] , \labels[7][94] , \labels[7][93] , 
	\labels[7][92] , \labels[7][91] , \labels[7][90] , \labels[7][89] , 
	\labels[7][88] , \labels[7][87] , \labels[7][86] , \labels[7][85] , 
	\labels[7][84] , \labels[7][83] , \labels[7][82] , \labels[7][81] , 
	\labels[7][80] , \labels[7][79] , \labels[7][78] , \labels[7][77] , 
	\labels[7][76] , \labels[7][75] , \labels[7][74] , \labels[7][73] , 
	\labels[7][72] , \labels[7][71] , \labels[7][70] , \labels[7][69] , 
	\labels[7][68] , \labels[7][67] , \labels[7][66] , \labels[7][65] , 
	\labels[7][64] , \labels[7][63] , \labels[7][62] , \labels[7][61] , 
	\labels[7][60] , \labels[7][59] , \labels[7][58] , \labels[7][57] , 
	\labels[7][56] , \labels[7][55] , \labels[7][54] , \labels[7][53] , 
	\labels[7][52] , \labels[7][51] , \labels[7][50] , \labels[7][49] , 
	\labels[7][48] , \labels[7][47] , \labels[7][46] , \labels[7][45] , 
	\labels[7][44] , \labels[7][43] , \labels[7][42] , \labels[7][41] , 
	\labels[7][40] , \labels[7][39] , \labels[7][38] , \labels[7][37] , 
	\labels[7][36] , \labels[7][35] , \labels[7][34] , \labels[7][33] , 
	\labels[7][32] , \labels[7][31] , \labels[7][30] , \labels[7][29] , 
	\labels[7][28] , \labels[7][27] , \labels[7][26] , \labels[7][25] , 
	\labels[7][24] , \labels[7][23] , \labels[7][22] , \labels[7][21] , 
	\labels[7][20] , \labels[7][19] , \labels[7][18] , \labels[7][17] , 
	\labels[7][16] , \labels[7][15] , \labels[7][14] , \labels[7][13] , 
	\labels[7][12] , \labels[7][11] , \labels[7][10] , \labels[7][9] , 
	\labels[7][8] , \labels[7][7] , \labels[7][6] , \labels[7][5] , 
	\labels[7][4] , \labels[7][3] , \labels[7][2] , \labels[7][1] , 
	\labels[7][0] , \labels[6][271] , \labels[6][270] , \labels[6][269] , 
	\labels[6][268] , \labels[6][267] , \labels[6][266] , 
	\labels[6][265] , \labels[6][264] , \labels[6][263] , 
	\labels[6][262] , \labels[6][261] , \labels[6][260] , 
	\labels[6][259] , \labels[6][258] , \labels[6][257] , 
	\labels[6][256] , \labels[6][255] , \labels[6][254] , 
	\labels[6][253] , \labels[6][252] , \labels[6][251] , 
	\labels[6][250] , \labels[6][249] , \labels[6][248] , 
	\labels[6][247] , \labels[6][246] , \labels[6][245] , 
	\labels[6][244] , \labels[6][243] , \labels[6][242] , 
	\labels[6][241] , \labels[6][240] , \labels[6][239] , 
	\labels[6][238] , \labels[6][237] , \labels[6][236] , 
	\labels[6][235] , \labels[6][234] , \labels[6][233] , 
	\labels[6][232] , \labels[6][231] , \labels[6][230] , 
	\labels[6][229] , \labels[6][228] , \labels[6][227] , 
	\labels[6][226] , \labels[6][225] , \labels[6][224] , 
	\labels[6][223] , \labels[6][222] , \labels[6][221] , 
	\labels[6][220] , \labels[6][219] , \labels[6][218] , 
	\labels[6][217] , \labels[6][216] , \labels[6][215] , 
	\labels[6][214] , \labels[6][213] , \labels[6][212] , 
	\labels[6][211] , \labels[6][210] , \labels[6][209] , 
	\labels[6][208] , \labels[6][207] , \labels[6][206] , 
	\labels[6][205] , \labels[6][204] , \labels[6][203] , 
	\labels[6][202] , \labels[6][201] , \labels[6][200] , 
	\labels[6][199] , \labels[6][198] , \labels[6][197] , 
	\labels[6][196] , \labels[6][195] , \labels[6][194] , 
	\labels[6][193] , \labels[6][192] , \labels[6][191] , 
	\labels[6][190] , \labels[6][189] , \labels[6][188] , 
	\labels[6][187] , \labels[6][186] , \labels[6][185] , 
	\labels[6][184] , \labels[6][183] , \labels[6][182] , 
	\labels[6][181] , \labels[6][180] , \labels[6][179] , 
	\labels[6][178] , \labels[6][177] , \labels[6][176] , 
	\labels[6][175] , \labels[6][174] , \labels[6][173] , 
	\labels[6][172] , \labels[6][171] , \labels[6][170] , 
	\labels[6][169] , \labels[6][168] , \labels[6][167] , 
	\labels[6][166] , \labels[6][165] , \labels[6][164] , 
	\labels[6][163] , \labels[6][162] , \labels[6][161] , 
	\labels[6][160] , \labels[6][159] , \labels[6][158] , 
	\labels[6][157] , \labels[6][156] , \labels[6][155] , 
	\labels[6][154] , \labels[6][153] , \labels[6][152] , 
	\labels[6][151] , \labels[6][150] , \labels[6][149] , 
	\labels[6][148] , \labels[6][147] , \labels[6][146] , 
	\labels[6][145] , \labels[6][144] , \labels[6][143] , 
	\labels[6][142] , \labels[6][141] , \labels[6][140] , 
	\labels[6][139] , \labels[6][138] , \labels[6][137] , 
	\labels[6][136] , \labels[6][135] , \labels[6][134] , 
	\labels[6][133] , \labels[6][132] , \labels[6][131] , 
	\labels[6][130] , \labels[6][129] , \labels[6][128] , 
	\labels[6][127] , \labels[6][126] , \labels[6][125] , 
	\labels[6][124] , \labels[6][123] , \labels[6][122] , 
	\labels[6][121] , \labels[6][120] , \labels[6][119] , 
	\labels[6][118] , \labels[6][117] , \labels[6][116] , 
	\labels[6][115] , \labels[6][114] , \labels[6][113] , 
	\labels[6][112] , \labels[6][111] , \labels[6][110] , 
	\labels[6][109] , \labels[6][108] , \labels[6][107] , 
	\labels[6][106] , \labels[6][105] , \labels[6][104] , 
	\labels[6][103] , \labels[6][102] , \labels[6][101] , 
	\labels[6][100] , \labels[6][99] , \labels[6][98] , \labels[6][97] , 
	\labels[6][96] , \labels[6][95] , \labels[6][94] , \labels[6][93] , 
	\labels[6][92] , \labels[6][91] , \labels[6][90] , \labels[6][89] , 
	\labels[6][88] , \labels[6][87] , \labels[6][86] , \labels[6][85] , 
	\labels[6][84] , \labels[6][83] , \labels[6][82] , \labels[6][81] , 
	\labels[6][80] , \labels[6][79] , \labels[6][78] , \labels[6][77] , 
	\labels[6][76] , \labels[6][75] , \labels[6][74] , \labels[6][73] , 
	\labels[6][72] , \labels[6][71] , \labels[6][70] , \labels[6][69] , 
	\labels[6][68] , \labels[6][67] , \labels[6][66] , \labels[6][65] , 
	\labels[6][64] , \labels[6][63] , \labels[6][62] , \labels[6][61] , 
	\labels[6][60] , \labels[6][59] , \labels[6][58] , \labels[6][57] , 
	\labels[6][56] , \labels[6][55] , \labels[6][54] , \labels[6][53] , 
	\labels[6][52] , \labels[6][51] , \labels[6][50] , \labels[6][49] , 
	\labels[6][48] , \labels[6][47] , \labels[6][46] , \labels[6][45] , 
	\labels[6][44] , \labels[6][43] , \labels[6][42] , \labels[6][41] , 
	\labels[6][40] , \labels[6][39] , \labels[6][38] , \labels[6][37] , 
	\labels[6][36] , \labels[6][35] , \labels[6][34] , \labels[6][33] , 
	\labels[6][32] , \labels[6][31] , \labels[6][30] , \labels[6][29] , 
	\labels[6][28] , \labels[6][27] , \labels[6][26] , \labels[6][25] , 
	\labels[6][24] , \labels[6][23] , \labels[6][22] , \labels[6][21] , 
	\labels[6][20] , \labels[6][19] , \labels[6][18] , \labels[6][17] , 
	\labels[6][16] , \labels[6][15] , \labels[6][14] , \labels[6][13] , 
	\labels[6][12] , \labels[6][11] , \labels[6][10] , \labels[6][9] , 
	\labels[6][8] , \labels[6][7] , \labels[6][6] , \labels[6][5] , 
	\labels[6][4] , \labels[6][3] , \labels[6][2] , \labels[6][1] , 
	\labels[6][0] , \labels[5][271] , \labels[5][270] , \labels[5][269] , 
	\labels[5][268] , \labels[5][267] , \labels[5][266] , 
	\labels[5][265] , \labels[5][264] , \labels[5][263] , 
	\labels[5][262] , \labels[5][261] , \labels[5][260] , 
	\labels[5][259] , \labels[5][258] , \labels[5][257] , 
	\labels[5][256] , \labels[5][255] , \labels[5][254] , 
	\labels[5][253] , \labels[5][252] , \labels[5][251] , 
	\labels[5][250] , \labels[5][249] , \labels[5][248] , 
	\labels[5][247] , \labels[5][246] , \labels[5][245] , 
	\labels[5][244] , \labels[5][243] , \labels[5][242] , 
	\labels[5][241] , \labels[5][240] , \labels[5][239] , 
	\labels[5][238] , \labels[5][237] , \labels[5][236] , 
	\labels[5][235] , \labels[5][234] , \labels[5][233] , 
	\labels[5][232] , \labels[5][231] , \labels[5][230] , 
	\labels[5][229] , \labels[5][228] , \labels[5][227] , 
	\labels[5][226] , \labels[5][225] , \labels[5][224] , 
	\labels[5][223] , \labels[5][222] , \labels[5][221] , 
	\labels[5][220] , \labels[5][219] , \labels[5][218] , 
	\labels[5][217] , \labels[5][216] , \labels[5][215] , 
	\labels[5][214] , \labels[5][213] , \labels[5][212] , 
	\labels[5][211] , \labels[5][210] , \labels[5][209] , 
	\labels[5][208] , \labels[5][207] , \labels[5][206] , 
	\labels[5][205] , \labels[5][204] , \labels[5][203] , 
	\labels[5][202] , \labels[5][201] , \labels[5][200] , 
	\labels[5][199] , \labels[5][198] , \labels[5][197] , 
	\labels[5][196] , \labels[5][195] , \labels[5][194] , 
	\labels[5][193] , \labels[5][192] , \labels[5][191] , 
	\labels[5][190] , \labels[5][189] , \labels[5][188] , 
	\labels[5][187] , \labels[5][186] , \labels[5][185] , 
	\labels[5][184] , \labels[5][183] , \labels[5][182] , 
	\labels[5][181] , \labels[5][180] , \labels[5][179] , 
	\labels[5][178] , \labels[5][177] , \labels[5][176] , 
	\labels[5][175] , \labels[5][174] , \labels[5][173] , 
	\labels[5][172] , \labels[5][171] , \labels[5][170] , 
	\labels[5][169] , \labels[5][168] , \labels[5][167] , 
	\labels[5][166] , \labels[5][165] , \labels[5][164] , 
	\labels[5][163] , \labels[5][162] , \labels[5][161] , 
	\labels[5][160] , \labels[5][159] , \labels[5][158] , 
	\labels[5][157] , \labels[5][156] , \labels[5][155] , 
	\labels[5][154] , \labels[5][153] , \labels[5][152] , 
	\labels[5][151] , \labels[5][150] , \labels[5][149] , 
	\labels[5][148] , \labels[5][147] , \labels[5][146] , 
	\labels[5][145] , \labels[5][144] , \labels[5][143] , 
	\labels[5][142] , \labels[5][141] , \labels[5][140] , 
	\labels[5][139] , \labels[5][138] , \labels[5][137] , 
	\labels[5][136] , \labels[5][135] , \labels[5][134] , 
	\labels[5][133] , \labels[5][132] , \labels[5][131] , 
	\labels[5][130] , \labels[5][129] , \labels[5][128] , 
	\labels[5][127] , \labels[5][126] , \labels[5][125] , 
	\labels[5][124] , \labels[5][123] , \labels[5][122] , 
	\labels[5][121] , \labels[5][120] , \labels[5][119] , 
	\labels[5][118] , \labels[5][117] , \labels[5][116] , 
	\labels[5][115] , \labels[5][114] , \labels[5][113] , 
	\labels[5][112] , \labels[5][111] , \labels[5][110] , 
	\labels[5][109] , \labels[5][108] , \labels[5][107] , 
	\labels[5][106] , \labels[5][105] , \labels[5][104] , 
	\labels[5][103] , \labels[5][102] , \labels[5][101] , 
	\labels[5][100] , \labels[5][99] , \labels[5][98] , \labels[5][97] , 
	\labels[5][96] , \labels[5][95] , \labels[5][94] , \labels[5][93] , 
	\labels[5][92] , \labels[5][91] , \labels[5][90] , \labels[5][89] , 
	\labels[5][88] , \labels[5][87] , \labels[5][86] , \labels[5][85] , 
	\labels[5][84] , \labels[5][83] , \labels[5][82] , \labels[5][81] , 
	\labels[5][80] , \labels[5][79] , \labels[5][78] , \labels[5][77] , 
	\labels[5][76] , \labels[5][75] , \labels[5][74] , \labels[5][73] , 
	\labels[5][72] , \labels[5][71] , \labels[5][70] , \labels[5][69] , 
	\labels[5][68] , \labels[5][67] , \labels[5][66] , \labels[5][65] , 
	\labels[5][64] , \labels[5][63] , \labels[5][62] , \labels[5][61] , 
	\labels[5][60] , \labels[5][59] , \labels[5][58] , \labels[5][57] , 
	\labels[5][56] , \labels[5][55] , \labels[5][54] , \labels[5][53] , 
	\labels[5][52] , \labels[5][51] , \labels[5][50] , \labels[5][49] , 
	\labels[5][48] , \labels[5][47] , \labels[5][46] , \labels[5][45] , 
	\labels[5][44] , \labels[5][43] , \labels[5][42] , \labels[5][41] , 
	\labels[5][40] , \labels[5][39] , \labels[5][38] , \labels[5][37] , 
	\labels[5][36] , \labels[5][35] , \labels[5][34] , \labels[5][33] , 
	\labels[5][32] , \labels[5][31] , \labels[5][30] , \labels[5][29] , 
	\labels[5][28] , \labels[5][27] , \labels[5][26] , \labels[5][25] , 
	\labels[5][24] , \labels[5][23] , \labels[5][22] , \labels[5][21] , 
	\labels[5][20] , \labels[5][19] , \labels[5][18] , \labels[5][17] , 
	\labels[5][16] , \labels[5][15] , \labels[5][14] , \labels[5][13] , 
	\labels[5][12] , \labels[5][11] , \labels[5][10] , \labels[5][9] , 
	\labels[5][8] , \labels[5][7] , \labels[5][6] , \labels[5][5] , 
	\labels[5][4] , \labels[5][3] , \labels[5][2] , \labels[5][1] , 
	\labels[5][0] , \labels[4][271] , \labels[4][270] , \labels[4][269] , 
	\labels[4][268] , \labels[4][267] , \labels[4][266] , 
	\labels[4][265] , \labels[4][264] , \labels[4][263] , 
	\labels[4][262] , \labels[4][261] , \labels[4][260] , 
	\labels[4][259] , \labels[4][258] , \labels[4][257] , 
	\labels[4][256] , \labels[4][255] , \labels[4][254] , 
	\labels[4][253] , \labels[4][252] , \labels[4][251] , 
	\labels[4][250] , \labels[4][249] , \labels[4][248] , 
	\labels[4][247] , \labels[4][246] , \labels[4][245] , 
	\labels[4][244] , \labels[4][243] , \labels[4][242] , 
	\labels[4][241] , \labels[4][240] , \labels[4][239] , 
	\labels[4][238] , \labels[4][237] , \labels[4][236] , 
	\labels[4][235] , \labels[4][234] , \labels[4][233] , 
	\labels[4][232] , \labels[4][231] , \labels[4][230] , 
	\labels[4][229] , \labels[4][228] , \labels[4][227] , 
	\labels[4][226] , \labels[4][225] , \labels[4][224] , 
	\labels[4][223] , \labels[4][222] , \labels[4][221] , 
	\labels[4][220] , \labels[4][219] , \labels[4][218] , 
	\labels[4][217] , \labels[4][216] , \labels[4][215] , 
	\labels[4][214] , \labels[4][213] , \labels[4][212] , 
	\labels[4][211] , \labels[4][210] , \labels[4][209] , 
	\labels[4][208] , \labels[4][207] , \labels[4][206] , 
	\labels[4][205] , \labels[4][204] , \labels[4][203] , 
	\labels[4][202] , \labels[4][201] , \labels[4][200] , 
	\labels[4][199] , \labels[4][198] , \labels[4][197] , 
	\labels[4][196] , \labels[4][195] , \labels[4][194] , 
	\labels[4][193] , \labels[4][192] , \labels[4][191] , 
	\labels[4][190] , \labels[4][189] , \labels[4][188] , 
	\labels[4][187] , \labels[4][186] , \labels[4][185] , 
	\labels[4][184] , \labels[4][183] , \labels[4][182] , 
	\labels[4][181] , \labels[4][180] , \labels[4][179] , 
	\labels[4][178] , \labels[4][177] , \labels[4][176] , 
	\labels[4][175] , \labels[4][174] , \labels[4][173] , 
	\labels[4][172] , \labels[4][171] , \labels[4][170] , 
	\labels[4][169] , \labels[4][168] , \labels[4][167] , 
	\labels[4][166] , \labels[4][165] , \labels[4][164] , 
	\labels[4][163] , \labels[4][162] , \labels[4][161] , 
	\labels[4][160] , \labels[4][159] , \labels[4][158] , 
	\labels[4][157] , \labels[4][156] , \labels[4][155] , 
	\labels[4][154] , \labels[4][153] , \labels[4][152] , 
	\labels[4][151] , \labels[4][150] , \labels[4][149] , 
	\labels[4][148] , \labels[4][147] , \labels[4][146] , 
	\labels[4][145] , \labels[4][144] , \labels[4][143] , 
	\labels[4][142] , \labels[4][141] , \labels[4][140] , 
	\labels[4][139] , \labels[4][138] , \labels[4][137] , 
	\labels[4][136] , \labels[4][135] , \labels[4][134] , 
	\labels[4][133] , \labels[4][132] , \labels[4][131] , 
	\labels[4][130] , \labels[4][129] , \labels[4][128] , 
	\labels[4][127] , \labels[4][126] , \labels[4][125] , 
	\labels[4][124] , \labels[4][123] , \labels[4][122] , 
	\labels[4][121] , \labels[4][120] , \labels[4][119] , 
	\labels[4][118] , \labels[4][117] , \labels[4][116] , 
	\labels[4][115] , \labels[4][114] , \labels[4][113] , 
	\labels[4][112] , \labels[4][111] , \labels[4][110] , 
	\labels[4][109] , \labels[4][108] , \labels[4][107] , 
	\labels[4][106] , \labels[4][105] , \labels[4][104] , 
	\labels[4][103] , \labels[4][102] , \labels[4][101] , 
	\labels[4][100] , \labels[4][99] , \labels[4][98] , \labels[4][97] , 
	\labels[4][96] , \labels[4][95] , \labels[4][94] , \labels[4][93] , 
	\labels[4][92] , \labels[4][91] , \labels[4][90] , \labels[4][89] , 
	\labels[4][88] , \labels[4][87] , \labels[4][86] , \labels[4][85] , 
	\labels[4][84] , \labels[4][83] , \labels[4][82] , \labels[4][81] , 
	\labels[4][80] , \labels[4][79] , \labels[4][78] , \labels[4][77] , 
	\labels[4][76] , \labels[4][75] , \labels[4][74] , \labels[4][73] , 
	\labels[4][72] , \labels[4][71] , \labels[4][70] , \labels[4][69] , 
	\labels[4][68] , \labels[4][67] , \labels[4][66] , \labels[4][65] , 
	\labels[4][64] , \labels[4][63] , \labels[4][62] , \labels[4][61] , 
	\labels[4][60] , \labels[4][59] , \labels[4][58] , \labels[4][57] , 
	\labels[4][56] , \labels[4][55] , \labels[4][54] , \labels[4][53] , 
	\labels[4][52] , \labels[4][51] , \labels[4][50] , \labels[4][49] , 
	\labels[4][48] , \labels[4][47] , \labels[4][46] , \labels[4][45] , 
	\labels[4][44] , \labels[4][43] , \labels[4][42] , \labels[4][41] , 
	\labels[4][40] , \labels[4][39] , \labels[4][38] , \labels[4][37] , 
	\labels[4][36] , \labels[4][35] , \labels[4][34] , \labels[4][33] , 
	\labels[4][32] , \labels[4][31] , \labels[4][30] , \labels[4][29] , 
	\labels[4][28] , \labels[4][27] , \labels[4][26] , \labels[4][25] , 
	\labels[4][24] , \labels[4][23] , \labels[4][22] , \labels[4][21] , 
	\labels[4][20] , \labels[4][19] , \labels[4][18] , \labels[4][17] , 
	\labels[4][16] , \labels[4][15] , \labels[4][14] , \labels[4][13] , 
	\labels[4][12] , \labels[4][11] , \labels[4][10] , \labels[4][9] , 
	\labels[4][8] , \labels[4][7] , \labels[4][6] , \labels[4][5] , 
	\labels[4][4] , \labels[4][3] , \labels[4][2] , \labels[4][1] , 
	\labels[4][0] , \labels[3][271] , \labels[3][270] , \labels[3][269] , 
	\labels[3][268] , \labels[3][267] , \labels[3][266] , 
	\labels[3][265] , \labels[3][264] , \labels[3][263] , 
	\labels[3][262] , \labels[3][261] , \labels[3][260] , 
	\labels[3][259] , \labels[3][258] , \labels[3][257] , 
	\labels[3][256] , \labels[3][255] , \labels[3][254] , 
	\labels[3][253] , \labels[3][252] , \labels[3][251] , 
	\labels[3][250] , \labels[3][249] , \labels[3][248] , 
	\labels[3][247] , \labels[3][246] , \labels[3][245] , 
	\labels[3][244] , \labels[3][243] , \labels[3][242] , 
	\labels[3][241] , \labels[3][240] , \labels[3][239] , 
	\labels[3][238] , \labels[3][237] , \labels[3][236] , 
	\labels[3][235] , \labels[3][234] , \labels[3][233] , 
	\labels[3][232] , \labels[3][231] , \labels[3][230] , 
	\labels[3][229] , \labels[3][228] , \labels[3][227] , 
	\labels[3][226] , \labels[3][225] , \labels[3][224] , 
	\labels[3][223] , \labels[3][222] , \labels[3][221] , 
	\labels[3][220] , \labels[3][219] , \labels[3][218] , 
	\labels[3][217] , \labels[3][216] , \labels[3][215] , 
	\labels[3][214] , \labels[3][213] , \labels[3][212] , 
	\labels[3][211] , \labels[3][210] , \labels[3][209] , 
	\labels[3][208] , \labels[3][207] , \labels[3][206] , 
	\labels[3][205] , \labels[3][204] , \labels[3][203] , 
	\labels[3][202] , \labels[3][201] , \labels[3][200] , 
	\labels[3][199] , \labels[3][198] , \labels[3][197] , 
	\labels[3][196] , \labels[3][195] , \labels[3][194] , 
	\labels[3][193] , \labels[3][192] , \labels[3][191] , 
	\labels[3][190] , \labels[3][189] , \labels[3][188] , 
	\labels[3][187] , \labels[3][186] , \labels[3][185] , 
	\labels[3][184] , \labels[3][183] , \labels[3][182] , 
	\labels[3][181] , \labels[3][180] , \labels[3][179] , 
	\labels[3][178] , \labels[3][177] , \labels[3][176] , 
	\labels[3][175] , \labels[3][174] , \labels[3][173] , 
	\labels[3][172] , \labels[3][171] , \labels[3][170] , 
	\labels[3][169] , \labels[3][168] , \labels[3][167] , 
	\labels[3][166] , \labels[3][165] , \labels[3][164] , 
	\labels[3][163] , \labels[3][162] , \labels[3][161] , 
	\labels[3][160] , \labels[3][159] , \labels[3][158] , 
	\labels[3][157] , \labels[3][156] , \labels[3][155] , 
	\labels[3][154] , \labels[3][153] , \labels[3][152] , 
	\labels[3][151] , \labels[3][150] , \labels[3][149] , 
	\labels[3][148] , \labels[3][147] , \labels[3][146] , 
	\labels[3][145] , \labels[3][144] , \labels[3][143] , 
	\labels[3][142] , \labels[3][141] , \labels[3][140] , 
	\labels[3][139] , \labels[3][138] , \labels[3][137] , 
	\labels[3][136] , \labels[3][135] , \labels[3][134] , 
	\labels[3][133] , \labels[3][132] , \labels[3][131] , 
	\labels[3][130] , \labels[3][129] , \labels[3][128] , 
	\labels[3][127] , \labels[3][126] , \labels[3][125] , 
	\labels[3][124] , \labels[3][123] , \labels[3][122] , 
	\labels[3][121] , \labels[3][120] , \labels[3][119] , 
	\labels[3][118] , \labels[3][117] , \labels[3][116] , 
	\labels[3][115] , \labels[3][114] , \labels[3][113] , 
	\labels[3][112] , \labels[3][111] , \labels[3][110] , 
	\labels[3][109] , \labels[3][108] , \labels[3][107] , 
	\labels[3][106] , \labels[3][105] , \labels[3][104] , 
	\labels[3][103] , \labels[3][102] , \labels[3][101] , 
	\labels[3][100] , \labels[3][99] , \labels[3][98] , \labels[3][97] , 
	\labels[3][96] , \labels[3][95] , \labels[3][94] , \labels[3][93] , 
	\labels[3][92] , \labels[3][91] , \labels[3][90] , \labels[3][89] , 
	\labels[3][88] , \labels[3][87] , \labels[3][86] , \labels[3][85] , 
	\labels[3][84] , \labels[3][83] , \labels[3][82] , \labels[3][81] , 
	\labels[3][80] , \labels[3][79] , \labels[3][78] , \labels[3][77] , 
	\labels[3][76] , \labels[3][75] , \labels[3][74] , \labels[3][73] , 
	\labels[3][72] , \labels[3][71] , \labels[3][70] , \labels[3][69] , 
	\labels[3][68] , \labels[3][67] , \labels[3][66] , \labels[3][65] , 
	\labels[3][64] , \labels[3][63] , \labels[3][62] , \labels[3][61] , 
	\labels[3][60] , \labels[3][59] , \labels[3][58] , \labels[3][57] , 
	\labels[3][56] , \labels[3][55] , \labels[3][54] , \labels[3][53] , 
	\labels[3][52] , \labels[3][51] , \labels[3][50] , \labels[3][49] , 
	\labels[3][48] , \labels[3][47] , \labels[3][46] , \labels[3][45] , 
	\labels[3][44] , \labels[3][43] , \labels[3][42] , \labels[3][41] , 
	\labels[3][40] , \labels[3][39] , \labels[3][38] , \labels[3][37] , 
	\labels[3][36] , \labels[3][35] , \labels[3][34] , \labels[3][33] , 
	\labels[3][32] , \labels[3][31] , \labels[3][30] , \labels[3][29] , 
	\labels[3][28] , \labels[3][27] , \labels[3][26] , \labels[3][25] , 
	\labels[3][24] , \labels[3][23] , \labels[3][22] , \labels[3][21] , 
	\labels[3][20] , \labels[3][19] , \labels[3][18] , \labels[3][17] , 
	\labels[3][16] , \labels[3][15] , \labels[3][14] , \labels[3][13] , 
	\labels[3][12] , \labels[3][11] , \labels[3][10] , \labels[3][9] , 
	\labels[3][8] , \labels[3][7] , \labels[3][6] , \labels[3][5] , 
	\labels[3][4] , \labels[3][3] , \labels[3][2] , \labels[3][1] , 
	\labels[3][0] , \labels[2][271] , \labels[2][270] , \labels[2][269] , 
	\labels[2][268] , \labels[2][267] , \labels[2][266] , 
	\labels[2][265] , \labels[2][264] , \labels[2][263] , 
	\labels[2][262] , \labels[2][261] , \labels[2][260] , 
	\labels[2][259] , \labels[2][258] , \labels[2][257] , 
	\labels[2][256] , \labels[2][255] , \labels[2][254] , 
	\labels[2][253] , \labels[2][252] , \labels[2][251] , 
	\labels[2][250] , \labels[2][249] , \labels[2][248] , 
	\labels[2][247] , \labels[2][246] , \labels[2][245] , 
	\labels[2][244] , \labels[2][243] , \labels[2][242] , 
	\labels[2][241] , \labels[2][240] , \labels[2][239] , 
	\labels[2][238] , \labels[2][237] , \labels[2][236] , 
	\labels[2][235] , \labels[2][234] , \labels[2][233] , 
	\labels[2][232] , \labels[2][231] , \labels[2][230] , 
	\labels[2][229] , \labels[2][228] , \labels[2][227] , 
	\labels[2][226] , \labels[2][225] , \labels[2][224] , 
	\labels[2][223] , \labels[2][222] , \labels[2][221] , 
	\labels[2][220] , \labels[2][219] , \labels[2][218] , 
	\labels[2][217] , \labels[2][216] , \labels[2][215] , 
	\labels[2][214] , \labels[2][213] , \labels[2][212] , 
	\labels[2][211] , \labels[2][210] , \labels[2][209] , 
	\labels[2][208] , \labels[2][207] , \labels[2][206] , 
	\labels[2][205] , \labels[2][204] , \labels[2][203] , 
	\labels[2][202] , \labels[2][201] , \labels[2][200] , 
	\labels[2][199] , \labels[2][198] , \labels[2][197] , 
	\labels[2][196] , \labels[2][195] , \labels[2][194] , 
	\labels[2][193] , \labels[2][192] , \labels[2][191] , 
	\labels[2][190] , \labels[2][189] , \labels[2][188] , 
	\labels[2][187] , \labels[2][186] , \labels[2][185] , 
	\labels[2][184] , \labels[2][183] , \labels[2][182] , 
	\labels[2][181] , \labels[2][180] , \labels[2][179] , 
	\labels[2][178] , \labels[2][177] , \labels[2][176] , 
	\labels[2][175] , \labels[2][174] , \labels[2][173] , 
	\labels[2][172] , \labels[2][171] , \labels[2][170] , 
	\labels[2][169] , \labels[2][168] , \labels[2][167] , 
	\labels[2][166] , \labels[2][165] , \labels[2][164] , 
	\labels[2][163] , \labels[2][162] , \labels[2][161] , 
	\labels[2][160] , \labels[2][159] , \labels[2][158] , 
	\labels[2][157] , \labels[2][156] , \labels[2][155] , 
	\labels[2][154] , \labels[2][153] , \labels[2][152] , 
	\labels[2][151] , \labels[2][150] , \labels[2][149] , 
	\labels[2][148] , \labels[2][147] , \labels[2][146] , 
	\labels[2][145] , \labels[2][144] , \labels[2][143] , 
	\labels[2][142] , \labels[2][141] , \labels[2][140] , 
	\labels[2][139] , \labels[2][138] , \labels[2][137] , 
	\labels[2][136] , \labels[2][135] , \labels[2][134] , 
	\labels[2][133] , \labels[2][132] , \labels[2][131] , 
	\labels[2][130] , \labels[2][129] , \labels[2][128] , 
	\labels[2][127] , \labels[2][126] , \labels[2][125] , 
	\labels[2][124] , \labels[2][123] , \labels[2][122] , 
	\labels[2][121] , \labels[2][120] , \labels[2][119] , 
	\labels[2][118] , \labels[2][117] , \labels[2][116] , 
	\labels[2][115] , \labels[2][114] , \labels[2][113] , 
	\labels[2][112] , \labels[2][111] , \labels[2][110] , 
	\labels[2][109] , \labels[2][108] , \labels[2][107] , 
	\labels[2][106] , \labels[2][105] , \labels[2][104] , 
	\labels[2][103] , \labels[2][102] , \labels[2][101] , 
	\labels[2][100] , \labels[2][99] , \labels[2][98] , \labels[2][97] , 
	\labels[2][96] , \labels[2][95] , \labels[2][94] , \labels[2][93] , 
	\labels[2][92] , \labels[2][91] , \labels[2][90] , \labels[2][89] , 
	\labels[2][88] , \labels[2][87] , \labels[2][86] , \labels[2][85] , 
	\labels[2][84] , \labels[2][83] , \labels[2][82] , \labels[2][81] , 
	\labels[2][80] , \labels[2][79] , \labels[2][78] , \labels[2][77] , 
	\labels[2][76] , \labels[2][75] , \labels[2][74] , \labels[2][73] , 
	\labels[2][72] , \labels[2][71] , \labels[2][70] , \labels[2][69] , 
	\labels[2][68] , \labels[2][67] , \labels[2][66] , \labels[2][65] , 
	\labels[2][64] , \labels[2][63] , \labels[2][62] , \labels[2][61] , 
	\labels[2][60] , \labels[2][59] , \labels[2][58] , \labels[2][57] , 
	\labels[2][56] , \labels[2][55] , \labels[2][54] , \labels[2][53] , 
	\labels[2][52] , \labels[2][51] , \labels[2][50] , \labels[2][49] , 
	\labels[2][48] , \labels[2][47] , \labels[2][46] , \labels[2][45] , 
	\labels[2][44] , \labels[2][43] , \labels[2][42] , \labels[2][41] , 
	\labels[2][40] , \labels[2][39] , \labels[2][38] , \labels[2][37] , 
	\labels[2][36] , \labels[2][35] , \labels[2][34] , \labels[2][33] , 
	\labels[2][32] , \labels[2][31] , \labels[2][30] , \labels[2][29] , 
	\labels[2][28] , \labels[2][27] , \labels[2][26] , \labels[2][25] , 
	\labels[2][24] , \labels[2][23] , \labels[2][22] , \labels[2][21] , 
	\labels[2][20] , \labels[2][19] , \labels[2][18] , \labels[2][17] , 
	\labels[2][16] , \labels[2][15] , \labels[2][14] , \labels[2][13] , 
	\labels[2][12] , \labels[2][11] , \labels[2][10] , \labels[2][9] , 
	\labels[2][8] , \labels[2][7] , \labels[2][6] , \labels[2][5] , 
	\labels[2][4] , \labels[2][3] , \labels[2][2] , \labels[2][1] , 
	\labels[2][0] , \labels[1][271] , \labels[1][270] , \labels[1][269] , 
	\labels[1][268] , \labels[1][267] , \labels[1][266] , 
	\labels[1][265] , \labels[1][264] , \labels[1][263] , 
	\labels[1][262] , \labels[1][261] , \labels[1][260] , 
	\labels[1][259] , \labels[1][258] , \labels[1][257] , 
	\labels[1][256] , \labels[1][255] , \labels[1][254] , 
	\labels[1][253] , \labels[1][252] , \labels[1][251] , 
	\labels[1][250] , \labels[1][249] , \labels[1][248] , 
	\labels[1][247] , \labels[1][246] , \labels[1][245] , 
	\labels[1][244] , \labels[1][243] , \labels[1][242] , 
	\labels[1][241] , \labels[1][240] , \labels[1][239] , 
	\labels[1][238] , \labels[1][237] , \labels[1][236] , 
	\labels[1][235] , \labels[1][234] , \labels[1][233] , 
	\labels[1][232] , \labels[1][231] , \labels[1][230] , 
	\labels[1][229] , \labels[1][228] , \labels[1][227] , 
	\labels[1][226] , \labels[1][225] , \labels[1][224] , 
	\labels[1][223] , \labels[1][222] , \labels[1][221] , 
	\labels[1][220] , \labels[1][219] , \labels[1][218] , 
	\labels[1][217] , \labels[1][216] , \labels[1][215] , 
	\labels[1][214] , \labels[1][213] , \labels[1][212] , 
	\labels[1][211] , \labels[1][210] , \labels[1][209] , 
	\labels[1][208] , \labels[1][207] , \labels[1][206] , 
	\labels[1][205] , \labels[1][204] , \labels[1][203] , 
	\labels[1][202] , \labels[1][201] , \labels[1][200] , 
	\labels[1][199] , \labels[1][198] , \labels[1][197] , 
	\labels[1][196] , \labels[1][195] , \labels[1][194] , 
	\labels[1][193] , \labels[1][192] , \labels[1][191] , 
	\labels[1][190] , \labels[1][189] , \labels[1][188] , 
	\labels[1][187] , \labels[1][186] , \labels[1][185] , 
	\labels[1][184] , \labels[1][183] , \labels[1][182] , 
	\labels[1][181] , \labels[1][180] , \labels[1][179] , 
	\labels[1][178] , \labels[1][177] , \labels[1][176] , 
	\labels[1][175] , \labels[1][174] , \labels[1][173] , 
	\labels[1][172] , \labels[1][171] , \labels[1][170] , 
	\labels[1][169] , \labels[1][168] , \labels[1][167] , 
	\labels[1][166] , \labels[1][165] , \labels[1][164] , 
	\labels[1][163] , \labels[1][162] , \labels[1][161] , 
	\labels[1][160] , \labels[1][159] , \labels[1][158] , 
	\labels[1][157] , \labels[1][156] , \labels[1][155] , 
	\labels[1][154] , \labels[1][153] , \labels[1][152] , 
	\labels[1][151] , \labels[1][150] , \labels[1][149] , 
	\labels[1][148] , \labels[1][147] , \labels[1][146] , 
	\labels[1][145] , \labels[1][144] , \labels[1][143] , 
	\labels[1][142] , \labels[1][141] , \labels[1][140] , 
	\labels[1][139] , \labels[1][138] , \labels[1][137] , 
	\labels[1][136] , \labels[1][135] , \labels[1][134] , 
	\labels[1][133] , \labels[1][132] , \labels[1][131] , 
	\labels[1][130] , \labels[1][129] , \labels[1][128] , 
	\labels[1][127] , \labels[1][126] , \labels[1][125] , 
	\labels[1][124] , \labels[1][123] , \labels[1][122] , 
	\labels[1][121] , \labels[1][120] , \labels[1][119] , 
	\labels[1][118] , \labels[1][117] , \labels[1][116] , 
	\labels[1][115] , \labels[1][114] , \labels[1][113] , 
	\labels[1][112] , \labels[1][111] , \labels[1][110] , 
	\labels[1][109] , \labels[1][108] , \labels[1][107] , 
	\labels[1][106] , \labels[1][105] , \labels[1][104] , 
	\labels[1][103] , \labels[1][102] , \labels[1][101] , 
	\labels[1][100] , \labels[1][99] , \labels[1][98] , \labels[1][97] , 
	\labels[1][96] , \labels[1][95] , \labels[1][94] , \labels[1][93] , 
	\labels[1][92] , \labels[1][91] , \labels[1][90] , \labels[1][89] , 
	\labels[1][88] , \labels[1][87] , \labels[1][86] , \labels[1][85] , 
	\labels[1][84] , \labels[1][83] , \labels[1][82] , \labels[1][81] , 
	\labels[1][80] , \labels[1][79] , \labels[1][78] , \labels[1][77] , 
	\labels[1][76] , \labels[1][75] , \labels[1][74] , \labels[1][73] , 
	\labels[1][72] , \labels[1][71] , \labels[1][70] , \labels[1][69] , 
	\labels[1][68] , \labels[1][67] , \labels[1][66] , \labels[1][65] , 
	\labels[1][64] , \labels[1][63] , \labels[1][62] , \labels[1][61] , 
	\labels[1][60] , \labels[1][59] , \labels[1][58] , \labels[1][57] , 
	\labels[1][56] , \labels[1][55] , \labels[1][54] , \labels[1][53] , 
	\labels[1][52] , \labels[1][51] , \labels[1][50] , \labels[1][49] , 
	\labels[1][48] , \labels[1][47] , \labels[1][46] , \labels[1][45] , 
	\labels[1][44] , \labels[1][43] , \labels[1][42] , \labels[1][41] , 
	\labels[1][40] , \labels[1][39] , \labels[1][38] , \labels[1][37] , 
	\labels[1][36] , \labels[1][35] , \labels[1][34] , \labels[1][33] , 
	\labels[1][32] , \labels[1][31] , \labels[1][30] , \labels[1][29] , 
	\labels[1][28] , \labels[1][27] , \labels[1][26] , \labels[1][25] , 
	\labels[1][24] , \labels[1][23] , \labels[1][22] , \labels[1][21] , 
	\labels[1][20] , \labels[1][19] , \labels[1][18] , \labels[1][17] , 
	\labels[1][16] , \labels[1][15] , \labels[1][14] , \labels[1][13] , 
	\labels[1][12] , \labels[1][11] , \labels[1][10] , \labels[1][9] , 
	\labels[1][8] , \labels[1][7] , \labels[1][6] , \labels[1][5] , 
	\labels[1][4] , \labels[1][3] , \labels[1][2] , \labels[1][1] , 
	\labels[1][0] , \labels[0][271] , \labels[0][270] , \labels[0][269] , 
	\labels[0][268] , \labels[0][267] , \labels[0][266] , 
	\labels[0][265] , \labels[0][264] , \labels[0][263] , 
	\labels[0][262] , \labels[0][261] , \labels[0][260] , 
	\labels[0][259] , \labels[0][258] , \labels[0][257] , 
	\labels[0][256] , \labels[0][255] , \labels[0][254] , 
	\labels[0][253] , \labels[0][252] , \labels[0][251] , 
	\labels[0][250] , \labels[0][249] , \labels[0][248] , 
	\labels[0][247] , \labels[0][246] , \labels[0][245] , 
	\labels[0][244] , \labels[0][243] , \labels[0][242] , 
	\labels[0][241] , \labels[0][240] , \labels[0][239] , 
	\labels[0][238] , \labels[0][237] , \labels[0][236] , 
	\labels[0][235] , \labels[0][234] , \labels[0][233] , 
	\labels[0][232] , \labels[0][231] , \labels[0][230] , 
	\labels[0][229] , \labels[0][228] , \labels[0][227] , 
	\labels[0][226] , \labels[0][225] , \labels[0][224] , 
	\labels[0][223] , \labels[0][222] , \labels[0][221] , 
	\labels[0][220] , \labels[0][219] , \labels[0][218] , 
	\labels[0][217] , \labels[0][216] , \labels[0][215] , 
	\labels[0][214] , \labels[0][213] , \labels[0][212] , 
	\labels[0][211] , \labels[0][210] , \labels[0][209] , 
	\labels[0][208] , \labels[0][207] , \labels[0][206] , 
	\labels[0][205] , \labels[0][204] , \labels[0][203] , 
	\labels[0][202] , \labels[0][201] , \labels[0][200] , 
	\labels[0][199] , \labels[0][198] , \labels[0][197] , 
	\labels[0][196] , \labels[0][195] , \labels[0][194] , 
	\labels[0][193] , \labels[0][192] , \labels[0][191] , 
	\labels[0][190] , \labels[0][189] , \labels[0][188] , 
	\labels[0][187] , \labels[0][186] , \labels[0][185] , 
	\labels[0][184] , \labels[0][183] , \labels[0][182] , 
	\labels[0][181] , \labels[0][180] , \labels[0][179] , 
	\labels[0][178] , \labels[0][177] , \labels[0][176] , 
	\labels[0][175] , \labels[0][174] , \labels[0][173] , 
	\labels[0][172] , \labels[0][171] , \labels[0][170] , 
	\labels[0][169] , \labels[0][168] , \labels[0][167] , 
	\labels[0][166] , \labels[0][165] , \labels[0][164] , 
	\labels[0][163] , \labels[0][162] , \labels[0][161] , 
	\labels[0][160] , \labels[0][159] , \labels[0][158] , 
	\labels[0][157] , \labels[0][156] , \labels[0][155] , 
	\labels[0][154] , \labels[0][153] , \labels[0][152] , 
	\labels[0][151] , \labels[0][150] , \labels[0][149] , 
	\labels[0][148] , \labels[0][147] , \labels[0][146] , 
	\labels[0][145] , \labels[0][144] , \labels[0][143] , 
	\labels[0][142] , \labels[0][141] , \labels[0][140] , 
	\labels[0][139] , \labels[0][138] , \labels[0][137] , 
	\labels[0][136] , \labels[0][135] , \labels[0][134] , 
	\labels[0][133] , \labels[0][132] , \labels[0][131] , 
	\labels[0][130] , \labels[0][129] , \labels[0][128] , 
	\labels[0][127] , \labels[0][126] , \labels[0][125] , 
	\labels[0][124] , \labels[0][123] , \labels[0][122] , 
	\labels[0][121] , \labels[0][120] , \labels[0][119] , 
	\labels[0][118] , \labels[0][117] , \labels[0][116] , 
	\labels[0][115] , \labels[0][114] , \labels[0][113] , 
	\labels[0][112] , \labels[0][111] , \labels[0][110] , 
	\labels[0][109] , \labels[0][108] , \labels[0][107] , 
	\labels[0][106] , \labels[0][105] , \labels[0][104] , 
	\labels[0][103] , \labels[0][102] , \labels[0][101] , 
	\labels[0][100] , \labels[0][99] , \labels[0][98] , \labels[0][97] , 
	\labels[0][96] , \labels[0][95] , \labels[0][94] , \labels[0][93] , 
	\labels[0][92] , \labels[0][91] , \labels[0][90] , \labels[0][89] , 
	\labels[0][88] , \labels[0][87] , \labels[0][86] , \labels[0][85] , 
	\labels[0][84] , \labels[0][83] , \labels[0][82] , \labels[0][81] , 
	\labels[0][80] , \labels[0][79] , \labels[0][78] , \labels[0][77] , 
	\labels[0][76] , \labels[0][75] , \labels[0][74] , \labels[0][73] , 
	\labels[0][72] , \labels[0][71] , \labels[0][70] , \labels[0][69] , 
	\labels[0][68] , \labels[0][67] , \labels[0][66] , \labels[0][65] , 
	\labels[0][64] , \labels[0][63] , \labels[0][62] , \labels[0][61] , 
	\labels[0][60] , \labels[0][59] , \labels[0][58] , \labels[0][57] , 
	\labels[0][56] , \labels[0][55] , \labels[0][54] , \labels[0][53] , 
	\labels[0][52] , \labels[0][51] , \labels[0][50] , \labels[0][49] , 
	\labels[0][48] , \labels[0][47] , \labels[0][46] , \labels[0][45] , 
	\labels[0][44] , \labels[0][43] , \labels[0][42] , \labels[0][41] , 
	\labels[0][40] , \labels[0][39] , \labels[0][38] , \labels[0][37] , 
	\labels[0][36] , \labels[0][35] , \labels[0][34] , \labels[0][33] , 
	\labels[0][32] , \labels[0][31] , \labels[0][30] , \labels[0][29] , 
	\labels[0][28] , \labels[0][27] , \labels[0][26] , \labels[0][25] , 
	\labels[0][24] , \labels[0][23] , \labels[0][22] , \labels[0][21] , 
	\labels[0][20] , \labels[0][19] , \labels[0][18] , \labels[0][17] , 
	\labels[0][16] , \labels[0][15] , \labels[0][14] , \labels[0][13] , 
	\labels[0][12] , \labels[0][11] , \labels[0][10] , \labels[0][9] , 
	\labels[0][8] , \labels[0][7] , \labels[0][6] , \labels[0][5] , 
	\labels[0][4] , \labels[0][3] , \labels[0][2] , \labels[0][1] , 
	\labels[0][0] }), .kme_internal_out( kme_internal_out[70:0]), 
	.kme_internal_out_valid( kme_internal_out_valid), 
	.gcm_cmd_in_stall( gcm_cmd_in_stall), .gcm_tag_data_in_stall( 
	gcm_tag_data_in_stall), .upsizer_inspector_stall( 
	upsizer_inspector_stall), .keyfilter_cmd_in_stall( 
	keyfilter_cmd_in_stall), .kdfstream_cmd_in_stall( 
	kdfstream_cmd_in_stall), .kdf_cmd_in_stall( kdf_cmd_in_stall), 
	.tlv_sb_data_in_stall( tlv_sb_data_in_stall));
cr_kme_kop_upsizer_x2_xcm72 upsizer ( .upsizer_in_stall( 
	upsizer_inspector_stall), .upsizer_out_valid( upsizer_gcm_valid), 
	.upsizer_out_eof( upsizer_gcm_eof), .upsizer_out_data( 
	upsizer_gcm_data[127:0]), .clk( clk), .rst_n( rst_n), 
	.in_upsizer_valid( inspector_upsizer_valid), .in_upsizer_eof( 
	inspector_upsizer_eof), .in_upsizer_data( 
	inspector_upsizer_data[63:0]), .out_upsizer_stall( gcm_upsizer_stall));
cr_kme_kop_gcm gcm ( .set_gcm_tag_fail_int( set_gcm_tag_fail_int), 
	.gcm_cmdfifo_ack( gcm_cmdfifo_ack), .gcm_upsizer_stall( 
	gcm_upsizer_stall), .gcm_tag_data_out_ack( gcm_tag_data_out_ack), 
	.gcm_kdf_valid( gcm_kdf_valid), .gcm_kdf_eof( gcm_kdf_eof), 
	.gcm_kdf_data( gcm_kdf_data[127:0]), .gcm_status_data_in_valid( 
	gcm_status_data_in_valid), .gcm_status_data_in( 
	_zy_simnet_gcm_status_data_in_5_w$), .clk( clk), .rst_n( rst_n), 
	.cmdfifo_gcm_valid( cmdfifo_gcm_valid), .cmdfifo_gcm_cmd( 
	cmdfifo_gcm_cmd[610:0]), .upsizer_gcm_valid( upsizer_gcm_valid), 
	.upsizer_gcm_eof( upsizer_gcm_eof), .upsizer_gcm_data( 
	upsizer_gcm_data[127:0]), .gcm_tag_data_out( 
	gcm_tag_data_out[95:0]), .gcm_tag_data_out_valid( 
	gcm_tag_data_out_valid), .kdf_gcm_stall( kdf_gcm_stall), 
	.gcm_status_data_in_stall( gcm_status_data_in_stall));
cr_kme_kop_kdf kdf ( .keyfilter_cmdfifo_ack( keyfilter_cmdfifo_ack), 
	.kdf_cmdfifo_ack( kdf_cmdfifo_ack), .kdfstream_cmdfifo_ack( 
	kdfstream_cmdfifo_ack), .kdf_gcm_stall( kdf_gcm_stall), 
	.kdf_keybuilder_data( kdf_keybuilder_data[63:0]), 
	.kdf_keybuilder_valid( kdf_keybuilder_valid), .clk( clk), .rst_n( 
	rst_n), .scan_en( scan_en), .scan_mode( scan_mode), .scan_rst_n( 
	scan_rst_n), .labels( { \labels[7][271] , \labels[7][270] , 
	\labels[7][269] , \labels[7][268] , \labels[7][267] , 
	\labels[7][266] , \labels[7][265] , \labels[7][264] , 
	\labels[7][263] , \labels[7][262] , \labels[7][261] , 
	\labels[7][260] , \labels[7][259] , \labels[7][258] , 
	\labels[7][257] , \labels[7][256] , \labels[7][255] , 
	\labels[7][254] , \labels[7][253] , \labels[7][252] , 
	\labels[7][251] , \labels[7][250] , \labels[7][249] , 
	\labels[7][248] , \labels[7][247] , \labels[7][246] , 
	\labels[7][245] , \labels[7][244] , \labels[7][243] , 
	\labels[7][242] , \labels[7][241] , \labels[7][240] , 
	\labels[7][239] , \labels[7][238] , \labels[7][237] , 
	\labels[7][236] , \labels[7][235] , \labels[7][234] , 
	\labels[7][233] , \labels[7][232] , \labels[7][231] , 
	\labels[7][230] , \labels[7][229] , \labels[7][228] , 
	\labels[7][227] , \labels[7][226] , \labels[7][225] , 
	\labels[7][224] , \labels[7][223] , \labels[7][222] , 
	\labels[7][221] , \labels[7][220] , \labels[7][219] , 
	\labels[7][218] , \labels[7][217] , \labels[7][216] , 
	\labels[7][215] , \labels[7][214] , \labels[7][213] , 
	\labels[7][212] , \labels[7][211] , \labels[7][210] , 
	\labels[7][209] , \labels[7][208] , \labels[7][207] , 
	\labels[7][206] , \labels[7][205] , \labels[7][204] , 
	\labels[7][203] , \labels[7][202] , \labels[7][201] , 
	\labels[7][200] , \labels[7][199] , \labels[7][198] , 
	\labels[7][197] , \labels[7][196] , \labels[7][195] , 
	\labels[7][194] , \labels[7][193] , \labels[7][192] , 
	\labels[7][191] , \labels[7][190] , \labels[7][189] , 
	\labels[7][188] , \labels[7][187] , \labels[7][186] , 
	\labels[7][185] , \labels[7][184] , \labels[7][183] , 
	\labels[7][182] , \labels[7][181] , \labels[7][180] , 
	\labels[7][179] , \labels[7][178] , \labels[7][177] , 
	\labels[7][176] , \labels[7][175] , \labels[7][174] , 
	\labels[7][173] , \labels[7][172] , \labels[7][171] , 
	\labels[7][170] , \labels[7][169] , \labels[7][168] , 
	\labels[7][167] , \labels[7][166] , \labels[7][165] , 
	\labels[7][164] , \labels[7][163] , \labels[7][162] , 
	\labels[7][161] , \labels[7][160] , \labels[7][159] , 
	\labels[7][158] , \labels[7][157] , \labels[7][156] , 
	\labels[7][155] , \labels[7][154] , \labels[7][153] , 
	\labels[7][152] , \labels[7][151] , \labels[7][150] , 
	\labels[7][149] , \labels[7][148] , \labels[7][147] , 
	\labels[7][146] , \labels[7][145] , \labels[7][144] , 
	\labels[7][143] , \labels[7][142] , \labels[7][141] , 
	\labels[7][140] , \labels[7][139] , \labels[7][138] , 
	\labels[7][137] , \labels[7][136] , \labels[7][135] , 
	\labels[7][134] , \labels[7][133] , \labels[7][132] , 
	\labels[7][131] , \labels[7][130] , \labels[7][129] , 
	\labels[7][128] , \labels[7][127] , \labels[7][126] , 
	\labels[7][125] , \labels[7][124] , \labels[7][123] , 
	\labels[7][122] , \labels[7][121] , \labels[7][120] , 
	\labels[7][119] , \labels[7][118] , \labels[7][117] , 
	\labels[7][116] , \labels[7][115] , \labels[7][114] , 
	\labels[7][113] , \labels[7][112] , \labels[7][111] , 
	\labels[7][110] , \labels[7][109] , \labels[7][108] , 
	\labels[7][107] , \labels[7][106] , \labels[7][105] , 
	\labels[7][104] , \labels[7][103] , \labels[7][102] , 
	\labels[7][101] , \labels[7][100] , \labels[7][99] , \labels[7][98] , 
	\labels[7][97] , \labels[7][96] , \labels[7][95] , \labels[7][94] , 
	\labels[7][93] , \labels[7][92] , \labels[7][91] , \labels[7][90] , 
	\labels[7][89] , \labels[7][88] , \labels[7][87] , \labels[7][86] , 
	\labels[7][85] , \labels[7][84] , \labels[7][83] , \labels[7][82] , 
	\labels[7][81] , \labels[7][80] , \labels[7][79] , \labels[7][78] , 
	\labels[7][77] , \labels[7][76] , \labels[7][75] , \labels[7][74] , 
	\labels[7][73] , \labels[7][72] , \labels[7][71] , \labels[7][70] , 
	\labels[7][69] , \labels[7][68] , \labels[7][67] , \labels[7][66] , 
	\labels[7][65] , \labels[7][64] , \labels[7][63] , \labels[7][62] , 
	\labels[7][61] , \labels[7][60] , \labels[7][59] , \labels[7][58] , 
	\labels[7][57] , \labels[7][56] , \labels[7][55] , \labels[7][54] , 
	\labels[7][53] , \labels[7][52] , \labels[7][51] , \labels[7][50] , 
	\labels[7][49] , \labels[7][48] , \labels[7][47] , \labels[7][46] , 
	\labels[7][45] , \labels[7][44] , \labels[7][43] , \labels[7][42] , 
	\labels[7][41] , \labels[7][40] , \labels[7][39] , \labels[7][38] , 
	\labels[7][37] , \labels[7][36] , \labels[7][35] , \labels[7][34] , 
	\labels[7][33] , \labels[7][32] , \labels[7][31] , \labels[7][30] , 
	\labels[7][29] , \labels[7][28] , \labels[7][27] , \labels[7][26] , 
	\labels[7][25] , \labels[7][24] , \labels[7][23] , \labels[7][22] , 
	\labels[7][21] , \labels[7][20] , \labels[7][19] , \labels[7][18] , 
	\labels[7][17] , \labels[7][16] , \labels[7][15] , \labels[7][14] , 
	\labels[7][13] , \labels[7][12] , \labels[7][11] , \labels[7][10] , 
	\labels[7][9] , \labels[7][8] , \labels[7][7] , \labels[7][6] , 
	\labels[7][5] , \labels[7][4] , \labels[7][3] , \labels[7][2] , 
	\labels[7][1] , \labels[7][0] , \labels[6][271] , \labels[6][270] , 
	\labels[6][269] , \labels[6][268] , \labels[6][267] , 
	\labels[6][266] , \labels[6][265] , \labels[6][264] , 
	\labels[6][263] , \labels[6][262] , \labels[6][261] , 
	\labels[6][260] , \labels[6][259] , \labels[6][258] , 
	\labels[6][257] , \labels[6][256] , \labels[6][255] , 
	\labels[6][254] , \labels[6][253] , \labels[6][252] , 
	\labels[6][251] , \labels[6][250] , \labels[6][249] , 
	\labels[6][248] , \labels[6][247] , \labels[6][246] , 
	\labels[6][245] , \labels[6][244] , \labels[6][243] , 
	\labels[6][242] , \labels[6][241] , \labels[6][240] , 
	\labels[6][239] , \labels[6][238] , \labels[6][237] , 
	\labels[6][236] , \labels[6][235] , \labels[6][234] , 
	\labels[6][233] , \labels[6][232] , \labels[6][231] , 
	\labels[6][230] , \labels[6][229] , \labels[6][228] , 
	\labels[6][227] , \labels[6][226] , \labels[6][225] , 
	\labels[6][224] , \labels[6][223] , \labels[6][222] , 
	\labels[6][221] , \labels[6][220] , \labels[6][219] , 
	\labels[6][218] , \labels[6][217] , \labels[6][216] , 
	\labels[6][215] , \labels[6][214] , \labels[6][213] , 
	\labels[6][212] , \labels[6][211] , \labels[6][210] , 
	\labels[6][209] , \labels[6][208] , \labels[6][207] , 
	\labels[6][206] , \labels[6][205] , \labels[6][204] , 
	\labels[6][203] , \labels[6][202] , \labels[6][201] , 
	\labels[6][200] , \labels[6][199] , \labels[6][198] , 
	\labels[6][197] , \labels[6][196] , \labels[6][195] , 
	\labels[6][194] , \labels[6][193] , \labels[6][192] , 
	\labels[6][191] , \labels[6][190] , \labels[6][189] , 
	\labels[6][188] , \labels[6][187] , \labels[6][186] , 
	\labels[6][185] , \labels[6][184] , \labels[6][183] , 
	\labels[6][182] , \labels[6][181] , \labels[6][180] , 
	\labels[6][179] , \labels[6][178] , \labels[6][177] , 
	\labels[6][176] , \labels[6][175] , \labels[6][174] , 
	\labels[6][173] , \labels[6][172] , \labels[6][171] , 
	\labels[6][170] , \labels[6][169] , \labels[6][168] , 
	\labels[6][167] , \labels[6][166] , \labels[6][165] , 
	\labels[6][164] , \labels[6][163] , \labels[6][162] , 
	\labels[6][161] , \labels[6][160] , \labels[6][159] , 
	\labels[6][158] , \labels[6][157] , \labels[6][156] , 
	\labels[6][155] , \labels[6][154] , \labels[6][153] , 
	\labels[6][152] , \labels[6][151] , \labels[6][150] , 
	\labels[6][149] , \labels[6][148] , \labels[6][147] , 
	\labels[6][146] , \labels[6][145] , \labels[6][144] , 
	\labels[6][143] , \labels[6][142] , \labels[6][141] , 
	\labels[6][140] , \labels[6][139] , \labels[6][138] , 
	\labels[6][137] , \labels[6][136] , \labels[6][135] , 
	\labels[6][134] , \labels[6][133] , \labels[6][132] , 
	\labels[6][131] , \labels[6][130] , \labels[6][129] , 
	\labels[6][128] , \labels[6][127] , \labels[6][126] , 
	\labels[6][125] , \labels[6][124] , \labels[6][123] , 
	\labels[6][122] , \labels[6][121] , \labels[6][120] , 
	\labels[6][119] , \labels[6][118] , \labels[6][117] , 
	\labels[6][116] , \labels[6][115] , \labels[6][114] , 
	\labels[6][113] , \labels[6][112] , \labels[6][111] , 
	\labels[6][110] , \labels[6][109] , \labels[6][108] , 
	\labels[6][107] , \labels[6][106] , \labels[6][105] , 
	\labels[6][104] , \labels[6][103] , \labels[6][102] , 
	\labels[6][101] , \labels[6][100] , \labels[6][99] , \labels[6][98] , 
	\labels[6][97] , \labels[6][96] , \labels[6][95] , \labels[6][94] , 
	\labels[6][93] , \labels[6][92] , \labels[6][91] , \labels[6][90] , 
	\labels[6][89] , \labels[6][88] , \labels[6][87] , \labels[6][86] , 
	\labels[6][85] , \labels[6][84] , \labels[6][83] , \labels[6][82] , 
	\labels[6][81] , \labels[6][80] , \labels[6][79] , \labels[6][78] , 
	\labels[6][77] , \labels[6][76] , \labels[6][75] , \labels[6][74] , 
	\labels[6][73] , \labels[6][72] , \labels[6][71] , \labels[6][70] , 
	\labels[6][69] , \labels[6][68] , \labels[6][67] , \labels[6][66] , 
	\labels[6][65] , \labels[6][64] , \labels[6][63] , \labels[6][62] , 
	\labels[6][61] , \labels[6][60] , \labels[6][59] , \labels[6][58] , 
	\labels[6][57] , \labels[6][56] , \labels[6][55] , \labels[6][54] , 
	\labels[6][53] , \labels[6][52] , \labels[6][51] , \labels[6][50] , 
	\labels[6][49] , \labels[6][48] , \labels[6][47] , \labels[6][46] , 
	\labels[6][45] , \labels[6][44] , \labels[6][43] , \labels[6][42] , 
	\labels[6][41] , \labels[6][40] , \labels[6][39] , \labels[6][38] , 
	\labels[6][37] , \labels[6][36] , \labels[6][35] , \labels[6][34] , 
	\labels[6][33] , \labels[6][32] , \labels[6][31] , \labels[6][30] , 
	\labels[6][29] , \labels[6][28] , \labels[6][27] , \labels[6][26] , 
	\labels[6][25] , \labels[6][24] , \labels[6][23] , \labels[6][22] , 
	\labels[6][21] , \labels[6][20] , \labels[6][19] , \labels[6][18] , 
	\labels[6][17] , \labels[6][16] , \labels[6][15] , \labels[6][14] , 
	\labels[6][13] , \labels[6][12] , \labels[6][11] , \labels[6][10] , 
	\labels[6][9] , \labels[6][8] , \labels[6][7] , \labels[6][6] , 
	\labels[6][5] , \labels[6][4] , \labels[6][3] , \labels[6][2] , 
	\labels[6][1] , \labels[6][0] , \labels[5][271] , \labels[5][270] , 
	\labels[5][269] , \labels[5][268] , \labels[5][267] , 
	\labels[5][266] , \labels[5][265] , \labels[5][264] , 
	\labels[5][263] , \labels[5][262] , \labels[5][261] , 
	\labels[5][260] , \labels[5][259] , \labels[5][258] , 
	\labels[5][257] , \labels[5][256] , \labels[5][255] , 
	\labels[5][254] , \labels[5][253] , \labels[5][252] , 
	\labels[5][251] , \labels[5][250] , \labels[5][249] , 
	\labels[5][248] , \labels[5][247] , \labels[5][246] , 
	\labels[5][245] , \labels[5][244] , \labels[5][243] , 
	\labels[5][242] , \labels[5][241] , \labels[5][240] , 
	\labels[5][239] , \labels[5][238] , \labels[5][237] , 
	\labels[5][236] , \labels[5][235] , \labels[5][234] , 
	\labels[5][233] , \labels[5][232] , \labels[5][231] , 
	\labels[5][230] , \labels[5][229] , \labels[5][228] , 
	\labels[5][227] , \labels[5][226] , \labels[5][225] , 
	\labels[5][224] , \labels[5][223] , \labels[5][222] , 
	\labels[5][221] , \labels[5][220] , \labels[5][219] , 
	\labels[5][218] , \labels[5][217] , \labels[5][216] , 
	\labels[5][215] , \labels[5][214] , \labels[5][213] , 
	\labels[5][212] , \labels[5][211] , \labels[5][210] , 
	\labels[5][209] , \labels[5][208] , \labels[5][207] , 
	\labels[5][206] , \labels[5][205] , \labels[5][204] , 
	\labels[5][203] , \labels[5][202] , \labels[5][201] , 
	\labels[5][200] , \labels[5][199] , \labels[5][198] , 
	\labels[5][197] , \labels[5][196] , \labels[5][195] , 
	\labels[5][194] , \labels[5][193] , \labels[5][192] , 
	\labels[5][191] , \labels[5][190] , \labels[5][189] , 
	\labels[5][188] , \labels[5][187] , \labels[5][186] , 
	\labels[5][185] , \labels[5][184] , \labels[5][183] , 
	\labels[5][182] , \labels[5][181] , \labels[5][180] , 
	\labels[5][179] , \labels[5][178] , \labels[5][177] , 
	\labels[5][176] , \labels[5][175] , \labels[5][174] , 
	\labels[5][173] , \labels[5][172] , \labels[5][171] , 
	\labels[5][170] , \labels[5][169] , \labels[5][168] , 
	\labels[5][167] , \labels[5][166] , \labels[5][165] , 
	\labels[5][164] , \labels[5][163] , \labels[5][162] , 
	\labels[5][161] , \labels[5][160] , \labels[5][159] , 
	\labels[5][158] , \labels[5][157] , \labels[5][156] , 
	\labels[5][155] , \labels[5][154] , \labels[5][153] , 
	\labels[5][152] , \labels[5][151] , \labels[5][150] , 
	\labels[5][149] , \labels[5][148] , \labels[5][147] , 
	\labels[5][146] , \labels[5][145] , \labels[5][144] , 
	\labels[5][143] , \labels[5][142] , \labels[5][141] , 
	\labels[5][140] , \labels[5][139] , \labels[5][138] , 
	\labels[5][137] , \labels[5][136] , \labels[5][135] , 
	\labels[5][134] , \labels[5][133] , \labels[5][132] , 
	\labels[5][131] , \labels[5][130] , \labels[5][129] , 
	\labels[5][128] , \labels[5][127] , \labels[5][126] , 
	\labels[5][125] , \labels[5][124] , \labels[5][123] , 
	\labels[5][122] , \labels[5][121] , \labels[5][120] , 
	\labels[5][119] , \labels[5][118] , \labels[5][117] , 
	\labels[5][116] , \labels[5][115] , \labels[5][114] , 
	\labels[5][113] , \labels[5][112] , \labels[5][111] , 
	\labels[5][110] , \labels[5][109] , \labels[5][108] , 
	\labels[5][107] , \labels[5][106] , \labels[5][105] , 
	\labels[5][104] , \labels[5][103] , \labels[5][102] , 
	\labels[5][101] , \labels[5][100] , \labels[5][99] , \labels[5][98] , 
	\labels[5][97] , \labels[5][96] , \labels[5][95] , \labels[5][94] , 
	\labels[5][93] , \labels[5][92] , \labels[5][91] , \labels[5][90] , 
	\labels[5][89] , \labels[5][88] , \labels[5][87] , \labels[5][86] , 
	\labels[5][85] , \labels[5][84] , \labels[5][83] , \labels[5][82] , 
	\labels[5][81] , \labels[5][80] , \labels[5][79] , \labels[5][78] , 
	\labels[5][77] , \labels[5][76] , \labels[5][75] , \labels[5][74] , 
	\labels[5][73] , \labels[5][72] , \labels[5][71] , \labels[5][70] , 
	\labels[5][69] , \labels[5][68] , \labels[5][67] , \labels[5][66] , 
	\labels[5][65] , \labels[5][64] , \labels[5][63] , \labels[5][62] , 
	\labels[5][61] , \labels[5][60] , \labels[5][59] , \labels[5][58] , 
	\labels[5][57] , \labels[5][56] , \labels[5][55] , \labels[5][54] , 
	\labels[5][53] , \labels[5][52] , \labels[5][51] , \labels[5][50] , 
	\labels[5][49] , \labels[5][48] , \labels[5][47] , \labels[5][46] , 
	\labels[5][45] , \labels[5][44] , \labels[5][43] , \labels[5][42] , 
	\labels[5][41] , \labels[5][40] , \labels[5][39] , \labels[5][38] , 
	\labels[5][37] , \labels[5][36] , \labels[5][35] , \labels[5][34] , 
	\labels[5][33] , \labels[5][32] , \labels[5][31] , \labels[5][30] , 
	\labels[5][29] , \labels[5][28] , \labels[5][27] , \labels[5][26] , 
	\labels[5][25] , \labels[5][24] , \labels[5][23] , \labels[5][22] , 
	\labels[5][21] , \labels[5][20] , \labels[5][19] , \labels[5][18] , 
	\labels[5][17] , \labels[5][16] , \labels[5][15] , \labels[5][14] , 
	\labels[5][13] , \labels[5][12] , \labels[5][11] , \labels[5][10] , 
	\labels[5][9] , \labels[5][8] , \labels[5][7] , \labels[5][6] , 
	\labels[5][5] , \labels[5][4] , \labels[5][3] , \labels[5][2] , 
	\labels[5][1] , \labels[5][0] , \labels[4][271] , \labels[4][270] , 
	\labels[4][269] , \labels[4][268] , \labels[4][267] , 
	\labels[4][266] , \labels[4][265] , \labels[4][264] , 
	\labels[4][263] , \labels[4][262] , \labels[4][261] , 
	\labels[4][260] , \labels[4][259] , \labels[4][258] , 
	\labels[4][257] , \labels[4][256] , \labels[4][255] , 
	\labels[4][254] , \labels[4][253] , \labels[4][252] , 
	\labels[4][251] , \labels[4][250] , \labels[4][249] , 
	\labels[4][248] , \labels[4][247] , \labels[4][246] , 
	\labels[4][245] , \labels[4][244] , \labels[4][243] , 
	\labels[4][242] , \labels[4][241] , \labels[4][240] , 
	\labels[4][239] , \labels[4][238] , \labels[4][237] , 
	\labels[4][236] , \labels[4][235] , \labels[4][234] , 
	\labels[4][233] , \labels[4][232] , \labels[4][231] , 
	\labels[4][230] , \labels[4][229] , \labels[4][228] , 
	\labels[4][227] , \labels[4][226] , \labels[4][225] , 
	\labels[4][224] , \labels[4][223] , \labels[4][222] , 
	\labels[4][221] , \labels[4][220] , \labels[4][219] , 
	\labels[4][218] , \labels[4][217] , \labels[4][216] , 
	\labels[4][215] , \labels[4][214] , \labels[4][213] , 
	\labels[4][212] , \labels[4][211] , \labels[4][210] , 
	\labels[4][209] , \labels[4][208] , \labels[4][207] , 
	\labels[4][206] , \labels[4][205] , \labels[4][204] , 
	\labels[4][203] , \labels[4][202] , \labels[4][201] , 
	\labels[4][200] , \labels[4][199] , \labels[4][198] , 
	\labels[4][197] , \labels[4][196] , \labels[4][195] , 
	\labels[4][194] , \labels[4][193] , \labels[4][192] , 
	\labels[4][191] , \labels[4][190] , \labels[4][189] , 
	\labels[4][188] , \labels[4][187] , \labels[4][186] , 
	\labels[4][185] , \labels[4][184] , \labels[4][183] , 
	\labels[4][182] , \labels[4][181] , \labels[4][180] , 
	\labels[4][179] , \labels[4][178] , \labels[4][177] , 
	\labels[4][176] , \labels[4][175] , \labels[4][174] , 
	\labels[4][173] , \labels[4][172] , \labels[4][171] , 
	\labels[4][170] , \labels[4][169] , \labels[4][168] , 
	\labels[4][167] , \labels[4][166] , \labels[4][165] , 
	\labels[4][164] , \labels[4][163] , \labels[4][162] , 
	\labels[4][161] , \labels[4][160] , \labels[4][159] , 
	\labels[4][158] , \labels[4][157] , \labels[4][156] , 
	\labels[4][155] , \labels[4][154] , \labels[4][153] , 
	\labels[4][152] , \labels[4][151] , \labels[4][150] , 
	\labels[4][149] , \labels[4][148] , \labels[4][147] , 
	\labels[4][146] , \labels[4][145] , \labels[4][144] , 
	\labels[4][143] , \labels[4][142] , \labels[4][141] , 
	\labels[4][140] , \labels[4][139] , \labels[4][138] , 
	\labels[4][137] , \labels[4][136] , \labels[4][135] , 
	\labels[4][134] , \labels[4][133] , \labels[4][132] , 
	\labels[4][131] , \labels[4][130] , \labels[4][129] , 
	\labels[4][128] , \labels[4][127] , \labels[4][126] , 
	\labels[4][125] , \labels[4][124] , \labels[4][123] , 
	\labels[4][122] , \labels[4][121] , \labels[4][120] , 
	\labels[4][119] , \labels[4][118] , \labels[4][117] , 
	\labels[4][116] , \labels[4][115] , \labels[4][114] , 
	\labels[4][113] , \labels[4][112] , \labels[4][111] , 
	\labels[4][110] , \labels[4][109] , \labels[4][108] , 
	\labels[4][107] , \labels[4][106] , \labels[4][105] , 
	\labels[4][104] , \labels[4][103] , \labels[4][102] , 
	\labels[4][101] , \labels[4][100] , \labels[4][99] , \labels[4][98] , 
	\labels[4][97] , \labels[4][96] , \labels[4][95] , \labels[4][94] , 
	\labels[4][93] , \labels[4][92] , \labels[4][91] , \labels[4][90] , 
	\labels[4][89] , \labels[4][88] , \labels[4][87] , \labels[4][86] , 
	\labels[4][85] , \labels[4][84] , \labels[4][83] , \labels[4][82] , 
	\labels[4][81] , \labels[4][80] , \labels[4][79] , \labels[4][78] , 
	\labels[4][77] , \labels[4][76] , \labels[4][75] , \labels[4][74] , 
	\labels[4][73] , \labels[4][72] , \labels[4][71] , \labels[4][70] , 
	\labels[4][69] , \labels[4][68] , \labels[4][67] , \labels[4][66] , 
	\labels[4][65] , \labels[4][64] , \labels[4][63] , \labels[4][62] , 
	\labels[4][61] , \labels[4][60] , \labels[4][59] , \labels[4][58] , 
	\labels[4][57] , \labels[4][56] , \labels[4][55] , \labels[4][54] , 
	\labels[4][53] , \labels[4][52] , \labels[4][51] , \labels[4][50] , 
	\labels[4][49] , \labels[4][48] , \labels[4][47] , \labels[4][46] , 
	\labels[4][45] , \labels[4][44] , \labels[4][43] , \labels[4][42] , 
	\labels[4][41] , \labels[4][40] , \labels[4][39] , \labels[4][38] , 
	\labels[4][37] , \labels[4][36] , \labels[4][35] , \labels[4][34] , 
	\labels[4][33] , \labels[4][32] , \labels[4][31] , \labels[4][30] , 
	\labels[4][29] , \labels[4][28] , \labels[4][27] , \labels[4][26] , 
	\labels[4][25] , \labels[4][24] , \labels[4][23] , \labels[4][22] , 
	\labels[4][21] , \labels[4][20] , \labels[4][19] , \labels[4][18] , 
	\labels[4][17] , \labels[4][16] , \labels[4][15] , \labels[4][14] , 
	\labels[4][13] , \labels[4][12] , \labels[4][11] , \labels[4][10] , 
	\labels[4][9] , \labels[4][8] , \labels[4][7] , \labels[4][6] , 
	\labels[4][5] , \labels[4][4] , \labels[4][3] , \labels[4][2] , 
	\labels[4][1] , \labels[4][0] , \labels[3][271] , \labels[3][270] , 
	\labels[3][269] , \labels[3][268] , \labels[3][267] , 
	\labels[3][266] , \labels[3][265] , \labels[3][264] , 
	\labels[3][263] , \labels[3][262] , \labels[3][261] , 
	\labels[3][260] , \labels[3][259] , \labels[3][258] , 
	\labels[3][257] , \labels[3][256] , \labels[3][255] , 
	\labels[3][254] , \labels[3][253] , \labels[3][252] , 
	\labels[3][251] , \labels[3][250] , \labels[3][249] , 
	\labels[3][248] , \labels[3][247] , \labels[3][246] , 
	\labels[3][245] , \labels[3][244] , \labels[3][243] , 
	\labels[3][242] , \labels[3][241] , \labels[3][240] , 
	\labels[3][239] , \labels[3][238] , \labels[3][237] , 
	\labels[3][236] , \labels[3][235] , \labels[3][234] , 
	\labels[3][233] , \labels[3][232] , \labels[3][231] , 
	\labels[3][230] , \labels[3][229] , \labels[3][228] , 
	\labels[3][227] , \labels[3][226] , \labels[3][225] , 
	\labels[3][224] , \labels[3][223] , \labels[3][222] , 
	\labels[3][221] , \labels[3][220] , \labels[3][219] , 
	\labels[3][218] , \labels[3][217] , \labels[3][216] , 
	\labels[3][215] , \labels[3][214] , \labels[3][213] , 
	\labels[3][212] , \labels[3][211] , \labels[3][210] , 
	\labels[3][209] , \labels[3][208] , \labels[3][207] , 
	\labels[3][206] , \labels[3][205] , \labels[3][204] , 
	\labels[3][203] , \labels[3][202] , \labels[3][201] , 
	\labels[3][200] , \labels[3][199] , \labels[3][198] , 
	\labels[3][197] , \labels[3][196] , \labels[3][195] , 
	\labels[3][194] , \labels[3][193] , \labels[3][192] , 
	\labels[3][191] , \labels[3][190] , \labels[3][189] , 
	\labels[3][188] , \labels[3][187] , \labels[3][186] , 
	\labels[3][185] , \labels[3][184] , \labels[3][183] , 
	\labels[3][182] , \labels[3][181] , \labels[3][180] , 
	\labels[3][179] , \labels[3][178] , \labels[3][177] , 
	\labels[3][176] , \labels[3][175] , \labels[3][174] , 
	\labels[3][173] , \labels[3][172] , \labels[3][171] , 
	\labels[3][170] , \labels[3][169] , \labels[3][168] , 
	\labels[3][167] , \labels[3][166] , \labels[3][165] , 
	\labels[3][164] , \labels[3][163] , \labels[3][162] , 
	\labels[3][161] , \labels[3][160] , \labels[3][159] , 
	\labels[3][158] , \labels[3][157] , \labels[3][156] , 
	\labels[3][155] , \labels[3][154] , \labels[3][153] , 
	\labels[3][152] , \labels[3][151] , \labels[3][150] , 
	\labels[3][149] , \labels[3][148] , \labels[3][147] , 
	\labels[3][146] , \labels[3][145] , \labels[3][144] , 
	\labels[3][143] , \labels[3][142] , \labels[3][141] , 
	\labels[3][140] , \labels[3][139] , \labels[3][138] , 
	\labels[3][137] , \labels[3][136] , \labels[3][135] , 
	\labels[3][134] , \labels[3][133] , \labels[3][132] , 
	\labels[3][131] , \labels[3][130] , \labels[3][129] , 
	\labels[3][128] , \labels[3][127] , \labels[3][126] , 
	\labels[3][125] , \labels[3][124] , \labels[3][123] , 
	\labels[3][122] , \labels[3][121] , \labels[3][120] , 
	\labels[3][119] , \labels[3][118] , \labels[3][117] , 
	\labels[3][116] , \labels[3][115] , \labels[3][114] , 
	\labels[3][113] , \labels[3][112] , \labels[3][111] , 
	\labels[3][110] , \labels[3][109] , \labels[3][108] , 
	\labels[3][107] , \labels[3][106] , \labels[3][105] , 
	\labels[3][104] , \labels[3][103] , \labels[3][102] , 
	\labels[3][101] , \labels[3][100] , \labels[3][99] , \labels[3][98] , 
	\labels[3][97] , \labels[3][96] , \labels[3][95] , \labels[3][94] , 
	\labels[3][93] , \labels[3][92] , \labels[3][91] , \labels[3][90] , 
	\labels[3][89] , \labels[3][88] , \labels[3][87] , \labels[3][86] , 
	\labels[3][85] , \labels[3][84] , \labels[3][83] , \labels[3][82] , 
	\labels[3][81] , \labels[3][80] , \labels[3][79] , \labels[3][78] , 
	\labels[3][77] , \labels[3][76] , \labels[3][75] , \labels[3][74] , 
	\labels[3][73] , \labels[3][72] , \labels[3][71] , \labels[3][70] , 
	\labels[3][69] , \labels[3][68] , \labels[3][67] , \labels[3][66] , 
	\labels[3][65] , \labels[3][64] , \labels[3][63] , \labels[3][62] , 
	\labels[3][61] , \labels[3][60] , \labels[3][59] , \labels[3][58] , 
	\labels[3][57] , \labels[3][56] , \labels[3][55] , \labels[3][54] , 
	\labels[3][53] , \labels[3][52] , \labels[3][51] , \labels[3][50] , 
	\labels[3][49] , \labels[3][48] , \labels[3][47] , \labels[3][46] , 
	\labels[3][45] , \labels[3][44] , \labels[3][43] , \labels[3][42] , 
	\labels[3][41] , \labels[3][40] , \labels[3][39] , \labels[3][38] , 
	\labels[3][37] , \labels[3][36] , \labels[3][35] , \labels[3][34] , 
	\labels[3][33] , \labels[3][32] , \labels[3][31] , \labels[3][30] , 
	\labels[3][29] , \labels[3][28] , \labels[3][27] , \labels[3][26] , 
	\labels[3][25] , \labels[3][24] , \labels[3][23] , \labels[3][22] , 
	\labels[3][21] , \labels[3][20] , \labels[3][19] , \labels[3][18] , 
	\labels[3][17] , \labels[3][16] , \labels[3][15] , \labels[3][14] , 
	\labels[3][13] , \labels[3][12] , \labels[3][11] , \labels[3][10] , 
	\labels[3][9] , \labels[3][8] , \labels[3][7] , \labels[3][6] , 
	\labels[3][5] , \labels[3][4] , \labels[3][3] , \labels[3][2] , 
	\labels[3][1] , \labels[3][0] , \labels[2][271] , \labels[2][270] , 
	\labels[2][269] , \labels[2][268] , \labels[2][267] , 
	\labels[2][266] , \labels[2][265] , \labels[2][264] , 
	\labels[2][263] , \labels[2][262] , \labels[2][261] , 
	\labels[2][260] , \labels[2][259] , \labels[2][258] , 
	\labels[2][257] , \labels[2][256] , \labels[2][255] , 
	\labels[2][254] , \labels[2][253] , \labels[2][252] , 
	\labels[2][251] , \labels[2][250] , \labels[2][249] , 
	\labels[2][248] , \labels[2][247] , \labels[2][246] , 
	\labels[2][245] , \labels[2][244] , \labels[2][243] , 
	\labels[2][242] , \labels[2][241] , \labels[2][240] , 
	\labels[2][239] , \labels[2][238] , \labels[2][237] , 
	\labels[2][236] , \labels[2][235] , \labels[2][234] , 
	\labels[2][233] , \labels[2][232] , \labels[2][231] , 
	\labels[2][230] , \labels[2][229] , \labels[2][228] , 
	\labels[2][227] , \labels[2][226] , \labels[2][225] , 
	\labels[2][224] , \labels[2][223] , \labels[2][222] , 
	\labels[2][221] , \labels[2][220] , \labels[2][219] , 
	\labels[2][218] , \labels[2][217] , \labels[2][216] , 
	\labels[2][215] , \labels[2][214] , \labels[2][213] , 
	\labels[2][212] , \labels[2][211] , \labels[2][210] , 
	\labels[2][209] , \labels[2][208] , \labels[2][207] , 
	\labels[2][206] , \labels[2][205] , \labels[2][204] , 
	\labels[2][203] , \labels[2][202] , \labels[2][201] , 
	\labels[2][200] , \labels[2][199] , \labels[2][198] , 
	\labels[2][197] , \labels[2][196] , \labels[2][195] , 
	\labels[2][194] , \labels[2][193] , \labels[2][192] , 
	\labels[2][191] , \labels[2][190] , \labels[2][189] , 
	\labels[2][188] , \labels[2][187] , \labels[2][186] , 
	\labels[2][185] , \labels[2][184] , \labels[2][183] , 
	\labels[2][182] , \labels[2][181] , \labels[2][180] , 
	\labels[2][179] , \labels[2][178] , \labels[2][177] , 
	\labels[2][176] , \labels[2][175] , \labels[2][174] , 
	\labels[2][173] , \labels[2][172] , \labels[2][171] , 
	\labels[2][170] , \labels[2][169] , \labels[2][168] , 
	\labels[2][167] , \labels[2][166] , \labels[2][165] , 
	\labels[2][164] , \labels[2][163] , \labels[2][162] , 
	\labels[2][161] , \labels[2][160] , \labels[2][159] , 
	\labels[2][158] , \labels[2][157] , \labels[2][156] , 
	\labels[2][155] , \labels[2][154] , \labels[2][153] , 
	\labels[2][152] , \labels[2][151] , \labels[2][150] , 
	\labels[2][149] , \labels[2][148] , \labels[2][147] , 
	\labels[2][146] , \labels[2][145] , \labels[2][144] , 
	\labels[2][143] , \labels[2][142] , \labels[2][141] , 
	\labels[2][140] , \labels[2][139] , \labels[2][138] , 
	\labels[2][137] , \labels[2][136] , \labels[2][135] , 
	\labels[2][134] , \labels[2][133] , \labels[2][132] , 
	\labels[2][131] , \labels[2][130] , \labels[2][129] , 
	\labels[2][128] , \labels[2][127] , \labels[2][126] , 
	\labels[2][125] , \labels[2][124] , \labels[2][123] , 
	\labels[2][122] , \labels[2][121] , \labels[2][120] , 
	\labels[2][119] , \labels[2][118] , \labels[2][117] , 
	\labels[2][116] , \labels[2][115] , \labels[2][114] , 
	\labels[2][113] , \labels[2][112] , \labels[2][111] , 
	\labels[2][110] , \labels[2][109] , \labels[2][108] , 
	\labels[2][107] , \labels[2][106] , \labels[2][105] , 
	\labels[2][104] , \labels[2][103] , \labels[2][102] , 
	\labels[2][101] , \labels[2][100] , \labels[2][99] , \labels[2][98] , 
	\labels[2][97] , \labels[2][96] , \labels[2][95] , \labels[2][94] , 
	\labels[2][93] , \labels[2][92] , \labels[2][91] , \labels[2][90] , 
	\labels[2][89] , \labels[2][88] , \labels[2][87] , \labels[2][86] , 
	\labels[2][85] , \labels[2][84] , \labels[2][83] , \labels[2][82] , 
	\labels[2][81] , \labels[2][80] , \labels[2][79] , \labels[2][78] , 
	\labels[2][77] , \labels[2][76] , \labels[2][75] , \labels[2][74] , 
	\labels[2][73] , \labels[2][72] , \labels[2][71] , \labels[2][70] , 
	\labels[2][69] , \labels[2][68] , \labels[2][67] , \labels[2][66] , 
	\labels[2][65] , \labels[2][64] , \labels[2][63] , \labels[2][62] , 
	\labels[2][61] , \labels[2][60] , \labels[2][59] , \labels[2][58] , 
	\labels[2][57] , \labels[2][56] , \labels[2][55] , \labels[2][54] , 
	\labels[2][53] , \labels[2][52] , \labels[2][51] , \labels[2][50] , 
	\labels[2][49] , \labels[2][48] , \labels[2][47] , \labels[2][46] , 
	\labels[2][45] , \labels[2][44] , \labels[2][43] , \labels[2][42] , 
	\labels[2][41] , \labels[2][40] , \labels[2][39] , \labels[2][38] , 
	\labels[2][37] , \labels[2][36] , \labels[2][35] , \labels[2][34] , 
	\labels[2][33] , \labels[2][32] , \labels[2][31] , \labels[2][30] , 
	\labels[2][29] , \labels[2][28] , \labels[2][27] , \labels[2][26] , 
	\labels[2][25] , \labels[2][24] , \labels[2][23] , \labels[2][22] , 
	\labels[2][21] , \labels[2][20] , \labels[2][19] , \labels[2][18] , 
	\labels[2][17] , \labels[2][16] , \labels[2][15] , \labels[2][14] , 
	\labels[2][13] , \labels[2][12] , \labels[2][11] , \labels[2][10] , 
	\labels[2][9] , \labels[2][8] , \labels[2][7] , \labels[2][6] , 
	\labels[2][5] , \labels[2][4] , \labels[2][3] , \labels[2][2] , 
	\labels[2][1] , \labels[2][0] , \labels[1][271] , \labels[1][270] , 
	\labels[1][269] , \labels[1][268] , \labels[1][267] , 
	\labels[1][266] , \labels[1][265] , \labels[1][264] , 
	\labels[1][263] , \labels[1][262] , \labels[1][261] , 
	\labels[1][260] , \labels[1][259] , \labels[1][258] , 
	\labels[1][257] , \labels[1][256] , \labels[1][255] , 
	\labels[1][254] , \labels[1][253] , \labels[1][252] , 
	\labels[1][251] , \labels[1][250] , \labels[1][249] , 
	\labels[1][248] , \labels[1][247] , \labels[1][246] , 
	\labels[1][245] , \labels[1][244] , \labels[1][243] , 
	\labels[1][242] , \labels[1][241] , \labels[1][240] , 
	\labels[1][239] , \labels[1][238] , \labels[1][237] , 
	\labels[1][236] , \labels[1][235] , \labels[1][234] , 
	\labels[1][233] , \labels[1][232] , \labels[1][231] , 
	\labels[1][230] , \labels[1][229] , \labels[1][228] , 
	\labels[1][227] , \labels[1][226] , \labels[1][225] , 
	\labels[1][224] , \labels[1][223] , \labels[1][222] , 
	\labels[1][221] , \labels[1][220] , \labels[1][219] , 
	\labels[1][218] , \labels[1][217] , \labels[1][216] , 
	\labels[1][215] , \labels[1][214] , \labels[1][213] , 
	\labels[1][212] , \labels[1][211] , \labels[1][210] , 
	\labels[1][209] , \labels[1][208] , \labels[1][207] , 
	\labels[1][206] , \labels[1][205] , \labels[1][204] , 
	\labels[1][203] , \labels[1][202] , \labels[1][201] , 
	\labels[1][200] , \labels[1][199] , \labels[1][198] , 
	\labels[1][197] , \labels[1][196] , \labels[1][195] , 
	\labels[1][194] , \labels[1][193] , \labels[1][192] , 
	\labels[1][191] , \labels[1][190] , \labels[1][189] , 
	\labels[1][188] , \labels[1][187] , \labels[1][186] , 
	\labels[1][185] , \labels[1][184] , \labels[1][183] , 
	\labels[1][182] , \labels[1][181] , \labels[1][180] , 
	\labels[1][179] , \labels[1][178] , \labels[1][177] , 
	\labels[1][176] , \labels[1][175] , \labels[1][174] , 
	\labels[1][173] , \labels[1][172] , \labels[1][171] , 
	\labels[1][170] , \labels[1][169] , \labels[1][168] , 
	\labels[1][167] , \labels[1][166] , \labels[1][165] , 
	\labels[1][164] , \labels[1][163] , \labels[1][162] , 
	\labels[1][161] , \labels[1][160] , \labels[1][159] , 
	\labels[1][158] , \labels[1][157] , \labels[1][156] , 
	\labels[1][155] , \labels[1][154] , \labels[1][153] , 
	\labels[1][152] , \labels[1][151] , \labels[1][150] , 
	\labels[1][149] , \labels[1][148] , \labels[1][147] , 
	\labels[1][146] , \labels[1][145] , \labels[1][144] , 
	\labels[1][143] , \labels[1][142] , \labels[1][141] , 
	\labels[1][140] , \labels[1][139] , \labels[1][138] , 
	\labels[1][137] , \labels[1][136] , \labels[1][135] , 
	\labels[1][134] , \labels[1][133] , \labels[1][132] , 
	\labels[1][131] , \labels[1][130] , \labels[1][129] , 
	\labels[1][128] , \labels[1][127] , \labels[1][126] , 
	\labels[1][125] , \labels[1][124] , \labels[1][123] , 
	\labels[1][122] , \labels[1][121] , \labels[1][120] , 
	\labels[1][119] , \labels[1][118] , \labels[1][117] , 
	\labels[1][116] , \labels[1][115] , \labels[1][114] , 
	\labels[1][113] , \labels[1][112] , \labels[1][111] , 
	\labels[1][110] , \labels[1][109] , \labels[1][108] , 
	\labels[1][107] , \labels[1][106] , \labels[1][105] , 
	\labels[1][104] , \labels[1][103] , \labels[1][102] , 
	\labels[1][101] , \labels[1][100] , \labels[1][99] , \labels[1][98] , 
	\labels[1][97] , \labels[1][96] , \labels[1][95] , \labels[1][94] , 
	\labels[1][93] , \labels[1][92] , \labels[1][91] , \labels[1][90] , 
	\labels[1][89] , \labels[1][88] , \labels[1][87] , \labels[1][86] , 
	\labels[1][85] , \labels[1][84] , \labels[1][83] , \labels[1][82] , 
	\labels[1][81] , \labels[1][80] , \labels[1][79] , \labels[1][78] , 
	\labels[1][77] , \labels[1][76] , \labels[1][75] , \labels[1][74] , 
	\labels[1][73] , \labels[1][72] , \labels[1][71] , \labels[1][70] , 
	\labels[1][69] , \labels[1][68] , \labels[1][67] , \labels[1][66] , 
	\labels[1][65] , \labels[1][64] , \labels[1][63] , \labels[1][62] , 
	\labels[1][61] , \labels[1][60] , \labels[1][59] , \labels[1][58] , 
	\labels[1][57] , \labels[1][56] , \labels[1][55] , \labels[1][54] , 
	\labels[1][53] , \labels[1][52] , \labels[1][51] , \labels[1][50] , 
	\labels[1][49] , \labels[1][48] , \labels[1][47] , \labels[1][46] , 
	\labels[1][45] , \labels[1][44] , \labels[1][43] , \labels[1][42] , 
	\labels[1][41] , \labels[1][40] , \labels[1][39] , \labels[1][38] , 
	\labels[1][37] , \labels[1][36] , \labels[1][35] , \labels[1][34] , 
	\labels[1][33] , \labels[1][32] , \labels[1][31] , \labels[1][30] , 
	\labels[1][29] , \labels[1][28] , \labels[1][27] , \labels[1][26] , 
	\labels[1][25] , \labels[1][24] , \labels[1][23] , \labels[1][22] , 
	\labels[1][21] , \labels[1][20] , \labels[1][19] , \labels[1][18] , 
	\labels[1][17] , \labels[1][16] , \labels[1][15] , \labels[1][14] , 
	\labels[1][13] , \labels[1][12] , \labels[1][11] , \labels[1][10] , 
	\labels[1][9] , \labels[1][8] , \labels[1][7] , \labels[1][6] , 
	\labels[1][5] , \labels[1][4] , \labels[1][3] , \labels[1][2] , 
	\labels[1][1] , \labels[1][0] , \labels[0][271] , \labels[0][270] , 
	\labels[0][269] , \labels[0][268] , \labels[0][267] , 
	\labels[0][266] , \labels[0][265] , \labels[0][264] , 
	\labels[0][263] , \labels[0][262] , \labels[0][261] , 
	\labels[0][260] , \labels[0][259] , \labels[0][258] , 
	\labels[0][257] , \labels[0][256] , \labels[0][255] , 
	\labels[0][254] , \labels[0][253] , \labels[0][252] , 
	\labels[0][251] , \labels[0][250] , \labels[0][249] , 
	\labels[0][248] , \labels[0][247] , \labels[0][246] , 
	\labels[0][245] , \labels[0][244] , \labels[0][243] , 
	\labels[0][242] , \labels[0][241] , \labels[0][240] , 
	\labels[0][239] , \labels[0][238] , \labels[0][237] , 
	\labels[0][236] , \labels[0][235] , \labels[0][234] , 
	\labels[0][233] , \labels[0][232] , \labels[0][231] , 
	\labels[0][230] , \labels[0][229] , \labels[0][228] , 
	\labels[0][227] , \labels[0][226] , \labels[0][225] , 
	\labels[0][224] , \labels[0][223] , \labels[0][222] , 
	\labels[0][221] , \labels[0][220] , \labels[0][219] , 
	\labels[0][218] , \labels[0][217] , \labels[0][216] , 
	\labels[0][215] , \labels[0][214] , \labels[0][213] , 
	\labels[0][212] , \labels[0][211] , \labels[0][210] , 
	\labels[0][209] , \labels[0][208] , \labels[0][207] , 
	\labels[0][206] , \labels[0][205] , \labels[0][204] , 
	\labels[0][203] , \labels[0][202] , \labels[0][201] , 
	\labels[0][200] , \labels[0][199] , \labels[0][198] , 
	\labels[0][197] , \labels[0][196] , \labels[0][195] , 
	\labels[0][194] , \labels[0][193] , \labels[0][192] , 
	\labels[0][191] , \labels[0][190] , \labels[0][189] , 
	\labels[0][188] , \labels[0][187] , \labels[0][186] , 
	\labels[0][185] , \labels[0][184] , \labels[0][183] , 
	\labels[0][182] , \labels[0][181] , \labels[0][180] , 
	\labels[0][179] , \labels[0][178] , \labels[0][177] , 
	\labels[0][176] , \labels[0][175] , \labels[0][174] , 
	\labels[0][173] , \labels[0][172] , \labels[0][171] , 
	\labels[0][170] , \labels[0][169] , \labels[0][168] , 
	\labels[0][167] , \labels[0][166] , \labels[0][165] , 
	\labels[0][164] , \labels[0][163] , \labels[0][162] , 
	\labels[0][161] , \labels[0][160] , \labels[0][159] , 
	\labels[0][158] , \labels[0][157] , \labels[0][156] , 
	\labels[0][155] , \labels[0][154] , \labels[0][153] , 
	\labels[0][152] , \labels[0][151] , \labels[0][150] , 
	\labels[0][149] , \labels[0][148] , \labels[0][147] , 
	\labels[0][146] , \labels[0][145] , \labels[0][144] , 
	\labels[0][143] , \labels[0][142] , \labels[0][141] , 
	\labels[0][140] , \labels[0][139] , \labels[0][138] , 
	\labels[0][137] , \labels[0][136] , \labels[0][135] , 
	\labels[0][134] , \labels[0][133] , \labels[0][132] , 
	\labels[0][131] , \labels[0][130] , \labels[0][129] , 
	\labels[0][128] , \labels[0][127] , \labels[0][126] , 
	\labels[0][125] , \labels[0][124] , \labels[0][123] , 
	\labels[0][122] , \labels[0][121] , \labels[0][120] , 
	\labels[0][119] , \labels[0][118] , \labels[0][117] , 
	\labels[0][116] , \labels[0][115] , \labels[0][114] , 
	\labels[0][113] , \labels[0][112] , \labels[0][111] , 
	\labels[0][110] , \labels[0][109] , \labels[0][108] , 
	\labels[0][107] , \labels[0][106] , \labels[0][105] , 
	\labels[0][104] , \labels[0][103] , \labels[0][102] , 
	\labels[0][101] , \labels[0][100] , \labels[0][99] , \labels[0][98] , 
	\labels[0][97] , \labels[0][96] , \labels[0][95] , \labels[0][94] , 
	\labels[0][93] , \labels[0][92] , \labels[0][91] , \labels[0][90] , 
	\labels[0][89] , \labels[0][88] , \labels[0][87] , \labels[0][86] , 
	\labels[0][85] , \labels[0][84] , \labels[0][83] , \labels[0][82] , 
	\labels[0][81] , \labels[0][80] , \labels[0][79] , \labels[0][78] , 
	\labels[0][77] , \labels[0][76] , \labels[0][75] , \labels[0][74] , 
	\labels[0][73] , \labels[0][72] , \labels[0][71] , \labels[0][70] , 
	\labels[0][69] , \labels[0][68] , \labels[0][67] , \labels[0][66] , 
	\labels[0][65] , \labels[0][64] , \labels[0][63] , \labels[0][62] , 
	\labels[0][61] , \labels[0][60] , \labels[0][59] , \labels[0][58] , 
	\labels[0][57] , \labels[0][56] , \labels[0][55] , \labels[0][54] , 
	\labels[0][53] , \labels[0][52] , \labels[0][51] , \labels[0][50] , 
	\labels[0][49] , \labels[0][48] , \labels[0][47] , \labels[0][46] , 
	\labels[0][45] , \labels[0][44] , \labels[0][43] , \labels[0][42] , 
	\labels[0][41] , \labels[0][40] , \labels[0][39] , \labels[0][38] , 
	\labels[0][37] , \labels[0][36] , \labels[0][35] , \labels[0][34] , 
	\labels[0][33] , \labels[0][32] , \labels[0][31] , \labels[0][30] , 
	\labels[0][29] , \labels[0][28] , \labels[0][27] , \labels[0][26] , 
	\labels[0][25] , \labels[0][24] , \labels[0][23] , \labels[0][22] , 
	\labels[0][21] , \labels[0][20] , \labels[0][19] , \labels[0][18] , 
	\labels[0][17] , \labels[0][16] , \labels[0][15] , \labels[0][14] , 
	\labels[0][13] , \labels[0][12] , \labels[0][11] , \labels[0][10] , 
	\labels[0][9] , \labels[0][8] , \labels[0][7] , \labels[0][6] , 
	\labels[0][5] , \labels[0][4] , \labels[0][3] , \labels[0][2] , 
	\labels[0][1] , \labels[0][0] }), .cmdfifo_keyfilter_valid( 
	cmdfifo_keyfilter_valid), .cmdfifo_keyfilter_cmd( 
	cmdfifo_keyfilter_cmd[0]), .cmdfifo_kdf_valid( cmdfifo_kdf_valid), 
	.cmdfifo_kdf_cmd( cmdfifo_kdf_cmd[3:0]), .cmdfifo_kdfstream_valid( 
	cmdfifo_kdfstream_valid), .cmdfifo_kdfstream_cmd( 
	cmdfifo_kdfstream_cmd[262:0]), .gcm_kdf_valid( gcm_kdf_valid), 
	.gcm_kdf_eof( gcm_kdf_eof), .gcm_kdf_data( gcm_kdf_data[127:0]), 
	.keybuilder_kdf_stall( keybuilder_kdf_stall), .kdf_test_key_size( 
	kdf_test_key_size[31:0]), .kdf_test_mode_en( kdf_test_mode_en));
cr_kme_kop_keybuilder key_builder ( .tlv_sb_data_out_ack( 
	tlv_sb_data_out_ack), .keybuilder_kdf_stall( keybuilder_kdf_stall), 
	.gcm_status_data_out_ack( gcm_status_data_out_ack), .key_tlv_ob_wr( 
	key_tlv_ob_wr), .key_tlv_ob_tlv( 
	_zy_simnet_key_tlv_ob_tlv_6_w$[0:105]), .clk( clk), .rst_n( rst_n), 
	.tlv_sb_data_out( tlv_sb_data_out[63:0]), .tlv_sb_data_out_valid( 
	tlv_sb_data_out_valid), .kdf_keybuilder_data( 
	kdf_keybuilder_data[63:0]), .kdf_keybuilder_valid( 
	kdf_keybuilder_valid), .gcm_status_data_out_valid( 
	gcm_status_data_out_valid), .gcm_status_data_out( 
	gcm_status_data_out[0]), .key_tlv_ob_full( key_tlv_ob_full), 
	.key_tlv_ob_afull( key_tlv_ob_afull));
cr_kme_fifo_xcm50 gcm_cmd_fifo ( .fifo_in_stall( gcm_cmd_in_stall), 
	.fifo_out( cmdfifo_gcm_cmd[610:0]), .fifo_out_valid( 
	cmdfifo_gcm_valid), .fifo_overflow( _zy_simnet_dio_7), 
	.fifo_underflow( _zy_simnet_dio_8), .clk( clk), .rst_n( rst_n), 
	.fifo_in( _zy_simnet_gcm_cmd_in_9_w$[0:610]), .fifo_in_valid( 
	gcm_cmd_in_valid), .fifo_out_ack( gcm_cmdfifo_ack), 
	.fifo_in_stall_override( kop_fifo_override[0]));
cr_kme_fifo_xcm49 keyfilter_cmd_fifo ( .fifo_in_stall( 
	keyfilter_cmd_in_stall), .fifo_out( cmdfifo_keyfilter_cmd[0]), 
	.fifo_out_valid( cmdfifo_keyfilter_valid), .fifo_overflow( 
	_zy_simnet_dio_10), .fifo_underflow( _zy_simnet_dio_11), .clk( clk), 
	.rst_n( rst_n), .fifo_in( _zy_simnet_keyfilter_cmd_in_12_w$), 
	.fifo_in_valid( keyfilter_cmd_in_valid), .fifo_out_ack( 
	keyfilter_cmdfifo_ack), .fifo_in_stall_override( 
	kop_fifo_override[2]));
cr_kme_fifo_xcm48 kdf_cmd_fifo ( .fifo_in_stall( kdf_cmd_in_stall), 
	.fifo_out( cmdfifo_kdf_cmd[3:0]), .fifo_out_valid( 
	cmdfifo_kdf_valid), .fifo_overflow( _zy_simnet_dio_13), 
	.fifo_underflow( _zy_simnet_dio_14), .clk( clk), .rst_n( rst_n), 
	.fifo_in( _zy_simnet_kdf_cmd_in_15_w$[0:3]), .fifo_in_valid( 
	kdf_cmd_in_valid), .fifo_out_ack( kdf_cmdfifo_ack), 
	.fifo_in_stall_override( kop_fifo_override[4]));
cr_kme_fifo_xcm47 kdfstream_cmd_fifo ( .fifo_in_stall( 
	kdfstream_cmd_in_stall), .fifo_out( cmdfifo_kdfstream_cmd[262:0]), 
	.fifo_out_valid( cmdfifo_kdfstream_valid), .fifo_overflow( 
	_zy_simnet_dio_16), .fifo_underflow( _zy_simnet_dio_17), .clk( clk), 
	.rst_n( rst_n), .fifo_in( _zy_simnet_kdfstream_cmd_in_18_w$[0:262]), 
	.fifo_in_valid( kdfstream_cmd_in_valid), .fifo_out_ack( 
	kdfstream_cmdfifo_ack), .fifo_in_stall_override( 
	kop_fifo_override[3]));
cr_kme_fifo_xcm46 tlv_sb_data_fifo ( .fifo_in_stall( tlv_sb_data_in_stall), 
	.fifo_out( tlv_sb_data_out[63:0]), .fifo_out_valid( 
	tlv_sb_data_out_valid), .fifo_overflow( _zy_simnet_dio_19), 
	.fifo_underflow( _zy_simnet_dio_20), .clk( clk), .rst_n( rst_n), 
	.fifo_in( tlv_sb_data_in[63:0]), .fifo_in_valid( 
	tlv_sb_data_in_valid), .fifo_out_ack( tlv_sb_data_out_ack), 
	.fifo_in_stall_override( kop_fifo_override[5]));
cr_kme_fifo_xcm45 gcm_tag_data_fifo ( .fifo_in_stall( gcm_tag_data_in_stall), 
	.fifo_out( gcm_tag_data_out[95:0]), .fifo_out_valid( 
	gcm_tag_data_out_valid), .fifo_overflow( _zy_simnet_dio_21), 
	.fifo_underflow( _zy_simnet_dio_22), .clk( clk), .rst_n( rst_n), 
	.fifo_in( gcm_tag_data_in[95:0]), .fifo_in_valid( 
	gcm_tag_data_in_valid), .fifo_out_ack( gcm_tag_data_out_ack), 
	.fifo_in_stall_override( kop_fifo_override[1]));
cr_kme_fifo_xcm49 gcm_status_data_fifo ( .fifo_in_stall( 
	gcm_status_data_in_stall), .fifo_out( gcm_status_data_out[0]), 
	.fifo_out_valid( gcm_status_data_out_valid), .fifo_overflow( 
	_zy_simnet_dio_23), .fifo_underflow( _zy_simnet_dio_24), .clk( clk), 
	.rst_n( rst_n), .fifo_in( _zy_simnet_gcm_status_data_in_25_w$), 
	.fifo_in_valid( gcm_status_data_in_valid), .fifo_out_ack( 
	gcm_status_data_out_ack), .fifo_in_stall_override( 
	kop_fifo_override[6]));
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "\key_tlv_ob_tlv.ordern  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m2 "\key_tlv_ob_tlv.typen  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m3 "\key_tlv_ob_tlv.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m4 "\key_tlv_ob_tlv.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m5 "\key_tlv_ob_tlv.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m6 "\key_tlv_ob_tlv.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m7 "\labels%s.guid_size  1 0 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m8 "\labels%s.label_size  1 5 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m9 "\labels%s.label  1 255 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m10 "\labels%s.delimiter_valid  1 0 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m11 "\labels%s.delimiter  1 7 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m12 "labels (2,0) 1 271 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m13 "\kme_internal_out.sot  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m14 "\kme_internal_out.eoi  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m15 "\kme_internal_out.eot  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m16 "\kme_internal_out.id  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m17 "\kme_internal_out.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m18 "\kop_fifo_override.r.part0  (1,0) 1 6 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m19 "\gcm_cmd_in.key0  (1,0) 1 255 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m20 "\gcm_cmd_in.key1  (1,0) 1 255 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m21 "\gcm_cmd_in.iv  (1,0) 1 95 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m22 "\gcm_cmd_in.op  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m23 "\gcm_status_data_in.tag_mismatch  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m24 "\kdf_cmd_in.kdf_dek_iter  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m25 "\kdf_cmd_in.combo_mode  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m26 "\kdf_cmd_in.dek_key_op  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m27 "\kdf_cmd_in.dak_key_op  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m28 "\kdfstream_cmd_in.combo_mode  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m29 "\kdfstream_cmd_in.skip  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m30 "\kdfstream_cmd_in.guid  (1,0) 1 255 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m31 "\kdfstream_cmd_in.label_index  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m32 "\kdfstream_cmd_in.num_iter  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m33 "\keyfilter_cmd_in.combo_mode  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "33"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r1 "key_tlv_ob_tlv 10 \key_tlv_ob_tlv.insert  \key_tlv_ob_tlv.ordern  \key_tlv_ob_tlv.typen  \key_tlv_ob_tlv.sot  \key_tlv_ob_tlv.eot  \key_tlv_ob_tlv.tlast  \key_tlv_ob_tlv.tid  \key_tlv_ob_tlv.tstrb  \key_tlv_ob_tlv.tuser  \key_tlv_ob_tlv.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r2 "labels%s 5 \labels%s.guid_size  \labels%s.label_size  \labels%s.label  \labels%s.delimiter_valid  \labels%s.delimiter "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r3 "kme_internal_out 5 \kme_internal_out.sot  \kme_internal_out.eoi  \kme_internal_out.eot  \kme_internal_out.id  \kme_internal_out.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r1 "kop_fifo_override 2 \kop_fifo_override.r  { \kop_fifo_override.r.part0  } \kop_fifo_override.f  { \kop_fifo_override.f.gcm_status_data_fifo  \kop_fifo_override.f.tlv_sb_data_fifo  \kop_fifo_override.f.kdf_cmd_fifo  \kop_fifo_override.f.kdfstream_cmd_fifo  \kop_fifo_override.f.keyfilter_cmd_fifo  \kop_fifo_override.f.gcm_tag_data_fifo  \kop_fifo_override.f.gcm_cmd_fifo  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r4 "gcm_cmd_in 4 \gcm_cmd_in.key0  \gcm_cmd_in.key1  \gcm_cmd_in.iv  \gcm_cmd_in.op "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r5 "gcm_status_data_in 1 \gcm_status_data_in.tag_mismatch "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r6 "kdf_cmd_in 4 \kdf_cmd_in.kdf_dek_iter  \kdf_cmd_in.combo_mode  \kdf_cmd_in.dek_key_op  \kdf_cmd_in.dak_key_op "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r7 "kdfstream_cmd_in 5 \kdfstream_cmd_in.combo_mode  \kdfstream_cmd_in.skip  \kdfstream_cmd_in.guid  \kdfstream_cmd_in.label_index  \kdfstream_cmd_in.num_iter "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r8 "keyfilter_cmd_in 1 \keyfilter_cmd_in.combo_mode "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_NUM "8"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_NUM "1"
endmodule
