
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module kme_tb ;
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
wire _zy_simnet_kme_apb_psel_0_w$;
wire _zy_simnet_kme_apb_penable_1_w$;
wire [0:19] _zy_simnet_kme_apb_paddr_2_w$;
wire [0:31] _zy_simnet_kme_apb_pwdata_3_w$;
wire _zy_simnet_kme_apb_pwrite_4_w$;
wire _zy_simnet_clk_5_w$;
wire _zy_simnet_rst_n_6_w$;
wire [0:31] _zy_simnet_kme_apb_prdata_7_w$;
wire _zy_simnet_kme_apb_pready_8_w$;
wire _zy_simnet_kme_apb_pslverr_9_w$;
wire _zy_simnet_dio_10;
wire _zy_simnet_kme_ib_tready_11_w$;
wire _zy_simnet_kme_ob_tvalid_12_w$;
wire _zy_simnet_kme_ob_tlast_13_w$;
wire _zy_simnet_kme_ob_tid_14_w$;
wire [0:7] _zy_simnet_kme_ob_tstrb_15_w$;
wire [0:7] _zy_simnet_kme_ob_tuser_16_w$;
wire [0:63] _zy_simnet_kme_ob_tdata_17_w$;
wire [0:31] _zy_simnet_kme_apb_prdata_18_w$;
wire _zy_simnet_kme_apb_pready_19_w$;
wire _zy_simnet_kme_apb_pslverr_20_w$;
wire _zy_simnet_dio_21;
wire _zy_simnet_clk_22_w$;
wire _zy_simnet_rst_n_23_w$;
wire _zy_simnet_cio_24;
wire _zy_simnet_cio_25;
wire _zy_simnet_cio_26;
wire _zy_simnet_cio_27;
wire _zy_simnet_cio_28;
wire _zy_simnet_cio_29;
wire _zy_simnet_cio_30;
wire _zy_simnet_cio_31;
wire _zy_simnet_kme_ib_tvalid_32_w$;
wire _zy_simnet_kme_ib_tlast_33_w$;
wire _zy_simnet_kme_ib_tid_34_w$;
wire [0:7] _zy_simnet_kme_ib_tstrb_35_w$;
wire [0:7] _zy_simnet_kme_ib_tuser_36_w$;
wire [0:63] _zy_simnet_kme_ib_tdata_37_w$;
wire _zy_simnet_kme_ob_tready_38_w$;
wire [0:15] _zy_simnet_kme_apb_paddr_39_w$;
wire _zy_simnet_kme_apb_psel_40_w$;
wire _zy_simnet_kme_apb_penable_41_w$;
wire _zy_simnet_kme_apb_pwrite_42_w$;
wire [0:31] _zy_simnet_kme_apb_pwdata_43_w$;
wire _zyixc_port_0_0_s2h;
wire _zyixc_port_0_0_s2hW;
wire _zySfifoF0_call;
wire _zySfifoF0_fen;
wire [31:0] _zySfifoF0_iarg;
wire [511:0] _zyGfifo_SiData;
wire [21:0] _zyGfifo_StId;
wire [511:0] _zyGfifo_SoData;
wire _zyGfifo_SoDataEn;
wire [3:0] _zyGfifo_SoDataLen;
wire _zySfifoF1_call;
wire _zySfifoF1_fen;
wire [71:0] _zySfifoF1_iarg;
wire _zySfifoF2_call;
wire _zySfifoF2_fen;
wire [31:0] _zySfifoF2_iarg;
wire _zySfifoF3_call;
wire _zySfifoF3_fen;
wire [135:0] _zySfifoF3_iarg;
wire _zySfifoF4_call;
wire _zySfifoF4_fen;
wire [31:0] _zySfifoF4_iarg;
wire _zySfifoF5_call;
wire _zySfifoF5_fen;
wire [135:0] _zySfifoF5_iarg;
wire _zyL94_iscX1c0_f;
wire [31:0] _zyL94_iscX1c0_o1;
wire _zyL94_iscX1c0_o2;
wire _zyL61_iscX2c0_f;
wire _zyL61_iscX2c0_o2;
wire _zyictd_finish_mgr;
wire _zyGfifo_mod2_dflt_ci;
wire _zyGfifo_mod2_dflt_co;
wire [26:0] _zyGfifo_dflt_ci;
wire [26:0] _zyGfifo_dflt_co;
wire _zyGfifo_SGFtsReq;
wire [19:0] _zyGfifo_SGFcbid;
wire [11:0] _zyGfifo_SGFlen;
wire [511:0] _zyGfifo_SGFidata;
wire _zyGfifo_SGFfull;
wire _zyGfifo_SLBreq;
wire [3:0] _zyGfifo_SLBrd;
wire [3:0] _zyGfifo_SLBwr;
wire _zyGfifo_SLBfull;
wire _zyGfifo_SRtkin;
wire _zyM2L324_pbcMevClk4;
wire _zyM2L324_pbcReq4;
wire _zyM2L324_pbcBusy4;
wire _zyM2L324_pbcWait4;
wire _zyM2L253_pbcMevClk12;
wire _zyM2L253_pbcReq12;
wire _zyM2L253_pbcBusy12;
wire _zyM2L253_pbcWait12;
wire _zzM2_bcBehEvalClk;
wire _zzM2_bcBehHalt;
wire _zzmdxOne;
wire _zzM2L306_mdxP0_EnNxt;
wire _zzM2L306_mdxP0_On;
wire _zzM2L324_mdxP2_EnNxt;
wire _zzM2L324_mdxP2_On;
wire _zzM2L368_mdxP3_EnNxt;
wire _zzM2L368_mdxP3_On;
wire _zzM2L439_mdxP4_EnNxt;
wire _zzM2L439_mdxP4_On;
wire _zzM2L253_mdxP5_EnNxt;
wire _zzM2L253_mdxP5_On;
wire _zyictd_finish_mgr_x$tbc;
wire [279:0] testname;
wire [279:0] seed;
wire [31:0] initial_seed;
`_2_ wire [31:0] error_cntr;
wire clk;
wire rst_n;
wire kme_ib_tready;
wire [0:0] kme_ib_tid;
wire [63:0] kme_ib_tdata;
wire [7:0] kme_ib_tstrb;
wire [7:0] kme_ib_tuser;
wire kme_ib_tvalid;
wire kme_ib_tlast;
wire kme_ob_tready;
wire [0:0] kme_ob_tid;
wire [63:0] kme_ob_tdata;
wire [7:0] kme_ob_tstrb;
wire [7:0] kme_ob_tuser;
wire kme_ob_tvalid;
wire kme_ob_tlast;
wire [19:0] kme_apb_paddr;
wire kme_apb_psel;
wire kme_apb_penable;
wire kme_apb_pwrite;
wire [31:0] kme_apb_pwdata;
wire [31:0] kme_apb_prdata;
wire kme_apb_pready;
wire kme_apb_pslverr;
wire my_clk;
wire config_done;
`_2_ wire [7:0] tstrb_ib;
`_2_ wire [63:0] tdata_ib;
`_2_ wire [31:0] tuser_string_ib;
`_2_ wire [31:0] str_get_ib;
wire [24:0] user_string_ib;
`_2_ wire [31:0] retval_ib;
wire ready_ib;
wire saw_mega;
wire saw_guid_tlv;
wire have_guid_tlv;
`_2_ wire [31:0] mega_tlv_word_count;
`_2_ wire [7:0] tstrb_ob;
`_2_ wire [63:0] tdata_ob;
`_2_ wire [31:0] tuser_string_ob;
wire [24:0] user_string_ob;
`_2_ wire [31:0] str_get_ob;
`_2_ wire [31:0] retval_ob;
wire ready_ob;
wire [7:0] tuser;
wire tlast;
wire saw_cqe;
wire saw_stats;
wire ignore_compare_result;
wire [31:0] watchdog_timer;
wire [31:0] returned_data;
wire response;
`_2_ wire [7:0] operation;
`_2_ wire [31:0] address;
`_2_ wire [31:0] data;
`_2_ wire [31:0] retval;
wire config_ready;
wire [31:0] _zz_58_258_2;
wire [31:0] _zz_58_264_3;
`_2_ wire [4:0] _zygsfis_get_config_data_wptr;
`_2_ wire [4:0] _zygsfis_get_config_data_rptr;
`_2_ wire [4:0] _zygsfis_get_config_data_req;
`_2_ wire [4:0] _zygsfis_get_config_data_ack;
`_2_ wire _zygsfis_get_config_data_eos;
`_2_ wire [4:0] _zygsfis_get_config_data_space;
`_2_ wire [4:0] _zygsfis_ib_service_data_wptr;
`_2_ wire [4:0] _zygsfis_ib_service_data_rptr;
`_2_ wire [4:0] _zygsfis_ib_service_data_req;
`_2_ wire [4:0] _zygsfis_ib_service_data_ack;
`_2_ wire _zygsfis_ib_service_data_eos;
`_2_ wire [4:0] _zygsfis_ib_service_data_space;
`_2_ wire [4:0] _zygsfis_ob_service_data_wptr;
`_2_ wire [4:0] _zygsfis_ob_service_data_rptr;
`_2_ wire [4:0] _zygsfis_ob_service_data_req;
`_2_ wire [4:0] _zygsfis_ob_service_data_ack;
`_2_ wire _zygsfis_ob_service_data_eos;
`_2_ wire [4:0] _zygsfis_ob_service_data_space;
`_2_ wire _zyixc_port_0_0_req;
`_2_ wire _zyixc_port_0_0_ack;
`_2_ wire _zyixc_port_0_0_isf;
`_2_ wire _zyixc_port_0_0_osf;
`_2_ wire [21:0] _zySfifoF0_get_config_data_zyackf_tid;
`_2_ wire [21:0] _zySfifoF1_get_config_data_zyputf_tid;
`_2_ wire [21:0] _zySfifoF2_ib_service_data_zyackf_tid;
`_2_ wire [21:0] _zySfifoF3_ib_service_data_zyputf_tid;
`_2_ wire [21:0] _zySfifoF4_ob_service_data_zyackf_tid;
`_2_ wire [21:0] _zySfifoF5_ob_service_data_zyputf_tid;
wire _zyL94_iscX1c0_s;
wire _zyL94_iscX1c0_n;
wire [63:0] _zyL94_iscX1c0_i0;
wire _zyL61_iscX2c0_s;
wire _zyL61_iscX2c0_n;
wire [63:0] _zyL61_iscX2c0_i0;
wire [31:0] _zyL61_iscX2c0_i1;
wire [24:0] _zyL372_tfiRv5;
wire [7:0] _zyL406_tfiRv6;
wire [24:0] _zyL443_tfiRv7;
wire [7:0] _zyL462_tfiRv8;
wire [279:0] _zyictd_sysfunc_36_L258_0;
wire [31:0] _zyictd_sysfunc_36_L258_1;
wire [31:0] _zyictd_sysfunc_11_L257_2;
wire [279:0] _zyictd_sysfunc_36_L264_3;
wire [31:0] _zyictd_sysfunc_36_L264_4;
wire [31:0] _zyictd_sysfunc_11_L263_5;
`_2_ wire _zyictd_finish_L320_0;
`_2_ wire _zyictd_finish_L338_1;
`_2_ wire _zyictd_finish_L454_2;
`_2_ wire [31:0] _zyL326_tfiRv17;
`_2_ wire [31:0] _zyL370_tfiRv18;
`_2_ wire [31:0] _zyL441_tfiRv19;
`_2_ wire [0:0] _zyGfifo_mod2_simData;
`_2_ wire _zyGfifo__gfdL435_34_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL435_34_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL513_33_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL513_33_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL316_32_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL316_32_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL318_31_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL318_31_P0_m2_cbid;
`_2_ wire _zyGfifo_get_config_data_2_zyprefetch_m2_gfOff;
`_2_ wire [19:0] _zyGfifo_get_config_data_2_zyprefetch_m2_cbid;
`_2_ wire _zyGfifo__gfdL327_30_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL327_30_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL330_29_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL330_29_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL334_28_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL334_28_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL336_27_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL336_27_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL341_26_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL341_26_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL351_25_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL351_25_P0_m2_cbid;
`_2_ wire _zyGfifo_ib_service_data_2_zyprefetch_m2_gfOff;
`_2_ wire [19:0] _zyGfifo_ib_service_data_2_zyprefetch_m2_cbid;
`_2_ wire _zyGfifo__gfdL519_24_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL519_24_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL522_23_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL522_23_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL373_22_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL373_22_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL375_21_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL375_21_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL381_20_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL381_20_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL390_19_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL390_19_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL530_18_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL530_18_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL412_17_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL412_17_P0_m2_cbid;
`_2_ wire _zyGfifo_ob_service_data_2_zyprefetch_m2_gfOff;
`_2_ wire [19:0] _zyGfifo_ob_service_data_2_zyprefetch_m2_cbid;
`_2_ wire _zyGfifo__gfdL519_16_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL519_16_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL522_15_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL522_15_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL444_14_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL444_14_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL446_13_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL446_13_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL460_12_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL460_12_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL530_11_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL530_11_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL480_10_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL480_10_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL482_9_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL482_9_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL487_8_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL487_8_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL491_7_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL491_7_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL496_6_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL496_6_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL265_5_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL265_5_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL268_4_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL268_4_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL271_3_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL271_3_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL276_2_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL276_2_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL289_1_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL289_1_P0_m2_cbid;
`_2_ wire _zyGfifo__gfdL365_0_P0_m2_gfOff;
`_2_ wire [19:0] _zyGfifo__gfdL365_0_P0_m2_cbid;
`_2_ wire _zyGfifoF0_L435_req_0;
`_2_ wire _zyGfifoF1_L513_req_0;
`_2_ wire _zyGfifoF0_L312_s2_req_0;
`_2_ wire [279:0] _zyGfifoF0_L312_s2_data_0;
`_2_ wire [19:0] _zyGfifoF0_L312_s2_cbid_0;
`_2_ wire _zyGfifoF0_L324_s3_req_1;
`_2_ wire [95:0] _zyGfifoF0_L324_s3_data_1;
`_2_ wire [19:0] _zyGfifoF0_L324_s3_cbid_1;
`_2_ wire [11:0] _zyGfifoF0_L324_s3_len_1;
`_2_ wire _zyGfifoF1_L324_s2_req_2;
`_2_ wire [31:0] _zyGfifoF1_L324_s2_data_2;
`_2_ wire [19:0] _zyGfifoF1_L324_s2_cbid_2;
`_2_ wire _zyGfifoF2_L324_s2_req_3;
`_2_ wire [71:0] _zyGfifoF2_L324_s2_data_3;
`_2_ wire [19:0] _zyGfifoF2_L324_s2_cbid_3;
`_2_ wire [11:0] _zyGfifoF2_L324_s2_len_3;
`_2_ wire _zyGfifoF11_L207_req_0;
`_2_ wire [31:0] _zyGfifoF11_L207_data_0;
`_2_ wire _zyGfifoF0_L368_s2_req_4;
`_2_ wire [19:0] _zyGfifoF0_L368_s2_cbid_4;
`_2_ wire _zyGfifoF14_L373_req_0;
`_2_ wire [31:0] _zyGfifoF14_L373_data_0;
`_2_ wire _zyGfifoF15_L375_req_0;
`_2_ wire [135:0] _zyGfifoF15_L375_data_0;
`_2_ wire _zyGfifoF16_L381_req_0;
`_2_ wire _zyGfifoF17_L390_req_0;
`_2_ wire [63:0] _zyGfifoF17_L390_data_0;
`_2_ wire _zyGfifoF18_L530_req_0;
`_2_ wire [31:0] _zyGfifoF18_L530_data_0;
`_2_ wire _zyGfifoF19_L412_req_0;
`_2_ wire [7:0] _zyGfifoF19_L412_data_0;
`_2_ wire _zyGfifoF20_L209_req_0;
`_2_ wire [31:0] _zyGfifoF20_L209_data_0;
`_2_ wire _zyGfifoF0_L439_s2_req_5;
`_2_ wire [19:0] _zyGfifoF0_L439_s2_cbid_5;
`_2_ wire _zyGfifoF23_L444_req_0;
`_2_ wire [31:0] _zyGfifoF23_L444_data_0;
`_2_ wire _zyGfifoF24_L446_req_0;
`_2_ wire [135:0] _zyGfifoF24_L446_data_0;
`_2_ wire _zyGfifoF25_L460_req_0;
`_2_ wire [63:0] _zyGfifoF25_L460_data_0;
`_2_ wire _zyGfifoF26_L530_req_0;
`_2_ wire [31:0] _zyGfifoF26_L530_data_0;
`_2_ wire _zyGfifoF27_L480_req_0;
`_2_ wire [7:0] _zyGfifoF27_L480_data_0;
`_2_ wire _zyGfifoF28_L482_req_0;
`_2_ wire [127:0] _zyGfifoF28_L482_data_0;
`_2_ wire _zyGfifoF29_L487_req_0;
`_2_ wire [15:0] _zyGfifoF29_L487_data_0;
`_2_ wire _zyGfifoF30_L491_req_0;
`_2_ wire [15:0] _zyGfifoF30_L491_data_0;
`_2_ wire _zyGfifoF31_L496_req_0;
`_2_ wire [15:0] _zyGfifoF31_L496_data_0;
`_2_ wire _zyGfifoF0_L253_s4_req_6;
`_2_ wire [559:0] _zyGfifoF0_L253_s4_data_6;
`_2_ wire [19:0] _zyGfifoF0_L253_s4_cbid_6;
`_2_ wire [11:0] _zyGfifoF0_L253_s4_len_6;
`_2_ wire _zyGfifoF1_L253_s2_req_7;
`_2_ wire [19:0] _zyGfifoF1_L253_s2_cbid_7;
`_2_ wire [7:0] _zyoperation_L206_tfiV0_M2_pbcG0;
`_2_ wire [31:0] _zyaddress_L206_tfiV1_M2_pbcG1;
`_2_ wire [31:0] _zydata_L206_tfiV2_M2_pbcG2;
`_2_ wire [31:0] _zyxr_L206_tfiV3_M2_pbcG3;
wire [31:0] _zyM2L273_pbcT0;
wire [31:0] _zyM2L286_pbcT1;
wire [31:0] _zyM2L292_pbcT2;
wire [31:0] _zyM2L299_pbcT3;
wire _zyM2L324_pbcCapEn0;
wire _zyM2L333_pbcCapEn1;
wire _zyM2L349_pbcCapEn2;
wire _zyM2L355_pbcCapEn3;
wire _zyM2L253_pbcCapEn5;
wire _zyM2L274_pbcCapEn6;
wire _zyM2L287_pbcCapEn7;
wire _zyM2L293_pbcCapEn8;
wire _zyM2L295_pbcCapEn9;
wire _zyM2L364_pbcCapEn10;
wire _zyM2L300_pbcCapEn11;
wire [2:0] _zyM2L324_pbcFsm0_s;
wire _zyM2L324_pbcEn13;
wire [2:0] _zyM2L253_pbcFsm2_s;
wire _zyM2L253_pbcEn14;
wire [0:0] _zyL306_meState0;
wire [0:0] _zyL312_meState2;
wire [0:0] _zyL368_meState4;
wire [1:0] _zyL439_meState8;
wire [31:0] _zzM2_bcBehEval;
wire _zzM2L36_kme_ib_tvalid_mdxTmp0;
wire _zzM2L37_kme_ib_tlast_mdxTmp1;
wire _zzM2L306_mdxP0_En;
wire _zzM2L306_mdxP0_kme_ib_tvalid_wr0;
wire _zzM2L306_mdxP0_kme_ib_tvalid_Dwen0;
wire _zzM2L306_mdxP0_kme_ib_tvalid_DwenOn0;
wire _zzM2L306_mdxP0_kme_ib_tlast_wr1;
wire _zzM2L306_mdxP0_kme_ib_tlast_Dwen1;
wire _zzM2L306_mdxP0_kme_ib_tlast_DwenOn1;
`_2_ wire [31:0] _zzM2L19_error_cntr_mdxTmp2;
wire _zzM2L324_mdxP2_En;
`_2_ wire [31:0] _zzM2L324_mdxP2_error_cntr_wr0;
wire _zzM2L324_mdxP2_error_cntr_Dwen0;
wire _zzM2L324_mdxP2_error_cntr_DwenOn0;
wire [63:0] _zzM2L33_kme_ib_tdata_mdxTmp3;
wire [7:0] _zzM2L34_kme_ib_tstrb_mdxTmp4;
wire [7:0] _zzM2L35_kme_ib_tuser_mdxTmp5;
wire _zzM2L368_mdxP3_En;
wire _zzM2L368_mdxP3_kme_ib_tvalid_wr0;
wire _zzM2L368_mdxP3_kme_ib_tvalid_Dwen0;
wire _zzM2L368_mdxP3_kme_ib_tvalid_DwenOn0;
wire _zzM2L368_mdxP3_kme_ib_tlast_wr1;
wire _zzM2L368_mdxP3_kme_ib_tlast_Dwen1;
wire _zzM2L368_mdxP3_kme_ib_tlast_DwenOn1;
wire [63:0] _zzM2L368_mdxP3_kme_ib_tdata_wr2;
wire _zzM2L368_mdxP3_kme_ib_tdata_Dwen2;
wire _zzM2L368_mdxP3_kme_ib_tdata_DwenOn2;
wire [7:0] _zzM2L368_mdxP3_kme_ib_tstrb_wr3;
wire _zzM2L368_mdxP3_kme_ib_tstrb_Dwen3;
wire _zzM2L368_mdxP3_kme_ib_tstrb_DwenOn3;
wire [7:0] _zzM2L368_mdxP3_kme_ib_tuser_wr4;
wire _zzM2L368_mdxP3_kme_ib_tuser_Dwen4;
wire _zzM2L368_mdxP3_kme_ib_tuser_DwenOn4;
wire _zzM2L439_mdxP4_En;
`_2_ wire [31:0] _zzM2L439_mdxP4_error_cntr_wr0;
wire _zzM2L439_mdxP4_error_cntr_Dwen0;
wire _zzM2L439_mdxP4_error_cntr_DwenOn0;
wire _zzM2L253_mdxP5_En;
`_2_ wire [31:0] _zzM2L253_mdxP5_error_cntr_wr0;
wire _zzM2L253_mdxP5_error_cntr_Dwen0;
wire _zzM2L253_mdxP5_error_cntr_DwenOn0;
wire _zzM2L253_mdxP5_kme_ib_tvalid_wr1;
wire _zzM2L253_mdxP5_kme_ib_tvalid_Dwen1;
wire _zzM2L253_mdxP5_kme_ib_tvalid_DwenOn1;
wire _zzM2L253_mdxP5_kme_ib_tlast_wr2;
wire _zzM2L253_mdxP5_kme_ib_tlast_Dwen2;
wire _zzM2L253_mdxP5_kme_ib_tlast_DwenOn2;
wire [63:0] _zzM2L253_mdxP5_kme_ib_tdata_wr3;
wire _zzM2L253_mdxP5_kme_ib_tdata_Dwen3;
wire _zzM2L253_mdxP5_kme_ib_tdata_DwenOn3;
wire [7:0] _zzM2L253_mdxP5_kme_ib_tstrb_wr4;
wire _zzM2L253_mdxP5_kme_ib_tstrb_Dwen4;
wire _zzM2L253_mdxP5_kme_ib_tstrb_DwenOn4;
wire [7:0] _zzM2L253_mdxP5_kme_ib_tuser_wr5;
wire _zzM2L253_mdxP5_kme_ib_tuser_Dwen5;
wire _zzM2L253_mdxP5_kme_ib_tuser_DwenOn5;
`_2_ wire [31:0] _zzerror_cntr_M2L19_mdxSvLt6;
wire _zzkme_ib_tvalid_M2L36_mdxSvLt7;
wire _zzkme_ib_tlast_M2L37_mdxSvLt8;
wire [63:0] _zzkme_ib_tdata_M2L33_mdxSvLt9;
wire [7:0] _zzkme_ib_tstrb_M2L34_mdxSvLt10;
wire [7:0] _zzkme_ib_tuser_M2L35_mdxSvLt11;
wire [7:0] \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytstrb_L207_tfiV7 ;
wire [31:0] \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 ;
wire [31:0] \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 ;
wire [63:0] \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 ;
wire [7:0] \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytstrb_L209_tfiV13 ;
wire [31:0] \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 ;
wire [31:0] \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 ;
wire [63:0] \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 ;
supply0 n59;
supply0 n60;
supply0 n61;
supply0 n62;
supply0 n63;
supply0 n64;
supply0 n65;
supply0 n66;
supply0 n67;
supply0 n68;
supply0 n69;
supply0 n126;
supply0 n127;
supply0 n128;
supply0 n129;
supply0 n130;
supply0 n131;
supply0 n132;
supply0 n133;
supply0 n134;
supply0 n135;
supply0 n136;
supply0 n137;
supply0 n138;
supply0 n152;
supply0 n153;
supply0 n157;
supply0 n158;
supply0 n159;
supply1 n160;
supply0 n161;
supply0 n162;
supply0 n163;
supply0 n164;
supply0 n165;
supply0 n166;
supply0 n167;
supply0 n168;
supply0 n169;
supply0 n170;
supply0 n171;
supply0 n172;
supply0 n173;
supply0 n174;
supply0 n175;
supply0 n176;
supply0 n177;
supply0 n178;
supply0 n179;
supply0 n180;
supply0 n181;
supply0 n182;
supply0 n183;
supply0 n184;
supply0 n185;
supply0 n186;
supply0 n187;
supply0 n188;
supply0 n189;
supply0 n190;
supply0 n191;
supply0 n192;
supply0 n193;
supply0 n194;
supply1 n195;
supply0 n196;
supply0 n197;
supply1 n198;
supply0 n199;
supply0 n200;
supply0 n201;
supply0 n202;
supply0 n203;
supply0 n204;
supply0 n205;
supply0 n206;
supply0 n207;
supply0 n208;
supply0 n209;
supply1 n210;
supply0 n211;
supply0 n212;
supply0 n213;
supply0 n214;
supply0 n215;
supply0 n216;
supply0 n217;
supply0 n218;
supply0 n219;
supply0 n220;
supply0 n221;
supply1 n222;
supply0 n223;
supply0 n224;
supply0 n225;
supply0 n226;
supply0 n227;
supply0 n228;
supply0 n229;
supply0 n230;
supply0 n231;
supply0 n232;
supply0 n233;
supply0 n234;
supply0 n235;
supply0 n236;
supply0 n237;
supply0 n238;
supply0 n239;
supply0 n240;
supply0 n241;
supply0 n242;
supply0 n243;
supply0 n244;
supply0 n245;
supply0 n246;
supply1 n247;
supply0 n248;
supply0 n249;
supply0 n250;
supply0 n251;
supply0 n252;
supply0 n253;
supply0 n254;
supply0 n255;
supply0 n256;
supply1 n257;
supply0 n258;
supply1 n259;
supply0 n260;
supply0 n261;
supply0 n262;
supply0 n263;
supply0 n264;
supply0 n265;
supply0 n266;
supply0 n267;
supply0 n268;
supply0 n269;
supply0 n270;
supply0 n271;
supply0 n272;
supply0 n273;
supply0 n274;
supply0 n275;
supply0 n276;
supply0 n277;
supply0 n278;
supply0 n279;
supply0 n280;
supply0 n281;
supply0 n282;
supply1 n283;
supply0 n284;
supply0 n285;
supply0 n286;
supply0 n287;
supply0 n288;
supply0 n289;
supply0 n290;
supply0 n291;
supply0 n292;
supply0 n293;
supply0 n294;
supply0 n295;
supply1 n296;
supply0 n297;
supply0 n298;
supply0 n299;
supply0 n300;
supply0 n301;
supply0 n302;
supply0 n303;
supply0 n304;
supply0 n305;
supply0 n306;
supply0 n307;
supply1 n308;
supply0 n309;
supply0 n310;
supply0 n311;
supply0 n312;
supply0 n313;
supply0 n314;
supply0 n315;
supply0 n316;
supply0 n317;
supply0 n318;
supply0 n319;
supply1 n320;
supply0 n321;
supply0 n322;
supply0 n323;
supply0 n324;
supply0 n325;
supply0 n326;
supply0 n327;
supply0 n328;
supply0 n329;
supply0 n330;
supply0 n331;
supply0 n332;
supply0 n333;
supply0 n334;
supply0 n335;
supply0 n336;
supply0 n337;
supply0 n338;
supply0 n339;
supply0 n340;
supply0 n341;
supply0 n342;
supply0 n343;
supply0 n344;
supply1 n345;
supply0 n346;
supply0 n347;
supply0 n348;
supply0 n349;
supply0 n350;
supply0 n351;
supply0 n352;
supply0 n353;
supply0 n354;
supply1 n355;
supply0 n356;
supply1 n357;
supply0 n358;
supply0 n359;
supply0 n360;
supply0 n361;
supply0 n362;
supply0 n363;
supply0 n364;
supply0 n365;
supply0 n366;
supply0 n367;
supply1 n368;
supply0 n369;
supply0 n370;
supply0 n371;
supply0 n372;
supply0 n373;
supply0 n374;
supply0 n375;
supply0 n376;
supply0 n377;
supply0 n378;
supply0 n379;
supply0 n380;
supply1 n381;
supply0 n382;
supply0 n383;
supply0 n384;
supply0 n385;
supply0 n386;
supply0 n387;
supply0 n388;
supply0 n389;
supply0 n390;
supply0 n391;
supply0 n392;
supply1 n393;
supply0 n394;
supply0 n395;
supply0 n396;
supply0 n397;
supply0 n398;
supply0 n399;
supply0 n400;
supply0 n401;
supply0 n402;
supply1 n403;
supply0 n404;
supply0 n405;
supply0 n406;
supply0 n407;
supply0 n408;
supply0 n409;
supply0 n410;
supply0 n411;
supply0 n412;
supply0 n413;
supply0 n414;
supply0 n415;
supply0 n416;
supply1 n417;
supply0 n418;
supply0 n419;
supply0 n420;
supply0 n421;
supply0 n422;
supply0 n423;
supply0 n424;
supply0 n425;
supply0 n426;
supply0 n427;
supply0 n428;
supply1 n429;
supply0 n430;
supply0 n431;
supply0 n432;
supply0 n433;
supply0 n434;
supply0 n435;
supply0 n436;
supply0 n437;
supply0 n438;
supply0 n439;
supply0 n440;
supply1 n441;
supply0 n1750;
supply1 n5382;
Q_BUF U0 ( .A(n1750), .Z(_zy_simnet_cio_31));
Q_BUF U1 ( .A(n1750), .Z(_zy_simnet_cio_30));
Q_BUF U2 ( .A(n1750), .Z(_zy_simnet_cio_29));
Q_BUF U3 ( .A(n1750), .Z(_zy_simnet_cio_28));
Q_BUF U4 ( .A(n5382), .Z(_zy_simnet_cio_27));
Q_BUF U5 ( .A(n1750), .Z(_zy_simnet_cio_26));
Q_BUF U6 ( .A(n1750), .Z(_zy_simnet_cio_25));
Q_BUF U7 ( .A(n1750), .Z(_zy_simnet_cio_24));
Q_AN02 U8 ( .A0(n591), .A1(n1123), .Z(n5886));
Q_AN02 U9 ( .A0(n585), .A1(n1123), .Z(n5885));
Q_AN02 U10 ( .A0(n579), .A1(n1134), .Z(n5884));
Q_AN02 U11 ( .A0(n1268), .A1(n1629), .Z(n5883));
Q_AN02 U12 ( .A0(n1262), .A1(n1629), .Z(n5882));
Q_AN02 U13 ( .A0(n1256), .A1(n1641), .Z(n5881));
Q_AN02 U14 ( .A0(n2389), .A1(n3534), .Z(n5880));
Q_AN02 U15 ( .A0(n2400), .A1(n3534), .Z(n5879));
Q_AN02 U16 ( .A0(n2905), .A1(n3549), .Z(n5878));
Q_AN02 U17 ( .A0(n2383), .A1(n3559), .Z(n5877));
Q_AN02 U18 ( .A0(n5455), .A1(n5457), .Z(n5876));
Q_OA21 U19 ( .A0(n2376), .A1(n2371), .B0(n2377), .Z(n3564));
Q_MX03 U20 ( .S0(n3556), .S1(n3283), .A0(error_cntr[0]), .A1(n2656), .A2(n5875), .Z(n3096));
Q_XOR2 U21 ( .A0(n3556), .A1(n2906), .Z(n5875));
Q_OR03 U22 ( .A0(n3721), .A1(n3719), .A2(_zyM2L253_pbcFsm2_s[0]), .Z(n5325));
Q_FDP0 U23 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[63]), .Q(n5874), .QN( ));
Q_FDP0 U24 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[62]), .Q(n5873), .QN( ));
Q_FDP0 U25 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[61]), .Q(n5872), .QN( ));
Q_FDP0 U26 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[60]), .Q(n5871), .QN( ));
Q_FDP0 U27 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[59]), .Q(n5870), .QN( ));
Q_FDP0 U28 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[58]), .Q(n5869), .QN( ));
Q_FDP0 U29 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[57]), .Q(n5868), .QN( ));
Q_FDP0 U30 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[56]), .Q(n5867), .QN( ));
Q_FDP0 U31 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[55]), .Q(n5866), .QN( ));
Q_FDP0 U32 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[54]), .Q(n5865), .QN( ));
Q_FDP0 U33 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[53]), .Q(n5864), .QN( ));
Q_FDP0 U34 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[52]), .Q(n5863), .QN( ));
Q_FDP0 U35 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[51]), .Q(n5862), .QN( ));
Q_FDP0 U36 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[50]), .Q(n5861), .QN( ));
Q_FDP0 U37 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[49]), .Q(n5860), .QN( ));
Q_FDP0 U38 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[48]), .Q(n5859), .QN( ));
Q_FDP0 U39 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[47]), .Q(n5858), .QN( ));
Q_FDP0 U40 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[46]), .Q(n5857), .QN( ));
Q_FDP0 U41 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[45]), .Q(n5856), .QN( ));
Q_FDP0 U42 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[44]), .Q(n5855), .QN( ));
Q_FDP0 U43 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[43]), .Q(n5854), .QN( ));
Q_FDP0 U44 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[42]), .Q(n5853), .QN( ));
Q_FDP0 U45 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[41]), .Q(n5852), .QN( ));
Q_FDP0 U46 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[40]), .Q(n5851), .QN( ));
Q_FDP0 U47 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[39]), .Q(n5850), .QN( ));
Q_FDP0 U48 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[38]), .Q(n5849), .QN( ));
Q_FDP0 U49 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[37]), .Q(n5848), .QN( ));
Q_FDP0 U50 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[36]), .Q(n5847), .QN( ));
Q_FDP0 U51 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[35]), .Q(n5846), .QN( ));
Q_FDP0 U52 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[34]), .Q(n5845), .QN( ));
Q_FDP0 U53 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[33]), .Q(n5844), .QN( ));
Q_FDP0 U54 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[32]), .Q(n5843), .QN( ));
Q_FDP0 U55 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[31]), .Q(n5842), .QN( ));
Q_FDP0 U56 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[30]), .Q(n5841), .QN( ));
Q_FDP0 U57 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[29]), .Q(n5840), .QN( ));
Q_FDP0 U58 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[28]), .Q(n5839), .QN( ));
Q_FDP0 U59 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[27]), .Q(n5838), .QN( ));
Q_FDP0 U60 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[26]), .Q(n5837), .QN( ));
Q_FDP0 U61 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[25]), .Q(n5836), .QN( ));
Q_FDP0 U62 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[24]), .Q(n5835), .QN( ));
Q_FDP0 U63 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[23]), .Q(n5834), .QN( ));
Q_FDP0 U64 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[22]), .Q(n5833), .QN( ));
Q_FDP0 U65 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[21]), .Q(n5832), .QN( ));
Q_FDP0 U66 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[20]), .Q(n5831), .QN( ));
Q_FDP0 U67 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[19]), .Q(n5830), .QN( ));
Q_FDP0 U68 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[18]), .Q(n5829), .QN( ));
Q_FDP0 U69 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[17]), .Q(n5828), .QN( ));
Q_FDP0 U70 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[16]), .Q(n5827), .QN( ));
Q_FDP0 U71 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[15]), .Q(n5826), .QN( ));
Q_FDP0 U72 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[14]), .Q(n5825), .QN( ));
Q_FDP0 U73 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[13]), .Q(n5824), .QN( ));
Q_FDP0 U74 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[12]), .Q(n5823), .QN( ));
Q_FDP0 U75 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[11]), .Q(n5822), .QN( ));
Q_FDP0 U76 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[10]), .Q(n5821), .QN( ));
Q_FDP0 U77 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[9]), .Q(n5820), .QN( ));
Q_FDP0 U78 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[8]), .Q(n5819), .QN( ));
Q_FDP0 U79 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[7]), .Q(n5818), .QN( ));
Q_FDP0 U80 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[6]), .Q(n5817), .QN( ));
Q_FDP0 U81 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[5]), .Q(n5816), .QN( ));
Q_FDP0 U82 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[4]), .Q(n5815), .QN( ));
Q_FDP0 U83 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[3]), .Q(n5814), .QN( ));
Q_FDP0 U84 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[2]), .Q(n5813), .QN( ));
Q_FDP0 U85 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[1]), .Q(n5812), .QN( ));
Q_FDP0 U86 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[0]), .Q(n5811), .QN( ));
Q_FDP0 U87 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[95]), .Q(n5810), .QN( ));
Q_FDP0 U88 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[94]), .Q(n5809), .QN( ));
Q_FDP0 U89 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[93]), .Q(n5808), .QN( ));
Q_FDP0 U90 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[92]), .Q(n5807), .QN( ));
Q_FDP0 U91 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[91]), .Q(n5806), .QN( ));
Q_FDP0 U92 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[90]), .Q(n5805), .QN( ));
Q_FDP0 U93 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[89]), .Q(n5804), .QN( ));
Q_FDP0 U94 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[88]), .Q(n5803), .QN( ));
Q_FDP0 U95 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[87]), .Q(n5802), .QN( ));
Q_FDP0 U96 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[86]), .Q(n5801), .QN( ));
Q_FDP0 U97 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[85]), .Q(n5800), .QN( ));
Q_FDP0 U98 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[84]), .Q(n5799), .QN( ));
Q_FDP0 U99 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[83]), .Q(n5798), .QN( ));
Q_FDP0 U100 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[82]), .Q(n5797), .QN( ));
Q_FDP0 U101 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[81]), .Q(n5796), .QN( ));
Q_FDP0 U102 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[80]), .Q(n5795), .QN( ));
Q_FDP0 U103 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[79]), .Q(n5794), .QN( ));
Q_FDP0 U104 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[78]), .Q(n5793), .QN( ));
Q_FDP0 U105 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[77]), .Q(n5792), .QN( ));
Q_FDP0 U106 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[76]), .Q(n5791), .QN( ));
Q_FDP0 U107 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[75]), .Q(n5790), .QN( ));
Q_FDP0 U108 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[74]), .Q(n5789), .QN( ));
Q_FDP0 U109 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[73]), .Q(n5788), .QN( ));
Q_FDP0 U110 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[72]), .Q(n5787), .QN( ));
Q_FDP0 U111 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[71]), .Q(n5786), .QN( ));
Q_FDP0 U112 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[70]), .Q(n5785), .QN( ));
Q_FDP0 U113 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[69]), .Q(n5784), .QN( ));
Q_FDP0 U114 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[68]), .Q(n5783), .QN( ));
Q_FDP0 U115 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[67]), .Q(n5782), .QN( ));
Q_FDP0 U116 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[66]), .Q(n5781), .QN( ));
Q_FDP0 U117 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[65]), .Q(n5780), .QN( ));
Q_FDP0 U118 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[64]), .Q(n5779), .QN( ));
Q_FDP0 U119 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[103]), .Q(n5778), .QN( ));
Q_FDP0 U120 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[102]), .Q(n5777), .QN( ));
Q_FDP0 U121 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[101]), .Q(n5776), .QN( ));
Q_FDP0 U122 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[100]), .Q(n5775), .QN( ));
Q_FDP0 U123 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[99]), .Q(n5774), .QN( ));
Q_FDP0 U124 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[98]), .Q(n5773), .QN( ));
Q_FDP0 U125 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[97]), .Q(n5772), .QN( ));
Q_FDP0 U126 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[96]), .Q(n5771), .QN( ));
Q_FDP0 U127 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[135]), .Q(n5770), .QN( ));
Q_FDP0 U128 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[134]), .Q(n5769), .QN( ));
Q_FDP0 U129 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[133]), .Q(n5768), .QN( ));
Q_FDP0 U130 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[132]), .Q(n5767), .QN( ));
Q_FDP0 U131 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[131]), .Q(n5766), .QN( ));
Q_FDP0 U132 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[130]), .Q(n5765), .QN( ));
Q_FDP0 U133 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[129]), .Q(n5764), .QN( ));
Q_FDP0 U134 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[128]), .Q(n5763), .QN( ));
Q_FDP0 U135 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[127]), .Q(n5762), .QN( ));
Q_FDP0 U136 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[126]), .Q(n5761), .QN( ));
Q_FDP0 U137 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[125]), .Q(n5760), .QN( ));
Q_FDP0 U138 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[124]), .Q(n5759), .QN( ));
Q_FDP0 U139 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[123]), .Q(n5758), .QN( ));
Q_FDP0 U140 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[122]), .Q(n5757), .QN( ));
Q_FDP0 U141 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[121]), .Q(n5756), .QN( ));
Q_FDP0 U142 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[120]), .Q(n5755), .QN( ));
Q_FDP0 U143 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[119]), .Q(n5754), .QN( ));
Q_FDP0 U144 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[118]), .Q(n5753), .QN( ));
Q_FDP0 U145 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[117]), .Q(n5752), .QN( ));
Q_FDP0 U146 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[116]), .Q(n5751), .QN( ));
Q_FDP0 U147 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[115]), .Q(n5750), .QN( ));
Q_FDP0 U148 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[114]), .Q(n5749), .QN( ));
Q_FDP0 U149 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[113]), .Q(n5748), .QN( ));
Q_FDP0 U150 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[112]), .Q(n5747), .QN( ));
Q_FDP0 U151 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[111]), .Q(n5746), .QN( ));
Q_FDP0 U152 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[110]), .Q(n5745), .QN( ));
Q_FDP0 U153 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[109]), .Q(n5744), .QN( ));
Q_FDP0 U154 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[108]), .Q(n5743), .QN( ));
Q_FDP0 U155 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[107]), .Q(n5742), .QN( ));
Q_FDP0 U156 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[106]), .Q(n5741), .QN( ));
Q_FDP0 U157 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[105]), .Q(n5740), .QN( ));
Q_FDP0 U158 ( .CK(_zySfifoF5_call), .D(_zySfifoF5_iarg[104]), .Q(n5739), .QN( ));
Q_FDP0 U159 ( .CK(_zySfifoF5_call), .D(_zygsfis_ob_service_data_wptr[4]), .Q(n5738), .QN( ));
Q_FDP0 U160 ( .CK(_zySfifoF5_call), .D(_zygsfis_ob_service_data_wptr[3]), .Q(n5737), .QN( ));
Q_FDP0 U161 ( .CK(_zySfifoF5_call), .D(_zygsfis_ob_service_data_wptr[2]), .Q(n5736), .QN( ));
Q_FDP0 U162 ( .CK(_zySfifoF5_call), .D(_zygsfis_ob_service_data_wptr[1]), .Q(n5735), .QN( ));
Q_FDP0 U163 ( .CK(_zySfifoF5_call), .D(_zygsfis_ob_service_data_wptr[0]), .Q(n5734), .QN( ));
Q_XOR2 U164 ( .A0(n5730), .A1(n5732), .Z(n5733));
// pragma CVAINTPROP NET n5730 _2_state_ 1
// pragma CVAINTPROP INSTANCE U164 NOBREAKS 1
Q_FDP0B U165 ( .D(n5730), .QTFCLK( ), .Q(n5732));
Q_FDP0 U166 ( .CK(_zySfifoF5_call), .D(n5731), .Q(n5730), .QN(n5731));
Q_FDP0 U167 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[63]), .Q(n5729), .QN( ));
Q_FDP0 U168 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[62]), .Q(n5728), .QN( ));
Q_FDP0 U169 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[61]), .Q(n5727), .QN( ));
Q_FDP0 U170 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[60]), .Q(n5726), .QN( ));
Q_FDP0 U171 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[59]), .Q(n5725), .QN( ));
Q_FDP0 U172 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[58]), .Q(n5724), .QN( ));
Q_FDP0 U173 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[57]), .Q(n5723), .QN( ));
Q_FDP0 U174 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[56]), .Q(n5722), .QN( ));
Q_FDP0 U175 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[55]), .Q(n5721), .QN( ));
Q_FDP0 U176 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[54]), .Q(n5720), .QN( ));
Q_FDP0 U177 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[53]), .Q(n5719), .QN( ));
Q_FDP0 U178 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[52]), .Q(n5718), .QN( ));
Q_FDP0 U179 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[51]), .Q(n5717), .QN( ));
Q_FDP0 U180 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[50]), .Q(n5716), .QN( ));
Q_FDP0 U181 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[49]), .Q(n5715), .QN( ));
Q_FDP0 U182 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[48]), .Q(n5714), .QN( ));
Q_FDP0 U183 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[47]), .Q(n5713), .QN( ));
Q_FDP0 U184 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[46]), .Q(n5712), .QN( ));
Q_FDP0 U185 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[45]), .Q(n5711), .QN( ));
Q_FDP0 U186 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[44]), .Q(n5710), .QN( ));
Q_FDP0 U187 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[43]), .Q(n5709), .QN( ));
Q_FDP0 U188 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[42]), .Q(n5708), .QN( ));
Q_FDP0 U189 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[41]), .Q(n5707), .QN( ));
Q_FDP0 U190 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[40]), .Q(n5706), .QN( ));
Q_FDP0 U191 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[39]), .Q(n5705), .QN( ));
Q_FDP0 U192 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[38]), .Q(n5704), .QN( ));
Q_FDP0 U193 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[37]), .Q(n5703), .QN( ));
Q_FDP0 U194 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[36]), .Q(n5702), .QN( ));
Q_FDP0 U195 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[35]), .Q(n5701), .QN( ));
Q_FDP0 U196 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[34]), .Q(n5700), .QN( ));
Q_FDP0 U197 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[33]), .Q(n5699), .QN( ));
Q_FDP0 U198 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[32]), .Q(n5698), .QN( ));
Q_FDP0 U199 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[31]), .Q(n5697), .QN( ));
Q_FDP0 U200 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[30]), .Q(n5696), .QN( ));
Q_FDP0 U201 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[29]), .Q(n5695), .QN( ));
Q_FDP0 U202 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[28]), .Q(n5694), .QN( ));
Q_FDP0 U203 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[27]), .Q(n5693), .QN( ));
Q_FDP0 U204 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[26]), .Q(n5692), .QN( ));
Q_FDP0 U205 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[25]), .Q(n5691), .QN( ));
Q_FDP0 U206 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[24]), .Q(n5690), .QN( ));
Q_FDP0 U207 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[23]), .Q(n5689), .QN( ));
Q_FDP0 U208 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[22]), .Q(n5688), .QN( ));
Q_FDP0 U209 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[21]), .Q(n5687), .QN( ));
Q_FDP0 U210 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[20]), .Q(n5686), .QN( ));
Q_FDP0 U211 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[19]), .Q(n5685), .QN( ));
Q_FDP0 U212 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[18]), .Q(n5684), .QN( ));
Q_FDP0 U213 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[17]), .Q(n5683), .QN( ));
Q_FDP0 U214 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[16]), .Q(n5682), .QN( ));
Q_FDP0 U215 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[15]), .Q(n5681), .QN( ));
Q_FDP0 U216 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[14]), .Q(n5680), .QN( ));
Q_FDP0 U217 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[13]), .Q(n5679), .QN( ));
Q_FDP0 U218 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[12]), .Q(n5678), .QN( ));
Q_FDP0 U219 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[11]), .Q(n5677), .QN( ));
Q_FDP0 U220 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[10]), .Q(n5676), .QN( ));
Q_FDP0 U221 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[9]), .Q(n5675), .QN( ));
Q_FDP0 U222 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[8]), .Q(n5674), .QN( ));
Q_FDP0 U223 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[7]), .Q(n5673), .QN( ));
Q_FDP0 U224 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[6]), .Q(n5672), .QN( ));
Q_FDP0 U225 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[5]), .Q(n5671), .QN( ));
Q_FDP0 U226 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[4]), .Q(n5670), .QN( ));
Q_FDP0 U227 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[3]), .Q(n5669), .QN( ));
Q_FDP0 U228 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[2]), .Q(n5668), .QN( ));
Q_FDP0 U229 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[1]), .Q(n5667), .QN( ));
Q_FDP0 U230 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[0]), .Q(n5666), .QN( ));
Q_FDP0 U231 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[95]), .Q(n5665), .QN( ));
Q_FDP0 U232 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[94]), .Q(n5664), .QN( ));
Q_FDP0 U233 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[93]), .Q(n5663), .QN( ));
Q_FDP0 U234 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[92]), .Q(n5662), .QN( ));
Q_FDP0 U235 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[91]), .Q(n5661), .QN( ));
Q_FDP0 U236 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[90]), .Q(n5660), .QN( ));
Q_FDP0 U237 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[89]), .Q(n5659), .QN( ));
Q_FDP0 U238 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[88]), .Q(n5658), .QN( ));
Q_FDP0 U239 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[87]), .Q(n5657), .QN( ));
Q_FDP0 U240 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[86]), .Q(n5656), .QN( ));
Q_FDP0 U241 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[85]), .Q(n5655), .QN( ));
Q_FDP0 U242 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[84]), .Q(n5654), .QN( ));
Q_FDP0 U243 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[83]), .Q(n5653), .QN( ));
Q_FDP0 U244 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[82]), .Q(n5652), .QN( ));
Q_FDP0 U245 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[81]), .Q(n5651), .QN( ));
Q_FDP0 U246 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[80]), .Q(n5650), .QN( ));
Q_FDP0 U247 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[79]), .Q(n5649), .QN( ));
Q_FDP0 U248 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[78]), .Q(n5648), .QN( ));
Q_FDP0 U249 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[77]), .Q(n5647), .QN( ));
Q_FDP0 U250 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[76]), .Q(n5646), .QN( ));
Q_FDP0 U251 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[75]), .Q(n5645), .QN( ));
Q_FDP0 U252 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[74]), .Q(n5644), .QN( ));
Q_FDP0 U253 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[73]), .Q(n5643), .QN( ));
Q_FDP0 U254 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[72]), .Q(n5642), .QN( ));
Q_FDP0 U255 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[71]), .Q(n5641), .QN( ));
Q_FDP0 U256 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[70]), .Q(n5640), .QN( ));
Q_FDP0 U257 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[69]), .Q(n5639), .QN( ));
Q_FDP0 U258 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[68]), .Q(n5638), .QN( ));
Q_FDP0 U259 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[67]), .Q(n5637), .QN( ));
Q_FDP0 U260 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[66]), .Q(n5636), .QN( ));
Q_FDP0 U261 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[65]), .Q(n5635), .QN( ));
Q_FDP0 U262 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[64]), .Q(n5634), .QN( ));
Q_FDP0 U263 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[103]), .Q(n5633), .QN( ));
Q_FDP0 U264 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[102]), .Q(n5632), .QN( ));
Q_FDP0 U265 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[101]), .Q(n5631), .QN( ));
Q_FDP0 U266 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[100]), .Q(n5630), .QN( ));
Q_FDP0 U267 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[99]), .Q(n5629), .QN( ));
Q_FDP0 U268 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[98]), .Q(n5628), .QN( ));
Q_FDP0 U269 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[97]), .Q(n5627), .QN( ));
Q_FDP0 U270 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[96]), .Q(n5626), .QN( ));
Q_FDP0 U271 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[135]), .Q(n5625), .QN( ));
Q_FDP0 U272 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[134]), .Q(n5624), .QN( ));
Q_FDP0 U273 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[133]), .Q(n5623), .QN( ));
Q_FDP0 U274 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[132]), .Q(n5622), .QN( ));
Q_FDP0 U275 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[131]), .Q(n5621), .QN( ));
Q_FDP0 U276 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[130]), .Q(n5620), .QN( ));
Q_FDP0 U277 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[129]), .Q(n5619), .QN( ));
Q_FDP0 U278 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[128]), .Q(n5618), .QN( ));
Q_FDP0 U279 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[127]), .Q(n5617), .QN( ));
Q_FDP0 U280 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[126]), .Q(n5616), .QN( ));
Q_FDP0 U281 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[125]), .Q(n5615), .QN( ));
Q_FDP0 U282 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[124]), .Q(n5614), .QN( ));
Q_FDP0 U283 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[123]), .Q(n5613), .QN( ));
Q_FDP0 U284 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[122]), .Q(n5612), .QN( ));
Q_FDP0 U285 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[121]), .Q(n5611), .QN( ));
Q_FDP0 U286 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[120]), .Q(n5610), .QN( ));
Q_FDP0 U287 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[119]), .Q(n5609), .QN( ));
Q_FDP0 U288 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[118]), .Q(n5608), .QN( ));
Q_FDP0 U289 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[117]), .Q(n5607), .QN( ));
Q_FDP0 U290 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[116]), .Q(n5606), .QN( ));
Q_FDP0 U291 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[115]), .Q(n5605), .QN( ));
Q_FDP0 U292 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[114]), .Q(n5604), .QN( ));
Q_FDP0 U293 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[113]), .Q(n5603), .QN( ));
Q_FDP0 U294 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[112]), .Q(n5602), .QN( ));
Q_FDP0 U295 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[111]), .Q(n5601), .QN( ));
Q_FDP0 U296 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[110]), .Q(n5600), .QN( ));
Q_FDP0 U297 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[109]), .Q(n5599), .QN( ));
Q_FDP0 U298 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[108]), .Q(n5598), .QN( ));
Q_FDP0 U299 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[107]), .Q(n5597), .QN( ));
Q_FDP0 U300 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[106]), .Q(n5596), .QN( ));
Q_FDP0 U301 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[105]), .Q(n5595), .QN( ));
Q_FDP0 U302 ( .CK(_zySfifoF3_call), .D(_zySfifoF3_iarg[104]), .Q(n5594), .QN( ));
Q_FDP0 U303 ( .CK(_zySfifoF3_call), .D(_zygsfis_ib_service_data_wptr[4]), .Q(n5593), .QN( ));
Q_FDP0 U304 ( .CK(_zySfifoF3_call), .D(_zygsfis_ib_service_data_wptr[3]), .Q(n5592), .QN( ));
Q_FDP0 U305 ( .CK(_zySfifoF3_call), .D(_zygsfis_ib_service_data_wptr[2]), .Q(n5591), .QN( ));
Q_FDP0 U306 ( .CK(_zySfifoF3_call), .D(_zygsfis_ib_service_data_wptr[1]), .Q(n5590), .QN( ));
Q_FDP0 U307 ( .CK(_zySfifoF3_call), .D(_zygsfis_ib_service_data_wptr[0]), .Q(n5589), .QN( ));
Q_XOR2 U308 ( .A0(n5585), .A1(n5587), .Z(n5588));
// pragma CVAINTPROP NET n5585 _2_state_ 1
// pragma CVAINTPROP INSTANCE U308 NOBREAKS 1
Q_FDP0B U309 ( .D(n5585), .QTFCLK( ), .Q(n5587));
Q_FDP0 U310 ( .CK(_zySfifoF3_call), .D(n5586), .Q(n5585), .QN(n5586));
Q_FDP0 U311 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[7]), .Q(n5584), .QN( ));
Q_FDP0 U312 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[6]), .Q(n5583), .QN( ));
Q_FDP0 U313 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[5]), .Q(n5582), .QN( ));
Q_FDP0 U314 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[4]), .Q(n5581), .QN( ));
Q_FDP0 U315 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[3]), .Q(n5580), .QN( ));
Q_FDP0 U316 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[2]), .Q(n5579), .QN( ));
Q_FDP0 U317 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[1]), .Q(n5578), .QN( ));
Q_FDP0 U318 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[0]), .Q(n5577), .QN( ));
Q_FDP0 U319 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[39]), .Q(n5576), .QN( ));
Q_FDP0 U320 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[38]), .Q(n5575), .QN( ));
Q_FDP0 U321 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[37]), .Q(n5574), .QN( ));
Q_FDP0 U322 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[36]), .Q(n5573), .QN( ));
Q_FDP0 U323 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[35]), .Q(n5572), .QN( ));
Q_FDP0 U324 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[34]), .Q(n5571), .QN( ));
Q_FDP0 U325 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[33]), .Q(n5570), .QN( ));
Q_FDP0 U326 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[32]), .Q(n5569), .QN( ));
Q_FDP0 U327 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[31]), .Q(n5568), .QN( ));
Q_FDP0 U328 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[30]), .Q(n5567), .QN( ));
Q_FDP0 U329 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[29]), .Q(n5566), .QN( ));
Q_FDP0 U330 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[28]), .Q(n5565), .QN( ));
Q_FDP0 U331 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[27]), .Q(n5564), .QN( ));
Q_FDP0 U332 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[26]), .Q(n5563), .QN( ));
Q_FDP0 U333 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[25]), .Q(n5562), .QN( ));
Q_FDP0 U334 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[24]), .Q(n5561), .QN( ));
Q_FDP0 U335 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[23]), .Q(n5560), .QN( ));
Q_FDP0 U336 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[22]), .Q(n5559), .QN( ));
Q_FDP0 U337 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[21]), .Q(n5558), .QN( ));
Q_FDP0 U338 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[20]), .Q(n5557), .QN( ));
Q_FDP0 U339 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[19]), .Q(n5556), .QN( ));
Q_FDP0 U340 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[18]), .Q(n5555), .QN( ));
Q_FDP0 U341 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[17]), .Q(n5554), .QN( ));
Q_FDP0 U342 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[16]), .Q(n5553), .QN( ));
Q_FDP0 U343 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[15]), .Q(n5552), .QN( ));
Q_FDP0 U344 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[14]), .Q(n5551), .QN( ));
Q_FDP0 U345 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[13]), .Q(n5550), .QN( ));
Q_FDP0 U346 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[12]), .Q(n5549), .QN( ));
Q_FDP0 U347 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[11]), .Q(n5548), .QN( ));
Q_FDP0 U348 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[10]), .Q(n5547), .QN( ));
Q_FDP0 U349 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[9]), .Q(n5546), .QN( ));
Q_FDP0 U350 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[8]), .Q(n5545), .QN( ));
Q_FDP0 U351 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[71]), .Q(n5544), .QN( ));
Q_FDP0 U352 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[70]), .Q(n5543), .QN( ));
Q_FDP0 U353 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[69]), .Q(n5542), .QN( ));
Q_FDP0 U354 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[68]), .Q(n5541), .QN( ));
Q_FDP0 U355 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[67]), .Q(n5540), .QN( ));
Q_FDP0 U356 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[66]), .Q(n5539), .QN( ));
Q_FDP0 U357 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[65]), .Q(n5538), .QN( ));
Q_FDP0 U358 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[64]), .Q(n5537), .QN( ));
Q_FDP0 U359 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[63]), .Q(n5536), .QN( ));
Q_FDP0 U360 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[62]), .Q(n5535), .QN( ));
Q_FDP0 U361 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[61]), .Q(n5534), .QN( ));
Q_FDP0 U362 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[60]), .Q(n5533), .QN( ));
Q_FDP0 U363 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[59]), .Q(n5532), .QN( ));
Q_FDP0 U364 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[58]), .Q(n5531), .QN( ));
Q_FDP0 U365 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[57]), .Q(n5530), .QN( ));
Q_FDP0 U366 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[56]), .Q(n5529), .QN( ));
Q_FDP0 U367 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[55]), .Q(n5528), .QN( ));
Q_FDP0 U368 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[54]), .Q(n5527), .QN( ));
Q_FDP0 U369 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[53]), .Q(n5526), .QN( ));
Q_FDP0 U370 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[52]), .Q(n5525), .QN( ));
Q_FDP0 U371 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[51]), .Q(n5524), .QN( ));
Q_FDP0 U372 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[50]), .Q(n5523), .QN( ));
Q_FDP0 U373 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[49]), .Q(n5522), .QN( ));
Q_FDP0 U374 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[48]), .Q(n5521), .QN( ));
Q_FDP0 U375 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[47]), .Q(n5520), .QN( ));
Q_FDP0 U376 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[46]), .Q(n5519), .QN( ));
Q_FDP0 U377 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[45]), .Q(n5518), .QN( ));
Q_FDP0 U378 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[44]), .Q(n5517), .QN( ));
Q_FDP0 U379 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[43]), .Q(n5516), .QN( ));
Q_FDP0 U380 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[42]), .Q(n5515), .QN( ));
Q_FDP0 U381 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[41]), .Q(n5514), .QN( ));
Q_FDP0 U382 ( .CK(_zySfifoF1_call), .D(_zySfifoF1_iarg[40]), .Q(n5513), .QN( ));
Q_FDP0 U383 ( .CK(_zySfifoF1_call), .D(_zygsfis_get_config_data_wptr[4]), .Q(n5512), .QN( ));
Q_FDP0 U384 ( .CK(_zySfifoF1_call), .D(_zygsfis_get_config_data_wptr[3]), .Q(n5511), .QN( ));
Q_FDP0 U385 ( .CK(_zySfifoF1_call), .D(_zygsfis_get_config_data_wptr[2]), .Q(n5510), .QN( ));
Q_FDP0 U386 ( .CK(_zySfifoF1_call), .D(_zygsfis_get_config_data_wptr[1]), .Q(n5509), .QN( ));
Q_FDP0 U387 ( .CK(_zySfifoF1_call), .D(_zygsfis_get_config_data_wptr[0]), .Q(n5508), .QN( ));
Q_XOR2 U388 ( .A0(n5504), .A1(n5506), .Z(n5507));
// pragma CVAINTPROP NET n5504 _2_state_ 1
// pragma CVAINTPROP INSTANCE U388 NOBREAKS 1
Q_FDP0B U389 ( .D(n5504), .QTFCLK( ), .Q(n5506));
Q_FDP0 U390 ( .CK(_zySfifoF1_call), .D(n5505), .Q(n5504), .QN(n5505));
Q_INV U391 ( .A(_zzM2L253_mdxP5_kme_ib_tuser_DwenOn5), .Z(n5502));
Q_AN02 U392 ( .A0(_zzM2L368_mdxP3_kme_ib_tuser_DwenOn4), .A1(n5502), .Z(n5503));
Q_LDP0 \kme_ib_tuser_REG[0] ( .G(_zzmdxOne), .D(_zzM2L35_kme_ib_tuser_mdxTmp5[0]), .Q(kme_ib_tuser[0]), .QN( ));
Q_LDP0 \kme_ib_tuser_REG[1] ( .G(_zzmdxOne), .D(_zzM2L35_kme_ib_tuser_mdxTmp5[1]), .Q(kme_ib_tuser[1]), .QN( ));
Q_LDP0 \kme_ib_tuser_REG[2] ( .G(_zzmdxOne), .D(_zzM2L35_kme_ib_tuser_mdxTmp5[2]), .Q(kme_ib_tuser[2]), .QN( ));
Q_LDP0 \kme_ib_tuser_REG[3] ( .G(_zzmdxOne), .D(_zzM2L35_kme_ib_tuser_mdxTmp5[3]), .Q(kme_ib_tuser[3]), .QN( ));
Q_LDP0 \kme_ib_tuser_REG[4] ( .G(_zzmdxOne), .D(_zzM2L35_kme_ib_tuser_mdxTmp5[4]), .Q(kme_ib_tuser[4]), .QN( ));
Q_LDP0 \kme_ib_tuser_REG[5] ( .G(_zzmdxOne), .D(_zzM2L35_kme_ib_tuser_mdxTmp5[5]), .Q(kme_ib_tuser[5]), .QN( ));
Q_LDP0 \kme_ib_tuser_REG[6] ( .G(_zzmdxOne), .D(_zzM2L35_kme_ib_tuser_mdxTmp5[6]), .Q(kme_ib_tuser[6]), .QN( ));
Q_LDP0 \kme_ib_tuser_REG[7] ( .G(_zzmdxOne), .D(_zzM2L35_kme_ib_tuser_mdxTmp5[7]), .Q(kme_ib_tuser[7]), .QN( ));
Q_MX03 U401 ( .S0(n5503), .S1(_zzM2L253_mdxP5_kme_ib_tuser_DwenOn5), .A0(_zzkme_ib_tuser_M2L35_mdxSvLt11[7]), .A1(_zzM2L368_mdxP3_kme_ib_tuser_wr4[7]), .A2(_zzM2L253_mdxP5_kme_ib_tuser_wr5[7]), .Z(_zzM2L35_kme_ib_tuser_mdxTmp5[7]));
Q_MX03 U402 ( .S0(n5503), .S1(_zzM2L253_mdxP5_kme_ib_tuser_DwenOn5), .A0(_zzkme_ib_tuser_M2L35_mdxSvLt11[6]), .A1(_zzM2L368_mdxP3_kme_ib_tuser_wr4[6]), .A2(_zzM2L253_mdxP5_kme_ib_tuser_wr5[6]), .Z(_zzM2L35_kme_ib_tuser_mdxTmp5[6]));
Q_MX03 U403 ( .S0(n5503), .S1(_zzM2L253_mdxP5_kme_ib_tuser_DwenOn5), .A0(_zzkme_ib_tuser_M2L35_mdxSvLt11[5]), .A1(_zzM2L368_mdxP3_kme_ib_tuser_wr4[5]), .A2(_zzM2L253_mdxP5_kme_ib_tuser_wr5[5]), .Z(_zzM2L35_kme_ib_tuser_mdxTmp5[5]));
Q_MX03 U404 ( .S0(n5503), .S1(_zzM2L253_mdxP5_kme_ib_tuser_DwenOn5), .A0(_zzkme_ib_tuser_M2L35_mdxSvLt11[4]), .A1(_zzM2L368_mdxP3_kme_ib_tuser_wr4[4]), .A2(_zzM2L253_mdxP5_kme_ib_tuser_wr5[4]), .Z(_zzM2L35_kme_ib_tuser_mdxTmp5[4]));
Q_MX03 U405 ( .S0(n5503), .S1(_zzM2L253_mdxP5_kme_ib_tuser_DwenOn5), .A0(_zzkme_ib_tuser_M2L35_mdxSvLt11[3]), .A1(_zzM2L368_mdxP3_kme_ib_tuser_wr4[3]), .A2(_zzM2L253_mdxP5_kme_ib_tuser_wr5[3]), .Z(_zzM2L35_kme_ib_tuser_mdxTmp5[3]));
Q_MX03 U406 ( .S0(n5503), .S1(_zzM2L253_mdxP5_kme_ib_tuser_DwenOn5), .A0(_zzkme_ib_tuser_M2L35_mdxSvLt11[2]), .A1(_zzM2L368_mdxP3_kme_ib_tuser_wr4[2]), .A2(_zzM2L253_mdxP5_kme_ib_tuser_wr5[2]), .Z(_zzM2L35_kme_ib_tuser_mdxTmp5[2]));
Q_MX03 U407 ( .S0(n5503), .S1(_zzM2L253_mdxP5_kme_ib_tuser_DwenOn5), .A0(_zzkme_ib_tuser_M2L35_mdxSvLt11[1]), .A1(_zzM2L368_mdxP3_kme_ib_tuser_wr4[1]), .A2(_zzM2L253_mdxP5_kme_ib_tuser_wr5[1]), .Z(_zzM2L35_kme_ib_tuser_mdxTmp5[1]));
Q_MX03 U408 ( .S0(n5503), .S1(_zzM2L253_mdxP5_kme_ib_tuser_DwenOn5), .A0(_zzkme_ib_tuser_M2L35_mdxSvLt11[0]), .A1(_zzM2L368_mdxP3_kme_ib_tuser_wr4[0]), .A2(_zzM2L253_mdxP5_kme_ib_tuser_wr5[0]), .Z(_zzM2L35_kme_ib_tuser_mdxTmp5[0]));
Q_AN02 U409 ( .A0(_zzM2L253_mdxP5_On), .A1(_zzM2L253_mdxP5_kme_ib_tuser_Dwen5), .Z(_zzM2L253_mdxP5_kme_ib_tuser_DwenOn5));
Q_AN02 U410 ( .A0(_zzM2L368_mdxP3_On), .A1(_zzM2L368_mdxP3_kme_ib_tuser_Dwen4), .Z(_zzM2L368_mdxP3_kme_ib_tuser_DwenOn4));
Q_INV U411 ( .A(_zzM2L253_mdxP5_kme_ib_tstrb_DwenOn4), .Z(n5500));
Q_AN02 U412 ( .A0(_zzM2L368_mdxP3_kme_ib_tstrb_DwenOn3), .A1(n5500), .Z(n5501));
Q_LDP0 \kme_ib_tstrb_REG[0] ( .G(_zzmdxOne), .D(_zzM2L34_kme_ib_tstrb_mdxTmp4[0]), .Q(kme_ib_tstrb[0]), .QN( ));
Q_LDP0 \kme_ib_tstrb_REG[1] ( .G(_zzmdxOne), .D(_zzM2L34_kme_ib_tstrb_mdxTmp4[1]), .Q(kme_ib_tstrb[1]), .QN( ));
Q_LDP0 \kme_ib_tstrb_REG[2] ( .G(_zzmdxOne), .D(_zzM2L34_kme_ib_tstrb_mdxTmp4[2]), .Q(kme_ib_tstrb[2]), .QN( ));
Q_LDP0 \kme_ib_tstrb_REG[3] ( .G(_zzmdxOne), .D(_zzM2L34_kme_ib_tstrb_mdxTmp4[3]), .Q(kme_ib_tstrb[3]), .QN( ));
Q_LDP0 \kme_ib_tstrb_REG[4] ( .G(_zzmdxOne), .D(_zzM2L34_kme_ib_tstrb_mdxTmp4[4]), .Q(kme_ib_tstrb[4]), .QN( ));
Q_LDP0 \kme_ib_tstrb_REG[5] ( .G(_zzmdxOne), .D(_zzM2L34_kme_ib_tstrb_mdxTmp4[5]), .Q(kme_ib_tstrb[5]), .QN( ));
Q_LDP0 \kme_ib_tstrb_REG[6] ( .G(_zzmdxOne), .D(_zzM2L34_kme_ib_tstrb_mdxTmp4[6]), .Q(kme_ib_tstrb[6]), .QN( ));
Q_LDP0 \kme_ib_tstrb_REG[7] ( .G(_zzmdxOne), .D(_zzM2L34_kme_ib_tstrb_mdxTmp4[7]), .Q(kme_ib_tstrb[7]), .QN( ));
Q_MX03 U421 ( .S0(n5501), .S1(_zzM2L253_mdxP5_kme_ib_tstrb_DwenOn4), .A0(_zzkme_ib_tstrb_M2L34_mdxSvLt10[7]), .A1(_zzM2L368_mdxP3_kme_ib_tstrb_wr3[7]), .A2(_zzM2L253_mdxP5_kme_ib_tstrb_wr4[7]), .Z(_zzM2L34_kme_ib_tstrb_mdxTmp4[7]));
Q_MX03 U422 ( .S0(n5501), .S1(_zzM2L253_mdxP5_kme_ib_tstrb_DwenOn4), .A0(_zzkme_ib_tstrb_M2L34_mdxSvLt10[6]), .A1(_zzM2L368_mdxP3_kme_ib_tstrb_wr3[6]), .A2(_zzM2L253_mdxP5_kme_ib_tstrb_wr4[6]), .Z(_zzM2L34_kme_ib_tstrb_mdxTmp4[6]));
Q_MX03 U423 ( .S0(n5501), .S1(_zzM2L253_mdxP5_kme_ib_tstrb_DwenOn4), .A0(_zzkme_ib_tstrb_M2L34_mdxSvLt10[5]), .A1(_zzM2L368_mdxP3_kme_ib_tstrb_wr3[5]), .A2(_zzM2L253_mdxP5_kme_ib_tstrb_wr4[5]), .Z(_zzM2L34_kme_ib_tstrb_mdxTmp4[5]));
Q_MX03 U424 ( .S0(n5501), .S1(_zzM2L253_mdxP5_kme_ib_tstrb_DwenOn4), .A0(_zzkme_ib_tstrb_M2L34_mdxSvLt10[4]), .A1(_zzM2L368_mdxP3_kme_ib_tstrb_wr3[4]), .A2(_zzM2L253_mdxP5_kme_ib_tstrb_wr4[4]), .Z(_zzM2L34_kme_ib_tstrb_mdxTmp4[4]));
Q_MX03 U425 ( .S0(n5501), .S1(_zzM2L253_mdxP5_kme_ib_tstrb_DwenOn4), .A0(_zzkme_ib_tstrb_M2L34_mdxSvLt10[3]), .A1(_zzM2L368_mdxP3_kme_ib_tstrb_wr3[3]), .A2(_zzM2L253_mdxP5_kme_ib_tstrb_wr4[3]), .Z(_zzM2L34_kme_ib_tstrb_mdxTmp4[3]));
Q_MX03 U426 ( .S0(n5501), .S1(_zzM2L253_mdxP5_kme_ib_tstrb_DwenOn4), .A0(_zzkme_ib_tstrb_M2L34_mdxSvLt10[2]), .A1(_zzM2L368_mdxP3_kme_ib_tstrb_wr3[2]), .A2(_zzM2L253_mdxP5_kme_ib_tstrb_wr4[2]), .Z(_zzM2L34_kme_ib_tstrb_mdxTmp4[2]));
Q_MX03 U427 ( .S0(n5501), .S1(_zzM2L253_mdxP5_kme_ib_tstrb_DwenOn4), .A0(_zzkme_ib_tstrb_M2L34_mdxSvLt10[1]), .A1(_zzM2L368_mdxP3_kme_ib_tstrb_wr3[1]), .A2(_zzM2L253_mdxP5_kme_ib_tstrb_wr4[1]), .Z(_zzM2L34_kme_ib_tstrb_mdxTmp4[1]));
Q_MX03 U428 ( .S0(n5501), .S1(_zzM2L253_mdxP5_kme_ib_tstrb_DwenOn4), .A0(_zzkme_ib_tstrb_M2L34_mdxSvLt10[0]), .A1(_zzM2L368_mdxP3_kme_ib_tstrb_wr3[0]), .A2(_zzM2L253_mdxP5_kme_ib_tstrb_wr4[0]), .Z(_zzM2L34_kme_ib_tstrb_mdxTmp4[0]));
Q_AN02 U429 ( .A0(_zzM2L253_mdxP5_On), .A1(_zzM2L253_mdxP5_kme_ib_tstrb_Dwen4), .Z(_zzM2L253_mdxP5_kme_ib_tstrb_DwenOn4));
Q_AN02 U430 ( .A0(_zzM2L368_mdxP3_On), .A1(_zzM2L368_mdxP3_kme_ib_tstrb_Dwen3), .Z(_zzM2L368_mdxP3_kme_ib_tstrb_DwenOn3));
Q_INV U431 ( .A(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .Z(n5498));
Q_AN02 U432 ( .A0(_zzM2L368_mdxP3_kme_ib_tdata_DwenOn2), .A1(n5498), .Z(n5499));
Q_LDP0 \kme_ib_tdata_REG[0] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[0]), .Q(kme_ib_tdata[0]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[1] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[1]), .Q(kme_ib_tdata[1]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[2] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[2]), .Q(kme_ib_tdata[2]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[3] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[3]), .Q(kme_ib_tdata[3]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[4] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[4]), .Q(kme_ib_tdata[4]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[5] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[5]), .Q(kme_ib_tdata[5]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[6] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[6]), .Q(kme_ib_tdata[6]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[7] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[7]), .Q(kme_ib_tdata[7]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[8] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[8]), .Q(kme_ib_tdata[8]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[9] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[9]), .Q(kme_ib_tdata[9]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[10] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[10]), .Q(kme_ib_tdata[10]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[11] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[11]), .Q(kme_ib_tdata[11]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[12] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[12]), .Q(kme_ib_tdata[12]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[13] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[13]), .Q(kme_ib_tdata[13]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[14] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[14]), .Q(kme_ib_tdata[14]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[15] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[15]), .Q(kme_ib_tdata[15]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[16] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[16]), .Q(kme_ib_tdata[16]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[17] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[17]), .Q(kme_ib_tdata[17]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[18] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[18]), .Q(kme_ib_tdata[18]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[19] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[19]), .Q(kme_ib_tdata[19]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[20] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[20]), .Q(kme_ib_tdata[20]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[21] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[21]), .Q(kme_ib_tdata[21]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[22] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[22]), .Q(kme_ib_tdata[22]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[23] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[23]), .Q(kme_ib_tdata[23]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[24] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[24]), .Q(kme_ib_tdata[24]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[25] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[25]), .Q(kme_ib_tdata[25]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[26] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[26]), .Q(kme_ib_tdata[26]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[27] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[27]), .Q(kme_ib_tdata[27]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[28] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[28]), .Q(kme_ib_tdata[28]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[29] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[29]), .Q(kme_ib_tdata[29]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[30] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[30]), .Q(kme_ib_tdata[30]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[31] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[31]), .Q(kme_ib_tdata[31]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[32] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[32]), .Q(kme_ib_tdata[32]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[33] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[33]), .Q(kme_ib_tdata[33]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[34] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[34]), .Q(kme_ib_tdata[34]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[35] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[35]), .Q(kme_ib_tdata[35]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[36] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[36]), .Q(kme_ib_tdata[36]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[37] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[37]), .Q(kme_ib_tdata[37]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[38] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[38]), .Q(kme_ib_tdata[38]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[39] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[39]), .Q(kme_ib_tdata[39]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[40] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[40]), .Q(kme_ib_tdata[40]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[41] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[41]), .Q(kme_ib_tdata[41]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[42] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[42]), .Q(kme_ib_tdata[42]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[43] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[43]), .Q(kme_ib_tdata[43]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[44] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[44]), .Q(kme_ib_tdata[44]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[45] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[45]), .Q(kme_ib_tdata[45]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[46] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[46]), .Q(kme_ib_tdata[46]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[47] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[47]), .Q(kme_ib_tdata[47]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[48] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[48]), .Q(kme_ib_tdata[48]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[49] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[49]), .Q(kme_ib_tdata[49]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[50] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[50]), .Q(kme_ib_tdata[50]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[51] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[51]), .Q(kme_ib_tdata[51]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[52] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[52]), .Q(kme_ib_tdata[52]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[53] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[53]), .Q(kme_ib_tdata[53]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[54] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[54]), .Q(kme_ib_tdata[54]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[55] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[55]), .Q(kme_ib_tdata[55]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[56] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[56]), .Q(kme_ib_tdata[56]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[57] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[57]), .Q(kme_ib_tdata[57]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[58] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[58]), .Q(kme_ib_tdata[58]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[59] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[59]), .Q(kme_ib_tdata[59]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[60] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[60]), .Q(kme_ib_tdata[60]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[61] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[61]), .Q(kme_ib_tdata[61]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[62] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[62]), .Q(kme_ib_tdata[62]), .QN( ));
Q_LDP0 \kme_ib_tdata_REG[63] ( .G(_zzmdxOne), .D(_zzM2L33_kme_ib_tdata_mdxTmp3[63]), .Q(kme_ib_tdata[63]), .QN( ));
Q_MX03 U497 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[63]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[63]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[63]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[63]));
Q_MX03 U498 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[62]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[62]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[62]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[62]));
Q_MX03 U499 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[61]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[61]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[61]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[61]));
Q_MX03 U500 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[60]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[60]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[60]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[60]));
Q_MX03 U501 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[59]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[59]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[59]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[59]));
Q_MX03 U502 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[58]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[58]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[58]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[58]));
Q_MX03 U503 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[57]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[57]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[57]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[57]));
Q_MX03 U504 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[56]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[56]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[56]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[56]));
Q_MX03 U505 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[55]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[55]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[55]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[55]));
Q_MX03 U506 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[54]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[54]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[54]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[54]));
Q_MX03 U507 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[53]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[53]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[53]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[53]));
Q_MX03 U508 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[52]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[52]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[52]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[52]));
Q_MX03 U509 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[51]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[51]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[51]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[51]));
Q_MX03 U510 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[50]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[50]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[50]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[50]));
Q_MX03 U511 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[49]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[49]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[49]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[49]));
Q_MX03 U512 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[48]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[48]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[48]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[48]));
Q_MX03 U513 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[47]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[47]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[47]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[47]));
Q_MX03 U514 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[46]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[46]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[46]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[46]));
Q_MX03 U515 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[45]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[45]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[45]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[45]));
Q_MX03 U516 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[44]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[44]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[44]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[44]));
Q_MX03 U517 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[43]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[43]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[43]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[43]));
Q_MX03 U518 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[42]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[42]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[42]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[42]));
Q_MX03 U519 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[41]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[41]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[41]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[41]));
Q_MX03 U520 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[40]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[40]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[40]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[40]));
Q_MX03 U521 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[39]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[39]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[39]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[39]));
Q_MX03 U522 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[38]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[38]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[38]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[38]));
Q_MX03 U523 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[37]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[37]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[37]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[37]));
Q_MX03 U524 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[36]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[36]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[36]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[36]));
Q_MX03 U525 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[35]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[35]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[35]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[35]));
Q_MX03 U526 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[34]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[34]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[34]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[34]));
Q_MX03 U527 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[33]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[33]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[33]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[33]));
Q_MX03 U528 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[32]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[32]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[32]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[32]));
Q_MX03 U529 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[31]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[31]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[31]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[31]));
Q_MX03 U530 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[30]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[30]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[30]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[30]));
Q_MX03 U531 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[29]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[29]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[29]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[29]));
Q_MX03 U532 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[28]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[28]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[28]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[28]));
Q_MX03 U533 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[27]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[27]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[27]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[27]));
Q_MX03 U534 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[26]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[26]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[26]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[26]));
Q_MX03 U535 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[25]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[25]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[25]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[25]));
Q_MX03 U536 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[24]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[24]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[24]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[24]));
Q_MX03 U537 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[23]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[23]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[23]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[23]));
Q_MX03 U538 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[22]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[22]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[22]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[22]));
Q_MX03 U539 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[21]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[21]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[21]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[21]));
Q_MX03 U540 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[20]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[20]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[20]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[20]));
Q_MX03 U541 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[19]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[19]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[19]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[19]));
Q_MX03 U542 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[18]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[18]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[18]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[18]));
Q_MX03 U543 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[17]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[17]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[17]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[17]));
Q_MX03 U544 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[16]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[16]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[16]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[16]));
Q_MX03 U545 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[15]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[15]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[15]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[15]));
Q_MX03 U546 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[14]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[14]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[14]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[14]));
Q_MX03 U547 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[13]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[13]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[13]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[13]));
Q_MX03 U548 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[12]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[12]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[12]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[12]));
Q_MX03 U549 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[11]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[11]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[11]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[11]));
Q_MX03 U550 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[10]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[10]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[10]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[10]));
Q_MX03 U551 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[9]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[9]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[9]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[9]));
Q_MX03 U552 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[8]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[8]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[8]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[8]));
Q_MX03 U553 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[7]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[7]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[7]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[7]));
Q_MX03 U554 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[6]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[6]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[6]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[6]));
Q_MX03 U555 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[5]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[5]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[5]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[5]));
Q_MX03 U556 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[4]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[4]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[4]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[4]));
Q_MX03 U557 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[3]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[3]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[3]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[3]));
Q_MX03 U558 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[2]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[2]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[2]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[2]));
Q_MX03 U559 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[1]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[1]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[1]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[1]));
Q_MX03 U560 ( .S0(n5499), .S1(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3), .A0(_zzkme_ib_tdata_M2L33_mdxSvLt9[0]), .A1(_zzM2L368_mdxP3_kme_ib_tdata_wr2[0]), .A2(_zzM2L253_mdxP5_kme_ib_tdata_wr3[0]), .Z(_zzM2L33_kme_ib_tdata_mdxTmp3[0]));
Q_AN02 U561 ( .A0(_zzM2L253_mdxP5_On), .A1(_zzM2L253_mdxP5_kme_ib_tdata_Dwen3), .Z(_zzM2L253_mdxP5_kme_ib_tdata_DwenOn3));
Q_AN02 U562 ( .A0(_zzM2L368_mdxP3_On), .A1(_zzM2L368_mdxP3_kme_ib_tdata_Dwen2), .Z(_zzM2L368_mdxP3_kme_ib_tdata_DwenOn2));
Q_OR02 U563 ( .A0(_zzM2L253_mdxP5_kme_ib_tlast_DwenOn2), .A1(_zzM2L368_mdxP3_kme_ib_tlast_DwenOn1), .Z(n5497));
Q_INV U564 ( .A(_zzM2L306_mdxP0_kme_ib_tlast_DwenOn1), .Z(n5495));
Q_NR02 U565 ( .A0(_zzM2L368_mdxP3_kme_ib_tlast_DwenOn1), .A1(n5495), .Z(n5494));
Q_OR02 U566 ( .A0(_zzM2L253_mdxP5_kme_ib_tlast_DwenOn2), .A1(n5494), .Z(n5496));
Q_LDP0 kme_ib_tlast_REG  ( .G(_zzmdxOne), .D(_zzM2L37_kme_ib_tlast_mdxTmp1), .Q(kme_ib_tlast), .QN( ));
Q_MX04 U568 ( .S0(n5496), .S1(n5497), .A0(_zzkme_ib_tlast_M2L37_mdxSvLt8), .A1(_zzM2L306_mdxP0_kme_ib_tlast_wr1), .A2(_zzM2L368_mdxP3_kme_ib_tlast_wr1), .A3(_zzM2L253_mdxP5_kme_ib_tlast_wr2), .Z(_zzM2L37_kme_ib_tlast_mdxTmp1));
Q_AN02 U569 ( .A0(_zzM2L253_mdxP5_On), .A1(_zzM2L253_mdxP5_kme_ib_tlast_Dwen2), .Z(_zzM2L253_mdxP5_kme_ib_tlast_DwenOn2));
Q_AN02 U570 ( .A0(_zzM2L368_mdxP3_On), .A1(_zzM2L368_mdxP3_kme_ib_tlast_Dwen1), .Z(_zzM2L368_mdxP3_kme_ib_tlast_DwenOn1));
Q_AN02 U571 ( .A0(_zzM2L306_mdxP0_On), .A1(_zzM2L306_mdxP0_kme_ib_tlast_Dwen1), .Z(_zzM2L306_mdxP0_kme_ib_tlast_DwenOn1));
Q_OR02 U572 ( .A0(_zzM2L253_mdxP5_kme_ib_tvalid_DwenOn1), .A1(_zzM2L368_mdxP3_kme_ib_tvalid_DwenOn0), .Z(n5493));
Q_INV U573 ( .A(_zzM2L306_mdxP0_kme_ib_tvalid_DwenOn0), .Z(n5491));
Q_NR02 U574 ( .A0(_zzM2L368_mdxP3_kme_ib_tvalid_DwenOn0), .A1(n5491), .Z(n5490));
Q_OR02 U575 ( .A0(_zzM2L253_mdxP5_kme_ib_tvalid_DwenOn1), .A1(n5490), .Z(n5492));
Q_LDP0 kme_ib_tvalid_REG  ( .G(_zzmdxOne), .D(_zzM2L36_kme_ib_tvalid_mdxTmp0), .Q(kme_ib_tvalid), .QN( ));
Q_MX04 U577 ( .S0(n5492), .S1(n5493), .A0(_zzkme_ib_tvalid_M2L36_mdxSvLt7), .A1(_zzM2L306_mdxP0_kme_ib_tvalid_wr0), .A2(_zzM2L368_mdxP3_kme_ib_tvalid_wr0), .A3(_zzM2L253_mdxP5_kme_ib_tvalid_wr1), .Z(_zzM2L36_kme_ib_tvalid_mdxTmp0));
Q_AN02 U578 ( .A0(_zzM2L253_mdxP5_On), .A1(_zzM2L253_mdxP5_kme_ib_tvalid_Dwen1), .Z(_zzM2L253_mdxP5_kme_ib_tvalid_DwenOn1));
Q_AN02 U579 ( .A0(_zzM2L368_mdxP3_On), .A1(_zzM2L368_mdxP3_kme_ib_tvalid_Dwen0), .Z(_zzM2L368_mdxP3_kme_ib_tvalid_DwenOn0));
Q_AN02 U580 ( .A0(_zzM2L306_mdxP0_On), .A1(_zzM2L306_mdxP0_kme_ib_tvalid_Dwen0), .Z(_zzM2L306_mdxP0_kme_ib_tvalid_DwenOn0));
Q_LDP0 \error_cntr_REG[0] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[0]), .Q(error_cntr[0]), .QN(n553));
Q_LDP0 \error_cntr_REG[1] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[1]), .Q(error_cntr[1]), .QN( ));
Q_LDP0 \error_cntr_REG[2] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[2]), .Q(error_cntr[2]), .QN( ));
Q_LDP0 \error_cntr_REG[3] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[3]), .Q(error_cntr[3]), .QN( ));
Q_LDP0 \error_cntr_REG[4] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[4]), .Q(error_cntr[4]), .QN( ));
Q_LDP0 \error_cntr_REG[5] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[5]), .Q(error_cntr[5]), .QN( ));
Q_LDP0 \error_cntr_REG[6] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[6]), .Q(error_cntr[6]), .QN( ));
Q_LDP0 \error_cntr_REG[7] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[7]), .Q(error_cntr[7]), .QN( ));
Q_LDP0 \error_cntr_REG[8] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[8]), .Q(error_cntr[8]), .QN( ));
Q_LDP0 \error_cntr_REG[9] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[9]), .Q(error_cntr[9]), .QN( ));
Q_LDP0 \error_cntr_REG[10] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[10]), .Q(error_cntr[10]), .QN( ));
Q_LDP0 \error_cntr_REG[11] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[11]), .Q(error_cntr[11]), .QN( ));
Q_LDP0 \error_cntr_REG[12] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[12]), .Q(error_cntr[12]), .QN( ));
Q_LDP0 \error_cntr_REG[13] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[13]), .Q(error_cntr[13]), .QN( ));
Q_LDP0 \error_cntr_REG[14] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[14]), .Q(error_cntr[14]), .QN( ));
Q_LDP0 \error_cntr_REG[15] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[15]), .Q(error_cntr[15]), .QN( ));
Q_LDP0 \error_cntr_REG[16] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[16]), .Q(error_cntr[16]), .QN( ));
Q_LDP0 \error_cntr_REG[17] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[17]), .Q(error_cntr[17]), .QN( ));
Q_LDP0 \error_cntr_REG[18] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[18]), .Q(error_cntr[18]), .QN( ));
Q_LDP0 \error_cntr_REG[19] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[19]), .Q(error_cntr[19]), .QN( ));
Q_LDP0 \error_cntr_REG[20] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[20]), .Q(error_cntr[20]), .QN( ));
Q_LDP0 \error_cntr_REG[21] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[21]), .Q(error_cntr[21]), .QN( ));
Q_LDP0 \error_cntr_REG[22] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[22]), .Q(error_cntr[22]), .QN( ));
Q_LDP0 \error_cntr_REG[23] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[23]), .Q(error_cntr[23]), .QN( ));
Q_LDP0 \error_cntr_REG[24] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[24]), .Q(error_cntr[24]), .QN( ));
Q_LDP0 \error_cntr_REG[25] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[25]), .Q(error_cntr[25]), .QN( ));
Q_LDP0 \error_cntr_REG[26] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[26]), .Q(error_cntr[26]), .QN( ));
Q_LDP0 \error_cntr_REG[27] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[27]), .Q(error_cntr[27]), .QN( ));
Q_LDP0 \error_cntr_REG[28] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[28]), .Q(error_cntr[28]), .QN( ));
Q_LDP0 \error_cntr_REG[29] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[29]), .Q(error_cntr[29]), .QN( ));
Q_LDP0 \error_cntr_REG[30] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[30]), .Q(error_cntr[30]), .QN( ));
Q_LDP0 \error_cntr_REG[31] ( .G(_zzmdxOne), .D(_zzM2L19_error_cntr_mdxTmp2[31]), .Q(error_cntr[31]), .QN( ));
Q_MX03 U613 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5489), .A1(_zzM2L439_mdxP4_error_cntr_wr0[31]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[31]), .Z(_zzM2L19_error_cntr_mdxTmp2[31]));
Q_MX03 U614 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5488), .A1(_zzM2L439_mdxP4_error_cntr_wr0[30]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[30]), .Z(_zzM2L19_error_cntr_mdxTmp2[30]));
Q_MX03 U615 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5487), .A1(_zzM2L439_mdxP4_error_cntr_wr0[29]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[29]), .Z(_zzM2L19_error_cntr_mdxTmp2[29]));
Q_MX03 U616 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5486), .A1(_zzM2L439_mdxP4_error_cntr_wr0[28]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[28]), .Z(_zzM2L19_error_cntr_mdxTmp2[28]));
Q_MX03 U617 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5485), .A1(_zzM2L439_mdxP4_error_cntr_wr0[27]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[27]), .Z(_zzM2L19_error_cntr_mdxTmp2[27]));
Q_MX03 U618 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5484), .A1(_zzM2L439_mdxP4_error_cntr_wr0[26]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[26]), .Z(_zzM2L19_error_cntr_mdxTmp2[26]));
Q_MX03 U619 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5483), .A1(_zzM2L439_mdxP4_error_cntr_wr0[25]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[25]), .Z(_zzM2L19_error_cntr_mdxTmp2[25]));
Q_MX03 U620 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5482), .A1(_zzM2L439_mdxP4_error_cntr_wr0[24]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[24]), .Z(_zzM2L19_error_cntr_mdxTmp2[24]));
Q_MX03 U621 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5481), .A1(_zzM2L439_mdxP4_error_cntr_wr0[23]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[23]), .Z(_zzM2L19_error_cntr_mdxTmp2[23]));
Q_MX03 U622 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5480), .A1(_zzM2L439_mdxP4_error_cntr_wr0[22]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[22]), .Z(_zzM2L19_error_cntr_mdxTmp2[22]));
Q_MX03 U623 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5479), .A1(_zzM2L439_mdxP4_error_cntr_wr0[21]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[21]), .Z(_zzM2L19_error_cntr_mdxTmp2[21]));
Q_MX03 U624 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5478), .A1(_zzM2L439_mdxP4_error_cntr_wr0[20]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[20]), .Z(_zzM2L19_error_cntr_mdxTmp2[20]));
Q_MX03 U625 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5477), .A1(_zzM2L439_mdxP4_error_cntr_wr0[19]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[19]), .Z(_zzM2L19_error_cntr_mdxTmp2[19]));
Q_MX03 U626 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5476), .A1(_zzM2L439_mdxP4_error_cntr_wr0[18]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[18]), .Z(_zzM2L19_error_cntr_mdxTmp2[18]));
Q_MX03 U627 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5475), .A1(_zzM2L439_mdxP4_error_cntr_wr0[17]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[17]), .Z(_zzM2L19_error_cntr_mdxTmp2[17]));
Q_MX03 U628 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5474), .A1(_zzM2L439_mdxP4_error_cntr_wr0[16]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[16]), .Z(_zzM2L19_error_cntr_mdxTmp2[16]));
Q_MX03 U629 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5473), .A1(_zzM2L439_mdxP4_error_cntr_wr0[15]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[15]), .Z(_zzM2L19_error_cntr_mdxTmp2[15]));
Q_MX03 U630 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5472), .A1(_zzM2L439_mdxP4_error_cntr_wr0[14]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[14]), .Z(_zzM2L19_error_cntr_mdxTmp2[14]));
Q_MX03 U631 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5471), .A1(_zzM2L439_mdxP4_error_cntr_wr0[13]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[13]), .Z(_zzM2L19_error_cntr_mdxTmp2[13]));
Q_MX03 U632 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5470), .A1(_zzM2L439_mdxP4_error_cntr_wr0[12]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[12]), .Z(_zzM2L19_error_cntr_mdxTmp2[12]));
Q_MX03 U633 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5469), .A1(_zzM2L439_mdxP4_error_cntr_wr0[11]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[11]), .Z(_zzM2L19_error_cntr_mdxTmp2[11]));
Q_MX03 U634 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5468), .A1(_zzM2L439_mdxP4_error_cntr_wr0[10]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[10]), .Z(_zzM2L19_error_cntr_mdxTmp2[10]));
Q_MX03 U635 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5467), .A1(_zzM2L439_mdxP4_error_cntr_wr0[9]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[9]), .Z(_zzM2L19_error_cntr_mdxTmp2[9]));
Q_MX03 U636 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5466), .A1(_zzM2L439_mdxP4_error_cntr_wr0[8]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[8]), .Z(_zzM2L19_error_cntr_mdxTmp2[8]));
Q_MX03 U637 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5465), .A1(_zzM2L439_mdxP4_error_cntr_wr0[7]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[7]), .Z(_zzM2L19_error_cntr_mdxTmp2[7]));
Q_MX03 U638 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5464), .A1(_zzM2L439_mdxP4_error_cntr_wr0[6]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[6]), .Z(_zzM2L19_error_cntr_mdxTmp2[6]));
Q_MX03 U639 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5463), .A1(_zzM2L439_mdxP4_error_cntr_wr0[5]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[5]), .Z(_zzM2L19_error_cntr_mdxTmp2[5]));
Q_MX03 U640 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5462), .A1(_zzM2L439_mdxP4_error_cntr_wr0[4]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[4]), .Z(_zzM2L19_error_cntr_mdxTmp2[4]));
Q_MX03 U641 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5461), .A1(_zzM2L439_mdxP4_error_cntr_wr0[3]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[3]), .Z(_zzM2L19_error_cntr_mdxTmp2[3]));
Q_MX03 U642 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5460), .A1(_zzM2L439_mdxP4_error_cntr_wr0[2]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[2]), .Z(_zzM2L19_error_cntr_mdxTmp2[2]));
Q_MX03 U643 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5459), .A1(_zzM2L439_mdxP4_error_cntr_wr0[1]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[1]), .Z(_zzM2L19_error_cntr_mdxTmp2[1]));
Q_MX03 U644 ( .S0(_zzM2L439_mdxP4_error_cntr_DwenOn0), .S1(_zzM2L253_mdxP5_error_cntr_DwenOn0), .A0(n5458), .A1(_zzM2L439_mdxP4_error_cntr_wr0[0]), .A2(_zzM2L253_mdxP5_error_cntr_wr0[0]), .Z(_zzM2L19_error_cntr_mdxTmp2[0]));
Q_AN02 U645 ( .A0(_zzM2L253_mdxP5_On), .A1(_zzM2L253_mdxP5_error_cntr_Dwen0), .Z(_zzM2L253_mdxP5_error_cntr_DwenOn0));
Q_AN02 U646 ( .A0(_zzM2L439_mdxP4_On), .A1(_zzM2L439_mdxP4_error_cntr_Dwen0), .Z(_zzM2L439_mdxP4_error_cntr_DwenOn0));
Q_MX02 U647 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[31]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[31]), .Z(n5489));
Q_MX02 U648 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[30]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[30]), .Z(n5488));
Q_MX02 U649 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[29]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[29]), .Z(n5487));
Q_MX02 U650 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[28]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[28]), .Z(n5486));
Q_MX02 U651 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[27]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[27]), .Z(n5485));
Q_MX02 U652 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[26]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[26]), .Z(n5484));
Q_MX02 U653 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[25]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[25]), .Z(n5483));
Q_MX02 U654 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[24]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[24]), .Z(n5482));
Q_MX02 U655 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[23]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[23]), .Z(n5481));
Q_MX02 U656 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[22]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[22]), .Z(n5480));
Q_MX02 U657 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[21]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[21]), .Z(n5479));
Q_MX02 U658 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[20]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[20]), .Z(n5478));
Q_MX02 U659 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[19]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[19]), .Z(n5477));
Q_MX02 U660 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[18]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[18]), .Z(n5476));
Q_MX02 U661 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[17]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[17]), .Z(n5475));
Q_MX02 U662 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[16]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[16]), .Z(n5474));
Q_MX02 U663 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[15]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[15]), .Z(n5473));
Q_MX02 U664 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[14]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[14]), .Z(n5472));
Q_MX02 U665 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[13]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[13]), .Z(n5471));
Q_MX02 U666 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[12]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[12]), .Z(n5470));
Q_MX02 U667 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[11]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[11]), .Z(n5469));
Q_MX02 U668 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[10]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[10]), .Z(n5468));
Q_MX02 U669 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[9]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[9]), .Z(n5467));
Q_MX02 U670 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[8]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[8]), .Z(n5466));
Q_MX02 U671 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[7]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[7]), .Z(n5465));
Q_MX02 U672 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[6]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[6]), .Z(n5464));
Q_MX02 U673 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[5]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[5]), .Z(n5463));
Q_MX02 U674 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[4]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[4]), .Z(n5462));
Q_MX02 U675 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[3]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[3]), .Z(n5461));
Q_MX02 U676 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[2]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[2]), .Z(n5460));
Q_MX02 U677 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[1]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[1]), .Z(n5459));
Q_MX02 U678 ( .S(_zzM2L324_mdxP2_error_cntr_DwenOn0), .A0(_zzerror_cntr_M2L19_mdxSvLt6[0]), .A1(_zzM2L324_mdxP2_error_cntr_wr0[0]), .Z(n5458));
Q_AN02 U679 ( .A0(_zzM2L324_mdxP2_On), .A1(_zzM2L324_mdxP2_error_cntr_Dwen0), .Z(_zzM2L324_mdxP2_error_cntr_DwenOn0));
Q_AN02 U680 ( .A0(n5456), .A1(n5397), .Z(n5457));
Q_AD01HF U681 ( .A0(_zzM2_bcBehEval[29]), .B0(n5453), .S(n5454), .CO(n5455));
Q_AD01HF U682 ( .A0(_zzM2_bcBehEval[28]), .B0(n5451), .S(n5452), .CO(n5453));
Q_AD01HF U683 ( .A0(_zzM2_bcBehEval[27]), .B0(n5449), .S(n5450), .CO(n5451));
Q_AD01HF U684 ( .A0(_zzM2_bcBehEval[26]), .B0(n5447), .S(n5448), .CO(n5449));
Q_AD01HF U685 ( .A0(_zzM2_bcBehEval[25]), .B0(n5445), .S(n5446), .CO(n5447));
Q_AD01HF U686 ( .A0(_zzM2_bcBehEval[24]), .B0(n5443), .S(n5444), .CO(n5445));
Q_AD01HF U687 ( .A0(_zzM2_bcBehEval[23]), .B0(n5441), .S(n5442), .CO(n5443));
Q_AD01HF U688 ( .A0(_zzM2_bcBehEval[22]), .B0(n5439), .S(n5440), .CO(n5441));
Q_AD01HF U689 ( .A0(_zzM2_bcBehEval[21]), .B0(n5437), .S(n5438), .CO(n5439));
Q_AD01HF U690 ( .A0(_zzM2_bcBehEval[20]), .B0(n5435), .S(n5436), .CO(n5437));
Q_AD01HF U691 ( .A0(_zzM2_bcBehEval[19]), .B0(n5433), .S(n5434), .CO(n5435));
Q_AD01HF U692 ( .A0(_zzM2_bcBehEval[18]), .B0(n5431), .S(n5432), .CO(n5433));
Q_AD01HF U693 ( .A0(_zzM2_bcBehEval[17]), .B0(n5429), .S(n5430), .CO(n5431));
Q_AD01HF U694 ( .A0(_zzM2_bcBehEval[16]), .B0(n5427), .S(n5428), .CO(n5429));
Q_AD01HF U695 ( .A0(_zzM2_bcBehEval[15]), .B0(n5425), .S(n5426), .CO(n5427));
Q_AD01HF U696 ( .A0(_zzM2_bcBehEval[14]), .B0(n5423), .S(n5424), .CO(n5425));
Q_AD01HF U697 ( .A0(_zzM2_bcBehEval[13]), .B0(n5421), .S(n5422), .CO(n5423));
Q_AD01HF U698 ( .A0(_zzM2_bcBehEval[12]), .B0(n5419), .S(n5420), .CO(n5421));
Q_AD01HF U699 ( .A0(_zzM2_bcBehEval[11]), .B0(n5417), .S(n5418), .CO(n5419));
Q_AD01HF U700 ( .A0(_zzM2_bcBehEval[10]), .B0(n5415), .S(n5416), .CO(n5417));
Q_AD01HF U701 ( .A0(_zzM2_bcBehEval[9]), .B0(n5413), .S(n5414), .CO(n5415));
Q_AD01HF U702 ( .A0(_zzM2_bcBehEval[8]), .B0(n5411), .S(n5412), .CO(n5413));
Q_AD01HF U703 ( .A0(_zzM2_bcBehEval[7]), .B0(n5409), .S(n5410), .CO(n5411));
Q_AD01HF U704 ( .A0(_zzM2_bcBehEval[6]), .B0(n5407), .S(n5408), .CO(n5409));
Q_AD01HF U705 ( .A0(_zzM2_bcBehEval[5]), .B0(n5405), .S(n5406), .CO(n5407));
Q_AD01HF U706 ( .A0(_zzM2_bcBehEval[4]), .B0(n5403), .S(n5404), .CO(n5405));
Q_AD01HF U707 ( .A0(_zzM2_bcBehEval[3]), .B0(n5401), .S(n5402), .CO(n5403));
Q_AD01HF U708 ( .A0(_zzM2_bcBehEval[2]), .B0(n5399), .S(n5400), .CO(n5401));
Q_AD01HF U709 ( .A0(_zzM2_bcBehEval[1]), .B0(_zzM2_bcBehEval[0]), .S(n5398), .CO(n5399));
Q_OR02 U710 ( .A0(_zyM2L324_pbcWait4), .A1(_zyM2L253_pbcWait12), .Z(n5456));
Q_ND03 U711 ( .A0(n5394), .A1(n5395), .A2(n5396), .Z(n5397));
Q_AN03 U712 ( .A0(n5391), .A1(n5392), .A2(n5393), .Z(n5396));
Q_AN03 U713 ( .A0(n5388), .A1(n5389), .A2(n5390), .Z(n5395));
Q_AN03 U714 ( .A0(n5385), .A1(n5386), .A2(n5387), .Z(n5394));
Q_AN03 U715 ( .A0(_zzM2_bcBehEval[0]), .A1(n5383), .A2(n5384), .Z(n5393));
Q_AN03 U716 ( .A0(_zzM2_bcBehEval[3]), .A1(_zzM2_bcBehEval[2]), .A2(_zzM2_bcBehEval[1]), .Z(n5392));
Q_AN03 U717 ( .A0(_zzM2_bcBehEval[6]), .A1(_zzM2_bcBehEval[5]), .A2(_zzM2_bcBehEval[4]), .Z(n5391));
Q_AN03 U718 ( .A0(_zzM2_bcBehEval[9]), .A1(_zzM2_bcBehEval[8]), .A2(_zzM2_bcBehEval[7]), .Z(n5390));
Q_AN03 U719 ( .A0(_zzM2_bcBehEval[12]), .A1(_zzM2_bcBehEval[11]), .A2(_zzM2_bcBehEval[10]), .Z(n5389));
Q_AN03 U720 ( .A0(_zzM2_bcBehEval[15]), .A1(_zzM2_bcBehEval[14]), .A2(_zzM2_bcBehEval[13]), .Z(n5388));
Q_AN03 U721 ( .A0(_zzM2_bcBehEval[18]), .A1(_zzM2_bcBehEval[17]), .A2(_zzM2_bcBehEval[16]), .Z(n5387));
Q_AN03 U722 ( .A0(_zzM2_bcBehEval[21]), .A1(_zzM2_bcBehEval[20]), .A2(_zzM2_bcBehEval[19]), .Z(n5386));
Q_AN03 U723 ( .A0(_zzM2_bcBehEval[24]), .A1(_zzM2_bcBehEval[23]), .A2(_zzM2_bcBehEval[22]), .Z(n5385));
Q_AN03 U724 ( .A0(_zzM2_bcBehEval[27]), .A1(_zzM2_bcBehEval[26]), .A2(_zzM2_bcBehEval[25]), .Z(n5384));
Q_AN03 U725 ( .A0(_zzM2_bcBehEval[30]), .A1(_zzM2_bcBehEval[29]), .A2(_zzM2_bcBehEval[28]), .Z(n5383));
Q_AD01HF U726 ( .A0(_zygsfis_ob_service_data_wptr[1]), .B0(_zygsfis_ob_service_data_wptr[0]), .S(n5380), .CO(n5379));
Q_AD01HF U727 ( .A0(_zygsfis_ob_service_data_wptr[2]), .B0(n5379), .S(n5378), .CO(n5377));
Q_AD01HF U728 ( .A0(_zygsfis_ob_service_data_wptr[3]), .B0(n5377), .S(n5376), .CO(n5375));
Q_FDP0 \_zygsfis_ob_service_data_wptr_REG[3] ( .CK(_zySfifoF5_call), .D(n5376), .Q(_zygsfis_ob_service_data_wptr[3]), .QN( ));
Q_FDP0 \_zygsfis_ob_service_data_wptr_REG[2] ( .CK(_zySfifoF5_call), .D(n5378), .Q(_zygsfis_ob_service_data_wptr[2]), .QN( ));
Q_FDP0 \_zygsfis_ob_service_data_wptr_REG[1] ( .CK(_zySfifoF5_call), .D(n5380), .Q(_zygsfis_ob_service_data_wptr[1]), .QN( ));
Q_FDP0 \_zygsfis_ob_service_data_wptr_REG[0] ( .CK(_zySfifoF5_call), .D(n5381), .Q(_zygsfis_ob_service_data_wptr[0]), .QN(n5381));
Q_AD01HF U733 ( .A0(_zygsfis_ob_service_data_ack[1]), .B0(_zygsfis_ob_service_data_ack[0]), .S(n5373), .CO(n5372));
Q_AD01HF U734 ( .A0(_zygsfis_ob_service_data_ack[2]), .B0(n5372), .S(n5371), .CO(n5370));
Q_AD01HF U735 ( .A0(_zygsfis_ob_service_data_ack[3]), .B0(n5370), .S(n5369), .CO(n5368));
Q_FDP0 \_zygsfis_ob_service_data_ack_REG[3] ( .CK(_zySfifoF4_call), .D(n5369), .Q(_zygsfis_ob_service_data_ack[3]), .QN( ));
Q_FDP0 \_zygsfis_ob_service_data_ack_REG[2] ( .CK(_zySfifoF4_call), .D(n5371), .Q(_zygsfis_ob_service_data_ack[2]), .QN( ));
Q_FDP0 \_zygsfis_ob_service_data_ack_REG[1] ( .CK(_zySfifoF4_call), .D(n5373), .Q(_zygsfis_ob_service_data_ack[1]), .QN( ));
Q_FDP0 \_zygsfis_ob_service_data_ack_REG[0] ( .CK(_zySfifoF4_call), .D(n5374), .Q(_zygsfis_ob_service_data_ack[0]), .QN(n5374));
Q_FDP0 _zygsfis_ob_service_data_eos_REG  ( .CK(_zySfifoF4_call), .D(_zySfifoF4_iarg[0]), .Q(_zygsfis_ob_service_data_eos), .QN( ));
Q_AD01HF U741 ( .A0(_zygsfis_ib_service_data_wptr[1]), .B0(_zygsfis_ib_service_data_wptr[0]), .S(n5366), .CO(n5365));
Q_AD01HF U742 ( .A0(_zygsfis_ib_service_data_wptr[2]), .B0(n5365), .S(n5364), .CO(n5363));
Q_AD01HF U743 ( .A0(_zygsfis_ib_service_data_wptr[3]), .B0(n5363), .S(n5362), .CO(n5361));
Q_FDP0 \_zygsfis_ib_service_data_wptr_REG[3] ( .CK(_zySfifoF3_call), .D(n5362), .Q(_zygsfis_ib_service_data_wptr[3]), .QN( ));
Q_FDP0 \_zygsfis_ib_service_data_wptr_REG[2] ( .CK(_zySfifoF3_call), .D(n5364), .Q(_zygsfis_ib_service_data_wptr[2]), .QN( ));
Q_FDP0 \_zygsfis_ib_service_data_wptr_REG[1] ( .CK(_zySfifoF3_call), .D(n5366), .Q(_zygsfis_ib_service_data_wptr[1]), .QN( ));
Q_FDP0 \_zygsfis_ib_service_data_wptr_REG[0] ( .CK(_zySfifoF3_call), .D(n5367), .Q(_zygsfis_ib_service_data_wptr[0]), .QN(n5367));
Q_AD01HF U748 ( .A0(_zygsfis_ib_service_data_ack[1]), .B0(_zygsfis_ib_service_data_ack[0]), .S(n5359), .CO(n5358));
Q_AD01HF U749 ( .A0(_zygsfis_ib_service_data_ack[2]), .B0(n5358), .S(n5357), .CO(n5356));
Q_AD01HF U750 ( .A0(_zygsfis_ib_service_data_ack[3]), .B0(n5356), .S(n5355), .CO(n5354));
Q_FDP0 \_zygsfis_ib_service_data_ack_REG[3] ( .CK(_zySfifoF2_call), .D(n5355), .Q(_zygsfis_ib_service_data_ack[3]), .QN( ));
Q_FDP0 \_zygsfis_ib_service_data_ack_REG[2] ( .CK(_zySfifoF2_call), .D(n5357), .Q(_zygsfis_ib_service_data_ack[2]), .QN( ));
Q_FDP0 \_zygsfis_ib_service_data_ack_REG[1] ( .CK(_zySfifoF2_call), .D(n5359), .Q(_zygsfis_ib_service_data_ack[1]), .QN( ));
Q_FDP0 \_zygsfis_ib_service_data_ack_REG[0] ( .CK(_zySfifoF2_call), .D(n5360), .Q(_zygsfis_ib_service_data_ack[0]), .QN(n5360));
Q_FDP0 _zygsfis_ib_service_data_eos_REG  ( .CK(_zySfifoF2_call), .D(_zySfifoF2_iarg[0]), .Q(_zygsfis_ib_service_data_eos), .QN( ));
Q_AD01HF U756 ( .A0(_zygsfis_get_config_data_wptr[1]), .B0(_zygsfis_get_config_data_wptr[0]), .S(n5352), .CO(n5351));
Q_AD01HF U757 ( .A0(_zygsfis_get_config_data_wptr[2]), .B0(n5351), .S(n5350), .CO(n5349));
Q_AD01HF U758 ( .A0(_zygsfis_get_config_data_wptr[3]), .B0(n5349), .S(n5348), .CO(n5347));
Q_FDP0 \_zygsfis_get_config_data_wptr_REG[3] ( .CK(_zySfifoF1_call), .D(n5348), .Q(_zygsfis_get_config_data_wptr[3]), .QN( ));
Q_FDP0 \_zygsfis_get_config_data_wptr_REG[2] ( .CK(_zySfifoF1_call), .D(n5350), .Q(_zygsfis_get_config_data_wptr[2]), .QN( ));
Q_FDP0 \_zygsfis_get_config_data_wptr_REG[1] ( .CK(_zySfifoF1_call), .D(n5352), .Q(_zygsfis_get_config_data_wptr[1]), .QN( ));
Q_FDP0 \_zygsfis_get_config_data_wptr_REG[0] ( .CK(_zySfifoF1_call), .D(n5353), .Q(_zygsfis_get_config_data_wptr[0]), .QN(n5353));
Q_AD01HF U763 ( .A0(_zygsfis_get_config_data_ack[1]), .B0(_zygsfis_get_config_data_ack[0]), .S(n5345), .CO(n5344));
Q_AD01HF U764 ( .A0(_zygsfis_get_config_data_ack[2]), .B0(n5344), .S(n5343), .CO(n5342));
Q_AD01HF U765 ( .A0(_zygsfis_get_config_data_ack[3]), .B0(n5342), .S(n5341), .CO(n5340));
Q_FDP0 \_zygsfis_get_config_data_ack_REG[3] ( .CK(_zySfifoF0_call), .D(n5341), .Q(_zygsfis_get_config_data_ack[3]), .QN( ));
Q_FDP0 \_zygsfis_get_config_data_ack_REG[2] ( .CK(_zySfifoF0_call), .D(n5343), .Q(_zygsfis_get_config_data_ack[2]), .QN( ));
Q_FDP0 \_zygsfis_get_config_data_ack_REG[1] ( .CK(_zySfifoF0_call), .D(n5345), .Q(_zygsfis_get_config_data_ack[1]), .QN( ));
Q_FDP0 \_zygsfis_get_config_data_ack_REG[0] ( .CK(_zySfifoF0_call), .D(n5346), .Q(_zygsfis_get_config_data_ack[0]), .QN(n5346));
Q_FDP0 _zygsfis_get_config_data_eos_REG  ( .CK(_zySfifoF0_call), .D(_zySfifoF0_iarg[0]), .Q(_zygsfis_get_config_data_eos), .QN( ));
Q_OR02 U771 ( .A0(n5330), .A1(_zyM2L253_pbcFsm2_s[0]), .Z(n5318));
Q_OR02 U772 ( .A0(_zyM2L253_pbcFsm2_s[1]), .A1(_zyM2L253_pbcFsm2_s[0]), .Z(n5294));
Q_INV U773 ( .A(n5294), .Z(n5317));
Q_MX02 U774 ( .S(_zyM2L253_pbcFsm2_s[2]), .A0(n5317), .A1(n5318), .Z(n5316));
Q_INV U775 ( .A(_zyM2L253_pbcFsm2_s[0]), .Z(n5326));
Q_OR02 U776 ( .A0(n5326), .A1(n5337), .Z(n5329));
Q_OR02 U777 ( .A0(n5296), .A1(n5329), .Z(n5315));
Q_INV U778 ( .A(n5315), .Z(n5320));
Q_INV U779 ( .A(n5305), .Z(n5321));
Q_AO21 U780 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n5337), .B0(_zyM2L253_pbcFsm2_s[1]), .Z(n5301));
Q_AN02 U781 ( .A0(_zyM2L253_pbcFsm2_s[2]), .A1(n5307), .Z(n5314));
Q_XOR2 U782 ( .A0(_zyM2L253_pbcFsm2_s[1]), .A1(n5326), .Z(n5286));
Q_OR02 U783 ( .A0(n5276), .A1(_zyM2L253_pbcFsm2_s[1]), .Z(n5313));
Q_OA21 U784 ( .A0(n5285), .A1(_zyM2L253_pbcFsm2_s[2]), .B0(n5293), .Z(n5312));
Q_INV U785 ( .A(n5338), .Z(n5311));
Q_OA21 U786 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n5311), .B0(_zyM2L253_pbcFsm2_s[1]), .Z(n5310));
Q_INV U787 ( .A(n5310), .Z(n5309));
Q_OR02 U788 ( .A0(_zyM2L253_pbcFsm2_s[2]), .A1(n5309), .Z(n5308));
Q_AN02 U789 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(_zyM2L253_pbcFsm2_s[1]), .Z(n5307));
Q_OR03 U790 ( .A0(n5307), .A1(n5275), .A2(_zyM2L253_pbcFsm2_s[2]), .Z(n5306));
Q_OR03 U791 ( .A0(n5330), .A1(n5325), .A2(n5276), .Z(n5272));
Q_OR02 U792 ( .A0(n5294), .A1(_zyM2L253_pbcFsm2_s[2]), .Z(n5305));
Q_AN02 U793 ( .A0(n5272), .A1(n5305), .Z(n5304));
Q_AO21 U794 ( .A0(n5328), .A1(_zyM2L253_pbcFsm2_s[1]), .B0(n5282), .Z(n5303));
Q_OR02 U795 ( .A0(_zyM2L253_pbcFsm2_s[2]), .A1(n5303), .Z(n5302));
Q_INV U796 ( .A(n5282), .Z(n5292));
Q_OR02 U797 ( .A0(n5301), .A1(_zyM2L253_pbcFsm2_s[2]), .Z(n5300));
Q_AN02 U798 ( .A0(n5291), .A1(n5300), .Z(n5299));
Q_INV U799 ( .A(n5272), .Z(n5336));
Q_INV U800 ( .A(n5333), .Z(n5298));
Q_OR02 U801 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n5298), .Z(n5288));
Q_OR02 U802 ( .A0(n5296), .A1(n5288), .Z(n5297));
Q_OR03 U803 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3968), .A2(n5296), .Z(n5295));
Q_OR02 U804 ( .A0(_zyM2L253_pbcFsm2_s[2]), .A1(_zyM2L253_pbcFsm2_s[1]), .Z(n5296));
Q_OR02 U805 ( .A0(n5276), .A1(n5294), .Z(n5293));
Q_INV U806 ( .A(n5293), .Z(n5335));
Q_OR02 U807 ( .A0(n5276), .A1(n5292), .Z(n5291));
Q_INV U808 ( .A(n5291), .Z(n5334));
Q_NR02 U809 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n5333), .Z(n5290));
Q_NR02 U810 ( .A0(_zyM2L253_pbcFsm2_s[2]), .A1(n5290), .Z(n5289));
Q_INV U811 ( .A(n5288), .Z(n5332));
Q_MX02 U812 ( .S(_zyM2L253_pbcFsm2_s[2]), .A0(n5290), .A1(_zyM2L253_pbcFsm2_s[0]), .Z(n5287));
Q_INV U813 ( .A(n5287), .Z(n5331));
Q_AN02 U814 ( .A0(n5276), .A1(n5285), .Z(n5324));
Q_OR02 U815 ( .A0(n5286), .A1(n5276), .Z(n5283));
Q_OR02 U816 ( .A0(n5327), .A1(n5330), .Z(n5285));
Q_ND02 U817 ( .A0(n5285), .A1(n54), .Z(n5284));
Q_OA21 U818 ( .A0(n5284), .A1(_zyM2L253_pbcFsm2_s[2]), .B0(n5283), .Z(n5323));
Q_AO21 U819 ( .A0(n5325), .A1(_zyM2L253_pbcFsm2_s[1]), .B0(n5282), .Z(n5281));
Q_AN02 U820 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n5330), .Z(n5282));
Q_AO21 U821 ( .A0(n5339), .A1(_zyM2L253_pbcFsm2_s[0]), .B0(n5280), .Z(n5279));
Q_INV U822 ( .A(n5328), .Z(n5280));
Q_MX02 U823 ( .S(_zyM2L253_pbcFsm2_s[1]), .A0(n5329), .A1(n5279), .Z(n5278));
Q_INV U824 ( .A(n5278), .Z(n5277));
Q_MX02 U825 ( .S(_zyM2L253_pbcFsm2_s[2]), .A0(n5277), .A1(n5281), .Z(n5322));
Q_OR02 U826 ( .A0(n5339), .A1(n5326), .Z(n5327));
Q_OR02 U827 ( .A0(n5338), .A1(_zyM2L253_pbcFsm2_s[0]), .Z(n5328));
Q_AN03 U828 ( .A0(n5327), .A1(n5328), .A2(_zyM2L253_pbcFsm2_s[1]), .Z(n5274));
Q_AN02 U829 ( .A0(n5329), .A1(n5330), .Z(n5275));
Q_OR03 U830 ( .A0(n5274), .A1(n5275), .A2(_zyM2L253_pbcFsm2_s[2]), .Z(n5273));
Q_ND02 U831 ( .A0(n5272), .A1(n5273), .Z(n5271));
Q_FDP0 _zzM2L253_mdxP5_kme_ib_tuser_Dwen5_REG  ( .CK(_zyM2L253_pbcMevClk12), .D(n5320), .Q(_zzM2L253_mdxP5_kme_ib_tuser_Dwen5), .QN( ));
Q_FDP0 _zzM2L253_mdxP5_kme_ib_tstrb_Dwen4_REG  ( .CK(_zyM2L253_pbcMevClk12), .D(n5320), .Q(_zzM2L253_mdxP5_kme_ib_tstrb_Dwen4), .QN( ));
Q_FDP0 _zzM2L253_mdxP5_kme_ib_tdata_Dwen3_REG  ( .CK(_zyM2L253_pbcMevClk12), .D(n5320), .Q(_zzM2L253_mdxP5_kme_ib_tdata_Dwen3), .QN( ));
Q_FDP0 _zzM2L253_mdxP5_kme_ib_tlast_Dwen2_REG  ( .CK(_zyM2L253_pbcMevClk12), .D(n5320), .Q(_zzM2L253_mdxP5_kme_ib_tlast_Dwen2), .QN( ));
Q_FDP0 _zzM2L253_mdxP5_kme_ib_tvalid_Dwen1_REG  ( .CK(_zyM2L253_pbcMevClk12), .D(n5320), .Q(_zzM2L253_mdxP5_kme_ib_tvalid_Dwen1), .QN( ));
Q_FDP0 _zzM2L253_mdxP5_error_cntr_Dwen0_REG  ( .CK(_zyM2L253_pbcMevClk12), .D(n5321), .Q(_zzM2L253_mdxP5_error_cntr_Dwen0), .QN( ));
Q_INV U838 ( .A(n5324), .Z(n5270));
Q_OR02 U839 ( .A0(n5323), .A1(n5270), .Z(n5265));
Q_INV U840 ( .A(n5323), .Z(n5269));
Q_OR02 U841 ( .A0(n5269), .A1(n5324), .Z(n5266));
Q_INV U842 ( .A(n5266), .Z(n5268));
Q_MX02 U843 ( .S(n5322), .A0(n5268), .A1(n5265), .Z(n5267));
Q_INV U844 ( .A(n5265), .Z(n5264));
Q_MX02 U845 ( .S(n5322), .A0(n5264), .A1(n5266), .Z(n5263));
Q_OA21 U846 ( .A0(n5323), .A1(n5324), .B0(n5261), .Z(n5262));
Q_INV U847 ( .A(n5322), .Z(n5261));
Q_AN02 U848 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3947), .Z(n5260));
Q_AN02 U849 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3945), .Z(n5259));
Q_AN02 U850 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3943), .Z(n5258));
Q_AN02 U851 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3941), .Z(n5257));
Q_AN02 U852 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3939), .Z(n5256));
Q_AN02 U853 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3937), .Z(n5255));
Q_AN02 U854 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3935), .Z(n5254));
Q_AN02 U855 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3933), .Z(n5253));
Q_AN02 U856 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3931), .Z(n5252));
Q_AN02 U857 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3929), .Z(n5251));
Q_AN02 U858 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3927), .Z(n5250));
Q_AN02 U859 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3925), .Z(n5249));
Q_AN02 U860 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3923), .Z(n5248));
Q_AN02 U861 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3921), .Z(n5247));
Q_AN02 U862 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3919), .Z(n5246));
Q_AN02 U863 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3917), .Z(n5245));
Q_AN02 U864 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3915), .Z(n5244));
Q_AN02 U865 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3913), .Z(n5243));
Q_AN02 U866 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3911), .Z(n5242));
Q_AN02 U867 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3909), .Z(n5241));
Q_AN02 U868 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3907), .Z(n5240));
Q_AN02 U869 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3905), .Z(n5239));
Q_AN02 U870 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3903), .Z(n5238));
Q_AN02 U871 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3901), .Z(n5237));
Q_AN02 U872 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3899), .Z(n5236));
Q_OR02 U873 ( .A0(n5228), .A1(n3897), .Z(n5235));
Q_OR02 U874 ( .A0(n5228), .A1(n3895), .Z(n5234));
Q_OR02 U875 ( .A0(n5228), .A1(n3893), .Z(n5233));
Q_OR02 U876 ( .A0(n5228), .A1(n3891), .Z(n5232));
Q_OR02 U877 ( .A0(n5228), .A1(n3889), .Z(n5231));
Q_AN02 U878 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3887), .Z(n5230));
Q_OR02 U879 ( .A0(n5228), .A1(n3886), .Z(n5229));
Q_INV U880 ( .A(_zyM2L253_pbcFsm2_s[0]), .Z(n5228));
Q_AN02 U881 ( .A0(n5326), .A1(n3865), .Z(n5227));
Q_AN02 U882 ( .A0(n5326), .A1(n3863), .Z(n5226));
Q_AN02 U883 ( .A0(n5326), .A1(n3861), .Z(n5225));
Q_AN02 U884 ( .A0(n5326), .A1(n3859), .Z(n5224));
Q_AN02 U885 ( .A0(n5326), .A1(n3857), .Z(n5223));
Q_AN02 U886 ( .A0(n5326), .A1(n3855), .Z(n5222));
Q_AN02 U887 ( .A0(n5326), .A1(n3853), .Z(n5221));
Q_AN02 U888 ( .A0(n5326), .A1(n3851), .Z(n5220));
Q_AN02 U889 ( .A0(n5326), .A1(n3849), .Z(n5219));
Q_AN02 U890 ( .A0(n5326), .A1(n3847), .Z(n5218));
Q_AN02 U891 ( .A0(n5326), .A1(n3845), .Z(n5217));
Q_AN02 U892 ( .A0(n5326), .A1(n3843), .Z(n5216));
Q_AN02 U893 ( .A0(n5326), .A1(n3841), .Z(n5215));
Q_AN02 U894 ( .A0(n5326), .A1(n3839), .Z(n5214));
Q_AN02 U895 ( .A0(n5326), .A1(n3837), .Z(n5213));
Q_AN02 U896 ( .A0(n5326), .A1(n3835), .Z(n5212));
Q_AN02 U897 ( .A0(n5326), .A1(n3833), .Z(n5211));
Q_AN02 U898 ( .A0(n5326), .A1(n3831), .Z(n5210));
Q_AN02 U899 ( .A0(n5326), .A1(n3829), .Z(n5209));
Q_AN02 U900 ( .A0(n5326), .A1(n3827), .Z(n5208));
Q_AN02 U901 ( .A0(n5326), .A1(n3825), .Z(n5207));
Q_AN02 U902 ( .A0(n5326), .A1(n3823), .Z(n5206));
Q_AN02 U903 ( .A0(n5326), .A1(n3821), .Z(n5205));
Q_AN02 U904 ( .A0(n5326), .A1(n3819), .Z(n5204));
Q_AN02 U905 ( .A0(n5326), .A1(n3817), .Z(n5203));
Q_AN02 U906 ( .A0(n5326), .A1(n3815), .Z(n5202));
Q_OR02 U907 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3813), .Z(n5201));
Q_OR02 U908 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3811), .Z(n5200));
Q_OR02 U909 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3809), .Z(n5199));
Q_OR02 U910 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3807), .Z(n5198));
Q_OR02 U911 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3805), .Z(n5197));
Q_OR02 U912 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3804), .Z(n5196));
Q_AN02 U913 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3783), .Z(n5195));
Q_AN02 U914 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3781), .Z(n5194));
Q_AN02 U915 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3779), .Z(n5193));
Q_AN02 U916 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3777), .Z(n5192));
Q_AN02 U917 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3775), .Z(n5191));
Q_AN02 U918 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3773), .Z(n5190));
Q_AN02 U919 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3771), .Z(n5189));
Q_AN02 U920 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3769), .Z(n5188));
Q_AN02 U921 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3767), .Z(n5187));
Q_AN02 U922 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3765), .Z(n5186));
Q_AN02 U923 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3763), .Z(n5185));
Q_AN02 U924 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3761), .Z(n5184));
Q_AN02 U925 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3759), .Z(n5183));
Q_AN02 U926 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3757), .Z(n5182));
Q_AN02 U927 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3755), .Z(n5181));
Q_AN02 U928 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3753), .Z(n5180));
Q_AN02 U929 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3751), .Z(n5179));
Q_AN02 U930 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3749), .Z(n5178));
Q_AN02 U931 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3747), .Z(n5177));
Q_AN02 U932 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3745), .Z(n5176));
Q_AN02 U933 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3743), .Z(n5175));
Q_AN02 U934 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3741), .Z(n5174));
Q_AN02 U935 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3739), .Z(n5173));
Q_AN02 U936 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3737), .Z(n5172));
Q_AN02 U937 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3735), .Z(n5171));
Q_OR02 U938 ( .A0(n5163), .A1(n3733), .Z(n5170));
Q_OR02 U939 ( .A0(n5163), .A1(n3731), .Z(n5169));
Q_OR02 U940 ( .A0(n5163), .A1(n3729), .Z(n5168));
Q_OR02 U941 ( .A0(n5163), .A1(n3727), .Z(n5167));
Q_OR02 U942 ( .A0(n5163), .A1(n3725), .Z(n5166));
Q_AN02 U943 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3723), .Z(n5165));
Q_OR02 U944 ( .A0(n5163), .A1(n3722), .Z(n5164));
Q_AN02 U945 ( .A0(n5326), .A1(n3701), .Z(n5162));
Q_AN02 U946 ( .A0(n5326), .A1(n3699), .Z(n5161));
Q_AN02 U947 ( .A0(n5326), .A1(n3697), .Z(n5160));
Q_AN02 U948 ( .A0(n5326), .A1(n3695), .Z(n5159));
Q_AN02 U949 ( .A0(n5326), .A1(n3693), .Z(n5158));
Q_AN02 U950 ( .A0(n5326), .A1(n3691), .Z(n5157));
Q_AN02 U951 ( .A0(n5326), .A1(n3689), .Z(n5156));
Q_AN02 U952 ( .A0(n5326), .A1(n3687), .Z(n5155));
Q_AN02 U953 ( .A0(n5326), .A1(n3685), .Z(n5154));
Q_AN02 U954 ( .A0(n5326), .A1(n3683), .Z(n5153));
Q_AN02 U955 ( .A0(n5326), .A1(n3681), .Z(n5152));
Q_AN02 U956 ( .A0(n5326), .A1(n3679), .Z(n5151));
Q_AN02 U957 ( .A0(n5326), .A1(n3677), .Z(n5150));
Q_AN02 U958 ( .A0(n5326), .A1(n3675), .Z(n5149));
Q_AN02 U959 ( .A0(n5326), .A1(n3673), .Z(n5148));
Q_AN02 U960 ( .A0(n5326), .A1(n3671), .Z(n5147));
Q_AN02 U961 ( .A0(n5326), .A1(n3669), .Z(n5146));
Q_AN02 U962 ( .A0(n5326), .A1(n3667), .Z(n5145));
Q_AN02 U963 ( .A0(n5326), .A1(n3665), .Z(n5144));
Q_AN02 U964 ( .A0(n5326), .A1(n3663), .Z(n5143));
Q_AN02 U965 ( .A0(n5326), .A1(n3661), .Z(n5142));
Q_AN02 U966 ( .A0(n5326), .A1(n3659), .Z(n5141));
Q_AN02 U967 ( .A0(n5326), .A1(n3657), .Z(n5140));
Q_AN02 U968 ( .A0(n5326), .A1(n3655), .Z(n5139));
Q_AN02 U969 ( .A0(n5326), .A1(n3653), .Z(n5138));
Q_AN02 U970 ( .A0(n5326), .A1(n3651), .Z(n5137));
Q_AN02 U971 ( .A0(n5326), .A1(n3649), .Z(n5136));
Q_AN02 U972 ( .A0(n5326), .A1(n3647), .Z(n5135));
Q_OR02 U973 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3645), .Z(n5134));
Q_OR02 U974 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3643), .Z(n5133));
Q_AN02 U975 ( .A0(n5326), .A1(n3641), .Z(n5132));
Q_OR02 U976 ( .A0(_zyM2L253_pbcFsm2_s[0]), .A1(n3640), .Z(n5131));
Q_AN02 U977 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[279]), .Z(n5130));
Q_AN02 U978 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[278]), .Z(n5129));
Q_AN02 U979 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[277]), .Z(n5128));
Q_AN02 U980 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[276]), .Z(n5127));
Q_AN02 U981 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[275]), .Z(n5126));
Q_AN02 U982 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[274]), .Z(n5125));
Q_AN02 U983 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[273]), .Z(n5124));
Q_AN02 U984 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[272]), .Z(n5123));
Q_AN02 U985 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[271]), .Z(n5122));
Q_AN02 U986 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[270]), .Z(n5121));
Q_AN02 U987 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[269]), .Z(n5120));
Q_AN02 U988 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[268]), .Z(n5119));
Q_AN02 U989 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[267]), .Z(n5118));
Q_AN02 U990 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[266]), .Z(n5117));
Q_AN02 U991 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[265]), .Z(n5116));
Q_AN02 U992 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[264]), .Z(n5115));
Q_AN02 U993 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[263]), .Z(n5114));
Q_AN02 U994 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[262]), .Z(n5113));
Q_AN02 U995 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[261]), .Z(n5112));
Q_AN02 U996 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[260]), .Z(n5111));
Q_AN02 U997 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[259]), .Z(n5110));
Q_AN02 U998 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[258]), .Z(n5109));
Q_AN02 U999 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[257]), .Z(n5108));
Q_AN02 U1000 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[256]), .Z(n5107));
Q_AN02 U1001 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[255]), .Z(n5106));
Q_AN02 U1002 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[254]), .Z(n5105));
Q_AN02 U1003 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[253]), .Z(n5104));
Q_AN02 U1004 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[252]), .Z(n5103));
Q_AN02 U1005 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[251]), .Z(n5102));
Q_AN02 U1006 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[250]), .Z(n5101));
Q_AN02 U1007 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[249]), .Z(n5100));
Q_AN02 U1008 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[248]), .Z(n5099));
Q_AN02 U1009 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[247]), .Z(n5098));
Q_AN02 U1010 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[246]), .Z(n5097));
Q_AN02 U1011 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[245]), .Z(n5096));
Q_AN02 U1012 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[244]), .Z(n5095));
Q_AN02 U1013 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[243]), .Z(n5094));
Q_AN02 U1014 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[242]), .Z(n5093));
Q_AN02 U1015 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[241]), .Z(n5092));
Q_AN02 U1016 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[240]), .Z(n5091));
Q_AN02 U1017 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[239]), .Z(n5090));
Q_AN02 U1018 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[238]), .Z(n5089));
Q_AN02 U1019 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[237]), .Z(n5088));
Q_AN02 U1020 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[236]), .Z(n5087));
Q_AN02 U1021 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[235]), .Z(n5086));
Q_AN02 U1022 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[234]), .Z(n5085));
Q_AN02 U1023 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[233]), .Z(n5084));
Q_AN02 U1024 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[232]), .Z(n5083));
Q_AN02 U1025 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[231]), .Z(n5082));
Q_AN02 U1026 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[230]), .Z(n5081));
Q_AN02 U1027 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[229]), .Z(n5080));
Q_AN02 U1028 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[228]), .Z(n5079));
Q_AN02 U1029 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[227]), .Z(n5078));
Q_AN02 U1030 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[226]), .Z(n5077));
Q_AN02 U1031 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[225]), .Z(n5076));
Q_AN02 U1032 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[224]), .Z(n5075));
Q_AN02 U1033 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[223]), .Z(n5074));
Q_AN02 U1034 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[222]), .Z(n5073));
Q_AN02 U1035 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[221]), .Z(n5072));
Q_AN02 U1036 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[220]), .Z(n5071));
Q_AN02 U1037 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[219]), .Z(n5070));
Q_AN02 U1038 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[218]), .Z(n5069));
Q_AN02 U1039 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[217]), .Z(n5068));
Q_AN02 U1040 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[216]), .Z(n5067));
Q_AN02 U1041 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[215]), .Z(n5066));
Q_AN02 U1042 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[214]), .Z(n5065));
Q_AN02 U1043 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[213]), .Z(n5064));
Q_AN02 U1044 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[212]), .Z(n5063));
Q_AN02 U1045 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[211]), .Z(n5062));
Q_AN02 U1046 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[210]), .Z(n5061));
Q_AN02 U1047 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[209]), .Z(n5060));
Q_AN02 U1048 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[208]), .Z(n5059));
Q_AN02 U1049 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[207]), .Z(n5058));
Q_AN02 U1050 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[206]), .Z(n5057));
Q_AN02 U1051 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[205]), .Z(n5056));
Q_AN02 U1052 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[204]), .Z(n5055));
Q_AN02 U1053 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[203]), .Z(n5054));
Q_AN02 U1054 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[202]), .Z(n5053));
Q_AN02 U1055 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[201]), .Z(n5052));
Q_AN02 U1056 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[200]), .Z(n5051));
Q_AN02 U1057 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[199]), .Z(n5050));
Q_AN02 U1058 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[198]), .Z(n5049));
Q_AN02 U1059 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[197]), .Z(n5048));
Q_AN02 U1060 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[196]), .Z(n5047));
Q_AN02 U1061 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[195]), .Z(n5046));
Q_AN02 U1062 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[194]), .Z(n5045));
Q_AN02 U1063 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[193]), .Z(n5044));
Q_AN02 U1064 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[192]), .Z(n5043));
Q_AN02 U1065 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[191]), .Z(n5042));
Q_AN02 U1066 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[190]), .Z(n5041));
Q_AN02 U1067 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[189]), .Z(n5040));
Q_AN02 U1068 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[188]), .Z(n5039));
Q_AN02 U1069 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[187]), .Z(n5038));
Q_AN02 U1070 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[186]), .Z(n5037));
Q_AN02 U1071 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[185]), .Z(n5036));
Q_AN02 U1072 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[184]), .Z(n5035));
Q_AN02 U1073 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[183]), .Z(n5034));
Q_AN02 U1074 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[182]), .Z(n5033));
Q_AN02 U1075 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[181]), .Z(n5032));
Q_AN02 U1076 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[180]), .Z(n5031));
Q_AN02 U1077 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[179]), .Z(n5030));
Q_AN02 U1078 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[178]), .Z(n5029));
Q_AN02 U1079 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[177]), .Z(n5028));
Q_AN02 U1080 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[176]), .Z(n5027));
Q_AN02 U1081 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[175]), .Z(n5026));
Q_AN02 U1082 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[174]), .Z(n5025));
Q_AN02 U1083 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[173]), .Z(n5024));
Q_AN02 U1084 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[172]), .Z(n5023));
Q_AN02 U1085 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[171]), .Z(n5022));
Q_AN02 U1086 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[170]), .Z(n5021));
Q_AN02 U1087 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[169]), .Z(n5020));
Q_AN02 U1088 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[168]), .Z(n5019));
Q_AN02 U1089 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[167]), .Z(n5018));
Q_AN02 U1090 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[166]), .Z(n5017));
Q_AN02 U1091 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[165]), .Z(n5016));
Q_AN02 U1092 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[164]), .Z(n5015));
Q_AN02 U1093 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[163]), .Z(n5014));
Q_AN02 U1094 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[162]), .Z(n5013));
Q_AN02 U1095 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[161]), .Z(n5012));
Q_AN02 U1096 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[160]), .Z(n5011));
Q_AN02 U1097 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[159]), .Z(n5010));
Q_AN02 U1098 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[158]), .Z(n5009));
Q_AN02 U1099 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[157]), .Z(n5008));
Q_AN02 U1100 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[156]), .Z(n5007));
Q_AN02 U1101 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[155]), .Z(n5006));
Q_AN02 U1102 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[154]), .Z(n5005));
Q_AN02 U1103 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[153]), .Z(n5004));
Q_AN02 U1104 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[152]), .Z(n5003));
Q_AN02 U1105 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[151]), .Z(n5002));
Q_AN02 U1106 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[150]), .Z(n5001));
Q_AN02 U1107 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[149]), .Z(n5000));
Q_AN02 U1108 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[148]), .Z(n4999));
Q_AN02 U1109 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[147]), .Z(n4998));
Q_AN02 U1110 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[146]), .Z(n4997));
Q_AN02 U1111 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[145]), .Z(n4996));
Q_AN02 U1112 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[144]), .Z(n4995));
Q_AN02 U1113 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[143]), .Z(n4994));
Q_AN02 U1114 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[142]), .Z(n4993));
Q_AN02 U1115 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[141]), .Z(n4992));
Q_AN02 U1116 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[140]), .Z(n4991));
Q_AN02 U1117 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[139]), .Z(n4990));
Q_AN02 U1118 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[138]), .Z(n4989));
Q_AN02 U1119 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[137]), .Z(n4988));
Q_AN02 U1120 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[136]), .Z(n4987));
Q_AN02 U1121 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[135]), .Z(n4986));
Q_AN02 U1122 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[134]), .Z(n4985));
Q_AN02 U1123 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[133]), .Z(n4984));
Q_AN02 U1124 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[132]), .Z(n4983));
Q_AN02 U1125 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[131]), .Z(n4982));
Q_AN02 U1126 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[130]), .Z(n4981));
Q_AN02 U1127 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[129]), .Z(n4980));
Q_AN02 U1128 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[128]), .Z(n4979));
Q_AN02 U1129 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[127]), .Z(n4978));
Q_AN02 U1130 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[126]), .Z(n4977));
Q_AN02 U1131 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[125]), .Z(n4976));
Q_AN02 U1132 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[124]), .Z(n4975));
Q_AN02 U1133 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[123]), .Z(n4974));
Q_AN02 U1134 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[122]), .Z(n4973));
Q_AN02 U1135 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[121]), .Z(n4972));
Q_AN02 U1136 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[120]), .Z(n4971));
Q_AN02 U1137 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[119]), .Z(n4970));
Q_AN02 U1138 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[118]), .Z(n4969));
Q_AN02 U1139 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[117]), .Z(n4968));
Q_AN02 U1140 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[116]), .Z(n4967));
Q_AN02 U1141 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[115]), .Z(n4966));
Q_AN02 U1142 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[114]), .Z(n4965));
Q_AN02 U1143 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[113]), .Z(n4964));
Q_AN02 U1144 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[112]), .Z(n4963));
Q_AN02 U1145 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[111]), .Z(n4962));
Q_AN02 U1146 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[110]), .Z(n4961));
Q_AN02 U1147 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[109]), .Z(n4960));
Q_AN02 U1148 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[108]), .Z(n4959));
Q_AN02 U1149 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[107]), .Z(n4958));
Q_AN02 U1150 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[106]), .Z(n4957));
Q_AN02 U1151 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[105]), .Z(n4956));
Q_AN02 U1152 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[104]), .Z(n4955));
Q_AN02 U1153 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[103]), .Z(n4954));
Q_AN02 U1154 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[102]), .Z(n4953));
Q_AN02 U1155 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[101]), .Z(n4952));
Q_AN02 U1156 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[100]), .Z(n4951));
Q_AN02 U1157 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[99]), .Z(n4950));
Q_AN02 U1158 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[98]), .Z(n4949));
Q_AN02 U1159 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[97]), .Z(n4948));
Q_AN02 U1160 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[96]), .Z(n4947));
Q_AN02 U1161 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[95]), .Z(n4946));
Q_AN02 U1162 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[94]), .Z(n4945));
Q_AN02 U1163 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[93]), .Z(n4944));
Q_AN02 U1164 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[92]), .Z(n4943));
Q_AN02 U1165 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[91]), .Z(n4942));
Q_AN02 U1166 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[90]), .Z(n4941));
Q_AN02 U1167 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[89]), .Z(n4940));
Q_AN02 U1168 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[88]), .Z(n4939));
Q_AN02 U1169 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[87]), .Z(n4938));
Q_AN02 U1170 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[86]), .Z(n4937));
Q_AN02 U1171 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[85]), .Z(n4936));
Q_AN02 U1172 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[84]), .Z(n4935));
Q_AN02 U1173 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[83]), .Z(n4934));
Q_AN02 U1174 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[82]), .Z(n4933));
Q_AN02 U1175 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[81]), .Z(n4932));
Q_AN02 U1176 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[80]), .Z(n4931));
Q_AN02 U1177 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[79]), .Z(n4930));
Q_AN02 U1178 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[78]), .Z(n4929));
Q_AN02 U1179 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[77]), .Z(n4928));
Q_AN02 U1180 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[76]), .Z(n4927));
Q_AN02 U1181 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[75]), .Z(n4926));
Q_AN02 U1182 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[74]), .Z(n4925));
Q_AN02 U1183 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[73]), .Z(n4924));
Q_AN02 U1184 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[72]), .Z(n4923));
Q_AN02 U1185 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[71]), .Z(n4922));
Q_AN02 U1186 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[70]), .Z(n4921));
Q_AN02 U1187 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[69]), .Z(n4920));
Q_AN02 U1188 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[68]), .Z(n4919));
Q_AN02 U1189 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[67]), .Z(n4918));
Q_AN02 U1190 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[66]), .Z(n4917));
Q_AN02 U1191 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[65]), .Z(n4916));
Q_AN02 U1192 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[64]), .Z(n4915));
Q_AN02 U1193 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[63]), .Z(n4914));
Q_AN02 U1194 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[62]), .Z(n4913));
Q_AN02 U1195 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[61]), .Z(n4912));
Q_AN02 U1196 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[60]), .Z(n4911));
Q_AN02 U1197 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[59]), .Z(n4910));
Q_AN02 U1198 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[58]), .Z(n4909));
Q_AN02 U1199 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[57]), .Z(n4908));
Q_AN02 U1200 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[56]), .Z(n4907));
Q_AN02 U1201 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[55]), .Z(n4906));
Q_OR02 U1202 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[54]), .Z(n4905));
Q_OR02 U1203 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[53]), .Z(n4904));
Q_OR02 U1204 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[52]), .Z(n4903));
Q_AN02 U1205 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[51]), .Z(n4902));
Q_OR02 U1206 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[50]), .Z(n4901));
Q_AN02 U1207 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[49]), .Z(n4900));
Q_OR02 U1208 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[48]), .Z(n4899));
Q_AN02 U1209 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[47]), .Z(n4898));
Q_OR02 U1210 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[46]), .Z(n4897));
Q_OR02 U1211 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[45]), .Z(n4896));
Q_AN02 U1212 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[44]), .Z(n4895));
Q_OR02 U1213 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[43]), .Z(n4894));
Q_OR02 U1214 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[42]), .Z(n4893));
Q_OR02 U1215 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[41]), .Z(n4892));
Q_AN02 U1216 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[40]), .Z(n4891));
Q_AN02 U1217 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[39]), .Z(n4890));
Q_OR02 U1218 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[38]), .Z(n4889));
Q_OR02 U1219 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[37]), .Z(n4888));
Q_AN02 U1220 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[36]), .Z(n4887));
Q_OR02 U1221 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[35]), .Z(n4886));
Q_AN02 U1222 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[34]), .Z(n4885));
Q_OR02 U1223 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[33]), .Z(n4884));
Q_OR02 U1224 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[32]), .Z(n4883));
Q_AN02 U1225 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[31]), .Z(n4882));
Q_OR02 U1226 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[30]), .Z(n4881));
Q_OR02 U1227 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[29]), .Z(n4880));
Q_AN02 U1228 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[28]), .Z(n4879));
Q_OR02 U1229 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[27]), .Z(n4878));
Q_OR02 U1230 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[26]), .Z(n4877));
Q_OR02 U1231 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[25]), .Z(n4876));
Q_AN02 U1232 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[24]), .Z(n4875));
Q_AN02 U1233 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[23]), .Z(n4874));
Q_OR02 U1234 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[22]), .Z(n4873));
Q_OR02 U1235 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[21]), .Z(n4872));
Q_AN02 U1236 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[20]), .Z(n4871));
Q_OR02 U1237 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[19]), .Z(n4870));
Q_OR02 U1238 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[18]), .Z(n4869));
Q_OR02 U1239 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[17]), .Z(n4868));
Q_OR02 U1240 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[16]), .Z(n4867));
Q_AN02 U1241 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[15]), .Z(n4866));
Q_OR02 U1242 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[14]), .Z(n4865));
Q_OR02 U1243 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[13]), .Z(n4864));
Q_OR02 U1244 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[12]), .Z(n4863));
Q_AN02 U1245 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[11]), .Z(n4862));
Q_OR02 U1246 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[10]), .Z(n4861));
Q_OR02 U1247 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[9]), .Z(n4860));
Q_OR02 U1248 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[8]), .Z(n4859));
Q_AN02 U1249 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[7]), .Z(n4858));
Q_OR02 U1250 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[6]), .Z(n4857));
Q_OR02 U1251 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[5]), .Z(n4856));
Q_AN02 U1252 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[4]), .Z(n4855));
Q_OR02 U1253 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[3]), .Z(n4854));
Q_OR02 U1254 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[2]), .Z(n4853));
Q_OR02 U1255 ( .A0(n5298), .A1(_zyictd_sysfunc_36_L264_3[1]), .Z(n4852));
Q_AN02 U1256 ( .A0(n5333), .A1(_zyictd_sysfunc_36_L264_3[0]), .Z(n4851));
Q_MX04 U1257 ( .S0(n5289), .S1(n5326), .A0(n3639), .A1(n3638), .A2(n3636), .A3(n3635), .Z(n4850));
Q_AN02 U1258 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[279]), .Z(n4849));
Q_AN02 U1259 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[278]), .Z(n4848));
Q_AN02 U1260 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[277]), .Z(n4847));
Q_AN02 U1261 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[276]), .Z(n4846));
Q_AN02 U1262 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[275]), .Z(n4845));
Q_AN02 U1263 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[274]), .Z(n4844));
Q_AN02 U1264 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[273]), .Z(n4843));
Q_AN02 U1265 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[272]), .Z(n4842));
Q_AN02 U1266 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[271]), .Z(n4841));
Q_AN02 U1267 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[270]), .Z(n4840));
Q_AN02 U1268 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[269]), .Z(n4839));
Q_AN02 U1269 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[268]), .Z(n4838));
Q_AN02 U1270 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[267]), .Z(n4837));
Q_AN02 U1271 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[266]), .Z(n4836));
Q_AN02 U1272 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[265]), .Z(n4835));
Q_AN02 U1273 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[264]), .Z(n4834));
Q_AN02 U1274 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[263]), .Z(n4833));
Q_AN02 U1275 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[262]), .Z(n4832));
Q_AN02 U1276 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[261]), .Z(n4831));
Q_AN02 U1277 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[260]), .Z(n4830));
Q_AN02 U1278 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[259]), .Z(n4829));
Q_AN02 U1279 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[258]), .Z(n4828));
Q_AN02 U1280 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[257]), .Z(n4827));
Q_AN02 U1281 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[256]), .Z(n4826));
Q_AN02 U1282 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[255]), .Z(n4825));
Q_AN02 U1283 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[254]), .Z(n4824));
Q_AN02 U1284 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[253]), .Z(n4823));
Q_AN02 U1285 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[252]), .Z(n4822));
Q_AN02 U1286 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[251]), .Z(n4821));
Q_AN02 U1287 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[250]), .Z(n4820));
Q_AN02 U1288 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[249]), .Z(n4819));
Q_AN02 U1289 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[248]), .Z(n4818));
Q_AN02 U1290 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[247]), .Z(n4817));
Q_AN02 U1291 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[246]), .Z(n4816));
Q_AN02 U1292 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[245]), .Z(n4815));
Q_AN02 U1293 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[244]), .Z(n4814));
Q_AN02 U1294 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[243]), .Z(n4813));
Q_AN02 U1295 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[242]), .Z(n4812));
Q_AN02 U1296 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[241]), .Z(n4811));
Q_AN02 U1297 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[240]), .Z(n4810));
Q_AN02 U1298 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[239]), .Z(n4809));
Q_AN02 U1299 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[238]), .Z(n4808));
Q_AN02 U1300 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[237]), .Z(n4807));
Q_AN02 U1301 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[236]), .Z(n4806));
Q_AN02 U1302 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[235]), .Z(n4805));
Q_AN02 U1303 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[234]), .Z(n4804));
Q_AN02 U1304 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[233]), .Z(n4803));
Q_AN02 U1305 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[232]), .Z(n4802));
Q_AN02 U1306 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[231]), .Z(n4801));
Q_AN02 U1307 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[230]), .Z(n4800));
Q_AN02 U1308 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[229]), .Z(n4799));
Q_AN02 U1309 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[228]), .Z(n4798));
Q_AN02 U1310 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[227]), .Z(n4797));
Q_AN02 U1311 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[226]), .Z(n4796));
Q_AN02 U1312 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[225]), .Z(n4795));
Q_AN02 U1313 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[224]), .Z(n4794));
Q_AN02 U1314 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[223]), .Z(n4793));
Q_AN02 U1315 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[222]), .Z(n4792));
Q_AN02 U1316 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[221]), .Z(n4791));
Q_AN02 U1317 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[220]), .Z(n4790));
Q_AN02 U1318 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[219]), .Z(n4789));
Q_AN02 U1319 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[218]), .Z(n4788));
Q_AN02 U1320 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[217]), .Z(n4787));
Q_AN02 U1321 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[216]), .Z(n4786));
Q_AN02 U1322 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[215]), .Z(n4785));
Q_AN02 U1323 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[214]), .Z(n4784));
Q_AN02 U1324 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[213]), .Z(n4783));
Q_AN02 U1325 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[212]), .Z(n4782));
Q_AN02 U1326 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[211]), .Z(n4781));
Q_AN02 U1327 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[210]), .Z(n4780));
Q_AN02 U1328 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[209]), .Z(n4779));
Q_AN02 U1329 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[208]), .Z(n4778));
Q_AN02 U1330 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[207]), .Z(n4777));
Q_AN02 U1331 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[206]), .Z(n4776));
Q_AN02 U1332 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[205]), .Z(n4775));
Q_AN02 U1333 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[204]), .Z(n4774));
Q_AN02 U1334 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[203]), .Z(n4773));
Q_AN02 U1335 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[202]), .Z(n4772));
Q_AN02 U1336 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[201]), .Z(n4771));
Q_AN02 U1337 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[200]), .Z(n4770));
Q_AN02 U1338 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[199]), .Z(n4769));
Q_AN02 U1339 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[198]), .Z(n4768));
Q_AN02 U1340 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[197]), .Z(n4767));
Q_AN02 U1341 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[196]), .Z(n4766));
Q_AN02 U1342 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[195]), .Z(n4765));
Q_AN02 U1343 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[194]), .Z(n4764));
Q_AN02 U1344 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[193]), .Z(n4763));
Q_AN02 U1345 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[192]), .Z(n4762));
Q_AN02 U1346 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[191]), .Z(n4761));
Q_AN02 U1347 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[190]), .Z(n4760));
Q_AN02 U1348 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[189]), .Z(n4759));
Q_AN02 U1349 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[188]), .Z(n4758));
Q_AN02 U1350 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[187]), .Z(n4757));
Q_AN02 U1351 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[186]), .Z(n4756));
Q_AN02 U1352 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[185]), .Z(n4755));
Q_AN02 U1353 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[184]), .Z(n4754));
Q_AN02 U1354 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[183]), .Z(n4753));
Q_AN02 U1355 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[182]), .Z(n4752));
Q_AN02 U1356 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[181]), .Z(n4751));
Q_AN02 U1357 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[180]), .Z(n4750));
Q_AN02 U1358 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[179]), .Z(n4749));
Q_AN02 U1359 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[178]), .Z(n4748));
Q_AN02 U1360 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[177]), .Z(n4747));
Q_AN02 U1361 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[176]), .Z(n4746));
Q_AN02 U1362 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[175]), .Z(n4745));
Q_AN02 U1363 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[174]), .Z(n4744));
Q_AN02 U1364 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[173]), .Z(n4743));
Q_AN02 U1365 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[172]), .Z(n4742));
Q_AN02 U1366 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[171]), .Z(n4741));
Q_AN02 U1367 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[170]), .Z(n4740));
Q_AN02 U1368 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[169]), .Z(n4739));
Q_AN02 U1369 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[168]), .Z(n4738));
Q_AN02 U1370 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[167]), .Z(n4737));
Q_AN02 U1371 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[166]), .Z(n4736));
Q_AN02 U1372 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[165]), .Z(n4735));
Q_AN02 U1373 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[164]), .Z(n4734));
Q_AN02 U1374 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[163]), .Z(n4733));
Q_AN02 U1375 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[162]), .Z(n4732));
Q_AN02 U1376 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[161]), .Z(n4731));
Q_AN02 U1377 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[160]), .Z(n4730));
Q_AN02 U1378 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[159]), .Z(n4729));
Q_AN02 U1379 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[158]), .Z(n4728));
Q_AN02 U1380 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[157]), .Z(n4727));
Q_AN02 U1381 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[156]), .Z(n4726));
Q_AN02 U1382 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[155]), .Z(n4725));
Q_AN02 U1383 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[154]), .Z(n4724));
Q_AN02 U1384 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[153]), .Z(n4723));
Q_AN02 U1385 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[152]), .Z(n4722));
Q_AN02 U1386 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[151]), .Z(n4721));
Q_AN02 U1387 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[150]), .Z(n4720));
Q_AN02 U1388 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[149]), .Z(n4719));
Q_AN02 U1389 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[148]), .Z(n4718));
Q_AN02 U1390 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[147]), .Z(n4717));
Q_AN02 U1391 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[146]), .Z(n4716));
Q_AN02 U1392 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[145]), .Z(n4715));
Q_AN02 U1393 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[144]), .Z(n4714));
Q_AN02 U1394 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[143]), .Z(n4713));
Q_AN02 U1395 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[142]), .Z(n4712));
Q_AN02 U1396 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[141]), .Z(n4711));
Q_AN02 U1397 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[140]), .Z(n4710));
Q_AN02 U1398 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[139]), .Z(n4709));
Q_AN02 U1399 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[138]), .Z(n4708));
Q_AN02 U1400 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[137]), .Z(n4707));
Q_AN02 U1401 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[136]), .Z(n4706));
Q_AN02 U1402 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[135]), .Z(n4705));
Q_AN02 U1403 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[134]), .Z(n4704));
Q_AN02 U1404 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[133]), .Z(n4703));
Q_AN02 U1405 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[132]), .Z(n4702));
Q_AN02 U1406 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[131]), .Z(n4701));
Q_AN02 U1407 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[130]), .Z(n4700));
Q_AN02 U1408 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[129]), .Z(n4699));
Q_AN02 U1409 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[128]), .Z(n4698));
Q_AN02 U1410 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[127]), .Z(n4697));
Q_AN02 U1411 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[126]), .Z(n4696));
Q_AN02 U1412 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[125]), .Z(n4695));
Q_AN02 U1413 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[124]), .Z(n4694));
Q_AN02 U1414 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[123]), .Z(n4693));
Q_AN02 U1415 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[122]), .Z(n4692));
Q_AN02 U1416 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[121]), .Z(n4691));
Q_AN02 U1417 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[120]), .Z(n4690));
Q_AN02 U1418 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[119]), .Z(n4689));
Q_AN02 U1419 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[118]), .Z(n4688));
Q_AN02 U1420 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[117]), .Z(n4687));
Q_AN02 U1421 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[116]), .Z(n4686));
Q_AN02 U1422 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[115]), .Z(n4685));
Q_AN02 U1423 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[114]), .Z(n4684));
Q_AN02 U1424 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[113]), .Z(n4683));
Q_AN02 U1425 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[112]), .Z(n4682));
Q_AN02 U1426 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[111]), .Z(n4681));
Q_AN02 U1427 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[110]), .Z(n4680));
Q_AN02 U1428 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[109]), .Z(n4679));
Q_AN02 U1429 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[108]), .Z(n4678));
Q_AN02 U1430 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[107]), .Z(n4677));
Q_AN02 U1431 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[106]), .Z(n4676));
Q_AN02 U1432 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[105]), .Z(n4675));
Q_AN02 U1433 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[104]), .Z(n4674));
Q_AN02 U1434 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[103]), .Z(n4673));
Q_AN02 U1435 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[102]), .Z(n4672));
Q_AN02 U1436 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[101]), .Z(n4671));
Q_AN02 U1437 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[100]), .Z(n4670));
Q_AN02 U1438 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[99]), .Z(n4669));
Q_AN02 U1439 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[98]), .Z(n4668));
Q_AN02 U1440 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[97]), .Z(n4667));
Q_AN02 U1441 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[96]), .Z(n4666));
Q_AN02 U1442 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[95]), .Z(n4665));
Q_AN02 U1443 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[94]), .Z(n4664));
Q_AN02 U1444 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[93]), .Z(n4663));
Q_AN02 U1445 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[92]), .Z(n4662));
Q_AN02 U1446 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[91]), .Z(n4661));
Q_AN02 U1447 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[90]), .Z(n4660));
Q_AN02 U1448 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[89]), .Z(n4659));
Q_AN02 U1449 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[88]), .Z(n4658));
Q_AN02 U1450 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[87]), .Z(n4657));
Q_AN02 U1451 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[86]), .Z(n4656));
Q_AN02 U1452 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[85]), .Z(n4655));
Q_AN02 U1453 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[84]), .Z(n4654));
Q_AN02 U1454 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[83]), .Z(n4653));
Q_AN02 U1455 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[82]), .Z(n4652));
Q_AN02 U1456 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[81]), .Z(n4651));
Q_AN02 U1457 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[80]), .Z(n4650));
Q_AN02 U1458 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[79]), .Z(n4649));
Q_AN02 U1459 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[78]), .Z(n4648));
Q_AN02 U1460 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[77]), .Z(n4647));
Q_AN02 U1461 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[76]), .Z(n4646));
Q_AN02 U1462 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[75]), .Z(n4645));
Q_AN02 U1463 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[74]), .Z(n4644));
Q_AN02 U1464 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[73]), .Z(n4643));
Q_AN02 U1465 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[72]), .Z(n4642));
Q_AN02 U1466 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[71]), .Z(n4641));
Q_AN02 U1467 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[70]), .Z(n4640));
Q_AN02 U1468 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[69]), .Z(n4639));
Q_AN02 U1469 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[68]), .Z(n4638));
Q_AN02 U1470 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[67]), .Z(n4637));
Q_AN02 U1471 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[66]), .Z(n4636));
Q_AN02 U1472 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[65]), .Z(n4635));
Q_AN02 U1473 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[64]), .Z(n4634));
Q_AN02 U1474 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[63]), .Z(n4633));
Q_AN02 U1475 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[62]), .Z(n4632));
Q_AN02 U1476 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[61]), .Z(n4631));
Q_AN02 U1477 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[60]), .Z(n4630));
Q_AN02 U1478 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[59]), .Z(n4629));
Q_AN02 U1479 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[58]), .Z(n4628));
Q_AN02 U1480 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[57]), .Z(n4627));
Q_AN02 U1481 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[56]), .Z(n4626));
Q_AN02 U1482 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[55]), .Z(n4625));
Q_MX02 U1483 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[54]), .A1(n5290), .Z(n4624));
Q_MX02 U1484 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[53]), .A1(n5290), .Z(n4623));
Q_MX02 U1485 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[52]), .A1(n5290), .Z(n4622));
Q_AN02 U1486 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[51]), .Z(n4621));
Q_MX02 U1487 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[50]), .A1(n5290), .Z(n4620));
Q_AN02 U1488 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[49]), .Z(n4619));
Q_MX02 U1489 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[48]), .A1(n5290), .Z(n4618));
Q_AN02 U1490 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[47]), .Z(n4617));
Q_MX02 U1491 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[46]), .A1(n5290), .Z(n4616));
Q_MX02 U1492 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[45]), .A1(n5290), .Z(n4615));
Q_AN02 U1493 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[44]), .Z(n4614));
Q_MX02 U1494 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[43]), .A1(n5290), .Z(n4613));
Q_MX02 U1495 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[42]), .A1(n5290), .Z(n4612));
Q_MX02 U1496 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[41]), .A1(n5290), .Z(n4611));
Q_AN02 U1497 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[40]), .Z(n4610));
Q_AN02 U1498 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[39]), .Z(n4609));
Q_MX02 U1499 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[38]), .A1(n5290), .Z(n4608));
Q_MX02 U1500 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[37]), .A1(n5290), .Z(n4607));
Q_AN02 U1501 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[36]), .Z(n4606));
Q_MX02 U1502 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[35]), .A1(n5290), .Z(n4605));
Q_AN02 U1503 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[34]), .Z(n4604));
Q_MX02 U1504 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[33]), .A1(n5290), .Z(n4603));
Q_MX02 U1505 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[32]), .A1(n5290), .Z(n4602));
Q_AN02 U1506 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[31]), .Z(n4601));
Q_MX02 U1507 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[30]), .A1(n5290), .Z(n4600));
Q_MX02 U1508 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[29]), .A1(n5290), .Z(n4599));
Q_AN02 U1509 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[28]), .Z(n4598));
Q_MX02 U1510 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[27]), .A1(n5290), .Z(n4597));
Q_MX02 U1511 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[26]), .A1(n5290), .Z(n4596));
Q_MX02 U1512 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[25]), .A1(n5290), .Z(n4595));
Q_AN02 U1513 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[24]), .Z(n4594));
Q_AN02 U1514 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[23]), .Z(n4593));
Q_MX02 U1515 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[22]), .A1(n5290), .Z(n4592));
Q_MX02 U1516 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[21]), .A1(n5290), .Z(n4591));
Q_AN02 U1517 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[20]), .Z(n4590));
Q_MX02 U1518 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[19]), .A1(n5290), .Z(n4589));
Q_MX02 U1519 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[18]), .A1(n5290), .Z(n4588));
Q_MX02 U1520 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[17]), .A1(n5290), .Z(n4587));
Q_MX02 U1521 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[16]), .A1(n5290), .Z(n4586));
Q_AN02 U1522 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[15]), .Z(n4585));
Q_MX02 U1523 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[14]), .A1(n5290), .Z(n4584));
Q_MX02 U1524 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[13]), .A1(n5290), .Z(n4583));
Q_MX02 U1525 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[12]), .A1(n5290), .Z(n4582));
Q_AN02 U1526 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[11]), .Z(n4581));
Q_MX02 U1527 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[10]), .A1(n5290), .Z(n4580));
Q_MX02 U1528 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[9]), .A1(n5290), .Z(n4579));
Q_MX02 U1529 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[8]), .A1(n5290), .Z(n4578));
Q_AN02 U1530 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[7]), .Z(n4577));
Q_MX02 U1531 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[6]), .A1(n5290), .Z(n4576));
Q_MX02 U1532 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[5]), .A1(n5290), .Z(n4575));
Q_AN02 U1533 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[4]), .Z(n4574));
Q_MX02 U1534 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[3]), .A1(n5290), .Z(n4573));
Q_MX02 U1535 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[2]), .A1(n5290), .Z(n4572));
Q_MX02 U1536 ( .S(n5288), .A0(_zyictd_sysfunc_36_L264_3[1]), .A1(n5290), .Z(n4571));
Q_AN02 U1537 ( .A0(n5332), .A1(_zyictd_sysfunc_36_L264_3[0]), .Z(n4570));
Q_AN02 U1538 ( .A0(n5326), .A1(n4248), .Z(n4569));
Q_AN02 U1539 ( .A0(n5326), .A1(n4247), .Z(n4568));
Q_AN02 U1540 ( .A0(n5326), .A1(n4246), .Z(n4567));
Q_AN02 U1541 ( .A0(n5326), .A1(n4245), .Z(n4566));
Q_AN02 U1542 ( .A0(n5326), .A1(n4244), .Z(n4565));
Q_AN02 U1543 ( .A0(n5326), .A1(n4243), .Z(n4564));
Q_AN02 U1544 ( .A0(n5326), .A1(n4242), .Z(n4563));
Q_AN02 U1545 ( .A0(n5326), .A1(n4241), .Z(n4562));
Q_AN02 U1546 ( .A0(n5326), .A1(n4240), .Z(n4561));
Q_AN02 U1547 ( .A0(n5326), .A1(n4239), .Z(n4560));
Q_AN02 U1548 ( .A0(n5326), .A1(n4238), .Z(n4559));
Q_AN02 U1549 ( .A0(n5326), .A1(n4237), .Z(n4558));
Q_AN02 U1550 ( .A0(n5326), .A1(n4236), .Z(n4557));
Q_AN02 U1551 ( .A0(n5326), .A1(n4235), .Z(n4556));
Q_AN02 U1552 ( .A0(n5326), .A1(n4234), .Z(n4555));
Q_AN02 U1553 ( .A0(n5326), .A1(n4233), .Z(n4554));
Q_AN02 U1554 ( .A0(n5326), .A1(n4232), .Z(n4553));
Q_AN02 U1555 ( .A0(n5326), .A1(n4231), .Z(n4552));
Q_AN02 U1556 ( .A0(n5326), .A1(n4230), .Z(n4551));
Q_AN02 U1557 ( .A0(n5326), .A1(n4229), .Z(n4550));
Q_AN02 U1558 ( .A0(n5326), .A1(n4228), .Z(n4549));
Q_AN02 U1559 ( .A0(n5326), .A1(n4227), .Z(n4548));
Q_AN02 U1560 ( .A0(n5326), .A1(n4226), .Z(n4547));
Q_AN02 U1561 ( .A0(n5326), .A1(n4225), .Z(n4546));
Q_AN02 U1562 ( .A0(n5326), .A1(n4224), .Z(n4545));
Q_AN02 U1563 ( .A0(n5326), .A1(n4223), .Z(n4544));
Q_AN02 U1564 ( .A0(n5326), .A1(n4222), .Z(n4543));
Q_AN02 U1565 ( .A0(n5326), .A1(n4221), .Z(n4542));
Q_AN02 U1566 ( .A0(n5326), .A1(n4220), .Z(n4541));
Q_AN02 U1567 ( .A0(n5326), .A1(n4219), .Z(n4540));
Q_AN02 U1568 ( .A0(n5326), .A1(n4218), .Z(n4539));
Q_AN02 U1569 ( .A0(n5326), .A1(n4217), .Z(n4538));
Q_AN02 U1570 ( .A0(n5326), .A1(n4216), .Z(n4537));
Q_AN02 U1571 ( .A0(n5326), .A1(n4215), .Z(n4536));
Q_AN02 U1572 ( .A0(n5326), .A1(n4214), .Z(n4535));
Q_AN02 U1573 ( .A0(n5326), .A1(n4213), .Z(n4534));
Q_AN02 U1574 ( .A0(n5326), .A1(n4212), .Z(n4533));
Q_AN02 U1575 ( .A0(n5326), .A1(n4211), .Z(n4532));
Q_AN02 U1576 ( .A0(n5326), .A1(n4210), .Z(n4531));
Q_AN02 U1577 ( .A0(n5326), .A1(n4209), .Z(n4530));
Q_AN02 U1578 ( .A0(n5326), .A1(n4208), .Z(n4529));
Q_AN02 U1579 ( .A0(n5326), .A1(n4207), .Z(n4528));
Q_AN02 U1580 ( .A0(n5326), .A1(n4206), .Z(n4527));
Q_AN02 U1581 ( .A0(n5326), .A1(n4205), .Z(n4526));
Q_AN02 U1582 ( .A0(n5326), .A1(n4204), .Z(n4525));
Q_AN02 U1583 ( .A0(n5326), .A1(n4203), .Z(n4524));
Q_AN02 U1584 ( .A0(n5326), .A1(n4202), .Z(n4523));
Q_AN02 U1585 ( .A0(n5326), .A1(n4201), .Z(n4522));
Q_AN02 U1586 ( .A0(n5326), .A1(n4200), .Z(n4521));
Q_AN02 U1587 ( .A0(n5326), .A1(n4199), .Z(n4520));
Q_AN02 U1588 ( .A0(n5326), .A1(n4198), .Z(n4519));
Q_AN02 U1589 ( .A0(n5326), .A1(n4197), .Z(n4518));
Q_AN02 U1590 ( .A0(n5326), .A1(n4196), .Z(n4517));
Q_AN02 U1591 ( .A0(n5326), .A1(n4195), .Z(n4516));
Q_AN02 U1592 ( .A0(n5326), .A1(n4194), .Z(n4515));
Q_AN02 U1593 ( .A0(n5326), .A1(n4193), .Z(n4514));
Q_AN02 U1594 ( .A0(n5326), .A1(n4192), .Z(n4513));
Q_AN02 U1595 ( .A0(n5326), .A1(n4191), .Z(n4512));
Q_AN02 U1596 ( .A0(n5326), .A1(n4190), .Z(n4511));
Q_AN02 U1597 ( .A0(n5326), .A1(n4189), .Z(n4510));
Q_AN02 U1598 ( .A0(n5326), .A1(n4188), .Z(n4509));
Q_AN02 U1599 ( .A0(n5326), .A1(n4187), .Z(n4508));
Q_AN02 U1600 ( .A0(n5326), .A1(n4186), .Z(n4507));
Q_AN02 U1601 ( .A0(n5326), .A1(n4185), .Z(n4506));
Q_AN02 U1602 ( .A0(n5326), .A1(n4184), .Z(n4505));
Q_AN02 U1603 ( .A0(n5326), .A1(n4183), .Z(n4504));
Q_AN02 U1604 ( .A0(n5326), .A1(n4182), .Z(n4503));
Q_AN02 U1605 ( .A0(n5326), .A1(n4181), .Z(n4502));
Q_AN02 U1606 ( .A0(n5326), .A1(n4180), .Z(n4501));
Q_AN02 U1607 ( .A0(n5326), .A1(n4179), .Z(n4500));
Q_AN02 U1608 ( .A0(n5326), .A1(n4178), .Z(n4499));
Q_AN02 U1609 ( .A0(n5326), .A1(n4177), .Z(n4498));
Q_AN02 U1610 ( .A0(n5326), .A1(n4176), .Z(n4497));
Q_AN02 U1611 ( .A0(n5326), .A1(n4175), .Z(n4496));
Q_AN02 U1612 ( .A0(n5326), .A1(n4174), .Z(n4495));
Q_AN02 U1613 ( .A0(n5326), .A1(n4173), .Z(n4494));
Q_AN02 U1614 ( .A0(n5326), .A1(n4172), .Z(n4493));
Q_AN02 U1615 ( .A0(n5326), .A1(n4171), .Z(n4492));
Q_AN02 U1616 ( .A0(n5326), .A1(n4170), .Z(n4491));
Q_AN02 U1617 ( .A0(n5326), .A1(n4169), .Z(n4490));
Q_AN02 U1618 ( .A0(n5326), .A1(n4168), .Z(n4489));
Q_AN02 U1619 ( .A0(n5326), .A1(n4167), .Z(n4488));
Q_AN02 U1620 ( .A0(n5326), .A1(n4166), .Z(n4487));
Q_AN02 U1621 ( .A0(n5326), .A1(n4165), .Z(n4486));
Q_AN02 U1622 ( .A0(n5326), .A1(n4164), .Z(n4485));
Q_AN02 U1623 ( .A0(n5326), .A1(n4163), .Z(n4484));
Q_AN02 U1624 ( .A0(n5326), .A1(n4162), .Z(n4483));
Q_AN02 U1625 ( .A0(n5326), .A1(n4161), .Z(n4482));
Q_AN02 U1626 ( .A0(n5326), .A1(n4160), .Z(n4481));
Q_AN02 U1627 ( .A0(n5326), .A1(n4159), .Z(n4480));
Q_AN02 U1628 ( .A0(n5326), .A1(n4158), .Z(n4479));
Q_AN02 U1629 ( .A0(n5326), .A1(n4157), .Z(n4478));
Q_AN02 U1630 ( .A0(n5326), .A1(n4156), .Z(n4477));
Q_AN02 U1631 ( .A0(n5326), .A1(n4155), .Z(n4476));
Q_AN02 U1632 ( .A0(n5326), .A1(n4154), .Z(n4475));
Q_AN02 U1633 ( .A0(n5326), .A1(n4153), .Z(n4474));
Q_AN02 U1634 ( .A0(n5326), .A1(n4152), .Z(n4473));
Q_AN02 U1635 ( .A0(n5326), .A1(n4151), .Z(n4472));
Q_AN02 U1636 ( .A0(n5326), .A1(n4150), .Z(n4471));
Q_AN02 U1637 ( .A0(n5326), .A1(n4149), .Z(n4470));
Q_AN02 U1638 ( .A0(n5326), .A1(n4148), .Z(n4469));
Q_AN02 U1639 ( .A0(n5326), .A1(n4147), .Z(n4468));
Q_AN02 U1640 ( .A0(n5326), .A1(n4146), .Z(n4467));
Q_AN02 U1641 ( .A0(n5326), .A1(n4145), .Z(n4466));
Q_AN02 U1642 ( .A0(n5326), .A1(n4144), .Z(n4465));
Q_AN02 U1643 ( .A0(n5326), .A1(n4143), .Z(n4464));
Q_AN02 U1644 ( .A0(n5326), .A1(n4142), .Z(n4463));
Q_AN02 U1645 ( .A0(n5326), .A1(n4141), .Z(n4462));
Q_AN02 U1646 ( .A0(n5326), .A1(n4140), .Z(n4461));
Q_AN02 U1647 ( .A0(n5326), .A1(n4139), .Z(n4460));
Q_AN02 U1648 ( .A0(n5326), .A1(n4138), .Z(n4459));
Q_AN02 U1649 ( .A0(n5326), .A1(n4137), .Z(n4458));
Q_AN02 U1650 ( .A0(n5326), .A1(n4136), .Z(n4457));
Q_AN02 U1651 ( .A0(n5326), .A1(n4135), .Z(n4456));
Q_AN02 U1652 ( .A0(n5326), .A1(n4134), .Z(n4455));
Q_AN02 U1653 ( .A0(n5326), .A1(n4133), .Z(n4454));
Q_AN02 U1654 ( .A0(n5326), .A1(n4132), .Z(n4453));
Q_AN02 U1655 ( .A0(n5326), .A1(n4131), .Z(n4452));
Q_AN02 U1656 ( .A0(n5326), .A1(n4130), .Z(n4451));
Q_AN02 U1657 ( .A0(n5326), .A1(n4129), .Z(n4450));
Q_AN02 U1658 ( .A0(n5326), .A1(n4128), .Z(n4449));
Q_AN02 U1659 ( .A0(n5326), .A1(n4127), .Z(n4448));
Q_AN02 U1660 ( .A0(n5326), .A1(n4126), .Z(n4447));
Q_AN02 U1661 ( .A0(n5326), .A1(n4125), .Z(n4446));
Q_AN02 U1662 ( .A0(n5326), .A1(n4124), .Z(n4445));
Q_AN02 U1663 ( .A0(n5326), .A1(n4123), .Z(n4444));
Q_AN02 U1664 ( .A0(n5326), .A1(n4122), .Z(n4443));
Q_AN02 U1665 ( .A0(n5326), .A1(n4121), .Z(n4442));
Q_AN02 U1666 ( .A0(n5326), .A1(n4120), .Z(n4441));
Q_AN02 U1667 ( .A0(n5326), .A1(n4119), .Z(n4440));
Q_AN02 U1668 ( .A0(n5326), .A1(n4118), .Z(n4439));
Q_AN02 U1669 ( .A0(n5326), .A1(n4117), .Z(n4438));
Q_AN02 U1670 ( .A0(n5326), .A1(n4116), .Z(n4437));
Q_AN02 U1671 ( .A0(n5326), .A1(n4115), .Z(n4436));
Q_AN02 U1672 ( .A0(n5326), .A1(n4114), .Z(n4435));
Q_AN02 U1673 ( .A0(n5326), .A1(n4113), .Z(n4434));
Q_AN02 U1674 ( .A0(n5326), .A1(n4112), .Z(n4433));
Q_AN02 U1675 ( .A0(n5326), .A1(n4111), .Z(n4432));
Q_AN02 U1676 ( .A0(n5326), .A1(n4110), .Z(n4431));
Q_AN02 U1677 ( .A0(n5326), .A1(n4109), .Z(n4430));
Q_AN02 U1678 ( .A0(n5326), .A1(n4108), .Z(n4429));
Q_AN02 U1679 ( .A0(n5326), .A1(n4107), .Z(n4428));
Q_AN02 U1680 ( .A0(n5326), .A1(n4106), .Z(n4427));
Q_AN02 U1681 ( .A0(n5326), .A1(n4105), .Z(n4426));
Q_AN02 U1682 ( .A0(n5326), .A1(n4104), .Z(n4425));
Q_AN02 U1683 ( .A0(n5326), .A1(n4103), .Z(n4424));
Q_AN02 U1684 ( .A0(n5326), .A1(n4102), .Z(n4423));
Q_AN02 U1685 ( .A0(n5326), .A1(n4101), .Z(n4422));
Q_AN02 U1686 ( .A0(n5326), .A1(n4100), .Z(n4421));
Q_AN02 U1687 ( .A0(n5326), .A1(n4099), .Z(n4420));
Q_AN02 U1688 ( .A0(n5326), .A1(n4098), .Z(n4419));
Q_AN02 U1689 ( .A0(n5326), .A1(n4097), .Z(n4418));
Q_AN02 U1690 ( .A0(n5326), .A1(n4096), .Z(n4417));
Q_AN02 U1691 ( .A0(n5326), .A1(n4095), .Z(n4416));
Q_AN02 U1692 ( .A0(n5326), .A1(n4094), .Z(n4415));
Q_AN02 U1693 ( .A0(n5326), .A1(n4093), .Z(n4414));
Q_AN02 U1694 ( .A0(n5326), .A1(n4092), .Z(n4413));
Q_AN02 U1695 ( .A0(n5326), .A1(n4091), .Z(n4412));
Q_AN02 U1696 ( .A0(n5326), .A1(n4090), .Z(n4411));
Q_AN02 U1697 ( .A0(n5326), .A1(n4089), .Z(n4410));
Q_AN02 U1698 ( .A0(n5326), .A1(n4088), .Z(n4409));
Q_AN02 U1699 ( .A0(n5326), .A1(n4087), .Z(n4408));
Q_AN02 U1700 ( .A0(n5326), .A1(n4086), .Z(n4407));
Q_AN02 U1701 ( .A0(n5326), .A1(n4085), .Z(n4406));
Q_AN02 U1702 ( .A0(n5326), .A1(n4084), .Z(n4405));
Q_AN02 U1703 ( .A0(n5326), .A1(n4083), .Z(n4404));
Q_AN02 U1704 ( .A0(n5326), .A1(n4082), .Z(n4403));
Q_AN02 U1705 ( .A0(n5326), .A1(n4081), .Z(n4402));
Q_AN02 U1706 ( .A0(n5326), .A1(n4080), .Z(n4401));
Q_AN02 U1707 ( .A0(n5326), .A1(n4079), .Z(n4400));
Q_AN02 U1708 ( .A0(n5326), .A1(n4078), .Z(n4399));
Q_AN02 U1709 ( .A0(n5326), .A1(n4077), .Z(n4398));
Q_AN02 U1710 ( .A0(n5326), .A1(n4076), .Z(n4397));
Q_AN02 U1711 ( .A0(n5326), .A1(n4075), .Z(n4396));
Q_AN02 U1712 ( .A0(n5326), .A1(n4074), .Z(n4395));
Q_AN02 U1713 ( .A0(n5326), .A1(n4073), .Z(n4394));
Q_AN02 U1714 ( .A0(n5326), .A1(n4072), .Z(n4393));
Q_AN02 U1715 ( .A0(n5326), .A1(n4071), .Z(n4392));
Q_AN02 U1716 ( .A0(n5326), .A1(n4070), .Z(n4391));
Q_AN02 U1717 ( .A0(n5326), .A1(n4069), .Z(n4390));
Q_AN02 U1718 ( .A0(n5326), .A1(n4068), .Z(n4389));
Q_AN02 U1719 ( .A0(n5326), .A1(n4067), .Z(n4388));
Q_AN02 U1720 ( .A0(n5326), .A1(n4066), .Z(n4387));
Q_AN02 U1721 ( .A0(n5326), .A1(n4065), .Z(n4386));
Q_AN02 U1722 ( .A0(n5326), .A1(n4064), .Z(n4385));
Q_AN02 U1723 ( .A0(n5326), .A1(n4063), .Z(n4384));
Q_AN02 U1724 ( .A0(n5326), .A1(n4062), .Z(n4383));
Q_AN02 U1725 ( .A0(n5326), .A1(n4061), .Z(n4382));
Q_AN02 U1726 ( .A0(n5326), .A1(n4060), .Z(n4381));
Q_AN02 U1727 ( .A0(n5326), .A1(n4059), .Z(n4380));
Q_AN02 U1728 ( .A0(n5326), .A1(n4058), .Z(n4379));
Q_AN02 U1729 ( .A0(n5326), .A1(n4057), .Z(n4378));
Q_AN02 U1730 ( .A0(n5326), .A1(n4056), .Z(n4377));
Q_AN02 U1731 ( .A0(n5326), .A1(n4055), .Z(n4376));
Q_AN02 U1732 ( .A0(n5326), .A1(n4054), .Z(n4375));
Q_AN02 U1733 ( .A0(n5326), .A1(n4053), .Z(n4374));
Q_AN02 U1734 ( .A0(n5326), .A1(n4052), .Z(n4373));
Q_AN02 U1735 ( .A0(n5326), .A1(n4051), .Z(n4372));
Q_AN02 U1736 ( .A0(n5326), .A1(n4050), .Z(n4371));
Q_AN02 U1737 ( .A0(n5326), .A1(n4049), .Z(n4370));
Q_AN02 U1738 ( .A0(n5326), .A1(n4048), .Z(n4369));
Q_AN02 U1739 ( .A0(n5326), .A1(n4047), .Z(n4368));
Q_AN02 U1740 ( .A0(n5326), .A1(n4046), .Z(n4367));
Q_AN02 U1741 ( .A0(n5326), .A1(n4045), .Z(n4366));
Q_AN02 U1742 ( .A0(n5326), .A1(n4044), .Z(n4365));
Q_AN02 U1743 ( .A0(n5326), .A1(n4043), .Z(n4364));
Q_AN02 U1744 ( .A0(n5326), .A1(n4042), .Z(n4363));
Q_AN02 U1745 ( .A0(n5326), .A1(n4041), .Z(n4362));
Q_AN02 U1746 ( .A0(n5326), .A1(n4040), .Z(n4361));
Q_AN02 U1747 ( .A0(n5326), .A1(n4039), .Z(n4360));
Q_AN02 U1748 ( .A0(n5326), .A1(n4038), .Z(n4359));
Q_AN02 U1749 ( .A0(n5326), .A1(n4037), .Z(n4358));
Q_AN02 U1750 ( .A0(n5326), .A1(n4036), .Z(n4357));
Q_AN02 U1751 ( .A0(n5326), .A1(n4035), .Z(n4356));
Q_AN02 U1752 ( .A0(n5326), .A1(n4034), .Z(n4355));
Q_AN02 U1753 ( .A0(n5326), .A1(n4033), .Z(n4354));
Q_AN02 U1754 ( .A0(n5326), .A1(n4032), .Z(n4353));
Q_AN02 U1755 ( .A0(n5326), .A1(n4031), .Z(n4352));
Q_AN02 U1756 ( .A0(n5326), .A1(n4030), .Z(n4351));
Q_AN02 U1757 ( .A0(n5326), .A1(n4029), .Z(n4350));
Q_AN02 U1758 ( .A0(n5326), .A1(n4028), .Z(n4349));
Q_AN02 U1759 ( .A0(n5326), .A1(n4027), .Z(n4348));
Q_AN02 U1760 ( .A0(n5326), .A1(n4026), .Z(n4347));
Q_AN02 U1761 ( .A0(n5326), .A1(n4025), .Z(n4346));
Q_AN02 U1762 ( .A0(n5326), .A1(n4024), .Z(n4345));
Q_AN02 U1763 ( .A0(n5326), .A1(n4023), .Z(n4344));
Q_AN02 U1764 ( .A0(n5326), .A1(n4022), .Z(n4343));
Q_AN02 U1765 ( .A0(n5326), .A1(n4021), .Z(n4342));
Q_AN02 U1766 ( .A0(n5326), .A1(n4020), .Z(n4341));
Q_AN02 U1767 ( .A0(n5326), .A1(n4019), .Z(n4340));
Q_AN02 U1768 ( .A0(n5326), .A1(n4018), .Z(n4339));
Q_AN02 U1769 ( .A0(n5326), .A1(n4017), .Z(n4338));
Q_AN02 U1770 ( .A0(n5326), .A1(n4016), .Z(n4337));
Q_AN02 U1771 ( .A0(n5326), .A1(n4015), .Z(n4336));
Q_AN02 U1772 ( .A0(n5326), .A1(n4014), .Z(n4335));
Q_AN02 U1773 ( .A0(n5326), .A1(n4013), .Z(n4334));
Q_AN02 U1774 ( .A0(n5326), .A1(n4012), .Z(n4333));
Q_AN02 U1775 ( .A0(n5326), .A1(n4011), .Z(n4332));
Q_AN02 U1776 ( .A0(n5326), .A1(n4010), .Z(n4331));
Q_AN02 U1777 ( .A0(n5326), .A1(n4009), .Z(n4330));
Q_AN02 U1778 ( .A0(n5326), .A1(n4008), .Z(n4329));
Q_AN02 U1779 ( .A0(n5326), .A1(n4007), .Z(n4328));
Q_AN02 U1780 ( .A0(n5326), .A1(n4006), .Z(n4327));
Q_AN02 U1781 ( .A0(n5326), .A1(n4005), .Z(n4326));
Q_AN02 U1782 ( .A0(n5326), .A1(n4004), .Z(n4325));
Q_AN02 U1783 ( .A0(n5326), .A1(n4003), .Z(n4324));
Q_AN02 U1784 ( .A0(n5326), .A1(n4002), .Z(n4323));
Q_AN02 U1785 ( .A0(n5326), .A1(n4001), .Z(n4322));
Q_AN02 U1786 ( .A0(n5326), .A1(n4000), .Z(n4321));
Q_AN02 U1787 ( .A0(n5326), .A1(n3999), .Z(n4320));
Q_AN02 U1788 ( .A0(n5326), .A1(n3998), .Z(n4319));
Q_AN02 U1789 ( .A0(n5326), .A1(n3997), .Z(n4318));
Q_AN02 U1790 ( .A0(n5326), .A1(n3996), .Z(n4317));
Q_AN02 U1791 ( .A0(n5326), .A1(n3995), .Z(n4316));
Q_AN02 U1792 ( .A0(n5326), .A1(n3994), .Z(n4315));
Q_AN02 U1793 ( .A0(n5326), .A1(n3993), .Z(n4314));
Q_AN02 U1794 ( .A0(n5326), .A1(n3992), .Z(n4313));
Q_AN02 U1795 ( .A0(n5326), .A1(n3991), .Z(n4312));
Q_AN02 U1796 ( .A0(n5326), .A1(n3990), .Z(n4311));
Q_AN02 U1797 ( .A0(n5326), .A1(n3989), .Z(n4310));
Q_AN02 U1798 ( .A0(n5326), .A1(n3988), .Z(n4309));
Q_AN02 U1799 ( .A0(n5326), .A1(n3987), .Z(n4308));
Q_AN02 U1800 ( .A0(n5326), .A1(n3986), .Z(n4307));
Q_AN02 U1801 ( .A0(n5326), .A1(n3985), .Z(n4306));
Q_AN02 U1802 ( .A0(n5326), .A1(n3984), .Z(n4305));
Q_AN02 U1803 ( .A0(n5326), .A1(n3983), .Z(n4304));
Q_AN02 U1804 ( .A0(n5326), .A1(n3982), .Z(n4303));
Q_AN02 U1805 ( .A0(n5326), .A1(n3981), .Z(n4302));
Q_AN02 U1806 ( .A0(n5326), .A1(n3980), .Z(n4301));
Q_AN02 U1807 ( .A0(n5326), .A1(n3979), .Z(n4300));
Q_AN02 U1808 ( .A0(n5326), .A1(n3978), .Z(n4299));
Q_AN02 U1809 ( .A0(n5326), .A1(n3977), .Z(n4298));
Q_AN02 U1810 ( .A0(n5326), .A1(n3976), .Z(n4297));
Q_AN02 U1811 ( .A0(n5326), .A1(n3975), .Z(n4296));
Q_AN02 U1812 ( .A0(n5326), .A1(n3974), .Z(n4295));
Q_AN02 U1813 ( .A0(n5326), .A1(n3973), .Z(n4294));
Q_AN02 U1814 ( .A0(n5326), .A1(n3972), .Z(n4293));
Q_AN02 U1815 ( .A0(n5326), .A1(n3971), .Z(n4292));
Q_AN02 U1816 ( .A0(n5326), .A1(n3970), .Z(n4291));
Q_AN02 U1817 ( .A0(n5326), .A1(n3969), .Z(n4290));
Q_MX04 U1818 ( .S0(n5331), .S1(n5326), .A0(_zyGfifo__gfdL365_0_P0_m2_cbid[19]), .A1(_zyGfifo__gfdL276_2_P0_m2_cbid[19]), .A2(_zyGfifo__gfdL268_4_P0_m2_cbid[19]), .A3(_zyGfifo__gfdL265_5_P0_m2_cbid[19]), .Z(n4289));
Q_MX04 U1819 ( .S0(n5331), .S1(n5326), .A0(_zyGfifo__gfdL365_0_P0_m2_cbid[18]), .A1(_zyGfifo__gfdL276_2_P0_m2_cbid[18]), .A2(_zyGfifo__gfdL268_4_P0_m2_cbid[18]), .A3(_zyGfifo__gfdL265_5_P0_m2_cbid[18]), .Z(n4288));
Q_MX04 U1820 ( .S0(n5331), .S1(n5326), .A0(_zyGfifo__gfdL365_0_P0_m2_cbid[17]), .A1(_zyGfifo__gfdL276_2_P0_m2_cbid[17]), .A2(_zyGfifo__gfdL268_4_P0_m2_cbid[17]), .A3(_zyGfifo__gfdL265_5_P0_m2_cbid[17]), .Z(n4287));
Q_MX04 U1821 ( .S0(n5331), .S1(n5326), .A0(_zyGfifo__gfdL365_0_P0_m2_cbid[16]), .A1(_zyGfifo__gfdL276_2_P0_m2_cbid[16]), .A2(_zyGfifo__gfdL268_4_P0_m2_cbid[16]), .A3(_zyGfifo__gfdL265_5_P0_m2_cbid[16]), .Z(n4286));
Q_MX04 U1822 ( .S0(n5331), .S1(n5326), .A0(_zyGfifo__gfdL365_0_P0_m2_cbid[15]), .A1(_zyGfifo__gfdL276_2_P0_m2_cbid[15]), .A2(_zyGfifo__gfdL268_4_P0_m2_cbid[15]), .A3(_zyGfifo__gfdL265_5_P0_m2_cbid[15]), .Z(n4285));
Q_MX04 U1823 ( .S0(n5331), .S1(n5326), .A0(_zyGfifo__gfdL365_0_P0_m2_cbid[14]), .A1(_zyGfifo__gfdL276_2_P0_m2_cbid[14]), .A2(_zyGfifo__gfdL268_4_P0_m2_cbid[14]), .A3(_zyGfifo__gfdL265_5_P0_m2_cbid[14]), .Z(n4284));
Q_MX04 U1824 ( .S0(n5331), .S1(n5326), .A0(_zyGfifo__gfdL365_0_P0_m2_cbid[13]), .A1(_zyGfifo__gfdL276_2_P0_m2_cbid[13]), .A2(_zyGfifo__gfdL268_4_P0_m2_cbid[13]), .A3(_zyGfifo__gfdL265_5_P0_m2_cbid[13]), .Z(n4283));
Q_MX04 U1825 ( .S0(n5331), .S1(n5326), .A0(_zyGfifo__gfdL365_0_P0_m2_cbid[12]), .A1(_zyGfifo__gfdL276_2_P0_m2_cbid[12]), .A2(_zyGfifo__gfdL268_4_P0_m2_cbid[12]), .A3(_zyGfifo__gfdL265_5_P0_m2_cbid[12]), .Z(n4282));
Q_MX04 U1826 ( .S0(n5331), .S1(n5326), .A0(_zyGfifo__gfdL365_0_P0_m2_cbid[11]), .A1(_zyGfifo__gfdL276_2_P0_m2_cbid[11]), .A2(_zyGfifo__gfdL268_4_P0_m2_cbid[11]), .A3(_zyGfifo__gfdL265_5_P0_m2_cbid[11]), .Z(n4281));
Q_MX04 U1827 ( .S0(n5331), .S1(n5326), .A0(_zyGfifo__gfdL365_0_P0_m2_cbid[10]), .A1(_zyGfifo__gfdL276_2_P0_m2_cbid[10]), .A2(_zyGfifo__gfdL268_4_P0_m2_cbid[10]), .A3(_zyGfifo__gfdL265_5_P0_m2_cbid[10]), .Z(n4280));
Q_MX04 U1828 ( .S0(n5331), .S1(n5326), .A0(_zyGfifo__gfdL365_0_P0_m2_cbid[9]), .A1(_zyGfifo__gfdL276_2_P0_m2_cbid[9]), .A2(_zyGfifo__gfdL268_4_P0_m2_cbid[9]), .A3(_zyGfifo__gfdL265_5_P0_m2_cbid[9]), .Z(n4279));
Q_MX04 U1829 ( .S0(n5331), .S1(n5326), .A0(_zyGfifo__gfdL365_0_P0_m2_cbid[8]), .A1(_zyGfifo__gfdL276_2_P0_m2_cbid[8]), .A2(_zyGfifo__gfdL268_4_P0_m2_cbid[8]), .A3(_zyGfifo__gfdL265_5_P0_m2_cbid[8]), .Z(n4278));
Q_MX04 U1830 ( .S0(n5331), .S1(n5326), .A0(_zyGfifo__gfdL365_0_P0_m2_cbid[7]), .A1(_zyGfifo__gfdL276_2_P0_m2_cbid[7]), .A2(_zyGfifo__gfdL268_4_P0_m2_cbid[7]), .A3(_zyGfifo__gfdL265_5_P0_m2_cbid[7]), .Z(n4277));
Q_MX04 U1831 ( .S0(n5331), .S1(n5326), .A0(_zyGfifo__gfdL365_0_P0_m2_cbid[6]), .A1(_zyGfifo__gfdL276_2_P0_m2_cbid[6]), .A2(_zyGfifo__gfdL268_4_P0_m2_cbid[6]), .A3(_zyGfifo__gfdL265_5_P0_m2_cbid[6]), .Z(n4276));
Q_MX04 U1832 ( .S0(n5331), .S1(n5326), .A0(_zyGfifo__gfdL365_0_P0_m2_cbid[5]), .A1(_zyGfifo__gfdL276_2_P0_m2_cbid[5]), .A2(_zyGfifo__gfdL268_4_P0_m2_cbid[5]), .A3(_zyGfifo__gfdL265_5_P0_m2_cbid[5]), .Z(n4275));
Q_MX04 U1833 ( .S0(n5331), .S1(n5326), .A0(_zyGfifo__gfdL365_0_P0_m2_cbid[4]), .A1(_zyGfifo__gfdL276_2_P0_m2_cbid[4]), .A2(_zyGfifo__gfdL268_4_P0_m2_cbid[4]), .A3(_zyGfifo__gfdL265_5_P0_m2_cbid[4]), .Z(n4274));
Q_MX04 U1834 ( .S0(n5331), .S1(n5326), .A0(_zyGfifo__gfdL365_0_P0_m2_cbid[3]), .A1(_zyGfifo__gfdL276_2_P0_m2_cbid[3]), .A2(_zyGfifo__gfdL268_4_P0_m2_cbid[3]), .A3(_zyGfifo__gfdL265_5_P0_m2_cbid[3]), .Z(n4273));
Q_MX04 U1835 ( .S0(n5331), .S1(n5326), .A0(_zyGfifo__gfdL365_0_P0_m2_cbid[2]), .A1(_zyGfifo__gfdL276_2_P0_m2_cbid[2]), .A2(_zyGfifo__gfdL268_4_P0_m2_cbid[2]), .A3(_zyGfifo__gfdL265_5_P0_m2_cbid[2]), .Z(n4272));
Q_MX04 U1836 ( .S0(n5331), .S1(n5326), .A0(_zyGfifo__gfdL365_0_P0_m2_cbid[1]), .A1(_zyGfifo__gfdL276_2_P0_m2_cbid[1]), .A2(_zyGfifo__gfdL268_4_P0_m2_cbid[1]), .A3(_zyGfifo__gfdL265_5_P0_m2_cbid[1]), .Z(n4271));
Q_MX04 U1837 ( .S0(n5331), .S1(n5326), .A0(_zyGfifo__gfdL365_0_P0_m2_cbid[0]), .A1(_zyGfifo__gfdL276_2_P0_m2_cbid[0]), .A2(_zyGfifo__gfdL268_4_P0_m2_cbid[0]), .A3(_zyGfifo__gfdL265_5_P0_m2_cbid[0]), .Z(n4270));
Q_MX02 U1838 ( .S(n5330), .A0(_zyGfifo__gfdL289_1_P0_m2_gfOff), .A1(_zyGfifo__gfdL271_3_P0_m2_gfOff), .Z(n3637));
Q_MX02 U1839 ( .S(n5330), .A0(_zyGfifo__gfdL289_1_P0_m2_cbid[19]), .A1(_zyGfifo__gfdL271_3_P0_m2_cbid[19]), .Z(n4268));
Q_MX02 U1840 ( .S(n5330), .A0(_zyGfifo__gfdL289_1_P0_m2_cbid[18]), .A1(_zyGfifo__gfdL271_3_P0_m2_cbid[18]), .Z(n4267));
Q_MX02 U1841 ( .S(n5330), .A0(_zyGfifo__gfdL289_1_P0_m2_cbid[17]), .A1(_zyGfifo__gfdL271_3_P0_m2_cbid[17]), .Z(n4266));
Q_MX02 U1842 ( .S(n5330), .A0(_zyGfifo__gfdL289_1_P0_m2_cbid[16]), .A1(_zyGfifo__gfdL271_3_P0_m2_cbid[16]), .Z(n4265));
Q_MX02 U1843 ( .S(n5330), .A0(_zyGfifo__gfdL289_1_P0_m2_cbid[15]), .A1(_zyGfifo__gfdL271_3_P0_m2_cbid[15]), .Z(n4264));
Q_MX02 U1844 ( .S(n5330), .A0(_zyGfifo__gfdL289_1_P0_m2_cbid[14]), .A1(_zyGfifo__gfdL271_3_P0_m2_cbid[14]), .Z(n4263));
Q_MX02 U1845 ( .S(n5330), .A0(_zyGfifo__gfdL289_1_P0_m2_cbid[13]), .A1(_zyGfifo__gfdL271_3_P0_m2_cbid[13]), .Z(n4262));
Q_MX02 U1846 ( .S(n5330), .A0(_zyGfifo__gfdL289_1_P0_m2_cbid[12]), .A1(_zyGfifo__gfdL271_3_P0_m2_cbid[12]), .Z(n4261));
Q_MX02 U1847 ( .S(n5330), .A0(_zyGfifo__gfdL289_1_P0_m2_cbid[11]), .A1(_zyGfifo__gfdL271_3_P0_m2_cbid[11]), .Z(n4260));
Q_MX02 U1848 ( .S(n5330), .A0(_zyGfifo__gfdL289_1_P0_m2_cbid[10]), .A1(_zyGfifo__gfdL271_3_P0_m2_cbid[10]), .Z(n4259));
Q_MX02 U1849 ( .S(n5330), .A0(_zyGfifo__gfdL289_1_P0_m2_cbid[9]), .A1(_zyGfifo__gfdL271_3_P0_m2_cbid[9]), .Z(n4258));
Q_MX02 U1850 ( .S(n5330), .A0(_zyGfifo__gfdL289_1_P0_m2_cbid[8]), .A1(_zyGfifo__gfdL271_3_P0_m2_cbid[8]), .Z(n4257));
Q_MX02 U1851 ( .S(n5330), .A0(_zyGfifo__gfdL289_1_P0_m2_cbid[7]), .A1(_zyGfifo__gfdL271_3_P0_m2_cbid[7]), .Z(n4256));
Q_MX02 U1852 ( .S(n5330), .A0(_zyGfifo__gfdL289_1_P0_m2_cbid[6]), .A1(_zyGfifo__gfdL271_3_P0_m2_cbid[6]), .Z(n4255));
Q_MX02 U1853 ( .S(n5330), .A0(_zyGfifo__gfdL289_1_P0_m2_cbid[5]), .A1(_zyGfifo__gfdL271_3_P0_m2_cbid[5]), .Z(n4254));
Q_MX02 U1854 ( .S(n5330), .A0(_zyGfifo__gfdL289_1_P0_m2_cbid[4]), .A1(_zyGfifo__gfdL271_3_P0_m2_cbid[4]), .Z(n4253));
Q_MX02 U1855 ( .S(n5330), .A0(_zyGfifo__gfdL289_1_P0_m2_cbid[3]), .A1(_zyGfifo__gfdL271_3_P0_m2_cbid[3]), .Z(n4252));
Q_MX02 U1856 ( .S(n5330), .A0(_zyGfifo__gfdL289_1_P0_m2_cbid[2]), .A1(_zyGfifo__gfdL271_3_P0_m2_cbid[2]), .Z(n4251));
Q_MX02 U1857 ( .S(n5330), .A0(_zyGfifo__gfdL289_1_P0_m2_cbid[1]), .A1(_zyGfifo__gfdL271_3_P0_m2_cbid[1]), .Z(n4250));
Q_MX02 U1858 ( .S(n5330), .A0(_zyGfifo__gfdL289_1_P0_m2_cbid[0]), .A1(_zyGfifo__gfdL271_3_P0_m2_cbid[0]), .Z(n4249));
Q_AN02 U1859 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[279]), .Z(n4248));
Q_AN02 U1860 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[278]), .Z(n4247));
Q_AN02 U1861 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[277]), .Z(n4246));
Q_AN02 U1862 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[276]), .Z(n4245));
Q_AN02 U1863 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[275]), .Z(n4244));
Q_AN02 U1864 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[274]), .Z(n4243));
Q_AN02 U1865 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[273]), .Z(n4242));
Q_AN02 U1866 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[272]), .Z(n4241));
Q_AN02 U1867 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[271]), .Z(n4240));
Q_AN02 U1868 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[270]), .Z(n4239));
Q_AN02 U1869 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[269]), .Z(n4238));
Q_AN02 U1870 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[268]), .Z(n4237));
Q_AN02 U1871 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[267]), .Z(n4236));
Q_AN02 U1872 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[266]), .Z(n4235));
Q_AN02 U1873 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[265]), .Z(n4234));
Q_AN02 U1874 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[264]), .Z(n4233));
Q_AN02 U1875 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[263]), .Z(n4232));
Q_AN02 U1876 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[262]), .Z(n4231));
Q_AN02 U1877 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[261]), .Z(n4230));
Q_AN02 U1878 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[260]), .Z(n4229));
Q_AN02 U1879 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[259]), .Z(n4228));
Q_AN02 U1880 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[258]), .Z(n4227));
Q_AN02 U1881 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[257]), .Z(n4226));
Q_AN02 U1882 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[256]), .Z(n4225));
Q_AN02 U1883 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[255]), .Z(n4224));
Q_AN02 U1884 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[254]), .Z(n4223));
Q_AN02 U1885 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[253]), .Z(n4222));
Q_AN02 U1886 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[252]), .Z(n4221));
Q_AN02 U1887 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[251]), .Z(n4220));
Q_AN02 U1888 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[250]), .Z(n4219));
Q_AN02 U1889 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[249]), .Z(n4218));
Q_AN02 U1890 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[248]), .Z(n4217));
Q_AN02 U1891 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[247]), .Z(n4216));
Q_AN02 U1892 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[246]), .Z(n4215));
Q_AN02 U1893 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[245]), .Z(n4214));
Q_AN02 U1894 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[244]), .Z(n4213));
Q_AN02 U1895 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[243]), .Z(n4212));
Q_AN02 U1896 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[242]), .Z(n4211));
Q_AN02 U1897 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[241]), .Z(n4210));
Q_AN02 U1898 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[240]), .Z(n4209));
Q_AN02 U1899 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[239]), .Z(n4208));
Q_AN02 U1900 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[238]), .Z(n4207));
Q_AN02 U1901 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[237]), .Z(n4206));
Q_AN02 U1902 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[236]), .Z(n4205));
Q_AN02 U1903 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[235]), .Z(n4204));
Q_AN02 U1904 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[234]), .Z(n4203));
Q_AN02 U1905 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[233]), .Z(n4202));
Q_AN02 U1906 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[232]), .Z(n4201));
Q_AN02 U1907 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[231]), .Z(n4200));
Q_AN02 U1908 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[230]), .Z(n4199));
Q_AN02 U1909 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[229]), .Z(n4198));
Q_AN02 U1910 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[228]), .Z(n4197));
Q_AN02 U1911 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[227]), .Z(n4196));
Q_AN02 U1912 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[226]), .Z(n4195));
Q_AN02 U1913 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[225]), .Z(n4194));
Q_AN02 U1914 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[224]), .Z(n4193));
Q_AN02 U1915 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[223]), .Z(n4192));
Q_AN02 U1916 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[222]), .Z(n4191));
Q_AN02 U1917 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[221]), .Z(n4190));
Q_AN02 U1918 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[220]), .Z(n4189));
Q_AN02 U1919 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[219]), .Z(n4188));
Q_AN02 U1920 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[218]), .Z(n4187));
Q_AN02 U1921 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[217]), .Z(n4186));
Q_AN02 U1922 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[216]), .Z(n4185));
Q_AN02 U1923 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[215]), .Z(n4184));
Q_AN02 U1924 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[214]), .Z(n4183));
Q_AN02 U1925 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[213]), .Z(n4182));
Q_AN02 U1926 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[212]), .Z(n4181));
Q_AN02 U1927 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[211]), .Z(n4180));
Q_AN02 U1928 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[210]), .Z(n4179));
Q_AN02 U1929 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[209]), .Z(n4178));
Q_AN02 U1930 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[208]), .Z(n4177));
Q_AN02 U1931 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[207]), .Z(n4176));
Q_AN02 U1932 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[206]), .Z(n4175));
Q_AN02 U1933 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[205]), .Z(n4174));
Q_AN02 U1934 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[204]), .Z(n4173));
Q_AN02 U1935 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[203]), .Z(n4172));
Q_AN02 U1936 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[202]), .Z(n4171));
Q_AN02 U1937 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[201]), .Z(n4170));
Q_AN02 U1938 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[200]), .Z(n4169));
Q_AN02 U1939 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[199]), .Z(n4168));
Q_AN02 U1940 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[198]), .Z(n4167));
Q_AN02 U1941 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[197]), .Z(n4166));
Q_AN02 U1942 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[196]), .Z(n4165));
Q_AN02 U1943 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[195]), .Z(n4164));
Q_AN02 U1944 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[194]), .Z(n4163));
Q_AN02 U1945 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[193]), .Z(n4162));
Q_AN02 U1946 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[192]), .Z(n4161));
Q_AN02 U1947 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[191]), .Z(n4160));
Q_AN02 U1948 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[190]), .Z(n4159));
Q_AN02 U1949 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[189]), .Z(n4158));
Q_AN02 U1950 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[188]), .Z(n4157));
Q_AN02 U1951 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[187]), .Z(n4156));
Q_AN02 U1952 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[186]), .Z(n4155));
Q_AN02 U1953 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[185]), .Z(n4154));
Q_AN02 U1954 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[184]), .Z(n4153));
Q_AN02 U1955 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[183]), .Z(n4152));
Q_AN02 U1956 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[182]), .Z(n4151));
Q_AN02 U1957 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[181]), .Z(n4150));
Q_AN02 U1958 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[180]), .Z(n4149));
Q_AN02 U1959 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[179]), .Z(n4148));
Q_AN02 U1960 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[178]), .Z(n4147));
Q_AN02 U1961 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[177]), .Z(n4146));
Q_AN02 U1962 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[176]), .Z(n4145));
Q_AN02 U1963 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[175]), .Z(n4144));
Q_AN02 U1964 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[174]), .Z(n4143));
Q_AN02 U1965 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[173]), .Z(n4142));
Q_AN02 U1966 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[172]), .Z(n4141));
Q_AN02 U1967 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[171]), .Z(n4140));
Q_AN02 U1968 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[170]), .Z(n4139));
Q_AN02 U1969 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[169]), .Z(n4138));
Q_AN02 U1970 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[168]), .Z(n4137));
Q_AN02 U1971 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[167]), .Z(n4136));
Q_AN02 U1972 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[166]), .Z(n4135));
Q_AN02 U1973 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[165]), .Z(n4134));
Q_AN02 U1974 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[164]), .Z(n4133));
Q_AN02 U1975 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[163]), .Z(n4132));
Q_AN02 U1976 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[162]), .Z(n4131));
Q_AN02 U1977 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[161]), .Z(n4130));
Q_AN02 U1978 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[160]), .Z(n4129));
Q_AN02 U1979 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[159]), .Z(n4128));
Q_AN02 U1980 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[158]), .Z(n4127));
Q_AN02 U1981 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[157]), .Z(n4126));
Q_AN02 U1982 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[156]), .Z(n4125));
Q_AN02 U1983 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[155]), .Z(n4124));
Q_AN02 U1984 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[154]), .Z(n4123));
Q_AN02 U1985 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[153]), .Z(n4122));
Q_AN02 U1986 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[152]), .Z(n4121));
Q_AN02 U1987 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[151]), .Z(n4120));
Q_AN02 U1988 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[150]), .Z(n4119));
Q_AN02 U1989 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[149]), .Z(n4118));
Q_AN02 U1990 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[148]), .Z(n4117));
Q_AN02 U1991 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[147]), .Z(n4116));
Q_AN02 U1992 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[146]), .Z(n4115));
Q_AN02 U1993 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[145]), .Z(n4114));
Q_AN02 U1994 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[144]), .Z(n4113));
Q_AN02 U1995 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[143]), .Z(n4112));
Q_AN02 U1996 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[142]), .Z(n4111));
Q_AN02 U1997 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[141]), .Z(n4110));
Q_AN02 U1998 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[140]), .Z(n4109));
Q_AN02 U1999 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[139]), .Z(n4108));
Q_AN02 U2000 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[138]), .Z(n4107));
Q_AN02 U2001 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[137]), .Z(n4106));
Q_AN02 U2002 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[136]), .Z(n4105));
Q_AN02 U2003 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[135]), .Z(n4104));
Q_AN02 U2004 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[134]), .Z(n4103));
Q_AN02 U2005 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[133]), .Z(n4102));
Q_AN02 U2006 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[132]), .Z(n4101));
Q_AN02 U2007 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[131]), .Z(n4100));
Q_AN02 U2008 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[130]), .Z(n4099));
Q_AN02 U2009 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[129]), .Z(n4098));
Q_AN02 U2010 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[128]), .Z(n4097));
Q_AN02 U2011 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[127]), .Z(n4096));
Q_AN02 U2012 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[126]), .Z(n4095));
Q_AN02 U2013 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[125]), .Z(n4094));
Q_AN02 U2014 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[124]), .Z(n4093));
Q_AN02 U2015 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[123]), .Z(n4092));
Q_AN02 U2016 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[122]), .Z(n4091));
Q_AN02 U2017 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[121]), .Z(n4090));
Q_AN02 U2018 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[120]), .Z(n4089));
Q_AN02 U2019 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[119]), .Z(n4088));
Q_AN02 U2020 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[118]), .Z(n4087));
Q_AN02 U2021 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[117]), .Z(n4086));
Q_AN02 U2022 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[116]), .Z(n4085));
Q_AN02 U2023 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[115]), .Z(n4084));
Q_AN02 U2024 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[114]), .Z(n4083));
Q_AN02 U2025 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[113]), .Z(n4082));
Q_AN02 U2026 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[112]), .Z(n4081));
Q_AN02 U2027 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[111]), .Z(n4080));
Q_AN02 U2028 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[110]), .Z(n4079));
Q_AN02 U2029 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[109]), .Z(n4078));
Q_AN02 U2030 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[108]), .Z(n4077));
Q_AN02 U2031 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[107]), .Z(n4076));
Q_AN02 U2032 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[106]), .Z(n4075));
Q_AN02 U2033 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[105]), .Z(n4074));
Q_AN02 U2034 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[104]), .Z(n4073));
Q_AN02 U2035 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[103]), .Z(n4072));
Q_AN02 U2036 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[102]), .Z(n4071));
Q_AN02 U2037 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[101]), .Z(n4070));
Q_AN02 U2038 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[100]), .Z(n4069));
Q_AN02 U2039 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[99]), .Z(n4068));
Q_AN02 U2040 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[98]), .Z(n4067));
Q_AN02 U2041 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[97]), .Z(n4066));
Q_AN02 U2042 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[96]), .Z(n4065));
Q_AN02 U2043 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[95]), .Z(n4064));
Q_AN02 U2044 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[94]), .Z(n4063));
Q_AN02 U2045 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[93]), .Z(n4062));
Q_AN02 U2046 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[92]), .Z(n4061));
Q_AN02 U2047 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[91]), .Z(n4060));
Q_AN02 U2048 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[90]), .Z(n4059));
Q_AN02 U2049 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[89]), .Z(n4058));
Q_AN02 U2050 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[88]), .Z(n4057));
Q_AN02 U2051 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[87]), .Z(n4056));
Q_AN02 U2052 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[86]), .Z(n4055));
Q_AN02 U2053 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[85]), .Z(n4054));
Q_AN02 U2054 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[84]), .Z(n4053));
Q_AN02 U2055 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[83]), .Z(n4052));
Q_AN02 U2056 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[82]), .Z(n4051));
Q_AN02 U2057 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[81]), .Z(n4050));
Q_AN02 U2058 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[80]), .Z(n4049));
Q_AN02 U2059 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[79]), .Z(n4048));
Q_AN02 U2060 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[78]), .Z(n4047));
Q_AN02 U2061 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[77]), .Z(n4046));
Q_AN02 U2062 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[76]), .Z(n4045));
Q_AN02 U2063 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[75]), .Z(n4044));
Q_AN02 U2064 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[74]), .Z(n4043));
Q_AN02 U2065 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[73]), .Z(n4042));
Q_AN02 U2066 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[72]), .Z(n4041));
Q_AN02 U2067 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[71]), .Z(n4040));
Q_AN02 U2068 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[70]), .Z(n4039));
Q_AN02 U2069 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[69]), .Z(n4038));
Q_AN02 U2070 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[68]), .Z(n4037));
Q_AN02 U2071 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[67]), .Z(n4036));
Q_AN02 U2072 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[66]), .Z(n4035));
Q_AN02 U2073 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[65]), .Z(n4034));
Q_AN02 U2074 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[64]), .Z(n4033));
Q_AN02 U2075 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[63]), .Z(n4032));
Q_AN02 U2076 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[62]), .Z(n4031));
Q_AN02 U2077 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[61]), .Z(n4030));
Q_AN02 U2078 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[60]), .Z(n4029));
Q_AN02 U2079 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[59]), .Z(n4028));
Q_AN02 U2080 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[58]), .Z(n4027));
Q_AN02 U2081 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[57]), .Z(n4026));
Q_AN02 U2082 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[56]), .Z(n4025));
Q_AN02 U2083 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[55]), .Z(n4024));
Q_AN02 U2084 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[54]), .Z(n4023));
Q_AN02 U2085 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[53]), .Z(n4022));
Q_AN02 U2086 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[52]), .Z(n4021));
Q_AN02 U2087 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[51]), .Z(n4020));
Q_AN02 U2088 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[50]), .Z(n4019));
Q_AN02 U2089 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[49]), .Z(n4018));
Q_AN02 U2090 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[48]), .Z(n4017));
Q_AN02 U2091 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[47]), .Z(n4016));
Q_AN02 U2092 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[46]), .Z(n4015));
Q_AN02 U2093 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[45]), .Z(n4014));
Q_AN02 U2094 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[44]), .Z(n4013));
Q_AN02 U2095 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[43]), .Z(n4012));
Q_AN02 U2096 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[42]), .Z(n4011));
Q_AN02 U2097 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[41]), .Z(n4010));
Q_AN02 U2098 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[40]), .Z(n4009));
Q_AN02 U2099 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[39]), .Z(n4008));
Q_AN02 U2100 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[38]), .Z(n4007));
Q_AN02 U2101 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[37]), .Z(n4006));
Q_AN02 U2102 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[36]), .Z(n4005));
Q_AN02 U2103 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[35]), .Z(n4004));
Q_AN02 U2104 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[34]), .Z(n4003));
Q_AN02 U2105 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[33]), .Z(n4002));
Q_AN02 U2106 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[32]), .Z(n4001));
Q_AN02 U2107 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[31]), .Z(n4000));
Q_AN02 U2108 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[30]), .Z(n3999));
Q_AN02 U2109 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[29]), .Z(n3998));
Q_AN02 U2110 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[28]), .Z(n3997));
Q_AN02 U2111 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[27]), .Z(n3996));
Q_AN02 U2112 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[26]), .Z(n3995));
Q_AN02 U2113 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[25]), .Z(n3994));
Q_AN02 U2114 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[24]), .Z(n3993));
Q_AN02 U2115 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[23]), .Z(n3992));
Q_AN02 U2116 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[22]), .Z(n3991));
Q_AN02 U2117 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[21]), .Z(n3990));
Q_AN02 U2118 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[20]), .Z(n3989));
Q_AN02 U2119 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[19]), .Z(n3988));
Q_AN02 U2120 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[18]), .Z(n3987));
Q_AN02 U2121 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[17]), .Z(n3986));
Q_AN02 U2122 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[16]), .Z(n3985));
Q_AN02 U2123 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[15]), .Z(n3984));
Q_AN02 U2124 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[14]), .Z(n3983));
Q_AN02 U2125 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[13]), .Z(n3982));
Q_AN02 U2126 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[12]), .Z(n3981));
Q_AN02 U2127 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[11]), .Z(n3980));
Q_AN02 U2128 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[10]), .Z(n3979));
Q_AN02 U2129 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[9]), .Z(n3978));
Q_AN02 U2130 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[8]), .Z(n3977));
Q_AN02 U2131 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[7]), .Z(n3976));
Q_AN02 U2132 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[6]), .Z(n3975));
Q_OR02 U2133 ( .A0(n3968), .A1(_zyictd_sysfunc_36_L258_0[5]), .Z(n3974));
Q_OR02 U2134 ( .A0(n3968), .A1(_zyictd_sysfunc_36_L258_0[4]), .Z(n3973));
Q_AN02 U2135 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[3]), .Z(n3972));
Q_AN02 U2136 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[2]), .Z(n3971));
Q_AN02 U2137 ( .A0(n5319), .A1(_zyictd_sysfunc_36_L258_0[1]), .Z(n3970));
Q_OR02 U2138 ( .A0(n3968), .A1(_zyictd_sysfunc_36_L258_0[0]), .Z(n3969));
Q_INV U2139 ( .A(n5319), .Z(n3968));
Q_OR03 U2140 ( .A0(n3967), .A1(n3966), .A2(n3965), .Z(n5337));
Q_OR03 U2141 ( .A0(n3949), .A1(n3951), .A2(n3964), .Z(n3965));
Q_OR03 U2142 ( .A0(n3963), .A1(n3962), .A2(n3961), .Z(n3966));
Q_OR02 U2143 ( .A0(n3891), .A1(n3889), .Z(n3963));
Q_OR02 U2144 ( .A0(n3887), .A1(n3886), .Z(n3962));
Q_OR03 U2145 ( .A0(n3899), .A1(n3897), .A2(n3960), .Z(n3961));
Q_OR02 U2146 ( .A0(n3895), .A1(n3893), .Z(n3960));
Q_OR03 U2147 ( .A0(n3959), .A1(n3958), .A2(n3957), .Z(n3967));
Q_OR02 U2148 ( .A0(n3907), .A1(n3905), .Z(n3959));
Q_OR02 U2149 ( .A0(n3903), .A1(n3901), .Z(n3958));
Q_OR03 U2150 ( .A0(n3915), .A1(n3913), .A2(n3956), .Z(n3957));
Q_OR02 U2151 ( .A0(n3911), .A1(n3909), .Z(n3956));
Q_OR03 U2152 ( .A0(n3955), .A1(n3954), .A2(n3953), .Z(n3964));
Q_OR02 U2153 ( .A0(n3923), .A1(n3921), .Z(n3955));
Q_OR02 U2154 ( .A0(n3919), .A1(n3917), .Z(n3954));
Q_OR03 U2155 ( .A0(n3931), .A1(n3929), .A2(n3952), .Z(n3953));
Q_OR02 U2156 ( .A0(n3927), .A1(n3925), .Z(n3952));
Q_OR03 U2157 ( .A0(n3939), .A1(n3937), .A2(n3950), .Z(n3951));
Q_OR02 U2158 ( .A0(n3935), .A1(n3933), .Z(n3950));
Q_OR03 U2159 ( .A0(n3947), .A1(n3945), .A2(n3948), .Z(n3949));
Q_OR02 U2160 ( .A0(n3943), .A1(n3941), .Z(n3948));
Q_XNR2 U2161 ( .A0(_zyM2L273_pbcT0[31]), .A1(n3946), .Z(n3947));
Q_OR02 U2162 ( .A0(_zyM2L273_pbcT0[30]), .A1(n3944), .Z(n3946));
Q_XNR2 U2163 ( .A0(_zyM2L273_pbcT0[30]), .A1(n3944), .Z(n3945));
Q_OR02 U2164 ( .A0(_zyM2L273_pbcT0[29]), .A1(n3942), .Z(n3944));
Q_XNR2 U2165 ( .A0(_zyM2L273_pbcT0[29]), .A1(n3942), .Z(n3943));
Q_OR02 U2166 ( .A0(_zyM2L273_pbcT0[28]), .A1(n3940), .Z(n3942));
Q_XNR2 U2167 ( .A0(_zyM2L273_pbcT0[28]), .A1(n3940), .Z(n3941));
Q_OR02 U2168 ( .A0(_zyM2L273_pbcT0[27]), .A1(n3938), .Z(n3940));
Q_XNR2 U2169 ( .A0(_zyM2L273_pbcT0[27]), .A1(n3938), .Z(n3939));
Q_OR02 U2170 ( .A0(_zyM2L273_pbcT0[26]), .A1(n3936), .Z(n3938));
Q_XNR2 U2171 ( .A0(_zyM2L273_pbcT0[26]), .A1(n3936), .Z(n3937));
Q_OR02 U2172 ( .A0(_zyM2L273_pbcT0[25]), .A1(n3934), .Z(n3936));
Q_XNR2 U2173 ( .A0(_zyM2L273_pbcT0[25]), .A1(n3934), .Z(n3935));
Q_OR02 U2174 ( .A0(_zyM2L273_pbcT0[24]), .A1(n3932), .Z(n3934));
Q_XNR2 U2175 ( .A0(_zyM2L273_pbcT0[24]), .A1(n3932), .Z(n3933));
Q_OR02 U2176 ( .A0(_zyM2L273_pbcT0[23]), .A1(n3930), .Z(n3932));
Q_XNR2 U2177 ( .A0(_zyM2L273_pbcT0[23]), .A1(n3930), .Z(n3931));
Q_OR02 U2178 ( .A0(_zyM2L273_pbcT0[22]), .A1(n3928), .Z(n3930));
Q_XNR2 U2179 ( .A0(_zyM2L273_pbcT0[22]), .A1(n3928), .Z(n3929));
Q_OR02 U2180 ( .A0(_zyM2L273_pbcT0[21]), .A1(n3926), .Z(n3928));
Q_XNR2 U2181 ( .A0(_zyM2L273_pbcT0[21]), .A1(n3926), .Z(n3927));
Q_OR02 U2182 ( .A0(_zyM2L273_pbcT0[20]), .A1(n3924), .Z(n3926));
Q_XNR2 U2183 ( .A0(_zyM2L273_pbcT0[20]), .A1(n3924), .Z(n3925));
Q_OR02 U2184 ( .A0(_zyM2L273_pbcT0[19]), .A1(n3922), .Z(n3924));
Q_XNR2 U2185 ( .A0(_zyM2L273_pbcT0[19]), .A1(n3922), .Z(n3923));
Q_OR02 U2186 ( .A0(_zyM2L273_pbcT0[18]), .A1(n3920), .Z(n3922));
Q_XNR2 U2187 ( .A0(_zyM2L273_pbcT0[18]), .A1(n3920), .Z(n3921));
Q_OR02 U2188 ( .A0(_zyM2L273_pbcT0[17]), .A1(n3918), .Z(n3920));
Q_XNR2 U2189 ( .A0(_zyM2L273_pbcT0[17]), .A1(n3918), .Z(n3919));
Q_OR02 U2190 ( .A0(_zyM2L273_pbcT0[16]), .A1(n3916), .Z(n3918));
Q_XNR2 U2191 ( .A0(_zyM2L273_pbcT0[16]), .A1(n3916), .Z(n3917));
Q_OR02 U2192 ( .A0(_zyM2L273_pbcT0[15]), .A1(n3914), .Z(n3916));
Q_XNR2 U2193 ( .A0(_zyM2L273_pbcT0[15]), .A1(n3914), .Z(n3915));
Q_OR02 U2194 ( .A0(_zyM2L273_pbcT0[14]), .A1(n3912), .Z(n3914));
Q_XNR2 U2195 ( .A0(_zyM2L273_pbcT0[14]), .A1(n3912), .Z(n3913));
Q_OR02 U2196 ( .A0(_zyM2L273_pbcT0[13]), .A1(n3910), .Z(n3912));
Q_XNR2 U2197 ( .A0(_zyM2L273_pbcT0[13]), .A1(n3910), .Z(n3911));
Q_OR02 U2198 ( .A0(_zyM2L273_pbcT0[12]), .A1(n3908), .Z(n3910));
Q_XNR2 U2199 ( .A0(_zyM2L273_pbcT0[12]), .A1(n3908), .Z(n3909));
Q_OR02 U2200 ( .A0(_zyM2L273_pbcT0[11]), .A1(n3906), .Z(n3908));
Q_XNR2 U2201 ( .A0(_zyM2L273_pbcT0[11]), .A1(n3906), .Z(n3907));
Q_OR02 U2202 ( .A0(_zyM2L273_pbcT0[10]), .A1(n3904), .Z(n3906));
Q_XNR2 U2203 ( .A0(_zyM2L273_pbcT0[10]), .A1(n3904), .Z(n3905));
Q_OR02 U2204 ( .A0(_zyM2L273_pbcT0[9]), .A1(n3902), .Z(n3904));
Q_XNR2 U2205 ( .A0(_zyM2L273_pbcT0[9]), .A1(n3902), .Z(n3903));
Q_OR02 U2206 ( .A0(_zyM2L273_pbcT0[8]), .A1(n3900), .Z(n3902));
Q_XNR2 U2207 ( .A0(_zyM2L273_pbcT0[8]), .A1(n3900), .Z(n3901));
Q_OR02 U2208 ( .A0(_zyM2L273_pbcT0[7]), .A1(n3898), .Z(n3900));
Q_XNR2 U2209 ( .A0(_zyM2L273_pbcT0[7]), .A1(n3898), .Z(n3899));
Q_OR02 U2210 ( .A0(_zyM2L273_pbcT0[6]), .A1(n3896), .Z(n3898));
Q_XNR2 U2211 ( .A0(_zyM2L273_pbcT0[6]), .A1(n3896), .Z(n3897));
Q_OR02 U2212 ( .A0(_zyM2L273_pbcT0[5]), .A1(n3894), .Z(n3896));
Q_XNR2 U2213 ( .A0(_zyM2L273_pbcT0[5]), .A1(n3894), .Z(n3895));
Q_OR02 U2214 ( .A0(_zyM2L273_pbcT0[4]), .A1(n3892), .Z(n3894));
Q_XNR2 U2215 ( .A0(_zyM2L273_pbcT0[4]), .A1(n3892), .Z(n3893));
Q_OR02 U2216 ( .A0(_zyM2L273_pbcT0[3]), .A1(n3890), .Z(n3892));
Q_XNR2 U2217 ( .A0(_zyM2L273_pbcT0[3]), .A1(n3890), .Z(n3891));
Q_OR02 U2218 ( .A0(_zyM2L273_pbcT0[2]), .A1(n3888), .Z(n3890));
Q_XNR2 U2219 ( .A0(_zyM2L273_pbcT0[2]), .A1(n3888), .Z(n3889));
Q_OR02 U2220 ( .A0(_zyM2L273_pbcT0[1]), .A1(_zyM2L273_pbcT0[0]), .Z(n3888));
Q_XNR2 U2221 ( .A0(_zyM2L273_pbcT0[1]), .A1(_zyM2L273_pbcT0[0]), .Z(n3887));
Q_OR03 U2222 ( .A0(n3885), .A1(n3884), .A2(n3883), .Z(n5338));
Q_OR03 U2223 ( .A0(n3867), .A1(n3869), .A2(n3882), .Z(n3883));
Q_OR03 U2224 ( .A0(n3881), .A1(n3880), .A2(n3879), .Z(n3884));
Q_OR02 U2225 ( .A0(n3809), .A1(n3807), .Z(n3881));
Q_OR02 U2226 ( .A0(n3805), .A1(n3804), .Z(n3880));
Q_OR03 U2227 ( .A0(n3817), .A1(n3815), .A2(n3878), .Z(n3879));
Q_OR02 U2228 ( .A0(n3813), .A1(n3811), .Z(n3878));
Q_OR03 U2229 ( .A0(n3877), .A1(n3876), .A2(n3875), .Z(n3885));
Q_OR02 U2230 ( .A0(n3825), .A1(n3823), .Z(n3877));
Q_OR02 U2231 ( .A0(n3821), .A1(n3819), .Z(n3876));
Q_OR03 U2232 ( .A0(n3833), .A1(n3831), .A2(n3874), .Z(n3875));
Q_OR02 U2233 ( .A0(n3829), .A1(n3827), .Z(n3874));
Q_OR03 U2234 ( .A0(n3873), .A1(n3872), .A2(n3871), .Z(n3882));
Q_OR02 U2235 ( .A0(n3841), .A1(n3839), .Z(n3873));
Q_OR02 U2236 ( .A0(n3837), .A1(n3835), .Z(n3872));
Q_OR03 U2237 ( .A0(n3849), .A1(n3847), .A2(n3870), .Z(n3871));
Q_OR02 U2238 ( .A0(n3845), .A1(n3843), .Z(n3870));
Q_OR03 U2239 ( .A0(n3857), .A1(n3855), .A2(n3868), .Z(n3869));
Q_OR02 U2240 ( .A0(n3853), .A1(n3851), .Z(n3868));
Q_OR03 U2241 ( .A0(n3865), .A1(n3863), .A2(n3866), .Z(n3867));
Q_OR02 U2242 ( .A0(n3861), .A1(n3859), .Z(n3866));
Q_XNR2 U2243 ( .A0(_zyM2L286_pbcT1[31]), .A1(n3864), .Z(n3865));
Q_OR02 U2244 ( .A0(_zyM2L286_pbcT1[30]), .A1(n3862), .Z(n3864));
Q_XNR2 U2245 ( .A0(_zyM2L286_pbcT1[30]), .A1(n3862), .Z(n3863));
Q_OR02 U2246 ( .A0(_zyM2L286_pbcT1[29]), .A1(n3860), .Z(n3862));
Q_XNR2 U2247 ( .A0(_zyM2L286_pbcT1[29]), .A1(n3860), .Z(n3861));
Q_OR02 U2248 ( .A0(_zyM2L286_pbcT1[28]), .A1(n3858), .Z(n3860));
Q_XNR2 U2249 ( .A0(_zyM2L286_pbcT1[28]), .A1(n3858), .Z(n3859));
Q_OR02 U2250 ( .A0(_zyM2L286_pbcT1[27]), .A1(n3856), .Z(n3858));
Q_XNR2 U2251 ( .A0(_zyM2L286_pbcT1[27]), .A1(n3856), .Z(n3857));
Q_OR02 U2252 ( .A0(_zyM2L286_pbcT1[26]), .A1(n3854), .Z(n3856));
Q_XNR2 U2253 ( .A0(_zyM2L286_pbcT1[26]), .A1(n3854), .Z(n3855));
Q_OR02 U2254 ( .A0(_zyM2L286_pbcT1[25]), .A1(n3852), .Z(n3854));
Q_XNR2 U2255 ( .A0(_zyM2L286_pbcT1[25]), .A1(n3852), .Z(n3853));
Q_OR02 U2256 ( .A0(_zyM2L286_pbcT1[24]), .A1(n3850), .Z(n3852));
Q_XNR2 U2257 ( .A0(_zyM2L286_pbcT1[24]), .A1(n3850), .Z(n3851));
Q_OR02 U2258 ( .A0(_zyM2L286_pbcT1[23]), .A1(n3848), .Z(n3850));
Q_XNR2 U2259 ( .A0(_zyM2L286_pbcT1[23]), .A1(n3848), .Z(n3849));
Q_OR02 U2260 ( .A0(_zyM2L286_pbcT1[22]), .A1(n3846), .Z(n3848));
Q_XNR2 U2261 ( .A0(_zyM2L286_pbcT1[22]), .A1(n3846), .Z(n3847));
Q_OR02 U2262 ( .A0(_zyM2L286_pbcT1[21]), .A1(n3844), .Z(n3846));
Q_XNR2 U2263 ( .A0(_zyM2L286_pbcT1[21]), .A1(n3844), .Z(n3845));
Q_OR02 U2264 ( .A0(_zyM2L286_pbcT1[20]), .A1(n3842), .Z(n3844));
Q_XNR2 U2265 ( .A0(_zyM2L286_pbcT1[20]), .A1(n3842), .Z(n3843));
Q_OR02 U2266 ( .A0(_zyM2L286_pbcT1[19]), .A1(n3840), .Z(n3842));
Q_XNR2 U2267 ( .A0(_zyM2L286_pbcT1[19]), .A1(n3840), .Z(n3841));
Q_OR02 U2268 ( .A0(_zyM2L286_pbcT1[18]), .A1(n3838), .Z(n3840));
Q_XNR2 U2269 ( .A0(_zyM2L286_pbcT1[18]), .A1(n3838), .Z(n3839));
Q_OR02 U2270 ( .A0(_zyM2L286_pbcT1[17]), .A1(n3836), .Z(n3838));
Q_XNR2 U2271 ( .A0(_zyM2L286_pbcT1[17]), .A1(n3836), .Z(n3837));
Q_OR02 U2272 ( .A0(_zyM2L286_pbcT1[16]), .A1(n3834), .Z(n3836));
Q_XNR2 U2273 ( .A0(_zyM2L286_pbcT1[16]), .A1(n3834), .Z(n3835));
Q_OR02 U2274 ( .A0(_zyM2L286_pbcT1[15]), .A1(n3832), .Z(n3834));
Q_XNR2 U2275 ( .A0(_zyM2L286_pbcT1[15]), .A1(n3832), .Z(n3833));
Q_OR02 U2276 ( .A0(_zyM2L286_pbcT1[14]), .A1(n3830), .Z(n3832));
Q_XNR2 U2277 ( .A0(_zyM2L286_pbcT1[14]), .A1(n3830), .Z(n3831));
Q_OR02 U2278 ( .A0(_zyM2L286_pbcT1[13]), .A1(n3828), .Z(n3830));
Q_XNR2 U2279 ( .A0(_zyM2L286_pbcT1[13]), .A1(n3828), .Z(n3829));
Q_OR02 U2280 ( .A0(_zyM2L286_pbcT1[12]), .A1(n3826), .Z(n3828));
Q_XNR2 U2281 ( .A0(_zyM2L286_pbcT1[12]), .A1(n3826), .Z(n3827));
Q_OR02 U2282 ( .A0(_zyM2L286_pbcT1[11]), .A1(n3824), .Z(n3826));
Q_XNR2 U2283 ( .A0(_zyM2L286_pbcT1[11]), .A1(n3824), .Z(n3825));
Q_OR02 U2284 ( .A0(_zyM2L286_pbcT1[10]), .A1(n3822), .Z(n3824));
Q_XNR2 U2285 ( .A0(_zyM2L286_pbcT1[10]), .A1(n3822), .Z(n3823));
Q_OR02 U2286 ( .A0(_zyM2L286_pbcT1[9]), .A1(n3820), .Z(n3822));
Q_XNR2 U2287 ( .A0(_zyM2L286_pbcT1[9]), .A1(n3820), .Z(n3821));
Q_OR02 U2288 ( .A0(_zyM2L286_pbcT1[8]), .A1(n3818), .Z(n3820));
Q_XNR2 U2289 ( .A0(_zyM2L286_pbcT1[8]), .A1(n3818), .Z(n3819));
Q_OR02 U2290 ( .A0(_zyM2L286_pbcT1[7]), .A1(n3816), .Z(n3818));
Q_XNR2 U2291 ( .A0(_zyM2L286_pbcT1[7]), .A1(n3816), .Z(n3817));
Q_OR02 U2292 ( .A0(_zyM2L286_pbcT1[6]), .A1(n3814), .Z(n3816));
Q_XNR2 U2293 ( .A0(_zyM2L286_pbcT1[6]), .A1(n3814), .Z(n3815));
Q_OR02 U2294 ( .A0(_zyM2L286_pbcT1[5]), .A1(n3812), .Z(n3814));
Q_XNR2 U2295 ( .A0(_zyM2L286_pbcT1[5]), .A1(n3812), .Z(n3813));
Q_OR02 U2296 ( .A0(_zyM2L286_pbcT1[4]), .A1(n3810), .Z(n3812));
Q_XNR2 U2297 ( .A0(_zyM2L286_pbcT1[4]), .A1(n3810), .Z(n3811));
Q_OR02 U2298 ( .A0(_zyM2L286_pbcT1[3]), .A1(n3808), .Z(n3810));
Q_XNR2 U2299 ( .A0(_zyM2L286_pbcT1[3]), .A1(n3808), .Z(n3809));
Q_OR02 U2300 ( .A0(_zyM2L286_pbcT1[2]), .A1(n3806), .Z(n3808));
Q_XNR2 U2301 ( .A0(_zyM2L286_pbcT1[2]), .A1(n3806), .Z(n3807));
Q_OR02 U2302 ( .A0(_zyM2L286_pbcT1[1]), .A1(_zyM2L286_pbcT1[0]), .Z(n3806));
Q_XNR2 U2303 ( .A0(_zyM2L286_pbcT1[1]), .A1(_zyM2L286_pbcT1[0]), .Z(n3805));
Q_OR03 U2304 ( .A0(n3803), .A1(n3802), .A2(n3801), .Z(n5339));
Q_OR03 U2305 ( .A0(n3785), .A1(n3787), .A2(n3800), .Z(n3801));
Q_OR03 U2306 ( .A0(n3799), .A1(n3798), .A2(n3797), .Z(n3802));
Q_OR02 U2307 ( .A0(n3727), .A1(n3725), .Z(n3799));
Q_OR02 U2308 ( .A0(n3723), .A1(n3722), .Z(n3798));
Q_OR03 U2309 ( .A0(n3735), .A1(n3733), .A2(n3796), .Z(n3797));
Q_OR02 U2310 ( .A0(n3731), .A1(n3729), .Z(n3796));
Q_OR03 U2311 ( .A0(n3795), .A1(n3794), .A2(n3793), .Z(n3803));
Q_OR02 U2312 ( .A0(n3743), .A1(n3741), .Z(n3795));
Q_OR02 U2313 ( .A0(n3739), .A1(n3737), .Z(n3794));
Q_OR03 U2314 ( .A0(n3751), .A1(n3749), .A2(n3792), .Z(n3793));
Q_OR02 U2315 ( .A0(n3747), .A1(n3745), .Z(n3792));
Q_OR03 U2316 ( .A0(n3791), .A1(n3790), .A2(n3789), .Z(n3800));
Q_OR02 U2317 ( .A0(n3759), .A1(n3757), .Z(n3791));
Q_OR02 U2318 ( .A0(n3755), .A1(n3753), .Z(n3790));
Q_OR03 U2319 ( .A0(n3767), .A1(n3765), .A2(n3788), .Z(n3789));
Q_OR02 U2320 ( .A0(n3763), .A1(n3761), .Z(n3788));
Q_OR03 U2321 ( .A0(n3775), .A1(n3773), .A2(n3786), .Z(n3787));
Q_OR02 U2322 ( .A0(n3771), .A1(n3769), .Z(n3786));
Q_OR03 U2323 ( .A0(n3783), .A1(n3781), .A2(n3784), .Z(n3785));
Q_OR02 U2324 ( .A0(n3779), .A1(n3777), .Z(n3784));
Q_XNR2 U2325 ( .A0(_zyM2L292_pbcT2[31]), .A1(n3782), .Z(n3783));
Q_OR02 U2326 ( .A0(_zyM2L292_pbcT2[30]), .A1(n3780), .Z(n3782));
Q_XNR2 U2327 ( .A0(_zyM2L292_pbcT2[30]), .A1(n3780), .Z(n3781));
Q_OR02 U2328 ( .A0(_zyM2L292_pbcT2[29]), .A1(n3778), .Z(n3780));
Q_XNR2 U2329 ( .A0(_zyM2L292_pbcT2[29]), .A1(n3778), .Z(n3779));
Q_OR02 U2330 ( .A0(_zyM2L292_pbcT2[28]), .A1(n3776), .Z(n3778));
Q_XNR2 U2331 ( .A0(_zyM2L292_pbcT2[28]), .A1(n3776), .Z(n3777));
Q_OR02 U2332 ( .A0(_zyM2L292_pbcT2[27]), .A1(n3774), .Z(n3776));
Q_XNR2 U2333 ( .A0(_zyM2L292_pbcT2[27]), .A1(n3774), .Z(n3775));
Q_OR02 U2334 ( .A0(_zyM2L292_pbcT2[26]), .A1(n3772), .Z(n3774));
Q_XNR2 U2335 ( .A0(_zyM2L292_pbcT2[26]), .A1(n3772), .Z(n3773));
Q_OR02 U2336 ( .A0(_zyM2L292_pbcT2[25]), .A1(n3770), .Z(n3772));
Q_XNR2 U2337 ( .A0(_zyM2L292_pbcT2[25]), .A1(n3770), .Z(n3771));
Q_OR02 U2338 ( .A0(_zyM2L292_pbcT2[24]), .A1(n3768), .Z(n3770));
Q_XNR2 U2339 ( .A0(_zyM2L292_pbcT2[24]), .A1(n3768), .Z(n3769));
Q_OR02 U2340 ( .A0(_zyM2L292_pbcT2[23]), .A1(n3766), .Z(n3768));
Q_XNR2 U2341 ( .A0(_zyM2L292_pbcT2[23]), .A1(n3766), .Z(n3767));
Q_OR02 U2342 ( .A0(_zyM2L292_pbcT2[22]), .A1(n3764), .Z(n3766));
Q_XNR2 U2343 ( .A0(_zyM2L292_pbcT2[22]), .A1(n3764), .Z(n3765));
Q_OR02 U2344 ( .A0(_zyM2L292_pbcT2[21]), .A1(n3762), .Z(n3764));
Q_XNR2 U2345 ( .A0(_zyM2L292_pbcT2[21]), .A1(n3762), .Z(n3763));
Q_OR02 U2346 ( .A0(_zyM2L292_pbcT2[20]), .A1(n3760), .Z(n3762));
Q_XNR2 U2347 ( .A0(_zyM2L292_pbcT2[20]), .A1(n3760), .Z(n3761));
Q_OR02 U2348 ( .A0(_zyM2L292_pbcT2[19]), .A1(n3758), .Z(n3760));
Q_XNR2 U2349 ( .A0(_zyM2L292_pbcT2[19]), .A1(n3758), .Z(n3759));
Q_OR02 U2350 ( .A0(_zyM2L292_pbcT2[18]), .A1(n3756), .Z(n3758));
Q_XNR2 U2351 ( .A0(_zyM2L292_pbcT2[18]), .A1(n3756), .Z(n3757));
Q_OR02 U2352 ( .A0(_zyM2L292_pbcT2[17]), .A1(n3754), .Z(n3756));
Q_XNR2 U2353 ( .A0(_zyM2L292_pbcT2[17]), .A1(n3754), .Z(n3755));
Q_OR02 U2354 ( .A0(_zyM2L292_pbcT2[16]), .A1(n3752), .Z(n3754));
Q_XNR2 U2355 ( .A0(_zyM2L292_pbcT2[16]), .A1(n3752), .Z(n3753));
Q_OR02 U2356 ( .A0(_zyM2L292_pbcT2[15]), .A1(n3750), .Z(n3752));
Q_XNR2 U2357 ( .A0(_zyM2L292_pbcT2[15]), .A1(n3750), .Z(n3751));
Q_OR02 U2358 ( .A0(_zyM2L292_pbcT2[14]), .A1(n3748), .Z(n3750));
Q_XNR2 U2359 ( .A0(_zyM2L292_pbcT2[14]), .A1(n3748), .Z(n3749));
Q_OR02 U2360 ( .A0(_zyM2L292_pbcT2[13]), .A1(n3746), .Z(n3748));
Q_XNR2 U2361 ( .A0(_zyM2L292_pbcT2[13]), .A1(n3746), .Z(n3747));
Q_OR02 U2362 ( .A0(_zyM2L292_pbcT2[12]), .A1(n3744), .Z(n3746));
Q_XNR2 U2363 ( .A0(_zyM2L292_pbcT2[12]), .A1(n3744), .Z(n3745));
Q_OR02 U2364 ( .A0(_zyM2L292_pbcT2[11]), .A1(n3742), .Z(n3744));
Q_XNR2 U2365 ( .A0(_zyM2L292_pbcT2[11]), .A1(n3742), .Z(n3743));
Q_OR02 U2366 ( .A0(_zyM2L292_pbcT2[10]), .A1(n3740), .Z(n3742));
Q_XNR2 U2367 ( .A0(_zyM2L292_pbcT2[10]), .A1(n3740), .Z(n3741));
Q_OR02 U2368 ( .A0(_zyM2L292_pbcT2[9]), .A1(n3738), .Z(n3740));
Q_XNR2 U2369 ( .A0(_zyM2L292_pbcT2[9]), .A1(n3738), .Z(n3739));
Q_OR02 U2370 ( .A0(_zyM2L292_pbcT2[8]), .A1(n3736), .Z(n3738));
Q_XNR2 U2371 ( .A0(_zyM2L292_pbcT2[8]), .A1(n3736), .Z(n3737));
Q_OR02 U2372 ( .A0(_zyM2L292_pbcT2[7]), .A1(n3734), .Z(n3736));
Q_XNR2 U2373 ( .A0(_zyM2L292_pbcT2[7]), .A1(n3734), .Z(n3735));
Q_OR02 U2374 ( .A0(_zyM2L292_pbcT2[6]), .A1(n3732), .Z(n3734));
Q_XNR2 U2375 ( .A0(_zyM2L292_pbcT2[6]), .A1(n3732), .Z(n3733));
Q_OR02 U2376 ( .A0(_zyM2L292_pbcT2[5]), .A1(n3730), .Z(n3732));
Q_XNR2 U2377 ( .A0(_zyM2L292_pbcT2[5]), .A1(n3730), .Z(n3731));
Q_OR02 U2378 ( .A0(_zyM2L292_pbcT2[4]), .A1(n3728), .Z(n3730));
Q_XNR2 U2379 ( .A0(_zyM2L292_pbcT2[4]), .A1(n3728), .Z(n3729));
Q_OR02 U2380 ( .A0(_zyM2L292_pbcT2[3]), .A1(n3726), .Z(n3728));
Q_XNR2 U2381 ( .A0(_zyM2L292_pbcT2[3]), .A1(n3726), .Z(n3727));
Q_OR02 U2382 ( .A0(_zyM2L292_pbcT2[2]), .A1(n3724), .Z(n3726));
Q_XNR2 U2383 ( .A0(_zyM2L292_pbcT2[2]), .A1(n3724), .Z(n3725));
Q_OR02 U2384 ( .A0(_zyM2L292_pbcT2[1]), .A1(_zyM2L292_pbcT2[0]), .Z(n3724));
Q_XNR2 U2385 ( .A0(_zyM2L292_pbcT2[1]), .A1(_zyM2L292_pbcT2[0]), .Z(n3723));
Q_OR03 U2386 ( .A0(n3711), .A1(n3713), .A2(n3720), .Z(n3721));
Q_OR03 U2387 ( .A0(n3703), .A1(n3705), .A2(n3718), .Z(n3719));
Q_OR03 U2388 ( .A0(n3717), .A1(n3716), .A2(n3715), .Z(n3720));
Q_OR02 U2389 ( .A0(n3645), .A1(n3643), .Z(n3717));
Q_OR02 U2390 ( .A0(n3641), .A1(n3640), .Z(n3716));
Q_OR03 U2391 ( .A0(n3653), .A1(n3651), .A2(n3714), .Z(n3715));
Q_OR02 U2392 ( .A0(n3649), .A1(n3647), .Z(n3714));
Q_OR03 U2393 ( .A0(n3661), .A1(n3659), .A2(n3712), .Z(n3713));
Q_OR02 U2394 ( .A0(n3657), .A1(n3655), .Z(n3712));
Q_OR03 U2395 ( .A0(n3669), .A1(n3667), .A2(n3710), .Z(n3711));
Q_OR02 U2396 ( .A0(n3665), .A1(n3663), .Z(n3710));
Q_OR03 U2397 ( .A0(n3709), .A1(n3708), .A2(n3707), .Z(n3718));
Q_OR02 U2398 ( .A0(n3677), .A1(n3675), .Z(n3709));
Q_OR02 U2399 ( .A0(n3673), .A1(n3671), .Z(n3708));
Q_OR03 U2400 ( .A0(n3685), .A1(n3683), .A2(n3706), .Z(n3707));
Q_OR02 U2401 ( .A0(n3681), .A1(n3679), .Z(n3706));
Q_OR03 U2402 ( .A0(n3693), .A1(n3691), .A2(n3704), .Z(n3705));
Q_OR02 U2403 ( .A0(n3689), .A1(n3687), .Z(n3704));
Q_OR03 U2404 ( .A0(n3701), .A1(n3699), .A2(n3702), .Z(n3703));
Q_OR02 U2405 ( .A0(n3697), .A1(n3695), .Z(n3702));
Q_XNR2 U2406 ( .A0(_zyM2L299_pbcT3[31]), .A1(n3700), .Z(n3701));
Q_OR02 U2407 ( .A0(_zyM2L299_pbcT3[30]), .A1(n3698), .Z(n3700));
Q_XNR2 U2408 ( .A0(_zyM2L299_pbcT3[30]), .A1(n3698), .Z(n3699));
Q_OR02 U2409 ( .A0(_zyM2L299_pbcT3[29]), .A1(n3696), .Z(n3698));
Q_XNR2 U2410 ( .A0(_zyM2L299_pbcT3[29]), .A1(n3696), .Z(n3697));
Q_OR02 U2411 ( .A0(_zyM2L299_pbcT3[28]), .A1(n3694), .Z(n3696));
Q_XNR2 U2412 ( .A0(_zyM2L299_pbcT3[28]), .A1(n3694), .Z(n3695));
Q_OR02 U2413 ( .A0(_zyM2L299_pbcT3[27]), .A1(n3692), .Z(n3694));
Q_XNR2 U2414 ( .A0(_zyM2L299_pbcT3[27]), .A1(n3692), .Z(n3693));
Q_OR02 U2415 ( .A0(_zyM2L299_pbcT3[26]), .A1(n3690), .Z(n3692));
Q_XNR2 U2416 ( .A0(_zyM2L299_pbcT3[26]), .A1(n3690), .Z(n3691));
Q_OR02 U2417 ( .A0(_zyM2L299_pbcT3[25]), .A1(n3688), .Z(n3690));
Q_XNR2 U2418 ( .A0(_zyM2L299_pbcT3[25]), .A1(n3688), .Z(n3689));
Q_OR02 U2419 ( .A0(_zyM2L299_pbcT3[24]), .A1(n3686), .Z(n3688));
Q_XNR2 U2420 ( .A0(_zyM2L299_pbcT3[24]), .A1(n3686), .Z(n3687));
Q_OR02 U2421 ( .A0(_zyM2L299_pbcT3[23]), .A1(n3684), .Z(n3686));
Q_XNR2 U2422 ( .A0(_zyM2L299_pbcT3[23]), .A1(n3684), .Z(n3685));
Q_OR02 U2423 ( .A0(_zyM2L299_pbcT3[22]), .A1(n3682), .Z(n3684));
Q_XNR2 U2424 ( .A0(_zyM2L299_pbcT3[22]), .A1(n3682), .Z(n3683));
Q_OR02 U2425 ( .A0(_zyM2L299_pbcT3[21]), .A1(n3680), .Z(n3682));
Q_XNR2 U2426 ( .A0(_zyM2L299_pbcT3[21]), .A1(n3680), .Z(n3681));
Q_OR02 U2427 ( .A0(_zyM2L299_pbcT3[20]), .A1(n3678), .Z(n3680));
Q_XNR2 U2428 ( .A0(_zyM2L299_pbcT3[20]), .A1(n3678), .Z(n3679));
Q_OR02 U2429 ( .A0(_zyM2L299_pbcT3[19]), .A1(n3676), .Z(n3678));
Q_XNR2 U2430 ( .A0(_zyM2L299_pbcT3[19]), .A1(n3676), .Z(n3677));
Q_OR02 U2431 ( .A0(_zyM2L299_pbcT3[18]), .A1(n3674), .Z(n3676));
Q_XNR2 U2432 ( .A0(_zyM2L299_pbcT3[18]), .A1(n3674), .Z(n3675));
Q_OR02 U2433 ( .A0(_zyM2L299_pbcT3[17]), .A1(n3672), .Z(n3674));
Q_XNR2 U2434 ( .A0(_zyM2L299_pbcT3[17]), .A1(n3672), .Z(n3673));
Q_OR02 U2435 ( .A0(_zyM2L299_pbcT3[16]), .A1(n3670), .Z(n3672));
Q_XNR2 U2436 ( .A0(_zyM2L299_pbcT3[16]), .A1(n3670), .Z(n3671));
Q_OR02 U2437 ( .A0(_zyM2L299_pbcT3[15]), .A1(n3668), .Z(n3670));
Q_XNR2 U2438 ( .A0(_zyM2L299_pbcT3[15]), .A1(n3668), .Z(n3669));
Q_OR02 U2439 ( .A0(_zyM2L299_pbcT3[14]), .A1(n3666), .Z(n3668));
Q_XNR2 U2440 ( .A0(_zyM2L299_pbcT3[14]), .A1(n3666), .Z(n3667));
Q_OR02 U2441 ( .A0(_zyM2L299_pbcT3[13]), .A1(n3664), .Z(n3666));
Q_XNR2 U2442 ( .A0(_zyM2L299_pbcT3[13]), .A1(n3664), .Z(n3665));
Q_OR02 U2443 ( .A0(_zyM2L299_pbcT3[12]), .A1(n3662), .Z(n3664));
Q_XNR2 U2444 ( .A0(_zyM2L299_pbcT3[12]), .A1(n3662), .Z(n3663));
Q_OR02 U2445 ( .A0(_zyM2L299_pbcT3[11]), .A1(n3660), .Z(n3662));
Q_XNR2 U2446 ( .A0(_zyM2L299_pbcT3[11]), .A1(n3660), .Z(n3661));
Q_OR02 U2447 ( .A0(_zyM2L299_pbcT3[10]), .A1(n3658), .Z(n3660));
Q_XNR2 U2448 ( .A0(_zyM2L299_pbcT3[10]), .A1(n3658), .Z(n3659));
Q_OR02 U2449 ( .A0(_zyM2L299_pbcT3[9]), .A1(n3656), .Z(n3658));
Q_XNR2 U2450 ( .A0(_zyM2L299_pbcT3[9]), .A1(n3656), .Z(n3657));
Q_OR02 U2451 ( .A0(_zyM2L299_pbcT3[8]), .A1(n3654), .Z(n3656));
Q_XNR2 U2452 ( .A0(_zyM2L299_pbcT3[8]), .A1(n3654), .Z(n3655));
Q_OR02 U2453 ( .A0(_zyM2L299_pbcT3[7]), .A1(n3652), .Z(n3654));
Q_XNR2 U2454 ( .A0(_zyM2L299_pbcT3[7]), .A1(n3652), .Z(n3653));
Q_OR02 U2455 ( .A0(_zyM2L299_pbcT3[6]), .A1(n3650), .Z(n3652));
Q_XNR2 U2456 ( .A0(_zyM2L299_pbcT3[6]), .A1(n3650), .Z(n3651));
Q_OR02 U2457 ( .A0(_zyM2L299_pbcT3[5]), .A1(n3648), .Z(n3650));
Q_XNR2 U2458 ( .A0(_zyM2L299_pbcT3[5]), .A1(n3648), .Z(n3649));
Q_OR02 U2459 ( .A0(_zyM2L299_pbcT3[4]), .A1(n3646), .Z(n3648));
Q_XNR2 U2460 ( .A0(_zyM2L299_pbcT3[4]), .A1(n3646), .Z(n3647));
Q_OR02 U2461 ( .A0(_zyM2L299_pbcT3[3]), .A1(n3644), .Z(n3646));
Q_XNR2 U2462 ( .A0(_zyM2L299_pbcT3[3]), .A1(n3644), .Z(n3645));
Q_OR02 U2463 ( .A0(_zyM2L299_pbcT3[2]), .A1(n3642), .Z(n3644));
Q_XNR2 U2464 ( .A0(_zyM2L299_pbcT3[2]), .A1(n3642), .Z(n3643));
Q_OR02 U2465 ( .A0(_zyM2L299_pbcT3[1]), .A1(_zyM2L299_pbcT3[0]), .Z(n3642));
Q_XNR2 U2466 ( .A0(_zyM2L299_pbcT3[1]), .A1(_zyM2L299_pbcT3[0]), .Z(n3641));
Q_XNR2 U2467 ( .A0(_zyGfifo__gfdL365_0_P0_m2_gfOff), .A1(_zyGfifoF0_L253_s4_req_6), .Z(n3639));
Q_XNR2 U2468 ( .A0(_zyGfifo__gfdL276_2_P0_m2_gfOff), .A1(_zyGfifoF0_L253_s4_req_6), .Z(n3638));
Q_XNR2 U2469 ( .A0(n3637), .A1(_zyGfifoF1_L253_s2_req_7), .Z(n4269));
Q_XNR2 U2470 ( .A0(_zyGfifo__gfdL268_4_P0_m2_gfOff), .A1(_zyGfifoF0_L253_s4_req_6), .Z(n3636));
Q_XNR2 U2471 ( .A0(_zyGfifo__gfdL265_5_P0_m2_gfOff), .A1(_zyGfifoF0_L253_s4_req_6), .Z(n3635));
Q_OR02 U2472 ( .A0(n3633), .A1(n3634), .Z(n5333));
Q_OR03 U2473 ( .A0(n3630), .A1(n3631), .A2(n3632), .Z(n3634));
Q_OR03 U2474 ( .A0(n3627), .A1(n3628), .A2(n3629), .Z(n3633));
Q_OR03 U2475 ( .A0(n3624), .A1(n3625), .A2(n3626), .Z(n3632));
Q_OR03 U2476 ( .A0(n3621), .A1(n3622), .A2(n3623), .Z(n3631));
Q_OR03 U2477 ( .A0(_zyictd_sysfunc_11_L263_5[1]), .A1(_zyictd_sysfunc_11_L263_5[0]), .A2(n3620), .Z(n3630));
Q_OR03 U2478 ( .A0(_zyictd_sysfunc_11_L263_5[4]), .A1(_zyictd_sysfunc_11_L263_5[3]), .A2(_zyictd_sysfunc_11_L263_5[2]), .Z(n3629));
Q_OR03 U2479 ( .A0(_zyictd_sysfunc_11_L263_5[7]), .A1(_zyictd_sysfunc_11_L263_5[6]), .A2(_zyictd_sysfunc_11_L263_5[5]), .Z(n3628));
Q_OR03 U2480 ( .A0(_zyictd_sysfunc_11_L263_5[10]), .A1(_zyictd_sysfunc_11_L263_5[9]), .A2(_zyictd_sysfunc_11_L263_5[8]), .Z(n3627));
Q_OR03 U2481 ( .A0(_zyictd_sysfunc_11_L263_5[13]), .A1(_zyictd_sysfunc_11_L263_5[12]), .A2(_zyictd_sysfunc_11_L263_5[11]), .Z(n3626));
Q_OR03 U2482 ( .A0(_zyictd_sysfunc_11_L263_5[16]), .A1(_zyictd_sysfunc_11_L263_5[15]), .A2(_zyictd_sysfunc_11_L263_5[14]), .Z(n3625));
Q_OR03 U2483 ( .A0(_zyictd_sysfunc_11_L263_5[19]), .A1(_zyictd_sysfunc_11_L263_5[18]), .A2(_zyictd_sysfunc_11_L263_5[17]), .Z(n3624));
Q_OR03 U2484 ( .A0(_zyictd_sysfunc_11_L263_5[22]), .A1(_zyictd_sysfunc_11_L263_5[21]), .A2(_zyictd_sysfunc_11_L263_5[20]), .Z(n3623));
Q_OR03 U2485 ( .A0(_zyictd_sysfunc_11_L263_5[25]), .A1(_zyictd_sysfunc_11_L263_5[24]), .A2(_zyictd_sysfunc_11_L263_5[23]), .Z(n3622));
Q_OR03 U2486 ( .A0(_zyictd_sysfunc_11_L263_5[28]), .A1(_zyictd_sysfunc_11_L263_5[27]), .A2(_zyictd_sysfunc_11_L263_5[26]), .Z(n3621));
Q_OR03 U2487 ( .A0(_zyictd_sysfunc_11_L263_5[31]), .A1(_zyictd_sysfunc_11_L263_5[30]), .A2(_zyictd_sysfunc_11_L263_5[29]), .Z(n3620));
Q_OR02 U2488 ( .A0(n3618), .A1(n3619), .Z(n5319));
Q_OR03 U2489 ( .A0(n3615), .A1(n3616), .A2(n3617), .Z(n3619));
Q_OR03 U2490 ( .A0(n3612), .A1(n3613), .A2(n3614), .Z(n3618));
Q_OR03 U2491 ( .A0(n3609), .A1(n3610), .A2(n3611), .Z(n3617));
Q_OR03 U2492 ( .A0(n3606), .A1(n3607), .A2(n3608), .Z(n3616));
Q_OR03 U2493 ( .A0(_zyictd_sysfunc_11_L257_2[1]), .A1(_zyictd_sysfunc_11_L257_2[0]), .A2(n3605), .Z(n3615));
Q_OR03 U2494 ( .A0(_zyictd_sysfunc_11_L257_2[4]), .A1(_zyictd_sysfunc_11_L257_2[3]), .A2(_zyictd_sysfunc_11_L257_2[2]), .Z(n3614));
Q_OR03 U2495 ( .A0(_zyictd_sysfunc_11_L257_2[7]), .A1(_zyictd_sysfunc_11_L257_2[6]), .A2(_zyictd_sysfunc_11_L257_2[5]), .Z(n3613));
Q_OR03 U2496 ( .A0(_zyictd_sysfunc_11_L257_2[10]), .A1(_zyictd_sysfunc_11_L257_2[9]), .A2(_zyictd_sysfunc_11_L257_2[8]), .Z(n3612));
Q_OR03 U2497 ( .A0(_zyictd_sysfunc_11_L257_2[13]), .A1(_zyictd_sysfunc_11_L257_2[12]), .A2(_zyictd_sysfunc_11_L257_2[11]), .Z(n3611));
Q_OR03 U2498 ( .A0(_zyictd_sysfunc_11_L257_2[16]), .A1(_zyictd_sysfunc_11_L257_2[15]), .A2(_zyictd_sysfunc_11_L257_2[14]), .Z(n3610));
Q_OR03 U2499 ( .A0(_zyictd_sysfunc_11_L257_2[19]), .A1(_zyictd_sysfunc_11_L257_2[18]), .A2(_zyictd_sysfunc_11_L257_2[17]), .Z(n3609));
Q_OR03 U2500 ( .A0(_zyictd_sysfunc_11_L257_2[22]), .A1(_zyictd_sysfunc_11_L257_2[21]), .A2(_zyictd_sysfunc_11_L257_2[20]), .Z(n3608));
Q_OR03 U2501 ( .A0(_zyictd_sysfunc_11_L257_2[25]), .A1(_zyictd_sysfunc_11_L257_2[24]), .A2(_zyictd_sysfunc_11_L257_2[23]), .Z(n3607));
Q_OR03 U2502 ( .A0(_zyictd_sysfunc_11_L257_2[28]), .A1(_zyictd_sysfunc_11_L257_2[27]), .A2(_zyictd_sysfunc_11_L257_2[26]), .Z(n3606));
Q_OR03 U2503 ( .A0(_zyictd_sysfunc_11_L257_2[31]), .A1(_zyictd_sysfunc_11_L257_2[30]), .A2(_zyictd_sysfunc_11_L257_2[29]), .Z(n3605));
Q_AN02 U2504 ( .A0(n446), .A1(n3094), .Z(n3603));
Q_OR02 U2505 ( .A0(n3558), .A1(n487), .Z(n3571));
Q_AN02 U2506 ( .A0(n446), .A1(n3000), .Z(n3570));
Q_OR02 U2507 ( .A0(n3291), .A1(n487), .Z(n3569));
Q_AN02 U2508 ( .A0(n446), .A1(n3554), .Z(n3568));
Q_INV U2509 ( .A(n3301), .Z(n3397));
Q_AN03 U2510 ( .A0(kme_ob_tvalid), .A1(n3543), .A2(n3298), .Z(n3396));
Q_MX02 U2511 ( .S(_zyL439_meState8[0]), .A0(n3396), .A1(n3397), .Z(n3395));
Q_INV U2512 ( .A(n3395), .Z(n3394));
Q_OR02 U2513 ( .A0(_zyL439_meState8[1]), .A1(n3394), .Z(n3393));
Q_INV U2514 ( .A(n3393), .Z(n3558));
Q_AN02 U2515 ( .A0(n3543), .A1(ready_ob), .Z(n3321));
Q_AO21 U2516 ( .A0(kme_ob_tvalid), .A1(n3321), .B0(_zyL439_meState8[0]), .Z(n3392));
Q_ND02 U2517 ( .A0(n3270), .A1(n3392), .Z(n3391));
Q_OR02 U2518 ( .A0(_zyL439_meState8[1]), .A1(n3391), .Z(n3390));
Q_OR03 U2519 ( .A0(user_string_ob[5]), .A1(n3389), .A2(n3387), .Z(n3385));
Q_OR02 U2520 ( .A0(user_string_ob[15]), .A1(n3388), .Z(n3387));
Q_ND02 U2521 ( .A0(user_string_ob[13]), .A1(user_string_ob[6]), .Z(n3386));
Q_OR03 U2522 ( .A0(user_string_ob[19]), .A1(user_string_ob[3]), .A2(n3386), .Z(n3384));
Q_OR03 U2523 ( .A0(n3384), .A1(n3385), .A2(n3381), .Z(n3334));
Q_ND02 U2524 ( .A0(user_string_ob[11]), .A1(user_string_ob[4]), .Z(n3383));
Q_OR03 U2525 ( .A0(user_string_ob[21]), .A1(user_string_ob[7]), .A2(n3383), .Z(n3382));
Q_OR02 U2526 ( .A0(user_string_ob[23]), .A1(n3382), .Z(n3381));
Q_OR03 U2527 ( .A0(user_string_ob[0]), .A1(n3549), .A2(n3380), .Z(n3379));
Q_OR02 U2528 ( .A0(n3336), .A1(user_string_ob[1]), .Z(n3380));
Q_OR02 U2529 ( .A0(n3548), .A1(n3335), .Z(n3378));
Q_OR03 U2530 ( .A0(user_string_ob[17]), .A1(n3378), .A2(n3379), .Z(n3377));
Q_OR02 U2531 ( .A0(n3332), .A1(user_string_ob[20]), .Z(n3376));
Q_OR03 U2532 ( .A0(n3375), .A1(n3376), .A2(n3377), .Z(n3374));
Q_OR02 U2533 ( .A0(n3564), .A1(user_string_ob[12]), .Z(n3375));
Q_OR03 U2534 ( .A0(n3374), .A1(n3334), .A2(n3372), .Z(n3371));
Q_ND02 U2535 ( .A0(user_string_ob[10]), .A1(n3216), .Z(n3373));
Q_OR03 U2536 ( .A0(n3330), .A1(n3373), .A2(user_string_ob[24]), .Z(n3372));
Q_OA21 U2537 ( .A0(n3371), .A1(n1885), .B0(n3366), .Z(n3368));
Q_OR03 U2538 ( .A0(n3548), .A1(n3549), .A2(n3370), .Z(n3369));
Q_OR02 U2539 ( .A0(n3563), .A1(n3564), .Z(n3370));
Q_OR02 U2540 ( .A0(n3369), .A1(n3562), .Z(n3366));
Q_MX02 U2541 ( .S(user_string_ob[18]), .A0(n3366), .A1(n3368), .Z(n3367));
Q_MX02 U2542 ( .S(n1774), .A0(n3367), .A1(n3366), .Z(n3365));
Q_MX02 U2543 ( .S(kme_ob_tvalid), .A0(n3564), .A1(n3365), .Z(n3364));
Q_OR02 U2544 ( .A0(n2130), .A1(n3537), .Z(n3248));
Q_INV U2545 ( .A(n3565), .Z(n3363));
Q_OR02 U2546 ( .A0(n3363), .A1(n3248), .Z(n3265));
Q_OR02 U2547 ( .A0(n2200), .A1(n3265), .Z(n3250));
Q_AN03 U2548 ( .A0(n2076), .A1(n3321), .A2(n3250), .Z(n3326));
Q_MX02 U2549 ( .S(n3540), .A0(n3326), .A1(n3321), .Z(n3362));
Q_MX02 U2550 ( .S(n2150), .A0(n3321), .A1(n3362), .Z(n3361));
Q_MX02 U2551 ( .S(n3207), .A0(n3321), .A1(n3361), .Z(n3360));
Q_AN02 U2552 ( .A0(kme_ob_tvalid), .A1(n3360), .Z(n3359));
Q_MX02 U2553 ( .S(_zyL439_meState8[0]), .A0(n3359), .A1(n3364), .Z(n3358));
Q_INV U2554 ( .A(n3358), .Z(n3357));
Q_OR02 U2555 ( .A0(_zyL439_meState8[1]), .A1(n3357), .Z(n3356));
Q_INV U2556 ( .A(n3356), .Z(n3551));
Q_OR02 U2557 ( .A0(n3315), .A1(n3566), .Z(n3271));
Q_OR02 U2558 ( .A0(n3543), .A1(n3271), .Z(n3355));
Q_MX02 U2559 ( .S(kme_ob_tvalid), .A0(n3355), .A1(n3271), .Z(n3354));
Q_NR02 U2560 ( .A0(_zyL439_meState8[0]), .A1(n3354), .Z(n3353));
Q_OA21 U2561 ( .A0(n3353), .A1(_zyL439_meState8[1]), .B0(n3267), .Z(n3352));
Q_AN02 U2562 ( .A0(kme_ob_tvalid), .A1(n3563), .Z(n3351));
Q_AN03 U2563 ( .A0(kme_ob_tvalid), .A1(n3561), .A2(n3321), .Z(n3289));
Q_MX02 U2564 ( .S(_zyL439_meState8[0]), .A0(n3289), .A1(n3351), .Z(n3350));
Q_INV U2565 ( .A(n3350), .Z(n3349));
Q_OR02 U2566 ( .A0(_zyL439_meState8[1]), .A1(n3349), .Z(n3348));
Q_AN02 U2567 ( .A0(kme_ob_tvalid), .A1(n3549), .Z(n3347));
Q_AN03 U2568 ( .A0(kme_ob_tvalid), .A1(n3542), .A2(n3321), .Z(n3346));
Q_MX02 U2569 ( .S(_zyL439_meState8[0]), .A0(n3346), .A1(n3347), .Z(n3345));
Q_INV U2570 ( .A(n3345), .Z(n3344));
Q_OR02 U2571 ( .A0(_zyL439_meState8[1]), .A1(n3344), .Z(n3343));
Q_AN02 U2572 ( .A0(kme_ob_tvalid), .A1(n3548), .Z(n3342));
Q_AN03 U2573 ( .A0(kme_ob_tvalid), .A1(n3540), .A2(n3321), .Z(n3341));
Q_MX02 U2574 ( .S(_zyL439_meState8[0]), .A0(n3341), .A1(n3342), .Z(n3340));
Q_INV U2575 ( .A(n3340), .Z(n3339));
Q_OR02 U2576 ( .A0(_zyL439_meState8[1]), .A1(n3339), .Z(n3338));
Q_OR03 U2577 ( .A0(user_string_ob[1]), .A1(user_string_ob[0]), .A2(n3337), .Z(n3333));
Q_ND02 U2578 ( .A0(user_string_ob[22]), .A1(user_string_ob[2]), .Z(n3337));
Q_OR02 U2579 ( .A0(n3333), .A1(n3334), .Z(n3306));
Q_OR03 U2580 ( .A0(user_string_ob[20]), .A1(user_string_ob[17]), .A2(n3307), .Z(n3331));
Q_OR02 U2581 ( .A0(user_string_ob[12]), .A1(n3332), .Z(n3307));
Q_OR03 U2582 ( .A0(n3259), .A1(n3331), .A2(n3306), .Z(n3309));
Q_ND02 U2583 ( .A0(user_string_ob[16]), .A1(n3567), .Z(n3330));
Q_OR03 U2584 ( .A0(user_string_ob[24]), .A1(n3330), .A2(n3309), .Z(n3266));
Q_AN02 U2585 ( .A0(n3562), .A1(n3266), .Z(n3329));
Q_MX02 U2586 ( .S(user_string_ob[18]), .A0(n3562), .A1(n3329), .Z(n3328));
Q_MX02 U2587 ( .S(n1774), .A0(n3328), .A1(n3562), .Z(n3547));
Q_AN02 U2588 ( .A0(kme_ob_tvalid), .A1(n3547), .Z(n3327));
Q_AN02 U2589 ( .A0(kme_ob_tvalid), .A1(n3326), .Z(n3325));
Q_MX02 U2590 ( .S(_zyL439_meState8[0]), .A0(n3325), .A1(n3327), .Z(n3324));
Q_INV U2591 ( .A(n3324), .Z(n3323));
Q_OR02 U2592 ( .A0(_zyL439_meState8[1]), .A1(n3323), .Z(n3322));
Q_INV U2593 ( .A(n3321), .Z(n3281));
Q_OR02 U2594 ( .A0(n3317), .A1(n3281), .Z(n3320));
Q_OR03 U2595 ( .A0(_zyL439_meState8[0]), .A1(n3315), .A2(_zyL439_meState8[1]), .Z(n3319));
Q_ND02 U2596 ( .A0(n2130), .A1(n2114), .Z(n3299));
Q_ND02 U2597 ( .A0(ready_ob), .A1(n3299), .Z(n3318));
Q_OR02 U2598 ( .A0(_zyL439_meState8[1]), .A1(_zyL439_meState8[0]), .Z(n3317));
Q_OR02 U2599 ( .A0(n3317), .A1(n3318), .Z(n3316));
Q_OR03 U2600 ( .A0(n3315), .A1(n3557), .A2(n3314), .Z(n3313));
Q_OR02 U2601 ( .A0(_zyL439_meState8[0]), .A1(n2432), .Z(n3314));
Q_OR02 U2602 ( .A0(_zyL439_meState8[1]), .A1(n3313), .Z(n3312));
Q_INV U2603 ( .A(n3312), .Z(n3559));
Q_ND02 U2604 ( .A0(_zyL439_meState8[0]), .A1(n3564), .Z(n3311));
Q_NR02 U2605 ( .A0(_zyL439_meState8[1]), .A1(n3311), .Z(n3310));
Q_OR02 U2606 ( .A0(user_string_ob[24]), .A1(n3258), .Z(n3305));
Q_OR02 U2607 ( .A0(n3305), .A1(n3309), .Z(n3264));
Q_ND02 U2608 ( .A0(user_string_ob[20]), .A1(user_string_ob[17]), .Z(n3308));
Q_OR03 U2609 ( .A0(n3307), .A1(n3308), .A2(n3306), .Z(n3257));
Q_OR03 U2610 ( .A0(n3259), .A1(n1778), .A2(n3305), .Z(n3304));
Q_OR02 U2611 ( .A0(n3304), .A1(n3257), .Z(n3303));
Q_MX02 U2612 ( .S(user_string_ob[18]), .A0(n3303), .A1(n3264), .Z(n3302));
Q_OR02 U2613 ( .A0(n3555), .A1(n1774), .Z(n3301));
Q_OR02 U2614 ( .A0(n3301), .A1(n3302), .Z(n3300));
Q_AN02 U2615 ( .A0(ready_ob), .A1(n3538), .Z(n3298));
Q_AN03 U2616 ( .A0(n3298), .A1(n3299), .A2(n3543), .Z(n3297));
Q_OA21 U2617 ( .A0(n3297), .A1(n1976), .B0(n3295), .Z(n3294));
Q_OR02 U2618 ( .A0(n2200), .A1(n3248), .Z(n3251));
Q_OR02 U2619 ( .A0(n3281), .A1(n3251), .Z(n3296));
Q_ND02 U2620 ( .A0(n3296), .A1(n1976), .Z(n3295));
Q_ND02 U2621 ( .A0(kme_ob_tvalid), .A1(n3294), .Z(n3293));
Q_MX02 U2622 ( .S(_zyL439_meState8[0]), .A0(n3293), .A1(n3300), .Z(n3292));
Q_NR02 U2623 ( .A0(_zyL439_meState8[1]), .A1(n3292), .Z(n3291));
Q_AO21 U2624 ( .A0(n3272), .A1(n3392), .B0(n487), .Z(n3604));
Q_OR02 U2625 ( .A0(n3560), .A1(n3557), .Z(n3290));
Q_INV U2626 ( .A(n3289), .Z(n3288));
Q_AO21 U2627 ( .A0(n3288), .A1(n3553), .B0(n3285), .Z(n3287));
Q_OR02 U2628 ( .A0(_zyL439_meState8[1]), .A1(n3287), .Z(n3286));
Q_AN02 U2629 ( .A0(_zyL439_meState8[0]), .A1(kme_ob_tvalid), .Z(n3285));
Q_INV U2630 ( .A(n3285), .Z(n3284));
Q_NR02 U2631 ( .A0(_zyL439_meState8[1]), .A1(n3284), .Z(n3283));
Q_ND02 U2632 ( .A0(kme_ob_tvalid), .A1(n3216), .Z(n3282));
Q_ND02 U2633 ( .A0(kme_ob_tvalid), .A1(n3207), .Z(n3280));
Q_NR02 U2634 ( .A0(n3280), .A1(n3281), .Z(n3279));
Q_MX02 U2635 ( .S(_zyL439_meState8[0]), .A0(n3279), .A1(n3282), .Z(n3278));
Q_INV U2636 ( .A(n3278), .Z(n3277));
Q_OR02 U2637 ( .A0(_zyL439_meState8[1]), .A1(n3277), .Z(n3276));
Q_INV U2638 ( .A(n3276), .Z(n3556));
Q_INV U2639 ( .A(kme_ob_tvalid), .Z(n3555));
Q_MX02 U2640 ( .S(_zyL439_meState8[0]), .A0(n3537), .A1(user_string_ob[17]), .Z(n3554));
Q_AO21 U2641 ( .A0(ready_ob), .A1(n3566), .B0(_zyL439_meState8[0]), .Z(n3275));
Q_ND02 U2642 ( .A0(n3270), .A1(n3275), .Z(n3274));
Q_NR02 U2643 ( .A0(_zyL439_meState8[1]), .A1(n3274), .Z(n3273));
Q_OR02 U2644 ( .A0(_zyL439_meState8[0]), .A1(n3272), .Z(n3267));
Q_OR02 U2645 ( .A0(kme_ob_tvalid), .A1(n3553), .Z(n3270));
Q_OA21 U2646 ( .A0(n3271), .A1(_zyL439_meState8[0]), .B0(n3270), .Z(n3269));
Q_INV U2647 ( .A(n3269), .Z(n3268));
Q_OA21 U2648 ( .A0(n3268), .A1(_zyL439_meState8[1]), .B0(n3267), .Z(n3552));
Q_OR02 U2649 ( .A0(n3263), .A1(n3266), .Z(n3261));
Q_AN02 U2650 ( .A0(_zyL439_meState8[0]), .A1(n3261), .Z(n3550));
Q_INV U2651 ( .A(_zyL439_meState8[0]), .Z(n3553));
Q_AN03 U2652 ( .A0(n3553), .A1(n3265), .A2(n3565), .Z(n2999));
Q_OR02 U2653 ( .A0(n3263), .A1(n3264), .Z(n3252));
Q_NR02 U2654 ( .A0(n1774), .A1(n3252), .Z(n3262));
Q_OR02 U2655 ( .A0(n1774), .A1(n3261), .Z(n3260));
Q_INV U2656 ( .A(n3546), .Z(n3217));
Q_ND02 U2657 ( .A0(user_string_ob[16]), .A1(user_string_ob[10]), .Z(n3256));
Q_OR02 U2658 ( .A0(n3256), .A1(n3257), .Z(n3254));
Q_OR03 U2659 ( .A0(user_string_ob[24]), .A1(n1782), .A2(user_string_ob[18]), .Z(n3255));
Q_NR02 U2660 ( .A0(n3255), .A1(n3254), .Z(n3544));
Q_OR03 U2661 ( .A0(user_string_ob[18]), .A1(user_string_ob[24]), .A2(n3254), .Z(n3253));
Q_INV U2662 ( .A(n3251), .Z(n3541));
Q_AN02 U2663 ( .A0(n2076), .A1(n3250), .Z(n3539));
Q_NR02 U2664 ( .A0(n2114), .A1(n1980), .Z(n3249));
Q_INV U2665 ( .A(n3248), .Z(n3536));
Q_MX02 U2666 ( .S(n3553), .A0(n3253), .A1(n2114), .Z(n3247));
Q_MX02 U2667 ( .S(n3553), .A0(n3252), .A1(n3248), .Z(n3246));
Q_MX02 U2668 ( .S(n3553), .A0(n3210), .A1(n3203), .Z(n3245));
Q_MX02 U2669 ( .S(n3553), .A0(n3209), .A1(n3202), .Z(n3244));
Q_AN02 U2670 ( .A0(_zyL439_meState8[0]), .A1(user_string_ob[24]), .Z(n3243));
Q_AN02 U2671 ( .A0(_zyL439_meState8[0]), .A1(user_string_ob[23]), .Z(n3242));
Q_MX02 U2672 ( .S(n3553), .A0(user_string_ob[22]), .A1(n3201), .Z(n3241));
Q_AN02 U2673 ( .A0(_zyL439_meState8[0]), .A1(user_string_ob[21]), .Z(n3240));
Q_MX02 U2674 ( .S(n3553), .A0(user_string_ob[20]), .A1(n3537), .Z(n3239));
Q_AN02 U2675 ( .A0(_zyL439_meState8[0]), .A1(user_string_ob[19]), .Z(n3238));
Q_MX02 U2676 ( .S(n3553), .A0(user_string_ob[18]), .A1(n3536), .Z(n3237));
Q_MX02 U2677 ( .S(n3553), .A0(user_string_ob[17]), .A1(n3537), .Z(n3236));
Q_MX02 U2678 ( .S(n3553), .A0(user_string_ob[16]), .A1(n3201), .Z(n3235));
Q_AN02 U2679 ( .A0(_zyL439_meState8[0]), .A1(user_string_ob[15]), .Z(n3234));
Q_MX02 U2680 ( .S(n3553), .A0(user_string_ob[14]), .A1(n3201), .Z(n3233));
Q_MX02 U2681 ( .S(n3553), .A0(user_string_ob[13]), .A1(n3201), .Z(n3232));
Q_AN02 U2682 ( .A0(_zyL439_meState8[0]), .A1(user_string_ob[12]), .Z(n3231));
Q_MX02 U2683 ( .S(n3553), .A0(user_string_ob[11]), .A1(n3201), .Z(n3230));
Q_MX02 U2684 ( .S(n3553), .A0(user_string_ob[10]), .A1(n3201), .Z(n3229));
Q_MX02 U2685 ( .S(n3553), .A0(user_string_ob[9]), .A1(n3201), .Z(n3228));
Q_MX02 U2686 ( .S(n3553), .A0(user_string_ob[8]), .A1(n3201), .Z(n3227));
Q_AN02 U2687 ( .A0(_zyL439_meState8[0]), .A1(user_string_ob[7]), .Z(n3226));
Q_MX02 U2688 ( .S(n3553), .A0(user_string_ob[6]), .A1(n3201), .Z(n3225));
Q_AN02 U2689 ( .A0(_zyL439_meState8[0]), .A1(user_string_ob[5]), .Z(n3224));
Q_MX02 U2690 ( .S(n3553), .A0(user_string_ob[4]), .A1(n3201), .Z(n3223));
Q_AN02 U2691 ( .A0(_zyL439_meState8[0]), .A1(user_string_ob[3]), .Z(n3222));
Q_MX02 U2692 ( .S(n3553), .A0(user_string_ob[2]), .A1(n3201), .Z(n3221));
Q_AN02 U2693 ( .A0(_zyL439_meState8[0]), .A1(user_string_ob[1]), .Z(n3220));
Q_AN02 U2694 ( .A0(_zyL439_meState8[0]), .A1(user_string_ob[0]), .Z(n3219));
Q_MX02 U2695 ( .S(_zyL439_meState8[0]), .A0(n3541), .A1(n3262), .Z(n3218));
Q_MX02 U2696 ( .S(_zyL439_meState8[0]), .A0(n3250), .A1(n3260), .Z(n3546));
Q_NR02 U2697 ( .A0(n1789), .A1(n3557), .Z(n3543));
Q_INV U2698 ( .A(n3216), .Z(n3563));
Q_XNR2 U2699 ( .A0(kme_ob_tlast), .A1(n3262), .Z(n3216));
Q_OR02 U2700 ( .A0(n3214), .A1(n3215), .Z(n3548));
Q_OR03 U2701 ( .A0(n3212), .A1(n3211), .A2(n3213), .Z(n3215));
Q_OR03 U2702 ( .A0(kme_ob_tuser[4]), .A1(kme_ob_tuser[3]), .A2(kme_ob_tuser[2]), .Z(n3214));
Q_OR03 U2703 ( .A0(kme_ob_tuser[7]), .A1(kme_ob_tuser[6]), .A2(kme_ob_tuser[5]), .Z(n3213));
Q_XOR2 U2704 ( .A0(kme_ob_tuser[1]), .A1(n3210), .Z(n3212));
Q_XOR2 U2705 ( .A0(kme_ob_tuser[0]), .A1(n3209), .Z(n3211));
Q_AN02 U2706 ( .A0(n3545), .A1(n3253), .Z(n3210));
Q_AN02 U2707 ( .A0(n3545), .A1(n3252), .Z(n3209));
Q_OR02 U2708 ( .A0(n3208), .A1(kme_ob_tvalid), .Z(n3566));
Q_INV U2709 ( .A(n3543), .Z(n3208));
Q_INV U2710 ( .A(n3207), .Z(n3561));
Q_XNR2 U2711 ( .A0(kme_ob_tlast), .A1(n3541), .Z(n3207));
Q_OR02 U2712 ( .A0(n3214), .A1(n3206), .Z(n3540));
Q_OR03 U2713 ( .A0(n3205), .A1(n3204), .A2(n3213), .Z(n3206));
Q_XOR2 U2714 ( .A0(kme_ob_tuser[1]), .A1(n3203), .Z(n3205));
Q_XOR2 U2715 ( .A0(kme_ob_tuser[0]), .A1(n3202), .Z(n3204));
Q_AN02 U2716 ( .A0(n3538), .A1(n2114), .Z(n3203));
Q_AN02 U2717 ( .A0(n3538), .A1(n3248), .Z(n3202));
Q_FDP0 _zzM2L439_mdxP4_error_cntr_Dwen0_REG  ( .CK(clk), .D(n3551), .Q(_zzM2L439_mdxP4_error_cntr_Dwen0), .QN( ));
Q_XNR2 U2719 ( .A0(n3536), .A1(n2114), .Z(n3201));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[0] ( .CK(clk), .D(n3097), .Q(_zzM2L439_mdxP4_error_cntr_wr0[0]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[1] ( .CK(clk), .D(n3100), .Q(_zzM2L439_mdxP4_error_cntr_wr0[1]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[2] ( .CK(clk), .D(n3103), .Q(_zzM2L439_mdxP4_error_cntr_wr0[2]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[3] ( .CK(clk), .D(n3106), .Q(_zzM2L439_mdxP4_error_cntr_wr0[3]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[4] ( .CK(clk), .D(n3109), .Q(_zzM2L439_mdxP4_error_cntr_wr0[4]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[5] ( .CK(clk), .D(n3112), .Q(_zzM2L439_mdxP4_error_cntr_wr0[5]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[6] ( .CK(clk), .D(n3115), .Q(_zzM2L439_mdxP4_error_cntr_wr0[6]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[7] ( .CK(clk), .D(n3118), .Q(_zzM2L439_mdxP4_error_cntr_wr0[7]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[8] ( .CK(clk), .D(n3121), .Q(_zzM2L439_mdxP4_error_cntr_wr0[8]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[9] ( .CK(clk), .D(n3124), .Q(_zzM2L439_mdxP4_error_cntr_wr0[9]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[10] ( .CK(clk), .D(n3127), .Q(_zzM2L439_mdxP4_error_cntr_wr0[10]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[11] ( .CK(clk), .D(n3130), .Q(_zzM2L439_mdxP4_error_cntr_wr0[11]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[12] ( .CK(clk), .D(n3133), .Q(_zzM2L439_mdxP4_error_cntr_wr0[12]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[13] ( .CK(clk), .D(n3136), .Q(_zzM2L439_mdxP4_error_cntr_wr0[13]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[14] ( .CK(clk), .D(n3139), .Q(_zzM2L439_mdxP4_error_cntr_wr0[14]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[15] ( .CK(clk), .D(n3142), .Q(_zzM2L439_mdxP4_error_cntr_wr0[15]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[16] ( .CK(clk), .D(n3145), .Q(_zzM2L439_mdxP4_error_cntr_wr0[16]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[17] ( .CK(clk), .D(n3148), .Q(_zzM2L439_mdxP4_error_cntr_wr0[17]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[18] ( .CK(clk), .D(n3151), .Q(_zzM2L439_mdxP4_error_cntr_wr0[18]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[19] ( .CK(clk), .D(n3154), .Q(_zzM2L439_mdxP4_error_cntr_wr0[19]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[20] ( .CK(clk), .D(n3157), .Q(_zzM2L439_mdxP4_error_cntr_wr0[20]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[21] ( .CK(clk), .D(n3160), .Q(_zzM2L439_mdxP4_error_cntr_wr0[21]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[22] ( .CK(clk), .D(n3163), .Q(_zzM2L439_mdxP4_error_cntr_wr0[22]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[23] ( .CK(clk), .D(n3166), .Q(_zzM2L439_mdxP4_error_cntr_wr0[23]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[24] ( .CK(clk), .D(n3169), .Q(_zzM2L439_mdxP4_error_cntr_wr0[24]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[25] ( .CK(clk), .D(n3172), .Q(_zzM2L439_mdxP4_error_cntr_wr0[25]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[26] ( .CK(clk), .D(n3175), .Q(_zzM2L439_mdxP4_error_cntr_wr0[26]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[27] ( .CK(clk), .D(n3178), .Q(_zzM2L439_mdxP4_error_cntr_wr0[27]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[28] ( .CK(clk), .D(n3181), .Q(_zzM2L439_mdxP4_error_cntr_wr0[28]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[29] ( .CK(clk), .D(n3184), .Q(_zzM2L439_mdxP4_error_cntr_wr0[29]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[30] ( .CK(clk), .D(n3187), .Q(_zzM2L439_mdxP4_error_cntr_wr0[30]), .QN( ));
Q_FDP0 \_zzM2L439_mdxP4_error_cntr_wr0_REG[31] ( .CK(clk), .D(n3190), .Q(_zzM2L439_mdxP4_error_cntr_wr0[31]), .QN( ));
Q_MX02 U2752 ( .S(n3290), .A0(n2431), .A1(n3199), .Z(n3200));
Q_AN02 U2753 ( .A0(n3557), .A1(n2394), .Z(n3199));
Q_MX02 U2754 ( .S(n3290), .A0(n2430), .A1(n3197), .Z(n3198));
Q_AN02 U2755 ( .A0(n3557), .A1(n2393), .Z(n3197));
Q_MX02 U2756 ( .S(n3290), .A0(n2429), .A1(n3195), .Z(n3196));
Q_AN02 U2757 ( .A0(n3557), .A1(n2392), .Z(n3195));
Q_MX02 U2758 ( .S(n3290), .A0(n2428), .A1(n3193), .Z(n3194));
Q_AN02 U2759 ( .A0(n3557), .A1(n2391), .Z(n3193));
Q_MX02 U2760 ( .S(n3290), .A0(n2427), .A1(n3191), .Z(n3192));
Q_AN02 U2761 ( .A0(n3557), .A1(n2390), .Z(n3191));
Q_MX02 U2762 ( .S(n3286), .A0(n3188), .A1(n3189), .Z(n3190));
Q_MX04 U2763 ( .S0(n3556), .S1(n3283), .A0(error_cntr[31]), .A1(n2687), .A2(n2937), .A3(n2998), .Z(n3189));
Q_MX02 U2764 ( .S(n3276), .A0(n2529), .A1(n2813), .Z(n3188));
Q_MX02 U2765 ( .S(n3286), .A0(n3185), .A1(n3186), .Z(n3187));
Q_MX04 U2766 ( .S0(n3556), .S1(n3283), .A0(error_cntr[30]), .A1(n2686), .A2(n2936), .A3(n2996), .Z(n3186));
Q_MX02 U2767 ( .S(n3276), .A0(n2527), .A1(n2811), .Z(n3185));
Q_MX02 U2768 ( .S(n3286), .A0(n3182), .A1(n3183), .Z(n3184));
Q_MX04 U2769 ( .S0(n3556), .S1(n3283), .A0(error_cntr[29]), .A1(n2685), .A2(n2935), .A3(n2994), .Z(n3183));
Q_MX02 U2770 ( .S(n3276), .A0(n2525), .A1(n2809), .Z(n3182));
Q_MX02 U2771 ( .S(n3286), .A0(n3179), .A1(n3180), .Z(n3181));
Q_MX04 U2772 ( .S0(n3556), .S1(n3283), .A0(error_cntr[28]), .A1(n2684), .A2(n2934), .A3(n2992), .Z(n3180));
Q_MX02 U2773 ( .S(n3276), .A0(n2523), .A1(n2807), .Z(n3179));
Q_MX02 U2774 ( .S(n3286), .A0(n3176), .A1(n3177), .Z(n3178));
Q_MX04 U2775 ( .S0(n3556), .S1(n3283), .A0(error_cntr[27]), .A1(n2683), .A2(n2933), .A3(n2990), .Z(n3177));
Q_MX02 U2776 ( .S(n3276), .A0(n2521), .A1(n2805), .Z(n3176));
Q_MX02 U2777 ( .S(n3286), .A0(n3173), .A1(n3174), .Z(n3175));
Q_MX04 U2778 ( .S0(n3556), .S1(n3283), .A0(error_cntr[26]), .A1(n2682), .A2(n2932), .A3(n2988), .Z(n3174));
Q_MX02 U2779 ( .S(n3276), .A0(n2519), .A1(n2803), .Z(n3173));
Q_MX02 U2780 ( .S(n3286), .A0(n3170), .A1(n3171), .Z(n3172));
Q_MX04 U2781 ( .S0(n3556), .S1(n3283), .A0(error_cntr[25]), .A1(n2681), .A2(n2931), .A3(n2986), .Z(n3171));
Q_MX02 U2782 ( .S(n3276), .A0(n2517), .A1(n2801), .Z(n3170));
Q_MX02 U2783 ( .S(n3286), .A0(n3167), .A1(n3168), .Z(n3169));
Q_MX04 U2784 ( .S0(n3556), .S1(n3283), .A0(error_cntr[24]), .A1(n2680), .A2(n2930), .A3(n2984), .Z(n3168));
Q_MX02 U2785 ( .S(n3276), .A0(n2515), .A1(n2799), .Z(n3167));
Q_MX02 U2786 ( .S(n3286), .A0(n3164), .A1(n3165), .Z(n3166));
Q_MX04 U2787 ( .S0(n3556), .S1(n3283), .A0(error_cntr[23]), .A1(n2679), .A2(n2929), .A3(n2982), .Z(n3165));
Q_MX02 U2788 ( .S(n3276), .A0(n2513), .A1(n2797), .Z(n3164));
Q_MX02 U2789 ( .S(n3286), .A0(n3161), .A1(n3162), .Z(n3163));
Q_MX04 U2790 ( .S0(n3556), .S1(n3283), .A0(error_cntr[22]), .A1(n2678), .A2(n2928), .A3(n2980), .Z(n3162));
Q_MX02 U2791 ( .S(n3276), .A0(n2511), .A1(n2795), .Z(n3161));
Q_MX02 U2792 ( .S(n3286), .A0(n3158), .A1(n3159), .Z(n3160));
Q_MX04 U2793 ( .S0(n3556), .S1(n3283), .A0(error_cntr[21]), .A1(n2677), .A2(n2927), .A3(n2978), .Z(n3159));
Q_MX02 U2794 ( .S(n3276), .A0(n2509), .A1(n2793), .Z(n3158));
Q_MX02 U2795 ( .S(n3286), .A0(n3155), .A1(n3156), .Z(n3157));
Q_MX04 U2796 ( .S0(n3556), .S1(n3283), .A0(error_cntr[20]), .A1(n2676), .A2(n2926), .A3(n2976), .Z(n3156));
Q_MX02 U2797 ( .S(n3276), .A0(n2507), .A1(n2791), .Z(n3155));
Q_MX02 U2798 ( .S(n3286), .A0(n3152), .A1(n3153), .Z(n3154));
Q_MX04 U2799 ( .S0(n3556), .S1(n3283), .A0(error_cntr[19]), .A1(n2675), .A2(n2925), .A3(n2974), .Z(n3153));
Q_MX02 U2800 ( .S(n3276), .A0(n2505), .A1(n2789), .Z(n3152));
Q_MX02 U2801 ( .S(n3286), .A0(n3149), .A1(n3150), .Z(n3151));
Q_MX04 U2802 ( .S0(n3556), .S1(n3283), .A0(error_cntr[18]), .A1(n2674), .A2(n2924), .A3(n2972), .Z(n3150));
Q_MX02 U2803 ( .S(n3276), .A0(n2503), .A1(n2787), .Z(n3149));
Q_MX02 U2804 ( .S(n3286), .A0(n3146), .A1(n3147), .Z(n3148));
Q_MX04 U2805 ( .S0(n3556), .S1(n3283), .A0(error_cntr[17]), .A1(n2673), .A2(n2923), .A3(n2970), .Z(n3147));
Q_MX02 U2806 ( .S(n3276), .A0(n2501), .A1(n2785), .Z(n3146));
Q_MX02 U2807 ( .S(n3286), .A0(n3143), .A1(n3144), .Z(n3145));
Q_MX04 U2808 ( .S0(n3556), .S1(n3283), .A0(error_cntr[16]), .A1(n2672), .A2(n2922), .A3(n2968), .Z(n3144));
Q_MX02 U2809 ( .S(n3276), .A0(n2499), .A1(n2783), .Z(n3143));
Q_MX02 U2810 ( .S(n3286), .A0(n3140), .A1(n3141), .Z(n3142));
Q_MX04 U2811 ( .S0(n3556), .S1(n3283), .A0(error_cntr[15]), .A1(n2671), .A2(n2921), .A3(n2966), .Z(n3141));
Q_MX02 U2812 ( .S(n3276), .A0(n2497), .A1(n2781), .Z(n3140));
Q_MX02 U2813 ( .S(n3286), .A0(n3137), .A1(n3138), .Z(n3139));
Q_MX04 U2814 ( .S0(n3556), .S1(n3283), .A0(error_cntr[14]), .A1(n2670), .A2(n2920), .A3(n2964), .Z(n3138));
Q_MX02 U2815 ( .S(n3276), .A0(n2495), .A1(n2779), .Z(n3137));
Q_MX02 U2816 ( .S(n3286), .A0(n3134), .A1(n3135), .Z(n3136));
Q_MX04 U2817 ( .S0(n3556), .S1(n3283), .A0(error_cntr[13]), .A1(n2669), .A2(n2919), .A3(n2962), .Z(n3135));
Q_MX02 U2818 ( .S(n3276), .A0(n2493), .A1(n2777), .Z(n3134));
Q_MX02 U2819 ( .S(n3286), .A0(n3131), .A1(n3132), .Z(n3133));
Q_MX04 U2820 ( .S0(n3556), .S1(n3283), .A0(error_cntr[12]), .A1(n2668), .A2(n2918), .A3(n2960), .Z(n3132));
Q_MX02 U2821 ( .S(n3276), .A0(n2491), .A1(n2775), .Z(n3131));
Q_MX02 U2822 ( .S(n3286), .A0(n3128), .A1(n3129), .Z(n3130));
Q_MX04 U2823 ( .S0(n3556), .S1(n3283), .A0(error_cntr[11]), .A1(n2667), .A2(n2917), .A3(n2958), .Z(n3129));
Q_MX02 U2824 ( .S(n3276), .A0(n2489), .A1(n2773), .Z(n3128));
Q_MX02 U2825 ( .S(n3286), .A0(n3125), .A1(n3126), .Z(n3127));
Q_MX04 U2826 ( .S0(n3556), .S1(n3283), .A0(error_cntr[10]), .A1(n2666), .A2(n2916), .A3(n2956), .Z(n3126));
Q_MX02 U2827 ( .S(n3276), .A0(n2487), .A1(n2771), .Z(n3125));
Q_MX02 U2828 ( .S(n3286), .A0(n3122), .A1(n3123), .Z(n3124));
Q_MX04 U2829 ( .S0(n3556), .S1(n3283), .A0(error_cntr[9]), .A1(n2665), .A2(n2915), .A3(n2954), .Z(n3123));
Q_MX02 U2830 ( .S(n3276), .A0(n2485), .A1(n2769), .Z(n3122));
Q_MX02 U2831 ( .S(n3286), .A0(n3119), .A1(n3120), .Z(n3121));
Q_MX04 U2832 ( .S0(n3556), .S1(n3283), .A0(error_cntr[8]), .A1(n2664), .A2(n2914), .A3(n2952), .Z(n3120));
Q_MX02 U2833 ( .S(n3276), .A0(n2483), .A1(n2767), .Z(n3119));
Q_MX02 U2834 ( .S(n3286), .A0(n3116), .A1(n3117), .Z(n3118));
Q_MX04 U2835 ( .S0(n3556), .S1(n3283), .A0(error_cntr[7]), .A1(n2663), .A2(n2913), .A3(n2950), .Z(n3117));
Q_MX02 U2836 ( .S(n3276), .A0(n2481), .A1(n2765), .Z(n3116));
Q_MX02 U2837 ( .S(n3286), .A0(n3113), .A1(n3114), .Z(n3115));
Q_MX04 U2838 ( .S0(n3556), .S1(n3283), .A0(error_cntr[6]), .A1(n2662), .A2(n2912), .A3(n2948), .Z(n3114));
Q_MX02 U2839 ( .S(n3276), .A0(n2479), .A1(n2763), .Z(n3113));
Q_MX02 U2840 ( .S(n3286), .A0(n3110), .A1(n3111), .Z(n3112));
Q_MX04 U2841 ( .S0(n3556), .S1(n3283), .A0(error_cntr[5]), .A1(n2661), .A2(n2911), .A3(n2946), .Z(n3111));
Q_MX02 U2842 ( .S(n3276), .A0(n2477), .A1(n2761), .Z(n3110));
Q_MX02 U2843 ( .S(n3286), .A0(n3107), .A1(n3108), .Z(n3109));
Q_MX04 U2844 ( .S0(n3556), .S1(n3283), .A0(error_cntr[4]), .A1(n2660), .A2(n2910), .A3(n2944), .Z(n3108));
Q_MX02 U2845 ( .S(n3276), .A0(n2475), .A1(n2759), .Z(n3107));
Q_MX02 U2846 ( .S(n3286), .A0(n3104), .A1(n3105), .Z(n3106));
Q_MX04 U2847 ( .S0(n3556), .S1(n3283), .A0(error_cntr[3]), .A1(n2659), .A2(n2909), .A3(n2942), .Z(n3105));
Q_MX02 U2848 ( .S(n3276), .A0(n2473), .A1(n2757), .Z(n3104));
Q_MX02 U2849 ( .S(n3286), .A0(n3101), .A1(n3102), .Z(n3103));
Q_MX04 U2850 ( .S0(n3556), .S1(n3283), .A0(error_cntr[2]), .A1(n2658), .A2(n2908), .A3(n2940), .Z(n3102));
Q_MX02 U2851 ( .S(n3276), .A0(n2471), .A1(n2755), .Z(n3101));
Q_MX02 U2852 ( .S(n3286), .A0(n3098), .A1(n3099), .Z(n3100));
Q_MX04 U2853 ( .S0(n3556), .S1(n3283), .A0(error_cntr[1]), .A1(n2657), .A2(n2907), .A3(n2938), .Z(n3099));
Q_MX02 U2854 ( .S(n3276), .A0(n2469), .A1(n2753), .Z(n3098));
Q_MX02 U2855 ( .S(n3286), .A0(n3095), .A1(n3096), .Z(n3097));
Q_MX02 U2856 ( .S(n3276), .A0(n2467), .A1(n2752), .Z(n3095));
Q_AN03 U2857 ( .A0(n3555), .A1(n2355), .A2(n446), .Z(n3572));
Q_AN03 U2858 ( .A0(n3555), .A1(n2353), .A2(n446), .Z(n3573));
Q_AN03 U2859 ( .A0(n3555), .A1(n2351), .A2(n446), .Z(n3574));
Q_AN03 U2860 ( .A0(n3555), .A1(n2349), .A2(n446), .Z(n3575));
Q_AN03 U2861 ( .A0(n3555), .A1(n2347), .A2(n446), .Z(n3576));
Q_AN03 U2862 ( .A0(n3555), .A1(n2345), .A2(n446), .Z(n3577));
Q_AN03 U2863 ( .A0(n3555), .A1(n2343), .A2(n446), .Z(n3578));
Q_AN03 U2864 ( .A0(n3555), .A1(n2341), .A2(n446), .Z(n3579));
Q_AN03 U2865 ( .A0(n3555), .A1(n2339), .A2(n446), .Z(n3580));
Q_AN03 U2866 ( .A0(n3555), .A1(n2337), .A2(n446), .Z(n3581));
Q_AN03 U2867 ( .A0(n3555), .A1(n2335), .A2(n446), .Z(n3582));
Q_AN03 U2868 ( .A0(n3555), .A1(n2333), .A2(n446), .Z(n3583));
Q_AN03 U2869 ( .A0(n3555), .A1(n2331), .A2(n446), .Z(n3584));
Q_AN03 U2870 ( .A0(n3555), .A1(n2329), .A2(n446), .Z(n3585));
Q_AN03 U2871 ( .A0(n3555), .A1(n2327), .A2(n446), .Z(n3586));
Q_AN03 U2872 ( .A0(n3555), .A1(n2325), .A2(n446), .Z(n3587));
Q_AN03 U2873 ( .A0(n3555), .A1(n2323), .A2(n446), .Z(n3588));
Q_AN03 U2874 ( .A0(n3555), .A1(n2321), .A2(n446), .Z(n3589));
Q_AN03 U2875 ( .A0(n3555), .A1(n2319), .A2(n446), .Z(n3590));
Q_AN03 U2876 ( .A0(n3555), .A1(n2317), .A2(n446), .Z(n3591));
Q_AN03 U2877 ( .A0(n3555), .A1(n2315), .A2(n446), .Z(n3592));
Q_AN03 U2878 ( .A0(n3555), .A1(n2313), .A2(n446), .Z(n3593));
Q_AN03 U2879 ( .A0(n3555), .A1(n2311), .A2(n446), .Z(n3594));
Q_AN03 U2880 ( .A0(n3555), .A1(n2309), .A2(n446), .Z(n3595));
Q_AN03 U2881 ( .A0(n3555), .A1(n2307), .A2(n446), .Z(n3596));
Q_AN03 U2882 ( .A0(n3555), .A1(n2305), .A2(n446), .Z(n3597));
Q_AN03 U2883 ( .A0(n3555), .A1(n2303), .A2(n446), .Z(n3598));
Q_AN03 U2884 ( .A0(n3555), .A1(n2301), .A2(n446), .Z(n3599));
Q_AN03 U2885 ( .A0(n3555), .A1(n2299), .A2(n446), .Z(n3600));
Q_AN03 U2886 ( .A0(n3555), .A1(n2297), .A2(n446), .Z(n3601));
Q_AN03 U2887 ( .A0(n3555), .A1(n2295), .A2(n446), .Z(n3602));
Q_NR02 U2888 ( .A0(kme_ob_tvalid), .A1(watchdog_timer[0]), .Z(n3094));
Q_MX02 U2889 ( .S(n2114), .A0(_zyGfifo__gfdL519_16_P0_m2_gfOff), .A1(_zyGfifo__gfdL522_15_P0_m2_gfOff), .Z(n1899));
Q_MX02 U2890 ( .S(n2114), .A0(_zyGfifo__gfdL519_16_P0_m2_cbid[19]), .A1(_zyGfifo__gfdL522_15_P0_m2_cbid[19]), .Z(n3092));
Q_MX02 U2891 ( .S(n2114), .A0(_zyGfifo__gfdL519_16_P0_m2_cbid[18]), .A1(_zyGfifo__gfdL522_15_P0_m2_cbid[18]), .Z(n3091));
Q_MX02 U2892 ( .S(n2114), .A0(_zyGfifo__gfdL519_16_P0_m2_cbid[17]), .A1(_zyGfifo__gfdL522_15_P0_m2_cbid[17]), .Z(n3090));
Q_MX02 U2893 ( .S(n2114), .A0(_zyGfifo__gfdL519_16_P0_m2_cbid[16]), .A1(_zyGfifo__gfdL522_15_P0_m2_cbid[16]), .Z(n3089));
Q_MX02 U2894 ( .S(n2114), .A0(_zyGfifo__gfdL519_16_P0_m2_cbid[15]), .A1(_zyGfifo__gfdL522_15_P0_m2_cbid[15]), .Z(n3088));
Q_MX02 U2895 ( .S(n2114), .A0(_zyGfifo__gfdL519_16_P0_m2_cbid[14]), .A1(_zyGfifo__gfdL522_15_P0_m2_cbid[14]), .Z(n3087));
Q_MX02 U2896 ( .S(n2114), .A0(_zyGfifo__gfdL519_16_P0_m2_cbid[13]), .A1(_zyGfifo__gfdL522_15_P0_m2_cbid[13]), .Z(n3086));
Q_MX02 U2897 ( .S(n2114), .A0(_zyGfifo__gfdL519_16_P0_m2_cbid[12]), .A1(_zyGfifo__gfdL522_15_P0_m2_cbid[12]), .Z(n3085));
Q_MX02 U2898 ( .S(n2114), .A0(_zyGfifo__gfdL519_16_P0_m2_cbid[11]), .A1(_zyGfifo__gfdL522_15_P0_m2_cbid[11]), .Z(n3084));
Q_MX02 U2899 ( .S(n2114), .A0(_zyGfifo__gfdL519_16_P0_m2_cbid[10]), .A1(_zyGfifo__gfdL522_15_P0_m2_cbid[10]), .Z(n3083));
Q_MX02 U2900 ( .S(n2114), .A0(_zyGfifo__gfdL519_16_P0_m2_cbid[9]), .A1(_zyGfifo__gfdL522_15_P0_m2_cbid[9]), .Z(n3082));
Q_MX02 U2901 ( .S(n2114), .A0(_zyGfifo__gfdL519_16_P0_m2_cbid[8]), .A1(_zyGfifo__gfdL522_15_P0_m2_cbid[8]), .Z(n3081));
Q_MX02 U2902 ( .S(n2114), .A0(_zyGfifo__gfdL519_16_P0_m2_cbid[7]), .A1(_zyGfifo__gfdL522_15_P0_m2_cbid[7]), .Z(n3080));
Q_MX02 U2903 ( .S(n2114), .A0(_zyGfifo__gfdL519_16_P0_m2_cbid[6]), .A1(_zyGfifo__gfdL522_15_P0_m2_cbid[6]), .Z(n3079));
Q_MX02 U2904 ( .S(n2114), .A0(_zyGfifo__gfdL519_16_P0_m2_cbid[5]), .A1(_zyGfifo__gfdL522_15_P0_m2_cbid[5]), .Z(n3078));
Q_MX02 U2905 ( .S(n2114), .A0(_zyGfifo__gfdL519_16_P0_m2_cbid[4]), .A1(_zyGfifo__gfdL522_15_P0_m2_cbid[4]), .Z(n3077));
Q_MX02 U2906 ( .S(n2114), .A0(_zyGfifo__gfdL519_16_P0_m2_cbid[3]), .A1(_zyGfifo__gfdL522_15_P0_m2_cbid[3]), .Z(n3076));
Q_MX02 U2907 ( .S(n2114), .A0(_zyGfifo__gfdL519_16_P0_m2_cbid[2]), .A1(_zyGfifo__gfdL522_15_P0_m2_cbid[2]), .Z(n3075));
Q_MX02 U2908 ( .S(n2114), .A0(_zyGfifo__gfdL519_16_P0_m2_cbid[1]), .A1(_zyGfifo__gfdL522_15_P0_m2_cbid[1]), .Z(n3074));
Q_MX02 U2909 ( .S(n2114), .A0(_zyGfifo__gfdL519_16_P0_m2_cbid[0]), .A1(_zyGfifo__gfdL522_15_P0_m2_cbid[0]), .Z(n3073));
Q_MX02 U2910 ( .S(n3553), .A0(tdata_ob[63]), .A1(n1972), .Z(n3072));
Q_MX02 U2911 ( .S(n3553), .A0(tdata_ob[62]), .A1(n1971), .Z(n3071));
Q_MX02 U2912 ( .S(n3553), .A0(tdata_ob[61]), .A1(n1970), .Z(n3070));
Q_MX02 U2913 ( .S(n3553), .A0(tdata_ob[60]), .A1(n1969), .Z(n3069));
Q_MX02 U2914 ( .S(n3553), .A0(tdata_ob[59]), .A1(n1968), .Z(n3068));
Q_MX02 U2915 ( .S(n3553), .A0(tdata_ob[58]), .A1(n1967), .Z(n3067));
Q_MX02 U2916 ( .S(n3553), .A0(tdata_ob[57]), .A1(n1966), .Z(n3066));
Q_MX02 U2917 ( .S(n3553), .A0(tdata_ob[56]), .A1(n1965), .Z(n3065));
Q_MX02 U2918 ( .S(n3553), .A0(tdata_ob[55]), .A1(n1964), .Z(n3064));
Q_MX02 U2919 ( .S(n3553), .A0(tdata_ob[54]), .A1(n1963), .Z(n3063));
Q_MX02 U2920 ( .S(n3553), .A0(tdata_ob[53]), .A1(n1962), .Z(n3062));
Q_MX02 U2921 ( .S(n3553), .A0(tdata_ob[52]), .A1(n1961), .Z(n3061));
Q_MX02 U2922 ( .S(n3553), .A0(tdata_ob[51]), .A1(n1960), .Z(n3060));
Q_MX02 U2923 ( .S(n3553), .A0(tdata_ob[50]), .A1(n1959), .Z(n3059));
Q_MX02 U2924 ( .S(n3553), .A0(tdata_ob[49]), .A1(n1958), .Z(n3058));
Q_MX02 U2925 ( .S(n3553), .A0(tdata_ob[48]), .A1(n1957), .Z(n3057));
Q_MX02 U2926 ( .S(n3553), .A0(tdata_ob[47]), .A1(n1956), .Z(n3056));
Q_MX02 U2927 ( .S(n3553), .A0(tdata_ob[46]), .A1(n1955), .Z(n3055));
Q_MX02 U2928 ( .S(n3553), .A0(tdata_ob[45]), .A1(n1954), .Z(n3054));
Q_MX02 U2929 ( .S(n3553), .A0(tdata_ob[44]), .A1(n1953), .Z(n3053));
Q_MX02 U2930 ( .S(n3553), .A0(tdata_ob[43]), .A1(n1952), .Z(n3052));
Q_MX02 U2931 ( .S(n3553), .A0(tdata_ob[42]), .A1(n1951), .Z(n3051));
Q_MX02 U2932 ( .S(n3553), .A0(tdata_ob[41]), .A1(n1950), .Z(n3050));
Q_MX02 U2933 ( .S(n3553), .A0(tdata_ob[40]), .A1(n1949), .Z(n3049));
Q_MX02 U2934 ( .S(n3553), .A0(tdata_ob[39]), .A1(n1948), .Z(n3048));
Q_MX02 U2935 ( .S(n3553), .A0(tdata_ob[38]), .A1(n1947), .Z(n3047));
Q_MX02 U2936 ( .S(n3553), .A0(tdata_ob[37]), .A1(n1946), .Z(n3046));
Q_MX02 U2937 ( .S(n3553), .A0(tdata_ob[36]), .A1(n1945), .Z(n3045));
Q_MX02 U2938 ( .S(n3553), .A0(tdata_ob[35]), .A1(n1944), .Z(n3044));
Q_MX02 U2939 ( .S(n3553), .A0(tdata_ob[34]), .A1(n1943), .Z(n3043));
Q_MX02 U2940 ( .S(n3553), .A0(tdata_ob[33]), .A1(n1942), .Z(n3042));
Q_MX02 U2941 ( .S(n3553), .A0(tdata_ob[32]), .A1(n1941), .Z(n3041));
Q_MX02 U2942 ( .S(n3553), .A0(tdata_ob[31]), .A1(n1940), .Z(n3040));
Q_MX02 U2943 ( .S(n3553), .A0(tdata_ob[30]), .A1(n1939), .Z(n3039));
Q_MX02 U2944 ( .S(n3553), .A0(tdata_ob[29]), .A1(n1938), .Z(n3038));
Q_MX02 U2945 ( .S(n3553), .A0(tdata_ob[28]), .A1(n1937), .Z(n3037));
Q_MX02 U2946 ( .S(n3553), .A0(tdata_ob[27]), .A1(n1936), .Z(n3036));
Q_MX02 U2947 ( .S(n3553), .A0(tdata_ob[26]), .A1(n1935), .Z(n3035));
Q_MX02 U2948 ( .S(n3553), .A0(tdata_ob[25]), .A1(n1934), .Z(n3034));
Q_MX02 U2949 ( .S(n3553), .A0(tdata_ob[24]), .A1(n1933), .Z(n3033));
Q_MX02 U2950 ( .S(n3553), .A0(tdata_ob[23]), .A1(n1932), .Z(n3032));
Q_MX02 U2951 ( .S(n3553), .A0(tdata_ob[22]), .A1(n1931), .Z(n3031));
Q_MX02 U2952 ( .S(n3553), .A0(tdata_ob[21]), .A1(n1930), .Z(n3030));
Q_MX02 U2953 ( .S(n3553), .A0(tdata_ob[20]), .A1(n1929), .Z(n3029));
Q_MX02 U2954 ( .S(n3553), .A0(tdata_ob[19]), .A1(n1928), .Z(n3028));
Q_MX02 U2955 ( .S(n3553), .A0(tdata_ob[18]), .A1(n1927), .Z(n3027));
Q_MX02 U2956 ( .S(n3553), .A0(tdata_ob[17]), .A1(n1926), .Z(n3026));
Q_MX02 U2957 ( .S(n3553), .A0(tdata_ob[16]), .A1(n1925), .Z(n3025));
Q_MX02 U2958 ( .S(n3553), .A0(tdata_ob[15]), .A1(n1924), .Z(n3024));
Q_MX02 U2959 ( .S(n3553), .A0(tdata_ob[14]), .A1(n1923), .Z(n3023));
Q_MX02 U2960 ( .S(n3553), .A0(tdata_ob[13]), .A1(n1922), .Z(n3022));
Q_MX02 U2961 ( .S(n3553), .A0(tdata_ob[12]), .A1(n1921), .Z(n3021));
Q_MX02 U2962 ( .S(n3553), .A0(tdata_ob[11]), .A1(n1920), .Z(n3020));
Q_MX02 U2963 ( .S(n3553), .A0(tdata_ob[10]), .A1(n1919), .Z(n3019));
Q_MX02 U2964 ( .S(n3553), .A0(tdata_ob[9]), .A1(n1918), .Z(n3018));
Q_MX02 U2965 ( .S(n3553), .A0(tdata_ob[8]), .A1(n1917), .Z(n3017));
Q_MX02 U2966 ( .S(n3553), .A0(tdata_ob[7]), .A1(n1916), .Z(n3016));
Q_MX02 U2967 ( .S(n3553), .A0(tdata_ob[6]), .A1(n1915), .Z(n3015));
Q_MX02 U2968 ( .S(n3553), .A0(tdata_ob[5]), .A1(n1914), .Z(n3014));
Q_MX02 U2969 ( .S(n3553), .A0(tdata_ob[4]), .A1(n1913), .Z(n3013));
Q_MX02 U2970 ( .S(n3553), .A0(tdata_ob[3]), .A1(n1912), .Z(n3012));
Q_MX02 U2971 ( .S(n3553), .A0(tdata_ob[2]), .A1(n1911), .Z(n3011));
Q_MX02 U2972 ( .S(n3553), .A0(tdata_ob[1]), .A1(n1910), .Z(n3010));
Q_MX02 U2973 ( .S(n3553), .A0(tdata_ob[0]), .A1(n1909), .Z(n3009));
Q_MX02 U2974 ( .S(_zyL439_meState8[0]), .A0(n2138), .A1(tstrb_ob[7]), .Z(n3008));
Q_MX02 U2975 ( .S(_zyL439_meState8[0]), .A0(n2137), .A1(tstrb_ob[6]), .Z(n3007));
Q_MX02 U2976 ( .S(_zyL439_meState8[0]), .A0(n2136), .A1(tstrb_ob[5]), .Z(n3006));
Q_MX02 U2977 ( .S(_zyL439_meState8[0]), .A0(n2135), .A1(tstrb_ob[4]), .Z(n3005));
Q_MX02 U2978 ( .S(_zyL439_meState8[0]), .A0(n2134), .A1(tstrb_ob[3]), .Z(n3004));
Q_MX02 U2979 ( .S(_zyL439_meState8[0]), .A0(n2133), .A1(tstrb_ob[2]), .Z(n3003));
Q_MX02 U2980 ( .S(_zyL439_meState8[0]), .A0(n2132), .A1(tstrb_ob[1]), .Z(n3002));
Q_MX02 U2981 ( .S(_zyL439_meState8[0]), .A0(n2131), .A1(tstrb_ob[0]), .Z(n3001));
Q_MX02 U2982 ( .S(n3550), .A0(n2999), .A1(n3567), .Z(n3000));
Q_XOR2 U2983 ( .A0(n2997), .A1(n2937), .Z(n2998));
Q_AD01HF U2984 ( .A0(n2995), .B0(n2936), .S(n2996), .CO(n2997));
Q_AD01HF U2985 ( .A0(n2993), .B0(n2935), .S(n2994), .CO(n2995));
Q_AD01HF U2986 ( .A0(n2991), .B0(n2934), .S(n2992), .CO(n2993));
Q_AD01HF U2987 ( .A0(n2989), .B0(n2933), .S(n2990), .CO(n2991));
Q_AD01HF U2988 ( .A0(n2987), .B0(n2932), .S(n2988), .CO(n2989));
Q_AD01HF U2989 ( .A0(n2985), .B0(n2931), .S(n2986), .CO(n2987));
Q_AD01HF U2990 ( .A0(n2983), .B0(n2930), .S(n2984), .CO(n2985));
Q_AD01HF U2991 ( .A0(n2981), .B0(n2929), .S(n2982), .CO(n2983));
Q_AD01HF U2992 ( .A0(n2979), .B0(n2928), .S(n2980), .CO(n2981));
Q_AD01HF U2993 ( .A0(n2977), .B0(n2927), .S(n2978), .CO(n2979));
Q_AD01HF U2994 ( .A0(n2975), .B0(n2926), .S(n2976), .CO(n2977));
Q_AD01HF U2995 ( .A0(n2973), .B0(n2925), .S(n2974), .CO(n2975));
Q_AD01HF U2996 ( .A0(n2971), .B0(n2924), .S(n2972), .CO(n2973));
Q_AD01HF U2997 ( .A0(n2969), .B0(n2923), .S(n2970), .CO(n2971));
Q_AD01HF U2998 ( .A0(n2967), .B0(n2922), .S(n2968), .CO(n2969));
Q_AD01HF U2999 ( .A0(n2965), .B0(n2921), .S(n2966), .CO(n2967));
Q_AD01HF U3000 ( .A0(n2963), .B0(n2920), .S(n2964), .CO(n2965));
Q_AD01HF U3001 ( .A0(n2961), .B0(n2919), .S(n2962), .CO(n2963));
Q_AD01HF U3002 ( .A0(n2959), .B0(n2918), .S(n2960), .CO(n2961));
Q_AD01HF U3003 ( .A0(n2957), .B0(n2917), .S(n2958), .CO(n2959));
Q_AD01HF U3004 ( .A0(n2955), .B0(n2916), .S(n2956), .CO(n2957));
Q_AD01HF U3005 ( .A0(n2953), .B0(n2915), .S(n2954), .CO(n2955));
Q_AD01HF U3006 ( .A0(n2951), .B0(n2914), .S(n2952), .CO(n2953));
Q_AD01HF U3007 ( .A0(n2949), .B0(n2913), .S(n2950), .CO(n2951));
Q_AD01HF U3008 ( .A0(n2947), .B0(n2912), .S(n2948), .CO(n2949));
Q_AD01HF U3009 ( .A0(n2945), .B0(n2911), .S(n2946), .CO(n2947));
Q_AD01HF U3010 ( .A0(n2943), .B0(n2910), .S(n2944), .CO(n2945));
Q_AD01HF U3011 ( .A0(n2941), .B0(n2909), .S(n2942), .CO(n2943));
Q_AD01HF U3012 ( .A0(n2939), .B0(n2908), .S(n2940), .CO(n2941));
Q_AD01HF U3013 ( .A0(n2906), .B0(n2907), .S(n2938), .CO(n2939));
Q_MX02 U3014 ( .S(n1897), .A0(n2904), .A1(n2844), .Z(n2936));
Q_MX02 U3015 ( .S(n1897), .A0(n2902), .A1(n2843), .Z(n2935));
Q_MX02 U3016 ( .S(n1897), .A0(n2900), .A1(n2842), .Z(n2934));
Q_MX02 U3017 ( .S(n1897), .A0(n2898), .A1(n2841), .Z(n2933));
Q_MX02 U3018 ( .S(n1897), .A0(n2896), .A1(n2840), .Z(n2932));
Q_MX02 U3019 ( .S(n1897), .A0(n2894), .A1(n2839), .Z(n2931));
Q_MX02 U3020 ( .S(n1897), .A0(n2892), .A1(n2838), .Z(n2930));
Q_MX02 U3021 ( .S(n1897), .A0(n2890), .A1(n2837), .Z(n2929));
Q_MX02 U3022 ( .S(n1897), .A0(n2888), .A1(n2836), .Z(n2928));
Q_MX02 U3023 ( .S(n1897), .A0(n2886), .A1(n2835), .Z(n2927));
Q_MX02 U3024 ( .S(n1897), .A0(n2884), .A1(n2834), .Z(n2926));
Q_MX02 U3025 ( .S(n1897), .A0(n2882), .A1(n2833), .Z(n2925));
Q_MX02 U3026 ( .S(n1897), .A0(n2880), .A1(n2832), .Z(n2924));
Q_MX02 U3027 ( .S(n1897), .A0(n2878), .A1(n2831), .Z(n2923));
Q_MX02 U3028 ( .S(n1897), .A0(n2876), .A1(n2830), .Z(n2922));
Q_MX02 U3029 ( .S(n1897), .A0(n2874), .A1(n2829), .Z(n2921));
Q_MX02 U3030 ( .S(n1897), .A0(n2872), .A1(n2828), .Z(n2920));
Q_MX02 U3031 ( .S(n1897), .A0(n2870), .A1(n2827), .Z(n2919));
Q_MX02 U3032 ( .S(n1897), .A0(n2868), .A1(n2826), .Z(n2918));
Q_MX02 U3033 ( .S(n1897), .A0(n2866), .A1(n2825), .Z(n2917));
Q_MX02 U3034 ( .S(n1897), .A0(n2864), .A1(n2824), .Z(n2916));
Q_MX02 U3035 ( .S(n1897), .A0(n2862), .A1(n2823), .Z(n2915));
Q_MX02 U3036 ( .S(n1897), .A0(n2860), .A1(n2822), .Z(n2914));
Q_MX02 U3037 ( .S(n1897), .A0(n2858), .A1(n2821), .Z(n2913));
Q_MX02 U3038 ( .S(n1897), .A0(n2856), .A1(n2820), .Z(n2912));
Q_MX02 U3039 ( .S(n1897), .A0(n2854), .A1(n2819), .Z(n2911));
Q_MX02 U3040 ( .S(n1897), .A0(n2852), .A1(n2818), .Z(n2910));
Q_MX02 U3041 ( .S(n1897), .A0(n2850), .A1(n2817), .Z(n2909));
Q_MX02 U3042 ( .S(n1897), .A0(n2848), .A1(n2816), .Z(n2908));
Q_MX02 U3043 ( .S(n1897), .A0(n2846), .A1(n2815), .Z(n2907));
Q_XOR2 U3044 ( .A0(n3549), .A1(n2814), .Z(n2906));
Q_XOR2 U3045 ( .A0(n5878), .A1(n2845), .Z(n2937));
Q_AD01HF U3046 ( .A0(n2903), .B0(n2844), .S(n2904), .CO(n2905));
Q_AD01HF U3047 ( .A0(n2901), .B0(n2843), .S(n2902), .CO(n2903));
Q_AD01HF U3048 ( .A0(n2899), .B0(n2842), .S(n2900), .CO(n2901));
Q_AD01HF U3049 ( .A0(n2897), .B0(n2841), .S(n2898), .CO(n2899));
Q_AD01HF U3050 ( .A0(n2895), .B0(n2840), .S(n2896), .CO(n2897));
Q_AD01HF U3051 ( .A0(n2893), .B0(n2839), .S(n2894), .CO(n2895));
Q_AD01HF U3052 ( .A0(n2891), .B0(n2838), .S(n2892), .CO(n2893));
Q_AD01HF U3053 ( .A0(n2889), .B0(n2837), .S(n2890), .CO(n2891));
Q_AD01HF U3054 ( .A0(n2887), .B0(n2836), .S(n2888), .CO(n2889));
Q_AD01HF U3055 ( .A0(n2885), .B0(n2835), .S(n2886), .CO(n2887));
Q_AD01HF U3056 ( .A0(n2883), .B0(n2834), .S(n2884), .CO(n2885));
Q_AD01HF U3057 ( .A0(n2881), .B0(n2833), .S(n2882), .CO(n2883));
Q_AD01HF U3058 ( .A0(n2879), .B0(n2832), .S(n2880), .CO(n2881));
Q_AD01HF U3059 ( .A0(n2877), .B0(n2831), .S(n2878), .CO(n2879));
Q_AD01HF U3060 ( .A0(n2875), .B0(n2830), .S(n2876), .CO(n2877));
Q_AD01HF U3061 ( .A0(n2873), .B0(n2829), .S(n2874), .CO(n2875));
Q_AD01HF U3062 ( .A0(n2871), .B0(n2828), .S(n2872), .CO(n2873));
Q_AD01HF U3063 ( .A0(n2869), .B0(n2827), .S(n2870), .CO(n2871));
Q_AD01HF U3064 ( .A0(n2867), .B0(n2826), .S(n2868), .CO(n2869));
Q_AD01HF U3065 ( .A0(n2865), .B0(n2825), .S(n2866), .CO(n2867));
Q_AD01HF U3066 ( .A0(n2863), .B0(n2824), .S(n2864), .CO(n2865));
Q_AD01HF U3067 ( .A0(n2861), .B0(n2823), .S(n2862), .CO(n2863));
Q_AD01HF U3068 ( .A0(n2859), .B0(n2822), .S(n2860), .CO(n2861));
Q_AD01HF U3069 ( .A0(n2857), .B0(n2821), .S(n2858), .CO(n2859));
Q_AD01HF U3070 ( .A0(n2855), .B0(n2820), .S(n2856), .CO(n2857));
Q_AD01HF U3071 ( .A0(n2853), .B0(n2819), .S(n2854), .CO(n2855));
Q_AD01HF U3072 ( .A0(n2851), .B0(n2818), .S(n2852), .CO(n2853));
Q_AD01HF U3073 ( .A0(n2849), .B0(n2817), .S(n2850), .CO(n2851));
Q_AD01HF U3074 ( .A0(n2847), .B0(n2816), .S(n2848), .CO(n2849));
Q_AD01HF U3075 ( .A0(n2814), .B0(n2815), .S(n2846), .CO(n2847));
Q_MX02 U3076 ( .S(n3548), .A0(n2719), .A1(n2813), .Z(n2845));
Q_MX02 U3077 ( .S(n3548), .A0(n2718), .A1(n2811), .Z(n2844));
Q_MX02 U3078 ( .S(n3548), .A0(n2717), .A1(n2809), .Z(n2843));
Q_MX02 U3079 ( .S(n3548), .A0(n2716), .A1(n2807), .Z(n2842));
Q_MX02 U3080 ( .S(n3548), .A0(n2715), .A1(n2805), .Z(n2841));
Q_MX02 U3081 ( .S(n3548), .A0(n2714), .A1(n2803), .Z(n2840));
Q_MX02 U3082 ( .S(n3548), .A0(n2713), .A1(n2801), .Z(n2839));
Q_MX02 U3083 ( .S(n3548), .A0(n2712), .A1(n2799), .Z(n2838));
Q_MX02 U3084 ( .S(n3548), .A0(n2711), .A1(n2797), .Z(n2837));
Q_MX02 U3085 ( .S(n3548), .A0(n2710), .A1(n2795), .Z(n2836));
Q_MX02 U3086 ( .S(n3548), .A0(n2709), .A1(n2793), .Z(n2835));
Q_MX02 U3087 ( .S(n3548), .A0(n2708), .A1(n2791), .Z(n2834));
Q_MX02 U3088 ( .S(n3548), .A0(n2707), .A1(n2789), .Z(n2833));
Q_MX02 U3089 ( .S(n3548), .A0(n2706), .A1(n2787), .Z(n2832));
Q_MX02 U3090 ( .S(n3548), .A0(n2705), .A1(n2785), .Z(n2831));
Q_MX02 U3091 ( .S(n3548), .A0(n2704), .A1(n2783), .Z(n2830));
Q_MX02 U3092 ( .S(n3548), .A0(n2703), .A1(n2781), .Z(n2829));
Q_MX02 U3093 ( .S(n3548), .A0(n2702), .A1(n2779), .Z(n2828));
Q_MX02 U3094 ( .S(n3548), .A0(n2701), .A1(n2777), .Z(n2827));
Q_MX02 U3095 ( .S(n3548), .A0(n2700), .A1(n2775), .Z(n2826));
Q_MX02 U3096 ( .S(n3548), .A0(n2699), .A1(n2773), .Z(n2825));
Q_MX02 U3097 ( .S(n3548), .A0(n2698), .A1(n2771), .Z(n2824));
Q_MX02 U3098 ( .S(n3548), .A0(n2697), .A1(n2769), .Z(n2823));
Q_MX02 U3099 ( .S(n3548), .A0(n2696), .A1(n2767), .Z(n2822));
Q_MX02 U3100 ( .S(n3548), .A0(n2695), .A1(n2765), .Z(n2821));
Q_MX02 U3101 ( .S(n3548), .A0(n2694), .A1(n2763), .Z(n2820));
Q_MX02 U3102 ( .S(n3548), .A0(n2693), .A1(n2761), .Z(n2819));
Q_MX02 U3103 ( .S(n3548), .A0(n2692), .A1(n2759), .Z(n2818));
Q_MX02 U3104 ( .S(n3548), .A0(n2691), .A1(n2757), .Z(n2817));
Q_MX02 U3105 ( .S(n3548), .A0(n2690), .A1(n2755), .Z(n2816));
Q_MX02 U3106 ( .S(n3548), .A0(n2689), .A1(n2753), .Z(n2815));
Q_MX02 U3107 ( .S(n3548), .A0(n2688), .A1(n2752), .Z(n2814));
Q_XOR2 U3108 ( .A0(n2812), .A1(n2751), .Z(n2813));
Q_AD01HF U3109 ( .A0(n2810), .B0(n2750), .S(n2811), .CO(n2812));
Q_AD01HF U3110 ( .A0(n2808), .B0(n2749), .S(n2809), .CO(n2810));
Q_AD01HF U3111 ( .A0(n2806), .B0(n2748), .S(n2807), .CO(n2808));
Q_AD01HF U3112 ( .A0(n2804), .B0(n2747), .S(n2805), .CO(n2806));
Q_AD01HF U3113 ( .A0(n2802), .B0(n2746), .S(n2803), .CO(n2804));
Q_AD01HF U3114 ( .A0(n2800), .B0(n2745), .S(n2801), .CO(n2802));
Q_AD01HF U3115 ( .A0(n2798), .B0(n2744), .S(n2799), .CO(n2800));
Q_AD01HF U3116 ( .A0(n2796), .B0(n2743), .S(n2797), .CO(n2798));
Q_AD01HF U3117 ( .A0(n2794), .B0(n2742), .S(n2795), .CO(n2796));
Q_AD01HF U3118 ( .A0(n2792), .B0(n2741), .S(n2793), .CO(n2794));
Q_AD01HF U3119 ( .A0(n2790), .B0(n2740), .S(n2791), .CO(n2792));
Q_AD01HF U3120 ( .A0(n2788), .B0(n2739), .S(n2789), .CO(n2790));
Q_AD01HF U3121 ( .A0(n2786), .B0(n2738), .S(n2787), .CO(n2788));
Q_AD01HF U3122 ( .A0(n2784), .B0(n2737), .S(n2785), .CO(n2786));
Q_AD01HF U3123 ( .A0(n2782), .B0(n2736), .S(n2783), .CO(n2784));
Q_AD01HF U3124 ( .A0(n2780), .B0(n2735), .S(n2781), .CO(n2782));
Q_AD01HF U3125 ( .A0(n2778), .B0(n2734), .S(n2779), .CO(n2780));
Q_AD01HF U3126 ( .A0(n2776), .B0(n2733), .S(n2777), .CO(n2778));
Q_AD01HF U3127 ( .A0(n2774), .B0(n2732), .S(n2775), .CO(n2776));
Q_AD01HF U3128 ( .A0(n2772), .B0(n2731), .S(n2773), .CO(n2774));
Q_AD01HF U3129 ( .A0(n2770), .B0(n2730), .S(n2771), .CO(n2772));
Q_AD01HF U3130 ( .A0(n2768), .B0(n2729), .S(n2769), .CO(n2770));
Q_AD01HF U3131 ( .A0(n2766), .B0(n2728), .S(n2767), .CO(n2768));
Q_AD01HF U3132 ( .A0(n2764), .B0(n2727), .S(n2765), .CO(n2766));
Q_AD01HF U3133 ( .A0(n2762), .B0(n2726), .S(n2763), .CO(n2764));
Q_AD01HF U3134 ( .A0(n2760), .B0(n2725), .S(n2761), .CO(n2762));
Q_AD01HF U3135 ( .A0(n2758), .B0(n2724), .S(n2759), .CO(n2760));
Q_AD01HF U3136 ( .A0(n2756), .B0(n2723), .S(n2757), .CO(n2758));
Q_AD01HF U3137 ( .A0(n2754), .B0(n2722), .S(n2755), .CO(n2756));
Q_AD01HF U3138 ( .A0(n2720), .B0(n2721), .S(n2753), .CO(n2754));
Q_INV U3139 ( .A(n2720), .Z(n2752));
Q_MX02 U3140 ( .S(_zyL439_meState8[0]), .A0(n2687), .A1(n2719), .Z(n2751));
Q_MX02 U3141 ( .S(_zyL439_meState8[0]), .A0(n2686), .A1(n2718), .Z(n2750));
Q_MX02 U3142 ( .S(_zyL439_meState8[0]), .A0(n2685), .A1(n2717), .Z(n2749));
Q_MX02 U3143 ( .S(_zyL439_meState8[0]), .A0(n2684), .A1(n2716), .Z(n2748));
Q_MX02 U3144 ( .S(_zyL439_meState8[0]), .A0(n2683), .A1(n2715), .Z(n2747));
Q_MX02 U3145 ( .S(_zyL439_meState8[0]), .A0(n2682), .A1(n2714), .Z(n2746));
Q_MX02 U3146 ( .S(_zyL439_meState8[0]), .A0(n2681), .A1(n2713), .Z(n2745));
Q_MX02 U3147 ( .S(_zyL439_meState8[0]), .A0(n2680), .A1(n2712), .Z(n2744));
Q_MX02 U3148 ( .S(_zyL439_meState8[0]), .A0(n2679), .A1(n2711), .Z(n2743));
Q_MX02 U3149 ( .S(_zyL439_meState8[0]), .A0(n2678), .A1(n2710), .Z(n2742));
Q_MX02 U3150 ( .S(_zyL439_meState8[0]), .A0(n2677), .A1(n2709), .Z(n2741));
Q_MX02 U3151 ( .S(_zyL439_meState8[0]), .A0(n2676), .A1(n2708), .Z(n2740));
Q_MX02 U3152 ( .S(_zyL439_meState8[0]), .A0(n2675), .A1(n2707), .Z(n2739));
Q_MX02 U3153 ( .S(_zyL439_meState8[0]), .A0(n2674), .A1(n2706), .Z(n2738));
Q_MX02 U3154 ( .S(_zyL439_meState8[0]), .A0(n2673), .A1(n2705), .Z(n2737));
Q_MX02 U3155 ( .S(_zyL439_meState8[0]), .A0(n2672), .A1(n2704), .Z(n2736));
Q_MX02 U3156 ( .S(_zyL439_meState8[0]), .A0(n2671), .A1(n2703), .Z(n2735));
Q_MX02 U3157 ( .S(_zyL439_meState8[0]), .A0(n2670), .A1(n2702), .Z(n2734));
Q_MX02 U3158 ( .S(_zyL439_meState8[0]), .A0(n2669), .A1(n2701), .Z(n2733));
Q_MX02 U3159 ( .S(_zyL439_meState8[0]), .A0(n2668), .A1(n2700), .Z(n2732));
Q_MX02 U3160 ( .S(_zyL439_meState8[0]), .A0(n2667), .A1(n2699), .Z(n2731));
Q_MX02 U3161 ( .S(_zyL439_meState8[0]), .A0(n2666), .A1(n2698), .Z(n2730));
Q_MX02 U3162 ( .S(_zyL439_meState8[0]), .A0(n2665), .A1(n2697), .Z(n2729));
Q_MX02 U3163 ( .S(_zyL439_meState8[0]), .A0(n2664), .A1(n2696), .Z(n2728));
Q_MX02 U3164 ( .S(_zyL439_meState8[0]), .A0(n2663), .A1(n2695), .Z(n2727));
Q_MX02 U3165 ( .S(_zyL439_meState8[0]), .A0(n2662), .A1(n2694), .Z(n2726));
Q_MX02 U3166 ( .S(_zyL439_meState8[0]), .A0(n2661), .A1(n2693), .Z(n2725));
Q_MX02 U3167 ( .S(_zyL439_meState8[0]), .A0(n2660), .A1(n2692), .Z(n2724));
Q_MX02 U3168 ( .S(_zyL439_meState8[0]), .A0(n2659), .A1(n2691), .Z(n2723));
Q_MX02 U3169 ( .S(_zyL439_meState8[0]), .A0(n2658), .A1(n2690), .Z(n2722));
Q_MX02 U3170 ( .S(_zyL439_meState8[0]), .A0(n2657), .A1(n2689), .Z(n2721));
Q_MX02 U3171 ( .S(_zyL439_meState8[0]), .A0(n2656), .A1(n2688), .Z(n2720));
Q_MX02 U3172 ( .S(n3547), .A0(n2529), .A1(n2655), .Z(n2719));
Q_MX02 U3173 ( .S(n3547), .A0(n2527), .A1(n2653), .Z(n2718));
Q_MX02 U3174 ( .S(n3547), .A0(n2525), .A1(n2651), .Z(n2717));
Q_MX02 U3175 ( .S(n3547), .A0(n2523), .A1(n2649), .Z(n2716));
Q_MX02 U3176 ( .S(n3547), .A0(n2521), .A1(n2647), .Z(n2715));
Q_MX02 U3177 ( .S(n3547), .A0(n2519), .A1(n2645), .Z(n2714));
Q_MX02 U3178 ( .S(n3547), .A0(n2517), .A1(n2643), .Z(n2713));
Q_MX02 U3179 ( .S(n3547), .A0(n2515), .A1(n2641), .Z(n2712));
Q_MX02 U3180 ( .S(n3547), .A0(n2513), .A1(n2639), .Z(n2711));
Q_MX02 U3181 ( .S(n3547), .A0(n2511), .A1(n2637), .Z(n2710));
Q_MX02 U3182 ( .S(n3547), .A0(n2509), .A1(n2635), .Z(n2709));
Q_MX02 U3183 ( .S(n3547), .A0(n2507), .A1(n2633), .Z(n2708));
Q_MX02 U3184 ( .S(n3547), .A0(n2505), .A1(n2631), .Z(n2707));
Q_MX02 U3185 ( .S(n3547), .A0(n2503), .A1(n2629), .Z(n2706));
Q_MX02 U3186 ( .S(n3547), .A0(n2501), .A1(n2627), .Z(n2705));
Q_MX02 U3187 ( .S(n3547), .A0(n2499), .A1(n2625), .Z(n2704));
Q_MX02 U3188 ( .S(n3547), .A0(n2497), .A1(n2623), .Z(n2703));
Q_MX02 U3189 ( .S(n3547), .A0(n2495), .A1(n2621), .Z(n2702));
Q_MX02 U3190 ( .S(n3547), .A0(n2493), .A1(n2619), .Z(n2701));
Q_MX02 U3191 ( .S(n3547), .A0(n2491), .A1(n2617), .Z(n2700));
Q_MX02 U3192 ( .S(n3547), .A0(n2489), .A1(n2615), .Z(n2699));
Q_MX02 U3193 ( .S(n3547), .A0(n2487), .A1(n2613), .Z(n2698));
Q_MX02 U3194 ( .S(n3547), .A0(n2485), .A1(n2611), .Z(n2697));
Q_MX02 U3195 ( .S(n3547), .A0(n2483), .A1(n2609), .Z(n2696));
Q_MX02 U3196 ( .S(n3547), .A0(n2481), .A1(n2607), .Z(n2695));
Q_MX02 U3197 ( .S(n3547), .A0(n2479), .A1(n2605), .Z(n2694));
Q_MX02 U3198 ( .S(n3547), .A0(n2477), .A1(n2603), .Z(n2693));
Q_MX02 U3199 ( .S(n3547), .A0(n2475), .A1(n2601), .Z(n2692));
Q_MX02 U3200 ( .S(n3547), .A0(n2473), .A1(n2599), .Z(n2691));
Q_MX02 U3201 ( .S(n3547), .A0(n2471), .A1(n2597), .Z(n2690));
Q_MX02 U3202 ( .S(n3547), .A0(n2469), .A1(n2595), .Z(n2689));
Q_MX02 U3203 ( .S(n3547), .A0(n2467), .A1(n2594), .Z(n2688));
Q_MX02 U3204 ( .S(n2150), .A0(n2655), .A1(n2561), .Z(n2687));
Q_MX02 U3205 ( .S(n2150), .A0(n2653), .A1(n2560), .Z(n2686));
Q_MX02 U3206 ( .S(n2150), .A0(n2651), .A1(n2559), .Z(n2685));
Q_MX02 U3207 ( .S(n2150), .A0(n2649), .A1(n2558), .Z(n2684));
Q_MX02 U3208 ( .S(n2150), .A0(n2647), .A1(n2557), .Z(n2683));
Q_MX02 U3209 ( .S(n2150), .A0(n2645), .A1(n2556), .Z(n2682));
Q_MX02 U3210 ( .S(n2150), .A0(n2643), .A1(n2555), .Z(n2681));
Q_MX02 U3211 ( .S(n2150), .A0(n2641), .A1(n2554), .Z(n2680));
Q_MX02 U3212 ( .S(n2150), .A0(n2639), .A1(n2553), .Z(n2679));
Q_MX02 U3213 ( .S(n2150), .A0(n2637), .A1(n2552), .Z(n2678));
Q_MX02 U3214 ( .S(n2150), .A0(n2635), .A1(n2551), .Z(n2677));
Q_MX02 U3215 ( .S(n2150), .A0(n2633), .A1(n2550), .Z(n2676));
Q_MX02 U3216 ( .S(n2150), .A0(n2631), .A1(n2549), .Z(n2675));
Q_MX02 U3217 ( .S(n2150), .A0(n2629), .A1(n2548), .Z(n2674));
Q_MX02 U3218 ( .S(n2150), .A0(n2627), .A1(n2547), .Z(n2673));
Q_MX02 U3219 ( .S(n2150), .A0(n2625), .A1(n2546), .Z(n2672));
Q_MX02 U3220 ( .S(n2150), .A0(n2623), .A1(n2545), .Z(n2671));
Q_MX02 U3221 ( .S(n2150), .A0(n2621), .A1(n2544), .Z(n2670));
Q_MX02 U3222 ( .S(n2150), .A0(n2619), .A1(n2543), .Z(n2669));
Q_MX02 U3223 ( .S(n2150), .A0(n2617), .A1(n2542), .Z(n2668));
Q_MX02 U3224 ( .S(n2150), .A0(n2615), .A1(n2541), .Z(n2667));
Q_MX02 U3225 ( .S(n2150), .A0(n2613), .A1(n2540), .Z(n2666));
Q_MX02 U3226 ( .S(n2150), .A0(n2611), .A1(n2539), .Z(n2665));
Q_MX02 U3227 ( .S(n2150), .A0(n2609), .A1(n2538), .Z(n2664));
Q_MX02 U3228 ( .S(n2150), .A0(n2607), .A1(n2537), .Z(n2663));
Q_MX02 U3229 ( .S(n2150), .A0(n2605), .A1(n2536), .Z(n2662));
Q_MX02 U3230 ( .S(n2150), .A0(n2603), .A1(n2535), .Z(n2661));
Q_MX02 U3231 ( .S(n2150), .A0(n2601), .A1(n2534), .Z(n2660));
Q_MX02 U3232 ( .S(n2150), .A0(n2599), .A1(n2533), .Z(n2659));
Q_MX02 U3233 ( .S(n2150), .A0(n2597), .A1(n2532), .Z(n2658));
Q_MX02 U3234 ( .S(n2150), .A0(n2595), .A1(n2531), .Z(n2657));
Q_MX02 U3235 ( .S(n2150), .A0(n2594), .A1(n2530), .Z(n2656));
Q_XOR2 U3236 ( .A0(n2654), .A1(n2593), .Z(n2655));
Q_AD01HF U3237 ( .A0(n2652), .B0(n2592), .S(n2653), .CO(n2654));
Q_AD01HF U3238 ( .A0(n2650), .B0(n2591), .S(n2651), .CO(n2652));
Q_AD01HF U3239 ( .A0(n2648), .B0(n2590), .S(n2649), .CO(n2650));
Q_AD01HF U3240 ( .A0(n2646), .B0(n2589), .S(n2647), .CO(n2648));
Q_AD01HF U3241 ( .A0(n2644), .B0(n2588), .S(n2645), .CO(n2646));
Q_AD01HF U3242 ( .A0(n2642), .B0(n2587), .S(n2643), .CO(n2644));
Q_AD01HF U3243 ( .A0(n2640), .B0(n2586), .S(n2641), .CO(n2642));
Q_AD01HF U3244 ( .A0(n2638), .B0(n2585), .S(n2639), .CO(n2640));
Q_AD01HF U3245 ( .A0(n2636), .B0(n2584), .S(n2637), .CO(n2638));
Q_AD01HF U3246 ( .A0(n2634), .B0(n2583), .S(n2635), .CO(n2636));
Q_AD01HF U3247 ( .A0(n2632), .B0(n2582), .S(n2633), .CO(n2634));
Q_AD01HF U3248 ( .A0(n2630), .B0(n2581), .S(n2631), .CO(n2632));
Q_AD01HF U3249 ( .A0(n2628), .B0(n2580), .S(n2629), .CO(n2630));
Q_AD01HF U3250 ( .A0(n2626), .B0(n2579), .S(n2627), .CO(n2628));
Q_AD01HF U3251 ( .A0(n2624), .B0(n2578), .S(n2625), .CO(n2626));
Q_AD01HF U3252 ( .A0(n2622), .B0(n2577), .S(n2623), .CO(n2624));
Q_AD01HF U3253 ( .A0(n2620), .B0(n2576), .S(n2621), .CO(n2622));
Q_AD01HF U3254 ( .A0(n2618), .B0(n2575), .S(n2619), .CO(n2620));
Q_AD01HF U3255 ( .A0(n2616), .B0(n2574), .S(n2617), .CO(n2618));
Q_AD01HF U3256 ( .A0(n2614), .B0(n2573), .S(n2615), .CO(n2616));
Q_AD01HF U3257 ( .A0(n2612), .B0(n2572), .S(n2613), .CO(n2614));
Q_AD01HF U3258 ( .A0(n2610), .B0(n2571), .S(n2611), .CO(n2612));
Q_AD01HF U3259 ( .A0(n2608), .B0(n2570), .S(n2609), .CO(n2610));
Q_AD01HF U3260 ( .A0(n2606), .B0(n2569), .S(n2607), .CO(n2608));
Q_AD01HF U3261 ( .A0(n2604), .B0(n2568), .S(n2605), .CO(n2606));
Q_AD01HF U3262 ( .A0(n2602), .B0(n2567), .S(n2603), .CO(n2604));
Q_AD01HF U3263 ( .A0(n2600), .B0(n2566), .S(n2601), .CO(n2602));
Q_AD01HF U3264 ( .A0(n2598), .B0(n2565), .S(n2599), .CO(n2600));
Q_AD01HF U3265 ( .A0(n2596), .B0(n2564), .S(n2597), .CO(n2598));
Q_AD01HF U3266 ( .A0(n2563), .B0(n2562), .S(n2595), .CO(n2596));
Q_INV U3267 ( .A(n2562), .Z(n2594));
Q_MX02 U3268 ( .S(_zyL439_meState8[0]), .A0(n2561), .A1(n2529), .Z(n2593));
Q_MX02 U3269 ( .S(_zyL439_meState8[0]), .A0(n2560), .A1(n2527), .Z(n2592));
Q_MX02 U3270 ( .S(_zyL439_meState8[0]), .A0(n2559), .A1(n2525), .Z(n2591));
Q_MX02 U3271 ( .S(_zyL439_meState8[0]), .A0(n2558), .A1(n2523), .Z(n2590));
Q_MX02 U3272 ( .S(_zyL439_meState8[0]), .A0(n2557), .A1(n2521), .Z(n2589));
Q_MX02 U3273 ( .S(_zyL439_meState8[0]), .A0(n2556), .A1(n2519), .Z(n2588));
Q_MX02 U3274 ( .S(_zyL439_meState8[0]), .A0(n2555), .A1(n2517), .Z(n2587));
Q_MX02 U3275 ( .S(_zyL439_meState8[0]), .A0(n2554), .A1(n2515), .Z(n2586));
Q_MX02 U3276 ( .S(_zyL439_meState8[0]), .A0(n2553), .A1(n2513), .Z(n2585));
Q_MX02 U3277 ( .S(_zyL439_meState8[0]), .A0(n2552), .A1(n2511), .Z(n2584));
Q_MX02 U3278 ( .S(_zyL439_meState8[0]), .A0(n2551), .A1(n2509), .Z(n2583));
Q_MX02 U3279 ( .S(_zyL439_meState8[0]), .A0(n2550), .A1(n2507), .Z(n2582));
Q_MX02 U3280 ( .S(_zyL439_meState8[0]), .A0(n2549), .A1(n2505), .Z(n2581));
Q_MX02 U3281 ( .S(_zyL439_meState8[0]), .A0(n2548), .A1(n2503), .Z(n2580));
Q_MX02 U3282 ( .S(_zyL439_meState8[0]), .A0(n2547), .A1(n2501), .Z(n2579));
Q_MX02 U3283 ( .S(_zyL439_meState8[0]), .A0(n2546), .A1(n2499), .Z(n2578));
Q_MX02 U3284 ( .S(_zyL439_meState8[0]), .A0(n2545), .A1(n2497), .Z(n2577));
Q_MX02 U3285 ( .S(_zyL439_meState8[0]), .A0(n2544), .A1(n2495), .Z(n2576));
Q_MX02 U3286 ( .S(_zyL439_meState8[0]), .A0(n2543), .A1(n2493), .Z(n2575));
Q_MX02 U3287 ( .S(_zyL439_meState8[0]), .A0(n2542), .A1(n2491), .Z(n2574));
Q_MX02 U3288 ( .S(_zyL439_meState8[0]), .A0(n2541), .A1(n2489), .Z(n2573));
Q_MX02 U3289 ( .S(_zyL439_meState8[0]), .A0(n2540), .A1(n2487), .Z(n2572));
Q_MX02 U3290 ( .S(_zyL439_meState8[0]), .A0(n2539), .A1(n2485), .Z(n2571));
Q_MX02 U3291 ( .S(_zyL439_meState8[0]), .A0(n2538), .A1(n2483), .Z(n2570));
Q_MX02 U3292 ( .S(_zyL439_meState8[0]), .A0(n2537), .A1(n2481), .Z(n2569));
Q_MX02 U3293 ( .S(_zyL439_meState8[0]), .A0(n2536), .A1(n2479), .Z(n2568));
Q_MX02 U3294 ( .S(_zyL439_meState8[0]), .A0(n2535), .A1(n2477), .Z(n2567));
Q_MX02 U3295 ( .S(_zyL439_meState8[0]), .A0(n2534), .A1(n2475), .Z(n2566));
Q_MX02 U3296 ( .S(_zyL439_meState8[0]), .A0(n2533), .A1(n2473), .Z(n2565));
Q_MX02 U3297 ( .S(_zyL439_meState8[0]), .A0(n2532), .A1(n2471), .Z(n2564));
Q_MX02 U3298 ( .S(_zyL439_meState8[0]), .A0(n2531), .A1(n2469), .Z(n2563));
Q_MX02 U3299 ( .S(_zyL439_meState8[0]), .A0(n2530), .A1(n2467), .Z(n2562));
Q_MX02 U3300 ( .S(n3540), .A0(n2293), .A1(n2529), .Z(n2561));
Q_MX02 U3301 ( .S(n3540), .A0(n2292), .A1(n2527), .Z(n2560));
Q_MX02 U3302 ( .S(n3540), .A0(n2291), .A1(n2525), .Z(n2559));
Q_MX02 U3303 ( .S(n3540), .A0(n2290), .A1(n2523), .Z(n2558));
Q_MX02 U3304 ( .S(n3540), .A0(n2289), .A1(n2521), .Z(n2557));
Q_MX02 U3305 ( .S(n3540), .A0(n2288), .A1(n2519), .Z(n2556));
Q_MX02 U3306 ( .S(n3540), .A0(n2287), .A1(n2517), .Z(n2555));
Q_MX02 U3307 ( .S(n3540), .A0(n2286), .A1(n2515), .Z(n2554));
Q_MX02 U3308 ( .S(n3540), .A0(n2285), .A1(n2513), .Z(n2553));
Q_MX02 U3309 ( .S(n3540), .A0(n2284), .A1(n2511), .Z(n2552));
Q_MX02 U3310 ( .S(n3540), .A0(n2283), .A1(n2509), .Z(n2551));
Q_MX02 U3311 ( .S(n3540), .A0(n2282), .A1(n2507), .Z(n2550));
Q_MX02 U3312 ( .S(n3540), .A0(n2281), .A1(n2505), .Z(n2549));
Q_MX02 U3313 ( .S(n3540), .A0(n2280), .A1(n2503), .Z(n2548));
Q_MX02 U3314 ( .S(n3540), .A0(n2279), .A1(n2501), .Z(n2547));
Q_MX02 U3315 ( .S(n3540), .A0(n2278), .A1(n2499), .Z(n2546));
Q_MX02 U3316 ( .S(n3540), .A0(n2277), .A1(n2497), .Z(n2545));
Q_MX02 U3317 ( .S(n3540), .A0(n2276), .A1(n2495), .Z(n2544));
Q_MX02 U3318 ( .S(n3540), .A0(n2275), .A1(n2493), .Z(n2543));
Q_MX02 U3319 ( .S(n3540), .A0(n2274), .A1(n2491), .Z(n2542));
Q_MX02 U3320 ( .S(n3540), .A0(n2273), .A1(n2489), .Z(n2541));
Q_MX02 U3321 ( .S(n3540), .A0(n2272), .A1(n2487), .Z(n2540));
Q_MX02 U3322 ( .S(n3540), .A0(n2271), .A1(n2485), .Z(n2539));
Q_MX02 U3323 ( .S(n3540), .A0(n2270), .A1(n2483), .Z(n2538));
Q_MX02 U3324 ( .S(n3540), .A0(n2269), .A1(n2481), .Z(n2537));
Q_MX02 U3325 ( .S(n3540), .A0(n2268), .A1(n2479), .Z(n2536));
Q_MX02 U3326 ( .S(n3540), .A0(n2267), .A1(n2477), .Z(n2535));
Q_MX02 U3327 ( .S(n3540), .A0(n2266), .A1(n2475), .Z(n2534));
Q_MX02 U3328 ( .S(n3540), .A0(n2265), .A1(n2473), .Z(n2533));
Q_MX02 U3329 ( .S(n3540), .A0(n2264), .A1(n2471), .Z(n2532));
Q_MX02 U3330 ( .S(n3540), .A0(n2263), .A1(n2469), .Z(n2531));
Q_MX02 U3331 ( .S(n3540), .A0(n2262), .A1(n2467), .Z(n2530));
Q_XOR2 U3332 ( .A0(n2528), .A1(n2464), .Z(n2529));
Q_AD01HF U3333 ( .A0(n2526), .B0(n2463), .S(n2527), .CO(n2528));
Q_AD01HF U3334 ( .A0(n2524), .B0(n2462), .S(n2525), .CO(n2526));
Q_AD01HF U3335 ( .A0(n2522), .B0(n2461), .S(n2523), .CO(n2524));
Q_AD01HF U3336 ( .A0(n2520), .B0(n2460), .S(n2521), .CO(n2522));
Q_AD01HF U3337 ( .A0(n2518), .B0(n2459), .S(n2519), .CO(n2520));
Q_AD01HF U3338 ( .A0(n2516), .B0(n2458), .S(n2517), .CO(n2518));
Q_AD01HF U3339 ( .A0(n2514), .B0(n2457), .S(n2515), .CO(n2516));
Q_AD01HF U3340 ( .A0(n2512), .B0(n2456), .S(n2513), .CO(n2514));
Q_AD01HF U3341 ( .A0(n2510), .B0(n2455), .S(n2511), .CO(n2512));
Q_AD01HF U3342 ( .A0(n2508), .B0(n2454), .S(n2509), .CO(n2510));
Q_AD01HF U3343 ( .A0(n2506), .B0(n2453), .S(n2507), .CO(n2508));
Q_AD01HF U3344 ( .A0(n2504), .B0(n2452), .S(n2505), .CO(n2506));
Q_AD01HF U3345 ( .A0(n2502), .B0(n2451), .S(n2503), .CO(n2504));
Q_AD01HF U3346 ( .A0(n2500), .B0(n2450), .S(n2501), .CO(n2502));
Q_AD01HF U3347 ( .A0(n2498), .B0(n2449), .S(n2499), .CO(n2500));
Q_AD01HF U3348 ( .A0(n2496), .B0(n2448), .S(n2497), .CO(n2498));
Q_AD01HF U3349 ( .A0(n2494), .B0(n2447), .S(n2495), .CO(n2496));
Q_AD01HF U3350 ( .A0(n2492), .B0(n2446), .S(n2493), .CO(n2494));
Q_AD01HF U3351 ( .A0(n2490), .B0(n2445), .S(n2491), .CO(n2492));
Q_AD01HF U3352 ( .A0(n2488), .B0(n2444), .S(n2489), .CO(n2490));
Q_AD01HF U3353 ( .A0(n2486), .B0(n2443), .S(n2487), .CO(n2488));
Q_AD01HF U3354 ( .A0(n2484), .B0(n2442), .S(n2485), .CO(n2486));
Q_AD01HF U3355 ( .A0(n2482), .B0(n2441), .S(n2483), .CO(n2484));
Q_AD01HF U3356 ( .A0(n2480), .B0(n2440), .S(n2481), .CO(n2482));
Q_AD01HF U3357 ( .A0(n2478), .B0(n2439), .S(n2479), .CO(n2480));
Q_AD01HF U3358 ( .A0(n2476), .B0(n2438), .S(n2477), .CO(n2478));
Q_AD01HF U3359 ( .A0(n2474), .B0(n2437), .S(n2475), .CO(n2476));
Q_AD01HF U3360 ( .A0(n2472), .B0(n2436), .S(n2473), .CO(n2474));
Q_AD01HF U3361 ( .A0(n2470), .B0(n2435), .S(n2471), .CO(n2472));
Q_AD01HF U3362 ( .A0(n2468), .B0(n2434), .S(n2469), .CO(n2470));
Q_AD01HF U3363 ( .A0(n2433), .B0(n2466), .S(n2467), .CO(n2468));
Q_OR02 U3364 ( .A0(n2465), .A1(n3564), .Z(n2466));
Q_MX02 U3365 ( .S(_zyL439_meState8[0]), .A0(n2293), .A1(error_cntr[31]), .Z(n2464));
Q_MX02 U3366 ( .S(_zyL439_meState8[0]), .A0(n2292), .A1(error_cntr[30]), .Z(n2463));
Q_MX02 U3367 ( .S(_zyL439_meState8[0]), .A0(n2291), .A1(error_cntr[29]), .Z(n2462));
Q_MX02 U3368 ( .S(_zyL439_meState8[0]), .A0(n2290), .A1(error_cntr[28]), .Z(n2461));
Q_MX02 U3369 ( .S(_zyL439_meState8[0]), .A0(n2289), .A1(error_cntr[27]), .Z(n2460));
Q_MX02 U3370 ( .S(_zyL439_meState8[0]), .A0(n2288), .A1(error_cntr[26]), .Z(n2459));
Q_MX02 U3371 ( .S(_zyL439_meState8[0]), .A0(n2287), .A1(error_cntr[25]), .Z(n2458));
Q_MX02 U3372 ( .S(_zyL439_meState8[0]), .A0(n2286), .A1(error_cntr[24]), .Z(n2457));
Q_MX02 U3373 ( .S(_zyL439_meState8[0]), .A0(n2285), .A1(error_cntr[23]), .Z(n2456));
Q_MX02 U3374 ( .S(_zyL439_meState8[0]), .A0(n2284), .A1(error_cntr[22]), .Z(n2455));
Q_MX02 U3375 ( .S(_zyL439_meState8[0]), .A0(n2283), .A1(error_cntr[21]), .Z(n2454));
Q_MX02 U3376 ( .S(_zyL439_meState8[0]), .A0(n2282), .A1(error_cntr[20]), .Z(n2453));
Q_MX02 U3377 ( .S(_zyL439_meState8[0]), .A0(n2281), .A1(error_cntr[19]), .Z(n2452));
Q_MX02 U3378 ( .S(_zyL439_meState8[0]), .A0(n2280), .A1(error_cntr[18]), .Z(n2451));
Q_MX02 U3379 ( .S(_zyL439_meState8[0]), .A0(n2279), .A1(error_cntr[17]), .Z(n2450));
Q_MX02 U3380 ( .S(_zyL439_meState8[0]), .A0(n2278), .A1(error_cntr[16]), .Z(n2449));
Q_MX02 U3381 ( .S(_zyL439_meState8[0]), .A0(n2277), .A1(error_cntr[15]), .Z(n2448));
Q_MX02 U3382 ( .S(_zyL439_meState8[0]), .A0(n2276), .A1(error_cntr[14]), .Z(n2447));
Q_MX02 U3383 ( .S(_zyL439_meState8[0]), .A0(n2275), .A1(error_cntr[13]), .Z(n2446));
Q_MX02 U3384 ( .S(_zyL439_meState8[0]), .A0(n2274), .A1(error_cntr[12]), .Z(n2445));
Q_MX02 U3385 ( .S(_zyL439_meState8[0]), .A0(n2273), .A1(error_cntr[11]), .Z(n2444));
Q_MX02 U3386 ( .S(_zyL439_meState8[0]), .A0(n2272), .A1(error_cntr[10]), .Z(n2443));
Q_MX02 U3387 ( .S(_zyL439_meState8[0]), .A0(n2271), .A1(error_cntr[9]), .Z(n2442));
Q_MX02 U3388 ( .S(_zyL439_meState8[0]), .A0(n2270), .A1(error_cntr[8]), .Z(n2441));
Q_MX02 U3389 ( .S(_zyL439_meState8[0]), .A0(n2269), .A1(error_cntr[7]), .Z(n2440));
Q_MX02 U3390 ( .S(_zyL439_meState8[0]), .A0(n2268), .A1(error_cntr[6]), .Z(n2439));
Q_MX02 U3391 ( .S(_zyL439_meState8[0]), .A0(n2267), .A1(error_cntr[5]), .Z(n2438));
Q_MX02 U3392 ( .S(_zyL439_meState8[0]), .A0(n2266), .A1(error_cntr[4]), .Z(n2437));
Q_MX02 U3393 ( .S(_zyL439_meState8[0]), .A0(n2265), .A1(error_cntr[3]), .Z(n2436));
Q_MX02 U3394 ( .S(_zyL439_meState8[0]), .A0(n2264), .A1(error_cntr[2]), .Z(n2435));
Q_MX02 U3395 ( .S(_zyL439_meState8[0]), .A0(n2263), .A1(error_cntr[1]), .Z(n2434));
Q_MX02 U3396 ( .S(_zyL439_meState8[0]), .A0(n2262), .A1(error_cntr[0]), .Z(n2433));
Q_INV U3397 ( .A(n2432), .Z(n3560));
Q_NR02 U3398 ( .A0(n2431), .A1(n2430), .Z(n2432));
Q_MX02 U3399 ( .S(n3535), .A0(n2394), .A1(n2423), .Z(n2431));
Q_MX02 U3400 ( .S(n3535), .A0(n2393), .A1(n2426), .Z(n2430));
Q_MX02 U3401 ( .S(n3535), .A0(n2392), .A1(n2425), .Z(n2429));
Q_MX02 U3402 ( .S(n3535), .A0(n2391), .A1(n2424), .Z(n2428));
Q_MX02 U3403 ( .S(n3535), .A0(n2390), .A1(n2416), .Z(n2427));
Q_INV U3404 ( .A(n2421), .Z(n2426));
Q_INV U3405 ( .A(n2420), .Z(n2425));
Q_INV U3406 ( .A(n2418), .Z(n2424));
Q_AD02 U3407 ( .CI(n2419), .A0(_zygsfis_ob_service_data_wptr[2]), .A1(_zygsfis_ob_service_data_wptr[3]), .B0(n2414), .B1(n2415), .S0(n2420), .S1(n2421), .CO(n2422));
Q_AD01 U3408 ( .CI(n2413), .A0(_zygsfis_ob_service_data_wptr[1]), .B0(n2417), .S(n2418), .CO(n2419));
Q_OR02 U3409 ( .A0(_zygsfis_ob_service_data_wptr[0]), .A1(n2412), .Z(n2417));
Q_XOR2 U3410 ( .A0(_zygsfis_ob_service_data_wptr[0]), .A1(n2412), .Z(n2416));
Q_XOR3 U3411 ( .A0(_zygsfis_ob_service_data_wptr[4]), .A1(n2405), .A2(n2422), .Z(n2423));
Q_INV U3412 ( .A(n2404), .Z(n2415));
Q_INV U3413 ( .A(n2403), .Z(n2414));
Q_INV U3414 ( .A(n2402), .Z(n2413));
Q_INV U3415 ( .A(n2401), .Z(n2412));
Q_AN02 U3416 ( .A0(n2411), .A1(_zygsfis_ob_service_data_eos), .Z(n3557));
Q_AN03 U3417 ( .A0(n2408), .A1(n2409), .A2(n2410), .Z(n2411));
Q_AN03 U3418 ( .A0(n2416), .A1(n2406), .A2(n2407), .Z(n2410));
Q_XNR2 U3419 ( .A0(n2405), .A1(_zygsfis_ob_service_data_wptr[4]), .Z(n2409));
Q_XNR2 U3420 ( .A0(n2404), .A1(_zygsfis_ob_service_data_wptr[3]), .Z(n2408));
Q_XNR2 U3421 ( .A0(n2403), .A1(_zygsfis_ob_service_data_wptr[2]), .Z(n2407));
Q_XNR2 U3422 ( .A0(n2402), .A1(_zygsfis_ob_service_data_wptr[1]), .Z(n2406));
Q_MX02 U3423 ( .S(n1789), .A0(n2399), .A1(_zygsfis_ob_service_data_rptr[3]), .Z(n2404));
Q_MX02 U3424 ( .S(n1789), .A0(n2397), .A1(_zygsfis_ob_service_data_rptr[2]), .Z(n2403));
Q_MX02 U3425 ( .S(n1789), .A0(n2395), .A1(_zygsfis_ob_service_data_rptr[1]), .Z(n2402));
Q_XOR2 U3426 ( .A0(n3534), .A1(_zygsfis_ob_service_data_rptr[0]), .Z(n2401));
Q_XOR2 U3427 ( .A0(_zygsfis_ob_service_data_rptr[4]), .A1(n5879), .Z(n2405));
Q_AD01HF U3428 ( .A0(_zygsfis_ob_service_data_rptr[3]), .B0(n2398), .S(n2399), .CO(n2400));
Q_AD01HF U3429 ( .A0(_zygsfis_ob_service_data_rptr[2]), .B0(n2396), .S(n2397), .CO(n2398));
Q_AD01HF U3430 ( .A0(_zygsfis_ob_service_data_rptr[1]), .B0(_zygsfis_ob_service_data_rptr[0]), .S(n2395), .CO(n2396));
Q_MX02 U3431 ( .S(n1789), .A0(n2388), .A1(_zygsfis_ob_service_data_space[3]), .Z(n2393));
Q_MX02 U3432 ( .S(n1789), .A0(n2386), .A1(_zygsfis_ob_service_data_space[2]), .Z(n2392));
Q_MX02 U3433 ( .S(n1789), .A0(n2384), .A1(_zygsfis_ob_service_data_space[1]), .Z(n2391));
Q_XOR2 U3434 ( .A0(n3534), .A1(_zygsfis_ob_service_data_space[0]), .Z(n2390));
Q_XOR2 U3435 ( .A0(_zygsfis_ob_service_data_space[4]), .A1(n5880), .Z(n2394));
Q_AD01HF U3436 ( .A0(_zygsfis_ob_service_data_space[3]), .B0(n2387), .S(n2388), .CO(n2389));
Q_AD01HF U3437 ( .A0(_zygsfis_ob_service_data_space[2]), .B0(n2385), .S(n2386), .CO(n2387));
Q_AD01HF U3438 ( .A0(_zygsfis_ob_service_data_space[1]), .B0(_zygsfis_ob_service_data_space[0]), .S(n2384), .CO(n2385));
Q_AD01HF U3439 ( .A0(_zygsfis_ob_service_data_req[3]), .B0(n2381), .S(n2382), .CO(n2383));
Q_AD01HF U3440 ( .A0(_zygsfis_ob_service_data_req[2]), .B0(n2379), .S(n2380), .CO(n2381));
Q_AD01HF U3441 ( .A0(_zygsfis_ob_service_data_req[1]), .B0(_zygsfis_ob_service_data_req[0]), .S(n2378), .CO(n2379));
Q_INV U3442 ( .A(n2355), .Z(n2377));
Q_OR03 U3443 ( .A0(n2365), .A1(n2375), .A2(n2374), .Z(n2376));
Q_AO21 U3444 ( .A0(n2372), .A1(n2368), .B0(n2373), .Z(n2374));
Q_AN03 U3445 ( .A0(n2372), .A1(n2301), .A2(n2369), .Z(n2373));
Q_AN02 U3446 ( .A0(n2319), .A1(n2366), .Z(n2372));
Q_OR03 U3447 ( .A0(n2357), .A1(n2359), .A2(n2370), .Z(n2371));
Q_OR03 U3448 ( .A0(n2297), .A1(n2295), .A2(n2294), .Z(n2369));
Q_OR03 U3449 ( .A0(n2305), .A1(n2303), .A2(n2367), .Z(n2368));
Q_AN02 U3450 ( .A0(n2301), .A1(n2299), .Z(n2367));
Q_AN03 U3451 ( .A0(n2366), .A1(n2307), .A2(n2319), .Z(n2375));
Q_AN03 U3452 ( .A0(n2313), .A1(n2311), .A2(n2309), .Z(n2366));
Q_AO21 U3453 ( .A0(n2319), .A1(n2364), .B0(n2321), .Z(n2365));
Q_OR02 U3454 ( .A0(n2317), .A1(n2315), .Z(n2364));
Q_OR03 U3455 ( .A0(n2363), .A1(n2362), .A2(n2361), .Z(n2370));
Q_OR02 U3456 ( .A0(n2329), .A1(n2327), .Z(n2363));
Q_OR02 U3457 ( .A0(n2325), .A1(n2323), .Z(n2362));
Q_OR03 U3458 ( .A0(n2337), .A1(n2335), .A2(n2360), .Z(n2361));
Q_OR02 U3459 ( .A0(n2333), .A1(n2331), .Z(n2360));
Q_OR03 U3460 ( .A0(n2345), .A1(n2343), .A2(n2358), .Z(n2359));
Q_OR02 U3461 ( .A0(n2341), .A1(n2339), .Z(n2358));
Q_OR03 U3462 ( .A0(n2353), .A1(n2351), .A2(n2356), .Z(n2357));
Q_OR02 U3463 ( .A0(n2349), .A1(n2347), .Z(n2356));
Q_XOR2 U3464 ( .A0(watchdog_timer[31]), .A1(n2354), .Z(n2355));
Q_AD01HF U3465 ( .A0(watchdog_timer[30]), .B0(n2352), .S(n2353), .CO(n2354));
Q_AD01HF U3466 ( .A0(watchdog_timer[29]), .B0(n2350), .S(n2351), .CO(n2352));
Q_AD01HF U3467 ( .A0(watchdog_timer[28]), .B0(n2348), .S(n2349), .CO(n2350));
Q_AD01HF U3468 ( .A0(watchdog_timer[27]), .B0(n2346), .S(n2347), .CO(n2348));
Q_AD01HF U3469 ( .A0(watchdog_timer[26]), .B0(n2344), .S(n2345), .CO(n2346));
Q_AD01HF U3470 ( .A0(watchdog_timer[25]), .B0(n2342), .S(n2343), .CO(n2344));
Q_AD01HF U3471 ( .A0(watchdog_timer[24]), .B0(n2340), .S(n2341), .CO(n2342));
Q_AD01HF U3472 ( .A0(watchdog_timer[23]), .B0(n2338), .S(n2339), .CO(n2340));
Q_AD01HF U3473 ( .A0(watchdog_timer[22]), .B0(n2336), .S(n2337), .CO(n2338));
Q_AD01HF U3474 ( .A0(watchdog_timer[21]), .B0(n2334), .S(n2335), .CO(n2336));
Q_AD01HF U3475 ( .A0(watchdog_timer[20]), .B0(n2332), .S(n2333), .CO(n2334));
Q_AD01HF U3476 ( .A0(watchdog_timer[19]), .B0(n2330), .S(n2331), .CO(n2332));
Q_AD01HF U3477 ( .A0(watchdog_timer[18]), .B0(n2328), .S(n2329), .CO(n2330));
Q_AD01HF U3478 ( .A0(watchdog_timer[17]), .B0(n2326), .S(n2327), .CO(n2328));
Q_AD01HF U3479 ( .A0(watchdog_timer[16]), .B0(n2324), .S(n2325), .CO(n2326));
Q_AD01HF U3480 ( .A0(watchdog_timer[15]), .B0(n2322), .S(n2323), .CO(n2324));
Q_AD01HF U3481 ( .A0(watchdog_timer[14]), .B0(n2320), .S(n2321), .CO(n2322));
Q_AD01HF U3482 ( .A0(watchdog_timer[13]), .B0(n2318), .S(n2319), .CO(n2320));
Q_AD01HF U3483 ( .A0(watchdog_timer[12]), .B0(n2316), .S(n2317), .CO(n2318));
Q_AD01HF U3484 ( .A0(watchdog_timer[11]), .B0(n2314), .S(n2315), .CO(n2316));
Q_AD01HF U3485 ( .A0(watchdog_timer[10]), .B0(n2312), .S(n2313), .CO(n2314));
Q_AD01HF U3486 ( .A0(watchdog_timer[9]), .B0(n2310), .S(n2311), .CO(n2312));
Q_AD01HF U3487 ( .A0(watchdog_timer[8]), .B0(n2308), .S(n2309), .CO(n2310));
Q_AD01HF U3488 ( .A0(watchdog_timer[7]), .B0(n2306), .S(n2307), .CO(n2308));
Q_AD01HF U3489 ( .A0(watchdog_timer[6]), .B0(n2304), .S(n2305), .CO(n2306));
Q_AD01HF U3490 ( .A0(watchdog_timer[5]), .B0(n2302), .S(n2303), .CO(n2304));
Q_AD01HF U3491 ( .A0(watchdog_timer[4]), .B0(n2300), .S(n2301), .CO(n2302));
Q_AD01HF U3492 ( .A0(watchdog_timer[3]), .B0(n2298), .S(n2299), .CO(n2300));
Q_AD01HF U3493 ( .A0(watchdog_timer[2]), .B0(n2296), .S(n2297), .CO(n2298));
Q_AD01HF U3494 ( .A0(watchdog_timer[1]), .B0(watchdog_timer[0]), .S(n2295), .CO(n2296));
Q_MX02 U3495 ( .S(n3539), .A0(error_cntr[31]), .A1(n2261), .Z(n2293));
Q_MX02 U3496 ( .S(n3539), .A0(error_cntr[30]), .A1(n2259), .Z(n2292));
Q_MX02 U3497 ( .S(n3539), .A0(error_cntr[29]), .A1(n2257), .Z(n2291));
Q_MX02 U3498 ( .S(n3539), .A0(error_cntr[28]), .A1(n2255), .Z(n2290));
Q_MX02 U3499 ( .S(n3539), .A0(error_cntr[27]), .A1(n2253), .Z(n2289));
Q_MX02 U3500 ( .S(n3539), .A0(error_cntr[26]), .A1(n2251), .Z(n2288));
Q_MX02 U3501 ( .S(n3539), .A0(error_cntr[25]), .A1(n2249), .Z(n2287));
Q_MX02 U3502 ( .S(n3539), .A0(error_cntr[24]), .A1(n2247), .Z(n2286));
Q_MX02 U3503 ( .S(n3539), .A0(error_cntr[23]), .A1(n2245), .Z(n2285));
Q_MX02 U3504 ( .S(n3539), .A0(error_cntr[22]), .A1(n2243), .Z(n2284));
Q_MX02 U3505 ( .S(n3539), .A0(error_cntr[21]), .A1(n2241), .Z(n2283));
Q_MX02 U3506 ( .S(n3539), .A0(error_cntr[20]), .A1(n2239), .Z(n2282));
Q_MX02 U3507 ( .S(n3539), .A0(error_cntr[19]), .A1(n2237), .Z(n2281));
Q_MX02 U3508 ( .S(n3539), .A0(error_cntr[18]), .A1(n2235), .Z(n2280));
Q_MX02 U3509 ( .S(n3539), .A0(error_cntr[17]), .A1(n2233), .Z(n2279));
Q_MX02 U3510 ( .S(n3539), .A0(error_cntr[16]), .A1(n2231), .Z(n2278));
Q_MX02 U3511 ( .S(n3539), .A0(error_cntr[15]), .A1(n2229), .Z(n2277));
Q_MX02 U3512 ( .S(n3539), .A0(error_cntr[14]), .A1(n2227), .Z(n2276));
Q_MX02 U3513 ( .S(n3539), .A0(error_cntr[13]), .A1(n2225), .Z(n2275));
Q_MX02 U3514 ( .S(n3539), .A0(error_cntr[12]), .A1(n2223), .Z(n2274));
Q_MX02 U3515 ( .S(n3539), .A0(error_cntr[11]), .A1(n2221), .Z(n2273));
Q_MX02 U3516 ( .S(n3539), .A0(error_cntr[10]), .A1(n2219), .Z(n2272));
Q_MX02 U3517 ( .S(n3539), .A0(error_cntr[9]), .A1(n2217), .Z(n2271));
Q_MX02 U3518 ( .S(n3539), .A0(error_cntr[8]), .A1(n2215), .Z(n2270));
Q_MX02 U3519 ( .S(n3539), .A0(error_cntr[7]), .A1(n2213), .Z(n2269));
Q_MX02 U3520 ( .S(n3539), .A0(error_cntr[6]), .A1(n2211), .Z(n2268));
Q_MX02 U3521 ( .S(n3539), .A0(error_cntr[5]), .A1(n2209), .Z(n2267));
Q_MX02 U3522 ( .S(n3539), .A0(error_cntr[4]), .A1(n2207), .Z(n2266));
Q_MX02 U3523 ( .S(n3539), .A0(error_cntr[3]), .A1(n2205), .Z(n2265));
Q_MX02 U3524 ( .S(n3539), .A0(error_cntr[2]), .A1(n2203), .Z(n2264));
Q_MX02 U3525 ( .S(n3539), .A0(error_cntr[1]), .A1(n2201), .Z(n2263));
Q_XOR2 U3526 ( .A0(n3539), .A1(error_cntr[0]), .Z(n2262));
Q_XOR2 U3527 ( .A0(error_cntr[31]), .A1(n2260), .Z(n2261));
Q_AD01HF U3528 ( .A0(error_cntr[30]), .B0(n2258), .S(n2259), .CO(n2260));
Q_AD01HF U3529 ( .A0(error_cntr[29]), .B0(n2256), .S(n2257), .CO(n2258));
Q_AD01HF U3530 ( .A0(error_cntr[28]), .B0(n2254), .S(n2255), .CO(n2256));
Q_AD01HF U3531 ( .A0(error_cntr[27]), .B0(n2252), .S(n2253), .CO(n2254));
Q_AD01HF U3532 ( .A0(error_cntr[26]), .B0(n2250), .S(n2251), .CO(n2252));
Q_AD01HF U3533 ( .A0(error_cntr[25]), .B0(n2248), .S(n2249), .CO(n2250));
Q_AD01HF U3534 ( .A0(error_cntr[24]), .B0(n2246), .S(n2247), .CO(n2248));
Q_AD01HF U3535 ( .A0(error_cntr[23]), .B0(n2244), .S(n2245), .CO(n2246));
Q_AD01HF U3536 ( .A0(error_cntr[22]), .B0(n2242), .S(n2243), .CO(n2244));
Q_AD01HF U3537 ( .A0(error_cntr[21]), .B0(n2240), .S(n2241), .CO(n2242));
Q_AD01HF U3538 ( .A0(error_cntr[20]), .B0(n2238), .S(n2239), .CO(n2240));
Q_AD01HF U3539 ( .A0(error_cntr[19]), .B0(n2236), .S(n2237), .CO(n2238));
Q_AD01HF U3540 ( .A0(error_cntr[18]), .B0(n2234), .S(n2235), .CO(n2236));
Q_AD01HF U3541 ( .A0(error_cntr[17]), .B0(n2232), .S(n2233), .CO(n2234));
Q_AD01HF U3542 ( .A0(error_cntr[16]), .B0(n2230), .S(n2231), .CO(n2232));
Q_AD01HF U3543 ( .A0(error_cntr[15]), .B0(n2228), .S(n2229), .CO(n2230));
Q_AD01HF U3544 ( .A0(error_cntr[14]), .B0(n2226), .S(n2227), .CO(n2228));
Q_AD01HF U3545 ( .A0(error_cntr[13]), .B0(n2224), .S(n2225), .CO(n2226));
Q_AD01HF U3546 ( .A0(error_cntr[12]), .B0(n2222), .S(n2223), .CO(n2224));
Q_AD01HF U3547 ( .A0(error_cntr[11]), .B0(n2220), .S(n2221), .CO(n2222));
Q_AD01HF U3548 ( .A0(error_cntr[10]), .B0(n2218), .S(n2219), .CO(n2220));
Q_AD01HF U3549 ( .A0(error_cntr[9]), .B0(n2216), .S(n2217), .CO(n2218));
Q_AD01HF U3550 ( .A0(error_cntr[8]), .B0(n2214), .S(n2215), .CO(n2216));
Q_AD01HF U3551 ( .A0(error_cntr[7]), .B0(n2212), .S(n2213), .CO(n2214));
Q_AD01HF U3552 ( .A0(error_cntr[6]), .B0(n2210), .S(n2211), .CO(n2212));
Q_AD01HF U3553 ( .A0(error_cntr[5]), .B0(n2208), .S(n2209), .CO(n2210));
Q_AD01HF U3554 ( .A0(error_cntr[4]), .B0(n2206), .S(n2207), .CO(n2208));
Q_AD01HF U3555 ( .A0(error_cntr[3]), .B0(n2204), .S(n2205), .CO(n2206));
Q_AD01HF U3556 ( .A0(error_cntr[2]), .B0(n2202), .S(n2203), .CO(n2204));
Q_AD01HF U3557 ( .A0(error_cntr[1]), .B0(error_cntr[0]), .S(n2201), .CO(n2202));
Q_OR02 U3558 ( .A0(n3544), .A1(saw_stats), .Z(n3567));
Q_OR02 U3559 ( .A0(n3249), .A1(saw_stats), .Z(n3565));
Q_INV U3560 ( .A(n2200), .Z(n3538));
Q_OR02 U3561 ( .A0(n2198), .A1(n2199), .Z(n2200));
Q_OR03 U3562 ( .A0(n2195), .A1(n2196), .A2(n2197), .Z(n2199));
Q_OR03 U3563 ( .A0(n2192), .A1(n2193), .A2(n2194), .Z(n2198));
Q_OR03 U3564 ( .A0(n2189), .A1(n2190), .A2(n2191), .Z(n2197));
Q_OR03 U3565 ( .A0(n2186), .A1(n2187), .A2(n2188), .Z(n2196));
Q_OR03 U3566 ( .A0(n2184), .A1(n2183), .A2(n2185), .Z(n2195));
Q_OR03 U3567 ( .A0(n2155), .A1(n2154), .A2(n2153), .Z(n2194));
Q_OR03 U3568 ( .A0(n2158), .A1(n2157), .A2(n2156), .Z(n2193));
Q_OR03 U3569 ( .A0(n2161), .A1(n2160), .A2(n2159), .Z(n2192));
Q_OR03 U3570 ( .A0(n2164), .A1(n2163), .A2(n2162), .Z(n2191));
Q_OR03 U3571 ( .A0(n2167), .A1(n2166), .A2(n2165), .Z(n2190));
Q_OR03 U3572 ( .A0(n2170), .A1(n2169), .A2(n2168), .Z(n2189));
Q_OR03 U3573 ( .A0(n2173), .A1(n2172), .A2(n2171), .Z(n2188));
Q_OR03 U3574 ( .A0(n2176), .A1(n2175), .A2(n2174), .Z(n2187));
Q_OR03 U3575 ( .A0(n2179), .A1(n2178), .A2(n2177), .Z(n2186));
Q_OR03 U3576 ( .A0(n2182), .A1(n2181), .A2(n2180), .Z(n2185));
Q_INV U3577 ( .A(n2152), .Z(n2184));
Q_INV U3578 ( .A(n2151), .Z(n2183));
Q_MX02 U3579 ( .S(n1789), .A0(n3502), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [31]), .Z(n2182));
Q_MX02 U3580 ( .S(n1789), .A0(n3503), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [30]), .Z(n2181));
Q_MX02 U3581 ( .S(n1789), .A0(n3504), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [29]), .Z(n2180));
Q_MX02 U3582 ( .S(n1789), .A0(n3505), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [28]), .Z(n2179));
Q_MX02 U3583 ( .S(n1789), .A0(n3506), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [27]), .Z(n2178));
Q_MX02 U3584 ( .S(n1789), .A0(n3507), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [26]), .Z(n2177));
Q_MX02 U3585 ( .S(n1789), .A0(n3508), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [25]), .Z(n2176));
Q_MX02 U3586 ( .S(n1789), .A0(n3509), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [24]), .Z(n2175));
Q_MX02 U3587 ( .S(n1789), .A0(n3510), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [23]), .Z(n2174));
Q_MX02 U3588 ( .S(n1789), .A0(n3511), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [22]), .Z(n2173));
Q_MX02 U3589 ( .S(n1789), .A0(n3512), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [21]), .Z(n2172));
Q_MX02 U3590 ( .S(n1789), .A0(n3513), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [20]), .Z(n2171));
Q_MX02 U3591 ( .S(n1789), .A0(n3514), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [19]), .Z(n2170));
Q_MX02 U3592 ( .S(n1789), .A0(n3515), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [18]), .Z(n2169));
Q_MX02 U3593 ( .S(n1789), .A0(n3516), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [17]), .Z(n2168));
Q_MX02 U3594 ( .S(n1789), .A0(n3517), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [16]), .Z(n2167));
Q_MX02 U3595 ( .S(n1789), .A0(n3518), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [15]), .Z(n2166));
Q_MX02 U3596 ( .S(n1789), .A0(n3519), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [14]), .Z(n2165));
Q_MX02 U3597 ( .S(n1789), .A0(n3520), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [13]), .Z(n2164));
Q_MX02 U3598 ( .S(n1789), .A0(n3521), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [12]), .Z(n2163));
Q_MX02 U3599 ( .S(n1789), .A0(n3522), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [11]), .Z(n2162));
Q_MX02 U3600 ( .S(n1789), .A0(n3523), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [10]), .Z(n2161));
Q_MX02 U3601 ( .S(n1789), .A0(n3524), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [9]), .Z(n2160));
Q_MX02 U3602 ( .S(n1789), .A0(n3525), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [8]), .Z(n2159));
Q_MX02 U3603 ( .S(n1789), .A0(n3526), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [7]), .Z(n2158));
Q_MX02 U3604 ( .S(n1789), .A0(n3527), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [6]), .Z(n2157));
Q_MX02 U3605 ( .S(n1789), .A0(n3528), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [5]), .Z(n2156));
Q_MX02 U3606 ( .S(n1789), .A0(n3529), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [4]), .Z(n2155));
Q_MX02 U3607 ( .S(n1789), .A0(n3530), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [3]), .Z(n2154));
Q_MX02 U3608 ( .S(n1789), .A0(n3531), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [2]), .Z(n2153));
Q_MX02 U3609 ( .S(n1789), .A0(n3532), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [1]), .Z(n2152));
Q_MX02 U3610 ( .S(n1789), .A0(n3533), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [0]), .Z(n2151));
Q_INV U3611 ( .A(n2150), .Z(n3542));
Q_AN02 U3612 ( .A0(n2148), .A1(n2149), .Z(n2150));
Q_AN03 U3613 ( .A0(n2140), .A1(n2139), .A2(n2147), .Z(n2149));
Q_AN03 U3614 ( .A0(n2143), .A1(n2142), .A2(n2141), .Z(n2148));
Q_AN03 U3615 ( .A0(n2146), .A1(n2145), .A2(n2144), .Z(n2147));
Q_XNR2 U3616 ( .A0(kme_ob_tstrb[7]), .A1(n2138), .Z(n2146));
Q_XNR2 U3617 ( .A0(kme_ob_tstrb[6]), .A1(n2137), .Z(n2145));
Q_XNR2 U3618 ( .A0(kme_ob_tstrb[5]), .A1(n2136), .Z(n2144));
Q_XNR2 U3619 ( .A0(kme_ob_tstrb[4]), .A1(n2135), .Z(n2143));
Q_XNR2 U3620 ( .A0(kme_ob_tstrb[3]), .A1(n2134), .Z(n2142));
Q_XNR2 U3621 ( .A0(kme_ob_tstrb[2]), .A1(n2133), .Z(n2141));
Q_XNR2 U3622 ( .A0(kme_ob_tstrb[1]), .A1(n2132), .Z(n2140));
Q_XNR2 U3623 ( .A0(kme_ob_tstrb[0]), .A1(n2131), .Z(n2139));
Q_MX02 U3624 ( .S(n1789), .A0(n3494), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytstrb_L209_tfiV13 [7]), .Z(n2138));
Q_MX02 U3625 ( .S(n1789), .A0(n3495), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytstrb_L209_tfiV13 [6]), .Z(n2137));
Q_MX02 U3626 ( .S(n1789), .A0(n3496), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytstrb_L209_tfiV13 [5]), .Z(n2136));
Q_MX02 U3627 ( .S(n1789), .A0(n3497), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytstrb_L209_tfiV13 [4]), .Z(n2135));
Q_MX02 U3628 ( .S(n1789), .A0(n3498), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytstrb_L209_tfiV13 [3]), .Z(n2134));
Q_MX02 U3629 ( .S(n1789), .A0(n3499), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytstrb_L209_tfiV13 [2]), .Z(n2133));
Q_MX02 U3630 ( .S(n1789), .A0(n3500), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytstrb_L209_tfiV13 [1]), .Z(n2132));
Q_MX02 U3631 ( .S(n1789), .A0(n3501), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytstrb_L209_tfiV13 [0]), .Z(n2131));
Q_OR02 U3632 ( .A0(n2128), .A1(n2129), .Z(n2130));
Q_OR03 U3633 ( .A0(n2125), .A1(n2126), .A2(n2127), .Z(n2129));
Q_OR03 U3634 ( .A0(n2122), .A1(n2123), .A2(n2124), .Z(n2128));
Q_OR03 U3635 ( .A0(n2119), .A1(n2120), .A2(n2121), .Z(n2127));
Q_OR03 U3636 ( .A0(n2116), .A1(n2117), .A2(n2118), .Z(n2126));
Q_OR03 U3637 ( .A0(n2110), .A1(n2077), .A2(n2115), .Z(n2125));
Q_OR03 U3638 ( .A0(n2081), .A1(n2111), .A2(n2079), .Z(n2124));
Q_OR03 U3639 ( .A0(n2084), .A1(n2083), .A2(n2082), .Z(n2123));
Q_OR03 U3640 ( .A0(n2087), .A1(n2086), .A2(n2085), .Z(n2122));
Q_OR03 U3641 ( .A0(n2090), .A1(n2089), .A2(n2088), .Z(n2121));
Q_OR03 U3642 ( .A0(n2093), .A1(n2092), .A2(n2091), .Z(n2120));
Q_OR03 U3643 ( .A0(n2096), .A1(n2095), .A2(n2094), .Z(n2119));
Q_OR03 U3644 ( .A0(n2099), .A1(n2098), .A2(n2097), .Z(n2118));
Q_OR03 U3645 ( .A0(n2102), .A1(n2101), .A2(n2100), .Z(n2117));
Q_OR03 U3646 ( .A0(n2105), .A1(n2104), .A2(n2103), .Z(n2116));
Q_OR03 U3647 ( .A0(n2108), .A1(n2107), .A2(n2106), .Z(n2115));
Q_INV U3648 ( .A(n2114), .Z(n3537));
Q_OR02 U3649 ( .A0(n2128), .A1(n2113), .Z(n2114));
Q_OR03 U3650 ( .A0(n2112), .A1(n2126), .A2(n2127), .Z(n2113));
Q_OR03 U3651 ( .A0(n2110), .A1(n2109), .A2(n2115), .Z(n2112));
Q_INV U3652 ( .A(n2080), .Z(n2111));
Q_INV U3653 ( .A(n2078), .Z(n2110));
Q_INV U3654 ( .A(n2077), .Z(n2109));
Q_MX02 U3655 ( .S(n1789), .A0(n3462), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [31]), .Z(n2108));
Q_MX02 U3656 ( .S(n1789), .A0(n3463), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [30]), .Z(n2107));
Q_MX02 U3657 ( .S(n1789), .A0(n3464), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [29]), .Z(n2106));
Q_MX02 U3658 ( .S(n1789), .A0(n3465), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [28]), .Z(n2105));
Q_MX02 U3659 ( .S(n1789), .A0(n3466), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [27]), .Z(n2104));
Q_MX02 U3660 ( .S(n1789), .A0(n3467), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [26]), .Z(n2103));
Q_MX02 U3661 ( .S(n1789), .A0(n3468), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [25]), .Z(n2102));
Q_MX02 U3662 ( .S(n1789), .A0(n3469), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [24]), .Z(n2101));
Q_MX02 U3663 ( .S(n1789), .A0(n3470), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [23]), .Z(n2100));
Q_MX02 U3664 ( .S(n1789), .A0(n3471), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [22]), .Z(n2099));
Q_MX02 U3665 ( .S(n1789), .A0(n3472), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [21]), .Z(n2098));
Q_MX02 U3666 ( .S(n1789), .A0(n3473), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [20]), .Z(n2097));
Q_MX02 U3667 ( .S(n1789), .A0(n3474), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [19]), .Z(n2096));
Q_MX02 U3668 ( .S(n1789), .A0(n3475), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [18]), .Z(n2095));
Q_MX02 U3669 ( .S(n1789), .A0(n3476), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [17]), .Z(n2094));
Q_MX02 U3670 ( .S(n1789), .A0(n3477), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [16]), .Z(n2093));
Q_MX02 U3671 ( .S(n1789), .A0(n3478), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [15]), .Z(n2092));
Q_MX02 U3672 ( .S(n1789), .A0(n3479), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [14]), .Z(n2091));
Q_MX02 U3673 ( .S(n1789), .A0(n3480), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [13]), .Z(n2090));
Q_MX02 U3674 ( .S(n1789), .A0(n3481), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [12]), .Z(n2089));
Q_MX02 U3675 ( .S(n1789), .A0(n3482), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [11]), .Z(n2088));
Q_MX02 U3676 ( .S(n1789), .A0(n3483), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [10]), .Z(n2087));
Q_MX02 U3677 ( .S(n1789), .A0(n3484), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [9]), .Z(n2086));
Q_MX02 U3678 ( .S(n1789), .A0(n3485), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [8]), .Z(n2085));
Q_MX02 U3679 ( .S(n1789), .A0(n3486), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [7]), .Z(n2084));
Q_MX02 U3680 ( .S(n1789), .A0(n3487), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [6]), .Z(n2083));
Q_MX02 U3681 ( .S(n1789), .A0(n3488), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [5]), .Z(n2082));
Q_MX02 U3682 ( .S(n1789), .A0(n3489), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [4]), .Z(n2081));
Q_MX02 U3683 ( .S(n1789), .A0(n3490), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [3]), .Z(n2080));
Q_MX02 U3684 ( .S(n1789), .A0(n3491), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [2]), .Z(n2079));
Q_MX02 U3685 ( .S(n1789), .A0(n3492), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [1]), .Z(n2078));
Q_MX02 U3686 ( .S(n1789), .A0(n3493), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [0]), .Z(n2077));
Q_ND02 U3687 ( .A0(n2074), .A1(n2075), .Z(n2076));
Q_AN03 U3688 ( .A0(n2071), .A1(n2072), .A2(n2073), .Z(n2075));
Q_AN03 U3689 ( .A0(n2068), .A1(n2069), .A2(n2070), .Z(n2074));
Q_AN03 U3690 ( .A0(n2065), .A1(n2066), .A2(n2067), .Z(n2073));
Q_AN03 U3691 ( .A0(n2062), .A1(n2063), .A2(n2064), .Z(n2072));
Q_AN03 U3692 ( .A0(n2059), .A1(n2060), .A2(n2061), .Z(n2071));
Q_AN03 U3693 ( .A0(n2056), .A1(n2057), .A2(n2058), .Z(n2070));
Q_AN03 U3694 ( .A0(n2053), .A1(n2054), .A2(n2055), .Z(n2069));
Q_AN03 U3695 ( .A0(n2050), .A1(n2051), .A2(n2052), .Z(n2068));
Q_AN03 U3696 ( .A0(n2047), .A1(n2048), .A2(n2049), .Z(n2067));
Q_AN03 U3697 ( .A0(n1981), .A1(n2045), .A2(n2046), .Z(n2066));
Q_AN03 U3698 ( .A0(n1984), .A1(n1983), .A2(n1982), .Z(n2065));
Q_AN03 U3699 ( .A0(n1987), .A1(n1986), .A2(n1985), .Z(n2064));
Q_AN03 U3700 ( .A0(n1990), .A1(n1989), .A2(n1988), .Z(n2063));
Q_AN03 U3701 ( .A0(n1993), .A1(n1992), .A2(n1991), .Z(n2062));
Q_AN03 U3702 ( .A0(n1996), .A1(n1995), .A2(n1994), .Z(n2061));
Q_AN03 U3703 ( .A0(n1999), .A1(n1998), .A2(n1997), .Z(n2060));
Q_AN03 U3704 ( .A0(n2002), .A1(n2001), .A2(n2000), .Z(n2059));
Q_AN03 U3705 ( .A0(n2005), .A1(n2004), .A2(n2003), .Z(n2058));
Q_AN03 U3706 ( .A0(n2008), .A1(n2007), .A2(n2006), .Z(n2057));
Q_AN03 U3707 ( .A0(n2011), .A1(n2010), .A2(n2009), .Z(n2056));
Q_AN03 U3708 ( .A0(n2014), .A1(n2013), .A2(n2012), .Z(n2055));
Q_AN03 U3709 ( .A0(n2017), .A1(n2016), .A2(n2015), .Z(n2054));
Q_AN03 U3710 ( .A0(n2020), .A1(n2019), .A2(n2018), .Z(n2053));
Q_AN03 U3711 ( .A0(n2023), .A1(n2022), .A2(n2021), .Z(n2052));
Q_AN03 U3712 ( .A0(n2026), .A1(n2025), .A2(n2024), .Z(n2051));
Q_AN03 U3713 ( .A0(n2029), .A1(n2028), .A2(n2027), .Z(n2050));
Q_AN03 U3714 ( .A0(n2032), .A1(n2031), .A2(n2030), .Z(n2049));
Q_AN03 U3715 ( .A0(n2035), .A1(n2034), .A2(n2033), .Z(n2048));
Q_AN03 U3716 ( .A0(n2038), .A1(n2037), .A2(n2036), .Z(n2047));
Q_AN03 U3717 ( .A0(n2041), .A1(n2040), .A2(n2039), .Z(n2046));
Q_AN03 U3718 ( .A0(n2044), .A1(n2043), .A2(n2042), .Z(n2045));
Q_XNR2 U3719 ( .A0(kme_ob_tdata[63]), .A1(n1972), .Z(n2044));
Q_XNR2 U3720 ( .A0(kme_ob_tdata[62]), .A1(n1971), .Z(n2043));
Q_XNR2 U3721 ( .A0(kme_ob_tdata[61]), .A1(n1970), .Z(n2042));
Q_XNR2 U3722 ( .A0(kme_ob_tdata[60]), .A1(n1969), .Z(n2041));
Q_XNR2 U3723 ( .A0(kme_ob_tdata[59]), .A1(n1968), .Z(n2040));
Q_XNR2 U3724 ( .A0(kme_ob_tdata[58]), .A1(n1967), .Z(n2039));
Q_XNR2 U3725 ( .A0(kme_ob_tdata[57]), .A1(n1966), .Z(n2038));
Q_XNR2 U3726 ( .A0(kme_ob_tdata[56]), .A1(n1965), .Z(n2037));
Q_XNR2 U3727 ( .A0(kme_ob_tdata[55]), .A1(n1964), .Z(n2036));
Q_XNR2 U3728 ( .A0(kme_ob_tdata[54]), .A1(n1963), .Z(n2035));
Q_XNR2 U3729 ( .A0(kme_ob_tdata[53]), .A1(n1962), .Z(n2034));
Q_XNR2 U3730 ( .A0(kme_ob_tdata[52]), .A1(n1961), .Z(n2033));
Q_XNR2 U3731 ( .A0(kme_ob_tdata[51]), .A1(n1960), .Z(n2032));
Q_XNR2 U3732 ( .A0(kme_ob_tdata[50]), .A1(n1959), .Z(n2031));
Q_XNR2 U3733 ( .A0(kme_ob_tdata[49]), .A1(n1958), .Z(n2030));
Q_XNR2 U3734 ( .A0(kme_ob_tdata[48]), .A1(n1957), .Z(n2029));
Q_XNR2 U3735 ( .A0(kme_ob_tdata[47]), .A1(n1956), .Z(n2028));
Q_XNR2 U3736 ( .A0(kme_ob_tdata[46]), .A1(n1955), .Z(n2027));
Q_XNR2 U3737 ( .A0(kme_ob_tdata[45]), .A1(n1954), .Z(n2026));
Q_XNR2 U3738 ( .A0(kme_ob_tdata[44]), .A1(n1953), .Z(n2025));
Q_XNR2 U3739 ( .A0(kme_ob_tdata[43]), .A1(n1952), .Z(n2024));
Q_XNR2 U3740 ( .A0(kme_ob_tdata[42]), .A1(n1951), .Z(n2023));
Q_XNR2 U3741 ( .A0(kme_ob_tdata[41]), .A1(n1950), .Z(n2022));
Q_XNR2 U3742 ( .A0(kme_ob_tdata[40]), .A1(n1949), .Z(n2021));
Q_XNR2 U3743 ( .A0(kme_ob_tdata[39]), .A1(n1948), .Z(n2020));
Q_XNR2 U3744 ( .A0(kme_ob_tdata[38]), .A1(n1947), .Z(n2019));
Q_XNR2 U3745 ( .A0(kme_ob_tdata[37]), .A1(n1946), .Z(n2018));
Q_XNR2 U3746 ( .A0(kme_ob_tdata[36]), .A1(n1945), .Z(n2017));
Q_XNR2 U3747 ( .A0(kme_ob_tdata[35]), .A1(n1944), .Z(n2016));
Q_XNR2 U3748 ( .A0(kme_ob_tdata[34]), .A1(n1943), .Z(n2015));
Q_XNR2 U3749 ( .A0(kme_ob_tdata[33]), .A1(n1942), .Z(n2014));
Q_XNR2 U3750 ( .A0(kme_ob_tdata[32]), .A1(n1941), .Z(n2013));
Q_XNR2 U3751 ( .A0(kme_ob_tdata[31]), .A1(n1940), .Z(n2012));
Q_XNR2 U3752 ( .A0(kme_ob_tdata[30]), .A1(n1939), .Z(n2011));
Q_XNR2 U3753 ( .A0(kme_ob_tdata[29]), .A1(n1938), .Z(n2010));
Q_XNR2 U3754 ( .A0(kme_ob_tdata[28]), .A1(n1937), .Z(n2009));
Q_XNR2 U3755 ( .A0(kme_ob_tdata[27]), .A1(n1936), .Z(n2008));
Q_XNR2 U3756 ( .A0(kme_ob_tdata[26]), .A1(n1935), .Z(n2007));
Q_XNR2 U3757 ( .A0(kme_ob_tdata[25]), .A1(n1934), .Z(n2006));
Q_XNR2 U3758 ( .A0(kme_ob_tdata[24]), .A1(n1933), .Z(n2005));
Q_XNR2 U3759 ( .A0(kme_ob_tdata[23]), .A1(n1932), .Z(n2004));
Q_XNR2 U3760 ( .A0(kme_ob_tdata[22]), .A1(n1931), .Z(n2003));
Q_XNR2 U3761 ( .A0(kme_ob_tdata[21]), .A1(n1930), .Z(n2002));
Q_XNR2 U3762 ( .A0(kme_ob_tdata[20]), .A1(n1929), .Z(n2001));
Q_XNR2 U3763 ( .A0(kme_ob_tdata[19]), .A1(n1928), .Z(n2000));
Q_XNR2 U3764 ( .A0(kme_ob_tdata[18]), .A1(n1927), .Z(n1999));
Q_XNR2 U3765 ( .A0(kme_ob_tdata[17]), .A1(n1926), .Z(n1998));
Q_XNR2 U3766 ( .A0(kme_ob_tdata[16]), .A1(n1925), .Z(n1997));
Q_XNR2 U3767 ( .A0(kme_ob_tdata[15]), .A1(n1924), .Z(n1996));
Q_XNR2 U3768 ( .A0(kme_ob_tdata[14]), .A1(n1923), .Z(n1995));
Q_XNR2 U3769 ( .A0(kme_ob_tdata[13]), .A1(n1922), .Z(n1994));
Q_XNR2 U3770 ( .A0(kme_ob_tdata[12]), .A1(n1921), .Z(n1993));
Q_XNR2 U3771 ( .A0(kme_ob_tdata[11]), .A1(n1920), .Z(n1992));
Q_XNR2 U3772 ( .A0(kme_ob_tdata[10]), .A1(n1919), .Z(n1991));
Q_XNR2 U3773 ( .A0(kme_ob_tdata[9]), .A1(n1918), .Z(n1990));
Q_XNR2 U3774 ( .A0(kme_ob_tdata[8]), .A1(n1917), .Z(n1989));
Q_XNR2 U3775 ( .A0(kme_ob_tdata[7]), .A1(n1916), .Z(n1988));
Q_XNR2 U3776 ( .A0(kme_ob_tdata[6]), .A1(n1915), .Z(n1987));
Q_XNR2 U3777 ( .A0(kme_ob_tdata[5]), .A1(n1914), .Z(n1986));
Q_XNR2 U3778 ( .A0(kme_ob_tdata[4]), .A1(n1913), .Z(n1985));
Q_XNR2 U3779 ( .A0(kme_ob_tdata[3]), .A1(n1912), .Z(n1984));
Q_XNR2 U3780 ( .A0(kme_ob_tdata[2]), .A1(n1911), .Z(n1983));
Q_XNR2 U3781 ( .A0(kme_ob_tdata[1]), .A1(n1910), .Z(n1982));
Q_XNR2 U3782 ( .A0(kme_ob_tdata[0]), .A1(n1909), .Z(n1981));
Q_OR02 U3783 ( .A0(n1978), .A1(n1979), .Z(n1980));
Q_OR03 U3784 ( .A0(n1910), .A1(n1909), .A2(n1977), .Z(n1979));
Q_OR03 U3785 ( .A0(n1913), .A1(n1974), .A2(n1911), .Z(n1978));
Q_OR03 U3786 ( .A0(n1916), .A1(n1915), .A2(n1914), .Z(n1977));
Q_OR02 U3787 ( .A0(n1978), .A1(n1975), .Z(n1976));
Q_OR03 U3788 ( .A0(n1910), .A1(n1973), .A2(n1977), .Z(n1975));
Q_INV U3789 ( .A(n1912), .Z(n1974));
Q_INV U3790 ( .A(n1909), .Z(n1973));
Q_MX02 U3791 ( .S(n1789), .A0(n3398), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [63]), .Z(n1972));
Q_MX02 U3792 ( .S(n1789), .A0(n3399), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [62]), .Z(n1971));
Q_MX02 U3793 ( .S(n1789), .A0(n3400), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [61]), .Z(n1970));
Q_MX02 U3794 ( .S(n1789), .A0(n3401), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [60]), .Z(n1969));
Q_MX02 U3795 ( .S(n1789), .A0(n3402), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [59]), .Z(n1968));
Q_MX02 U3796 ( .S(n1789), .A0(n3403), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [58]), .Z(n1967));
Q_MX02 U3797 ( .S(n1789), .A0(n3404), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [57]), .Z(n1966));
Q_MX02 U3798 ( .S(n1789), .A0(n3405), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [56]), .Z(n1965));
Q_MX02 U3799 ( .S(n1789), .A0(n3406), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [55]), .Z(n1964));
Q_MX02 U3800 ( .S(n1789), .A0(n3407), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [54]), .Z(n1963));
Q_MX02 U3801 ( .S(n1789), .A0(n3408), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [53]), .Z(n1962));
Q_MX02 U3802 ( .S(n1789), .A0(n3409), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [52]), .Z(n1961));
Q_MX02 U3803 ( .S(n1789), .A0(n3410), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [51]), .Z(n1960));
Q_MX02 U3804 ( .S(n1789), .A0(n3411), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [50]), .Z(n1959));
Q_MX02 U3805 ( .S(n1789), .A0(n3412), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [49]), .Z(n1958));
Q_MX02 U3806 ( .S(n1789), .A0(n3413), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [48]), .Z(n1957));
Q_MX02 U3807 ( .S(n1789), .A0(n3414), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [47]), .Z(n1956));
Q_MX02 U3808 ( .S(n1789), .A0(n3415), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [46]), .Z(n1955));
Q_MX02 U3809 ( .S(n1789), .A0(n3416), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [45]), .Z(n1954));
Q_MX02 U3810 ( .S(n1789), .A0(n3417), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [44]), .Z(n1953));
Q_MX02 U3811 ( .S(n1789), .A0(n3418), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [43]), .Z(n1952));
Q_MX02 U3812 ( .S(n1789), .A0(n3419), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [42]), .Z(n1951));
Q_MX02 U3813 ( .S(n1789), .A0(n3420), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [41]), .Z(n1950));
Q_MX02 U3814 ( .S(n1789), .A0(n3421), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [40]), .Z(n1949));
Q_MX02 U3815 ( .S(n1789), .A0(n3422), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [39]), .Z(n1948));
Q_MX02 U3816 ( .S(n1789), .A0(n3423), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [38]), .Z(n1947));
Q_MX02 U3817 ( .S(n1789), .A0(n3424), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [37]), .Z(n1946));
Q_MX02 U3818 ( .S(n1789), .A0(n3425), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [36]), .Z(n1945));
Q_MX02 U3819 ( .S(n1789), .A0(n3426), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [35]), .Z(n1944));
Q_MX02 U3820 ( .S(n1789), .A0(n3427), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [34]), .Z(n1943));
Q_MX02 U3821 ( .S(n1789), .A0(n3428), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [33]), .Z(n1942));
Q_MX02 U3822 ( .S(n1789), .A0(n3429), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [32]), .Z(n1941));
Q_MX02 U3823 ( .S(n1789), .A0(n3430), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [31]), .Z(n1940));
Q_MX02 U3824 ( .S(n1789), .A0(n3431), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [30]), .Z(n1939));
Q_MX02 U3825 ( .S(n1789), .A0(n3432), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [29]), .Z(n1938));
Q_MX02 U3826 ( .S(n1789), .A0(n3433), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [28]), .Z(n1937));
Q_MX02 U3827 ( .S(n1789), .A0(n3434), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [27]), .Z(n1936));
Q_MX02 U3828 ( .S(n1789), .A0(n3435), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [26]), .Z(n1935));
Q_MX02 U3829 ( .S(n1789), .A0(n3436), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [25]), .Z(n1934));
Q_MX02 U3830 ( .S(n1789), .A0(n3437), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [24]), .Z(n1933));
Q_MX02 U3831 ( .S(n1789), .A0(n3438), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [23]), .Z(n1932));
Q_MX02 U3832 ( .S(n1789), .A0(n3439), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [22]), .Z(n1931));
Q_MX02 U3833 ( .S(n1789), .A0(n3440), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [21]), .Z(n1930));
Q_MX02 U3834 ( .S(n1789), .A0(n3441), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [20]), .Z(n1929));
Q_MX02 U3835 ( .S(n1789), .A0(n3442), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [19]), .Z(n1928));
Q_MX02 U3836 ( .S(n1789), .A0(n3443), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [18]), .Z(n1927));
Q_MX02 U3837 ( .S(n1789), .A0(n3444), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [17]), .Z(n1926));
Q_MX02 U3838 ( .S(n1789), .A0(n3445), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [16]), .Z(n1925));
Q_MX02 U3839 ( .S(n1789), .A0(n3446), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [15]), .Z(n1924));
Q_MX02 U3840 ( .S(n1789), .A0(n3447), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [14]), .Z(n1923));
Q_MX02 U3841 ( .S(n1789), .A0(n3448), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [13]), .Z(n1922));
Q_MX02 U3842 ( .S(n1789), .A0(n3449), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [12]), .Z(n1921));
Q_MX02 U3843 ( .S(n1789), .A0(n3450), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [11]), .Z(n1920));
Q_MX02 U3844 ( .S(n1789), .A0(n3451), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [10]), .Z(n1919));
Q_MX02 U3845 ( .S(n1789), .A0(n3452), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [9]), .Z(n1918));
Q_MX02 U3846 ( .S(n1789), .A0(n3453), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [8]), .Z(n1917));
Q_MX02 U3847 ( .S(n1789), .A0(n3454), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [7]), .Z(n1916));
Q_MX02 U3848 ( .S(n1789), .A0(n3455), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [6]), .Z(n1915));
Q_MX02 U3849 ( .S(n1789), .A0(n3456), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [5]), .Z(n1914));
Q_MX02 U3850 ( .S(n1789), .A0(n3457), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [4]), .Z(n1913));
Q_MX02 U3851 ( .S(n1789), .A0(n3458), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [3]), .Z(n1912));
Q_MX02 U3852 ( .S(n1789), .A0(n3459), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [2]), .Z(n1911));
Q_MX02 U3853 ( .S(n1789), .A0(n3460), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [1]), .Z(n1910));
Q_MX02 U3854 ( .S(n1789), .A0(n3461), .A1(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [0]), .Z(n1909));
Q_XNR2 U3855 ( .A0(_zyGfifo__gfdL496_6_P0_m2_gfOff), .A1(_zyGfifoF31_L496_req_0), .Z(n1908));
Q_XNR2 U3856 ( .A0(_zyGfifo__gfdL491_7_P0_m2_gfOff), .A1(_zyGfifoF30_L491_req_0), .Z(n1907));
Q_XNR2 U3857 ( .A0(_zyGfifo__gfdL487_8_P0_m2_gfOff), .A1(_zyGfifoF29_L487_req_0), .Z(n1906));
Q_XNR2 U3858 ( .A0(_zyGfifo__gfdL482_9_P0_m2_gfOff), .A1(_zyGfifoF28_L482_req_0), .Z(n1905));
Q_XNR2 U3859 ( .A0(_zyGfifo__gfdL480_10_P0_m2_gfOff), .A1(_zyGfifoF27_L480_req_0), .Z(n1904));
Q_XNR2 U3860 ( .A0(_zyGfifo__gfdL530_11_P0_m2_gfOff), .A1(_zyGfifoF26_L530_req_0), .Z(n1903));
Q_XNR2 U3861 ( .A0(_zyGfifo__gfdL460_12_P0_m2_gfOff), .A1(_zyGfifoF25_L460_req_0), .Z(n1902));
Q_XNR2 U3862 ( .A0(_zyGfifo__gfdL446_13_P0_m2_gfOff), .A1(_zyGfifoF24_L446_req_0), .Z(n1901));
Q_XNR2 U3863 ( .A0(_zyGfifo__gfdL444_14_P0_m2_gfOff), .A1(_zyGfifoF23_L444_req_0), .Z(n1900));
Q_XNR2 U3864 ( .A0(n1899), .A1(_zyGfifoF0_L439_s2_req_5), .Z(n3093));
Q_XNR2 U3865 ( .A0(_zyGfifo_ob_service_data_2_zyprefetch_m2_gfOff), .A1(_zyGfifoF20_L209_req_0), .Z(n1898));
Q_INV U3866 ( .A(n1897), .Z(n3549));
Q_AN02 U3867 ( .A0(n1895), .A1(n1896), .Z(n1897));
Q_AN03 U3868 ( .A0(n1887), .A1(n1886), .A2(n1894), .Z(n1896));
Q_AN03 U3869 ( .A0(n1890), .A1(n1889), .A2(n1888), .Z(n1895));
Q_AN03 U3870 ( .A0(n1893), .A1(n1892), .A2(n1891), .Z(n1894));
Q_XNR2 U3871 ( .A0(kme_ob_tstrb[7]), .A1(tstrb_ob[7]), .Z(n1893));
Q_XNR2 U3872 ( .A0(kme_ob_tstrb[6]), .A1(tstrb_ob[6]), .Z(n1892));
Q_XNR2 U3873 ( .A0(kme_ob_tstrb[5]), .A1(tstrb_ob[5]), .Z(n1891));
Q_XNR2 U3874 ( .A0(kme_ob_tstrb[4]), .A1(tstrb_ob[4]), .Z(n1890));
Q_XNR2 U3875 ( .A0(kme_ob_tstrb[3]), .A1(tstrb_ob[3]), .Z(n1889));
Q_XNR2 U3876 ( .A0(kme_ob_tstrb[2]), .A1(tstrb_ob[2]), .Z(n1888));
Q_XNR2 U3877 ( .A0(kme_ob_tstrb[1]), .A1(tstrb_ob[1]), .Z(n1887));
Q_XNR2 U3878 ( .A0(kme_ob_tstrb[0]), .A1(tstrb_ob[0]), .Z(n1886));
Q_INV U3879 ( .A(n1885), .Z(n3562));
Q_AN02 U3880 ( .A0(n1883), .A1(n1884), .Z(n1885));
Q_AN03 U3881 ( .A0(n1880), .A1(n1881), .A2(n1882), .Z(n1884));
Q_AN03 U3882 ( .A0(n1877), .A1(n1878), .A2(n1879), .Z(n1883));
Q_AN03 U3883 ( .A0(n1874), .A1(n1875), .A2(n1876), .Z(n1882));
Q_AN03 U3884 ( .A0(n1871), .A1(n1872), .A2(n1873), .Z(n1881));
Q_AN03 U3885 ( .A0(n1868), .A1(n1869), .A2(n1870), .Z(n1880));
Q_AN03 U3886 ( .A0(n1865), .A1(n1866), .A2(n1867), .Z(n1879));
Q_AN03 U3887 ( .A0(n1862), .A1(n1863), .A2(n1864), .Z(n1878));
Q_AN03 U3888 ( .A0(n1859), .A1(n1860), .A2(n1861), .Z(n1877));
Q_AN03 U3889 ( .A0(n1856), .A1(n1857), .A2(n1858), .Z(n1876));
Q_AN03 U3890 ( .A0(n1790), .A1(n1854), .A2(n1855), .Z(n1875));
Q_AN03 U3891 ( .A0(n1793), .A1(n1792), .A2(n1791), .Z(n1874));
Q_AN03 U3892 ( .A0(n1796), .A1(n1795), .A2(n1794), .Z(n1873));
Q_AN03 U3893 ( .A0(n1799), .A1(n1798), .A2(n1797), .Z(n1872));
Q_AN03 U3894 ( .A0(n1802), .A1(n1801), .A2(n1800), .Z(n1871));
Q_AN03 U3895 ( .A0(n1805), .A1(n1804), .A2(n1803), .Z(n1870));
Q_AN03 U3896 ( .A0(n1808), .A1(n1807), .A2(n1806), .Z(n1869));
Q_AN03 U3897 ( .A0(n1811), .A1(n1810), .A2(n1809), .Z(n1868));
Q_AN03 U3898 ( .A0(n1814), .A1(n1813), .A2(n1812), .Z(n1867));
Q_AN03 U3899 ( .A0(n1817), .A1(n1816), .A2(n1815), .Z(n1866));
Q_AN03 U3900 ( .A0(n1820), .A1(n1819), .A2(n1818), .Z(n1865));
Q_AN03 U3901 ( .A0(n1823), .A1(n1822), .A2(n1821), .Z(n1864));
Q_AN03 U3902 ( .A0(n1826), .A1(n1825), .A2(n1824), .Z(n1863));
Q_AN03 U3903 ( .A0(n1829), .A1(n1828), .A2(n1827), .Z(n1862));
Q_AN03 U3904 ( .A0(n1832), .A1(n1831), .A2(n1830), .Z(n1861));
Q_AN03 U3905 ( .A0(n1835), .A1(n1834), .A2(n1833), .Z(n1860));
Q_AN03 U3906 ( .A0(n1838), .A1(n1837), .A2(n1836), .Z(n1859));
Q_AN03 U3907 ( .A0(n1841), .A1(n1840), .A2(n1839), .Z(n1858));
Q_AN03 U3908 ( .A0(n1844), .A1(n1843), .A2(n1842), .Z(n1857));
Q_AN03 U3909 ( .A0(n1847), .A1(n1846), .A2(n1845), .Z(n1856));
Q_AN03 U3910 ( .A0(n1850), .A1(n1849), .A2(n1848), .Z(n1855));
Q_AN03 U3911 ( .A0(n1853), .A1(n1852), .A2(n1851), .Z(n1854));
Q_XNR2 U3912 ( .A0(kme_ob_tdata[63]), .A1(tdata_ob[63]), .Z(n1853));
Q_XNR2 U3913 ( .A0(kme_ob_tdata[62]), .A1(tdata_ob[62]), .Z(n1852));
Q_XNR2 U3914 ( .A0(kme_ob_tdata[61]), .A1(tdata_ob[61]), .Z(n1851));
Q_XNR2 U3915 ( .A0(kme_ob_tdata[60]), .A1(tdata_ob[60]), .Z(n1850));
Q_XNR2 U3916 ( .A0(kme_ob_tdata[59]), .A1(tdata_ob[59]), .Z(n1849));
Q_XNR2 U3917 ( .A0(kme_ob_tdata[58]), .A1(tdata_ob[58]), .Z(n1848));
Q_XNR2 U3918 ( .A0(kme_ob_tdata[57]), .A1(tdata_ob[57]), .Z(n1847));
Q_XNR2 U3919 ( .A0(kme_ob_tdata[56]), .A1(tdata_ob[56]), .Z(n1846));
Q_XNR2 U3920 ( .A0(kme_ob_tdata[55]), .A1(tdata_ob[55]), .Z(n1845));
Q_XNR2 U3921 ( .A0(kme_ob_tdata[54]), .A1(tdata_ob[54]), .Z(n1844));
Q_XNR2 U3922 ( .A0(kme_ob_tdata[53]), .A1(tdata_ob[53]), .Z(n1843));
Q_XNR2 U3923 ( .A0(kme_ob_tdata[52]), .A1(tdata_ob[52]), .Z(n1842));
Q_XNR2 U3924 ( .A0(kme_ob_tdata[51]), .A1(tdata_ob[51]), .Z(n1841));
Q_XNR2 U3925 ( .A0(kme_ob_tdata[50]), .A1(tdata_ob[50]), .Z(n1840));
Q_XNR2 U3926 ( .A0(kme_ob_tdata[49]), .A1(tdata_ob[49]), .Z(n1839));
Q_XNR2 U3927 ( .A0(kme_ob_tdata[48]), .A1(tdata_ob[48]), .Z(n1838));
Q_XNR2 U3928 ( .A0(kme_ob_tdata[47]), .A1(tdata_ob[47]), .Z(n1837));
Q_XNR2 U3929 ( .A0(kme_ob_tdata[46]), .A1(tdata_ob[46]), .Z(n1836));
Q_XNR2 U3930 ( .A0(kme_ob_tdata[45]), .A1(tdata_ob[45]), .Z(n1835));
Q_XNR2 U3931 ( .A0(kme_ob_tdata[44]), .A1(tdata_ob[44]), .Z(n1834));
Q_XNR2 U3932 ( .A0(kme_ob_tdata[43]), .A1(tdata_ob[43]), .Z(n1833));
Q_XNR2 U3933 ( .A0(kme_ob_tdata[42]), .A1(tdata_ob[42]), .Z(n1832));
Q_XNR2 U3934 ( .A0(kme_ob_tdata[41]), .A1(tdata_ob[41]), .Z(n1831));
Q_XNR2 U3935 ( .A0(kme_ob_tdata[40]), .A1(tdata_ob[40]), .Z(n1830));
Q_XNR2 U3936 ( .A0(kme_ob_tdata[39]), .A1(tdata_ob[39]), .Z(n1829));
Q_XNR2 U3937 ( .A0(kme_ob_tdata[38]), .A1(tdata_ob[38]), .Z(n1828));
Q_XNR2 U3938 ( .A0(kme_ob_tdata[37]), .A1(tdata_ob[37]), .Z(n1827));
Q_XNR2 U3939 ( .A0(kme_ob_tdata[36]), .A1(tdata_ob[36]), .Z(n1826));
Q_XNR2 U3940 ( .A0(kme_ob_tdata[35]), .A1(tdata_ob[35]), .Z(n1825));
Q_XNR2 U3941 ( .A0(kme_ob_tdata[34]), .A1(tdata_ob[34]), .Z(n1824));
Q_XNR2 U3942 ( .A0(kme_ob_tdata[33]), .A1(tdata_ob[33]), .Z(n1823));
Q_XNR2 U3943 ( .A0(kme_ob_tdata[32]), .A1(tdata_ob[32]), .Z(n1822));
Q_XNR2 U3944 ( .A0(kme_ob_tdata[31]), .A1(tdata_ob[31]), .Z(n1821));
Q_XNR2 U3945 ( .A0(kme_ob_tdata[30]), .A1(tdata_ob[30]), .Z(n1820));
Q_XNR2 U3946 ( .A0(kme_ob_tdata[29]), .A1(tdata_ob[29]), .Z(n1819));
Q_XNR2 U3947 ( .A0(kme_ob_tdata[28]), .A1(tdata_ob[28]), .Z(n1818));
Q_XNR2 U3948 ( .A0(kme_ob_tdata[27]), .A1(tdata_ob[27]), .Z(n1817));
Q_XNR2 U3949 ( .A0(kme_ob_tdata[26]), .A1(tdata_ob[26]), .Z(n1816));
Q_XNR2 U3950 ( .A0(kme_ob_tdata[25]), .A1(tdata_ob[25]), .Z(n1815));
Q_XNR2 U3951 ( .A0(kme_ob_tdata[24]), .A1(tdata_ob[24]), .Z(n1814));
Q_XNR2 U3952 ( .A0(kme_ob_tdata[23]), .A1(tdata_ob[23]), .Z(n1813));
Q_XNR2 U3953 ( .A0(kme_ob_tdata[22]), .A1(tdata_ob[22]), .Z(n1812));
Q_XNR2 U3954 ( .A0(kme_ob_tdata[21]), .A1(tdata_ob[21]), .Z(n1811));
Q_XNR2 U3955 ( .A0(kme_ob_tdata[20]), .A1(tdata_ob[20]), .Z(n1810));
Q_XNR2 U3956 ( .A0(kme_ob_tdata[19]), .A1(tdata_ob[19]), .Z(n1809));
Q_XNR2 U3957 ( .A0(kme_ob_tdata[18]), .A1(tdata_ob[18]), .Z(n1808));
Q_XNR2 U3958 ( .A0(kme_ob_tdata[17]), .A1(tdata_ob[17]), .Z(n1807));
Q_XNR2 U3959 ( .A0(kme_ob_tdata[16]), .A1(tdata_ob[16]), .Z(n1806));
Q_XNR2 U3960 ( .A0(kme_ob_tdata[15]), .A1(tdata_ob[15]), .Z(n1805));
Q_XNR2 U3961 ( .A0(kme_ob_tdata[14]), .A1(tdata_ob[14]), .Z(n1804));
Q_XNR2 U3962 ( .A0(kme_ob_tdata[13]), .A1(tdata_ob[13]), .Z(n1803));
Q_XNR2 U3963 ( .A0(kme_ob_tdata[12]), .A1(tdata_ob[12]), .Z(n1802));
Q_XNR2 U3964 ( .A0(kme_ob_tdata[11]), .A1(tdata_ob[11]), .Z(n1801));
Q_XNR2 U3965 ( .A0(kme_ob_tdata[10]), .A1(tdata_ob[10]), .Z(n1800));
Q_XNR2 U3966 ( .A0(kme_ob_tdata[9]), .A1(tdata_ob[9]), .Z(n1799));
Q_XNR2 U3967 ( .A0(kme_ob_tdata[8]), .A1(tdata_ob[8]), .Z(n1798));
Q_XNR2 U3968 ( .A0(kme_ob_tdata[7]), .A1(tdata_ob[7]), .Z(n1797));
Q_XNR2 U3969 ( .A0(kme_ob_tdata[6]), .A1(tdata_ob[6]), .Z(n1796));
Q_XNR2 U3970 ( .A0(kme_ob_tdata[5]), .A1(tdata_ob[5]), .Z(n1795));
Q_XNR2 U3971 ( .A0(kme_ob_tdata[4]), .A1(tdata_ob[4]), .Z(n1794));
Q_XNR2 U3972 ( .A0(kme_ob_tdata[3]), .A1(tdata_ob[3]), .Z(n1793));
Q_XNR2 U3973 ( .A0(kme_ob_tdata[2]), .A1(tdata_ob[2]), .Z(n1792));
Q_XNR2 U3974 ( .A0(kme_ob_tdata[1]), .A1(tdata_ob[1]), .Z(n1791));
Q_XNR2 U3975 ( .A0(kme_ob_tdata[0]), .A1(tdata_ob[0]), .Z(n1790));
Q_INV U3976 ( .A(n1789), .Z(n3534));
Q_AN03 U3977 ( .A0(n1784), .A1(n1783), .A2(n1788), .Z(n1789));
Q_AN03 U3978 ( .A0(n1787), .A1(n1786), .A2(n1785), .Z(n1788));
Q_XNR2 U3979 ( .A0(_zygsfis_ob_service_data_rptr[4]), .A1(_zygsfis_ob_service_data_wptr[4]), .Z(n1787));
Q_XNR2 U3980 ( .A0(_zygsfis_ob_service_data_rptr[3]), .A1(_zygsfis_ob_service_data_wptr[3]), .Z(n1786));
Q_XNR2 U3981 ( .A0(_zygsfis_ob_service_data_rptr[2]), .A1(_zygsfis_ob_service_data_wptr[2]), .Z(n1785));
Q_XNR2 U3982 ( .A0(_zygsfis_ob_service_data_rptr[1]), .A1(_zygsfis_ob_service_data_wptr[1]), .Z(n1784));
Q_XNR2 U3983 ( .A0(_zygsfis_ob_service_data_rptr[0]), .A1(_zygsfis_ob_service_data_wptr[0]), .Z(n1783));
Q_OR02 U3984 ( .A0(n1780), .A1(n1781), .Z(n1782));
Q_OR03 U3985 ( .A0(tdata_ob[1]), .A1(tdata_ob[0]), .A2(n1779), .Z(n1781));
Q_OR03 U3986 ( .A0(tdata_ob[4]), .A1(n1776), .A2(tdata_ob[2]), .Z(n1780));
Q_OR03 U3987 ( .A0(tdata_ob[7]), .A1(tdata_ob[6]), .A2(tdata_ob[5]), .Z(n1779));
Q_OR02 U3988 ( .A0(n1780), .A1(n1777), .Z(n1778));
Q_OR03 U3989 ( .A0(tdata_ob[1]), .A1(n1775), .A2(n1779), .Z(n1777));
Q_INV U3990 ( .A(n1774), .Z(n3545));
Q_OR02 U3991 ( .A0(n1772), .A1(n1773), .Z(n1774));
Q_OR03 U3992 ( .A0(n1769), .A1(n1770), .A2(n1771), .Z(n1773));
Q_OR03 U3993 ( .A0(n1766), .A1(n1767), .A2(n1768), .Z(n1772));
Q_OR03 U3994 ( .A0(n1763), .A1(n1764), .A2(n1765), .Z(n1771));
Q_OR03 U3995 ( .A0(n1760), .A1(n1761), .A2(n1762), .Z(n1770));
Q_OR03 U3996 ( .A0(n1758), .A1(n1757), .A2(n1759), .Z(n1769));
Q_OR03 U3997 ( .A0(str_get_ob[4]), .A1(str_get_ob[3]), .A2(str_get_ob[2]), .Z(n1768));
Q_OR03 U3998 ( .A0(str_get_ob[7]), .A1(str_get_ob[6]), .A2(str_get_ob[5]), .Z(n1767));
Q_OR03 U3999 ( .A0(str_get_ob[10]), .A1(str_get_ob[9]), .A2(str_get_ob[8]), .Z(n1766));
Q_OR03 U4000 ( .A0(str_get_ob[13]), .A1(str_get_ob[12]), .A2(str_get_ob[11]), .Z(n1765));
Q_OR03 U4001 ( .A0(str_get_ob[16]), .A1(str_get_ob[15]), .A2(str_get_ob[14]), .Z(n1764));
Q_OR03 U4002 ( .A0(str_get_ob[19]), .A1(str_get_ob[18]), .A2(str_get_ob[17]), .Z(n1763));
Q_OR03 U4003 ( .A0(str_get_ob[22]), .A1(str_get_ob[21]), .A2(str_get_ob[20]), .Z(n1762));
Q_OR03 U4004 ( .A0(str_get_ob[25]), .A1(str_get_ob[24]), .A2(str_get_ob[23]), .Z(n1761));
Q_OR03 U4005 ( .A0(str_get_ob[28]), .A1(str_get_ob[27]), .A2(str_get_ob[26]), .Z(n1760));
Q_OR03 U4006 ( .A0(str_get_ob[31]), .A1(str_get_ob[30]), .A2(str_get_ob[29]), .Z(n1759));
Q_AN03 U4007 ( .A0(n1752), .A1(n1751), .A2(n1756), .Z(n3535));
Q_AN03 U4008 ( .A0(n1755), .A1(n1754), .A2(n1753), .Z(n1756));
Q_XNR2 U4009 ( .A0(_zygsfis_ob_service_data_req[4]), .A1(_zygsfis_ob_service_data_ack[4]), .Z(n1755));
Q_XNR2 U4010 ( .A0(_zygsfis_ob_service_data_req[3]), .A1(_zygsfis_ob_service_data_ack[3]), .Z(n1754));
Q_XNR2 U4011 ( .A0(_zygsfis_ob_service_data_req[2]), .A1(_zygsfis_ob_service_data_ack[2]), .Z(n1753));
Q_XNR2 U4012 ( .A0(_zygsfis_ob_service_data_req[1]), .A1(_zygsfis_ob_service_data_ack[1]), .Z(n1752));
Q_XNR2 U4013 ( .A0(_zygsfis_ob_service_data_req[0]), .A1(_zygsfis_ob_service_data_ack[0]), .Z(n1751));
Q_OR02 U4014 ( .A0(n1481), .A1(n445), .Z(n1749));
Q_NR02 U4015 ( .A0(n445), .A1(mega_tlv_word_count[0]), .Z(n1748));
Q_AN02 U4016 ( .A0(n442), .A1(n1173), .Z(n1746));
Q_AN02 U4017 ( .A0(n442), .A1(n1175), .Z(n1745));
Q_AN02 U4018 ( .A0(n442), .A1(n1177), .Z(n1744));
Q_AN02 U4019 ( .A0(n442), .A1(n1179), .Z(n1743));
Q_AN02 U4020 ( .A0(n442), .A1(n1181), .Z(n1742));
Q_AN02 U4021 ( .A0(n442), .A1(n1183), .Z(n1741));
Q_AN02 U4022 ( .A0(n442), .A1(n1185), .Z(n1740));
Q_AN02 U4023 ( .A0(n442), .A1(n1187), .Z(n1739));
Q_AN02 U4024 ( .A0(n442), .A1(n1189), .Z(n1738));
Q_AN02 U4025 ( .A0(n442), .A1(n1191), .Z(n1737));
Q_AN02 U4026 ( .A0(n442), .A1(n1193), .Z(n1736));
Q_AN02 U4027 ( .A0(n442), .A1(n1195), .Z(n1735));
Q_AN02 U4028 ( .A0(n442), .A1(n1197), .Z(n1734));
Q_AN02 U4029 ( .A0(n442), .A1(n1199), .Z(n1733));
Q_AN02 U4030 ( .A0(n442), .A1(n1201), .Z(n1732));
Q_AN02 U4031 ( .A0(n442), .A1(n1203), .Z(n1731));
Q_AN02 U4032 ( .A0(n442), .A1(n1205), .Z(n1730));
Q_AN02 U4033 ( .A0(n442), .A1(n1207), .Z(n1729));
Q_AN02 U4034 ( .A0(n442), .A1(n1209), .Z(n1728));
Q_AN02 U4035 ( .A0(n442), .A1(n1211), .Z(n1727));
Q_AN02 U4036 ( .A0(n442), .A1(n1213), .Z(n1726));
Q_AN02 U4037 ( .A0(n442), .A1(n1215), .Z(n1725));
Q_AN02 U4038 ( .A0(n442), .A1(n1217), .Z(n1724));
Q_AN02 U4039 ( .A0(n442), .A1(n1219), .Z(n1723));
Q_AN02 U4040 ( .A0(n442), .A1(n1221), .Z(n1722));
Q_AN02 U4041 ( .A0(n442), .A1(n1223), .Z(n1721));
Q_AN02 U4042 ( .A0(n442), .A1(n1225), .Z(n1720));
Q_AN02 U4043 ( .A0(n442), .A1(n1227), .Z(n1719));
Q_AN02 U4044 ( .A0(n442), .A1(n1229), .Z(n1718));
Q_AN02 U4045 ( .A0(n442), .A1(n1231), .Z(n1717));
Q_AN02 U4046 ( .A0(n442), .A1(n1233), .Z(n1716));
Q_OR02 U4047 ( .A0(n1640), .A1(n445), .Z(n1715));
Q_AN02 U4048 ( .A0(n442), .A1(n1711), .Z(n1714));
Q_AN02 U4049 ( .A0(n442), .A1(n1433), .Z(n1713));
Q_AN02 U4050 ( .A0(n442), .A1(n1434), .Z(n1712));
Q_OR02 U4051 ( .A0(n1492), .A1(_zyL368_meState4[0]), .Z(n1484));
Q_ND02 U4052 ( .A0(n1643), .A1(kme_ib_tready), .Z(n1491));
Q_INV U4053 ( .A(n1643), .Z(n1487));
Q_OR02 U4054 ( .A0(n1491), .A1(n1484), .Z(n1490));
Q_OR02 U4055 ( .A0(n1432), .A1(n1490), .Z(n1482));
Q_INV U4056 ( .A(n1482), .Z(n1640));
Q_INV U4057 ( .A(n1490), .Z(n1635));
Q_OR03 U4058 ( .A0(n1474), .A1(n1250), .A2(n1482), .Z(n1489));
Q_INV U4059 ( .A(n1709), .Z(n1474));
Q_OR02 U4060 ( .A0(n1633), .A1(n1482), .Z(n1488));
Q_NR02 U4061 ( .A0(n1487), .A1(n1484), .Z(n1638));
Q_OR02 U4062 ( .A0(n1374), .A1(n1484), .Z(n1486));
Q_MX02 U4063 ( .S(n1358), .A0(n1484), .A1(n1486), .Z(n1485));
Q_OR03 U4064 ( .A0(n1305), .A1(n1639), .A2(n1484), .Z(n1483));
Q_INV U4065 ( .A(n1483), .Z(n1641));
Q_NR02 U4066 ( .A0(n1474), .A1(n1482), .Z(n1481));
Q_OR02 U4067 ( .A0(n1642), .A1(n1639), .Z(n1480));
Q_NR02 U4068 ( .A0(n1374), .A1(n1432), .Z(n1479));
Q_ND02 U4069 ( .A0(n1358), .A1(n1479), .Z(n1477));
Q_OR02 U4070 ( .A0(n1711), .A1(n1477), .Z(n1478));
Q_INV U4071 ( .A(n1710), .Z(n1473));
Q_OR02 U4072 ( .A0(n1473), .A1(n1477), .Z(n1476));
Q_MX02 U4073 ( .S(n1709), .A0(n1476), .A1(n1478), .Z(n1475));
Q_INV U4074 ( .A(n1475), .Z(n1637));
Q_OR02 U4075 ( .A0(n1632), .A1(n1374), .Z(n1471));
Q_OA21 U4076 ( .A0(n1474), .A1(n1471), .B0(n1709), .Z(n1434));
Q_OR02 U4077 ( .A0(n1709), .A1(n1473), .Z(n1472));
Q_OA21 U4078 ( .A0(n1472), .A1(n1471), .B0(n1710), .Z(n1433));
Q_INV U4079 ( .A(n1471), .Z(n1631));
Q_AN03 U4080 ( .A0(n1649), .A1(n1644), .A2(n1709), .Z(n1470));
Q_NR02 U4081 ( .A0(n1320), .A1(n1358), .Z(n1469));
Q_INV U4082 ( .A(n1469), .Z(n1633));
Q_AN02 U4083 ( .A0(n1636), .A1(n1358), .Z(n1468));
Q_AN02 U4084 ( .A0(n1636), .A1(n1471), .Z(n1467));
Q_NR02 U4085 ( .A0(n1164), .A1(n1639), .Z(n1643));
Q_FDP0 _zzM2L368_mdxP3_kme_ib_tuser_Dwen4_REG  ( .CK(clk), .D(n1635), .Q(_zzM2L368_mdxP3_kme_ib_tuser_Dwen4), .QN( ));
Q_FDP0 _zzM2L368_mdxP3_kme_ib_tstrb_Dwen3_REG  ( .CK(clk), .D(n1635), .Q(_zzM2L368_mdxP3_kme_ib_tstrb_Dwen3), .QN( ));
Q_FDP0 _zzM2L368_mdxP3_kme_ib_tdata_Dwen2_REG  ( .CK(clk), .D(n1635), .Q(_zzM2L368_mdxP3_kme_ib_tdata_Dwen2), .QN( ));
Q_FDP0 _zzM2L368_mdxP3_kme_ib_tlast_Dwen1_REG  ( .CK(clk), .D(n1635), .Q(_zzM2L368_mdxP3_kme_ib_tlast_Dwen1), .QN( ));
Q_FDP0 _zzM2L368_mdxP3_kme_ib_tvalid_Dwen0_REG  ( .CK(clk), .D(n1635), .Q(_zzM2L368_mdxP3_kme_ib_tvalid_Dwen0), .QN( ));
Q_FDP0 \_zyL368_meState4_REG[0] ( .CK(clk), .D(n1638), .Q(_zyL368_meState4[0]), .QN( ));
Q_XNR2 U4092 ( .A0(n1631), .A1(n1358), .Z(n1466));
Q_MX02 U4093 ( .S(n1480), .A0(n1304), .A1(n1464), .Z(n1465));
Q_AN02 U4094 ( .A0(n1639), .A1(n1299), .Z(n1464));
Q_MX02 U4095 ( .S(n1480), .A0(n1303), .A1(n1462), .Z(n1463));
Q_AN02 U4096 ( .A0(n1639), .A1(n1298), .Z(n1462));
Q_MX02 U4097 ( .S(n1480), .A0(n1302), .A1(n1460), .Z(n1461));
Q_AN02 U4098 ( .A0(n1639), .A1(n1297), .Z(n1460));
Q_MX02 U4099 ( .S(n1480), .A0(n1301), .A1(n1458), .Z(n1459));
Q_AN02 U4100 ( .A0(n1639), .A1(n1296), .Z(n1458));
Q_MX02 U4101 ( .S(n1480), .A0(n1300), .A1(n1456), .Z(n1457));
Q_AN02 U4102 ( .A0(n1639), .A1(n1295), .Z(n1456));
Q_MX02 U4103 ( .S(n1358), .A0(_zyGfifo__gfdL519_24_P0_m2_gfOff), .A1(_zyGfifo__gfdL522_23_P0_m2_gfOff), .Z(n1166));
Q_MX02 U4104 ( .S(n1358), .A0(_zyGfifo__gfdL519_24_P0_m2_cbid[19]), .A1(_zyGfifo__gfdL522_23_P0_m2_cbid[19]), .Z(n1454));
Q_MX02 U4105 ( .S(n1358), .A0(_zyGfifo__gfdL519_24_P0_m2_cbid[18]), .A1(_zyGfifo__gfdL522_23_P0_m2_cbid[18]), .Z(n1453));
Q_MX02 U4106 ( .S(n1358), .A0(_zyGfifo__gfdL519_24_P0_m2_cbid[17]), .A1(_zyGfifo__gfdL522_23_P0_m2_cbid[17]), .Z(n1452));
Q_MX02 U4107 ( .S(n1358), .A0(_zyGfifo__gfdL519_24_P0_m2_cbid[16]), .A1(_zyGfifo__gfdL522_23_P0_m2_cbid[16]), .Z(n1451));
Q_MX02 U4108 ( .S(n1358), .A0(_zyGfifo__gfdL519_24_P0_m2_cbid[15]), .A1(_zyGfifo__gfdL522_23_P0_m2_cbid[15]), .Z(n1450));
Q_MX02 U4109 ( .S(n1358), .A0(_zyGfifo__gfdL519_24_P0_m2_cbid[14]), .A1(_zyGfifo__gfdL522_23_P0_m2_cbid[14]), .Z(n1449));
Q_MX02 U4110 ( .S(n1358), .A0(_zyGfifo__gfdL519_24_P0_m2_cbid[13]), .A1(_zyGfifo__gfdL522_23_P0_m2_cbid[13]), .Z(n1448));
Q_MX02 U4111 ( .S(n1358), .A0(_zyGfifo__gfdL519_24_P0_m2_cbid[12]), .A1(_zyGfifo__gfdL522_23_P0_m2_cbid[12]), .Z(n1447));
Q_MX02 U4112 ( .S(n1358), .A0(_zyGfifo__gfdL519_24_P0_m2_cbid[11]), .A1(_zyGfifo__gfdL522_23_P0_m2_cbid[11]), .Z(n1446));
Q_MX02 U4113 ( .S(n1358), .A0(_zyGfifo__gfdL519_24_P0_m2_cbid[10]), .A1(_zyGfifo__gfdL522_23_P0_m2_cbid[10]), .Z(n1445));
Q_MX02 U4114 ( .S(n1358), .A0(_zyGfifo__gfdL519_24_P0_m2_cbid[9]), .A1(_zyGfifo__gfdL522_23_P0_m2_cbid[9]), .Z(n1444));
Q_MX02 U4115 ( .S(n1358), .A0(_zyGfifo__gfdL519_24_P0_m2_cbid[8]), .A1(_zyGfifo__gfdL522_23_P0_m2_cbid[8]), .Z(n1443));
Q_MX02 U4116 ( .S(n1358), .A0(_zyGfifo__gfdL519_24_P0_m2_cbid[7]), .A1(_zyGfifo__gfdL522_23_P0_m2_cbid[7]), .Z(n1442));
Q_MX02 U4117 ( .S(n1358), .A0(_zyGfifo__gfdL519_24_P0_m2_cbid[6]), .A1(_zyGfifo__gfdL522_23_P0_m2_cbid[6]), .Z(n1441));
Q_MX02 U4118 ( .S(n1358), .A0(_zyGfifo__gfdL519_24_P0_m2_cbid[5]), .A1(_zyGfifo__gfdL522_23_P0_m2_cbid[5]), .Z(n1440));
Q_MX02 U4119 ( .S(n1358), .A0(_zyGfifo__gfdL519_24_P0_m2_cbid[4]), .A1(_zyGfifo__gfdL522_23_P0_m2_cbid[4]), .Z(n1439));
Q_MX02 U4120 ( .S(n1358), .A0(_zyGfifo__gfdL519_24_P0_m2_cbid[3]), .A1(_zyGfifo__gfdL522_23_P0_m2_cbid[3]), .Z(n1438));
Q_MX02 U4121 ( .S(n1358), .A0(_zyGfifo__gfdL519_24_P0_m2_cbid[2]), .A1(_zyGfifo__gfdL522_23_P0_m2_cbid[2]), .Z(n1437));
Q_MX02 U4122 ( .S(n1358), .A0(_zyGfifo__gfdL519_24_P0_m2_cbid[1]), .A1(_zyGfifo__gfdL522_23_P0_m2_cbid[1]), .Z(n1436));
Q_MX02 U4123 ( .S(n1358), .A0(_zyGfifo__gfdL519_24_P0_m2_cbid[0]), .A1(_zyGfifo__gfdL522_23_P0_m2_cbid[0]), .Z(n1435));
Q_OR02 U4124 ( .A0(n1470), .A1(have_guid_tlv), .Z(n1711));
Q_OR02 U4125 ( .A0(n1634), .A1(saw_guid_tlv), .Z(n1710));
Q_OR02 U4126 ( .A0(n1469), .A1(saw_mega), .Z(n1709));
Q_INV U4127 ( .A(n1432), .Z(n1636));
Q_OR02 U4128 ( .A0(n1430), .A1(n1431), .Z(n1432));
Q_OR03 U4129 ( .A0(n1427), .A1(n1428), .A2(n1429), .Z(n1431));
Q_OR03 U4130 ( .A0(n1424), .A1(n1425), .A2(n1426), .Z(n1430));
Q_OR03 U4131 ( .A0(n1421), .A1(n1422), .A2(n1423), .Z(n1429));
Q_OR03 U4132 ( .A0(n1418), .A1(n1419), .A2(n1420), .Z(n1428));
Q_OR03 U4133 ( .A0(n1416), .A1(n1415), .A2(n1417), .Z(n1427));
Q_OR03 U4134 ( .A0(n1387), .A1(n1386), .A2(n1385), .Z(n1426));
Q_OR03 U4135 ( .A0(n1390), .A1(n1389), .A2(n1388), .Z(n1425));
Q_OR03 U4136 ( .A0(n1393), .A1(n1392), .A2(n1391), .Z(n1424));
Q_OR03 U4137 ( .A0(n1396), .A1(n1395), .A2(n1394), .Z(n1423));
Q_OR03 U4138 ( .A0(n1399), .A1(n1398), .A2(n1397), .Z(n1422));
Q_OR03 U4139 ( .A0(n1402), .A1(n1401), .A2(n1400), .Z(n1421));
Q_OR03 U4140 ( .A0(n1405), .A1(n1404), .A2(n1403), .Z(n1420));
Q_OR03 U4141 ( .A0(n1408), .A1(n1407), .A2(n1406), .Z(n1419));
Q_OR03 U4142 ( .A0(n1411), .A1(n1410), .A2(n1409), .Z(n1418));
Q_OR03 U4143 ( .A0(n1414), .A1(n1413), .A2(n1412), .Z(n1417));
Q_INV U4144 ( .A(n1384), .Z(n1416));
Q_INV U4145 ( .A(n1383), .Z(n1415));
Q_MX02 U4146 ( .S(n1164), .A0(n1597), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [31]), .Z(n1414));
Q_MX02 U4147 ( .S(n1164), .A0(n1598), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [30]), .Z(n1413));
Q_MX02 U4148 ( .S(n1164), .A0(n1599), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [29]), .Z(n1412));
Q_MX02 U4149 ( .S(n1164), .A0(n1600), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [28]), .Z(n1411));
Q_MX02 U4150 ( .S(n1164), .A0(n1601), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [27]), .Z(n1410));
Q_MX02 U4151 ( .S(n1164), .A0(n1602), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [26]), .Z(n1409));
Q_MX02 U4152 ( .S(n1164), .A0(n1603), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [25]), .Z(n1408));
Q_MX02 U4153 ( .S(n1164), .A0(n1604), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [24]), .Z(n1407));
Q_MX02 U4154 ( .S(n1164), .A0(n1605), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [23]), .Z(n1406));
Q_MX02 U4155 ( .S(n1164), .A0(n1606), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [22]), .Z(n1405));
Q_MX02 U4156 ( .S(n1164), .A0(n1607), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [21]), .Z(n1404));
Q_MX02 U4157 ( .S(n1164), .A0(n1608), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [20]), .Z(n1403));
Q_MX02 U4158 ( .S(n1164), .A0(n1609), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [19]), .Z(n1402));
Q_MX02 U4159 ( .S(n1164), .A0(n1610), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [18]), .Z(n1401));
Q_MX02 U4160 ( .S(n1164), .A0(n1611), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [17]), .Z(n1400));
Q_MX02 U4161 ( .S(n1164), .A0(n1612), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [16]), .Z(n1399));
Q_MX02 U4162 ( .S(n1164), .A0(n1613), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [15]), .Z(n1398));
Q_MX02 U4163 ( .S(n1164), .A0(n1614), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [14]), .Z(n1397));
Q_MX02 U4164 ( .S(n1164), .A0(n1615), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [13]), .Z(n1396));
Q_MX02 U4165 ( .S(n1164), .A0(n1616), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [12]), .Z(n1395));
Q_MX02 U4166 ( .S(n1164), .A0(n1617), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [11]), .Z(n1394));
Q_MX02 U4167 ( .S(n1164), .A0(n1618), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [10]), .Z(n1393));
Q_MX02 U4168 ( .S(n1164), .A0(n1619), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [9]), .Z(n1392));
Q_MX02 U4169 ( .S(n1164), .A0(n1620), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [8]), .Z(n1391));
Q_MX02 U4170 ( .S(n1164), .A0(n1621), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [7]), .Z(n1390));
Q_MX02 U4171 ( .S(n1164), .A0(n1622), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [6]), .Z(n1389));
Q_MX02 U4172 ( .S(n1164), .A0(n1623), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [5]), .Z(n1388));
Q_MX02 U4173 ( .S(n1164), .A0(n1624), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [4]), .Z(n1387));
Q_MX02 U4174 ( .S(n1164), .A0(n1625), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [3]), .Z(n1386));
Q_MX02 U4175 ( .S(n1164), .A0(n1626), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [2]), .Z(n1385));
Q_MX02 U4176 ( .S(n1164), .A0(n1627), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [1]), .Z(n1384));
Q_MX02 U4177 ( .S(n1164), .A0(n1628), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [0]), .Z(n1383));
Q_MX02 U4178 ( .S(n1164), .A0(n1589), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytstrb_L207_tfiV7 [7]), .Z(n1382));
Q_MX02 U4179 ( .S(n1164), .A0(n1590), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytstrb_L207_tfiV7 [6]), .Z(n1381));
Q_MX02 U4180 ( .S(n1164), .A0(n1591), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytstrb_L207_tfiV7 [5]), .Z(n1380));
Q_MX02 U4181 ( .S(n1164), .A0(n1592), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytstrb_L207_tfiV7 [4]), .Z(n1379));
Q_MX02 U4182 ( .S(n1164), .A0(n1593), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytstrb_L207_tfiV7 [3]), .Z(n1378));
Q_MX02 U4183 ( .S(n1164), .A0(n1594), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytstrb_L207_tfiV7 [2]), .Z(n1377));
Q_MX02 U4184 ( .S(n1164), .A0(n1595), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytstrb_L207_tfiV7 [1]), .Z(n1376));
Q_MX02 U4185 ( .S(n1164), .A0(n1596), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytstrb_L207_tfiV7 [0]), .Z(n1375));
Q_OR02 U4186 ( .A0(n1372), .A1(n1373), .Z(n1374));
Q_OR03 U4187 ( .A0(n1369), .A1(n1370), .A2(n1371), .Z(n1373));
Q_OR03 U4188 ( .A0(n1366), .A1(n1367), .A2(n1368), .Z(n1372));
Q_OR03 U4189 ( .A0(n1363), .A1(n1364), .A2(n1365), .Z(n1371));
Q_OR03 U4190 ( .A0(n1360), .A1(n1361), .A2(n1362), .Z(n1370));
Q_OR03 U4191 ( .A0(n1354), .A1(n1321), .A2(n1359), .Z(n1369));
Q_OR03 U4192 ( .A0(n1325), .A1(n1355), .A2(n1323), .Z(n1368));
Q_OR03 U4193 ( .A0(n1328), .A1(n1327), .A2(n1326), .Z(n1367));
Q_OR03 U4194 ( .A0(n1331), .A1(n1330), .A2(n1329), .Z(n1366));
Q_OR03 U4195 ( .A0(n1334), .A1(n1333), .A2(n1332), .Z(n1365));
Q_OR03 U4196 ( .A0(n1337), .A1(n1336), .A2(n1335), .Z(n1364));
Q_OR03 U4197 ( .A0(n1340), .A1(n1339), .A2(n1338), .Z(n1363));
Q_OR03 U4198 ( .A0(n1343), .A1(n1342), .A2(n1341), .Z(n1362));
Q_OR03 U4199 ( .A0(n1346), .A1(n1345), .A2(n1344), .Z(n1361));
Q_OR03 U4200 ( .A0(n1349), .A1(n1348), .A2(n1347), .Z(n1360));
Q_OR03 U4201 ( .A0(n1352), .A1(n1351), .A2(n1350), .Z(n1359));
Q_INV U4202 ( .A(n1358), .Z(n1632));
Q_OR02 U4203 ( .A0(n1372), .A1(n1357), .Z(n1358));
Q_OR03 U4204 ( .A0(n1356), .A1(n1370), .A2(n1371), .Z(n1357));
Q_OR03 U4205 ( .A0(n1354), .A1(n1353), .A2(n1359), .Z(n1356));
Q_INV U4206 ( .A(n1324), .Z(n1355));
Q_INV U4207 ( .A(n1322), .Z(n1354));
Q_INV U4208 ( .A(n1321), .Z(n1353));
Q_MX02 U4209 ( .S(n1164), .A0(n1557), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [31]), .Z(n1352));
Q_MX02 U4210 ( .S(n1164), .A0(n1558), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [30]), .Z(n1351));
Q_MX02 U4211 ( .S(n1164), .A0(n1559), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [29]), .Z(n1350));
Q_MX02 U4212 ( .S(n1164), .A0(n1560), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [28]), .Z(n1349));
Q_MX02 U4213 ( .S(n1164), .A0(n1561), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [27]), .Z(n1348));
Q_MX02 U4214 ( .S(n1164), .A0(n1562), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [26]), .Z(n1347));
Q_MX02 U4215 ( .S(n1164), .A0(n1563), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [25]), .Z(n1346));
Q_MX02 U4216 ( .S(n1164), .A0(n1564), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [24]), .Z(n1345));
Q_MX02 U4217 ( .S(n1164), .A0(n1565), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [23]), .Z(n1344));
Q_MX02 U4218 ( .S(n1164), .A0(n1566), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [22]), .Z(n1343));
Q_MX02 U4219 ( .S(n1164), .A0(n1567), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [21]), .Z(n1342));
Q_MX02 U4220 ( .S(n1164), .A0(n1568), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [20]), .Z(n1341));
Q_MX02 U4221 ( .S(n1164), .A0(n1569), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [19]), .Z(n1340));
Q_MX02 U4222 ( .S(n1164), .A0(n1570), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [18]), .Z(n1339));
Q_MX02 U4223 ( .S(n1164), .A0(n1571), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [17]), .Z(n1338));
Q_MX02 U4224 ( .S(n1164), .A0(n1572), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [16]), .Z(n1337));
Q_MX02 U4225 ( .S(n1164), .A0(n1573), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [15]), .Z(n1336));
Q_MX02 U4226 ( .S(n1164), .A0(n1574), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [14]), .Z(n1335));
Q_MX02 U4227 ( .S(n1164), .A0(n1575), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [13]), .Z(n1334));
Q_MX02 U4228 ( .S(n1164), .A0(n1576), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [12]), .Z(n1333));
Q_MX02 U4229 ( .S(n1164), .A0(n1577), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [11]), .Z(n1332));
Q_MX02 U4230 ( .S(n1164), .A0(n1578), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [10]), .Z(n1331));
Q_MX02 U4231 ( .S(n1164), .A0(n1579), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [9]), .Z(n1330));
Q_MX02 U4232 ( .S(n1164), .A0(n1580), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [8]), .Z(n1329));
Q_MX02 U4233 ( .S(n1164), .A0(n1581), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [7]), .Z(n1328));
Q_MX02 U4234 ( .S(n1164), .A0(n1582), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [6]), .Z(n1327));
Q_MX02 U4235 ( .S(n1164), .A0(n1583), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [5]), .Z(n1326));
Q_MX02 U4236 ( .S(n1164), .A0(n1584), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [4]), .Z(n1325));
Q_MX02 U4237 ( .S(n1164), .A0(n1585), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [3]), .Z(n1324));
Q_MX02 U4238 ( .S(n1164), .A0(n1586), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [2]), .Z(n1323));
Q_MX02 U4239 ( .S(n1164), .A0(n1587), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [1]), .Z(n1322));
Q_MX02 U4240 ( .S(n1164), .A0(n1588), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [0]), .Z(n1321));
Q_AO21 U4241 ( .A0(n1314), .A1(n1319), .B0(n1315), .Z(n1320));
Q_NR02 U4242 ( .A0(n1648), .A1(n1647), .Z(n1318));
Q_AO21 U4243 ( .A0(n1317), .A1(n1316), .B0(n1318), .Z(n1319));
Q_NR02 U4244 ( .A0(n1648), .A1(n1646), .Z(n1317));
Q_INV U4245 ( .A(n1645), .Z(n1316));
Q_AN02 U4246 ( .A0(n1314), .A1(n1312), .Z(n1315));
Q_AN02 U4247 ( .A0(n1313), .A1(n1311), .Z(n1314));
Q_NR02 U4248 ( .A0(n1652), .A1(n1651), .Z(n1313));
Q_INV U4249 ( .A(n1649), .Z(n1312));
Q_INV U4250 ( .A(n1650), .Z(n1311));
Q_NR03 U4251 ( .A0(n1309), .A1(n1310), .A2(n1469), .Z(n1634));
Q_OR03 U4252 ( .A0(n1306), .A1(n1645), .A2(n1308), .Z(n1310));
Q_OR03 U4253 ( .A0(n1649), .A1(n1307), .A2(n1647), .Z(n1309));
Q_OR03 U4254 ( .A0(n1652), .A1(n1651), .A2(n1650), .Z(n1308));
Q_INV U4255 ( .A(n1648), .Z(n1307));
Q_INV U4256 ( .A(n1646), .Z(n1306));
Q_MX02 U4257 ( .S(n1164), .A0(n1493), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [63]), .Z(n1708));
Q_MX02 U4258 ( .S(n1164), .A0(n1494), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [62]), .Z(n1707));
Q_MX02 U4259 ( .S(n1164), .A0(n1495), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [61]), .Z(n1706));
Q_MX02 U4260 ( .S(n1164), .A0(n1496), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [60]), .Z(n1705));
Q_MX02 U4261 ( .S(n1164), .A0(n1497), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [59]), .Z(n1704));
Q_MX02 U4262 ( .S(n1164), .A0(n1498), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [58]), .Z(n1703));
Q_MX02 U4263 ( .S(n1164), .A0(n1499), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [57]), .Z(n1702));
Q_MX02 U4264 ( .S(n1164), .A0(n1500), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [56]), .Z(n1701));
Q_MX02 U4265 ( .S(n1164), .A0(n1501), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [55]), .Z(n1700));
Q_MX02 U4266 ( .S(n1164), .A0(n1502), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [54]), .Z(n1699));
Q_MX02 U4267 ( .S(n1164), .A0(n1503), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [53]), .Z(n1698));
Q_MX02 U4268 ( .S(n1164), .A0(n1504), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [52]), .Z(n1697));
Q_MX02 U4269 ( .S(n1164), .A0(n1505), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [51]), .Z(n1696));
Q_MX02 U4270 ( .S(n1164), .A0(n1506), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [50]), .Z(n1695));
Q_MX02 U4271 ( .S(n1164), .A0(n1507), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [49]), .Z(n1694));
Q_MX02 U4272 ( .S(n1164), .A0(n1508), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [48]), .Z(n1693));
Q_MX02 U4273 ( .S(n1164), .A0(n1509), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [47]), .Z(n1692));
Q_MX02 U4274 ( .S(n1164), .A0(n1510), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [46]), .Z(n1691));
Q_MX02 U4275 ( .S(n1164), .A0(n1511), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [45]), .Z(n1690));
Q_MX02 U4276 ( .S(n1164), .A0(n1512), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [44]), .Z(n1689));
Q_MX02 U4277 ( .S(n1164), .A0(n1513), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [43]), .Z(n1688));
Q_MX02 U4278 ( .S(n1164), .A0(n1514), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [42]), .Z(n1687));
Q_MX02 U4279 ( .S(n1164), .A0(n1515), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [41]), .Z(n1686));
Q_MX02 U4280 ( .S(n1164), .A0(n1516), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [40]), .Z(n1685));
Q_MX02 U4281 ( .S(n1164), .A0(n1517), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [39]), .Z(n1684));
Q_MX02 U4282 ( .S(n1164), .A0(n1518), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [38]), .Z(n1683));
Q_MX02 U4283 ( .S(n1164), .A0(n1519), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [37]), .Z(n1682));
Q_MX02 U4284 ( .S(n1164), .A0(n1520), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [36]), .Z(n1681));
Q_MX02 U4285 ( .S(n1164), .A0(n1521), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [35]), .Z(n1680));
Q_MX02 U4286 ( .S(n1164), .A0(n1522), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [34]), .Z(n1679));
Q_MX02 U4287 ( .S(n1164), .A0(n1523), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [33]), .Z(n1678));
Q_MX02 U4288 ( .S(n1164), .A0(n1524), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [32]), .Z(n1677));
Q_MX02 U4289 ( .S(n1164), .A0(n1525), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [31]), .Z(n1676));
Q_MX02 U4290 ( .S(n1164), .A0(n1526), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [30]), .Z(n1675));
Q_MX02 U4291 ( .S(n1164), .A0(n1527), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [29]), .Z(n1674));
Q_MX02 U4292 ( .S(n1164), .A0(n1528), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [28]), .Z(n1673));
Q_MX02 U4293 ( .S(n1164), .A0(n1529), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [27]), .Z(n1672));
Q_MX02 U4294 ( .S(n1164), .A0(n1530), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [26]), .Z(n1671));
Q_MX02 U4295 ( .S(n1164), .A0(n1531), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [25]), .Z(n1670));
Q_MX02 U4296 ( .S(n1164), .A0(n1532), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [24]), .Z(n1669));
Q_MX02 U4297 ( .S(n1164), .A0(n1533), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [23]), .Z(n1668));
Q_MX02 U4298 ( .S(n1164), .A0(n1534), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [22]), .Z(n1667));
Q_MX02 U4299 ( .S(n1164), .A0(n1535), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [21]), .Z(n1666));
Q_MX02 U4300 ( .S(n1164), .A0(n1536), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [20]), .Z(n1665));
Q_MX02 U4301 ( .S(n1164), .A0(n1537), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [19]), .Z(n1664));
Q_MX02 U4302 ( .S(n1164), .A0(n1538), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [18]), .Z(n1663));
Q_MX02 U4303 ( .S(n1164), .A0(n1539), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [17]), .Z(n1662));
Q_MX02 U4304 ( .S(n1164), .A0(n1540), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [16]), .Z(n1661));
Q_MX02 U4305 ( .S(n1164), .A0(n1541), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [15]), .Z(n1660));
Q_MX02 U4306 ( .S(n1164), .A0(n1542), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [14]), .Z(n1659));
Q_MX02 U4307 ( .S(n1164), .A0(n1543), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [13]), .Z(n1658));
Q_MX02 U4308 ( .S(n1164), .A0(n1544), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [12]), .Z(n1657));
Q_MX02 U4309 ( .S(n1164), .A0(n1545), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [11]), .Z(n1656));
Q_MX02 U4310 ( .S(n1164), .A0(n1546), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [10]), .Z(n1655));
Q_MX02 U4311 ( .S(n1164), .A0(n1547), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [9]), .Z(n1654));
Q_MX02 U4312 ( .S(n1164), .A0(n1548), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [8]), .Z(n1653));
Q_MX02 U4313 ( .S(n1164), .A0(n1549), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [7]), .Z(n1652));
Q_MX02 U4314 ( .S(n1164), .A0(n1550), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [6]), .Z(n1651));
Q_MX02 U4315 ( .S(n1164), .A0(n1551), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [5]), .Z(n1650));
Q_MX02 U4316 ( .S(n1164), .A0(n1552), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [4]), .Z(n1649));
Q_MX02 U4317 ( .S(n1164), .A0(n1553), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [3]), .Z(n1648));
Q_MX02 U4318 ( .S(n1164), .A0(n1554), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [2]), .Z(n1647));
Q_MX02 U4319 ( .S(n1164), .A0(n1555), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [1]), .Z(n1646));
Q_MX02 U4320 ( .S(n1164), .A0(n1556), .A1(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [0]), .Z(n1645));
Q_INV U4321 ( .A(n1305), .Z(n1642));
Q_NR02 U4322 ( .A0(n1304), .A1(n1303), .Z(n1305));
Q_MX02 U4323 ( .S(n1630), .A0(n1299), .A1(n1291), .Z(n1304));
Q_MX02 U4324 ( .S(n1630), .A0(n1298), .A1(n1294), .Z(n1303));
Q_MX02 U4325 ( .S(n1630), .A0(n1297), .A1(n1293), .Z(n1302));
Q_MX02 U4326 ( .S(n1630), .A0(n1296), .A1(n1292), .Z(n1301));
Q_MX02 U4327 ( .S(n1630), .A0(n1295), .A1(n1284), .Z(n1300));
Q_MX02 U4328 ( .S(n1164), .A0(n1261), .A1(_zygsfis_ib_service_data_space[3]), .Z(n1298));
Q_MX02 U4329 ( .S(n1164), .A0(n1259), .A1(_zygsfis_ib_service_data_space[2]), .Z(n1297));
Q_MX02 U4330 ( .S(n1164), .A0(n1257), .A1(_zygsfis_ib_service_data_space[1]), .Z(n1296));
Q_XOR2 U4331 ( .A0(n1629), .A1(_zygsfis_ib_service_data_space[0]), .Z(n1295));
Q_INV U4332 ( .A(n1289), .Z(n1294));
Q_INV U4333 ( .A(n1288), .Z(n1293));
Q_INV U4334 ( .A(n1286), .Z(n1292));
Q_AD02 U4335 ( .CI(n1287), .A0(_zygsfis_ib_service_data_wptr[2]), .A1(_zygsfis_ib_service_data_wptr[3]), .B0(n1282), .B1(n1283), .S0(n1288), .S1(n1289), .CO(n1290));
Q_AD01 U4336 ( .CI(n1281), .A0(_zygsfis_ib_service_data_wptr[1]), .B0(n1285), .S(n1286), .CO(n1287));
Q_OR02 U4337 ( .A0(_zygsfis_ib_service_data_wptr[0]), .A1(n1280), .Z(n1285));
Q_XOR2 U4338 ( .A0(_zygsfis_ib_service_data_wptr[0]), .A1(n1280), .Z(n1284));
Q_XOR3 U4339 ( .A0(_zygsfis_ib_service_data_wptr[4]), .A1(n1273), .A2(n1290), .Z(n1291));
Q_INV U4340 ( .A(n1272), .Z(n1283));
Q_INV U4341 ( .A(n1271), .Z(n1282));
Q_INV U4342 ( .A(n1270), .Z(n1281));
Q_INV U4343 ( .A(n1269), .Z(n1280));
Q_AN02 U4344 ( .A0(n1279), .A1(_zygsfis_ib_service_data_eos), .Z(n1639));
Q_AN03 U4345 ( .A0(n1276), .A1(n1277), .A2(n1278), .Z(n1279));
Q_AN03 U4346 ( .A0(n1284), .A1(n1274), .A2(n1275), .Z(n1278));
Q_XNR2 U4347 ( .A0(n1273), .A1(_zygsfis_ib_service_data_wptr[4]), .Z(n1277));
Q_XNR2 U4348 ( .A0(n1272), .A1(_zygsfis_ib_service_data_wptr[3]), .Z(n1276));
Q_XNR2 U4349 ( .A0(n1271), .A1(_zygsfis_ib_service_data_wptr[2]), .Z(n1275));
Q_XNR2 U4350 ( .A0(n1270), .A1(_zygsfis_ib_service_data_wptr[1]), .Z(n1274));
Q_MX02 U4351 ( .S(n1164), .A0(n1267), .A1(_zygsfis_ib_service_data_rptr[3]), .Z(n1272));
Q_MX02 U4352 ( .S(n1164), .A0(n1265), .A1(_zygsfis_ib_service_data_rptr[2]), .Z(n1271));
Q_MX02 U4353 ( .S(n1164), .A0(n1263), .A1(_zygsfis_ib_service_data_rptr[1]), .Z(n1270));
Q_XOR2 U4354 ( .A0(n1629), .A1(_zygsfis_ib_service_data_rptr[0]), .Z(n1269));
Q_XOR2 U4355 ( .A0(_zygsfis_ib_service_data_rptr[4]), .A1(n5883), .Z(n1273));
Q_AD01HF U4356 ( .A0(_zygsfis_ib_service_data_rptr[3]), .B0(n1266), .S(n1267), .CO(n1268));
Q_AD01HF U4357 ( .A0(_zygsfis_ib_service_data_rptr[2]), .B0(n1264), .S(n1265), .CO(n1266));
Q_AD01HF U4358 ( .A0(_zygsfis_ib_service_data_rptr[1]), .B0(_zygsfis_ib_service_data_rptr[0]), .S(n1263), .CO(n1264));
Q_XOR2 U4359 ( .A0(_zygsfis_ib_service_data_space[4]), .A1(n5882), .Z(n1299));
Q_AD01HF U4360 ( .A0(_zygsfis_ib_service_data_space[3]), .B0(n1260), .S(n1261), .CO(n1262));
Q_AD01HF U4361 ( .A0(_zygsfis_ib_service_data_space[2]), .B0(n1258), .S(n1259), .CO(n1260));
Q_AD01HF U4362 ( .A0(_zygsfis_ib_service_data_space[1]), .B0(_zygsfis_ib_service_data_space[0]), .S(n1257), .CO(n1258));
Q_AD01HF U4363 ( .A0(_zygsfis_ib_service_data_req[3]), .B0(n1254), .S(n1255), .CO(n1256));
Q_AD01HF U4364 ( .A0(_zygsfis_ib_service_data_req[2]), .B0(n1252), .S(n1253), .CO(n1254));
Q_AD01HF U4365 ( .A0(_zygsfis_ib_service_data_req[1]), .B0(_zygsfis_ib_service_data_req[0]), .S(n1251), .CO(n1252));
Q_INV U4366 ( .A(n1250), .Z(n1644));
Q_OR02 U4367 ( .A0(n1248), .A1(n1249), .Z(n1250));
Q_OR03 U4368 ( .A0(n1245), .A1(n1246), .A2(n1247), .Z(n1249));
Q_OR03 U4369 ( .A0(n1242), .A1(n1243), .A2(n1244), .Z(n1248));
Q_OR03 U4370 ( .A0(n1239), .A1(n1240), .A2(n1241), .Z(n1247));
Q_OR03 U4371 ( .A0(n1236), .A1(n1237), .A2(n1238), .Z(n1246));
Q_OR03 U4372 ( .A0(n1231), .A1(n1233), .A2(n1235), .Z(n1245));
Q_OR03 U4373 ( .A0(n1225), .A1(n1227), .A2(n1229), .Z(n1244));
Q_OR03 U4374 ( .A0(n1219), .A1(n1221), .A2(n1223), .Z(n1243));
Q_OR03 U4375 ( .A0(n1213), .A1(n1215), .A2(n1217), .Z(n1242));
Q_OR03 U4376 ( .A0(n1207), .A1(n1209), .A2(n1211), .Z(n1241));
Q_OR03 U4377 ( .A0(n1201), .A1(n1203), .A2(n1205), .Z(n1240));
Q_OR03 U4378 ( .A0(n1195), .A1(n1197), .A2(n1199), .Z(n1239));
Q_OR03 U4379 ( .A0(n1189), .A1(n1191), .A2(n1193), .Z(n1238));
Q_OR03 U4380 ( .A0(n1183), .A1(n1185), .A2(n1187), .Z(n1237));
Q_OR03 U4381 ( .A0(n1177), .A1(n1179), .A2(n1181), .Z(n1236));
Q_OR03 U4382 ( .A0(n1747), .A1(n1234), .A2(n1175), .Z(n1235));
Q_INV U4383 ( .A(n1173), .Z(n1234));
Q_XOR2 U4384 ( .A0(mega_tlv_word_count[31]), .A1(n1232), .Z(n1233));
Q_AD01HF U4385 ( .A0(mega_tlv_word_count[30]), .B0(n1230), .S(n1231), .CO(n1232));
Q_AD01HF U4386 ( .A0(mega_tlv_word_count[29]), .B0(n1228), .S(n1229), .CO(n1230));
Q_AD01HF U4387 ( .A0(mega_tlv_word_count[28]), .B0(n1226), .S(n1227), .CO(n1228));
Q_AD01HF U4388 ( .A0(mega_tlv_word_count[27]), .B0(n1224), .S(n1225), .CO(n1226));
Q_AD01HF U4389 ( .A0(mega_tlv_word_count[26]), .B0(n1222), .S(n1223), .CO(n1224));
Q_AD01HF U4390 ( .A0(mega_tlv_word_count[25]), .B0(n1220), .S(n1221), .CO(n1222));
Q_AD01HF U4391 ( .A0(mega_tlv_word_count[24]), .B0(n1218), .S(n1219), .CO(n1220));
Q_AD01HF U4392 ( .A0(mega_tlv_word_count[23]), .B0(n1216), .S(n1217), .CO(n1218));
Q_AD01HF U4393 ( .A0(mega_tlv_word_count[22]), .B0(n1214), .S(n1215), .CO(n1216));
Q_AD01HF U4394 ( .A0(mega_tlv_word_count[21]), .B0(n1212), .S(n1213), .CO(n1214));
Q_AD01HF U4395 ( .A0(mega_tlv_word_count[20]), .B0(n1210), .S(n1211), .CO(n1212));
Q_AD01HF U4396 ( .A0(mega_tlv_word_count[19]), .B0(n1208), .S(n1209), .CO(n1210));
Q_AD01HF U4397 ( .A0(mega_tlv_word_count[18]), .B0(n1206), .S(n1207), .CO(n1208));
Q_AD01HF U4398 ( .A0(mega_tlv_word_count[17]), .B0(n1204), .S(n1205), .CO(n1206));
Q_AD01HF U4399 ( .A0(mega_tlv_word_count[16]), .B0(n1202), .S(n1203), .CO(n1204));
Q_AD01HF U4400 ( .A0(mega_tlv_word_count[15]), .B0(n1200), .S(n1201), .CO(n1202));
Q_AD01HF U4401 ( .A0(mega_tlv_word_count[14]), .B0(n1198), .S(n1199), .CO(n1200));
Q_AD01HF U4402 ( .A0(mega_tlv_word_count[13]), .B0(n1196), .S(n1197), .CO(n1198));
Q_AD01HF U4403 ( .A0(mega_tlv_word_count[12]), .B0(n1194), .S(n1195), .CO(n1196));
Q_AD01HF U4404 ( .A0(mega_tlv_word_count[11]), .B0(n1192), .S(n1193), .CO(n1194));
Q_AD01HF U4405 ( .A0(mega_tlv_word_count[10]), .B0(n1190), .S(n1191), .CO(n1192));
Q_AD01HF U4406 ( .A0(mega_tlv_word_count[9]), .B0(n1188), .S(n1189), .CO(n1190));
Q_AD01HF U4407 ( .A0(mega_tlv_word_count[8]), .B0(n1186), .S(n1187), .CO(n1188));
Q_AD01HF U4408 ( .A0(mega_tlv_word_count[7]), .B0(n1184), .S(n1185), .CO(n1186));
Q_AD01HF U4409 ( .A0(mega_tlv_word_count[6]), .B0(n1182), .S(n1183), .CO(n1184));
Q_AD01HF U4410 ( .A0(mega_tlv_word_count[5]), .B0(n1180), .S(n1181), .CO(n1182));
Q_AD01HF U4411 ( .A0(mega_tlv_word_count[4]), .B0(n1178), .S(n1179), .CO(n1180));
Q_AD01HF U4412 ( .A0(mega_tlv_word_count[3]), .B0(n1176), .S(n1177), .CO(n1178));
Q_AD01HF U4413 ( .A0(mega_tlv_word_count[2]), .B0(n1174), .S(n1175), .CO(n1176));
Q_AD01HF U4414 ( .A0(mega_tlv_word_count[1]), .B0(mega_tlv_word_count[0]), .S(n1173), .CO(n1174));
Q_XNR2 U4415 ( .A0(_zyGfifo__gfdL412_17_P0_m2_gfOff), .A1(_zyGfifoF19_L412_req_0), .Z(n1172));
Q_XNR2 U4416 ( .A0(_zyGfifo__gfdL530_18_P0_m2_gfOff), .A1(_zyGfifoF18_L530_req_0), .Z(n1171));
Q_XNR2 U4417 ( .A0(_zyGfifo__gfdL390_19_P0_m2_gfOff), .A1(_zyGfifoF17_L390_req_0), .Z(n1170));
Q_XNR2 U4418 ( .A0(_zyGfifo__gfdL381_20_P0_m2_gfOff), .A1(_zyGfifoF16_L381_req_0), .Z(n1169));
Q_XNR2 U4419 ( .A0(_zyGfifo__gfdL375_21_P0_m2_gfOff), .A1(_zyGfifoF15_L375_req_0), .Z(n1168));
Q_XNR2 U4420 ( .A0(_zyGfifo__gfdL373_22_P0_m2_gfOff), .A1(_zyGfifoF14_L373_req_0), .Z(n1167));
Q_XNR2 U4421 ( .A0(n1166), .A1(_zyGfifoF0_L368_s2_req_4), .Z(n1455));
Q_XNR2 U4422 ( .A0(_zyGfifo_ib_service_data_2_zyprefetch_m2_gfOff), .A1(_zyGfifoF11_L207_req_0), .Z(n1165));
Q_INV U4423 ( .A(n1164), .Z(n1629));
Q_AN03 U4424 ( .A0(n1159), .A1(n1158), .A2(n1163), .Z(n1164));
Q_AN03 U4425 ( .A0(n1162), .A1(n1161), .A2(n1160), .Z(n1163));
Q_XNR2 U4426 ( .A0(_zygsfis_ib_service_data_rptr[4]), .A1(_zygsfis_ib_service_data_wptr[4]), .Z(n1162));
Q_XNR2 U4427 ( .A0(_zygsfis_ib_service_data_rptr[3]), .A1(_zygsfis_ib_service_data_wptr[3]), .Z(n1161));
Q_XNR2 U4428 ( .A0(_zygsfis_ib_service_data_rptr[2]), .A1(_zygsfis_ib_service_data_wptr[2]), .Z(n1160));
Q_XNR2 U4429 ( .A0(_zygsfis_ib_service_data_rptr[1]), .A1(_zygsfis_ib_service_data_wptr[1]), .Z(n1159));
Q_XNR2 U4430 ( .A0(_zygsfis_ib_service_data_rptr[0]), .A1(_zygsfis_ib_service_data_wptr[0]), .Z(n1158));
Q_AN03 U4431 ( .A0(n1153), .A1(n1152), .A2(n1157), .Z(n1630));
Q_AN03 U4432 ( .A0(n1156), .A1(n1155), .A2(n1154), .Z(n1157));
Q_XNR2 U4433 ( .A0(_zygsfis_ib_service_data_req[4]), .A1(_zygsfis_ib_service_data_ack[4]), .Z(n1156));
Q_XNR2 U4434 ( .A0(_zygsfis_ib_service_data_req[3]), .A1(_zygsfis_ib_service_data_ack[3]), .Z(n1155));
Q_XNR2 U4435 ( .A0(_zygsfis_ib_service_data_req[2]), .A1(_zygsfis_ib_service_data_ack[2]), .Z(n1154));
Q_XNR2 U4436 ( .A0(_zygsfis_ib_service_data_req[1]), .A1(_zygsfis_ib_service_data_ack[1]), .Z(n1153));
Q_XNR2 U4437 ( .A0(_zygsfis_ib_service_data_req[0]), .A1(_zygsfis_ib_service_data_ack[0]), .Z(n1152));
Q_OR02 U4438 ( .A0(_zyM2L324_pbcFsm0_s[1]), .A1(_zyM2L324_pbcFsm0_s[2]), .Z(n1009));
Q_OR02 U4439 ( .A0(n1129), .A1(_zyM2L324_pbcFsm0_s[2]), .Z(n1037));
Q_AN02 U4440 ( .A0(n1008), .A1(n1049), .Z(n1050));
Q_OR03 U4441 ( .A0(_zyM2L324_pbcFsm0_s[1]), .A1(n1023), .A2(_zyM2L324_pbcFsm0_s[0]), .Z(n1027));
Q_OR03 U4442 ( .A0(_zyM2L324_pbcFsm0_s[2]), .A1(n548), .A2(_zyM2L324_pbcFsm0_s[1]), .Z(n1034));
Q_INV U4443 ( .A(n1031), .Z(n1126));
Q_OA21 U4444 ( .A0(_zyM2L324_pbcFsm0_s[2]), .A1(n1130), .B0(n1049), .Z(n1048));
Q_OR02 U4445 ( .A0(n1037), .A1(_zyM2L324_pbcFsm0_s[0]), .Z(n1049));
Q_ND02 U4446 ( .A0(n1148), .A1(n1145), .Z(n1047));
Q_OR03 U4447 ( .A0(n1046), .A1(n1147), .A2(n1047), .Z(n1044));
Q_INV U4448 ( .A(n1150), .Z(n1046));
Q_OR03 U4449 ( .A0(n1045), .A1(n1151), .A2(n1024), .Z(n1043));
Q_INV U4450 ( .A(n1142), .Z(n1045));
Q_OR02 U4451 ( .A0(n1043), .A1(n1044), .Z(n1039));
Q_INV U4452 ( .A(n1146), .Z(n1042));
Q_OR02 U4453 ( .A0(n1042), .A1(n1039), .Z(n1005));
Q_INV U4454 ( .A(n1144), .Z(n1004));
Q_OR02 U4455 ( .A0(n1004), .A1(n1005), .Z(n1001));
Q_OR02 U4456 ( .A0(_zyM2L324_pbcFsm0_s[2]), .A1(n1001), .Z(n1014));
Q_MX02 U4457 ( .S(_zyM2L324_pbcFsm0_s[1]), .A0(n1014), .A1(_zyM2L324_pbcFsm0_s[2]), .Z(n1041));
Q_OR02 U4458 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(n1041), .Z(n1040));
Q_OR02 U4459 ( .A0(n1146), .A1(n1039), .Z(n1003));
Q_OR02 U4460 ( .A0(n1144), .A1(n1003), .Z(n999));
Q_OR03 U4461 ( .A0(n1009), .A1(n999), .A2(_zyM2L324_pbcFsm0_s[0]), .Z(n1012));
Q_AN02 U4462 ( .A0(n1008), .A1(n1012), .Z(n1038));
Q_OA21 U4463 ( .A0(n1037), .A1(n1130), .B0(n1036), .Z(n1035));
Q_OR02 U4464 ( .A0(n1009), .A1(_zyM2L324_pbcFsm0_s[0]), .Z(n1036));
Q_OR02 U4465 ( .A0(n1034), .A1(n1130), .Z(n1031));
Q_ND02 U4466 ( .A0(config_ready), .A1(n1142), .Z(n1033));
Q_OR03 U4467 ( .A0(n1009), .A1(n1033), .A2(_zyM2L324_pbcFsm0_s[0]), .Z(n1032));
Q_AN02 U4468 ( .A0(n1031), .A1(n1032), .Z(n1030));
Q_INV U4469 ( .A(n1030), .Z(n1139));
Q_INV U4470 ( .A(_zyL94_iscX1c0_o2), .Z(n1029));
Q_OR03 U4471 ( .A0(_zyM2L324_pbcFsm0_s[2]), .A1(n1029), .A2(_zyM2L324_pbcFsm0_s[1]), .Z(n1028));
Q_OA21 U4472 ( .A0(n1028), .A1(n1130), .B0(n1027), .Z(n1026));
Q_INV U4473 ( .A(_zyL61_iscX2c0_o2), .Z(n1025));
Q_OR02 U4474 ( .A0(_zyM2L324_pbcFsm0_s[2]), .A1(n1025), .Z(n1017));
Q_OR03 U4475 ( .A0(n1133), .A1(n628), .A2(n1023), .Z(n1011));
Q_OR02 U4476 ( .A0(_zyM2L324_pbcFsm0_s[2]), .A1(n1024), .Z(n1023));
Q_MX02 U4477 ( .S(_zyM2L324_pbcFsm0_s[1]), .A0(n1011), .A1(n1017), .Z(n1022));
Q_OA21 U4478 ( .A0(n1022), .A1(_zyM2L324_pbcFsm0_s[0]), .B0(n1008), .Z(n1021));
Q_INV U4479 ( .A(n1021), .Z(n1138));
Q_NR02 U4480 ( .A0(_zyL94_iscX1c0_o2), .A1(n1020), .Z(n1019));
Q_OR02 U4481 ( .A0(n1009), .A1(n1019), .Z(n1018));
Q_OR02 U4482 ( .A0(n1129), .A1(n1017), .Z(n1016));
Q_MX02 U4483 ( .S(_zyM2L324_pbcFsm0_s[0]), .A0(n1016), .A1(n1018), .Z(n1015));
Q_INV U4484 ( .A(n1015), .Z(n1137));
Q_OR02 U4485 ( .A0(n1006), .A1(n1014), .Z(n1013));
Q_INV U4486 ( .A(n1013), .Z(n1136));
Q_INV U4487 ( .A(n1012), .Z(n1135));
Q_OR02 U4488 ( .A0(n1006), .A1(n1011), .Z(n1010));
Q_INV U4489 ( .A(n1010), .Z(n1134));
Q_OR02 U4490 ( .A0(n1130), .A1(n1009), .Z(n1008));
Q_OR02 U4491 ( .A0(n1133), .A1(n1141), .Z(n1007));
Q_OR02 U4492 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(_zyM2L324_pbcFsm0_s[1]), .Z(n1006));
Q_INV U4493 ( .A(n1006), .Z(n1132));
Q_MX02 U4494 ( .S(n1144), .A0(n1003), .A1(n1005), .Z(n1125));
Q_OR02 U4495 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(n1125), .Z(n1131));
Q_XNR2 U4496 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(n1129), .Z(n1002));
Q_AO21 U4497 ( .A0(n1129), .A1(n1001), .B0(_zyM2L324_pbcFsm0_s[0]), .Z(n1000));
Q_ND02 U4498 ( .A0(n997), .A1(n1000), .Z(n1128));
Q_OR02 U4499 ( .A0(_zyM2L324_pbcFsm0_s[1]), .A1(n1130), .Z(n997));
Q_AO21 U4500 ( .A0(n1129), .A1(n999), .B0(_zyM2L324_pbcFsm0_s[0]), .Z(n998));
Q_ND02 U4501 ( .A0(n997), .A1(n998), .Z(n1127));
Q_AN02 U4502 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[31]), .Z(n996));
Q_AN02 U4503 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[30]), .Z(n995));
Q_AN02 U4504 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[29]), .Z(n994));
Q_AN02 U4505 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[28]), .Z(n993));
Q_AN02 U4506 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[27]), .Z(n992));
Q_AN02 U4507 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[26]), .Z(n991));
Q_AN02 U4508 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[25]), .Z(n990));
Q_AN02 U4509 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[24]), .Z(n989));
Q_AN02 U4510 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[23]), .Z(n988));
Q_AN02 U4511 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[22]), .Z(n987));
Q_AN02 U4512 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[21]), .Z(n986));
Q_AN02 U4513 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[20]), .Z(n985));
Q_AN02 U4514 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[19]), .Z(n984));
Q_AN02 U4515 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[18]), .Z(n983));
Q_AN02 U4516 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[17]), .Z(n982));
Q_AN02 U4517 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[16]), .Z(n981));
Q_AN02 U4518 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[15]), .Z(n980));
Q_AN02 U4519 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[14]), .Z(n979));
Q_AN02 U4520 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[13]), .Z(n978));
Q_AN02 U4521 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[12]), .Z(n977));
Q_AN02 U4522 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[11]), .Z(n976));
Q_AN02 U4523 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[10]), .Z(n975));
Q_AN02 U4524 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[9]), .Z(n974));
Q_AN02 U4525 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[8]), .Z(n973));
Q_AN02 U4526 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[7]), .Z(n972));
Q_AN02 U4527 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[6]), .Z(n971));
Q_AN02 U4528 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[5]), .Z(n970));
Q_AN02 U4529 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[4]), .Z(n969));
Q_AN02 U4530 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[3]), .Z(n968));
Q_AN02 U4531 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[2]), .Z(n967));
Q_MX02 U4532 ( .S(_zyM2L324_pbcFsm0_s[0]), .A0(n1133), .A1(address[1]), .Z(n966));
Q_MX02 U4533 ( .S(_zyM2L324_pbcFsm0_s[0]), .A0(n1123), .A1(address[0]), .Z(n965));
Q_NR02 U4534 ( .A0(n500), .A1(n1133), .Z(n1142));
Q_FDP0 _zzM2L324_mdxP2_error_cntr_Dwen0_REG  ( .CK(_zyM2L324_pbcMevClk4), .D(n1126), .Q(_zzM2L324_mdxP2_error_cntr_Dwen0), .QN( ));
Q_FDP0 \_zyM2L324_pbcFsm0_s_REG[2] ( .CK(_zyM2L324_pbcMevClk4), .D(_zyM2L324_pbcFsm0_s[2]), .Q(_zyM2L324_pbcFsm0_s[2]), .QN(n1140));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[0] ( .CK(_zyM2L324_pbcMevClk4), .D(n923), .Q(_zzM2L324_mdxP2_error_cntr_wr0[0]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[1] ( .CK(_zyM2L324_pbcMevClk4), .D(n924), .Q(_zzM2L324_mdxP2_error_cntr_wr0[1]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[2] ( .CK(_zyM2L324_pbcMevClk4), .D(n925), .Q(_zzM2L324_mdxP2_error_cntr_wr0[2]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[3] ( .CK(_zyM2L324_pbcMevClk4), .D(n926), .Q(_zzM2L324_mdxP2_error_cntr_wr0[3]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[4] ( .CK(_zyM2L324_pbcMevClk4), .D(n927), .Q(_zzM2L324_mdxP2_error_cntr_wr0[4]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[5] ( .CK(_zyM2L324_pbcMevClk4), .D(n928), .Q(_zzM2L324_mdxP2_error_cntr_wr0[5]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[6] ( .CK(_zyM2L324_pbcMevClk4), .D(n929), .Q(_zzM2L324_mdxP2_error_cntr_wr0[6]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[7] ( .CK(_zyM2L324_pbcMevClk4), .D(n930), .Q(_zzM2L324_mdxP2_error_cntr_wr0[7]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[8] ( .CK(_zyM2L324_pbcMevClk4), .D(n931), .Q(_zzM2L324_mdxP2_error_cntr_wr0[8]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[9] ( .CK(_zyM2L324_pbcMevClk4), .D(n932), .Q(_zzM2L324_mdxP2_error_cntr_wr0[9]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[10] ( .CK(_zyM2L324_pbcMevClk4), .D(n933), .Q(_zzM2L324_mdxP2_error_cntr_wr0[10]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[11] ( .CK(_zyM2L324_pbcMevClk4), .D(n934), .Q(_zzM2L324_mdxP2_error_cntr_wr0[11]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[12] ( .CK(_zyM2L324_pbcMevClk4), .D(n935), .Q(_zzM2L324_mdxP2_error_cntr_wr0[12]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[13] ( .CK(_zyM2L324_pbcMevClk4), .D(n936), .Q(_zzM2L324_mdxP2_error_cntr_wr0[13]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[14] ( .CK(_zyM2L324_pbcMevClk4), .D(n937), .Q(_zzM2L324_mdxP2_error_cntr_wr0[14]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[15] ( .CK(_zyM2L324_pbcMevClk4), .D(n938), .Q(_zzM2L324_mdxP2_error_cntr_wr0[15]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[16] ( .CK(_zyM2L324_pbcMevClk4), .D(n939), .Q(_zzM2L324_mdxP2_error_cntr_wr0[16]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[17] ( .CK(_zyM2L324_pbcMevClk4), .D(n940), .Q(_zzM2L324_mdxP2_error_cntr_wr0[17]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[18] ( .CK(_zyM2L324_pbcMevClk4), .D(n941), .Q(_zzM2L324_mdxP2_error_cntr_wr0[18]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[19] ( .CK(_zyM2L324_pbcMevClk4), .D(n942), .Q(_zzM2L324_mdxP2_error_cntr_wr0[19]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[20] ( .CK(_zyM2L324_pbcMevClk4), .D(n943), .Q(_zzM2L324_mdxP2_error_cntr_wr0[20]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[21] ( .CK(_zyM2L324_pbcMevClk4), .D(n944), .Q(_zzM2L324_mdxP2_error_cntr_wr0[21]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[22] ( .CK(_zyM2L324_pbcMevClk4), .D(n945), .Q(_zzM2L324_mdxP2_error_cntr_wr0[22]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[23] ( .CK(_zyM2L324_pbcMevClk4), .D(n946), .Q(_zzM2L324_mdxP2_error_cntr_wr0[23]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[24] ( .CK(_zyM2L324_pbcMevClk4), .D(n947), .Q(_zzM2L324_mdxP2_error_cntr_wr0[24]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[25] ( .CK(_zyM2L324_pbcMevClk4), .D(n948), .Q(_zzM2L324_mdxP2_error_cntr_wr0[25]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[26] ( .CK(_zyM2L324_pbcMevClk4), .D(n949), .Q(_zzM2L324_mdxP2_error_cntr_wr0[26]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[27] ( .CK(_zyM2L324_pbcMevClk4), .D(n950), .Q(_zzM2L324_mdxP2_error_cntr_wr0[27]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[28] ( .CK(_zyM2L324_pbcMevClk4), .D(n951), .Q(_zzM2L324_mdxP2_error_cntr_wr0[28]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[29] ( .CK(_zyM2L324_pbcMevClk4), .D(n952), .Q(_zzM2L324_mdxP2_error_cntr_wr0[29]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[30] ( .CK(_zyM2L324_pbcMevClk4), .D(n953), .Q(_zzM2L324_mdxP2_error_cntr_wr0[30]), .QN( ));
Q_FDP0 \_zzM2L324_mdxP2_error_cntr_wr0_REG[31] ( .CK(_zyM2L324_pbcMevClk4), .D(n954), .Q(_zzM2L324_mdxP2_error_cntr_wr0[31]), .QN( ));
Q_MX02 U4569 ( .S(n1007), .A0(n627), .A1(n963), .Z(n964));
Q_AN02 U4570 ( .A0(n1133), .A1(n622), .Z(n963));
Q_MX02 U4571 ( .S(n1007), .A0(n626), .A1(n961), .Z(n962));
Q_AN02 U4572 ( .A0(n1133), .A1(n621), .Z(n961));
Q_MX02 U4573 ( .S(n1007), .A0(n625), .A1(n959), .Z(n960));
Q_AN02 U4574 ( .A0(n1133), .A1(n620), .Z(n959));
Q_MX02 U4575 ( .S(n1007), .A0(n624), .A1(n957), .Z(n958));
Q_AN02 U4576 ( .A0(n1133), .A1(n619), .Z(n957));
Q_MX02 U4577 ( .S(n1007), .A0(n623), .A1(n955), .Z(n956));
Q_AN02 U4578 ( .A0(n1133), .A1(n618), .Z(n955));
Q_MX02 U4579 ( .S(n1031), .A0(n2261), .A1(error_cntr[31]), .Z(n954));
Q_MX02 U4580 ( .S(n1031), .A0(n2259), .A1(error_cntr[30]), .Z(n953));
Q_MX02 U4581 ( .S(n1031), .A0(n2257), .A1(error_cntr[29]), .Z(n952));
Q_MX02 U4582 ( .S(n1031), .A0(n2255), .A1(error_cntr[28]), .Z(n951));
Q_MX02 U4583 ( .S(n1031), .A0(n2253), .A1(error_cntr[27]), .Z(n950));
Q_MX02 U4584 ( .S(n1031), .A0(n2251), .A1(error_cntr[26]), .Z(n949));
Q_MX02 U4585 ( .S(n1031), .A0(n2249), .A1(error_cntr[25]), .Z(n948));
Q_MX02 U4586 ( .S(n1031), .A0(n2247), .A1(error_cntr[24]), .Z(n947));
Q_MX02 U4587 ( .S(n1031), .A0(n2245), .A1(error_cntr[23]), .Z(n946));
Q_MX02 U4588 ( .S(n1031), .A0(n2243), .A1(error_cntr[22]), .Z(n945));
Q_MX02 U4589 ( .S(n1031), .A0(n2241), .A1(error_cntr[21]), .Z(n944));
Q_MX02 U4590 ( .S(n1031), .A0(n2239), .A1(error_cntr[20]), .Z(n943));
Q_MX02 U4591 ( .S(n1031), .A0(n2237), .A1(error_cntr[19]), .Z(n942));
Q_MX02 U4592 ( .S(n1031), .A0(n2235), .A1(error_cntr[18]), .Z(n941));
Q_MX02 U4593 ( .S(n1031), .A0(n2233), .A1(error_cntr[17]), .Z(n940));
Q_MX02 U4594 ( .S(n1031), .A0(n2231), .A1(error_cntr[16]), .Z(n939));
Q_MX02 U4595 ( .S(n1031), .A0(n2229), .A1(error_cntr[15]), .Z(n938));
Q_MX02 U4596 ( .S(n1031), .A0(n2227), .A1(error_cntr[14]), .Z(n937));
Q_MX02 U4597 ( .S(n1031), .A0(n2225), .A1(error_cntr[13]), .Z(n936));
Q_MX02 U4598 ( .S(n1031), .A0(n2223), .A1(error_cntr[12]), .Z(n935));
Q_MX02 U4599 ( .S(n1031), .A0(n2221), .A1(error_cntr[11]), .Z(n934));
Q_MX02 U4600 ( .S(n1031), .A0(n2219), .A1(error_cntr[10]), .Z(n933));
Q_MX02 U4601 ( .S(n1031), .A0(n2217), .A1(error_cntr[9]), .Z(n932));
Q_MX02 U4602 ( .S(n1031), .A0(n2215), .A1(error_cntr[8]), .Z(n931));
Q_MX02 U4603 ( .S(n1031), .A0(n2213), .A1(error_cntr[7]), .Z(n930));
Q_MX02 U4604 ( .S(n1031), .A0(n2211), .A1(error_cntr[6]), .Z(n929));
Q_MX02 U4605 ( .S(n1031), .A0(n2209), .A1(error_cntr[5]), .Z(n928));
Q_MX02 U4606 ( .S(n1031), .A0(n2207), .A1(error_cntr[4]), .Z(n927));
Q_MX02 U4607 ( .S(n1031), .A0(n2205), .A1(error_cntr[3]), .Z(n926));
Q_MX02 U4608 ( .S(n1031), .A0(n2203), .A1(error_cntr[2]), .Z(n925));
Q_MX02 U4609 ( .S(n1031), .A0(n2201), .A1(error_cntr[1]), .Z(n924));
Q_XOR2 U4610 ( .A0(n1126), .A1(error_cntr[0]), .Z(n923));
Q_MX02 U4611 ( .S(n1006), .A0(n549), .A1(n921), .Z(n922));
Q_MX02 U4612 ( .S(_zyM2L324_pbcFsm0_s[0]), .A0(_zyGfifo__gfdL351_25_P0_m2_gfOff), .A1(_zyGfifo__gfdL334_28_P0_m2_gfOff), .Z(n552));
Q_AN02 U4613 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[1]), .Z(n920));
Q_AN02 U4614 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(address[0]), .Z(n919));
Q_AN02 U4615 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[31]), .Z(n918));
Q_AN02 U4616 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[30]), .Z(n917));
Q_AN02 U4617 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[29]), .Z(n916));
Q_AN02 U4618 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[28]), .Z(n915));
Q_AN02 U4619 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[27]), .Z(n914));
Q_AN02 U4620 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[26]), .Z(n913));
Q_AN02 U4621 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[25]), .Z(n912));
Q_AN02 U4622 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[24]), .Z(n911));
Q_AN02 U4623 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[23]), .Z(n910));
Q_AN02 U4624 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[22]), .Z(n909));
Q_AN02 U4625 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[21]), .Z(n908));
Q_AN02 U4626 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[20]), .Z(n907));
Q_AN02 U4627 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[19]), .Z(n906));
Q_AN02 U4628 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[18]), .Z(n905));
Q_AN02 U4629 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[17]), .Z(n904));
Q_AN02 U4630 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[16]), .Z(n903));
Q_AN02 U4631 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[15]), .Z(n902));
Q_AN02 U4632 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[14]), .Z(n901));
Q_AN02 U4633 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[13]), .Z(n900));
Q_AN02 U4634 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[12]), .Z(n899));
Q_AN02 U4635 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[11]), .Z(n898));
Q_AN02 U4636 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[10]), .Z(n897));
Q_AN02 U4637 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[9]), .Z(n896));
Q_AN02 U4638 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[8]), .Z(n895));
Q_AN02 U4639 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[7]), .Z(n894));
Q_AN02 U4640 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[6]), .Z(n893));
Q_AN02 U4641 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[5]), .Z(n892));
Q_AN02 U4642 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[4]), .Z(n891));
Q_AN02 U4643 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[3]), .Z(n890));
Q_AN02 U4644 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[2]), .Z(n889));
Q_AN02 U4645 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[1]), .Z(n888));
Q_AN02 U4646 ( .A0(_zyM2L324_pbcFsm0_s[0]), .A1(data[0]), .Z(n887));
Q_MX02 U4647 ( .S(_zyM2L324_pbcFsm0_s[1]), .A0(n885), .A1(address[31]), .Z(n886));
Q_AN02 U4648 ( .A0(n1006), .A1(_zyL94_iscX1c0_o1[31]), .Z(n885));
Q_MX02 U4649 ( .S(_zyM2L324_pbcFsm0_s[1]), .A0(n883), .A1(address[30]), .Z(n884));
Q_AN02 U4650 ( .A0(n1006), .A1(_zyL94_iscX1c0_o1[30]), .Z(n883));
Q_MX02 U4651 ( .S(_zyM2L324_pbcFsm0_s[1]), .A0(n881), .A1(address[29]), .Z(n882));
Q_AN02 U4652 ( .A0(n1006), .A1(_zyL94_iscX1c0_o1[29]), .Z(n881));
Q_MX02 U4653 ( .S(_zyM2L324_pbcFsm0_s[1]), .A0(n879), .A1(address[28]), .Z(n880));
Q_AN02 U4654 ( .A0(n1006), .A1(_zyL94_iscX1c0_o1[28]), .Z(n879));
Q_MX02 U4655 ( .S(_zyM2L324_pbcFsm0_s[1]), .A0(n877), .A1(address[27]), .Z(n878));
Q_AN02 U4656 ( .A0(n1006), .A1(_zyL94_iscX1c0_o1[27]), .Z(n877));
Q_MX02 U4657 ( .S(_zyM2L324_pbcFsm0_s[1]), .A0(n875), .A1(address[26]), .Z(n876));
Q_AN02 U4658 ( .A0(n1006), .A1(_zyL94_iscX1c0_o1[26]), .Z(n875));
Q_MX02 U4659 ( .S(_zyM2L324_pbcFsm0_s[1]), .A0(n873), .A1(address[25]), .Z(n874));
Q_AN02 U4660 ( .A0(n1006), .A1(_zyL94_iscX1c0_o1[25]), .Z(n873));
Q_MX02 U4661 ( .S(_zyM2L324_pbcFsm0_s[1]), .A0(n871), .A1(address[24]), .Z(n872));
Q_AN02 U4662 ( .A0(n1006), .A1(_zyL94_iscX1c0_o1[24]), .Z(n871));
Q_MX02 U4663 ( .S(_zyM2L324_pbcFsm0_s[1]), .A0(n869), .A1(address[23]), .Z(n870));
Q_AN02 U4664 ( .A0(n1006), .A1(_zyL94_iscX1c0_o1[23]), .Z(n869));
Q_MX02 U4665 ( .S(_zyM2L324_pbcFsm0_s[1]), .A0(n867), .A1(address[22]), .Z(n868));
Q_AN02 U4666 ( .A0(n1006), .A1(_zyL94_iscX1c0_o1[22]), .Z(n867));
Q_MX02 U4667 ( .S(_zyM2L324_pbcFsm0_s[1]), .A0(n865), .A1(address[21]), .Z(n866));
Q_AN02 U4668 ( .A0(n1006), .A1(_zyL94_iscX1c0_o1[21]), .Z(n865));
Q_MX02 U4669 ( .S(_zyM2L324_pbcFsm0_s[1]), .A0(n863), .A1(address[20]), .Z(n864));
Q_AN02 U4670 ( .A0(n1006), .A1(_zyL94_iscX1c0_o1[20]), .Z(n863));
Q_MX02 U4671 ( .S(_zyM2L324_pbcFsm0_s[1]), .A0(n861), .A1(address[19]), .Z(n862));
Q_AN02 U4672 ( .A0(n1006), .A1(_zyL94_iscX1c0_o1[19]), .Z(n861));
Q_MX02 U4673 ( .S(_zyM2L324_pbcFsm0_s[1]), .A0(n859), .A1(address[18]), .Z(n860));
Q_AN02 U4674 ( .A0(n1006), .A1(_zyL94_iscX1c0_o1[18]), .Z(n859));
Q_MX02 U4675 ( .S(_zyM2L324_pbcFsm0_s[1]), .A0(n857), .A1(address[17]), .Z(n858));
Q_AN02 U4676 ( .A0(n1006), .A1(_zyL94_iscX1c0_o1[17]), .Z(n857));
Q_MX02 U4677 ( .S(_zyM2L324_pbcFsm0_s[1]), .A0(n855), .A1(address[16]), .Z(n856));
Q_AN02 U4678 ( .A0(n1006), .A1(_zyL94_iscX1c0_o1[16]), .Z(n855));
Q_MX02 U4679 ( .S(_zyM2L324_pbcFsm0_s[1]), .A0(n853), .A1(address[15]), .Z(n854));
Q_AN02 U4680 ( .A0(n1006), .A1(_zyL94_iscX1c0_o1[15]), .Z(n853));
Q_MX02 U4681 ( .S(_zyM2L324_pbcFsm0_s[1]), .A0(n851), .A1(address[14]), .Z(n852));
Q_AN02 U4682 ( .A0(n1006), .A1(_zyL94_iscX1c0_o1[14]), .Z(n851));
Q_MX02 U4683 ( .S(_zyM2L324_pbcFsm0_s[1]), .A0(n849), .A1(address[13]), .Z(n850));
Q_AN02 U4684 ( .A0(n1006), .A1(_zyL94_iscX1c0_o1[13]), .Z(n849));
Q_MX02 U4685 ( .S(_zyM2L324_pbcFsm0_s[1]), .A0(n847), .A1(address[12]), .Z(n848));
Q_AN02 U4686 ( .A0(n1006), .A1(_zyL94_iscX1c0_o1[12]), .Z(n847));
Q_MX02 U4687 ( .S(_zyM2L324_pbcFsm0_s[1]), .A0(n845), .A1(address[11]), .Z(n846));
Q_AN02 U4688 ( .A0(n1006), .A1(_zyL94_iscX1c0_o1[11]), .Z(n845));
Q_MX02 U4689 ( .S(_zyM2L324_pbcFsm0_s[1]), .A0(n843), .A1(address[10]), .Z(n844));
Q_AN02 U4690 ( .A0(n1006), .A1(_zyL94_iscX1c0_o1[10]), .Z(n843));
Q_MX02 U4691 ( .S(_zyM2L324_pbcFsm0_s[1]), .A0(n841), .A1(address[9]), .Z(n842));
Q_AN02 U4692 ( .A0(n1006), .A1(_zyL94_iscX1c0_o1[9]), .Z(n841));
Q_MX02 U4693 ( .S(_zyM2L324_pbcFsm0_s[1]), .A0(n839), .A1(address[8]), .Z(n840));
Q_AN02 U4694 ( .A0(n1006), .A1(_zyL94_iscX1c0_o1[8]), .Z(n839));
Q_MX02 U4695 ( .S(_zyM2L324_pbcFsm0_s[1]), .A0(n837), .A1(address[7]), .Z(n838));
Q_AN02 U4696 ( .A0(n1006), .A1(_zyL94_iscX1c0_o1[7]), .Z(n837));
Q_MX02 U4697 ( .S(_zyM2L324_pbcFsm0_s[1]), .A0(n835), .A1(address[6]), .Z(n836));
Q_AN02 U4698 ( .A0(n1006), .A1(_zyL94_iscX1c0_o1[6]), .Z(n835));
Q_MX02 U4699 ( .S(_zyM2L324_pbcFsm0_s[1]), .A0(n833), .A1(address[5]), .Z(n834));
Q_AN02 U4700 ( .A0(n1006), .A1(_zyL94_iscX1c0_o1[5]), .Z(n833));
Q_MX03 U4701 ( .S0(n1132), .S1(_zyM2L324_pbcFsm0_s[1]), .A0(_zyL94_iscX1c0_o1[4]), .A1(n627), .A2(address[4]), .Z(n832));
Q_MX03 U4702 ( .S0(n1132), .S1(_zyM2L324_pbcFsm0_s[1]), .A0(_zyL94_iscX1c0_o1[3]), .A1(n626), .A2(address[3]), .Z(n831));
Q_MX03 U4703 ( .S0(n1132), .S1(_zyM2L324_pbcFsm0_s[1]), .A0(_zyL94_iscX1c0_o1[2]), .A1(n625), .A2(address[2]), .Z(n830));
Q_MX03 U4704 ( .S0(n1132), .S1(_zyM2L324_pbcFsm0_s[1]), .A0(_zyL94_iscX1c0_o1[1]), .A1(n624), .A2(address[1]), .Z(n829));
Q_MX03 U4705 ( .S0(n1132), .S1(_zyM2L324_pbcFsm0_s[1]), .A0(_zyL94_iscX1c0_o1[0]), .A1(n623), .A2(address[0]), .Z(n828));
Q_MX03 U4706 ( .S0(_zyM2L324_pbcFsm0_s[0]), .S1(n1132), .A0(_zyGfifo__gfdL351_25_P0_m2_cbid[19]), .A1(_zyGfifo__gfdL334_28_P0_m2_cbid[19]), .A2(_zyGfifo_get_config_data_2_zyprefetch_m2_cbid[19]), .Z(n827));
Q_MX03 U4707 ( .S0(_zyM2L324_pbcFsm0_s[0]), .S1(n1132), .A0(_zyGfifo__gfdL351_25_P0_m2_cbid[18]), .A1(_zyGfifo__gfdL334_28_P0_m2_cbid[18]), .A2(_zyGfifo_get_config_data_2_zyprefetch_m2_cbid[18]), .Z(n826));
Q_MX03 U4708 ( .S0(_zyM2L324_pbcFsm0_s[0]), .S1(n1132), .A0(_zyGfifo__gfdL351_25_P0_m2_cbid[17]), .A1(_zyGfifo__gfdL334_28_P0_m2_cbid[17]), .A2(_zyGfifo_get_config_data_2_zyprefetch_m2_cbid[17]), .Z(n825));
Q_MX03 U4709 ( .S0(_zyM2L324_pbcFsm0_s[0]), .S1(n1132), .A0(_zyGfifo__gfdL351_25_P0_m2_cbid[16]), .A1(_zyGfifo__gfdL334_28_P0_m2_cbid[16]), .A2(_zyGfifo_get_config_data_2_zyprefetch_m2_cbid[16]), .Z(n824));
Q_MX03 U4710 ( .S0(_zyM2L324_pbcFsm0_s[0]), .S1(n1132), .A0(_zyGfifo__gfdL351_25_P0_m2_cbid[15]), .A1(_zyGfifo__gfdL334_28_P0_m2_cbid[15]), .A2(_zyGfifo_get_config_data_2_zyprefetch_m2_cbid[15]), .Z(n823));
Q_MX03 U4711 ( .S0(_zyM2L324_pbcFsm0_s[0]), .S1(n1132), .A0(_zyGfifo__gfdL351_25_P0_m2_cbid[14]), .A1(_zyGfifo__gfdL334_28_P0_m2_cbid[14]), .A2(_zyGfifo_get_config_data_2_zyprefetch_m2_cbid[14]), .Z(n822));
Q_MX03 U4712 ( .S0(_zyM2L324_pbcFsm0_s[0]), .S1(n1132), .A0(_zyGfifo__gfdL351_25_P0_m2_cbid[13]), .A1(_zyGfifo__gfdL334_28_P0_m2_cbid[13]), .A2(_zyGfifo_get_config_data_2_zyprefetch_m2_cbid[13]), .Z(n821));
Q_MX03 U4713 ( .S0(_zyM2L324_pbcFsm0_s[0]), .S1(n1132), .A0(_zyGfifo__gfdL351_25_P0_m2_cbid[12]), .A1(_zyGfifo__gfdL334_28_P0_m2_cbid[12]), .A2(_zyGfifo_get_config_data_2_zyprefetch_m2_cbid[12]), .Z(n820));
Q_MX03 U4714 ( .S0(_zyM2L324_pbcFsm0_s[0]), .S1(n1132), .A0(_zyGfifo__gfdL351_25_P0_m2_cbid[11]), .A1(_zyGfifo__gfdL334_28_P0_m2_cbid[11]), .A2(_zyGfifo_get_config_data_2_zyprefetch_m2_cbid[11]), .Z(n819));
Q_MX03 U4715 ( .S0(_zyM2L324_pbcFsm0_s[0]), .S1(n1132), .A0(_zyGfifo__gfdL351_25_P0_m2_cbid[10]), .A1(_zyGfifo__gfdL334_28_P0_m2_cbid[10]), .A2(_zyGfifo_get_config_data_2_zyprefetch_m2_cbid[10]), .Z(n818));
Q_MX03 U4716 ( .S0(_zyM2L324_pbcFsm0_s[0]), .S1(n1132), .A0(_zyGfifo__gfdL351_25_P0_m2_cbid[9]), .A1(_zyGfifo__gfdL334_28_P0_m2_cbid[9]), .A2(_zyGfifo_get_config_data_2_zyprefetch_m2_cbid[9]), .Z(n817));
Q_MX03 U4717 ( .S0(_zyM2L324_pbcFsm0_s[0]), .S1(n1132), .A0(_zyGfifo__gfdL351_25_P0_m2_cbid[8]), .A1(_zyGfifo__gfdL334_28_P0_m2_cbid[8]), .A2(_zyGfifo_get_config_data_2_zyprefetch_m2_cbid[8]), .Z(n816));
Q_MX03 U4718 ( .S0(_zyM2L324_pbcFsm0_s[0]), .S1(n1132), .A0(_zyGfifo__gfdL351_25_P0_m2_cbid[7]), .A1(_zyGfifo__gfdL334_28_P0_m2_cbid[7]), .A2(_zyGfifo_get_config_data_2_zyprefetch_m2_cbid[7]), .Z(n815));
Q_MX03 U4719 ( .S0(_zyM2L324_pbcFsm0_s[0]), .S1(n1132), .A0(_zyGfifo__gfdL351_25_P0_m2_cbid[6]), .A1(_zyGfifo__gfdL334_28_P0_m2_cbid[6]), .A2(_zyGfifo_get_config_data_2_zyprefetch_m2_cbid[6]), .Z(n814));
Q_MX03 U4720 ( .S0(_zyM2L324_pbcFsm0_s[0]), .S1(n1132), .A0(_zyGfifo__gfdL351_25_P0_m2_cbid[5]), .A1(_zyGfifo__gfdL334_28_P0_m2_cbid[5]), .A2(_zyGfifo_get_config_data_2_zyprefetch_m2_cbid[5]), .Z(n813));
Q_MX03 U4721 ( .S0(_zyM2L324_pbcFsm0_s[0]), .S1(n1132), .A0(_zyGfifo__gfdL351_25_P0_m2_cbid[4]), .A1(_zyGfifo__gfdL334_28_P0_m2_cbid[4]), .A2(_zyGfifo_get_config_data_2_zyprefetch_m2_cbid[4]), .Z(n812));
Q_MX03 U4722 ( .S0(_zyM2L324_pbcFsm0_s[0]), .S1(n1132), .A0(_zyGfifo__gfdL351_25_P0_m2_cbid[3]), .A1(_zyGfifo__gfdL334_28_P0_m2_cbid[3]), .A2(_zyGfifo_get_config_data_2_zyprefetch_m2_cbid[3]), .Z(n811));
Q_MX03 U4723 ( .S0(_zyM2L324_pbcFsm0_s[0]), .S1(n1132), .A0(_zyGfifo__gfdL351_25_P0_m2_cbid[2]), .A1(_zyGfifo__gfdL334_28_P0_m2_cbid[2]), .A2(_zyGfifo_get_config_data_2_zyprefetch_m2_cbid[2]), .Z(n810));
Q_MX03 U4724 ( .S0(_zyM2L324_pbcFsm0_s[0]), .S1(n1132), .A0(_zyGfifo__gfdL351_25_P0_m2_cbid[1]), .A1(_zyGfifo__gfdL334_28_P0_m2_cbid[1]), .A2(_zyGfifo_get_config_data_2_zyprefetch_m2_cbid[1]), .Z(n809));
Q_MX03 U4725 ( .S0(_zyM2L324_pbcFsm0_s[0]), .S1(n1132), .A0(_zyGfifo__gfdL351_25_P0_m2_cbid[0]), .A1(_zyGfifo__gfdL334_28_P0_m2_cbid[0]), .A2(_zyGfifo_get_config_data_2_zyprefetch_m2_cbid[0]), .Z(n808));
Q_MX02 U4726 ( .S(n1130), .A0(_zyGfifo__gfdL336_27_P0_m2_gfOff), .A1(_zyGfifo__gfdL327_30_P0_m2_gfOff), .Z(n550));
Q_MX02 U4727 ( .S(n1130), .A0(_zyGfifo__gfdL336_27_P0_m2_cbid[19]), .A1(_zyGfifo__gfdL327_30_P0_m2_cbid[19]), .Z(n806));
Q_MX02 U4728 ( .S(n1130), .A0(_zyGfifo__gfdL336_27_P0_m2_cbid[18]), .A1(_zyGfifo__gfdL327_30_P0_m2_cbid[18]), .Z(n805));
Q_MX02 U4729 ( .S(n1130), .A0(_zyGfifo__gfdL336_27_P0_m2_cbid[17]), .A1(_zyGfifo__gfdL327_30_P0_m2_cbid[17]), .Z(n804));
Q_MX02 U4730 ( .S(n1130), .A0(_zyGfifo__gfdL336_27_P0_m2_cbid[16]), .A1(_zyGfifo__gfdL327_30_P0_m2_cbid[16]), .Z(n803));
Q_MX02 U4731 ( .S(n1130), .A0(_zyGfifo__gfdL336_27_P0_m2_cbid[15]), .A1(_zyGfifo__gfdL327_30_P0_m2_cbid[15]), .Z(n802));
Q_MX02 U4732 ( .S(n1130), .A0(_zyGfifo__gfdL336_27_P0_m2_cbid[14]), .A1(_zyGfifo__gfdL327_30_P0_m2_cbid[14]), .Z(n801));
Q_MX02 U4733 ( .S(n1130), .A0(_zyGfifo__gfdL336_27_P0_m2_cbid[13]), .A1(_zyGfifo__gfdL327_30_P0_m2_cbid[13]), .Z(n800));
Q_MX02 U4734 ( .S(n1130), .A0(_zyGfifo__gfdL336_27_P0_m2_cbid[12]), .A1(_zyGfifo__gfdL327_30_P0_m2_cbid[12]), .Z(n799));
Q_MX02 U4735 ( .S(n1130), .A0(_zyGfifo__gfdL336_27_P0_m2_cbid[11]), .A1(_zyGfifo__gfdL327_30_P0_m2_cbid[11]), .Z(n798));
Q_MX02 U4736 ( .S(n1130), .A0(_zyGfifo__gfdL336_27_P0_m2_cbid[10]), .A1(_zyGfifo__gfdL327_30_P0_m2_cbid[10]), .Z(n797));
Q_MX02 U4737 ( .S(n1130), .A0(_zyGfifo__gfdL336_27_P0_m2_cbid[9]), .A1(_zyGfifo__gfdL327_30_P0_m2_cbid[9]), .Z(n796));
Q_MX02 U4738 ( .S(n1130), .A0(_zyGfifo__gfdL336_27_P0_m2_cbid[8]), .A1(_zyGfifo__gfdL327_30_P0_m2_cbid[8]), .Z(n795));
Q_MX02 U4739 ( .S(n1130), .A0(_zyGfifo__gfdL336_27_P0_m2_cbid[7]), .A1(_zyGfifo__gfdL327_30_P0_m2_cbid[7]), .Z(n794));
Q_MX02 U4740 ( .S(n1130), .A0(_zyGfifo__gfdL336_27_P0_m2_cbid[6]), .A1(_zyGfifo__gfdL327_30_P0_m2_cbid[6]), .Z(n793));
Q_MX02 U4741 ( .S(n1130), .A0(_zyGfifo__gfdL336_27_P0_m2_cbid[5]), .A1(_zyGfifo__gfdL327_30_P0_m2_cbid[5]), .Z(n792));
Q_MX02 U4742 ( .S(n1130), .A0(_zyGfifo__gfdL336_27_P0_m2_cbid[4]), .A1(_zyGfifo__gfdL327_30_P0_m2_cbid[4]), .Z(n791));
Q_MX02 U4743 ( .S(n1130), .A0(_zyGfifo__gfdL336_27_P0_m2_cbid[3]), .A1(_zyGfifo__gfdL327_30_P0_m2_cbid[3]), .Z(n790));
Q_MX02 U4744 ( .S(n1130), .A0(_zyGfifo__gfdL336_27_P0_m2_cbid[2]), .A1(_zyGfifo__gfdL327_30_P0_m2_cbid[2]), .Z(n789));
Q_MX02 U4745 ( .S(n1130), .A0(_zyGfifo__gfdL336_27_P0_m2_cbid[1]), .A1(_zyGfifo__gfdL327_30_P0_m2_cbid[1]), .Z(n788));
Q_MX02 U4746 ( .S(n1130), .A0(_zyGfifo__gfdL336_27_P0_m2_cbid[0]), .A1(_zyGfifo__gfdL327_30_P0_m2_cbid[0]), .Z(n787));
Q_MX02 U4747 ( .S(n1130), .A0(_zyGfifo__gfdL341_26_P0_m2_gfOff), .A1(_zyGfifo__gfdL330_29_P0_m2_gfOff), .Z(n551));
Q_AN02 U4748 ( .A0(n1130), .A1(n1151), .Z(n785));
Q_AN02 U4749 ( .A0(n1130), .A1(n1150), .Z(n784));
Q_AN02 U4750 ( .A0(n1130), .A1(n1149), .Z(n783));
Q_AN02 U4751 ( .A0(n1130), .A1(n1148), .Z(n782));
Q_AN02 U4752 ( .A0(n1130), .A1(n1147), .Z(n781));
Q_AN02 U4753 ( .A0(n1130), .A1(n1146), .Z(n780));
Q_AN02 U4754 ( .A0(n1130), .A1(n1145), .Z(n779));
Q_AN02 U4755 ( .A0(n1130), .A1(n1144), .Z(n778));
Q_MX02 U4756 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[31]), .A1(n660), .Z(n777));
Q_MX02 U4757 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[30]), .A1(n659), .Z(n776));
Q_MX02 U4758 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[29]), .A1(n658), .Z(n775));
Q_MX02 U4759 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[28]), .A1(n657), .Z(n774));
Q_MX02 U4760 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[27]), .A1(n656), .Z(n773));
Q_MX02 U4761 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[26]), .A1(n655), .Z(n772));
Q_MX02 U4762 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[25]), .A1(n654), .Z(n771));
Q_MX02 U4763 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[24]), .A1(n653), .Z(n770));
Q_MX02 U4764 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[23]), .A1(n652), .Z(n769));
Q_MX02 U4765 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[22]), .A1(n651), .Z(n768));
Q_MX02 U4766 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[21]), .A1(n650), .Z(n767));
Q_MX02 U4767 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[20]), .A1(n649), .Z(n766));
Q_MX02 U4768 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[19]), .A1(n648), .Z(n765));
Q_MX02 U4769 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[18]), .A1(n647), .Z(n764));
Q_MX02 U4770 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[17]), .A1(n646), .Z(n763));
Q_MX02 U4771 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[16]), .A1(n645), .Z(n762));
Q_MX02 U4772 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[15]), .A1(n644), .Z(n761));
Q_MX02 U4773 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[14]), .A1(n643), .Z(n760));
Q_MX02 U4774 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[13]), .A1(n642), .Z(n759));
Q_MX02 U4775 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[12]), .A1(n641), .Z(n758));
Q_MX02 U4776 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[11]), .A1(n640), .Z(n757));
Q_MX02 U4777 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[10]), .A1(n639), .Z(n756));
Q_MX02 U4778 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[9]), .A1(n638), .Z(n755));
Q_MX02 U4779 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[8]), .A1(n637), .Z(n754));
Q_MX02 U4780 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[7]), .A1(n636), .Z(n753));
Q_MX02 U4781 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[6]), .A1(n635), .Z(n752));
Q_MX02 U4782 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[5]), .A1(n634), .Z(n751));
Q_MX02 U4783 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[4]), .A1(n633), .Z(n750));
Q_MX02 U4784 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[3]), .A1(n632), .Z(n749));
Q_MX02 U4785 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[2]), .A1(n631), .Z(n748));
Q_MX02 U4786 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[1]), .A1(n630), .Z(n747));
Q_MX02 U4787 ( .S(n1130), .A0(_zyL94_iscX1c0_o1[0]), .A1(n629), .Z(n746));
Q_MX02 U4788 ( .S(n1130), .A0(data[31]), .A1(n692), .Z(n745));
Q_MX02 U4789 ( .S(n1130), .A0(data[30]), .A1(n691), .Z(n744));
Q_MX02 U4790 ( .S(n1130), .A0(data[29]), .A1(n690), .Z(n743));
Q_MX02 U4791 ( .S(n1130), .A0(data[28]), .A1(n689), .Z(n742));
Q_MX02 U4792 ( .S(n1130), .A0(data[27]), .A1(n688), .Z(n741));
Q_MX02 U4793 ( .S(n1130), .A0(data[26]), .A1(n687), .Z(n740));
Q_MX02 U4794 ( .S(n1130), .A0(data[25]), .A1(n686), .Z(n739));
Q_MX02 U4795 ( .S(n1130), .A0(data[24]), .A1(n685), .Z(n738));
Q_MX02 U4796 ( .S(n1130), .A0(data[23]), .A1(n684), .Z(n737));
Q_MX02 U4797 ( .S(n1130), .A0(data[22]), .A1(n683), .Z(n736));
Q_MX02 U4798 ( .S(n1130), .A0(data[21]), .A1(n682), .Z(n735));
Q_MX02 U4799 ( .S(n1130), .A0(data[20]), .A1(n681), .Z(n734));
Q_MX02 U4800 ( .S(n1130), .A0(data[19]), .A1(n680), .Z(n733));
Q_MX02 U4801 ( .S(n1130), .A0(data[18]), .A1(n679), .Z(n732));
Q_MX02 U4802 ( .S(n1130), .A0(data[17]), .A1(n678), .Z(n731));
Q_MX02 U4803 ( .S(n1130), .A0(data[16]), .A1(n677), .Z(n730));
Q_MX02 U4804 ( .S(n1130), .A0(data[15]), .A1(n676), .Z(n729));
Q_MX02 U4805 ( .S(n1130), .A0(data[14]), .A1(n675), .Z(n728));
Q_MX02 U4806 ( .S(n1130), .A0(data[13]), .A1(n674), .Z(n727));
Q_MX02 U4807 ( .S(n1130), .A0(data[12]), .A1(n673), .Z(n726));
Q_MX02 U4808 ( .S(n1130), .A0(data[11]), .A1(n672), .Z(n725));
Q_MX02 U4809 ( .S(n1130), .A0(data[10]), .A1(n671), .Z(n724));
Q_MX02 U4810 ( .S(n1130), .A0(data[9]), .A1(n670), .Z(n723));
Q_MX02 U4811 ( .S(n1130), .A0(data[8]), .A1(n669), .Z(n722));
Q_MX02 U4812 ( .S(n1130), .A0(data[7]), .A1(n668), .Z(n721));
Q_MX02 U4813 ( .S(n1130), .A0(data[6]), .A1(n667), .Z(n720));
Q_MX02 U4814 ( .S(n1130), .A0(data[5]), .A1(n666), .Z(n719));
Q_MX02 U4815 ( .S(n1130), .A0(data[4]), .A1(n665), .Z(n718));
Q_MX02 U4816 ( .S(n1130), .A0(data[3]), .A1(n664), .Z(n717));
Q_MX02 U4817 ( .S(n1130), .A0(data[2]), .A1(n663), .Z(n716));
Q_MX02 U4818 ( .S(n1130), .A0(data[1]), .A1(n662), .Z(n715));
Q_MX02 U4819 ( .S(n1130), .A0(data[0]), .A1(n661), .Z(n714));
Q_MX02 U4820 ( .S(n1130), .A0(_zyGfifo__gfdL341_26_P0_m2_cbid[19]), .A1(_zyGfifo__gfdL330_29_P0_m2_cbid[19]), .Z(n713));
Q_MX02 U4821 ( .S(n1130), .A0(_zyGfifo__gfdL341_26_P0_m2_cbid[18]), .A1(_zyGfifo__gfdL330_29_P0_m2_cbid[18]), .Z(n712));
Q_MX02 U4822 ( .S(n1130), .A0(_zyGfifo__gfdL341_26_P0_m2_cbid[17]), .A1(_zyGfifo__gfdL330_29_P0_m2_cbid[17]), .Z(n711));
Q_MX02 U4823 ( .S(n1130), .A0(_zyGfifo__gfdL341_26_P0_m2_cbid[16]), .A1(_zyGfifo__gfdL330_29_P0_m2_cbid[16]), .Z(n710));
Q_MX02 U4824 ( .S(n1130), .A0(_zyGfifo__gfdL341_26_P0_m2_cbid[15]), .A1(_zyGfifo__gfdL330_29_P0_m2_cbid[15]), .Z(n709));
Q_MX02 U4825 ( .S(n1130), .A0(_zyGfifo__gfdL341_26_P0_m2_cbid[14]), .A1(_zyGfifo__gfdL330_29_P0_m2_cbid[14]), .Z(n708));
Q_MX02 U4826 ( .S(n1130), .A0(_zyGfifo__gfdL341_26_P0_m2_cbid[13]), .A1(_zyGfifo__gfdL330_29_P0_m2_cbid[13]), .Z(n707));
Q_MX02 U4827 ( .S(n1130), .A0(_zyGfifo__gfdL341_26_P0_m2_cbid[12]), .A1(_zyGfifo__gfdL330_29_P0_m2_cbid[12]), .Z(n706));
Q_MX02 U4828 ( .S(n1130), .A0(_zyGfifo__gfdL341_26_P0_m2_cbid[11]), .A1(_zyGfifo__gfdL330_29_P0_m2_cbid[11]), .Z(n705));
Q_MX02 U4829 ( .S(n1130), .A0(_zyGfifo__gfdL341_26_P0_m2_cbid[10]), .A1(_zyGfifo__gfdL330_29_P0_m2_cbid[10]), .Z(n704));
Q_MX02 U4830 ( .S(n1130), .A0(_zyGfifo__gfdL341_26_P0_m2_cbid[9]), .A1(_zyGfifo__gfdL330_29_P0_m2_cbid[9]), .Z(n703));
Q_MX02 U4831 ( .S(n1130), .A0(_zyGfifo__gfdL341_26_P0_m2_cbid[8]), .A1(_zyGfifo__gfdL330_29_P0_m2_cbid[8]), .Z(n702));
Q_MX02 U4832 ( .S(n1130), .A0(_zyGfifo__gfdL341_26_P0_m2_cbid[7]), .A1(_zyGfifo__gfdL330_29_P0_m2_cbid[7]), .Z(n701));
Q_MX02 U4833 ( .S(n1130), .A0(_zyGfifo__gfdL341_26_P0_m2_cbid[6]), .A1(_zyGfifo__gfdL330_29_P0_m2_cbid[6]), .Z(n700));
Q_MX02 U4834 ( .S(n1130), .A0(_zyGfifo__gfdL341_26_P0_m2_cbid[5]), .A1(_zyGfifo__gfdL330_29_P0_m2_cbid[5]), .Z(n699));
Q_MX02 U4835 ( .S(n1130), .A0(_zyGfifo__gfdL341_26_P0_m2_cbid[4]), .A1(_zyGfifo__gfdL330_29_P0_m2_cbid[4]), .Z(n698));
Q_MX02 U4836 ( .S(n1130), .A0(_zyGfifo__gfdL341_26_P0_m2_cbid[3]), .A1(_zyGfifo__gfdL330_29_P0_m2_cbid[3]), .Z(n697));
Q_MX02 U4837 ( .S(n1130), .A0(_zyGfifo__gfdL341_26_P0_m2_cbid[2]), .A1(_zyGfifo__gfdL330_29_P0_m2_cbid[2]), .Z(n696));
Q_MX02 U4838 ( .S(n1130), .A0(_zyGfifo__gfdL341_26_P0_m2_cbid[1]), .A1(_zyGfifo__gfdL330_29_P0_m2_cbid[1]), .Z(n695));
Q_MX02 U4839 ( .S(n1130), .A0(_zyGfifo__gfdL341_26_P0_m2_cbid[0]), .A1(_zyGfifo__gfdL330_29_P0_m2_cbid[0]), .Z(n694));
Q_MX02 U4840 ( .S(_zyM2L324_pbcFsm0_s[0]), .A0(_zyL61_iscX2c0_o2), .A1(_zyL94_iscX1c0_o2), .Z(n693));
Q_MX02 U4841 ( .S(n500), .A0(n1091), .A1(_zydata_L206_tfiV2_M2_pbcG2[31]), .Z(n692));
Q_MX02 U4842 ( .S(n500), .A0(n1092), .A1(_zydata_L206_tfiV2_M2_pbcG2[30]), .Z(n691));
Q_MX02 U4843 ( .S(n500), .A0(n1093), .A1(_zydata_L206_tfiV2_M2_pbcG2[29]), .Z(n690));
Q_MX02 U4844 ( .S(n500), .A0(n1094), .A1(_zydata_L206_tfiV2_M2_pbcG2[28]), .Z(n689));
Q_MX02 U4845 ( .S(n500), .A0(n1095), .A1(_zydata_L206_tfiV2_M2_pbcG2[27]), .Z(n688));
Q_MX02 U4846 ( .S(n500), .A0(n1096), .A1(_zydata_L206_tfiV2_M2_pbcG2[26]), .Z(n687));
Q_MX02 U4847 ( .S(n500), .A0(n1097), .A1(_zydata_L206_tfiV2_M2_pbcG2[25]), .Z(n686));
Q_MX02 U4848 ( .S(n500), .A0(n1098), .A1(_zydata_L206_tfiV2_M2_pbcG2[24]), .Z(n685));
Q_MX02 U4849 ( .S(n500), .A0(n1099), .A1(_zydata_L206_tfiV2_M2_pbcG2[23]), .Z(n684));
Q_MX02 U4850 ( .S(n500), .A0(n1100), .A1(_zydata_L206_tfiV2_M2_pbcG2[22]), .Z(n683));
Q_MX02 U4851 ( .S(n500), .A0(n1101), .A1(_zydata_L206_tfiV2_M2_pbcG2[21]), .Z(n682));
Q_MX02 U4852 ( .S(n500), .A0(n1102), .A1(_zydata_L206_tfiV2_M2_pbcG2[20]), .Z(n681));
Q_MX02 U4853 ( .S(n500), .A0(n1103), .A1(_zydata_L206_tfiV2_M2_pbcG2[19]), .Z(n680));
Q_MX02 U4854 ( .S(n500), .A0(n1104), .A1(_zydata_L206_tfiV2_M2_pbcG2[18]), .Z(n679));
Q_MX02 U4855 ( .S(n500), .A0(n1105), .A1(_zydata_L206_tfiV2_M2_pbcG2[17]), .Z(n678));
Q_MX02 U4856 ( .S(n500), .A0(n1106), .A1(_zydata_L206_tfiV2_M2_pbcG2[16]), .Z(n677));
Q_MX02 U4857 ( .S(n500), .A0(n1107), .A1(_zydata_L206_tfiV2_M2_pbcG2[15]), .Z(n676));
Q_MX02 U4858 ( .S(n500), .A0(n1108), .A1(_zydata_L206_tfiV2_M2_pbcG2[14]), .Z(n675));
Q_MX02 U4859 ( .S(n500), .A0(n1109), .A1(_zydata_L206_tfiV2_M2_pbcG2[13]), .Z(n674));
Q_MX02 U4860 ( .S(n500), .A0(n1110), .A1(_zydata_L206_tfiV2_M2_pbcG2[12]), .Z(n673));
Q_MX02 U4861 ( .S(n500), .A0(n1111), .A1(_zydata_L206_tfiV2_M2_pbcG2[11]), .Z(n672));
Q_MX02 U4862 ( .S(n500), .A0(n1112), .A1(_zydata_L206_tfiV2_M2_pbcG2[10]), .Z(n671));
Q_MX02 U4863 ( .S(n500), .A0(n1113), .A1(_zydata_L206_tfiV2_M2_pbcG2[9]), .Z(n670));
Q_MX02 U4864 ( .S(n500), .A0(n1114), .A1(_zydata_L206_tfiV2_M2_pbcG2[8]), .Z(n669));
Q_MX02 U4865 ( .S(n500), .A0(n1115), .A1(_zydata_L206_tfiV2_M2_pbcG2[7]), .Z(n668));
Q_MX02 U4866 ( .S(n500), .A0(n1116), .A1(_zydata_L206_tfiV2_M2_pbcG2[6]), .Z(n667));
Q_MX02 U4867 ( .S(n500), .A0(n1117), .A1(_zydata_L206_tfiV2_M2_pbcG2[5]), .Z(n666));
Q_MX02 U4868 ( .S(n500), .A0(n1118), .A1(_zydata_L206_tfiV2_M2_pbcG2[4]), .Z(n665));
Q_MX02 U4869 ( .S(n500), .A0(n1119), .A1(_zydata_L206_tfiV2_M2_pbcG2[3]), .Z(n664));
Q_MX02 U4870 ( .S(n500), .A0(n1120), .A1(_zydata_L206_tfiV2_M2_pbcG2[2]), .Z(n663));
Q_MX02 U4871 ( .S(n500), .A0(n1121), .A1(_zydata_L206_tfiV2_M2_pbcG2[1]), .Z(n662));
Q_MX02 U4872 ( .S(n500), .A0(n1122), .A1(_zydata_L206_tfiV2_M2_pbcG2[0]), .Z(n661));
Q_MX02 U4873 ( .S(n500), .A0(n1059), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[31]), .Z(n660));
Q_MX02 U4874 ( .S(n500), .A0(n1060), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[30]), .Z(n659));
Q_MX02 U4875 ( .S(n500), .A0(n1061), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[29]), .Z(n658));
Q_MX02 U4876 ( .S(n500), .A0(n1062), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[28]), .Z(n657));
Q_MX02 U4877 ( .S(n500), .A0(n1063), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[27]), .Z(n656));
Q_MX02 U4878 ( .S(n500), .A0(n1064), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[26]), .Z(n655));
Q_MX02 U4879 ( .S(n500), .A0(n1065), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[25]), .Z(n654));
Q_MX02 U4880 ( .S(n500), .A0(n1066), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[24]), .Z(n653));
Q_MX02 U4881 ( .S(n500), .A0(n1067), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[23]), .Z(n652));
Q_MX02 U4882 ( .S(n500), .A0(n1068), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[22]), .Z(n651));
Q_MX02 U4883 ( .S(n500), .A0(n1069), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[21]), .Z(n650));
Q_MX02 U4884 ( .S(n500), .A0(n1070), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[20]), .Z(n649));
Q_MX02 U4885 ( .S(n500), .A0(n1071), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[19]), .Z(n648));
Q_MX02 U4886 ( .S(n500), .A0(n1072), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[18]), .Z(n647));
Q_MX02 U4887 ( .S(n500), .A0(n1073), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[17]), .Z(n646));
Q_MX02 U4888 ( .S(n500), .A0(n1074), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[16]), .Z(n645));
Q_MX02 U4889 ( .S(n500), .A0(n1075), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[15]), .Z(n644));
Q_MX02 U4890 ( .S(n500), .A0(n1076), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[14]), .Z(n643));
Q_MX02 U4891 ( .S(n500), .A0(n1077), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[13]), .Z(n642));
Q_MX02 U4892 ( .S(n500), .A0(n1078), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[12]), .Z(n641));
Q_MX02 U4893 ( .S(n500), .A0(n1079), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[11]), .Z(n640));
Q_MX02 U4894 ( .S(n500), .A0(n1080), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[10]), .Z(n639));
Q_MX02 U4895 ( .S(n500), .A0(n1081), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[9]), .Z(n638));
Q_MX02 U4896 ( .S(n500), .A0(n1082), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[8]), .Z(n637));
Q_MX02 U4897 ( .S(n500), .A0(n1083), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[7]), .Z(n636));
Q_MX02 U4898 ( .S(n500), .A0(n1084), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[6]), .Z(n635));
Q_MX02 U4899 ( .S(n500), .A0(n1085), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[5]), .Z(n634));
Q_MX02 U4900 ( .S(n500), .A0(n1086), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[4]), .Z(n633));
Q_MX02 U4901 ( .S(n500), .A0(n1087), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[3]), .Z(n632));
Q_MX02 U4902 ( .S(n500), .A0(n1088), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[2]), .Z(n631));
Q_MX02 U4903 ( .S(n500), .A0(n1089), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[1]), .Z(n630));
Q_MX02 U4904 ( .S(n500), .A0(n1090), .A1(_zyaddress_L206_tfiV1_M2_pbcG1[0]), .Z(n629));
Q_MX02 U4905 ( .S(n500), .A0(n1051), .A1(_zyoperation_L206_tfiV0_M2_pbcG0[7]), .Z(n1151));
Q_MX02 U4906 ( .S(n500), .A0(n1052), .A1(_zyoperation_L206_tfiV0_M2_pbcG0[6]), .Z(n1150));
Q_MX02 U4907 ( .S(n500), .A0(n1053), .A1(_zyoperation_L206_tfiV0_M2_pbcG0[5]), .Z(n1149));
Q_MX02 U4908 ( .S(n500), .A0(n1054), .A1(_zyoperation_L206_tfiV0_M2_pbcG0[4]), .Z(n1148));
Q_MX02 U4909 ( .S(n500), .A0(n1055), .A1(_zyoperation_L206_tfiV0_M2_pbcG0[3]), .Z(n1147));
Q_MX02 U4910 ( .S(n500), .A0(n1056), .A1(_zyoperation_L206_tfiV0_M2_pbcG0[2]), .Z(n1146));
Q_MX02 U4911 ( .S(n500), .A0(n1057), .A1(_zyoperation_L206_tfiV0_M2_pbcG0[1]), .Z(n1145));
Q_MX02 U4912 ( .S(n500), .A0(n1058), .A1(_zyoperation_L206_tfiV0_M2_pbcG0[0]), .Z(n1144));
Q_INV U4913 ( .A(n628), .Z(n1141));
Q_NR02 U4914 ( .A0(n627), .A1(n626), .Z(n628));
Q_MX02 U4915 ( .S(n1124), .A0(n622), .A1(n614), .Z(n627));
Q_MX02 U4916 ( .S(n1124), .A0(n621), .A1(n617), .Z(n626));
Q_MX02 U4917 ( .S(n1124), .A0(n620), .A1(n616), .Z(n625));
Q_MX02 U4918 ( .S(n1124), .A0(n619), .A1(n615), .Z(n624));
Q_MX02 U4919 ( .S(n1124), .A0(n618), .A1(n607), .Z(n623));
Q_MX02 U4920 ( .S(n500), .A0(n584), .A1(_zygsfis_get_config_data_space[3]), .Z(n621));
Q_MX02 U4921 ( .S(n500), .A0(n582), .A1(_zygsfis_get_config_data_space[2]), .Z(n620));
Q_MX02 U4922 ( .S(n500), .A0(n580), .A1(_zygsfis_get_config_data_space[1]), .Z(n619));
Q_XOR2 U4923 ( .A0(n1123), .A1(_zygsfis_get_config_data_space[0]), .Z(n618));
Q_INV U4924 ( .A(n612), .Z(n617));
Q_INV U4925 ( .A(n611), .Z(n616));
Q_INV U4926 ( .A(n609), .Z(n615));
Q_AD02 U4927 ( .CI(n610), .A0(_zygsfis_get_config_data_wptr[2]), .A1(_zygsfis_get_config_data_wptr[3]), .B0(n605), .B1(n606), .S0(n611), .S1(n612), .CO(n613));
Q_AD01 U4928 ( .CI(n604), .A0(_zygsfis_get_config_data_wptr[1]), .B0(n608), .S(n609), .CO(n610));
Q_OR02 U4929 ( .A0(_zygsfis_get_config_data_wptr[0]), .A1(n603), .Z(n608));
Q_XOR2 U4930 ( .A0(_zygsfis_get_config_data_wptr[0]), .A1(n603), .Z(n607));
Q_XOR3 U4931 ( .A0(_zygsfis_get_config_data_wptr[4]), .A1(n596), .A2(n613), .Z(n614));
Q_INV U4932 ( .A(n595), .Z(n606));
Q_INV U4933 ( .A(n594), .Z(n605));
Q_INV U4934 ( .A(n593), .Z(n604));
Q_INV U4935 ( .A(n592), .Z(n603));
Q_AN02 U4936 ( .A0(n602), .A1(_zygsfis_get_config_data_eos), .Z(n1133));
Q_AN03 U4937 ( .A0(n599), .A1(n600), .A2(n601), .Z(n602));
Q_AN03 U4938 ( .A0(n607), .A1(n597), .A2(n598), .Z(n601));
Q_XNR2 U4939 ( .A0(n596), .A1(_zygsfis_get_config_data_wptr[4]), .Z(n600));
Q_XNR2 U4940 ( .A0(n595), .A1(_zygsfis_get_config_data_wptr[3]), .Z(n599));
Q_XNR2 U4941 ( .A0(n594), .A1(_zygsfis_get_config_data_wptr[2]), .Z(n598));
Q_XNR2 U4942 ( .A0(n593), .A1(_zygsfis_get_config_data_wptr[1]), .Z(n597));
Q_MX02 U4943 ( .S(n500), .A0(n590), .A1(_zygsfis_get_config_data_rptr[3]), .Z(n595));
Q_MX02 U4944 ( .S(n500), .A0(n588), .A1(_zygsfis_get_config_data_rptr[2]), .Z(n594));
Q_MX02 U4945 ( .S(n500), .A0(n586), .A1(_zygsfis_get_config_data_rptr[1]), .Z(n593));
Q_XOR2 U4946 ( .A0(n1123), .A1(_zygsfis_get_config_data_rptr[0]), .Z(n592));
Q_XOR2 U4947 ( .A0(_zygsfis_get_config_data_rptr[4]), .A1(n5886), .Z(n596));
Q_AD01HF U4948 ( .A0(_zygsfis_get_config_data_rptr[3]), .B0(n589), .S(n590), .CO(n591));
Q_AD01HF U4949 ( .A0(_zygsfis_get_config_data_rptr[2]), .B0(n587), .S(n588), .CO(n589));
Q_AD01HF U4950 ( .A0(_zygsfis_get_config_data_rptr[1]), .B0(_zygsfis_get_config_data_rptr[0]), .S(n586), .CO(n587));
Q_XOR2 U4951 ( .A0(_zygsfis_get_config_data_space[4]), .A1(n5885), .Z(n622));
Q_AD01HF U4952 ( .A0(_zygsfis_get_config_data_space[3]), .B0(n583), .S(n584), .CO(n585));
Q_AD01HF U4953 ( .A0(_zygsfis_get_config_data_space[2]), .B0(n581), .S(n582), .CO(n583));
Q_AD01HF U4954 ( .A0(_zygsfis_get_config_data_space[1]), .B0(_zygsfis_get_config_data_space[0]), .S(n580), .CO(n581));
Q_AD01HF U4955 ( .A0(_zygsfis_get_config_data_req[3]), .B0(n577), .S(n578), .CO(n579));
Q_AD01HF U4956 ( .A0(_zygsfis_get_config_data_req[2]), .B0(n575), .S(n576), .CO(n577));
Q_AD01HF U4957 ( .A0(_zygsfis_get_config_data_req[1]), .B0(_zygsfis_get_config_data_req[0]), .S(n574), .CO(n575));
Q_AN03 U4958 ( .A0(n572), .A1(n573), .A2(n1143), .Z(n1020));
Q_INV U4959 ( .A(n2261), .Z(n573));
Q_OR03 U4960 ( .A0(n571), .A1(n570), .A2(n569), .Z(n572));
Q_AO21 U4961 ( .A0(n2205), .A1(n567), .B0(n566), .Z(n570));
Q_OR03 U4962 ( .A0(n555), .A1(n557), .A2(n568), .Z(n569));
Q_AO21 U4963 ( .A0(n2201), .A1(n553), .B0(n2203), .Z(n567));
Q_OR03 U4964 ( .A0(n2211), .A1(n2209), .A2(n2207), .Z(n566));
Q_OR03 U4965 ( .A0(n565), .A1(n564), .A2(n563), .Z(n571));
Q_OR02 U4966 ( .A0(n2219), .A1(n2217), .Z(n565));
Q_OR02 U4967 ( .A0(n2215), .A1(n2213), .Z(n564));
Q_OR03 U4968 ( .A0(n2227), .A1(n2225), .A2(n562), .Z(n563));
Q_OR02 U4969 ( .A0(n2223), .A1(n2221), .Z(n562));
Q_OR03 U4970 ( .A0(n561), .A1(n560), .A2(n559), .Z(n568));
Q_OR02 U4971 ( .A0(n2235), .A1(n2233), .Z(n561));
Q_OR02 U4972 ( .A0(n2231), .A1(n2229), .Z(n560));
Q_OR03 U4973 ( .A0(n2243), .A1(n2241), .A2(n558), .Z(n559));
Q_OR02 U4974 ( .A0(n2239), .A1(n2237), .Z(n558));
Q_OR03 U4975 ( .A0(n2251), .A1(n2249), .A2(n556), .Z(n557));
Q_OR02 U4976 ( .A0(n2247), .A1(n2245), .Z(n556));
Q_OR03 U4977 ( .A0(n2259), .A1(n2257), .A2(n554), .Z(n555));
Q_OR02 U4978 ( .A0(n2255), .A1(n2253), .Z(n554));
Q_XNR2 U4979 ( .A0(n552), .A1(_zyGfifoF0_L324_s3_req_1), .Z(n921));
Q_XNR2 U4980 ( .A0(n551), .A1(_zyGfifoF2_L324_s2_req_3), .Z(n786));
Q_XNR2 U4981 ( .A0(n550), .A1(_zyGfifoF1_L324_s2_req_2), .Z(n807));
Q_XNR2 U4982 ( .A0(_zyGfifo_get_config_data_2_zyprefetch_m2_gfOff), .A1(_zyGfifoF0_L324_s3_req_1), .Z(n549));
Q_INV U4983 ( .A(n548), .Z(n1143));
Q_AN02 U4984 ( .A0(n546), .A1(n547), .Z(n548));
Q_AN03 U4985 ( .A0(n543), .A1(n544), .A2(n545), .Z(n547));
Q_AN03 U4986 ( .A0(n540), .A1(n541), .A2(n542), .Z(n546));
Q_AN03 U4987 ( .A0(n537), .A1(n538), .A2(n539), .Z(n545));
Q_AN03 U4988 ( .A0(n534), .A1(n535), .A2(n536), .Z(n544));
Q_AN03 U4989 ( .A0(n502), .A1(n501), .A2(n533), .Z(n543));
Q_AN03 U4990 ( .A0(n505), .A1(n504), .A2(n503), .Z(n542));
Q_AN03 U4991 ( .A0(n508), .A1(n507), .A2(n506), .Z(n541));
Q_AN03 U4992 ( .A0(n511), .A1(n510), .A2(n509), .Z(n540));
Q_AN03 U4993 ( .A0(n514), .A1(n513), .A2(n512), .Z(n539));
Q_AN03 U4994 ( .A0(n517), .A1(n516), .A2(n515), .Z(n538));
Q_AN03 U4995 ( .A0(n520), .A1(n519), .A2(n518), .Z(n537));
Q_AN03 U4996 ( .A0(n523), .A1(n522), .A2(n521), .Z(n536));
Q_AN03 U4997 ( .A0(n526), .A1(n525), .A2(n524), .Z(n535));
Q_AN03 U4998 ( .A0(n529), .A1(n528), .A2(n527), .Z(n534));
Q_AN03 U4999 ( .A0(n532), .A1(n531), .A2(n530), .Z(n533));
Q_XNR2 U5000 ( .A0(_zyL94_iscX1c0_o1[31]), .A1(data[31]), .Z(n532));
Q_XNR2 U5001 ( .A0(_zyL94_iscX1c0_o1[30]), .A1(data[30]), .Z(n531));
Q_XNR2 U5002 ( .A0(_zyL94_iscX1c0_o1[29]), .A1(data[29]), .Z(n530));
Q_XNR2 U5003 ( .A0(_zyL94_iscX1c0_o1[28]), .A1(data[28]), .Z(n529));
Q_XNR2 U5004 ( .A0(_zyL94_iscX1c0_o1[27]), .A1(data[27]), .Z(n528));
Q_XNR2 U5005 ( .A0(_zyL94_iscX1c0_o1[26]), .A1(data[26]), .Z(n527));
Q_XNR2 U5006 ( .A0(_zyL94_iscX1c0_o1[25]), .A1(data[25]), .Z(n526));
Q_XNR2 U5007 ( .A0(_zyL94_iscX1c0_o1[24]), .A1(data[24]), .Z(n525));
Q_XNR2 U5008 ( .A0(_zyL94_iscX1c0_o1[23]), .A1(data[23]), .Z(n524));
Q_XNR2 U5009 ( .A0(_zyL94_iscX1c0_o1[22]), .A1(data[22]), .Z(n523));
Q_XNR2 U5010 ( .A0(_zyL94_iscX1c0_o1[21]), .A1(data[21]), .Z(n522));
Q_XNR2 U5011 ( .A0(_zyL94_iscX1c0_o1[20]), .A1(data[20]), .Z(n521));
Q_XNR2 U5012 ( .A0(_zyL94_iscX1c0_o1[19]), .A1(data[19]), .Z(n520));
Q_XNR2 U5013 ( .A0(_zyL94_iscX1c0_o1[18]), .A1(data[18]), .Z(n519));
Q_XNR2 U5014 ( .A0(_zyL94_iscX1c0_o1[17]), .A1(data[17]), .Z(n518));
Q_XNR2 U5015 ( .A0(_zyL94_iscX1c0_o1[16]), .A1(data[16]), .Z(n517));
Q_XNR2 U5016 ( .A0(_zyL94_iscX1c0_o1[15]), .A1(data[15]), .Z(n516));
Q_XNR2 U5017 ( .A0(_zyL94_iscX1c0_o1[14]), .A1(data[14]), .Z(n515));
Q_XNR2 U5018 ( .A0(_zyL94_iscX1c0_o1[13]), .A1(data[13]), .Z(n514));
Q_XNR2 U5019 ( .A0(_zyL94_iscX1c0_o1[12]), .A1(data[12]), .Z(n513));
Q_XNR2 U5020 ( .A0(_zyL94_iscX1c0_o1[11]), .A1(data[11]), .Z(n512));
Q_XNR2 U5021 ( .A0(_zyL94_iscX1c0_o1[10]), .A1(data[10]), .Z(n511));
Q_XNR2 U5022 ( .A0(_zyL94_iscX1c0_o1[9]), .A1(data[9]), .Z(n510));
Q_XNR2 U5023 ( .A0(_zyL94_iscX1c0_o1[8]), .A1(data[8]), .Z(n509));
Q_XNR2 U5024 ( .A0(_zyL94_iscX1c0_o1[7]), .A1(data[7]), .Z(n508));
Q_XNR2 U5025 ( .A0(_zyL94_iscX1c0_o1[6]), .A1(data[6]), .Z(n507));
Q_XNR2 U5026 ( .A0(_zyL94_iscX1c0_o1[5]), .A1(data[5]), .Z(n506));
Q_XNR2 U5027 ( .A0(_zyL94_iscX1c0_o1[4]), .A1(data[4]), .Z(n505));
Q_XNR2 U5028 ( .A0(_zyL94_iscX1c0_o1[3]), .A1(data[3]), .Z(n504));
Q_XNR2 U5029 ( .A0(_zyL94_iscX1c0_o1[2]), .A1(data[2]), .Z(n503));
Q_XNR2 U5030 ( .A0(_zyL94_iscX1c0_o1[1]), .A1(data[1]), .Z(n502));
Q_XNR2 U5031 ( .A0(_zyL94_iscX1c0_o1[0]), .A1(data[0]), .Z(n501));
Q_INV U5032 ( .A(n500), .Z(n1123));
Q_AN03 U5033 ( .A0(n495), .A1(n494), .A2(n499), .Z(n500));
Q_AN03 U5034 ( .A0(n498), .A1(n497), .A2(n496), .Z(n499));
Q_XNR2 U5035 ( .A0(_zygsfis_get_config_data_rptr[4]), .A1(_zygsfis_get_config_data_wptr[4]), .Z(n498));
Q_XNR2 U5036 ( .A0(_zygsfis_get_config_data_rptr[3]), .A1(_zygsfis_get_config_data_wptr[3]), .Z(n497));
Q_XNR2 U5037 ( .A0(_zygsfis_get_config_data_rptr[2]), .A1(_zygsfis_get_config_data_wptr[2]), .Z(n496));
Q_XNR2 U5038 ( .A0(_zygsfis_get_config_data_rptr[1]), .A1(_zygsfis_get_config_data_wptr[1]), .Z(n495));
Q_XNR2 U5039 ( .A0(_zygsfis_get_config_data_rptr[0]), .A1(_zygsfis_get_config_data_wptr[0]), .Z(n494));
Q_AN03 U5040 ( .A0(n489), .A1(n488), .A2(n493), .Z(n1124));
Q_AN03 U5041 ( .A0(n492), .A1(n491), .A2(n490), .Z(n493));
Q_XNR2 U5042 ( .A0(_zygsfis_get_config_data_req[4]), .A1(_zygsfis_get_config_data_ack[4]), .Z(n492));
Q_XNR2 U5043 ( .A0(_zygsfis_get_config_data_req[3]), .A1(_zygsfis_get_config_data_ack[3]), .Z(n491));
Q_XNR2 U5044 ( .A0(_zygsfis_get_config_data_req[2]), .A1(_zygsfis_get_config_data_ack[2]), .Z(n490));
Q_XNR2 U5045 ( .A0(_zygsfis_get_config_data_req[1]), .A1(_zygsfis_get_config_data_ack[1]), .Z(n489));
Q_XNR2 U5046 ( .A0(_zygsfis_get_config_data_req[0]), .A1(_zygsfis_get_config_data_ack[0]), .Z(n488));
Q_AN02 U5047 ( .A0(n485), .A1(config_done), .Z(n487));
Q_FDP0 \_zyL312_meState2_REG[0] ( .CK(clk), .D(n487), .Q(_zyL312_meState2[0]), .QN(n485));
Q_MX02 U5049 ( .S(n486), .A0(_zyGfifo__gfdL318_31_P0_m2_gfOff), .A1(_zyGfifo__gfdL316_32_P0_m2_gfOff), .Z(n463));
Q_MX02 U5050 ( .S(n486), .A0(_zyGfifo__gfdL318_31_P0_m2_cbid[19]), .A1(_zyGfifo__gfdL316_32_P0_m2_cbid[19]), .Z(n483));
Q_MX02 U5051 ( .S(n486), .A0(_zyGfifo__gfdL318_31_P0_m2_cbid[18]), .A1(_zyGfifo__gfdL316_32_P0_m2_cbid[18]), .Z(n482));
Q_MX02 U5052 ( .S(n486), .A0(_zyGfifo__gfdL318_31_P0_m2_cbid[17]), .A1(_zyGfifo__gfdL316_32_P0_m2_cbid[17]), .Z(n481));
Q_MX02 U5053 ( .S(n486), .A0(_zyGfifo__gfdL318_31_P0_m2_cbid[16]), .A1(_zyGfifo__gfdL316_32_P0_m2_cbid[16]), .Z(n480));
Q_MX02 U5054 ( .S(n486), .A0(_zyGfifo__gfdL318_31_P0_m2_cbid[15]), .A1(_zyGfifo__gfdL316_32_P0_m2_cbid[15]), .Z(n479));
Q_MX02 U5055 ( .S(n486), .A0(_zyGfifo__gfdL318_31_P0_m2_cbid[14]), .A1(_zyGfifo__gfdL316_32_P0_m2_cbid[14]), .Z(n478));
Q_MX02 U5056 ( .S(n486), .A0(_zyGfifo__gfdL318_31_P0_m2_cbid[13]), .A1(_zyGfifo__gfdL316_32_P0_m2_cbid[13]), .Z(n477));
Q_MX02 U5057 ( .S(n486), .A0(_zyGfifo__gfdL318_31_P0_m2_cbid[12]), .A1(_zyGfifo__gfdL316_32_P0_m2_cbid[12]), .Z(n476));
Q_MX02 U5058 ( .S(n486), .A0(_zyGfifo__gfdL318_31_P0_m2_cbid[11]), .A1(_zyGfifo__gfdL316_32_P0_m2_cbid[11]), .Z(n475));
Q_MX02 U5059 ( .S(n486), .A0(_zyGfifo__gfdL318_31_P0_m2_cbid[10]), .A1(_zyGfifo__gfdL316_32_P0_m2_cbid[10]), .Z(n474));
Q_MX02 U5060 ( .S(n486), .A0(_zyGfifo__gfdL318_31_P0_m2_cbid[9]), .A1(_zyGfifo__gfdL316_32_P0_m2_cbid[9]), .Z(n473));
Q_MX02 U5061 ( .S(n486), .A0(_zyGfifo__gfdL318_31_P0_m2_cbid[8]), .A1(_zyGfifo__gfdL316_32_P0_m2_cbid[8]), .Z(n472));
Q_MX02 U5062 ( .S(n486), .A0(_zyGfifo__gfdL318_31_P0_m2_cbid[7]), .A1(_zyGfifo__gfdL316_32_P0_m2_cbid[7]), .Z(n471));
Q_MX02 U5063 ( .S(n486), .A0(_zyGfifo__gfdL318_31_P0_m2_cbid[6]), .A1(_zyGfifo__gfdL316_32_P0_m2_cbid[6]), .Z(n470));
Q_MX02 U5064 ( .S(n486), .A0(_zyGfifo__gfdL318_31_P0_m2_cbid[5]), .A1(_zyGfifo__gfdL316_32_P0_m2_cbid[5]), .Z(n469));
Q_MX02 U5065 ( .S(n486), .A0(_zyGfifo__gfdL318_31_P0_m2_cbid[4]), .A1(_zyGfifo__gfdL316_32_P0_m2_cbid[4]), .Z(n468));
Q_MX02 U5066 ( .S(n486), .A0(_zyGfifo__gfdL318_31_P0_m2_cbid[3]), .A1(_zyGfifo__gfdL316_32_P0_m2_cbid[3]), .Z(n467));
Q_MX02 U5067 ( .S(n486), .A0(_zyGfifo__gfdL318_31_P0_m2_cbid[2]), .A1(_zyGfifo__gfdL316_32_P0_m2_cbid[2]), .Z(n466));
Q_MX02 U5068 ( .S(n486), .A0(_zyGfifo__gfdL318_31_P0_m2_cbid[1]), .A1(_zyGfifo__gfdL316_32_P0_m2_cbid[1]), .Z(n465));
Q_MX02 U5069 ( .S(n486), .A0(_zyGfifo__gfdL318_31_P0_m2_cbid[0]), .A1(_zyGfifo__gfdL316_32_P0_m2_cbid[0]), .Z(n464));
Q_XNR2 U5070 ( .A0(n463), .A1(_zyGfifoF0_L312_s2_req_0), .Z(n484));
Q_XNR2 U5071 ( .A0(_zyGfifo__gfdL513_33_P0_m2_gfOff), .A1(_zyGfifoF1_L513_req_0), .Z(n462));
Q_OR02 U5072 ( .A0(n460), .A1(n461), .Z(n486));
Q_OR03 U5073 ( .A0(n457), .A1(n458), .A2(n459), .Z(n461));
Q_OR03 U5074 ( .A0(n454), .A1(n455), .A2(n456), .Z(n460));
Q_OR03 U5075 ( .A0(n451), .A1(n452), .A2(n453), .Z(n459));
Q_OR03 U5076 ( .A0(n448), .A1(n449), .A2(n450), .Z(n458));
Q_OR03 U5077 ( .A0(error_cntr[1]), .A1(error_cntr[0]), .A2(n447), .Z(n457));
Q_OR03 U5078 ( .A0(error_cntr[4]), .A1(error_cntr[3]), .A2(error_cntr[2]), .Z(n456));
Q_OR03 U5079 ( .A0(error_cntr[7]), .A1(error_cntr[6]), .A2(error_cntr[5]), .Z(n455));
Q_OR03 U5080 ( .A0(error_cntr[10]), .A1(error_cntr[9]), .A2(error_cntr[8]), .Z(n454));
Q_OR03 U5081 ( .A0(error_cntr[13]), .A1(error_cntr[12]), .A2(error_cntr[11]), .Z(n453));
Q_OR03 U5082 ( .A0(error_cntr[16]), .A1(error_cntr[15]), .A2(error_cntr[14]), .Z(n452));
Q_OR03 U5083 ( .A0(error_cntr[19]), .A1(error_cntr[18]), .A2(error_cntr[17]), .Z(n451));
Q_OR03 U5084 ( .A0(error_cntr[22]), .A1(error_cntr[21]), .A2(error_cntr[20]), .Z(n450));
Q_OR03 U5085 ( .A0(error_cntr[25]), .A1(error_cntr[24]), .A2(error_cntr[23]), .Z(n449));
Q_OR03 U5086 ( .A0(error_cntr[28]), .A1(error_cntr[27]), .A2(error_cntr[26]), .Z(n448));
Q_OR03 U5087 ( .A0(error_cntr[31]), .A1(error_cntr[30]), .A2(error_cntr[29]), .Z(n447));
Q_INV U5088 ( .A(n487), .Z(n446));
Q_AN02 U5089 ( .A0(n444), .A1(config_done), .Z(n445));
Q_FDP0 _zzM2L306_mdxP0_kme_ib_tlast_Dwen1_REG  ( .CK(clk), .D(n445), .Q(_zzM2L306_mdxP0_kme_ib_tlast_Dwen1), .QN( ));
Q_FDP0 _zzM2L306_mdxP0_kme_ib_tvalid_Dwen0_REG  ( .CK(clk), .D(n445), .Q(_zzM2L306_mdxP0_kme_ib_tvalid_Dwen0), .QN( ));
Q_FDP0 \_zyL306_meState0_REG[0] ( .CK(clk), .D(n445), .Q(_zyL306_meState0[0]), .QN(n444));
Q_XNR2 U5093 ( .A0(_zyGfifo__gfdL435_34_P0_m2_gfOff), .A1(_zyGfifoF0_L435_req_0), .Z(n443));
Q_INV U5094 ( .A(n445), .Z(n442));
Q_NOT_TOUCH _zzqnt ( .sig());
ixc_assign _zz_strnp_0 ( clk, my_clk);
ixc_assign _zz_strnp_1 ( kme_apb_psel, _zy_simnet_kme_apb_psel_0_w$);
ixc_assign _zz_strnp_2 ( kme_apb_penable, _zy_simnet_kme_apb_penable_1_w$);
ixc_assign_20 _zz_strnp_3 ( kme_apb_paddr[19:0], 
	_zy_simnet_kme_apb_paddr_2_w$[0:19]);
ixc_assign_32 _zz_strnp_4 ( kme_apb_pwdata[31:0], 
	_zy_simnet_kme_apb_pwdata_3_w$[0:31]);
ixc_assign _zz_strnp_5 ( kme_apb_pwrite, _zy_simnet_kme_apb_pwrite_4_w$);
ixc_assign _zz_strnp_6 ( _zy_simnet_clk_5_w$, clk);
ixc_assign _zz_strnp_7 ( _zy_simnet_rst_n_6_w$, rst_n);
ixc_assign_32 _zz_strnp_8 ( _zy_simnet_kme_apb_prdata_7_w$[0:31], 
	kme_apb_prdata[31:0]);
ixc_assign _zz_strnp_9 ( _zy_simnet_kme_apb_pready_8_w$, kme_apb_pready);
ixc_assign _zz_strnp_10 ( _zy_simnet_kme_apb_pslverr_9_w$, kme_apb_pslverr);
ixc_assign _zz_strnp_11 ( kme_ib_tready, _zy_simnet_kme_ib_tready_11_w$);
ixc_assign _zz_strnp_12 ( kme_ob_tvalid, _zy_simnet_kme_ob_tvalid_12_w$);
ixc_assign _zz_strnp_13 ( kme_ob_tlast, _zy_simnet_kme_ob_tlast_13_w$);
ixc_assign _zz_strnp_14 ( kme_ob_tid[0], _zy_simnet_kme_ob_tid_14_w$);
ixc_assign_8 _zz_strnp_15 ( kme_ob_tstrb[7:0], 
	_zy_simnet_kme_ob_tstrb_15_w$[0:7]);
ixc_assign_8 _zz_strnp_16 ( kme_ob_tuser[7:0], 
	_zy_simnet_kme_ob_tuser_16_w$[0:7]);
ixc_assign_64 _zz_strnp_17 ( kme_ob_tdata[63:0], 
	_zy_simnet_kme_ob_tdata_17_w$[0:63]);
ixc_assign_32 _zz_strnp_18 ( kme_apb_prdata[31:0], 
	_zy_simnet_kme_apb_prdata_18_w$[0:31]);
ixc_assign _zz_strnp_19 ( kme_apb_pready, _zy_simnet_kme_apb_pready_19_w$);
ixc_assign _zz_strnp_20 ( kme_apb_pslverr, _zy_simnet_kme_apb_pslverr_20_w$);
ixc_assign _zz_strnp_21 ( _zy_simnet_clk_22_w$, clk);
ixc_assign _zz_strnp_22 ( _zy_simnet_rst_n_23_w$, rst_n);
ixc_assign _zz_strnp_23 ( _zy_simnet_kme_ib_tvalid_32_w$, kme_ib_tvalid);
ixc_assign _zz_strnp_24 ( _zy_simnet_kme_ib_tlast_33_w$, kme_ib_tlast);
ixc_assign _zz_strnp_25 ( _zy_simnet_kme_ib_tid_34_w$, kme_ib_tid[0]);
ixc_assign_8 _zz_strnp_26 ( _zy_simnet_kme_ib_tstrb_35_w$[0:7], 
	kme_ib_tstrb[7:0]);
ixc_assign_8 _zz_strnp_27 ( _zy_simnet_kme_ib_tuser_36_w$[0:7], 
	kme_ib_tuser[7:0]);
ixc_assign_64 _zz_strnp_28 ( _zy_simnet_kme_ib_tdata_37_w$[0:63], 
	kme_ib_tdata[63:0]);
ixc_assign _zz_strnp_29 ( _zy_simnet_kme_ob_tready_38_w$, kme_ob_tready);
ixc_assign_16 _zz_strnp_30 ( _zy_simnet_kme_apb_paddr_39_w$[0:15], 
	kme_apb_paddr[15:0]);
ixc_assign _zz_strnp_31 ( _zy_simnet_kme_apb_psel_40_w$, kme_apb_psel);
ixc_assign _zz_strnp_32 ( _zy_simnet_kme_apb_penable_41_w$, kme_apb_penable);
ixc_assign _zz_strnp_33 ( _zy_simnet_kme_apb_pwrite_42_w$, kme_apb_pwrite);
ixc_assign_32 _zz_strnp_34 ( _zy_simnet_kme_apb_pwdata_43_w$[0:31], 
	kme_apb_pwdata[31:0]);
ixc_mem_call_0_0 _zzixc_tfport_0_0 ( _zyixc_port_0_0_req, _zyixc_port_0_0_s2h, 
	_zyixc_port_0_0_isf, _zyixc_port_0_0_ack, n59, _zyixc_port_0_0_osf, 
	n60, n61);
ixc_sfifo_port_32_0 _zzSfifoF0_L206_p ( _zySfifoF0_call, 
	_zySfifoF0_iarg[31:0], n62, 
	_zySfifoF0_get_config_data_zyackf_tid[21:0], _zySfifoF0_fen, 
	_zyGfifo_SiData[511:0], _zyGfifo_StId[21:0], 
	_zyGfifo_SoData[511:0], _zyGfifo_SoDataEn, _zyGfifo_SoDataLen[3:0]);
ixc_sfifo_port_72_0 _zzSfifoF1_L206_p ( _zySfifoF1_call, 
	_zySfifoF1_iarg[71:0], n63, 
	_zySfifoF1_get_config_data_zyputf_tid[21:0], _zySfifoF1_fen, 
	_zyGfifo_SiData[511:0], _zyGfifo_StId[21:0], 
	_zyGfifo_SoData[511:0], _zyGfifo_SoDataEn, _zyGfifo_SoDataLen[3:0]);
ixc_sfifo_port_32_0 _zzSfifoF2_L207_p ( _zySfifoF2_call, 
	_zySfifoF2_iarg[31:0], n64, 
	_zySfifoF2_ib_service_data_zyackf_tid[21:0], _zySfifoF2_fen, 
	_zyGfifo_SiData[511:0], _zyGfifo_StId[21:0], 
	_zyGfifo_SoData[511:0], _zyGfifo_SoDataEn, _zyGfifo_SoDataLen[3:0]);
ixc_sfifo_port_136_0 _zzSfifoF3_L207_p ( _zySfifoF3_call, 
	_zySfifoF3_iarg[135:0], n65, 
	_zySfifoF3_ib_service_data_zyputf_tid[21:0], _zySfifoF3_fen, 
	_zyGfifo_SiData[511:0], _zyGfifo_StId[21:0], 
	_zyGfifo_SoData[511:0], _zyGfifo_SoDataEn, _zyGfifo_SoDataLen[3:0]);
ixc_sfifo_port_32_0 _zzSfifoF4_L209_p ( _zySfifoF4_call, 
	_zySfifoF4_iarg[31:0], n66, 
	_zySfifoF4_ob_service_data_zyackf_tid[21:0], _zySfifoF4_fen, 
	_zyGfifo_SiData[511:0], _zyGfifo_StId[21:0], 
	_zyGfifo_SoData[511:0], _zyGfifo_SoDataEn, _zyGfifo_SoDataLen[3:0]);
ixc_sfifo_port_136_0 _zzSfifoF5_L209_p ( _zySfifoF5_call, 
	_zySfifoF5_iarg[135:0], n67, 
	_zySfifoF5_ob_service_data_zyputf_tid[21:0], _zySfifoF5_fen, 
	_zyGfifo_SiData[511:0], _zyGfifo_StId[21:0], 
	_zyGfifo_SoData[511:0], _zyGfifo_SoDataEn, _zyGfifo_SoDataLen[3:0]);
ixc_assign _zz_strnp_35 ( apb_xactor._zyL94_iscX1c0_s, _zyL94_iscX1c0_s);
ixc_assign _zz_strnp_36 ( _zyL94_iscX1c0_f, apb_xactor._zyL94_iscX1c0_f);
ixc_assign_64 _zz_strnp_37 ( apb_xactor._zyL94_iscX1c0_i0[63:0], 
	_zyL94_iscX1c0_i0[63:0]);
ixc_assign_32 _zz_strnp_38 ( _zyL94_iscX1c0_o1[31:0], 
	apb_xactor._zyL94_iscX1c0_o1[31:0]);
ixc_assign _zz_strnp_39 ( _zyL94_iscX1c0_o2, apb_xactor._zyL94_iscX1c0_o2);
ixc_assign _zz_strnp_40 ( apb_xactor._zyL61_iscX2c0_s, _zyL61_iscX2c0_s);
ixc_assign _zz_strnp_41 ( _zyL61_iscX2c0_f, apb_xactor._zyL61_iscX2c0_f);
ixc_assign_64 _zz_strnp_42 ( apb_xactor._zyL61_iscX2c0_i0[63:0], 
	_zyL61_iscX2c0_i0[63:0]);
ixc_assign_32 _zz_strnp_43 ( apb_xactor._zyL61_iscX2c0_i1[31:0], 
	_zyL61_iscX2c0_i1[31:0]);
ixc_assign _zz_strnp_44 ( _zyL61_iscX2c0_o2, apb_xactor._zyL61_iscX2c0_o2);
axis_tbcall_2 _zz_zzictd_finishT_L10_0TbcP_L10 ( _zyictd_finish_mgr, n68, 
	_zyictd_finish_mgr_x$tbc, n69);
Q_OR03 U5149 ( .A0(_zyictd_finish_L454_2), .A1(_zyictd_finish_L320_0), .A2(_zyictd_finish_L338_1), .Z(_zyictd_finish_mgr));
ixc_assign _zz_strnp_45 ( _zyGfifo_dflt_ci[0], _zyGfifo_mod2_dflt_ci);
Q_OR02 U5151 ( .A0(_zyGfifo_dflt_co[0]), .A1(_zyGfifo_mod2_dflt_ci), .Z(_zyGfifo_dflt_ci[1]));
Q_OR03 U5152 ( .A0(_zyGfifo_dflt_co[0]), .A1(_zyGfifo_dflt_co[1]), .A2(_zyGfifo_mod2_dflt_ci), .Z(_zyGfifo_dflt_ci[2]));
Q_OR02 U5153 ( .A0(n147), .A1(_zyGfifo_mod2_dflt_ci), .Z(_zyGfifo_dflt_ci[3]));
Q_OR03 U5154 ( .A0(_zyGfifo_dflt_co[0]), .A1(n109), .A2(_zyGfifo_mod2_dflt_ci), .Z(_zyGfifo_dflt_ci[4]));
Q_OR03 U5155 ( .A0(_zyGfifo_dflt_co[1]), .A1(_zyGfifo_dflt_co[0]), .A2(n121), .Z(n70));
Q_OR02 U5156 ( .A0(n70), .A1(_zyGfifo_mod2_dflt_ci), .Z(_zyGfifo_dflt_ci[5]));
Q_OR03 U5157 ( .A0(n146), .A1(n147), .A2(_zyGfifo_mod2_dflt_ci), .Z(_zyGfifo_dflt_ci[6]));
Q_OR03 U5158 ( .A0(_zyGfifo_dflt_co[0]), .A1(n108), .A2(n109), .Z(n71));
Q_OR02 U5159 ( .A0(n71), .A1(_zyGfifo_mod2_dflt_ci), .Z(_zyGfifo_dflt_ci[7]));
Q_OR03 U5160 ( .A0(_zyGfifo_dflt_co[1]), .A1(_zyGfifo_dflt_co[0]), .A2(n120), .Z(n72));
Q_OR03 U5161 ( .A0(n121), .A1(n72), .A2(_zyGfifo_mod2_dflt_ci), .Z(_zyGfifo_dflt_ci[8]));
Q_OR02 U5162 ( .A0(n150), .A1(_zyGfifo_mod2_dflt_ci), .Z(_zyGfifo_dflt_ci[9]));
Q_OR03 U5163 ( .A0(_zyGfifo_dflt_co[0]), .A1(n107), .A2(n108), .Z(n73));
Q_OR03 U5164 ( .A0(n109), .A1(n73), .A2(_zyGfifo_mod2_dflt_ci), .Z(_zyGfifo_dflt_ci[10]));
Q_OR03 U5165 ( .A0(_zyGfifo_dflt_co[1]), .A1(_zyGfifo_dflt_co[0]), .A2(n119), .Z(n74));
Q_OR03 U5166 ( .A0(n120), .A1(n121), .A2(n74), .Z(n75));
Q_OR02 U5167 ( .A0(n75), .A1(_zyGfifo_mod2_dflt_ci), .Z(_zyGfifo_dflt_ci[11]));
Q_OR03 U5168 ( .A0(n147), .A1(n90), .A2(_zyGfifo_mod2_dflt_ci), .Z(_zyGfifo_dflt_ci[12]));
Q_OR03 U5169 ( .A0(_zyGfifo_dflt_co[0]), .A1(n106), .A2(n107), .Z(n76));
Q_OR03 U5170 ( .A0(n108), .A1(n109), .A2(n76), .Z(n77));
Q_OR02 U5171 ( .A0(n77), .A1(_zyGfifo_mod2_dflt_ci), .Z(_zyGfifo_dflt_ci[13]));
Q_OR03 U5172 ( .A0(_zyGfifo_dflt_co[1]), .A1(_zyGfifo_dflt_co[0]), .A2(n118), .Z(n78));
Q_OR03 U5173 ( .A0(n78), .A1(n97), .A2(_zyGfifo_mod2_dflt_ci), .Z(_zyGfifo_dflt_ci[14]));
Q_OR03 U5174 ( .A0(n146), .A1(n147), .A2(n100), .Z(n79));
Q_OR02 U5175 ( .A0(n79), .A1(_zyGfifo_mod2_dflt_ci), .Z(_zyGfifo_dflt_ci[15]));
Q_OR03 U5176 ( .A0(_zyGfifo_dflt_co[0]), .A1(n105), .A2(n106), .Z(n80));
Q_OR03 U5177 ( .A0(n80), .A1(n112), .A2(_zyGfifo_mod2_dflt_ci), .Z(_zyGfifo_dflt_ci[16]));
Q_OR03 U5178 ( .A0(_zyGfifo_dflt_co[1]), .A1(_zyGfifo_dflt_co[0]), .A2(n117), .Z(n81));
Q_OR03 U5179 ( .A0(n121), .A1(n81), .A2(n124), .Z(n82));
Q_OR02 U5180 ( .A0(n82), .A1(_zyGfifo_mod2_dflt_ci), .Z(_zyGfifo_dflt_ci[17]));
Q_OR03 U5181 ( .A0(n149), .A1(n150), .A2(_zyGfifo_mod2_dflt_ci), .Z(_zyGfifo_dflt_ci[18]));
Q_OR03 U5182 ( .A0(_zyGfifo_dflt_co[0]), .A1(n104), .A2(n105), .Z(n83));
Q_OR03 U5183 ( .A0(n106), .A1(n107), .A2(n108), .Z(n84));
Q_OR03 U5184 ( .A0(n109), .A1(n83), .A2(n84), .Z(n85));
Q_OR02 U5185 ( .A0(n85), .A1(_zyGfifo_mod2_dflt_ci), .Z(_zyGfifo_dflt_ci[19]));
Q_OR03 U5186 ( .A0(_zyGfifo_dflt_co[1]), .A1(_zyGfifo_dflt_co[0]), .A2(n116), .Z(n86));
Q_OR03 U5187 ( .A0(n117), .A1(n118), .A2(n119), .Z(n87));
Q_OR03 U5188 ( .A0(n120), .A1(n121), .A2(n86), .Z(n88));
Q_OR03 U5189 ( .A0(n87), .A1(n88), .A2(_zyGfifo_mod2_dflt_ci), .Z(_zyGfifo_dflt_ci[20]));
Q_OR03 U5190 ( .A0(n141), .A1(n142), .A2(n143), .Z(n89));
Q_OR03 U5191 ( .A0(n144), .A1(n145), .A2(n146), .Z(n90));
Q_OR03 U5192 ( .A0(n147), .A1(n89), .A2(n90), .Z(n91));
Q_OR02 U5193 ( .A0(n91), .A1(_zyGfifo_mod2_dflt_ci), .Z(_zyGfifo_dflt_ci[21]));
Q_OR03 U5194 ( .A0(_zyGfifo_dflt_co[0]), .A1(n103), .A2(n104), .Z(n92));
Q_OR03 U5195 ( .A0(n105), .A1(n106), .A2(n107), .Z(n93));
Q_OR03 U5196 ( .A0(n108), .A1(n109), .A2(n92), .Z(n94));
Q_OR03 U5197 ( .A0(n93), .A1(n94), .A2(_zyGfifo_mod2_dflt_ci), .Z(_zyGfifo_dflt_ci[22]));
Q_OR03 U5198 ( .A0(_zyGfifo_dflt_co[1]), .A1(_zyGfifo_dflt_co[0]), .A2(n115), .Z(n95));
Q_OR03 U5199 ( .A0(n116), .A1(n117), .A2(n118), .Z(n96));
Q_OR03 U5200 ( .A0(n119), .A1(n120), .A2(n121), .Z(n97));
Q_OR03 U5201 ( .A0(n95), .A1(n96), .A2(n97), .Z(n98));
Q_OR02 U5202 ( .A0(n98), .A1(_zyGfifo_mod2_dflt_ci), .Z(_zyGfifo_dflt_ci[23]));
Q_OR03 U5203 ( .A0(n140), .A1(n141), .A2(n142), .Z(n99));
Q_OR03 U5204 ( .A0(n143), .A1(n144), .A2(n145), .Z(n100));
Q_OR03 U5205 ( .A0(n146), .A1(n147), .A2(n99), .Z(n101));
Q_OR03 U5206 ( .A0(n100), .A1(n101), .A2(_zyGfifo_mod2_dflt_ci), .Z(_zyGfifo_dflt_ci[24]));
Q_OR03 U5207 ( .A0(_zyGfifo_dflt_co[24]), .A1(_zyGfifo_dflt_co[23]), .A2(_zyGfifo_dflt_co[22]), .Z(n102));
Q_OR03 U5208 ( .A0(_zyGfifo_dflt_co[21]), .A1(_zyGfifo_dflt_co[20]), .A2(_zyGfifo_dflt_co[19]), .Z(n103));
Q_OR03 U5209 ( .A0(_zyGfifo_dflt_co[18]), .A1(_zyGfifo_dflt_co[17]), .A2(_zyGfifo_dflt_co[16]), .Z(n104));
Q_OR03 U5210 ( .A0(_zyGfifo_dflt_co[15]), .A1(_zyGfifo_dflt_co[14]), .A2(_zyGfifo_dflt_co[13]), .Z(n105));
Q_OR03 U5211 ( .A0(_zyGfifo_dflt_co[12]), .A1(_zyGfifo_dflt_co[11]), .A2(_zyGfifo_dflt_co[10]), .Z(n106));
Q_OR03 U5212 ( .A0(_zyGfifo_dflt_co[9]), .A1(_zyGfifo_dflt_co[8]), .A2(_zyGfifo_dflt_co[7]), .Z(n107));
Q_OR03 U5213 ( .A0(_zyGfifo_dflt_co[6]), .A1(_zyGfifo_dflt_co[5]), .A2(_zyGfifo_dflt_co[4]), .Z(n108));
Q_OR03 U5214 ( .A0(_zyGfifo_dflt_co[3]), .A1(_zyGfifo_dflt_co[2]), .A2(_zyGfifo_dflt_co[1]), .Z(n109));
Q_OR03 U5215 ( .A0(_zyGfifo_dflt_co[0]), .A1(n102), .A2(n103), .Z(n110));
Q_OR03 U5216 ( .A0(n104), .A1(n105), .A2(n106), .Z(n111));
Q_OR03 U5217 ( .A0(n107), .A1(n108), .A2(n109), .Z(n112));
Q_OR03 U5218 ( .A0(n110), .A1(n111), .A2(n112), .Z(n113));
Q_OR02 U5219 ( .A0(n113), .A1(_zyGfifo_mod2_dflt_ci), .Z(_zyGfifo_dflt_ci[25]));
Q_OR03 U5220 ( .A0(_zyGfifo_dflt_co[25]), .A1(_zyGfifo_dflt_co[24]), .A2(_zyGfifo_dflt_co[23]), .Z(n114));
Q_OR03 U5221 ( .A0(_zyGfifo_dflt_co[22]), .A1(_zyGfifo_dflt_co[21]), .A2(_zyGfifo_dflt_co[20]), .Z(n115));
Q_OR03 U5222 ( .A0(_zyGfifo_dflt_co[19]), .A1(_zyGfifo_dflt_co[18]), .A2(_zyGfifo_dflt_co[17]), .Z(n116));
Q_OR03 U5223 ( .A0(_zyGfifo_dflt_co[16]), .A1(_zyGfifo_dflt_co[15]), .A2(_zyGfifo_dflt_co[14]), .Z(n117));
Q_OR03 U5224 ( .A0(_zyGfifo_dflt_co[13]), .A1(_zyGfifo_dflt_co[12]), .A2(_zyGfifo_dflt_co[11]), .Z(n118));
Q_OR03 U5225 ( .A0(_zyGfifo_dflt_co[10]), .A1(_zyGfifo_dflt_co[9]), .A2(_zyGfifo_dflt_co[8]), .Z(n119));
Q_OR03 U5226 ( .A0(_zyGfifo_dflt_co[7]), .A1(_zyGfifo_dflt_co[6]), .A2(_zyGfifo_dflt_co[5]), .Z(n120));
Q_OR03 U5227 ( .A0(_zyGfifo_dflt_co[4]), .A1(_zyGfifo_dflt_co[3]), .A2(_zyGfifo_dflt_co[2]), .Z(n121));
Q_OR03 U5228 ( .A0(_zyGfifo_dflt_co[1]), .A1(_zyGfifo_dflt_co[0]), .A2(n114), .Z(n122));
Q_OR03 U5229 ( .A0(n115), .A1(n116), .A2(n117), .Z(n123));
Q_OR03 U5230 ( .A0(n118), .A1(n119), .A2(n120), .Z(n124));
Q_OR03 U5231 ( .A0(n121), .A1(n122), .A2(n123), .Z(n125));
Q_OR03 U5232 ( .A0(n124), .A1(n125), .A2(_zyGfifo_mod2_dflt_ci), .Z(_zyGfifo_dflt_ci[26]));
ixc_gfifo_port_1_2_0 _zzGfifoF1_L253_s2_p_7 ( _zyGfifo_dflt_co[26], 
	_zyGfifo_dflt_ci[26], _zyGfifoF1_L253_s2_req_7, 
	_zyGfifoF1_L253_s2_cbid_7[19:0], { n126, n127, n128, n129, n130, n131, 
	n132, n133, n134, n135, n136, n137}, n138, _zyGfifo_SGFtsReq, 
	_zyGfifo_SGFcbid[19:0], _zyGfifo_SGFlen[11:0], 
	_zyGfifo_SGFidata[511:0], _zyGfifo_SGFfull, _zyGfifo_SLBreq, 
	_zyGfifo_SLBrd[3:0], _zyGfifo_SLBwr[3:0], _zyGfifo_SLBfull, 
	_zyGfifo_SRtkin);
Q_OR03 U5234 ( .A0(_zyGfifo_dflt_co[26]), .A1(_zyGfifo_dflt_co[25]), .A2(_zyGfifo_dflt_co[24]), .Z(n139));
Q_OR03 U5235 ( .A0(_zyGfifo_dflt_co[23]), .A1(_zyGfifo_dflt_co[22]), .A2(_zyGfifo_dflt_co[21]), .Z(n140));
Q_OR03 U5236 ( .A0(_zyGfifo_dflt_co[20]), .A1(_zyGfifo_dflt_co[19]), .A2(_zyGfifo_dflt_co[18]), .Z(n141));
Q_OR03 U5237 ( .A0(_zyGfifo_dflt_co[17]), .A1(_zyGfifo_dflt_co[16]), .A2(_zyGfifo_dflt_co[15]), .Z(n142));
Q_OR03 U5238 ( .A0(_zyGfifo_dflt_co[14]), .A1(_zyGfifo_dflt_co[13]), .A2(_zyGfifo_dflt_co[12]), .Z(n143));
Q_OR03 U5239 ( .A0(_zyGfifo_dflt_co[11]), .A1(_zyGfifo_dflt_co[10]), .A2(_zyGfifo_dflt_co[9]), .Z(n144));
Q_OR03 U5240 ( .A0(_zyGfifo_dflt_co[8]), .A1(_zyGfifo_dflt_co[7]), .A2(_zyGfifo_dflt_co[6]), .Z(n145));
Q_OR03 U5241 ( .A0(_zyGfifo_dflt_co[5]), .A1(_zyGfifo_dflt_co[4]), .A2(_zyGfifo_dflt_co[3]), .Z(n146));
Q_OR03 U5242 ( .A0(_zyGfifo_dflt_co[2]), .A1(_zyGfifo_dflt_co[1]), .A2(_zyGfifo_dflt_co[0]), .Z(n147));
Q_OR03 U5243 ( .A0(n139), .A1(n140), .A2(n141), .Z(n148));
Q_OR03 U5244 ( .A0(n142), .A1(n143), .A2(n144), .Z(n149));
Q_OR03 U5245 ( .A0(n145), .A1(n146), .A2(n147), .Z(n150));
Q_OR03 U5246 ( .A0(n148), .A1(n149), .A2(n150), .Z(_zyGfifo_mod2_dflt_co));
Q_OR02 U5247 ( .A0(_zyM2L324_pbcCapEn0), .A1(_zyM2L355_pbcCapEn3), .Z(n151));
ixc_mevClk_3_0_0_4_0_3 _zzM2L324_pbcMevClk4 ( _zyM2L324_pbcMevClk4, { clk, 
	_zyL94_iscX1c0_f, _zyL61_iscX2c0_f}, { n151, _zyM2L333_pbcCapEn1, 
	_zyM2L349_pbcCapEn2}, n152, n153, _zyM2L324_pbcReq4, 
	_zyM2L324_pbcBusy4, _zyM2L324_pbcWait4);
Q_OR03 U5249 ( .A0(_zyM2L300_pbcCapEn11), .A1(_zyM2L364_pbcCapEn10), .A2(_zyM2L295_pbcCapEn9), .Z(n154));
Q_OR03 U5250 ( .A0(_zyM2L293_pbcCapEn8), .A1(_zyM2L287_pbcCapEn7), .A2(_zyM2L274_pbcCapEn6), .Z(n155));
Q_OR02 U5251 ( .A0(n154), .A1(n155), .Z(n156));
ixc_mevClk_2_0_0_1 _zzM2L253_pbcMevClk12 ( _zyM2L253_pbcMevClk12, { 
	_zyixc_port_0_0_req, clk}, { _zyM2L253_pbcCapEn5, n156}, n157, n158, 
	_zyM2L253_pbcReq12, _zyM2L253_pbcBusy12, _zyM2L253_pbcWait12);
ixc_capLoopXp _zzM2L10_bcBehEvalP0 ( _zzM2_bcBehEvalClk, n159,, 
	_zzM2_bcBehHalt);
ixc_mdrOn _zzM2L306_mdxP0_OnP ( _zzM2L306_mdxP0_On, _zzM2L306_mdxP0_EnNxt, 
	_zzM2L306_mdxP0_En);
ixc_mdrOn _zzM2L324_mdxP2_OnP ( _zzM2L324_mdxP2_On, _zzM2L324_mdxP2_EnNxt, 
	_zzM2L324_mdxP2_En);
ixc_mdrOn _zzM2L368_mdxP3_OnP ( _zzM2L368_mdxP3_On, _zzM2L368_mdxP3_EnNxt, 
	_zzM2L368_mdxP3_En);
ixc_mdrOn _zzM2L439_mdxP4_OnP ( _zzM2L439_mdxP4_On, _zzM2L439_mdxP4_EnNxt, 
	_zzM2L439_mdxP4_En);
ixc_mdrOn _zzM2L253_mdxP5_OnP ( _zzM2L253_mdxP5_On, _zzM2L253_mdxP5_EnNxt, 
	_zzM2L253_mdxP5_En);
ixc_sampleLT _zzkme_ib_tvalid_M2L36_mdxSpLt7 ( 
	_zzkme_ib_tvalid_M2L36_mdxSvLt7, kme_ib_tvalid);
ixc_sampleLT _zzkme_ib_tlast_M2L37_mdxSpLt8 ( _zzkme_ib_tlast_M2L37_mdxSvLt8, 
	kme_ib_tlast);
ixc_sampleLT_64 _zzkme_ib_tdata_M2L33_mdxSpLt9 ( 
	_zzkme_ib_tdata_M2L33_mdxSvLt9[63:0], kme_ib_tdata[63:0]);
ixc_sampleLT_8 _zzkme_ib_tstrb_M2L34_mdxSpLt10 ( 
	_zzkme_ib_tstrb_M2L34_mdxSvLt10[7:0], kme_ib_tstrb[7:0]);
ixc_sampleLT_8 _zzkme_ib_tuser_M2L35_mdxSpLt11 ( 
	_zzkme_ib_tuser_M2L35_mdxSvLt11[7:0], kme_ib_tuser[7:0]);
apb_xactor apb_xactor ( .psel( _zy_simnet_kme_apb_psel_0_w$), .penable( 
	_zy_simnet_kme_apb_penable_1_w$), .paddr( 
	_zy_simnet_kme_apb_paddr_2_w$[0:19]), .pwdata( 
	_zy_simnet_kme_apb_pwdata_3_w$[0:31]), .pwrite( 
	_zy_simnet_kme_apb_pwrite_4_w$), .clk( _zy_simnet_clk_5_w$), 
	.reset_n( _zy_simnet_rst_n_6_w$), .prdata( 
	_zy_simnet_kme_apb_prdata_7_w$[0:31]), .pready( 
	_zy_simnet_kme_apb_pready_8_w$), .pslverr( 
	_zy_simnet_kme_apb_pslverr_9_w$));
cr_kme kme_dut ( .kme_interrupt( _zy_simnet_dio_10), .kme_ib_tready( 
	_zy_simnet_kme_ib_tready_11_w$), .kme_cceip0_ob_tvalid( 
	_zy_simnet_kme_ob_tvalid_12_w$), .kme_cceip0_ob_tlast( 
	_zy_simnet_kme_ob_tlast_13_w$), .kme_cceip0_ob_tid( 
	_zy_simnet_kme_ob_tid_14_w$), .kme_cceip0_ob_tstrb( 
	_zy_simnet_kme_ob_tstrb_15_w$[0:7]), .kme_cceip0_ob_tuser( 
	_zy_simnet_kme_ob_tuser_16_w$[0:7]), .kme_cceip0_ob_tdata( 
	_zy_simnet_kme_ob_tdata_17_w$[0:63]), .apb_prdata( 
	_zy_simnet_kme_apb_prdata_18_w$[0:31]), .apb_pready( 
	_zy_simnet_kme_apb_pready_19_w$), .apb_pslverr( 
	_zy_simnet_kme_apb_pslverr_20_w$), .kme_idle( _zy_simnet_dio_21), 
	.clk( _zy_simnet_clk_22_w$), .rst_n( _zy_simnet_rst_n_23_w$), 
	.scan_en( _zy_simnet_cio_24), .scan_mode( _zy_simnet_cio_25), 
	.scan_rst_n( _zy_simnet_cio_26), .ovstb( _zy_simnet_cio_27), .lvm( 
	_zy_simnet_cio_28), .mlvm( _zy_simnet_cio_29), .disable_debug_cmd( 
	_zy_simnet_cio_30), .disable_unencrypted_keys( _zy_simnet_cio_31), 
	.kme_ib_tvalid( _zy_simnet_kme_ib_tvalid_32_w$), .kme_ib_tlast( 
	_zy_simnet_kme_ib_tlast_33_w$), .kme_ib_tid( 
	_zy_simnet_kme_ib_tid_34_w$), .kme_ib_tstrb( 
	_zy_simnet_kme_ib_tstrb_35_w$[0:7]), .kme_ib_tuser( 
	_zy_simnet_kme_ib_tuser_36_w$[0:7]), .kme_ib_tdata( 
	_zy_simnet_kme_ib_tdata_37_w$[0:63]), .kme_cceip0_ob_tready( 
	_zy_simnet_kme_ob_tready_38_w$), .apb_paddr( 
	_zy_simnet_kme_apb_paddr_39_w$[0:15]), .apb_psel( 
	_zy_simnet_kme_apb_psel_40_w$), .apb_penable( 
	_zy_simnet_kme_apb_penable_41_w$), .apb_pwrite( 
	_zy_simnet_kme_apb_pwrite_42_w$), .apb_pwdata( 
	_zy_simnet_kme_apb_pwdata_43_w$[0:31]));
ixc_assign _zzmdx1 ( _zzmdxOne, n160);
ixc_gfifo_port_1 _zzGfifoF0_L435_p_0 ( _zyGfifo_dflt_co[0], 
	_zyGfifo_dflt_ci[0], _zyGfifoF0_L435_req_0, 
	_zyGfifo__gfdL435_34_P0_m2_cbid[19:0], { n161, n162, n163, n164, n165, 
	n166, n167, n168, n169, n170, n171, n172}, n173, _zyGfifo_SGFtsReq, 
	_zyGfifo_SGFcbid[19:0], _zyGfifo_SGFlen[11:0], 
	_zyGfifo_SGFidata[511:0], _zyGfifo_SGFfull, _zyGfifo_SLBreq, 
	_zyGfifo_SLBrd[3:0], _zyGfifo_SLBwr[3:0], _zyGfifo_SLBfull, 
	_zyGfifo_SRtkin);
ixc_gfifo_port_1 _zzGfifoF1_L513_p_0 ( _zyGfifo_dflt_co[1], 
	_zyGfifo_dflt_ci[1], _zyGfifoF1_L513_req_0, 
	_zyGfifo__gfdL513_33_P0_m2_cbid[19:0], { n174, n175, n176, n177, n178, 
	n179, n180, n181, n182, n183, n184, n185}, n186, _zyGfifo_SGFtsReq, 
	_zyGfifo_SGFcbid[19:0], _zyGfifo_SGFlen[11:0], 
	_zyGfifo_SGFidata[511:0], _zyGfifo_SGFfull, _zyGfifo_SLBreq, 
	_zyGfifo_SLBrd[3:0], _zyGfifo_SLBwr[3:0], _zyGfifo_SLBfull, 
	_zyGfifo_SRtkin);
ixc_gfifo_port_280_2_0 _zzGfifoF0_L312_s2_p_0 ( _zyGfifo_dflt_co[2], 
	_zyGfifo_dflt_ci[2], _zyGfifoF0_L312_s2_req_0, 
	_zyGfifoF0_L312_s2_cbid_0[19:0], { n187, n188, n189, n190, n191, n192, 
	n193, n194, n195, n196, n197, n198}, 
	_zyGfifoF0_L312_s2_data_0[279:0], _zyGfifo_SGFtsReq, 
	_zyGfifo_SGFcbid[19:0], _zyGfifo_SGFlen[11:0], 
	_zyGfifo_SGFidata[511:0], _zyGfifo_SGFfull, _zyGfifo_SLBreq, 
	_zyGfifo_SLBrd[3:0], _zyGfifo_SLBwr[3:0], _zyGfifo_SLBfull, 
	_zyGfifo_SRtkin);
ixc_gfifo_port_96_3 _zzGfifoF0_L324_s3_p_1 ( _zyGfifo_dflt_co[3], 
	_zyGfifo_dflt_ci[3], _zyGfifoF0_L324_s3_req_1, 
	_zyGfifoF0_L324_s3_cbid_1[19:0], _zyGfifoF0_L324_s3_len_1[11:0], 
	_zyGfifoF0_L324_s3_data_1[95:0], _zyGfifo_SGFtsReq, 
	_zyGfifo_SGFcbid[19:0], _zyGfifo_SGFlen[11:0], 
	_zyGfifo_SGFidata[511:0], _zyGfifo_SGFfull, _zyGfifo_SLBreq, 
	_zyGfifo_SLBrd[3:0], _zyGfifo_SLBwr[3:0], _zyGfifo_SLBfull, 
	_zyGfifo_SRtkin);
ixc_gfifo_port_32_2 _zzGfifoF1_L324_s2_p_2 ( _zyGfifo_dflt_co[4], 
	_zyGfifo_dflt_ci[4], _zyGfifoF1_L324_s2_req_2, 
	_zyGfifoF1_L324_s2_cbid_2[19:0], { n199, n200, n201, n202, n203, n204, 
	n205, n206, n207, n208, n209, n210}, 
	_zyGfifoF1_L324_s2_data_2[31:0], _zyGfifo_SGFtsReq, 
	_zyGfifo_SGFcbid[19:0], _zyGfifo_SGFlen[11:0], 
	_zyGfifo_SGFidata[511:0], _zyGfifo_SGFfull, _zyGfifo_SLBreq, 
	_zyGfifo_SLBrd[3:0], _zyGfifo_SLBwr[3:0], _zyGfifo_SLBfull, 
	_zyGfifo_SRtkin);
ixc_gfifo_port_72_3 _zzGfifoF2_L324_s2_p_3 ( _zyGfifo_dflt_co[5], 
	_zyGfifo_dflt_ci[5], _zyGfifoF2_L324_s2_req_3, 
	_zyGfifoF2_L324_s2_cbid_3[19:0], _zyGfifoF2_L324_s2_len_3[11:0], 
	_zyGfifoF2_L324_s2_data_3[71:0], _zyGfifo_SGFtsReq, 
	_zyGfifo_SGFcbid[19:0], _zyGfifo_SGFlen[11:0], 
	_zyGfifo_SGFidata[511:0], _zyGfifo_SGFfull, _zyGfifo_SLBreq, 
	_zyGfifo_SLBrd[3:0], _zyGfifo_SLBwr[3:0], _zyGfifo_SLBfull, 
	_zyGfifo_SRtkin);
ixc_gfifo_port_32_0_0 _zzGfifoF11_L207_p_0 ( _zyGfifo_dflt_co[6], 
	_zyGfifo_dflt_ci[6], _zyGfifoF11_L207_req_0, 
	_zyGfifo_ib_service_data_2_zyprefetch_m2_cbid[19:0], { n211, n212, 
	n213, n214, n215, n216, n217, n218, n219, n220, n221, n222}, 
	_zyGfifoF11_L207_data_0[31:0], _zyGfifo_SGFtsReq, 
	_zyGfifo_SGFcbid[19:0], _zyGfifo_SGFlen[11:0], 
	_zyGfifo_SGFidata[511:0], _zyGfifo_SGFfull, _zyGfifo_SLBreq, 
	_zyGfifo_SLBrd[3:0], _zyGfifo_SLBwr[3:0], _zyGfifo_SLBfull, 
	_zyGfifo_SRtkin);
ixc_gfifo_port_1_2_0 _zzGfifoF0_L368_s2_p_4 ( _zyGfifo_dflt_co[7], 
	_zyGfifo_dflt_ci[7], _zyGfifoF0_L368_s2_req_4, 
	_zyGfifoF0_L368_s2_cbid_4[19:0], { n223, n224, n225, n226, n227, n228, 
	n229, n230, n231, n232, n233, n234}, n235, _zyGfifo_SGFtsReq, 
	_zyGfifo_SGFcbid[19:0], _zyGfifo_SGFlen[11:0], 
	_zyGfifo_SGFidata[511:0], _zyGfifo_SGFfull, _zyGfifo_SLBreq, 
	_zyGfifo_SLBrd[3:0], _zyGfifo_SLBwr[3:0], _zyGfifo_SLBfull, 
	_zyGfifo_SRtkin);
ixc_gfifo_port_32_0_0 _zzGfifoF14_L373_p_0 ( _zyGfifo_dflt_co[8], 
	_zyGfifo_dflt_ci[8], _zyGfifoF14_L373_req_0, 
	_zyGfifo__gfdL373_22_P0_m2_cbid[19:0], { n236, n237, n238, n239, n240, 
	n241, n242, n243, n244, n245, n246, n247}, 
	_zyGfifoF14_L373_data_0[31:0], _zyGfifo_SGFtsReq, 
	_zyGfifo_SGFcbid[19:0], _zyGfifo_SGFlen[11:0], 
	_zyGfifo_SGFidata[511:0], _zyGfifo_SGFfull, _zyGfifo_SLBreq, 
	_zyGfifo_SLBrd[3:0], _zyGfifo_SLBwr[3:0], _zyGfifo_SLBfull, 
	_zyGfifo_SRtkin);
ixc_gfifo_port_136_0_0 _zzGfifoF15_L375_p_0 ( _zyGfifo_dflt_co[9], 
	_zyGfifo_dflt_ci[9], _zyGfifoF15_L375_req_0, 
	_zyGfifo__gfdL375_21_P0_m2_cbid[19:0], { n248, n249, n250, n251, n252, 
	n253, n254, n255, n256, n257, n258, n259}, 
	_zyGfifoF15_L375_data_0[135:0], _zyGfifo_SGFtsReq, 
	_zyGfifo_SGFcbid[19:0], _zyGfifo_SGFlen[11:0], 
	_zyGfifo_SGFidata[511:0], _zyGfifo_SGFfull, _zyGfifo_SLBreq, 
	_zyGfifo_SLBrd[3:0], _zyGfifo_SLBwr[3:0], _zyGfifo_SLBfull, 
	_zyGfifo_SRtkin);
ixc_gfifo_port_1_0_0 _zzGfifoF16_L381_p_0 ( _zyGfifo_dflt_co[10], 
	_zyGfifo_dflt_ci[10], _zyGfifoF16_L381_req_0, 
	_zyGfifo__gfdL381_20_P0_m2_cbid[19:0], { n260, n261, n262, n263, n264, 
	n265, n266, n267, n268, n269, n270, n271}, n272, _zyGfifo_SGFtsReq, 
	_zyGfifo_SGFcbid[19:0], _zyGfifo_SGFlen[11:0], 
	_zyGfifo_SGFidata[511:0], _zyGfifo_SGFfull, _zyGfifo_SLBreq, 
	_zyGfifo_SLBrd[3:0], _zyGfifo_SLBwr[3:0], _zyGfifo_SLBfull, 
	_zyGfifo_SRtkin);
ixc_gfifo_port_64_0_0 _zzGfifoF17_L390_p_0 ( _zyGfifo_dflt_co[11], 
	_zyGfifo_dflt_ci[11], _zyGfifoF17_L390_req_0, 
	_zyGfifo__gfdL390_19_P0_m2_cbid[19:0], { n273, n274, n275, n276, n277, 
	n278, n279, n280, n281, n282, n283, n284}, 
	_zyGfifoF17_L390_data_0[63:0], _zyGfifo_SGFtsReq, 
	_zyGfifo_SGFcbid[19:0], _zyGfifo_SGFlen[11:0], 
	_zyGfifo_SGFidata[511:0], _zyGfifo_SGFfull, _zyGfifo_SLBreq, 
	_zyGfifo_SLBrd[3:0], _zyGfifo_SLBwr[3:0], _zyGfifo_SLBfull, 
	_zyGfifo_SRtkin);
ixc_gfifo_port_32_0_0 _zzGfifoF18_L530_p_0 ( _zyGfifo_dflt_co[12], 
	_zyGfifo_dflt_ci[12], _zyGfifoF18_L530_req_0, 
	_zyGfifo__gfdL530_18_P0_m2_cbid[19:0], { n285, n286, n287, n288, n289, 
	n290, n291, n292, n293, n294, n295, n296}, 
	_zyGfifoF18_L530_data_0[31:0], _zyGfifo_SGFtsReq, 
	_zyGfifo_SGFcbid[19:0], _zyGfifo_SGFlen[11:0], 
	_zyGfifo_SGFidata[511:0], _zyGfifo_SGFfull, _zyGfifo_SLBreq, 
	_zyGfifo_SLBrd[3:0], _zyGfifo_SLBwr[3:0], _zyGfifo_SLBfull, 
	_zyGfifo_SRtkin);
ixc_gfifo_port_8_0_0 _zzGfifoF19_L412_p_0 ( _zyGfifo_dflt_co[13], 
	_zyGfifo_dflt_ci[13], _zyGfifoF19_L412_req_0, 
	_zyGfifo__gfdL412_17_P0_m2_cbid[19:0], { n297, n298, n299, n300, n301, 
	n302, n303, n304, n305, n306, n307, n308}, 
	_zyGfifoF19_L412_data_0[7:0], _zyGfifo_SGFtsReq, 
	_zyGfifo_SGFcbid[19:0], _zyGfifo_SGFlen[11:0], 
	_zyGfifo_SGFidata[511:0], _zyGfifo_SGFfull, _zyGfifo_SLBreq, 
	_zyGfifo_SLBrd[3:0], _zyGfifo_SLBwr[3:0], _zyGfifo_SLBfull, 
	_zyGfifo_SRtkin);
ixc_gfifo_port_32_0_0 _zzGfifoF20_L209_p_0 ( _zyGfifo_dflt_co[14], 
	_zyGfifo_dflt_ci[14], _zyGfifoF20_L209_req_0, 
	_zyGfifo_ob_service_data_2_zyprefetch_m2_cbid[19:0], { n309, n310, 
	n311, n312, n313, n314, n315, n316, n317, n318, n319, n320}, 
	_zyGfifoF20_L209_data_0[31:0], _zyGfifo_SGFtsReq, 
	_zyGfifo_SGFcbid[19:0], _zyGfifo_SGFlen[11:0], 
	_zyGfifo_SGFidata[511:0], _zyGfifo_SGFfull, _zyGfifo_SLBreq, 
	_zyGfifo_SLBrd[3:0], _zyGfifo_SLBwr[3:0], _zyGfifo_SLBfull, 
	_zyGfifo_SRtkin);
ixc_gfifo_port_1_2_0 _zzGfifoF0_L439_s2_p_5 ( _zyGfifo_dflt_co[15], 
	_zyGfifo_dflt_ci[15], _zyGfifoF0_L439_s2_req_5, 
	_zyGfifoF0_L439_s2_cbid_5[19:0], { n321, n322, n323, n324, n325, n326, 
	n327, n328, n329, n330, n331, n332}, n333, _zyGfifo_SGFtsReq, 
	_zyGfifo_SGFcbid[19:0], _zyGfifo_SGFlen[11:0], 
	_zyGfifo_SGFidata[511:0], _zyGfifo_SGFfull, _zyGfifo_SLBreq, 
	_zyGfifo_SLBrd[3:0], _zyGfifo_SLBwr[3:0], _zyGfifo_SLBfull, 
	_zyGfifo_SRtkin);
ixc_gfifo_port_32_0_0 _zzGfifoF23_L444_p_0 ( _zyGfifo_dflt_co[16], 
	_zyGfifo_dflt_ci[16], _zyGfifoF23_L444_req_0, 
	_zyGfifo__gfdL444_14_P0_m2_cbid[19:0], { n334, n335, n336, n337, n338, 
	n339, n340, n341, n342, n343, n344, n345}, 
	_zyGfifoF23_L444_data_0[31:0], _zyGfifo_SGFtsReq, 
	_zyGfifo_SGFcbid[19:0], _zyGfifo_SGFlen[11:0], 
	_zyGfifo_SGFidata[511:0], _zyGfifo_SGFfull, _zyGfifo_SLBreq, 
	_zyGfifo_SLBrd[3:0], _zyGfifo_SLBwr[3:0], _zyGfifo_SLBfull, 
	_zyGfifo_SRtkin);
ixc_gfifo_port_136_0_0 _zzGfifoF24_L446_p_0 ( _zyGfifo_dflt_co[17], 
	_zyGfifo_dflt_ci[17], _zyGfifoF24_L446_req_0, 
	_zyGfifo__gfdL446_13_P0_m2_cbid[19:0], { n346, n347, n348, n349, n350, 
	n351, n352, n353, n354, n355, n356, n357}, 
	_zyGfifoF24_L446_data_0[135:0], _zyGfifo_SGFtsReq, 
	_zyGfifo_SGFcbid[19:0], _zyGfifo_SGFlen[11:0], 
	_zyGfifo_SGFidata[511:0], _zyGfifo_SGFfull, _zyGfifo_SLBreq, 
	_zyGfifo_SLBrd[3:0], _zyGfifo_SLBwr[3:0], _zyGfifo_SLBfull, 
	_zyGfifo_SRtkin);
ixc_gfifo_port_64 _zzGfifoF25_L460_p_0 ( _zyGfifo_dflt_co[18], 
	_zyGfifo_dflt_ci[18], _zyGfifoF25_L460_req_0, 
	_zyGfifo__gfdL460_12_P0_m2_cbid[19:0], { n358, n359, n360, n361, n362, 
	n363, n364, n365, n366, n367, n368, n369}, 
	_zyGfifoF25_L460_data_0[63:0], _zyGfifo_SGFtsReq, 
	_zyGfifo_SGFcbid[19:0], _zyGfifo_SGFlen[11:0], 
	_zyGfifo_SGFidata[511:0], _zyGfifo_SGFfull, _zyGfifo_SLBreq, 
	_zyGfifo_SLBrd[3:0], _zyGfifo_SLBwr[3:0], _zyGfifo_SLBfull, 
	_zyGfifo_SRtkin);
ixc_gfifo_port_32_0_0 _zzGfifoF26_L530_p_0 ( _zyGfifo_dflt_co[19], 
	_zyGfifo_dflt_ci[19], _zyGfifoF26_L530_req_0, 
	_zyGfifo__gfdL530_11_P0_m2_cbid[19:0], { n370, n371, n372, n373, n374, 
	n375, n376, n377, n378, n379, n380, n381}, 
	_zyGfifoF26_L530_data_0[31:0], _zyGfifo_SGFtsReq, 
	_zyGfifo_SGFcbid[19:0], _zyGfifo_SGFlen[11:0], 
	_zyGfifo_SGFidata[511:0], _zyGfifo_SGFfull, _zyGfifo_SLBreq, 
	_zyGfifo_SLBrd[3:0], _zyGfifo_SLBwr[3:0], _zyGfifo_SLBfull, 
	_zyGfifo_SRtkin);
ixc_gfifo_port_8_0_0 _zzGfifoF27_L480_p_0 ( _zyGfifo_dflt_co[20], 
	_zyGfifo_dflt_ci[20], _zyGfifoF27_L480_req_0, 
	_zyGfifo__gfdL480_10_P0_m2_cbid[19:0], { n382, n383, n384, n385, n386, 
	n387, n388, n389, n390, n391, n392, n393}, 
	_zyGfifoF27_L480_data_0[7:0], _zyGfifo_SGFtsReq, 
	_zyGfifo_SGFcbid[19:0], _zyGfifo_SGFlen[11:0], 
	_zyGfifo_SGFidata[511:0], _zyGfifo_SGFfull, _zyGfifo_SLBreq, 
	_zyGfifo_SLBrd[3:0], _zyGfifo_SLBwr[3:0], _zyGfifo_SLBfull, 
	_zyGfifo_SRtkin);
ixc_gfifo_port_128 _zzGfifoF28_L482_p_0 ( _zyGfifo_dflt_co[21], 
	_zyGfifo_dflt_ci[21], _zyGfifoF28_L482_req_0, 
	_zyGfifo__gfdL482_9_P0_m2_cbid[19:0], { n394, n395, n396, n397, n398, 
	n399, n400, n401, n402, n403, n404, n405}, 
	_zyGfifoF28_L482_data_0[127:0], _zyGfifo_SGFtsReq, 
	_zyGfifo_SGFcbid[19:0], _zyGfifo_SGFlen[11:0], 
	_zyGfifo_SGFidata[511:0], _zyGfifo_SGFfull, _zyGfifo_SLBreq, 
	_zyGfifo_SLBrd[3:0], _zyGfifo_SLBwr[3:0], _zyGfifo_SLBfull, 
	_zyGfifo_SRtkin);
ixc_gfifo_port_16 _zzGfifoF29_L487_p_0 ( _zyGfifo_dflt_co[22], 
	_zyGfifo_dflt_ci[22], _zyGfifoF29_L487_req_0, 
	_zyGfifo__gfdL487_8_P0_m2_cbid[19:0], { n406, n407, n408, n409, n410, 
	n411, n412, n413, n414, n415, n416, n417}, 
	_zyGfifoF29_L487_data_0[15:0], _zyGfifo_SGFtsReq, 
	_zyGfifo_SGFcbid[19:0], _zyGfifo_SGFlen[11:0], 
	_zyGfifo_SGFidata[511:0], _zyGfifo_SGFfull, _zyGfifo_SLBreq, 
	_zyGfifo_SLBrd[3:0], _zyGfifo_SLBwr[3:0], _zyGfifo_SLBfull, 
	_zyGfifo_SRtkin);
ixc_gfifo_port_16 _zzGfifoF30_L491_p_0 ( _zyGfifo_dflt_co[23], 
	_zyGfifo_dflt_ci[23], _zyGfifoF30_L491_req_0, 
	_zyGfifo__gfdL491_7_P0_m2_cbid[19:0], { n418, n419, n420, n421, n422, 
	n423, n424, n425, n426, n427, n428, n429}, 
	_zyGfifoF30_L491_data_0[15:0], _zyGfifo_SGFtsReq, 
	_zyGfifo_SGFcbid[19:0], _zyGfifo_SGFlen[11:0], 
	_zyGfifo_SGFidata[511:0], _zyGfifo_SGFfull, _zyGfifo_SLBreq, 
	_zyGfifo_SLBrd[3:0], _zyGfifo_SLBwr[3:0], _zyGfifo_SLBfull, 
	_zyGfifo_SRtkin);
ixc_gfifo_port_16 _zzGfifoF31_L496_p_0 ( _zyGfifo_dflt_co[24], 
	_zyGfifo_dflt_ci[24], _zyGfifoF31_L496_req_0, 
	_zyGfifo__gfdL496_6_P0_m2_cbid[19:0], { n430, n431, n432, n433, n434, 
	n435, n436, n437, n438, n439, n440, n441}, 
	_zyGfifoF31_L496_data_0[15:0], _zyGfifo_SGFtsReq, 
	_zyGfifo_SGFcbid[19:0], _zyGfifo_SGFlen[11:0], 
	_zyGfifo_SGFidata[511:0], _zyGfifo_SGFfull, _zyGfifo_SLBreq, 
	_zyGfifo_SLBrd[3:0], _zyGfifo_SLBwr[3:0], _zyGfifo_SLBfull, 
	_zyGfifo_SRtkin);
ixc_gfifo_port_560_3 _zzGfifoF0_L253_s4_p_6 ( _zyGfifo_dflt_co[25], 
	_zyGfifo_dflt_ci[25], _zyGfifoF0_L253_s4_req_6, 
	_zyGfifoF0_L253_s4_cbid_6[19:0], _zyGfifoF0_L253_s4_len_6[11:0], 
	_zyGfifoF0_L253_s4_data_6[559:0], _zyGfifo_SGFtsReq, 
	_zyGfifo_SGFcbid[19:0], _zyGfifo_SGFlen[11:0], 
	_zyGfifo_SGFidata[511:0], _zyGfifo_SGFfull, _zyGfifo_SLBreq, 
	_zyGfifo_SLBrd[3:0], _zyGfifo_SLBwr[3:0], _zyGfifo_SLBfull, 
	_zyGfifo_SRtkin);
ixc_sampleLT_32 _zzerror_cntr_M2L19_mdxSpLt6 ( 
	_zzerror_cntr_M2L19_mdxSvLt6[31:0], error_cntr[31:0]);
Q_INV U5294 ( .A(n5275), .Z(n54));
Q_FDP4EP ready_ib_REG  ( .CK(clk), .CE(n445), .R(n1750), .D(n5382), .Q(ready_ib));
Q_INV U5296 ( .A(ready_ib), .Z(n1492));
Q_FDP4EP saw_mega_REG  ( .CK(clk), .CE(n1715), .R(n1750), .D(n1712), .Q(saw_mega));
Q_FDP4EP saw_guid_tlv_REG  ( .CK(clk), .CE(n1715), .R(n1750), .D(n1713), .Q(saw_guid_tlv));
Q_FDP4EP have_guid_tlv_REG  ( .CK(clk), .CE(n1715), .R(n1750), .D(n1714), .Q(have_guid_tlv));
Q_FDP4EP \mega_tlv_word_count_REG[31] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1716), .Q(mega_tlv_word_count[31]));
Q_FDP4EP \mega_tlv_word_count_REG[30] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1717), .Q(mega_tlv_word_count[30]));
Q_FDP4EP \mega_tlv_word_count_REG[29] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1718), .Q(mega_tlv_word_count[29]));
Q_FDP4EP \mega_tlv_word_count_REG[28] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1719), .Q(mega_tlv_word_count[28]));
Q_FDP4EP \mega_tlv_word_count_REG[27] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1720), .Q(mega_tlv_word_count[27]));
Q_FDP4EP \mega_tlv_word_count_REG[26] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1721), .Q(mega_tlv_word_count[26]));
Q_FDP4EP \mega_tlv_word_count_REG[25] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1722), .Q(mega_tlv_word_count[25]));
Q_FDP4EP \mega_tlv_word_count_REG[24] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1723), .Q(mega_tlv_word_count[24]));
Q_FDP4EP \mega_tlv_word_count_REG[23] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1724), .Q(mega_tlv_word_count[23]));
Q_FDP4EP \mega_tlv_word_count_REG[22] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1725), .Q(mega_tlv_word_count[22]));
Q_FDP4EP \mega_tlv_word_count_REG[21] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1726), .Q(mega_tlv_word_count[21]));
Q_FDP4EP \mega_tlv_word_count_REG[20] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1727), .Q(mega_tlv_word_count[20]));
Q_FDP4EP \mega_tlv_word_count_REG[19] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1728), .Q(mega_tlv_word_count[19]));
Q_FDP4EP \mega_tlv_word_count_REG[18] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1729), .Q(mega_tlv_word_count[18]));
Q_FDP4EP \mega_tlv_word_count_REG[17] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1730), .Q(mega_tlv_word_count[17]));
Q_FDP4EP \mega_tlv_word_count_REG[16] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1731), .Q(mega_tlv_word_count[16]));
Q_FDP4EP \mega_tlv_word_count_REG[15] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1732), .Q(mega_tlv_word_count[15]));
Q_FDP4EP \mega_tlv_word_count_REG[14] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1733), .Q(mega_tlv_word_count[14]));
Q_FDP4EP \mega_tlv_word_count_REG[13] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1734), .Q(mega_tlv_word_count[13]));
Q_FDP4EP \mega_tlv_word_count_REG[12] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1735), .Q(mega_tlv_word_count[12]));
Q_FDP4EP \mega_tlv_word_count_REG[11] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1736), .Q(mega_tlv_word_count[11]));
Q_FDP4EP \mega_tlv_word_count_REG[10] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1737), .Q(mega_tlv_word_count[10]));
Q_FDP4EP \mega_tlv_word_count_REG[9] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1738), .Q(mega_tlv_word_count[9]));
Q_FDP4EP \mega_tlv_word_count_REG[8] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1739), .Q(mega_tlv_word_count[8]));
Q_FDP4EP \mega_tlv_word_count_REG[7] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1740), .Q(mega_tlv_word_count[7]));
Q_FDP4EP \mega_tlv_word_count_REG[6] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1741), .Q(mega_tlv_word_count[6]));
Q_FDP4EP \mega_tlv_word_count_REG[5] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1742), .Q(mega_tlv_word_count[5]));
Q_FDP4EP \mega_tlv_word_count_REG[4] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1743), .Q(mega_tlv_word_count[4]));
Q_FDP4EP \mega_tlv_word_count_REG[3] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1744), .Q(mega_tlv_word_count[3]));
Q_FDP4EP \mega_tlv_word_count_REG[2] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1745), .Q(mega_tlv_word_count[2]));
Q_FDP4EP \mega_tlv_word_count_REG[1] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1746), .Q(mega_tlv_word_count[1]));
Q_FDP4EP \mega_tlv_word_count_REG[0] ( .CK(clk), .CE(n1749), .R(n1750), .D(n1748), .Q(mega_tlv_word_count[0]));
Q_INV U5332 ( .A(mega_tlv_word_count[0]), .Z(n1747));
Q_FDP4EP _zzM2L306_mdxP0_En_REG  ( .CK(clk), .CE(n445), .R(n1750), .D(_zzM2L306_mdxP0_EnNxt), .Q(_zzM2L306_mdxP0_En));
Q_FDP4EP _zzM2L306_mdxP0_kme_ib_tvalid_wr0_REG  ( .CK(clk), .CE(n445), .R(n1750), .D(n1750), .Q(_zzM2L306_mdxP0_kme_ib_tvalid_wr0));
Q_FDP4EP _zzM2L306_mdxP0_kme_ib_tlast_wr1_REG  ( .CK(clk), .CE(n445), .R(n1750), .D(n1750), .Q(_zzM2L306_mdxP0_kme_ib_tlast_wr1));
Q_FDP4EP _zyGfifoF0_L435_req_0_REG  ( .CK(clk), .CE(_zyL306_meState0[0]), .R(n1750), .D(n443), .Q(_zyGfifoF0_L435_req_0));
Q_FDP4EP ready_ob_REG  ( .CK(clk), .CE(n487), .R(n1750), .D(n5382), .Q(ready_ob));
Q_INV U5338 ( .A(ready_ob), .Z(n3315));
Q_FDP4EP saw_cqe_REG  ( .CK(clk), .CE(n3569), .R(n1750), .D(n3568), .Q(saw_cqe));
Q_FDP4EP saw_stats_REG  ( .CK(clk), .CE(n3571), .R(n1750), .D(n3570), .Q(saw_stats));
Q_FDP4EP \watchdog_timer_REG[31] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3572), .Q(watchdog_timer[31]));
Q_FDP4EP \watchdog_timer_REG[30] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3573), .Q(watchdog_timer[30]));
Q_FDP4EP \watchdog_timer_REG[29] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3574), .Q(watchdog_timer[29]));
Q_FDP4EP \watchdog_timer_REG[28] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3575), .Q(watchdog_timer[28]));
Q_FDP4EP \watchdog_timer_REG[27] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3576), .Q(watchdog_timer[27]));
Q_FDP4EP \watchdog_timer_REG[26] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3577), .Q(watchdog_timer[26]));
Q_FDP4EP \watchdog_timer_REG[25] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3578), .Q(watchdog_timer[25]));
Q_FDP4EP \watchdog_timer_REG[24] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3579), .Q(watchdog_timer[24]));
Q_FDP4EP \watchdog_timer_REG[23] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3580), .Q(watchdog_timer[23]));
Q_FDP4EP \watchdog_timer_REG[22] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3581), .Q(watchdog_timer[22]));
Q_FDP4EP \watchdog_timer_REG[21] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3582), .Q(watchdog_timer[21]));
Q_FDP4EP \watchdog_timer_REG[20] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3583), .Q(watchdog_timer[20]));
Q_FDP4EP \watchdog_timer_REG[19] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3584), .Q(watchdog_timer[19]));
Q_FDP4EP \watchdog_timer_REG[18] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3585), .Q(watchdog_timer[18]));
Q_FDP4EP \watchdog_timer_REG[17] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3586), .Q(watchdog_timer[17]));
Q_FDP4EP \watchdog_timer_REG[16] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3587), .Q(watchdog_timer[16]));
Q_FDP4EP \watchdog_timer_REG[15] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3588), .Q(watchdog_timer[15]));
Q_FDP4EP \watchdog_timer_REG[14] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3589), .Q(watchdog_timer[14]));
Q_FDP4EP \watchdog_timer_REG[13] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3590), .Q(watchdog_timer[13]));
Q_FDP4EP \watchdog_timer_REG[12] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3591), .Q(watchdog_timer[12]));
Q_FDP4EP \watchdog_timer_REG[11] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3592), .Q(watchdog_timer[11]));
Q_FDP4EP \watchdog_timer_REG[10] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3593), .Q(watchdog_timer[10]));
Q_FDP4EP \watchdog_timer_REG[9] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3594), .Q(watchdog_timer[9]));
Q_FDP4EP \watchdog_timer_REG[8] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3595), .Q(watchdog_timer[8]));
Q_FDP4EP \watchdog_timer_REG[7] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3596), .Q(watchdog_timer[7]));
Q_FDP4EP \watchdog_timer_REG[6] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3597), .Q(watchdog_timer[6]));
Q_FDP4EP \watchdog_timer_REG[5] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3598), .Q(watchdog_timer[5]));
Q_FDP4EP \watchdog_timer_REG[4] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3599), .Q(watchdog_timer[4]));
Q_FDP4EP \watchdog_timer_REG[3] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3600), .Q(watchdog_timer[3]));
Q_FDP4EP \watchdog_timer_REG[2] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3601), .Q(watchdog_timer[2]));
Q_FDP4EP \watchdog_timer_REG[1] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3602), .Q(watchdog_timer[1]));
Q_FDP4EP \watchdog_timer_REG[0] ( .CK(clk), .CE(n3604), .R(n1750), .D(n3603), .Q(watchdog_timer[0]));
Q_INV U5373 ( .A(watchdog_timer[0]), .Z(n2294));
Q_FDP4EP _zyictd_finish_L320_0_REG  ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(n5382), .Q(_zyictd_finish_L320_0));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[279] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[279]), .Q(_zyGfifoF0_L312_s2_data_0[279]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[278] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[278]), .Q(_zyGfifoF0_L312_s2_data_0[278]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[277] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[277]), .Q(_zyGfifoF0_L312_s2_data_0[277]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[276] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[276]), .Q(_zyGfifoF0_L312_s2_data_0[276]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[275] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[275]), .Q(_zyGfifoF0_L312_s2_data_0[275]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[274] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[274]), .Q(_zyGfifoF0_L312_s2_data_0[274]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[273] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[273]), .Q(_zyGfifoF0_L312_s2_data_0[273]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[272] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[272]), .Q(_zyGfifoF0_L312_s2_data_0[272]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[271] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[271]), .Q(_zyGfifoF0_L312_s2_data_0[271]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[270] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[270]), .Q(_zyGfifoF0_L312_s2_data_0[270]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[269] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[269]), .Q(_zyGfifoF0_L312_s2_data_0[269]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[268] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[268]), .Q(_zyGfifoF0_L312_s2_data_0[268]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[267] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[267]), .Q(_zyGfifoF0_L312_s2_data_0[267]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[266] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[266]), .Q(_zyGfifoF0_L312_s2_data_0[266]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[265] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[265]), .Q(_zyGfifoF0_L312_s2_data_0[265]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[264] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[264]), .Q(_zyGfifoF0_L312_s2_data_0[264]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[263] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[263]), .Q(_zyGfifoF0_L312_s2_data_0[263]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[262] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[262]), .Q(_zyGfifoF0_L312_s2_data_0[262]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[261] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[261]), .Q(_zyGfifoF0_L312_s2_data_0[261]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[260] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[260]), .Q(_zyGfifoF0_L312_s2_data_0[260]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[259] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[259]), .Q(_zyGfifoF0_L312_s2_data_0[259]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[258] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[258]), .Q(_zyGfifoF0_L312_s2_data_0[258]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[257] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[257]), .Q(_zyGfifoF0_L312_s2_data_0[257]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[256] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[256]), .Q(_zyGfifoF0_L312_s2_data_0[256]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[255] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[255]), .Q(_zyGfifoF0_L312_s2_data_0[255]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[254] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[254]), .Q(_zyGfifoF0_L312_s2_data_0[254]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[253] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[253]), .Q(_zyGfifoF0_L312_s2_data_0[253]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[252] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[252]), .Q(_zyGfifoF0_L312_s2_data_0[252]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[251] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[251]), .Q(_zyGfifoF0_L312_s2_data_0[251]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[250] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[250]), .Q(_zyGfifoF0_L312_s2_data_0[250]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[249] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[249]), .Q(_zyGfifoF0_L312_s2_data_0[249]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[248] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[248]), .Q(_zyGfifoF0_L312_s2_data_0[248]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[247] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[247]), .Q(_zyGfifoF0_L312_s2_data_0[247]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[246] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[246]), .Q(_zyGfifoF0_L312_s2_data_0[246]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[245] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[245]), .Q(_zyGfifoF0_L312_s2_data_0[245]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[244] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[244]), .Q(_zyGfifoF0_L312_s2_data_0[244]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[243] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[243]), .Q(_zyGfifoF0_L312_s2_data_0[243]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[242] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[242]), .Q(_zyGfifoF0_L312_s2_data_0[242]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[241] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[241]), .Q(_zyGfifoF0_L312_s2_data_0[241]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[240] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[240]), .Q(_zyGfifoF0_L312_s2_data_0[240]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[239] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[239]), .Q(_zyGfifoF0_L312_s2_data_0[239]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[238] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[238]), .Q(_zyGfifoF0_L312_s2_data_0[238]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[237] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[237]), .Q(_zyGfifoF0_L312_s2_data_0[237]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[236] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[236]), .Q(_zyGfifoF0_L312_s2_data_0[236]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[235] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[235]), .Q(_zyGfifoF0_L312_s2_data_0[235]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[234] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[234]), .Q(_zyGfifoF0_L312_s2_data_0[234]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[233] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[233]), .Q(_zyGfifoF0_L312_s2_data_0[233]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[232] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[232]), .Q(_zyGfifoF0_L312_s2_data_0[232]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[231] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[231]), .Q(_zyGfifoF0_L312_s2_data_0[231]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[230] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[230]), .Q(_zyGfifoF0_L312_s2_data_0[230]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[229] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[229]), .Q(_zyGfifoF0_L312_s2_data_0[229]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[228] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[228]), .Q(_zyGfifoF0_L312_s2_data_0[228]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[227] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[227]), .Q(_zyGfifoF0_L312_s2_data_0[227]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[226] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[226]), .Q(_zyGfifoF0_L312_s2_data_0[226]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[225] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[225]), .Q(_zyGfifoF0_L312_s2_data_0[225]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[224] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[224]), .Q(_zyGfifoF0_L312_s2_data_0[224]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[223] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[223]), .Q(_zyGfifoF0_L312_s2_data_0[223]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[222] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[222]), .Q(_zyGfifoF0_L312_s2_data_0[222]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[221] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[221]), .Q(_zyGfifoF0_L312_s2_data_0[221]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[220] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[220]), .Q(_zyGfifoF0_L312_s2_data_0[220]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[219] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[219]), .Q(_zyGfifoF0_L312_s2_data_0[219]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[218] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[218]), .Q(_zyGfifoF0_L312_s2_data_0[218]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[217] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[217]), .Q(_zyGfifoF0_L312_s2_data_0[217]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[216] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[216]), .Q(_zyGfifoF0_L312_s2_data_0[216]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[215] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[215]), .Q(_zyGfifoF0_L312_s2_data_0[215]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[214] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[214]), .Q(_zyGfifoF0_L312_s2_data_0[214]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[213] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[213]), .Q(_zyGfifoF0_L312_s2_data_0[213]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[212] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[212]), .Q(_zyGfifoF0_L312_s2_data_0[212]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[211] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[211]), .Q(_zyGfifoF0_L312_s2_data_0[211]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[210] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[210]), .Q(_zyGfifoF0_L312_s2_data_0[210]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[209] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[209]), .Q(_zyGfifoF0_L312_s2_data_0[209]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[208] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[208]), .Q(_zyGfifoF0_L312_s2_data_0[208]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[207] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[207]), .Q(_zyGfifoF0_L312_s2_data_0[207]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[206] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[206]), .Q(_zyGfifoF0_L312_s2_data_0[206]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[205] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[205]), .Q(_zyGfifoF0_L312_s2_data_0[205]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[204] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[204]), .Q(_zyGfifoF0_L312_s2_data_0[204]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[203] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[203]), .Q(_zyGfifoF0_L312_s2_data_0[203]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[202] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[202]), .Q(_zyGfifoF0_L312_s2_data_0[202]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[201] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[201]), .Q(_zyGfifoF0_L312_s2_data_0[201]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[200] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[200]), .Q(_zyGfifoF0_L312_s2_data_0[200]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[199] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[199]), .Q(_zyGfifoF0_L312_s2_data_0[199]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[198] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[198]), .Q(_zyGfifoF0_L312_s2_data_0[198]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[197] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[197]), .Q(_zyGfifoF0_L312_s2_data_0[197]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[196] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[196]), .Q(_zyGfifoF0_L312_s2_data_0[196]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[195] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[195]), .Q(_zyGfifoF0_L312_s2_data_0[195]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[194] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[194]), .Q(_zyGfifoF0_L312_s2_data_0[194]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[193] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[193]), .Q(_zyGfifoF0_L312_s2_data_0[193]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[192] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[192]), .Q(_zyGfifoF0_L312_s2_data_0[192]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[191] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[191]), .Q(_zyGfifoF0_L312_s2_data_0[191]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[190] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[190]), .Q(_zyGfifoF0_L312_s2_data_0[190]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[189] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[189]), .Q(_zyGfifoF0_L312_s2_data_0[189]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[188] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[188]), .Q(_zyGfifoF0_L312_s2_data_0[188]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[187] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[187]), .Q(_zyGfifoF0_L312_s2_data_0[187]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[186] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[186]), .Q(_zyGfifoF0_L312_s2_data_0[186]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[185] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[185]), .Q(_zyGfifoF0_L312_s2_data_0[185]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[184] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[184]), .Q(_zyGfifoF0_L312_s2_data_0[184]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[183] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[183]), .Q(_zyGfifoF0_L312_s2_data_0[183]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[182] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[182]), .Q(_zyGfifoF0_L312_s2_data_0[182]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[181] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[181]), .Q(_zyGfifoF0_L312_s2_data_0[181]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[180] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[180]), .Q(_zyGfifoF0_L312_s2_data_0[180]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[179] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[179]), .Q(_zyGfifoF0_L312_s2_data_0[179]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[178] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[178]), .Q(_zyGfifoF0_L312_s2_data_0[178]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[177] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[177]), .Q(_zyGfifoF0_L312_s2_data_0[177]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[176] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[176]), .Q(_zyGfifoF0_L312_s2_data_0[176]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[175] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[175]), .Q(_zyGfifoF0_L312_s2_data_0[175]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[174] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[174]), .Q(_zyGfifoF0_L312_s2_data_0[174]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[173] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[173]), .Q(_zyGfifoF0_L312_s2_data_0[173]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[172] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[172]), .Q(_zyGfifoF0_L312_s2_data_0[172]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[171] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[171]), .Q(_zyGfifoF0_L312_s2_data_0[171]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[170] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[170]), .Q(_zyGfifoF0_L312_s2_data_0[170]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[169] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[169]), .Q(_zyGfifoF0_L312_s2_data_0[169]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[168] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[168]), .Q(_zyGfifoF0_L312_s2_data_0[168]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[167] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[167]), .Q(_zyGfifoF0_L312_s2_data_0[167]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[166] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[166]), .Q(_zyGfifoF0_L312_s2_data_0[166]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[165] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[165]), .Q(_zyGfifoF0_L312_s2_data_0[165]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[164] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[164]), .Q(_zyGfifoF0_L312_s2_data_0[164]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[163] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[163]), .Q(_zyGfifoF0_L312_s2_data_0[163]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[162] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[162]), .Q(_zyGfifoF0_L312_s2_data_0[162]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[161] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[161]), .Q(_zyGfifoF0_L312_s2_data_0[161]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[160] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[160]), .Q(_zyGfifoF0_L312_s2_data_0[160]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[159] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[159]), .Q(_zyGfifoF0_L312_s2_data_0[159]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[158] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[158]), .Q(_zyGfifoF0_L312_s2_data_0[158]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[157] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[157]), .Q(_zyGfifoF0_L312_s2_data_0[157]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[156] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[156]), .Q(_zyGfifoF0_L312_s2_data_0[156]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[155] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[155]), .Q(_zyGfifoF0_L312_s2_data_0[155]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[154] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[154]), .Q(_zyGfifoF0_L312_s2_data_0[154]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[153] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[153]), .Q(_zyGfifoF0_L312_s2_data_0[153]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[152] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[152]), .Q(_zyGfifoF0_L312_s2_data_0[152]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[151] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[151]), .Q(_zyGfifoF0_L312_s2_data_0[151]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[150] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[150]), .Q(_zyGfifoF0_L312_s2_data_0[150]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[149] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[149]), .Q(_zyGfifoF0_L312_s2_data_0[149]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[148] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[148]), .Q(_zyGfifoF0_L312_s2_data_0[148]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[147] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[147]), .Q(_zyGfifoF0_L312_s2_data_0[147]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[146] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[146]), .Q(_zyGfifoF0_L312_s2_data_0[146]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[145] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[145]), .Q(_zyGfifoF0_L312_s2_data_0[145]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[144] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[144]), .Q(_zyGfifoF0_L312_s2_data_0[144]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[143] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[143]), .Q(_zyGfifoF0_L312_s2_data_0[143]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[142] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[142]), .Q(_zyGfifoF0_L312_s2_data_0[142]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[141] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[141]), .Q(_zyGfifoF0_L312_s2_data_0[141]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[140] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[140]), .Q(_zyGfifoF0_L312_s2_data_0[140]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[139] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[139]), .Q(_zyGfifoF0_L312_s2_data_0[139]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[138] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[138]), .Q(_zyGfifoF0_L312_s2_data_0[138]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[137] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[137]), .Q(_zyGfifoF0_L312_s2_data_0[137]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[136] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[136]), .Q(_zyGfifoF0_L312_s2_data_0[136]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[135] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[135]), .Q(_zyGfifoF0_L312_s2_data_0[135]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[134] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[134]), .Q(_zyGfifoF0_L312_s2_data_0[134]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[133] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[133]), .Q(_zyGfifoF0_L312_s2_data_0[133]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[132] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[132]), .Q(_zyGfifoF0_L312_s2_data_0[132]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[131] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[131]), .Q(_zyGfifoF0_L312_s2_data_0[131]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[130] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[130]), .Q(_zyGfifoF0_L312_s2_data_0[130]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[129] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[129]), .Q(_zyGfifoF0_L312_s2_data_0[129]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[128] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[128]), .Q(_zyGfifoF0_L312_s2_data_0[128]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[127] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[127]), .Q(_zyGfifoF0_L312_s2_data_0[127]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[126] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[126]), .Q(_zyGfifoF0_L312_s2_data_0[126]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[125] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[125]), .Q(_zyGfifoF0_L312_s2_data_0[125]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[124] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[124]), .Q(_zyGfifoF0_L312_s2_data_0[124]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[123] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[123]), .Q(_zyGfifoF0_L312_s2_data_0[123]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[122] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[122]), .Q(_zyGfifoF0_L312_s2_data_0[122]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[121] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[121]), .Q(_zyGfifoF0_L312_s2_data_0[121]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[120] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[120]), .Q(_zyGfifoF0_L312_s2_data_0[120]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[119] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[119]), .Q(_zyGfifoF0_L312_s2_data_0[119]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[118] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[118]), .Q(_zyGfifoF0_L312_s2_data_0[118]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[117] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[117]), .Q(_zyGfifoF0_L312_s2_data_0[117]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[116] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[116]), .Q(_zyGfifoF0_L312_s2_data_0[116]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[115] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[115]), .Q(_zyGfifoF0_L312_s2_data_0[115]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[114] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[114]), .Q(_zyGfifoF0_L312_s2_data_0[114]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[113] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[113]), .Q(_zyGfifoF0_L312_s2_data_0[113]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[112] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[112]), .Q(_zyGfifoF0_L312_s2_data_0[112]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[111] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[111]), .Q(_zyGfifoF0_L312_s2_data_0[111]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[110] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[110]), .Q(_zyGfifoF0_L312_s2_data_0[110]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[109] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[109]), .Q(_zyGfifoF0_L312_s2_data_0[109]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[108] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[108]), .Q(_zyGfifoF0_L312_s2_data_0[108]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[107] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[107]), .Q(_zyGfifoF0_L312_s2_data_0[107]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[106] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[106]), .Q(_zyGfifoF0_L312_s2_data_0[106]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[105] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[105]), .Q(_zyGfifoF0_L312_s2_data_0[105]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[104] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[104]), .Q(_zyGfifoF0_L312_s2_data_0[104]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[103] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[103]), .Q(_zyGfifoF0_L312_s2_data_0[103]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[102] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[102]), .Q(_zyGfifoF0_L312_s2_data_0[102]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[101] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[101]), .Q(_zyGfifoF0_L312_s2_data_0[101]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[100] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[100]), .Q(_zyGfifoF0_L312_s2_data_0[100]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[99] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[99]), .Q(_zyGfifoF0_L312_s2_data_0[99]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[98] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[98]), .Q(_zyGfifoF0_L312_s2_data_0[98]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[97] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[97]), .Q(_zyGfifoF0_L312_s2_data_0[97]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[96] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[96]), .Q(_zyGfifoF0_L312_s2_data_0[96]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[95] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[95]), .Q(_zyGfifoF0_L312_s2_data_0[95]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[94] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[94]), .Q(_zyGfifoF0_L312_s2_data_0[94]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[93] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[93]), .Q(_zyGfifoF0_L312_s2_data_0[93]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[92] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[92]), .Q(_zyGfifoF0_L312_s2_data_0[92]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[91] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[91]), .Q(_zyGfifoF0_L312_s2_data_0[91]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[90] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[90]), .Q(_zyGfifoF0_L312_s2_data_0[90]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[89] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[89]), .Q(_zyGfifoF0_L312_s2_data_0[89]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[88] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[88]), .Q(_zyGfifoF0_L312_s2_data_0[88]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[87] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[87]), .Q(_zyGfifoF0_L312_s2_data_0[87]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[86] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[86]), .Q(_zyGfifoF0_L312_s2_data_0[86]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[85] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[85]), .Q(_zyGfifoF0_L312_s2_data_0[85]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[84] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[84]), .Q(_zyGfifoF0_L312_s2_data_0[84]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[83] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[83]), .Q(_zyGfifoF0_L312_s2_data_0[83]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[82] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[82]), .Q(_zyGfifoF0_L312_s2_data_0[82]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[81] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[81]), .Q(_zyGfifoF0_L312_s2_data_0[81]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[80] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[80]), .Q(_zyGfifoF0_L312_s2_data_0[80]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[79] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[79]), .Q(_zyGfifoF0_L312_s2_data_0[79]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[78] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[78]), .Q(_zyGfifoF0_L312_s2_data_0[78]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[77] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[77]), .Q(_zyGfifoF0_L312_s2_data_0[77]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[76] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[76]), .Q(_zyGfifoF0_L312_s2_data_0[76]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[75] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[75]), .Q(_zyGfifoF0_L312_s2_data_0[75]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[74] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[74]), .Q(_zyGfifoF0_L312_s2_data_0[74]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[73] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[73]), .Q(_zyGfifoF0_L312_s2_data_0[73]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[72] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[72]), .Q(_zyGfifoF0_L312_s2_data_0[72]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[71] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[71]), .Q(_zyGfifoF0_L312_s2_data_0[71]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[70] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[70]), .Q(_zyGfifoF0_L312_s2_data_0[70]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[69] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[69]), .Q(_zyGfifoF0_L312_s2_data_0[69]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[68] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[68]), .Q(_zyGfifoF0_L312_s2_data_0[68]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[67] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[67]), .Q(_zyGfifoF0_L312_s2_data_0[67]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[66] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[66]), .Q(_zyGfifoF0_L312_s2_data_0[66]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[65] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[65]), .Q(_zyGfifoF0_L312_s2_data_0[65]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[64] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[64]), .Q(_zyGfifoF0_L312_s2_data_0[64]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[63] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[63]), .Q(_zyGfifoF0_L312_s2_data_0[63]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[62] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[62]), .Q(_zyGfifoF0_L312_s2_data_0[62]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[61] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[61]), .Q(_zyGfifoF0_L312_s2_data_0[61]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[60] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[60]), .Q(_zyGfifoF0_L312_s2_data_0[60]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[59] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[59]), .Q(_zyGfifoF0_L312_s2_data_0[59]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[58] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[58]), .Q(_zyGfifoF0_L312_s2_data_0[58]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[57] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[57]), .Q(_zyGfifoF0_L312_s2_data_0[57]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[56] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[56]), .Q(_zyGfifoF0_L312_s2_data_0[56]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[55] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[55]), .Q(_zyGfifoF0_L312_s2_data_0[55]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[54] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[54]), .Q(_zyGfifoF0_L312_s2_data_0[54]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[53] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[53]), .Q(_zyGfifoF0_L312_s2_data_0[53]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[52] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[52]), .Q(_zyGfifoF0_L312_s2_data_0[52]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[51] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[51]), .Q(_zyGfifoF0_L312_s2_data_0[51]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[50] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[50]), .Q(_zyGfifoF0_L312_s2_data_0[50]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[49] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[49]), .Q(_zyGfifoF0_L312_s2_data_0[49]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[48] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[48]), .Q(_zyGfifoF0_L312_s2_data_0[48]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[47] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[47]), .Q(_zyGfifoF0_L312_s2_data_0[47]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[46] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[46]), .Q(_zyGfifoF0_L312_s2_data_0[46]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[45] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[45]), .Q(_zyGfifoF0_L312_s2_data_0[45]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[44] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[44]), .Q(_zyGfifoF0_L312_s2_data_0[44]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[43] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[43]), .Q(_zyGfifoF0_L312_s2_data_0[43]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[42] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[42]), .Q(_zyGfifoF0_L312_s2_data_0[42]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[41] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[41]), .Q(_zyGfifoF0_L312_s2_data_0[41]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[40] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[40]), .Q(_zyGfifoF0_L312_s2_data_0[40]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[39] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[39]), .Q(_zyGfifoF0_L312_s2_data_0[39]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[38] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[38]), .Q(_zyGfifoF0_L312_s2_data_0[38]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[37] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[37]), .Q(_zyGfifoF0_L312_s2_data_0[37]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[36] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[36]), .Q(_zyGfifoF0_L312_s2_data_0[36]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[35] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[35]), .Q(_zyGfifoF0_L312_s2_data_0[35]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[34] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[34]), .Q(_zyGfifoF0_L312_s2_data_0[34]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[33] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[33]), .Q(_zyGfifoF0_L312_s2_data_0[33]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[32] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[32]), .Q(_zyGfifoF0_L312_s2_data_0[32]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[31] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[31]), .Q(_zyGfifoF0_L312_s2_data_0[31]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[30] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[30]), .Q(_zyGfifoF0_L312_s2_data_0[30]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[29] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[29]), .Q(_zyGfifoF0_L312_s2_data_0[29]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[28] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[28]), .Q(_zyGfifoF0_L312_s2_data_0[28]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[27] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[27]), .Q(_zyGfifoF0_L312_s2_data_0[27]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[26] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[26]), .Q(_zyGfifoF0_L312_s2_data_0[26]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[25] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[25]), .Q(_zyGfifoF0_L312_s2_data_0[25]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[24] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[24]), .Q(_zyGfifoF0_L312_s2_data_0[24]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[23] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[23]), .Q(_zyGfifoF0_L312_s2_data_0[23]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[22] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[22]), .Q(_zyGfifoF0_L312_s2_data_0[22]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[21] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[21]), .Q(_zyGfifoF0_L312_s2_data_0[21]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[20] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[20]), .Q(_zyGfifoF0_L312_s2_data_0[20]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[19] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[19]), .Q(_zyGfifoF0_L312_s2_data_0[19]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[18] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[18]), .Q(_zyGfifoF0_L312_s2_data_0[18]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[17] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[17]), .Q(_zyGfifoF0_L312_s2_data_0[17]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[16] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[16]), .Q(_zyGfifoF0_L312_s2_data_0[16]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[15] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[15]), .Q(_zyGfifoF0_L312_s2_data_0[15]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[14] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[14]), .Q(_zyGfifoF0_L312_s2_data_0[14]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[13] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[13]), .Q(_zyGfifoF0_L312_s2_data_0[13]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[12] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[12]), .Q(_zyGfifoF0_L312_s2_data_0[12]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[11] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[11]), .Q(_zyGfifoF0_L312_s2_data_0[11]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[10] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[10]), .Q(_zyGfifoF0_L312_s2_data_0[10]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[9] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[9]), .Q(_zyGfifoF0_L312_s2_data_0[9]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[8] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[8]), .Q(_zyGfifoF0_L312_s2_data_0[8]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[7] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[7]), .Q(_zyGfifoF0_L312_s2_data_0[7]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[6] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[6]), .Q(_zyGfifoF0_L312_s2_data_0[6]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[5] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[5]), .Q(_zyGfifoF0_L312_s2_data_0[5]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[4] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[4]), .Q(_zyGfifoF0_L312_s2_data_0[4]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[3] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[3]), .Q(_zyGfifoF0_L312_s2_data_0[3]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[2] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[2]), .Q(_zyGfifoF0_L312_s2_data_0[2]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[1] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[1]), .Q(_zyGfifoF0_L312_s2_data_0[1]));
Q_FDP4EP \_zyGfifoF0_L312_s2_data_0_REG[0] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(testname[0]), .Q(_zyGfifoF0_L312_s2_data_0[0]));
Q_FDP4EP _zyGfifoF1_L513_req_0_REG  ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(n462), .Q(_zyGfifoF1_L513_req_0));
Q_FDP4EP _zyGfifoF0_L312_s2_req_0_REG  ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(n484), .Q(_zyGfifoF0_L312_s2_req_0));
Q_FDP4EP \_zyGfifoF0_L312_s2_cbid_0_REG[19] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(n483), .Q(_zyGfifoF0_L312_s2_cbid_0[19]));
Q_FDP4EP \_zyGfifoF0_L312_s2_cbid_0_REG[18] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(n482), .Q(_zyGfifoF0_L312_s2_cbid_0[18]));
Q_FDP4EP \_zyGfifoF0_L312_s2_cbid_0_REG[17] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(n481), .Q(_zyGfifoF0_L312_s2_cbid_0[17]));
Q_FDP4EP \_zyGfifoF0_L312_s2_cbid_0_REG[16] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(n480), .Q(_zyGfifoF0_L312_s2_cbid_0[16]));
Q_FDP4EP \_zyGfifoF0_L312_s2_cbid_0_REG[15] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(n479), .Q(_zyGfifoF0_L312_s2_cbid_0[15]));
Q_FDP4EP \_zyGfifoF0_L312_s2_cbid_0_REG[14] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(n478), .Q(_zyGfifoF0_L312_s2_cbid_0[14]));
Q_FDP4EP \_zyGfifoF0_L312_s2_cbid_0_REG[13] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(n477), .Q(_zyGfifoF0_L312_s2_cbid_0[13]));
Q_FDP4EP \_zyGfifoF0_L312_s2_cbid_0_REG[12] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(n476), .Q(_zyGfifoF0_L312_s2_cbid_0[12]));
Q_FDP4EP \_zyGfifoF0_L312_s2_cbid_0_REG[11] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(n475), .Q(_zyGfifoF0_L312_s2_cbid_0[11]));
Q_FDP4EP \_zyGfifoF0_L312_s2_cbid_0_REG[10] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(n474), .Q(_zyGfifoF0_L312_s2_cbid_0[10]));
Q_FDP4EP \_zyGfifoF0_L312_s2_cbid_0_REG[9] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(n473), .Q(_zyGfifoF0_L312_s2_cbid_0[9]));
Q_FDP4EP \_zyGfifoF0_L312_s2_cbid_0_REG[8] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(n472), .Q(_zyGfifoF0_L312_s2_cbid_0[8]));
Q_FDP4EP \_zyGfifoF0_L312_s2_cbid_0_REG[7] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(n471), .Q(_zyGfifoF0_L312_s2_cbid_0[7]));
Q_FDP4EP \_zyGfifoF0_L312_s2_cbid_0_REG[6] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(n470), .Q(_zyGfifoF0_L312_s2_cbid_0[6]));
Q_FDP4EP \_zyGfifoF0_L312_s2_cbid_0_REG[5] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(n469), .Q(_zyGfifoF0_L312_s2_cbid_0[5]));
Q_FDP4EP \_zyGfifoF0_L312_s2_cbid_0_REG[4] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(n468), .Q(_zyGfifoF0_L312_s2_cbid_0[4]));
Q_FDP4EP \_zyGfifoF0_L312_s2_cbid_0_REG[3] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(n467), .Q(_zyGfifoF0_L312_s2_cbid_0[3]));
Q_FDP4EP \_zyGfifoF0_L312_s2_cbid_0_REG[2] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(n466), .Q(_zyGfifoF0_L312_s2_cbid_0[2]));
Q_FDP4EP \_zyGfifoF0_L312_s2_cbid_0_REG[1] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(n465), .Q(_zyGfifoF0_L312_s2_cbid_0[1]));
Q_FDP4EP \_zyGfifoF0_L312_s2_cbid_0_REG[0] ( .CK(clk), .CE(_zyL312_meState2[0]), .R(n1750), .D(n464), .Q(_zyGfifoF0_L312_s2_cbid_0[0]));
Q_FDP4EP _zyL94_iscX1c0_s_REG  ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(_zyL94_iscX1c0_n), .Q(_zyL94_iscX1c0_s));
Q_FDP4EP _zyL61_iscX2c0_s_REG  ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(_zyL61_iscX2c0_n), .Q(_zyL61_iscX2c0_s));
Q_FDP4EP _zyictd_finish_L338_1_REG  ( .CK(_zyM2L324_pbcMevClk4), .CE(n1137), .R(n1750), .D(n5382), .Q(_zyictd_finish_L338_1));
Q_FDP4EP _zzM2L324_mdxP2_En_REG  ( .CK(_zyM2L324_pbcMevClk4), .CE(n1126), .R(n1750), .D(_zzM2L324_mdxP2_EnNxt), .Q(_zzM2L324_mdxP2_En));
Q_INV U5681 ( .A(n1008), .Z(n53));
Q_FDP4EP \returned_data_REG[31] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[31]), .Q(returned_data[31]));
Q_FDP4EP \returned_data_REG[30] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[30]), .Q(returned_data[30]));
Q_FDP4EP \returned_data_REG[29] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[29]), .Q(returned_data[29]));
Q_FDP4EP \returned_data_REG[28] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[28]), .Q(returned_data[28]));
Q_FDP4EP \returned_data_REG[27] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[27]), .Q(returned_data[27]));
Q_FDP4EP \returned_data_REG[26] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[26]), .Q(returned_data[26]));
Q_FDP4EP \returned_data_REG[25] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[25]), .Q(returned_data[25]));
Q_FDP4EP \returned_data_REG[24] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[24]), .Q(returned_data[24]));
Q_FDP4EP \returned_data_REG[23] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[23]), .Q(returned_data[23]));
Q_FDP4EP \returned_data_REG[22] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[22]), .Q(returned_data[22]));
Q_FDP4EP \returned_data_REG[21] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[21]), .Q(returned_data[21]));
Q_FDP4EP \returned_data_REG[20] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[20]), .Q(returned_data[20]));
Q_FDP4EP \returned_data_REG[19] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[19]), .Q(returned_data[19]));
Q_FDP4EP \returned_data_REG[18] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[18]), .Q(returned_data[18]));
Q_FDP4EP \returned_data_REG[17] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[17]), .Q(returned_data[17]));
Q_FDP4EP \returned_data_REG[16] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[16]), .Q(returned_data[16]));
Q_FDP4EP \returned_data_REG[15] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[15]), .Q(returned_data[15]));
Q_FDP4EP \returned_data_REG[14] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[14]), .Q(returned_data[14]));
Q_FDP4EP \returned_data_REG[13] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[13]), .Q(returned_data[13]));
Q_FDP4EP \returned_data_REG[12] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[12]), .Q(returned_data[12]));
Q_FDP4EP \returned_data_REG[11] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[11]), .Q(returned_data[11]));
Q_FDP4EP \returned_data_REG[10] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[10]), .Q(returned_data[10]));
Q_FDP4EP \returned_data_REG[9] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[9]), .Q(returned_data[9]));
Q_FDP4EP \returned_data_REG[8] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[8]), .Q(returned_data[8]));
Q_FDP4EP \returned_data_REG[7] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[7]), .Q(returned_data[7]));
Q_FDP4EP \returned_data_REG[6] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[6]), .Q(returned_data[6]));
Q_FDP4EP \returned_data_REG[5] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[5]), .Q(returned_data[5]));
Q_FDP4EP \returned_data_REG[4] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[4]), .Q(returned_data[4]));
Q_FDP4EP \returned_data_REG[3] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[3]), .Q(returned_data[3]));
Q_FDP4EP \returned_data_REG[2] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[2]), .Q(returned_data[2]));
Q_FDP4EP \returned_data_REG[1] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[1]), .Q(returned_data[1]));
Q_FDP4EP \returned_data_REG[0] ( .CK(_zyM2L324_pbcMevClk4), .CE(n53), .R(n1750), .D(_zyL94_iscX1c0_o1[0]), .Q(returned_data[0]));
Q_INV U5714 ( .A(_zygsfis_get_config_data_req[4]), .Z(n52));
Q_FDP4EP \_zygsfis_get_config_data_req_REG[4] ( .CK(_zyM2L324_pbcMevClk4), .CE(n5884), .R(n1750), .D(n52), .Q(_zygsfis_get_config_data_req[4]));
Q_FDP4EP \_zygsfis_get_config_data_req_REG[3] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1134), .R(n1750), .D(n578), .Q(_zygsfis_get_config_data_req[3]));
Q_FDP4EP \_zygsfis_get_config_data_req_REG[2] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1134), .R(n1750), .D(n576), .Q(_zygsfis_get_config_data_req[2]));
Q_FDP4EP \_zygsfis_get_config_data_req_REG[1] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1134), .R(n1750), .D(n574), .Q(_zygsfis_get_config_data_req[1]));
Q_INV U5719 ( .A(_zygsfis_get_config_data_req[0]), .Z(n51));
Q_FDP4EP \_zygsfis_get_config_data_req_REG[0] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1134), .R(n1750), .D(n51), .Q(_zygsfis_get_config_data_req[0]));
Q_INV U5721 ( .A(_zyL94_iscX1c0_n), .Z(n50));
Q_FDP4EP _zyL94_iscX1c0_n_REG  ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n50), .Q(_zyL94_iscX1c0_n));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[63] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[63]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[62] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[62]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[61] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[61]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[60] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[60]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[59] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[59]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[58] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[58]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[57] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[57]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[56] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[56]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[55] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[55]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[54] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[54]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[53] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[53]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[52] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[52]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[51] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[51]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[50] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[50]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[49] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[49]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[48] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[48]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[47] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[47]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[46] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[46]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[45] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[45]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[44] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[44]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[43] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[43]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[42] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[42]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[41] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[41]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[40] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[40]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[39] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[39]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[38] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[38]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[37] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[37]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[36] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[36]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[35] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[35]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[34] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[34]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[33] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[33]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[32] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n1750), .Q(_zyL94_iscX1c0_i0[32]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[31] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n660), .Q(_zyL94_iscX1c0_i0[31]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[30] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n659), .Q(_zyL94_iscX1c0_i0[30]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[29] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n658), .Q(_zyL94_iscX1c0_i0[29]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[28] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n657), .Q(_zyL94_iscX1c0_i0[28]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[27] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n656), .Q(_zyL94_iscX1c0_i0[27]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[26] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n655), .Q(_zyL94_iscX1c0_i0[26]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[25] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n654), .Q(_zyL94_iscX1c0_i0[25]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[24] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n653), .Q(_zyL94_iscX1c0_i0[24]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[23] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n652), .Q(_zyL94_iscX1c0_i0[23]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[22] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n651), .Q(_zyL94_iscX1c0_i0[22]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[21] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n650), .Q(_zyL94_iscX1c0_i0[21]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[20] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n649), .Q(_zyL94_iscX1c0_i0[20]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[19] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n648), .Q(_zyL94_iscX1c0_i0[19]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[18] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n647), .Q(_zyL94_iscX1c0_i0[18]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[17] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n646), .Q(_zyL94_iscX1c0_i0[17]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[16] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n645), .Q(_zyL94_iscX1c0_i0[16]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[15] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n644), .Q(_zyL94_iscX1c0_i0[15]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[14] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n643), .Q(_zyL94_iscX1c0_i0[14]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[13] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n642), .Q(_zyL94_iscX1c0_i0[13]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[12] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n641), .Q(_zyL94_iscX1c0_i0[12]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[11] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n640), .Q(_zyL94_iscX1c0_i0[11]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[10] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n639), .Q(_zyL94_iscX1c0_i0[10]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[9] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n638), .Q(_zyL94_iscX1c0_i0[9]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[8] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n637), .Q(_zyL94_iscX1c0_i0[8]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[7] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n636), .Q(_zyL94_iscX1c0_i0[7]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[6] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n635), .Q(_zyL94_iscX1c0_i0[6]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[5] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n634), .Q(_zyL94_iscX1c0_i0[5]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[4] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n633), .Q(_zyL94_iscX1c0_i0[4]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[3] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n632), .Q(_zyL94_iscX1c0_i0[3]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[2] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n631), .Q(_zyL94_iscX1c0_i0[2]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[1] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n630), .Q(_zyL94_iscX1c0_i0[1]));
Q_FDP4EP \_zyL94_iscX1c0_i0_REG[0] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1135), .R(n1750), .D(n629), .Q(_zyL94_iscX1c0_i0[0]));
Q_INV U5787 ( .A(_zyL61_iscX2c0_n), .Z(n49));
Q_FDP4EP _zyL61_iscX2c0_n_REG  ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n49), .Q(_zyL61_iscX2c0_n));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[63] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[63]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[62] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[62]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[61] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[61]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[60] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[60]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[59] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[59]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[58] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[58]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[57] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[57]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[56] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[56]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[55] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[55]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[54] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[54]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[53] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[53]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[52] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[52]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[51] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[51]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[50] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[50]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[49] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[49]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[48] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[48]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[47] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[47]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[46] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[46]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[45] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[45]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[44] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[44]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[43] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[43]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[42] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[42]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[41] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[41]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[40] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[40]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[39] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[39]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[38] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[38]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[37] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[37]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[36] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[36]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[35] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[35]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[34] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[34]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[33] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[33]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[32] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n1750), .Q(_zyL61_iscX2c0_i0[32]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[31] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n660), .Q(_zyL61_iscX2c0_i0[31]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[30] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n659), .Q(_zyL61_iscX2c0_i0[30]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[29] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n658), .Q(_zyL61_iscX2c0_i0[29]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[28] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n657), .Q(_zyL61_iscX2c0_i0[28]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[27] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n656), .Q(_zyL61_iscX2c0_i0[27]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[26] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n655), .Q(_zyL61_iscX2c0_i0[26]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[25] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n654), .Q(_zyL61_iscX2c0_i0[25]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[24] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n653), .Q(_zyL61_iscX2c0_i0[24]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[23] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n652), .Q(_zyL61_iscX2c0_i0[23]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[22] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n651), .Q(_zyL61_iscX2c0_i0[22]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[21] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n650), .Q(_zyL61_iscX2c0_i0[21]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[20] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n649), .Q(_zyL61_iscX2c0_i0[20]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[19] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n648), .Q(_zyL61_iscX2c0_i0[19]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[18] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n647), .Q(_zyL61_iscX2c0_i0[18]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[17] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n646), .Q(_zyL61_iscX2c0_i0[17]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[16] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n645), .Q(_zyL61_iscX2c0_i0[16]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[15] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n644), .Q(_zyL61_iscX2c0_i0[15]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[14] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n643), .Q(_zyL61_iscX2c0_i0[14]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[13] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n642), .Q(_zyL61_iscX2c0_i0[13]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[12] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n641), .Q(_zyL61_iscX2c0_i0[12]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[11] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n640), .Q(_zyL61_iscX2c0_i0[11]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[10] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n639), .Q(_zyL61_iscX2c0_i0[10]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[9] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n638), .Q(_zyL61_iscX2c0_i0[9]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[8] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n637), .Q(_zyL61_iscX2c0_i0[8]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[7] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n636), .Q(_zyL61_iscX2c0_i0[7]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[6] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n635), .Q(_zyL61_iscX2c0_i0[6]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[5] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n634), .Q(_zyL61_iscX2c0_i0[5]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[4] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n633), .Q(_zyL61_iscX2c0_i0[4]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[3] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n632), .Q(_zyL61_iscX2c0_i0[3]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[2] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n631), .Q(_zyL61_iscX2c0_i0[2]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[1] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n630), .Q(_zyL61_iscX2c0_i0[1]));
Q_FDP4EP \_zyL61_iscX2c0_i0_REG[0] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n629), .Q(_zyL61_iscX2c0_i0[0]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[31] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n692), .Q(_zyL61_iscX2c0_i1[31]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[30] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n691), .Q(_zyL61_iscX2c0_i1[30]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[29] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n690), .Q(_zyL61_iscX2c0_i1[29]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[28] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n689), .Q(_zyL61_iscX2c0_i1[28]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[27] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n688), .Q(_zyL61_iscX2c0_i1[27]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[26] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n687), .Q(_zyL61_iscX2c0_i1[26]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[25] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n686), .Q(_zyL61_iscX2c0_i1[25]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[24] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n685), .Q(_zyL61_iscX2c0_i1[24]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[23] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n684), .Q(_zyL61_iscX2c0_i1[23]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[22] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n683), .Q(_zyL61_iscX2c0_i1[22]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[21] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n682), .Q(_zyL61_iscX2c0_i1[21]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[20] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n681), .Q(_zyL61_iscX2c0_i1[20]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[19] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n680), .Q(_zyL61_iscX2c0_i1[19]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[18] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n679), .Q(_zyL61_iscX2c0_i1[18]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[17] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n678), .Q(_zyL61_iscX2c0_i1[17]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[16] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n677), .Q(_zyL61_iscX2c0_i1[16]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[15] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n676), .Q(_zyL61_iscX2c0_i1[15]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[14] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n675), .Q(_zyL61_iscX2c0_i1[14]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[13] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n674), .Q(_zyL61_iscX2c0_i1[13]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[12] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n673), .Q(_zyL61_iscX2c0_i1[12]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[11] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n672), .Q(_zyL61_iscX2c0_i1[11]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[10] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n671), .Q(_zyL61_iscX2c0_i1[10]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[9] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n670), .Q(_zyL61_iscX2c0_i1[9]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[8] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n669), .Q(_zyL61_iscX2c0_i1[8]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[7] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n668), .Q(_zyL61_iscX2c0_i1[7]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[6] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n667), .Q(_zyL61_iscX2c0_i1[6]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[5] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n666), .Q(_zyL61_iscX2c0_i1[5]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[4] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n665), .Q(_zyL61_iscX2c0_i1[4]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[3] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n664), .Q(_zyL61_iscX2c0_i1[3]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[2] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n663), .Q(_zyL61_iscX2c0_i1[2]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[1] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n662), .Q(_zyL61_iscX2c0_i1[1]));
Q_FDP4EP \_zyL61_iscX2c0_i1_REG[0] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1136), .R(n1750), .D(n661), .Q(_zyL61_iscX2c0_i1[0]));
Q_FDP4EP _zyGfifoF0_L324_s3_req_1_REG  ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n922), .Q(_zyGfifoF0_L324_s3_req_1));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[95] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n996), .Q(_zyGfifoF0_L324_s3_data_1[95]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[94] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n995), .Q(_zyGfifoF0_L324_s3_data_1[94]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[93] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n994), .Q(_zyGfifoF0_L324_s3_data_1[93]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[92] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n993), .Q(_zyGfifoF0_L324_s3_data_1[92]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[91] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n992), .Q(_zyGfifoF0_L324_s3_data_1[91]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[90] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n991), .Q(_zyGfifoF0_L324_s3_data_1[90]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[89] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n990), .Q(_zyGfifoF0_L324_s3_data_1[89]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[88] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n989), .Q(_zyGfifoF0_L324_s3_data_1[88]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[87] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n988), .Q(_zyGfifoF0_L324_s3_data_1[87]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[86] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n987), .Q(_zyGfifoF0_L324_s3_data_1[86]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[85] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n986), .Q(_zyGfifoF0_L324_s3_data_1[85]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[84] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n985), .Q(_zyGfifoF0_L324_s3_data_1[84]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[83] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n984), .Q(_zyGfifoF0_L324_s3_data_1[83]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[82] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n983), .Q(_zyGfifoF0_L324_s3_data_1[82]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[81] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n982), .Q(_zyGfifoF0_L324_s3_data_1[81]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[80] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n981), .Q(_zyGfifoF0_L324_s3_data_1[80]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[79] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n980), .Q(_zyGfifoF0_L324_s3_data_1[79]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[78] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n979), .Q(_zyGfifoF0_L324_s3_data_1[78]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[77] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n978), .Q(_zyGfifoF0_L324_s3_data_1[77]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[76] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n977), .Q(_zyGfifoF0_L324_s3_data_1[76]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[75] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n976), .Q(_zyGfifoF0_L324_s3_data_1[75]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[74] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n975), .Q(_zyGfifoF0_L324_s3_data_1[74]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[73] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n974), .Q(_zyGfifoF0_L324_s3_data_1[73]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[72] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n973), .Q(_zyGfifoF0_L324_s3_data_1[72]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[71] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n972), .Q(_zyGfifoF0_L324_s3_data_1[71]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[70] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n971), .Q(_zyGfifoF0_L324_s3_data_1[70]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[69] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n970), .Q(_zyGfifoF0_L324_s3_data_1[69]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[68] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n969), .Q(_zyGfifoF0_L324_s3_data_1[68]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[67] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n968), .Q(_zyGfifoF0_L324_s3_data_1[67]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[66] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n967), .Q(_zyGfifoF0_L324_s3_data_1[66]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[65] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n920), .Q(_zyGfifoF0_L324_s3_data_1[65]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[64] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n919), .Q(_zyGfifoF0_L324_s3_data_1[64]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[63] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n918), .Q(_zyGfifoF0_L324_s3_data_1[63]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[62] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n917), .Q(_zyGfifoF0_L324_s3_data_1[62]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[61] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n916), .Q(_zyGfifoF0_L324_s3_data_1[61]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[60] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n915), .Q(_zyGfifoF0_L324_s3_data_1[60]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[59] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n914), .Q(_zyGfifoF0_L324_s3_data_1[59]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[58] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n913), .Q(_zyGfifoF0_L324_s3_data_1[58]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[57] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n912), .Q(_zyGfifoF0_L324_s3_data_1[57]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[56] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n911), .Q(_zyGfifoF0_L324_s3_data_1[56]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[55] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n910), .Q(_zyGfifoF0_L324_s3_data_1[55]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[54] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n909), .Q(_zyGfifoF0_L324_s3_data_1[54]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[53] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n908), .Q(_zyGfifoF0_L324_s3_data_1[53]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[52] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n907), .Q(_zyGfifoF0_L324_s3_data_1[52]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[51] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n906), .Q(_zyGfifoF0_L324_s3_data_1[51]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[50] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n905), .Q(_zyGfifoF0_L324_s3_data_1[50]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[49] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n904), .Q(_zyGfifoF0_L324_s3_data_1[49]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[48] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n903), .Q(_zyGfifoF0_L324_s3_data_1[48]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[47] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n902), .Q(_zyGfifoF0_L324_s3_data_1[47]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[46] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n901), .Q(_zyGfifoF0_L324_s3_data_1[46]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[45] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n900), .Q(_zyGfifoF0_L324_s3_data_1[45]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[44] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n899), .Q(_zyGfifoF0_L324_s3_data_1[44]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[43] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n898), .Q(_zyGfifoF0_L324_s3_data_1[43]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[42] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n897), .Q(_zyGfifoF0_L324_s3_data_1[42]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[41] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n896), .Q(_zyGfifoF0_L324_s3_data_1[41]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[40] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n895), .Q(_zyGfifoF0_L324_s3_data_1[40]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[39] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n894), .Q(_zyGfifoF0_L324_s3_data_1[39]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[38] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n893), .Q(_zyGfifoF0_L324_s3_data_1[38]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[37] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n892), .Q(_zyGfifoF0_L324_s3_data_1[37]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[36] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n891), .Q(_zyGfifoF0_L324_s3_data_1[36]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[35] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n890), .Q(_zyGfifoF0_L324_s3_data_1[35]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[34] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n889), .Q(_zyGfifoF0_L324_s3_data_1[34]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[33] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n888), .Q(_zyGfifoF0_L324_s3_data_1[33]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[32] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n887), .Q(_zyGfifoF0_L324_s3_data_1[32]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[31] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n886), .Q(_zyGfifoF0_L324_s3_data_1[31]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[30] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n884), .Q(_zyGfifoF0_L324_s3_data_1[30]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[29] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n882), .Q(_zyGfifoF0_L324_s3_data_1[29]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[28] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n880), .Q(_zyGfifoF0_L324_s3_data_1[28]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[27] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n878), .Q(_zyGfifoF0_L324_s3_data_1[27]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[26] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n876), .Q(_zyGfifoF0_L324_s3_data_1[26]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[25] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n874), .Q(_zyGfifoF0_L324_s3_data_1[25]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[24] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n872), .Q(_zyGfifoF0_L324_s3_data_1[24]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[23] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n870), .Q(_zyGfifoF0_L324_s3_data_1[23]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[22] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n868), .Q(_zyGfifoF0_L324_s3_data_1[22]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[21] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n866), .Q(_zyGfifoF0_L324_s3_data_1[21]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[20] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n864), .Q(_zyGfifoF0_L324_s3_data_1[20]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[19] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n862), .Q(_zyGfifoF0_L324_s3_data_1[19]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[18] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n860), .Q(_zyGfifoF0_L324_s3_data_1[18]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[17] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n858), .Q(_zyGfifoF0_L324_s3_data_1[17]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[16] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n856), .Q(_zyGfifoF0_L324_s3_data_1[16]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[15] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n854), .Q(_zyGfifoF0_L324_s3_data_1[15]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[14] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n852), .Q(_zyGfifoF0_L324_s3_data_1[14]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[13] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n850), .Q(_zyGfifoF0_L324_s3_data_1[13]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[12] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n848), .Q(_zyGfifoF0_L324_s3_data_1[12]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[11] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n846), .Q(_zyGfifoF0_L324_s3_data_1[11]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[10] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n844), .Q(_zyGfifoF0_L324_s3_data_1[10]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[9] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n842), .Q(_zyGfifoF0_L324_s3_data_1[9]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[8] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n840), .Q(_zyGfifoF0_L324_s3_data_1[8]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[7] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n838), .Q(_zyGfifoF0_L324_s3_data_1[7]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[6] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n836), .Q(_zyGfifoF0_L324_s3_data_1[6]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[5] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n834), .Q(_zyGfifoF0_L324_s3_data_1[5]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[4] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n832), .Q(_zyGfifoF0_L324_s3_data_1[4]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[3] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n831), .Q(_zyGfifoF0_L324_s3_data_1[3]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[2] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n830), .Q(_zyGfifoF0_L324_s3_data_1[2]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[1] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n829), .Q(_zyGfifoF0_L324_s3_data_1[1]));
Q_FDP4EP \_zyGfifoF0_L324_s3_data_1_REG[0] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n828), .Q(_zyGfifoF0_L324_s3_data_1[0]));
Q_FDP4EP \_zyGfifoF0_L324_s3_cbid_1_REG[19] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n827), .Q(_zyGfifoF0_L324_s3_cbid_1[19]));
Q_FDP4EP \_zyGfifoF0_L324_s3_cbid_1_REG[18] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n826), .Q(_zyGfifoF0_L324_s3_cbid_1[18]));
Q_FDP4EP \_zyGfifoF0_L324_s3_cbid_1_REG[17] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n825), .Q(_zyGfifoF0_L324_s3_cbid_1[17]));
Q_FDP4EP \_zyGfifoF0_L324_s3_cbid_1_REG[16] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n824), .Q(_zyGfifoF0_L324_s3_cbid_1[16]));
Q_FDP4EP \_zyGfifoF0_L324_s3_cbid_1_REG[15] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n823), .Q(_zyGfifoF0_L324_s3_cbid_1[15]));
Q_FDP4EP \_zyGfifoF0_L324_s3_cbid_1_REG[14] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n822), .Q(_zyGfifoF0_L324_s3_cbid_1[14]));
Q_FDP4EP \_zyGfifoF0_L324_s3_cbid_1_REG[13] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n821), .Q(_zyGfifoF0_L324_s3_cbid_1[13]));
Q_FDP4EP \_zyGfifoF0_L324_s3_cbid_1_REG[12] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n820), .Q(_zyGfifoF0_L324_s3_cbid_1[12]));
Q_FDP4EP \_zyGfifoF0_L324_s3_cbid_1_REG[11] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n819), .Q(_zyGfifoF0_L324_s3_cbid_1[11]));
Q_FDP4EP \_zyGfifoF0_L324_s3_cbid_1_REG[10] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n818), .Q(_zyGfifoF0_L324_s3_cbid_1[10]));
Q_FDP4EP \_zyGfifoF0_L324_s3_cbid_1_REG[9] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n817), .Q(_zyGfifoF0_L324_s3_cbid_1[9]));
Q_FDP4EP \_zyGfifoF0_L324_s3_cbid_1_REG[8] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n816), .Q(_zyGfifoF0_L324_s3_cbid_1[8]));
Q_FDP4EP \_zyGfifoF0_L324_s3_cbid_1_REG[7] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n815), .Q(_zyGfifoF0_L324_s3_cbid_1[7]));
Q_FDP4EP \_zyGfifoF0_L324_s3_cbid_1_REG[6] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n814), .Q(_zyGfifoF0_L324_s3_cbid_1[6]));
Q_FDP4EP \_zyGfifoF0_L324_s3_cbid_1_REG[5] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n813), .Q(_zyGfifoF0_L324_s3_cbid_1[5]));
Q_FDP4EP \_zyGfifoF0_L324_s3_cbid_1_REG[4] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n812), .Q(_zyGfifoF0_L324_s3_cbid_1[4]));
Q_FDP4EP \_zyGfifoF0_L324_s3_cbid_1_REG[3] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n811), .Q(_zyGfifoF0_L324_s3_cbid_1[3]));
Q_FDP4EP \_zyGfifoF0_L324_s3_cbid_1_REG[2] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n810), .Q(_zyGfifoF0_L324_s3_cbid_1[2]));
Q_FDP4EP \_zyGfifoF0_L324_s3_cbid_1_REG[1] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n809), .Q(_zyGfifoF0_L324_s3_cbid_1[1]));
Q_FDP4EP \_zyGfifoF0_L324_s3_cbid_1_REG[0] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n808), .Q(_zyGfifoF0_L324_s3_cbid_1[0]));
Q_INV U6002 ( .A(n1026), .Z(n48));
Q_FDP4EP _zyGfifoF1_L324_s2_req_2_REG  ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n807), .Q(_zyGfifoF1_L324_s2_req_2));
Q_FDP4EP \_zyGfifoF1_L324_s2_cbid_2_REG[19] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n806), .Q(_zyGfifoF1_L324_s2_cbid_2[19]));
Q_FDP4EP \_zyGfifoF1_L324_s2_cbid_2_REG[18] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n805), .Q(_zyGfifoF1_L324_s2_cbid_2[18]));
Q_FDP4EP \_zyGfifoF1_L324_s2_cbid_2_REG[17] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n804), .Q(_zyGfifoF1_L324_s2_cbid_2[17]));
Q_FDP4EP \_zyGfifoF1_L324_s2_cbid_2_REG[16] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n803), .Q(_zyGfifoF1_L324_s2_cbid_2[16]));
Q_FDP4EP \_zyGfifoF1_L324_s2_cbid_2_REG[15] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n802), .Q(_zyGfifoF1_L324_s2_cbid_2[15]));
Q_FDP4EP \_zyGfifoF1_L324_s2_cbid_2_REG[14] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n801), .Q(_zyGfifoF1_L324_s2_cbid_2[14]));
Q_FDP4EP \_zyGfifoF1_L324_s2_cbid_2_REG[13] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n800), .Q(_zyGfifoF1_L324_s2_cbid_2[13]));
Q_FDP4EP \_zyGfifoF1_L324_s2_cbid_2_REG[12] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n799), .Q(_zyGfifoF1_L324_s2_cbid_2[12]));
Q_FDP4EP \_zyGfifoF1_L324_s2_cbid_2_REG[11] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n798), .Q(_zyGfifoF1_L324_s2_cbid_2[11]));
Q_FDP4EP \_zyGfifoF1_L324_s2_cbid_2_REG[10] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n797), .Q(_zyGfifoF1_L324_s2_cbid_2[10]));
Q_FDP4EP \_zyGfifoF1_L324_s2_cbid_2_REG[9] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n796), .Q(_zyGfifoF1_L324_s2_cbid_2[9]));
Q_FDP4EP \_zyGfifoF1_L324_s2_cbid_2_REG[8] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n795), .Q(_zyGfifoF1_L324_s2_cbid_2[8]));
Q_FDP4EP \_zyGfifoF1_L324_s2_cbid_2_REG[7] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n794), .Q(_zyGfifoF1_L324_s2_cbid_2[7]));
Q_FDP4EP \_zyGfifoF1_L324_s2_cbid_2_REG[6] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n793), .Q(_zyGfifoF1_L324_s2_cbid_2[6]));
Q_FDP4EP \_zyGfifoF1_L324_s2_cbid_2_REG[5] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n792), .Q(_zyGfifoF1_L324_s2_cbid_2[5]));
Q_FDP4EP \_zyGfifoF1_L324_s2_cbid_2_REG[4] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n791), .Q(_zyGfifoF1_L324_s2_cbid_2[4]));
Q_FDP4EP \_zyGfifoF1_L324_s2_cbid_2_REG[3] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n790), .Q(_zyGfifoF1_L324_s2_cbid_2[3]));
Q_FDP4EP \_zyGfifoF1_L324_s2_cbid_2_REG[2] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n789), .Q(_zyGfifoF1_L324_s2_cbid_2[2]));
Q_FDP4EP \_zyGfifoF1_L324_s2_cbid_2_REG[1] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n788), .Q(_zyGfifoF1_L324_s2_cbid_2[1]));
Q_FDP4EP \_zyGfifoF1_L324_s2_cbid_2_REG[0] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n787), .Q(_zyGfifoF1_L324_s2_cbid_2[0]));
Q_FDP4EP _zyGfifoF2_L324_s2_req_3_REG  ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n786), .Q(_zyGfifoF2_L324_s2_req_3));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[71] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n785), .Q(_zyGfifoF2_L324_s2_data_3[71]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[70] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n784), .Q(_zyGfifoF2_L324_s2_data_3[70]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[69] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n783), .Q(_zyGfifoF2_L324_s2_data_3[69]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[68] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n782), .Q(_zyGfifoF2_L324_s2_data_3[68]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[67] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n781), .Q(_zyGfifoF2_L324_s2_data_3[67]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[66] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n780), .Q(_zyGfifoF2_L324_s2_data_3[66]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[65] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n779), .Q(_zyGfifoF2_L324_s2_data_3[65]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[64] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n778), .Q(_zyGfifoF2_L324_s2_data_3[64]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[63] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n777), .Q(_zyGfifoF2_L324_s2_data_3[63]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[62] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n776), .Q(_zyGfifoF2_L324_s2_data_3[62]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[61] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n775), .Q(_zyGfifoF2_L324_s2_data_3[61]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[60] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n774), .Q(_zyGfifoF2_L324_s2_data_3[60]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[59] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n773), .Q(_zyGfifoF2_L324_s2_data_3[59]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[58] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n772), .Q(_zyGfifoF2_L324_s2_data_3[58]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[57] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n771), .Q(_zyGfifoF2_L324_s2_data_3[57]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[56] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n770), .Q(_zyGfifoF2_L324_s2_data_3[56]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[55] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n769), .Q(_zyGfifoF2_L324_s2_data_3[55]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[54] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n768), .Q(_zyGfifoF2_L324_s2_data_3[54]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[53] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n767), .Q(_zyGfifoF2_L324_s2_data_3[53]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[52] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n766), .Q(_zyGfifoF2_L324_s2_data_3[52]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[51] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n765), .Q(_zyGfifoF2_L324_s2_data_3[51]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[50] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n764), .Q(_zyGfifoF2_L324_s2_data_3[50]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[49] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n763), .Q(_zyGfifoF2_L324_s2_data_3[49]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[48] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n762), .Q(_zyGfifoF2_L324_s2_data_3[48]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[47] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n761), .Q(_zyGfifoF2_L324_s2_data_3[47]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[46] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n760), .Q(_zyGfifoF2_L324_s2_data_3[46]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[45] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n759), .Q(_zyGfifoF2_L324_s2_data_3[45]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[44] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n758), .Q(_zyGfifoF2_L324_s2_data_3[44]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[43] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n757), .Q(_zyGfifoF2_L324_s2_data_3[43]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[42] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n756), .Q(_zyGfifoF2_L324_s2_data_3[42]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[41] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n755), .Q(_zyGfifoF2_L324_s2_data_3[41]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[40] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n754), .Q(_zyGfifoF2_L324_s2_data_3[40]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[39] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n753), .Q(_zyGfifoF2_L324_s2_data_3[39]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[38] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n752), .Q(_zyGfifoF2_L324_s2_data_3[38]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[37] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n751), .Q(_zyGfifoF2_L324_s2_data_3[37]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[36] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n750), .Q(_zyGfifoF2_L324_s2_data_3[36]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[35] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n749), .Q(_zyGfifoF2_L324_s2_data_3[35]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[34] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n748), .Q(_zyGfifoF2_L324_s2_data_3[34]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[33] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n747), .Q(_zyGfifoF2_L324_s2_data_3[33]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[32] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n746), .Q(_zyGfifoF2_L324_s2_data_3[32]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[31] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n745), .Q(_zyGfifoF2_L324_s2_data_3[31]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[30] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n744), .Q(_zyGfifoF2_L324_s2_data_3[30]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[29] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n743), .Q(_zyGfifoF2_L324_s2_data_3[29]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[28] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n742), .Q(_zyGfifoF2_L324_s2_data_3[28]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[27] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n741), .Q(_zyGfifoF2_L324_s2_data_3[27]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[26] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n740), .Q(_zyGfifoF2_L324_s2_data_3[26]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[25] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n739), .Q(_zyGfifoF2_L324_s2_data_3[25]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[24] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n738), .Q(_zyGfifoF2_L324_s2_data_3[24]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[23] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n737), .Q(_zyGfifoF2_L324_s2_data_3[23]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[22] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n736), .Q(_zyGfifoF2_L324_s2_data_3[22]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[21] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n735), .Q(_zyGfifoF2_L324_s2_data_3[21]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[20] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n734), .Q(_zyGfifoF2_L324_s2_data_3[20]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[19] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n733), .Q(_zyGfifoF2_L324_s2_data_3[19]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[18] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n732), .Q(_zyGfifoF2_L324_s2_data_3[18]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[17] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n731), .Q(_zyGfifoF2_L324_s2_data_3[17]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[16] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n730), .Q(_zyGfifoF2_L324_s2_data_3[16]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[15] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n729), .Q(_zyGfifoF2_L324_s2_data_3[15]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[14] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n728), .Q(_zyGfifoF2_L324_s2_data_3[14]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[13] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n727), .Q(_zyGfifoF2_L324_s2_data_3[13]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[12] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n726), .Q(_zyGfifoF2_L324_s2_data_3[12]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[11] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n725), .Q(_zyGfifoF2_L324_s2_data_3[11]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[10] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n724), .Q(_zyGfifoF2_L324_s2_data_3[10]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[9] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n723), .Q(_zyGfifoF2_L324_s2_data_3[9]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[8] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n722), .Q(_zyGfifoF2_L324_s2_data_3[8]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[7] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n721), .Q(_zyGfifoF2_L324_s2_data_3[7]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[6] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n720), .Q(_zyGfifoF2_L324_s2_data_3[6]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[5] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n719), .Q(_zyGfifoF2_L324_s2_data_3[5]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[4] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n718), .Q(_zyGfifoF2_L324_s2_data_3[4]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[3] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n717), .Q(_zyGfifoF2_L324_s2_data_3[3]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[2] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n716), .Q(_zyGfifoF2_L324_s2_data_3[2]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[1] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n715), .Q(_zyGfifoF2_L324_s2_data_3[1]));
Q_FDP4EP \_zyGfifoF2_L324_s2_data_3_REG[0] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n714), .Q(_zyGfifoF2_L324_s2_data_3[0]));
Q_FDP4EP \_zyGfifoF2_L324_s2_cbid_3_REG[19] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n713), .Q(_zyGfifoF2_L324_s2_cbid_3[19]));
Q_FDP4EP \_zyGfifoF2_L324_s2_cbid_3_REG[18] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n712), .Q(_zyGfifoF2_L324_s2_cbid_3[18]));
Q_FDP4EP \_zyGfifoF2_L324_s2_cbid_3_REG[17] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n711), .Q(_zyGfifoF2_L324_s2_cbid_3[17]));
Q_FDP4EP \_zyGfifoF2_L324_s2_cbid_3_REG[16] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n710), .Q(_zyGfifoF2_L324_s2_cbid_3[16]));
Q_FDP4EP \_zyGfifoF2_L324_s2_cbid_3_REG[15] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n709), .Q(_zyGfifoF2_L324_s2_cbid_3[15]));
Q_FDP4EP \_zyGfifoF2_L324_s2_cbid_3_REG[14] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n708), .Q(_zyGfifoF2_L324_s2_cbid_3[14]));
Q_FDP4EP \_zyGfifoF2_L324_s2_cbid_3_REG[13] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n707), .Q(_zyGfifoF2_L324_s2_cbid_3[13]));
Q_FDP4EP \_zyGfifoF2_L324_s2_cbid_3_REG[12] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n706), .Q(_zyGfifoF2_L324_s2_cbid_3[12]));
Q_FDP4EP \_zyGfifoF2_L324_s2_cbid_3_REG[11] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n705), .Q(_zyGfifoF2_L324_s2_cbid_3[11]));
Q_FDP4EP \_zyGfifoF2_L324_s2_cbid_3_REG[10] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n704), .Q(_zyGfifoF2_L324_s2_cbid_3[10]));
Q_FDP4EP \_zyGfifoF2_L324_s2_cbid_3_REG[9] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n703), .Q(_zyGfifoF2_L324_s2_cbid_3[9]));
Q_FDP4EP \_zyGfifoF2_L324_s2_cbid_3_REG[8] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n702), .Q(_zyGfifoF2_L324_s2_cbid_3[8]));
Q_FDP4EP \_zyGfifoF2_L324_s2_cbid_3_REG[7] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n701), .Q(_zyGfifoF2_L324_s2_cbid_3[7]));
Q_FDP4EP \_zyGfifoF2_L324_s2_cbid_3_REG[6] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n700), .Q(_zyGfifoF2_L324_s2_cbid_3[6]));
Q_FDP4EP \_zyGfifoF2_L324_s2_cbid_3_REG[5] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n699), .Q(_zyGfifoF2_L324_s2_cbid_3[5]));
Q_FDP4EP \_zyGfifoF2_L324_s2_cbid_3_REG[4] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n698), .Q(_zyGfifoF2_L324_s2_cbid_3[4]));
Q_FDP4EP \_zyGfifoF2_L324_s2_cbid_3_REG[3] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n697), .Q(_zyGfifoF2_L324_s2_cbid_3[3]));
Q_FDP4EP \_zyGfifoF2_L324_s2_cbid_3_REG[2] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n696), .Q(_zyGfifoF2_L324_s2_cbid_3[2]));
Q_FDP4EP \_zyGfifoF2_L324_s2_cbid_3_REG[1] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n695), .Q(_zyGfifoF2_L324_s2_cbid_3[1]));
Q_FDP4EP \_zyGfifoF2_L324_s2_cbid_3_REG[0] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n694), .Q(_zyGfifoF2_L324_s2_cbid_3[0]));
Q_INV U6117 ( .A(n1027), .Z(n47));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[1] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1133), .Q(_zyxr_L206_tfiV3_M2_pbcG3[1]));
Q_INV U6119 ( .A(n1050), .Z(n46));
Q_FDP4EP response_REG  ( .CK(_zyM2L324_pbcMevClk4), .CE(n46), .R(n1750), .D(n693), .Q(response));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[31] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n660), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[31]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[30] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n659), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[30]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[29] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n658), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[29]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[28] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n657), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[28]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[27] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n656), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[27]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[26] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n655), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[26]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[25] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n654), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[25]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[24] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n653), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[24]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[23] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n652), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[23]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[22] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n651), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[22]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[21] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n650), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[21]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[20] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n649), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[20]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[19] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n648), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[19]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[18] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n647), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[18]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[17] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n646), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[17]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[16] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n645), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[16]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[15] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n644), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[15]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[14] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n643), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[14]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[13] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n642), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[13]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[12] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n641), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[12]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[11] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n640), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[11]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[10] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n639), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[10]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[9] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n638), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[9]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[8] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n637), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[8]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[7] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n636), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[7]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[6] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n635), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[6]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[5] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n634), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[5]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[4] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n633), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[4]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[3] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n632), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[3]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[2] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n631), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[2]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[1] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n630), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[1]));
Q_FDP4EP \_zyaddress_L206_tfiV1_M2_pbcG1_REG[0] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n629), .Q(_zyaddress_L206_tfiV1_M2_pbcG1[0]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[31] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n692), .Q(_zydata_L206_tfiV2_M2_pbcG2[31]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[30] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n691), .Q(_zydata_L206_tfiV2_M2_pbcG2[30]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[29] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n690), .Q(_zydata_L206_tfiV2_M2_pbcG2[29]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[28] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n689), .Q(_zydata_L206_tfiV2_M2_pbcG2[28]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[27] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n688), .Q(_zydata_L206_tfiV2_M2_pbcG2[27]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[26] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n687), .Q(_zydata_L206_tfiV2_M2_pbcG2[26]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[25] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n686), .Q(_zydata_L206_tfiV2_M2_pbcG2[25]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[24] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n685), .Q(_zydata_L206_tfiV2_M2_pbcG2[24]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[23] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n684), .Q(_zydata_L206_tfiV2_M2_pbcG2[23]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[22] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n683), .Q(_zydata_L206_tfiV2_M2_pbcG2[22]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[21] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n682), .Q(_zydata_L206_tfiV2_M2_pbcG2[21]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[20] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n681), .Q(_zydata_L206_tfiV2_M2_pbcG2[20]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[19] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n680), .Q(_zydata_L206_tfiV2_M2_pbcG2[19]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[18] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n679), .Q(_zydata_L206_tfiV2_M2_pbcG2[18]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[17] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n678), .Q(_zydata_L206_tfiV2_M2_pbcG2[17]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[16] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n677), .Q(_zydata_L206_tfiV2_M2_pbcG2[16]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[15] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n676), .Q(_zydata_L206_tfiV2_M2_pbcG2[15]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[14] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n675), .Q(_zydata_L206_tfiV2_M2_pbcG2[14]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[13] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n674), .Q(_zydata_L206_tfiV2_M2_pbcG2[13]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[12] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n673), .Q(_zydata_L206_tfiV2_M2_pbcG2[12]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[11] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n672), .Q(_zydata_L206_tfiV2_M2_pbcG2[11]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[10] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n671), .Q(_zydata_L206_tfiV2_M2_pbcG2[10]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[9] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n670), .Q(_zydata_L206_tfiV2_M2_pbcG2[9]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[8] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n669), .Q(_zydata_L206_tfiV2_M2_pbcG2[8]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[7] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n668), .Q(_zydata_L206_tfiV2_M2_pbcG2[7]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[6] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n667), .Q(_zydata_L206_tfiV2_M2_pbcG2[6]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[5] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n666), .Q(_zydata_L206_tfiV2_M2_pbcG2[5]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[4] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n665), .Q(_zydata_L206_tfiV2_M2_pbcG2[4]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[3] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n664), .Q(_zydata_L206_tfiV2_M2_pbcG2[3]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[2] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n663), .Q(_zydata_L206_tfiV2_M2_pbcG2[2]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[1] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n662), .Q(_zydata_L206_tfiV2_M2_pbcG2[1]));
Q_FDP4EP \_zydata_L206_tfiV2_M2_pbcG2_REG[0] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n661), .Q(_zydata_L206_tfiV2_M2_pbcG2[0]));
Q_FDP4EP \address_REG[31] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n660), .Q(address[31]));
Q_FDP4EP \address_REG[30] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n659), .Q(address[30]));
Q_FDP4EP \address_REG[29] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n658), .Q(address[29]));
Q_FDP4EP \address_REG[28] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n657), .Q(address[28]));
Q_FDP4EP \address_REG[27] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n656), .Q(address[27]));
Q_FDP4EP \address_REG[26] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n655), .Q(address[26]));
Q_FDP4EP \address_REG[25] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n654), .Q(address[25]));
Q_FDP4EP \address_REG[24] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n653), .Q(address[24]));
Q_FDP4EP \address_REG[23] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n652), .Q(address[23]));
Q_FDP4EP \address_REG[22] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n651), .Q(address[22]));
Q_FDP4EP \address_REG[21] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n650), .Q(address[21]));
Q_FDP4EP \address_REG[20] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n649), .Q(address[20]));
Q_FDP4EP \address_REG[19] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n648), .Q(address[19]));
Q_FDP4EP \address_REG[18] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n647), .Q(address[18]));
Q_FDP4EP \address_REG[17] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n646), .Q(address[17]));
Q_FDP4EP \address_REG[16] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n645), .Q(address[16]));
Q_FDP4EP \address_REG[15] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n644), .Q(address[15]));
Q_FDP4EP \address_REG[14] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n643), .Q(address[14]));
Q_FDP4EP \address_REG[13] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n642), .Q(address[13]));
Q_FDP4EP \address_REG[12] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n641), .Q(address[12]));
Q_FDP4EP \address_REG[11] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n640), .Q(address[11]));
Q_FDP4EP \address_REG[10] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n639), .Q(address[10]));
Q_FDP4EP \address_REG[9] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n638), .Q(address[9]));
Q_FDP4EP \address_REG[8] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n637), .Q(address[8]));
Q_FDP4EP \address_REG[7] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n636), .Q(address[7]));
Q_FDP4EP \address_REG[6] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n635), .Q(address[6]));
Q_FDP4EP \address_REG[5] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n634), .Q(address[5]));
Q_FDP4EP \address_REG[4] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n633), .Q(address[4]));
Q_FDP4EP \address_REG[3] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n632), .Q(address[3]));
Q_FDP4EP \address_REG[2] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n631), .Q(address[2]));
Q_FDP4EP \address_REG[1] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n630), .Q(address[1]));
Q_FDP4EP \address_REG[0] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n629), .Q(address[0]));
Q_FDP4EP \data_REG[31] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n692), .Q(data[31]));
Q_FDP4EP \data_REG[30] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n691), .Q(data[30]));
Q_FDP4EP \data_REG[29] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n690), .Q(data[29]));
Q_FDP4EP \data_REG[28] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n689), .Q(data[28]));
Q_FDP4EP \data_REG[27] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n688), .Q(data[27]));
Q_FDP4EP \data_REG[26] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n687), .Q(data[26]));
Q_FDP4EP \data_REG[25] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n686), .Q(data[25]));
Q_FDP4EP \data_REG[24] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n685), .Q(data[24]));
Q_FDP4EP \data_REG[23] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n684), .Q(data[23]));
Q_FDP4EP \data_REG[22] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n683), .Q(data[22]));
Q_FDP4EP \data_REG[21] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n682), .Q(data[21]));
Q_FDP4EP \data_REG[20] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n681), .Q(data[20]));
Q_FDP4EP \data_REG[19] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n680), .Q(data[19]));
Q_FDP4EP \data_REG[18] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n679), .Q(data[18]));
Q_FDP4EP \data_REG[17] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n678), .Q(data[17]));
Q_FDP4EP \data_REG[16] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n677), .Q(data[16]));
Q_FDP4EP \data_REG[15] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n676), .Q(data[15]));
Q_FDP4EP \data_REG[14] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n675), .Q(data[14]));
Q_FDP4EP \data_REG[13] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n674), .Q(data[13]));
Q_FDP4EP \data_REG[12] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n673), .Q(data[12]));
Q_FDP4EP \data_REG[11] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n672), .Q(data[11]));
Q_FDP4EP \data_REG[10] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n671), .Q(data[10]));
Q_FDP4EP \data_REG[9] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n670), .Q(data[9]));
Q_FDP4EP \data_REG[8] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n669), .Q(data[8]));
Q_FDP4EP \data_REG[7] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n668), .Q(data[7]));
Q_FDP4EP \data_REG[6] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n667), .Q(data[6]));
Q_FDP4EP \data_REG[5] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n666), .Q(data[5]));
Q_FDP4EP \data_REG[4] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n665), .Q(data[4]));
Q_FDP4EP \data_REG[3] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n664), .Q(data[3]));
Q_FDP4EP \data_REG[2] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n663), .Q(data[2]));
Q_FDP4EP \data_REG[1] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n662), .Q(data[1]));
Q_FDP4EP \data_REG[0] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n661), .Q(data[0]));
Q_FDP4EP \_zyoperation_L206_tfiV0_M2_pbcG0_REG[7] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1151), .Q(_zyoperation_L206_tfiV0_M2_pbcG0[7]));
Q_FDP4EP \_zyoperation_L206_tfiV0_M2_pbcG0_REG[6] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1150), .Q(_zyoperation_L206_tfiV0_M2_pbcG0[6]));
Q_FDP4EP \_zyoperation_L206_tfiV0_M2_pbcG0_REG[5] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1149), .Q(_zyoperation_L206_tfiV0_M2_pbcG0[5]));
Q_FDP4EP \_zyoperation_L206_tfiV0_M2_pbcG0_REG[4] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1148), .Q(_zyoperation_L206_tfiV0_M2_pbcG0[4]));
Q_FDP4EP \_zyoperation_L206_tfiV0_M2_pbcG0_REG[3] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1147), .Q(_zyoperation_L206_tfiV0_M2_pbcG0[3]));
Q_FDP4EP \_zyoperation_L206_tfiV0_M2_pbcG0_REG[2] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1146), .Q(_zyoperation_L206_tfiV0_M2_pbcG0[2]));
Q_FDP4EP \_zyoperation_L206_tfiV0_M2_pbcG0_REG[1] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1145), .Q(_zyoperation_L206_tfiV0_M2_pbcG0[1]));
Q_FDP4EP \_zyoperation_L206_tfiV0_M2_pbcG0_REG[0] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1144), .Q(_zyoperation_L206_tfiV0_M2_pbcG0[0]));
Q_FDP4EP \operation_REG[7] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1151), .Q(operation[7]));
Q_FDP4EP \operation_REG[6] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1150), .Q(operation[6]));
Q_FDP4EP \operation_REG[5] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1149), .Q(operation[5]));
Q_FDP4EP \operation_REG[4] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1148), .Q(operation[4]));
Q_FDP4EP \operation_REG[3] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1147), .Q(operation[3]));
Q_FDP4EP \operation_REG[2] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1146), .Q(operation[2]));
Q_FDP4EP \operation_REG[1] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1145), .Q(operation[1]));
Q_FDP4EP \operation_REG[0] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1144), .Q(operation[0]));
Q_FDP4EP \_zygsfis_get_config_data_rptr_REG[4] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n596), .Q(_zygsfis_get_config_data_rptr[4]));
Q_FDP4EP \_zygsfis_get_config_data_rptr_REG[3] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n595), .Q(_zygsfis_get_config_data_rptr[3]));
Q_FDP4EP \_zygsfis_get_config_data_rptr_REG[2] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n594), .Q(_zygsfis_get_config_data_rptr[2]));
Q_FDP4EP \_zygsfis_get_config_data_rptr_REG[1] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n593), .Q(_zygsfis_get_config_data_rptr[1]));
Q_FDP4EP \_zygsfis_get_config_data_rptr_REG[0] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n592), .Q(_zygsfis_get_config_data_rptr[0]));
Q_FDP4EP \_zygsfis_get_config_data_space_REG[4] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n964), .Q(_zygsfis_get_config_data_space[4]));
Q_FDP4EP \_zygsfis_get_config_data_space_REG[3] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n962), .Q(_zygsfis_get_config_data_space[3]));
Q_FDP4EP \_zygsfis_get_config_data_space_REG[2] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n960), .Q(_zygsfis_get_config_data_space[2]));
Q_FDP4EP \_zygsfis_get_config_data_space_REG[1] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n958), .Q(_zygsfis_get_config_data_space[1]));
Q_FDP4EP \_zygsfis_get_config_data_space_REG[0] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n956), .Q(_zygsfis_get_config_data_space[0]));
Q_FDP4EP \_zyGfifoF0_L324_s3_len_1_REG[11] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n1750), .Q(_zyGfifoF0_L324_s3_len_1[11]));
Q_FDP4EP \_zyGfifoF0_L324_s3_len_1_REG[10] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n1750), .Q(_zyGfifoF0_L324_s3_len_1[10]));
Q_FDP4EP \_zyGfifoF0_L324_s3_len_1_REG[9] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n1750), .Q(_zyGfifoF0_L324_s3_len_1[9]));
Q_FDP4EP \_zyGfifoF0_L324_s3_len_1_REG[8] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n1750), .Q(_zyGfifoF0_L324_s3_len_1[8]));
Q_FDP4EP \_zyGfifoF0_L324_s3_len_1_REG[7] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n1750), .Q(_zyGfifoF0_L324_s3_len_1[7]));
Q_FDP4EP \_zyGfifoF0_L324_s3_len_1_REG[6] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n1750), .Q(_zyGfifoF0_L324_s3_len_1[6]));
Q_FDP4EP \_zyGfifoF0_L324_s3_len_1_REG[5] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n1750), .Q(_zyGfifoF0_L324_s3_len_1[5]));
Q_FDP4EP \_zyGfifoF0_L324_s3_len_1_REG[4] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n1750), .Q(_zyGfifoF0_L324_s3_len_1[4]));
Q_FDP4EP \_zyGfifoF0_L324_s3_len_1_REG[3] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n1750), .Q(_zyGfifoF0_L324_s3_len_1[3]));
Q_FDP4EP \_zyGfifoF0_L324_s3_len_1_REG[2] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n1750), .Q(_zyGfifoF0_L324_s3_len_1[2]));
Q_FDP4EP \_zyGfifoF0_L324_s3_len_1_REG[1] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(_zyM2L324_pbcFsm0_s[0]), .Q(_zyGfifoF0_L324_s3_len_1[1]));
Q_FDP4EP \_zyGfifoF0_L324_s3_len_1_REG[0] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1138), .R(n1750), .D(n5382), .Q(_zyGfifoF0_L324_s3_len_1[0]));
Q_FDP4EP \_zyGfifoF2_L324_s2_len_3_REG[11] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n1750), .Q(_zyGfifoF2_L324_s2_len_3[11]));
Q_FDP4EP \_zyGfifoF2_L324_s2_len_3_REG[10] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n1750), .Q(_zyGfifoF2_L324_s2_len_3[10]));
Q_FDP4EP \_zyGfifoF2_L324_s2_len_3_REG[9] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n1750), .Q(_zyGfifoF2_L324_s2_len_3[9]));
Q_FDP4EP \_zyGfifoF2_L324_s2_len_3_REG[8] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n1750), .Q(_zyGfifoF2_L324_s2_len_3[8]));
Q_FDP4EP \_zyGfifoF2_L324_s2_len_3_REG[7] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n1750), .Q(_zyGfifoF2_L324_s2_len_3[7]));
Q_FDP4EP \_zyGfifoF2_L324_s2_len_3_REG[6] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n1750), .Q(_zyGfifoF2_L324_s2_len_3[6]));
Q_FDP4EP \_zyGfifoF2_L324_s2_len_3_REG[5] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n1750), .Q(_zyGfifoF2_L324_s2_len_3[5]));
Q_FDP4EP \_zyGfifoF2_L324_s2_len_3_REG[4] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n1750), .Q(_zyGfifoF2_L324_s2_len_3[4]));
Q_FDP4EP \_zyGfifoF2_L324_s2_len_3_REG[3] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n1750), .Q(_zyGfifoF2_L324_s2_len_3[3]));
Q_FDP4EP \_zyGfifoF2_L324_s2_len_3_REG[2] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n1750), .Q(_zyGfifoF2_L324_s2_len_3[2]));
Q_FDP4EP \_zyGfifoF2_L324_s2_len_3_REG[1] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n5382), .Q(_zyGfifoF2_L324_s2_len_3[1]));
Q_FDP4EP \_zyGfifoF2_L324_s2_len_3_REG[0] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1139), .R(n1750), .D(n1130), .Q(_zyGfifoF2_L324_s2_len_3[0]));
Q_INV U6299 ( .A(n1035), .Z(n45));
Q_FDP4EP _zyM2L324_pbcCapEn0_REG  ( .CK(_zyM2L324_pbcMevClk4), .CE(n45), .R(n1750), .D(n1131), .Q(_zyM2L324_pbcCapEn0));
Q_INV U6301 ( .A(n1038), .Z(n44));
Q_FDP4EP _zyM2L333_pbcCapEn1_REG  ( .CK(_zyM2L324_pbcMevClk4), .CE(n44), .R(n1750), .D(n1130), .Q(_zyM2L333_pbcCapEn1));
Q_INV U6303 ( .A(n1040), .Z(n43));
Q_FDP4EP _zyM2L349_pbcCapEn2_REG  ( .CK(_zyM2L324_pbcMevClk4), .CE(n43), .R(n1750), .D(n1129), .Q(_zyM2L349_pbcCapEn2));
Q_INV U6305 ( .A(n1048), .Z(n42));
Q_FDP4EP _zyM2L355_pbcCapEn3_REG  ( .CK(_zyM2L324_pbcMevClk4), .CE(n42), .R(n1750), .D(n1002), .Q(_zyM2L355_pbcCapEn3));
Q_FDP4EP \_zyM2L324_pbcFsm0_s_REG[1] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1140), .R(n1750), .D(n1128), .Q(_zyM2L324_pbcFsm0_s[1]));
Q_INV U6308 ( .A(_zyM2L324_pbcFsm0_s[1]), .Z(n1129));
Q_FDP4EP \_zyM2L324_pbcFsm0_s_REG[0] ( .CK(_zyM2L324_pbcMevClk4), .CE(n1140), .R(n1750), .D(n1127), .Q(_zyM2L324_pbcFsm0_s[0]));
Q_INV U6310 ( .A(_zyM2L324_pbcFsm0_s[0]), .Z(n1130));
Q_INV U6311 ( .A(n1036), .Z(n41));
Q_FDP4EP _zyM2L324_pbcEn13_REG  ( .CK(_zyM2L324_pbcMevClk4), .CE(n41), .R(n1750), .D(n1125), .Q(_zyM2L324_pbcEn13));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[0] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1123), .Q(_zyxr_L206_tfiV3_M2_pbcG3[0]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[31] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[31]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[30] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[30]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[29] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[29]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[28] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[28]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[27] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[27]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[26] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[26]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[25] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[25]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[24] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[24]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[23] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[23]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[22] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[22]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[21] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[21]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[20] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[20]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[19] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[19]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[18] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[18]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[17] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[17]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[16] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[16]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[15] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[15]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[14] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[14]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[13] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[13]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[12] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[12]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[11] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[11]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[10] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[10]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[9] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[9]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[8] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[8]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[7] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[7]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[6] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[6]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[5] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[5]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[4] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[4]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[3] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[3]));
Q_FDP4EP \_zyxr_L206_tfiV3_M2_pbcG3_REG[2] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyxr_L206_tfiV3_M2_pbcG3[2]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[31] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n996), .Q(_zyGfifoF1_L324_s2_data_2[31]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[30] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n995), .Q(_zyGfifoF1_L324_s2_data_2[30]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[29] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n994), .Q(_zyGfifoF1_L324_s2_data_2[29]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[28] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n993), .Q(_zyGfifoF1_L324_s2_data_2[28]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[27] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n992), .Q(_zyGfifoF1_L324_s2_data_2[27]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[26] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n991), .Q(_zyGfifoF1_L324_s2_data_2[26]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[25] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n990), .Q(_zyGfifoF1_L324_s2_data_2[25]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[24] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n989), .Q(_zyGfifoF1_L324_s2_data_2[24]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[23] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n988), .Q(_zyGfifoF1_L324_s2_data_2[23]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[22] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n987), .Q(_zyGfifoF1_L324_s2_data_2[22]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[21] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n986), .Q(_zyGfifoF1_L324_s2_data_2[21]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[20] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n985), .Q(_zyGfifoF1_L324_s2_data_2[20]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[19] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n984), .Q(_zyGfifoF1_L324_s2_data_2[19]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[18] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n983), .Q(_zyGfifoF1_L324_s2_data_2[18]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[17] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n982), .Q(_zyGfifoF1_L324_s2_data_2[17]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[16] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n981), .Q(_zyGfifoF1_L324_s2_data_2[16]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[15] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n980), .Q(_zyGfifoF1_L324_s2_data_2[15]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[14] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n979), .Q(_zyGfifoF1_L324_s2_data_2[14]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[13] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n978), .Q(_zyGfifoF1_L324_s2_data_2[13]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[12] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n977), .Q(_zyGfifoF1_L324_s2_data_2[12]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[11] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n976), .Q(_zyGfifoF1_L324_s2_data_2[11]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[10] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n975), .Q(_zyGfifoF1_L324_s2_data_2[10]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[9] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n974), .Q(_zyGfifoF1_L324_s2_data_2[9]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[8] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n973), .Q(_zyGfifoF1_L324_s2_data_2[8]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[7] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n972), .Q(_zyGfifoF1_L324_s2_data_2[7]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[6] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n971), .Q(_zyGfifoF1_L324_s2_data_2[6]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[5] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n970), .Q(_zyGfifoF1_L324_s2_data_2[5]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[4] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n969), .Q(_zyGfifoF1_L324_s2_data_2[4]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[3] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n968), .Q(_zyGfifoF1_L324_s2_data_2[3]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[2] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n967), .Q(_zyGfifoF1_L324_s2_data_2[2]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[1] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n966), .Q(_zyGfifoF1_L324_s2_data_2[1]));
Q_FDP4EP \_zyGfifoF1_L324_s2_data_2_REG[0] ( .CK(_zyM2L324_pbcMevClk4), .CE(n48), .R(n1750), .D(n965), .Q(_zyGfifoF1_L324_s2_data_2[0]));
Q_FDP4EP \_zyL326_tfiRv17_REG[31] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[31]));
Q_FDP4EP \_zyL326_tfiRv17_REG[30] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[30]));
Q_FDP4EP \_zyL326_tfiRv17_REG[29] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[29]));
Q_FDP4EP \_zyL326_tfiRv17_REG[28] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[28]));
Q_FDP4EP \_zyL326_tfiRv17_REG[27] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[27]));
Q_FDP4EP \_zyL326_tfiRv17_REG[26] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[26]));
Q_FDP4EP \_zyL326_tfiRv17_REG[25] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[25]));
Q_FDP4EP \_zyL326_tfiRv17_REG[24] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[24]));
Q_FDP4EP \_zyL326_tfiRv17_REG[23] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[23]));
Q_FDP4EP \_zyL326_tfiRv17_REG[22] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[22]));
Q_FDP4EP \_zyL326_tfiRv17_REG[21] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[21]));
Q_FDP4EP \_zyL326_tfiRv17_REG[20] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[20]));
Q_FDP4EP \_zyL326_tfiRv17_REG[19] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[19]));
Q_FDP4EP \_zyL326_tfiRv17_REG[18] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[18]));
Q_FDP4EP \_zyL326_tfiRv17_REG[17] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[17]));
Q_FDP4EP \_zyL326_tfiRv17_REG[16] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[16]));
Q_FDP4EP \_zyL326_tfiRv17_REG[15] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[15]));
Q_FDP4EP \_zyL326_tfiRv17_REG[14] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[14]));
Q_FDP4EP \_zyL326_tfiRv17_REG[13] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[13]));
Q_FDP4EP \_zyL326_tfiRv17_REG[12] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[12]));
Q_FDP4EP \_zyL326_tfiRv17_REG[11] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[11]));
Q_FDP4EP \_zyL326_tfiRv17_REG[10] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[10]));
Q_FDP4EP \_zyL326_tfiRv17_REG[9] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[9]));
Q_FDP4EP \_zyL326_tfiRv17_REG[8] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[8]));
Q_FDP4EP \_zyL326_tfiRv17_REG[7] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[7]));
Q_FDP4EP \_zyL326_tfiRv17_REG[6] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[6]));
Q_FDP4EP \_zyL326_tfiRv17_REG[5] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[5]));
Q_FDP4EP \_zyL326_tfiRv17_REG[4] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[4]));
Q_FDP4EP \_zyL326_tfiRv17_REG[3] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[3]));
Q_FDP4EP \_zyL326_tfiRv17_REG[2] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(_zyL326_tfiRv17[2]));
Q_FDP4EP \_zyL326_tfiRv17_REG[1] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1133), .Q(_zyL326_tfiRv17[1]));
Q_FDP4EP \_zyL326_tfiRv17_REG[0] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1123), .Q(_zyL326_tfiRv17[0]));
Q_FDP4EP \retval_REG[31] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[31]));
Q_FDP4EP \retval_REG[30] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[30]));
Q_FDP4EP \retval_REG[29] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[29]));
Q_FDP4EP \retval_REG[28] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[28]));
Q_FDP4EP \retval_REG[27] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[27]));
Q_FDP4EP \retval_REG[26] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[26]));
Q_FDP4EP \retval_REG[25] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[25]));
Q_FDP4EP \retval_REG[24] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[24]));
Q_FDP4EP \retval_REG[23] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[23]));
Q_FDP4EP \retval_REG[22] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[22]));
Q_FDP4EP \retval_REG[21] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[21]));
Q_FDP4EP \retval_REG[20] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[20]));
Q_FDP4EP \retval_REG[19] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[19]));
Q_FDP4EP \retval_REG[18] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[18]));
Q_FDP4EP \retval_REG[17] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[17]));
Q_FDP4EP \retval_REG[16] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[16]));
Q_FDP4EP \retval_REG[15] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[15]));
Q_FDP4EP \retval_REG[14] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[14]));
Q_FDP4EP \retval_REG[13] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[13]));
Q_FDP4EP \retval_REG[12] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[12]));
Q_FDP4EP \retval_REG[11] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[11]));
Q_FDP4EP \retval_REG[10] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[10]));
Q_FDP4EP \retval_REG[9] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[9]));
Q_FDP4EP \retval_REG[8] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[8]));
Q_FDP4EP \retval_REG[7] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[7]));
Q_FDP4EP \retval_REG[6] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[6]));
Q_FDP4EP \retval_REG[5] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[5]));
Q_FDP4EP \retval_REG[4] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[4]));
Q_FDP4EP \retval_REG[3] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[3]));
Q_FDP4EP \retval_REG[2] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1750), .Q(retval[2]));
Q_FDP4EP \retval_REG[1] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1133), .Q(retval[1]));
Q_FDP4EP \retval_REG[0] ( .CK(_zyM2L324_pbcMevClk4), .CE(n47), .R(n1750), .D(n1123), .Q(retval[0]));
Q_FDP4EP _zzM2L368_mdxP3_En_REG  ( .CK(clk), .CE(n1635), .R(n1750), .D(_zzM2L368_mdxP3_EnNxt), .Q(_zzM2L368_mdxP3_En));
Q_FDP4EP _zzM2L368_mdxP3_kme_ib_tvalid_wr0_REG  ( .CK(clk), .CE(n1635), .R(n1750), .D(n5382), .Q(_zzM2L368_mdxP3_kme_ib_tvalid_wr0));
Q_INV U6442 ( .A(_zygsfis_ib_service_data_req[4]), .Z(n40));
Q_FDP4EP \_zygsfis_ib_service_data_req_REG[4] ( .CK(clk), .CE(n5881), .R(n1750), .D(n40), .Q(_zygsfis_ib_service_data_req[4]));
Q_FDP4EP \_zygsfis_ib_service_data_req_REG[3] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1255), .Q(_zygsfis_ib_service_data_req[3]));
Q_FDP4EP \_zygsfis_ib_service_data_req_REG[2] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1253), .Q(_zygsfis_ib_service_data_req[2]));
Q_FDP4EP \_zygsfis_ib_service_data_req_REG[1] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1251), .Q(_zygsfis_ib_service_data_req[1]));
Q_INV U6447 ( .A(_zygsfis_ib_service_data_req[0]), .Z(n39));
Q_FDP4EP \_zygsfis_ib_service_data_req_REG[0] ( .CK(clk), .CE(n1641), .R(n1750), .D(n39), .Q(_zygsfis_ib_service_data_req[0]));
Q_FDP4EP _zyGfifoF11_L207_req_0_REG  ( .CK(clk), .CE(n1641), .R(n1750), .D(n1165), .Q(_zyGfifoF11_L207_req_0));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[31] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1750), .Q(_zyGfifoF11_L207_data_0[31]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[30] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1750), .Q(_zyGfifoF11_L207_data_0[30]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[29] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1750), .Q(_zyGfifoF11_L207_data_0[29]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[28] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1750), .Q(_zyGfifoF11_L207_data_0[28]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[27] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1750), .Q(_zyGfifoF11_L207_data_0[27]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[26] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1750), .Q(_zyGfifoF11_L207_data_0[26]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[25] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1750), .Q(_zyGfifoF11_L207_data_0[25]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[24] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1750), .Q(_zyGfifoF11_L207_data_0[24]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[23] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1750), .Q(_zyGfifoF11_L207_data_0[23]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[22] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1750), .Q(_zyGfifoF11_L207_data_0[22]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[21] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1750), .Q(_zyGfifoF11_L207_data_0[21]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[20] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1750), .Q(_zyGfifoF11_L207_data_0[20]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[19] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1750), .Q(_zyGfifoF11_L207_data_0[19]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[18] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1750), .Q(_zyGfifoF11_L207_data_0[18]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[17] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1750), .Q(_zyGfifoF11_L207_data_0[17]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[16] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1750), .Q(_zyGfifoF11_L207_data_0[16]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[15] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1750), .Q(_zyGfifoF11_L207_data_0[15]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[14] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1750), .Q(_zyGfifoF11_L207_data_0[14]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[13] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1750), .Q(_zyGfifoF11_L207_data_0[13]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[12] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1750), .Q(_zyGfifoF11_L207_data_0[12]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[11] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1750), .Q(_zyGfifoF11_L207_data_0[11]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[10] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1750), .Q(_zyGfifoF11_L207_data_0[10]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[9] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1750), .Q(_zyGfifoF11_L207_data_0[9]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[8] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1750), .Q(_zyGfifoF11_L207_data_0[8]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[7] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1750), .Q(_zyGfifoF11_L207_data_0[7]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[6] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1750), .Q(_zyGfifoF11_L207_data_0[6]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[5] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1750), .Q(_zyGfifoF11_L207_data_0[5]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[4] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1304), .Q(_zyGfifoF11_L207_data_0[4]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[3] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1303), .Q(_zyGfifoF11_L207_data_0[3]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[2] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1302), .Q(_zyGfifoF11_L207_data_0[2]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[1] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1301), .Q(_zyGfifoF11_L207_data_0[1]));
Q_FDP4EP \_zyGfifoF11_L207_data_0_REG[0] ( .CK(clk), .CE(n1641), .R(n1750), .D(n1300), .Q(_zyGfifoF11_L207_data_0[0]));
Q_INV U6482 ( .A(n1485), .Z(n38));
Q_FDP4EP _zyGfifoF0_L368_s2_req_4_REG  ( .CK(clk), .CE(n38), .R(n1750), .D(n1455), .Q(_zyGfifoF0_L368_s2_req_4));
Q_FDP4EP \_zyGfifoF0_L368_s2_cbid_4_REG[19] ( .CK(clk), .CE(n38), .R(n1750), .D(n1454), .Q(_zyGfifoF0_L368_s2_cbid_4[19]));
Q_FDP4EP \_zyGfifoF0_L368_s2_cbid_4_REG[18] ( .CK(clk), .CE(n38), .R(n1750), .D(n1453), .Q(_zyGfifoF0_L368_s2_cbid_4[18]));
Q_FDP4EP \_zyGfifoF0_L368_s2_cbid_4_REG[17] ( .CK(clk), .CE(n38), .R(n1750), .D(n1452), .Q(_zyGfifoF0_L368_s2_cbid_4[17]));
Q_FDP4EP \_zyGfifoF0_L368_s2_cbid_4_REG[16] ( .CK(clk), .CE(n38), .R(n1750), .D(n1451), .Q(_zyGfifoF0_L368_s2_cbid_4[16]));
Q_FDP4EP \_zyGfifoF0_L368_s2_cbid_4_REG[15] ( .CK(clk), .CE(n38), .R(n1750), .D(n1450), .Q(_zyGfifoF0_L368_s2_cbid_4[15]));
Q_FDP4EP \_zyGfifoF0_L368_s2_cbid_4_REG[14] ( .CK(clk), .CE(n38), .R(n1750), .D(n1449), .Q(_zyGfifoF0_L368_s2_cbid_4[14]));
Q_FDP4EP \_zyGfifoF0_L368_s2_cbid_4_REG[13] ( .CK(clk), .CE(n38), .R(n1750), .D(n1448), .Q(_zyGfifoF0_L368_s2_cbid_4[13]));
Q_FDP4EP \_zyGfifoF0_L368_s2_cbid_4_REG[12] ( .CK(clk), .CE(n38), .R(n1750), .D(n1447), .Q(_zyGfifoF0_L368_s2_cbid_4[12]));
Q_FDP4EP \_zyGfifoF0_L368_s2_cbid_4_REG[11] ( .CK(clk), .CE(n38), .R(n1750), .D(n1446), .Q(_zyGfifoF0_L368_s2_cbid_4[11]));
Q_FDP4EP \_zyGfifoF0_L368_s2_cbid_4_REG[10] ( .CK(clk), .CE(n38), .R(n1750), .D(n1445), .Q(_zyGfifoF0_L368_s2_cbid_4[10]));
Q_FDP4EP \_zyGfifoF0_L368_s2_cbid_4_REG[9] ( .CK(clk), .CE(n38), .R(n1750), .D(n1444), .Q(_zyGfifoF0_L368_s2_cbid_4[9]));
Q_FDP4EP \_zyGfifoF0_L368_s2_cbid_4_REG[8] ( .CK(clk), .CE(n38), .R(n1750), .D(n1443), .Q(_zyGfifoF0_L368_s2_cbid_4[8]));
Q_FDP4EP \_zyGfifoF0_L368_s2_cbid_4_REG[7] ( .CK(clk), .CE(n38), .R(n1750), .D(n1442), .Q(_zyGfifoF0_L368_s2_cbid_4[7]));
Q_FDP4EP \_zyGfifoF0_L368_s2_cbid_4_REG[6] ( .CK(clk), .CE(n38), .R(n1750), .D(n1441), .Q(_zyGfifoF0_L368_s2_cbid_4[6]));
Q_FDP4EP \_zyGfifoF0_L368_s2_cbid_4_REG[5] ( .CK(clk), .CE(n38), .R(n1750), .D(n1440), .Q(_zyGfifoF0_L368_s2_cbid_4[5]));
Q_FDP4EP \_zyGfifoF0_L368_s2_cbid_4_REG[4] ( .CK(clk), .CE(n38), .R(n1750), .D(n1439), .Q(_zyGfifoF0_L368_s2_cbid_4[4]));
Q_FDP4EP \_zyGfifoF0_L368_s2_cbid_4_REG[3] ( .CK(clk), .CE(n38), .R(n1750), .D(n1438), .Q(_zyGfifoF0_L368_s2_cbid_4[3]));
Q_FDP4EP \_zyGfifoF0_L368_s2_cbid_4_REG[2] ( .CK(clk), .CE(n38), .R(n1750), .D(n1437), .Q(_zyGfifoF0_L368_s2_cbid_4[2]));
Q_FDP4EP \_zyGfifoF0_L368_s2_cbid_4_REG[1] ( .CK(clk), .CE(n38), .R(n1750), .D(n1436), .Q(_zyGfifoF0_L368_s2_cbid_4[1]));
Q_FDP4EP \_zyGfifoF0_L368_s2_cbid_4_REG[0] ( .CK(clk), .CE(n38), .R(n1750), .D(n1435), .Q(_zyGfifoF0_L368_s2_cbid_4[0]));
Q_INV U6504 ( .A(n1484), .Z(n37));
Q_FDP4EP _zyGfifoF14_L373_req_0_REG  ( .CK(clk), .CE(n37), .R(n1750), .D(n1167), .Q(_zyGfifoF14_L373_req_0));
Q_FDP4EP _zyGfifoF15_L375_req_0_REG  ( .CK(clk), .CE(n1638), .R(n1750), .D(n1168), .Q(_zyGfifoF15_L375_req_0));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[135] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1708), .Q(_zyGfifoF15_L375_data_0[135]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[134] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1707), .Q(_zyGfifoF15_L375_data_0[134]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[133] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1706), .Q(_zyGfifoF15_L375_data_0[133]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[132] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1705), .Q(_zyGfifoF15_L375_data_0[132]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[131] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1704), .Q(_zyGfifoF15_L375_data_0[131]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[130] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1703), .Q(_zyGfifoF15_L375_data_0[130]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[129] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1702), .Q(_zyGfifoF15_L375_data_0[129]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[128] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1701), .Q(_zyGfifoF15_L375_data_0[128]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[127] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1700), .Q(_zyGfifoF15_L375_data_0[127]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[126] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1699), .Q(_zyGfifoF15_L375_data_0[126]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[125] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1698), .Q(_zyGfifoF15_L375_data_0[125]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[124] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1697), .Q(_zyGfifoF15_L375_data_0[124]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[123] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1696), .Q(_zyGfifoF15_L375_data_0[123]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[122] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1695), .Q(_zyGfifoF15_L375_data_0[122]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[121] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1694), .Q(_zyGfifoF15_L375_data_0[121]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[120] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1693), .Q(_zyGfifoF15_L375_data_0[120]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[119] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1692), .Q(_zyGfifoF15_L375_data_0[119]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[118] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1691), .Q(_zyGfifoF15_L375_data_0[118]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[117] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1690), .Q(_zyGfifoF15_L375_data_0[117]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[116] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1689), .Q(_zyGfifoF15_L375_data_0[116]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[115] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1688), .Q(_zyGfifoF15_L375_data_0[115]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[114] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1687), .Q(_zyGfifoF15_L375_data_0[114]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[113] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1686), .Q(_zyGfifoF15_L375_data_0[113]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[112] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1685), .Q(_zyGfifoF15_L375_data_0[112]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[111] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1684), .Q(_zyGfifoF15_L375_data_0[111]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[110] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1683), .Q(_zyGfifoF15_L375_data_0[110]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[109] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1682), .Q(_zyGfifoF15_L375_data_0[109]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[108] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1681), .Q(_zyGfifoF15_L375_data_0[108]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[107] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1680), .Q(_zyGfifoF15_L375_data_0[107]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[106] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1679), .Q(_zyGfifoF15_L375_data_0[106]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[105] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1678), .Q(_zyGfifoF15_L375_data_0[105]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[104] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1677), .Q(_zyGfifoF15_L375_data_0[104]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[103] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1676), .Q(_zyGfifoF15_L375_data_0[103]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[102] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1675), .Q(_zyGfifoF15_L375_data_0[102]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[101] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1674), .Q(_zyGfifoF15_L375_data_0[101]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[100] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1673), .Q(_zyGfifoF15_L375_data_0[100]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[99] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1672), .Q(_zyGfifoF15_L375_data_0[99]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[98] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1671), .Q(_zyGfifoF15_L375_data_0[98]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[97] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1670), .Q(_zyGfifoF15_L375_data_0[97]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[96] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1669), .Q(_zyGfifoF15_L375_data_0[96]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[95] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1668), .Q(_zyGfifoF15_L375_data_0[95]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[94] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1667), .Q(_zyGfifoF15_L375_data_0[94]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[93] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1666), .Q(_zyGfifoF15_L375_data_0[93]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[92] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1665), .Q(_zyGfifoF15_L375_data_0[92]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[91] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1664), .Q(_zyGfifoF15_L375_data_0[91]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[90] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1663), .Q(_zyGfifoF15_L375_data_0[90]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[89] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1662), .Q(_zyGfifoF15_L375_data_0[89]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[88] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1661), .Q(_zyGfifoF15_L375_data_0[88]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[87] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1660), .Q(_zyGfifoF15_L375_data_0[87]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[86] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1659), .Q(_zyGfifoF15_L375_data_0[86]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[85] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1658), .Q(_zyGfifoF15_L375_data_0[85]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[84] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1657), .Q(_zyGfifoF15_L375_data_0[84]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[83] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1656), .Q(_zyGfifoF15_L375_data_0[83]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[82] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1655), .Q(_zyGfifoF15_L375_data_0[82]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[81] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1654), .Q(_zyGfifoF15_L375_data_0[81]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[80] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1653), .Q(_zyGfifoF15_L375_data_0[80]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[79] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1652), .Q(_zyGfifoF15_L375_data_0[79]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[78] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1651), .Q(_zyGfifoF15_L375_data_0[78]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[77] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1650), .Q(_zyGfifoF15_L375_data_0[77]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[76] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1649), .Q(_zyGfifoF15_L375_data_0[76]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[75] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1648), .Q(_zyGfifoF15_L375_data_0[75]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[74] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1647), .Q(_zyGfifoF15_L375_data_0[74]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[73] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1646), .Q(_zyGfifoF15_L375_data_0[73]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[72] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1645), .Q(_zyGfifoF15_L375_data_0[72]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[71] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1352), .Q(_zyGfifoF15_L375_data_0[71]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[70] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1351), .Q(_zyGfifoF15_L375_data_0[70]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[69] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1350), .Q(_zyGfifoF15_L375_data_0[69]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[68] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1349), .Q(_zyGfifoF15_L375_data_0[68]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[67] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1348), .Q(_zyGfifoF15_L375_data_0[67]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[66] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1347), .Q(_zyGfifoF15_L375_data_0[66]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[65] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1346), .Q(_zyGfifoF15_L375_data_0[65]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[64] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1345), .Q(_zyGfifoF15_L375_data_0[64]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[63] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1344), .Q(_zyGfifoF15_L375_data_0[63]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[62] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1343), .Q(_zyGfifoF15_L375_data_0[62]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[61] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1342), .Q(_zyGfifoF15_L375_data_0[61]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[60] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1341), .Q(_zyGfifoF15_L375_data_0[60]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[59] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1340), .Q(_zyGfifoF15_L375_data_0[59]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[58] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1339), .Q(_zyGfifoF15_L375_data_0[58]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[57] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1338), .Q(_zyGfifoF15_L375_data_0[57]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[56] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1337), .Q(_zyGfifoF15_L375_data_0[56]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[55] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1336), .Q(_zyGfifoF15_L375_data_0[55]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[54] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1335), .Q(_zyGfifoF15_L375_data_0[54]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[53] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1334), .Q(_zyGfifoF15_L375_data_0[53]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[52] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1333), .Q(_zyGfifoF15_L375_data_0[52]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[51] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1332), .Q(_zyGfifoF15_L375_data_0[51]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[50] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1331), .Q(_zyGfifoF15_L375_data_0[50]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[49] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1330), .Q(_zyGfifoF15_L375_data_0[49]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[48] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1329), .Q(_zyGfifoF15_L375_data_0[48]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[47] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1328), .Q(_zyGfifoF15_L375_data_0[47]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[46] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1327), .Q(_zyGfifoF15_L375_data_0[46]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[45] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1326), .Q(_zyGfifoF15_L375_data_0[45]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[44] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1325), .Q(_zyGfifoF15_L375_data_0[44]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[43] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1324), .Q(_zyGfifoF15_L375_data_0[43]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[42] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1323), .Q(_zyGfifoF15_L375_data_0[42]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[41] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1322), .Q(_zyGfifoF15_L375_data_0[41]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[40] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1321), .Q(_zyGfifoF15_L375_data_0[40]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[39] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1382), .Q(_zyGfifoF15_L375_data_0[39]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[38] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1381), .Q(_zyGfifoF15_L375_data_0[38]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[37] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1380), .Q(_zyGfifoF15_L375_data_0[37]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[36] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1379), .Q(_zyGfifoF15_L375_data_0[36]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[35] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1378), .Q(_zyGfifoF15_L375_data_0[35]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[34] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1377), .Q(_zyGfifoF15_L375_data_0[34]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[33] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1376), .Q(_zyGfifoF15_L375_data_0[33]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[32] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1375), .Q(_zyGfifoF15_L375_data_0[32]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[31] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1414), .Q(_zyGfifoF15_L375_data_0[31]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[30] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1413), .Q(_zyGfifoF15_L375_data_0[30]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[29] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1412), .Q(_zyGfifoF15_L375_data_0[29]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[28] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1411), .Q(_zyGfifoF15_L375_data_0[28]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[27] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1410), .Q(_zyGfifoF15_L375_data_0[27]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[26] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1409), .Q(_zyGfifoF15_L375_data_0[26]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[25] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1408), .Q(_zyGfifoF15_L375_data_0[25]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[24] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1407), .Q(_zyGfifoF15_L375_data_0[24]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[23] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1406), .Q(_zyGfifoF15_L375_data_0[23]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[22] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1405), .Q(_zyGfifoF15_L375_data_0[22]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[21] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1404), .Q(_zyGfifoF15_L375_data_0[21]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[20] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1403), .Q(_zyGfifoF15_L375_data_0[20]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[19] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1402), .Q(_zyGfifoF15_L375_data_0[19]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[18] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1401), .Q(_zyGfifoF15_L375_data_0[18]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[17] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1400), .Q(_zyGfifoF15_L375_data_0[17]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[16] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1399), .Q(_zyGfifoF15_L375_data_0[16]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[15] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1398), .Q(_zyGfifoF15_L375_data_0[15]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[14] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1397), .Q(_zyGfifoF15_L375_data_0[14]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[13] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1396), .Q(_zyGfifoF15_L375_data_0[13]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[12] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1395), .Q(_zyGfifoF15_L375_data_0[12]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[11] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1394), .Q(_zyGfifoF15_L375_data_0[11]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[10] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1393), .Q(_zyGfifoF15_L375_data_0[10]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[9] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1392), .Q(_zyGfifoF15_L375_data_0[9]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[8] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1391), .Q(_zyGfifoF15_L375_data_0[8]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[7] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1390), .Q(_zyGfifoF15_L375_data_0[7]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[6] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1389), .Q(_zyGfifoF15_L375_data_0[6]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[5] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1388), .Q(_zyGfifoF15_L375_data_0[5]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[4] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1387), .Q(_zyGfifoF15_L375_data_0[4]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[3] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1386), .Q(_zyGfifoF15_L375_data_0[3]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[2] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1385), .Q(_zyGfifoF15_L375_data_0[2]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[1] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1384), .Q(_zyGfifoF15_L375_data_0[1]));
Q_FDP4EP \_zyGfifoF15_L375_data_0_REG[0] ( .CK(clk), .CE(n1638), .R(n1750), .D(n1383), .Q(_zyGfifoF15_L375_data_0[0]));
Q_INV U6643 ( .A(n1488), .Z(n36));
Q_FDP4EP _zyGfifoF16_L381_req_0_REG  ( .CK(clk), .CE(n36), .R(n1750), .D(n1169), .Q(_zyGfifoF16_L381_req_0));
Q_INV U6645 ( .A(n1489), .Z(n35));
Q_FDP4EP _zyGfifoF17_L390_req_0_REG  ( .CK(clk), .CE(n35), .R(n1750), .D(n1170), .Q(_zyGfifoF17_L390_req_0));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[63] ( .CK(clk), .CE(n35), .R(n1750), .D(n1708), .Q(_zyGfifoF17_L390_data_0[63]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[62] ( .CK(clk), .CE(n35), .R(n1750), .D(n1707), .Q(_zyGfifoF17_L390_data_0[62]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[61] ( .CK(clk), .CE(n35), .R(n1750), .D(n1706), .Q(_zyGfifoF17_L390_data_0[61]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[60] ( .CK(clk), .CE(n35), .R(n1750), .D(n1705), .Q(_zyGfifoF17_L390_data_0[60]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[59] ( .CK(clk), .CE(n35), .R(n1750), .D(n1704), .Q(_zyGfifoF17_L390_data_0[59]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[58] ( .CK(clk), .CE(n35), .R(n1750), .D(n1703), .Q(_zyGfifoF17_L390_data_0[58]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[57] ( .CK(clk), .CE(n35), .R(n1750), .D(n1702), .Q(_zyGfifoF17_L390_data_0[57]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[56] ( .CK(clk), .CE(n35), .R(n1750), .D(n1701), .Q(_zyGfifoF17_L390_data_0[56]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[55] ( .CK(clk), .CE(n35), .R(n1750), .D(n1700), .Q(_zyGfifoF17_L390_data_0[55]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[54] ( .CK(clk), .CE(n35), .R(n1750), .D(n1699), .Q(_zyGfifoF17_L390_data_0[54]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[53] ( .CK(clk), .CE(n35), .R(n1750), .D(n1698), .Q(_zyGfifoF17_L390_data_0[53]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[52] ( .CK(clk), .CE(n35), .R(n1750), .D(n1697), .Q(_zyGfifoF17_L390_data_0[52]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[51] ( .CK(clk), .CE(n35), .R(n1750), .D(n1696), .Q(_zyGfifoF17_L390_data_0[51]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[50] ( .CK(clk), .CE(n35), .R(n1750), .D(n1695), .Q(_zyGfifoF17_L390_data_0[50]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[49] ( .CK(clk), .CE(n35), .R(n1750), .D(n1694), .Q(_zyGfifoF17_L390_data_0[49]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[48] ( .CK(clk), .CE(n35), .R(n1750), .D(n1693), .Q(_zyGfifoF17_L390_data_0[48]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[47] ( .CK(clk), .CE(n35), .R(n1750), .D(n1692), .Q(_zyGfifoF17_L390_data_0[47]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[46] ( .CK(clk), .CE(n35), .R(n1750), .D(n1691), .Q(_zyGfifoF17_L390_data_0[46]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[45] ( .CK(clk), .CE(n35), .R(n1750), .D(n1690), .Q(_zyGfifoF17_L390_data_0[45]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[44] ( .CK(clk), .CE(n35), .R(n1750), .D(n1689), .Q(_zyGfifoF17_L390_data_0[44]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[43] ( .CK(clk), .CE(n35), .R(n1750), .D(n1688), .Q(_zyGfifoF17_L390_data_0[43]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[42] ( .CK(clk), .CE(n35), .R(n1750), .D(n1687), .Q(_zyGfifoF17_L390_data_0[42]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[41] ( .CK(clk), .CE(n35), .R(n1750), .D(n1686), .Q(_zyGfifoF17_L390_data_0[41]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[40] ( .CK(clk), .CE(n35), .R(n1750), .D(n1685), .Q(_zyGfifoF17_L390_data_0[40]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[39] ( .CK(clk), .CE(n35), .R(n1750), .D(n1684), .Q(_zyGfifoF17_L390_data_0[39]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[38] ( .CK(clk), .CE(n35), .R(n1750), .D(n1683), .Q(_zyGfifoF17_L390_data_0[38]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[37] ( .CK(clk), .CE(n35), .R(n1750), .D(n1682), .Q(_zyGfifoF17_L390_data_0[37]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[36] ( .CK(clk), .CE(n35), .R(n1750), .D(n1681), .Q(_zyGfifoF17_L390_data_0[36]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[35] ( .CK(clk), .CE(n35), .R(n1750), .D(n1680), .Q(_zyGfifoF17_L390_data_0[35]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[34] ( .CK(clk), .CE(n35), .R(n1750), .D(n1679), .Q(_zyGfifoF17_L390_data_0[34]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[33] ( .CK(clk), .CE(n35), .R(n1750), .D(n1678), .Q(_zyGfifoF17_L390_data_0[33]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[32] ( .CK(clk), .CE(n35), .R(n1750), .D(n1677), .Q(_zyGfifoF17_L390_data_0[32]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[31] ( .CK(clk), .CE(n35), .R(n1750), .D(n1676), .Q(_zyGfifoF17_L390_data_0[31]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[30] ( .CK(clk), .CE(n35), .R(n1750), .D(n1675), .Q(_zyGfifoF17_L390_data_0[30]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[29] ( .CK(clk), .CE(n35), .R(n1750), .D(n1674), .Q(_zyGfifoF17_L390_data_0[29]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[28] ( .CK(clk), .CE(n35), .R(n1750), .D(n1673), .Q(_zyGfifoF17_L390_data_0[28]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[27] ( .CK(clk), .CE(n35), .R(n1750), .D(n1672), .Q(_zyGfifoF17_L390_data_0[27]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[26] ( .CK(clk), .CE(n35), .R(n1750), .D(n1671), .Q(_zyGfifoF17_L390_data_0[26]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[25] ( .CK(clk), .CE(n35), .R(n1750), .D(n1670), .Q(_zyGfifoF17_L390_data_0[25]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[24] ( .CK(clk), .CE(n35), .R(n1750), .D(n1669), .Q(_zyGfifoF17_L390_data_0[24]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[23] ( .CK(clk), .CE(n35), .R(n1750), .D(n1668), .Q(_zyGfifoF17_L390_data_0[23]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[22] ( .CK(clk), .CE(n35), .R(n1750), .D(n1667), .Q(_zyGfifoF17_L390_data_0[22]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[21] ( .CK(clk), .CE(n35), .R(n1750), .D(n1666), .Q(_zyGfifoF17_L390_data_0[21]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[20] ( .CK(clk), .CE(n35), .R(n1750), .D(n1665), .Q(_zyGfifoF17_L390_data_0[20]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[19] ( .CK(clk), .CE(n35), .R(n1750), .D(n1664), .Q(_zyGfifoF17_L390_data_0[19]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[18] ( .CK(clk), .CE(n35), .R(n1750), .D(n1663), .Q(_zyGfifoF17_L390_data_0[18]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[17] ( .CK(clk), .CE(n35), .R(n1750), .D(n1662), .Q(_zyGfifoF17_L390_data_0[17]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[16] ( .CK(clk), .CE(n35), .R(n1750), .D(n1661), .Q(_zyGfifoF17_L390_data_0[16]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[15] ( .CK(clk), .CE(n35), .R(n1750), .D(n1660), .Q(_zyGfifoF17_L390_data_0[15]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[14] ( .CK(clk), .CE(n35), .R(n1750), .D(n1659), .Q(_zyGfifoF17_L390_data_0[14]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[13] ( .CK(clk), .CE(n35), .R(n1750), .D(n1658), .Q(_zyGfifoF17_L390_data_0[13]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[12] ( .CK(clk), .CE(n35), .R(n1750), .D(n1657), .Q(_zyGfifoF17_L390_data_0[12]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[11] ( .CK(clk), .CE(n35), .R(n1750), .D(n1656), .Q(_zyGfifoF17_L390_data_0[11]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[10] ( .CK(clk), .CE(n35), .R(n1750), .D(n1655), .Q(_zyGfifoF17_L390_data_0[10]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[9] ( .CK(clk), .CE(n35), .R(n1750), .D(n1654), .Q(_zyGfifoF17_L390_data_0[9]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[8] ( .CK(clk), .CE(n35), .R(n1750), .D(n1653), .Q(_zyGfifoF17_L390_data_0[8]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[7] ( .CK(clk), .CE(n35), .R(n1750), .D(n1652), .Q(_zyGfifoF17_L390_data_0[7]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[6] ( .CK(clk), .CE(n35), .R(n1750), .D(n1651), .Q(_zyGfifoF17_L390_data_0[6]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[5] ( .CK(clk), .CE(n35), .R(n1750), .D(n1650), .Q(_zyGfifoF17_L390_data_0[5]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[4] ( .CK(clk), .CE(n35), .R(n1750), .D(n1649), .Q(_zyGfifoF17_L390_data_0[4]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[3] ( .CK(clk), .CE(n35), .R(n1750), .D(n1648), .Q(_zyGfifoF17_L390_data_0[3]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[2] ( .CK(clk), .CE(n35), .R(n1750), .D(n1647), .Q(_zyGfifoF17_L390_data_0[2]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[1] ( .CK(clk), .CE(n35), .R(n1750), .D(n1646), .Q(_zyGfifoF17_L390_data_0[1]));
Q_FDP4EP \_zyGfifoF17_L390_data_0_REG[0] ( .CK(clk), .CE(n35), .R(n1750), .D(n1645), .Q(_zyGfifoF17_L390_data_0[0]));
Q_FDP4EP _zyGfifoF18_L530_req_0_REG  ( .CK(clk), .CE(n1640), .R(n1750), .D(n1171), .Q(_zyGfifoF18_L530_req_0));
Q_FDP4EP _zyGfifoF19_L412_req_0_REG  ( .CK(clk), .CE(n1635), .R(n1750), .D(n1172), .Q(_zyGfifoF19_L412_req_0));
Q_FDP4EP \_zyGfifoF19_L412_data_0_REG[7] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1382), .Q(_zyGfifoF19_L412_data_0[7]));
Q_FDP4EP \_zyGfifoF19_L412_data_0_REG[6] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1381), .Q(_zyGfifoF19_L412_data_0[6]));
Q_FDP4EP \_zyGfifoF19_L412_data_0_REG[5] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1380), .Q(_zyGfifoF19_L412_data_0[5]));
Q_FDP4EP \_zyGfifoF19_L412_data_0_REG[4] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1379), .Q(_zyGfifoF19_L412_data_0[4]));
Q_FDP4EP \_zyGfifoF19_L412_data_0_REG[3] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1378), .Q(_zyGfifoF19_L412_data_0[3]));
Q_FDP4EP \_zyGfifoF19_L412_data_0_REG[2] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1377), .Q(_zyGfifoF19_L412_data_0[2]));
Q_FDP4EP \_zyGfifoF19_L412_data_0_REG[1] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1376), .Q(_zyGfifoF19_L412_data_0[1]));
Q_FDP4EP \_zyGfifoF19_L412_data_0_REG[0] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1375), .Q(_zyGfifoF19_L412_data_0[0]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[63] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1708), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[63]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[62] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1707), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[62]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[61] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1706), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[61]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[60] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1705), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[60]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[59] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1704), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[59]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[58] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1703), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[58]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[57] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1702), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[57]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[56] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1701), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[56]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[55] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1700), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[55]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[54] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1699), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[54]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[53] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1698), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[53]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[52] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1697), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[52]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[51] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1696), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[51]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[50] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1695), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[50]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[49] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1694), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[49]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[48] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1693), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[48]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[47] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1692), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[47]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[46] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1691), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[46]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[45] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1690), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[45]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[44] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1689), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[44]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[43] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1688), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[43]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[42] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1687), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[42]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[41] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1686), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[41]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[40] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1685), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[40]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[39] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1684), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[39]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[38] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1683), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[38]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[37] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1682), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[37]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[36] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1681), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[36]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[35] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1680), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[35]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[34] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1679), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[34]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[33] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1678), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[33]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[32] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1677), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[32]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[31] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1676), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[31]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[30] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1675), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[30]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[29] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1674), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[29]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[28] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1673), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[28]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[27] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1672), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[27]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[26] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1671), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[26]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[25] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1670), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[25]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[24] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1669), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[24]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[23] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1668), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[23]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[22] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1667), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[22]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[21] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1666), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[21]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[20] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1665), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[20]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[19] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1664), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[19]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[18] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1663), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[18]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[17] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1662), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[17]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[16] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1661), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[16]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[15] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1660), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[15]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[14] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1659), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[14]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[13] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1658), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[13]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[12] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1657), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[12]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[11] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1656), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[11]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[10] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1655), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[10]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[9] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1654), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[9]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[8] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1653), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[8]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[7] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1652), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[7]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[6] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1651), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[6]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[5] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1650), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[5]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[4] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1649), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[4]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[3] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1648), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[3]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[2] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1647), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[2]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[1] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1646), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[1]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tdata_wr2_REG[0] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1645), .Q(_zzM2L368_mdxP3_kme_ib_tdata_wr2[0]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tstrb_wr3_REG[7] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1382), .Q(_zzM2L368_mdxP3_kme_ib_tstrb_wr3[7]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tstrb_wr3_REG[6] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1381), .Q(_zzM2L368_mdxP3_kme_ib_tstrb_wr3[6]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tstrb_wr3_REG[5] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1380), .Q(_zzM2L368_mdxP3_kme_ib_tstrb_wr3[5]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tstrb_wr3_REG[4] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1379), .Q(_zzM2L368_mdxP3_kme_ib_tstrb_wr3[4]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tstrb_wr3_REG[3] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1378), .Q(_zzM2L368_mdxP3_kme_ib_tstrb_wr3[3]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tstrb_wr3_REG[2] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1377), .Q(_zzM2L368_mdxP3_kme_ib_tstrb_wr3[2]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tstrb_wr3_REG[1] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1376), .Q(_zzM2L368_mdxP3_kme_ib_tstrb_wr3[1]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tstrb_wr3_REG[0] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1375), .Q(_zzM2L368_mdxP3_kme_ib_tstrb_wr3[0]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[63] ( .CK(clk), .CE(n37), .R(n1750), .D(n1708), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [63]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[62] ( .CK(clk), .CE(n37), .R(n1750), .D(n1707), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [62]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[61] ( .CK(clk), .CE(n37), .R(n1750), .D(n1706), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [61]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[60] ( .CK(clk), .CE(n37), .R(n1750), .D(n1705), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [60]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[59] ( .CK(clk), .CE(n37), .R(n1750), .D(n1704), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [59]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[58] ( .CK(clk), .CE(n37), .R(n1750), .D(n1703), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [58]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[57] ( .CK(clk), .CE(n37), .R(n1750), .D(n1702), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [57]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[56] ( .CK(clk), .CE(n37), .R(n1750), .D(n1701), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [56]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[55] ( .CK(clk), .CE(n37), .R(n1750), .D(n1700), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [55]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[54] ( .CK(clk), .CE(n37), .R(n1750), .D(n1699), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [54]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[53] ( .CK(clk), .CE(n37), .R(n1750), .D(n1698), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [53]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[52] ( .CK(clk), .CE(n37), .R(n1750), .D(n1697), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [52]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[51] ( .CK(clk), .CE(n37), .R(n1750), .D(n1696), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [51]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[50] ( .CK(clk), .CE(n37), .R(n1750), .D(n1695), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [50]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[49] ( .CK(clk), .CE(n37), .R(n1750), .D(n1694), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [49]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[48] ( .CK(clk), .CE(n37), .R(n1750), .D(n1693), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [48]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[47] ( .CK(clk), .CE(n37), .R(n1750), .D(n1692), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [47]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[46] ( .CK(clk), .CE(n37), .R(n1750), .D(n1691), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [46]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[45] ( .CK(clk), .CE(n37), .R(n1750), .D(n1690), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [45]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[44] ( .CK(clk), .CE(n37), .R(n1750), .D(n1689), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [44]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[43] ( .CK(clk), .CE(n37), .R(n1750), .D(n1688), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [43]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[42] ( .CK(clk), .CE(n37), .R(n1750), .D(n1687), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [42]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[41] ( .CK(clk), .CE(n37), .R(n1750), .D(n1686), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [41]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[40] ( .CK(clk), .CE(n37), .R(n1750), .D(n1685), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [40]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[39] ( .CK(clk), .CE(n37), .R(n1750), .D(n1684), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [39]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[38] ( .CK(clk), .CE(n37), .R(n1750), .D(n1683), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [38]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[37] ( .CK(clk), .CE(n37), .R(n1750), .D(n1682), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [37]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[36] ( .CK(clk), .CE(n37), .R(n1750), .D(n1681), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [36]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[35] ( .CK(clk), .CE(n37), .R(n1750), .D(n1680), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [35]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[34] ( .CK(clk), .CE(n37), .R(n1750), .D(n1679), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [34]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[33] ( .CK(clk), .CE(n37), .R(n1750), .D(n1678), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [33]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[32] ( .CK(clk), .CE(n37), .R(n1750), .D(n1677), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [32]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[31] ( .CK(clk), .CE(n37), .R(n1750), .D(n1676), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [31]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[30] ( .CK(clk), .CE(n37), .R(n1750), .D(n1675), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [30]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[29] ( .CK(clk), .CE(n37), .R(n1750), .D(n1674), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [29]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[28] ( .CK(clk), .CE(n37), .R(n1750), .D(n1673), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [28]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[27] ( .CK(clk), .CE(n37), .R(n1750), .D(n1672), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [27]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[26] ( .CK(clk), .CE(n37), .R(n1750), .D(n1671), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [26]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[25] ( .CK(clk), .CE(n37), .R(n1750), .D(n1670), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [25]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[24] ( .CK(clk), .CE(n37), .R(n1750), .D(n1669), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [24]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[23] ( .CK(clk), .CE(n37), .R(n1750), .D(n1668), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [23]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[22] ( .CK(clk), .CE(n37), .R(n1750), .D(n1667), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [22]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[21] ( .CK(clk), .CE(n37), .R(n1750), .D(n1666), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [21]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[20] ( .CK(clk), .CE(n37), .R(n1750), .D(n1665), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [20]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[19] ( .CK(clk), .CE(n37), .R(n1750), .D(n1664), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [19]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[18] ( .CK(clk), .CE(n37), .R(n1750), .D(n1663), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [18]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[17] ( .CK(clk), .CE(n37), .R(n1750), .D(n1662), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [17]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[16] ( .CK(clk), .CE(n37), .R(n1750), .D(n1661), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [16]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[15] ( .CK(clk), .CE(n37), .R(n1750), .D(n1660), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [15]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[14] ( .CK(clk), .CE(n37), .R(n1750), .D(n1659), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [14]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[13] ( .CK(clk), .CE(n37), .R(n1750), .D(n1658), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [13]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[12] ( .CK(clk), .CE(n37), .R(n1750), .D(n1657), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [12]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[11] ( .CK(clk), .CE(n37), .R(n1750), .D(n1656), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [11]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[10] ( .CK(clk), .CE(n37), .R(n1750), .D(n1655), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [10]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[9] ( .CK(clk), .CE(n37), .R(n1750), .D(n1654), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [9]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[8] ( .CK(clk), .CE(n37), .R(n1750), .D(n1653), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [8]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[7] ( .CK(clk), .CE(n37), .R(n1750), .D(n1652), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [7]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[6] ( .CK(clk), .CE(n37), .R(n1750), .D(n1651), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [6]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[5] ( .CK(clk), .CE(n37), .R(n1750), .D(n1650), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [5]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[4] ( .CK(clk), .CE(n37), .R(n1750), .D(n1649), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [4]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[3] ( .CK(clk), .CE(n37), .R(n1750), .D(n1648), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [3]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[2] ( .CK(clk), .CE(n37), .R(n1750), .D(n1647), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [2]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[1] ( .CK(clk), .CE(n37), .R(n1750), .D(n1646), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [1]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5_REG[0] ( .CK(clk), .CE(n37), .R(n1750), .D(n1645), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytdata_L207_tfiV5 [0]));
Q_FDP4EP \tdata_ib_REG[63] ( .CK(clk), .CE(n37), .R(n1750), .D(n1708), .Q(tdata_ib[63]));
Q_FDP4EP \tdata_ib_REG[62] ( .CK(clk), .CE(n37), .R(n1750), .D(n1707), .Q(tdata_ib[62]));
Q_FDP4EP \tdata_ib_REG[61] ( .CK(clk), .CE(n37), .R(n1750), .D(n1706), .Q(tdata_ib[61]));
Q_FDP4EP \tdata_ib_REG[60] ( .CK(clk), .CE(n37), .R(n1750), .D(n1705), .Q(tdata_ib[60]));
Q_FDP4EP \tdata_ib_REG[59] ( .CK(clk), .CE(n37), .R(n1750), .D(n1704), .Q(tdata_ib[59]));
Q_FDP4EP \tdata_ib_REG[58] ( .CK(clk), .CE(n37), .R(n1750), .D(n1703), .Q(tdata_ib[58]));
Q_FDP4EP \tdata_ib_REG[57] ( .CK(clk), .CE(n37), .R(n1750), .D(n1702), .Q(tdata_ib[57]));
Q_FDP4EP \tdata_ib_REG[56] ( .CK(clk), .CE(n37), .R(n1750), .D(n1701), .Q(tdata_ib[56]));
Q_FDP4EP \tdata_ib_REG[55] ( .CK(clk), .CE(n37), .R(n1750), .D(n1700), .Q(tdata_ib[55]));
Q_FDP4EP \tdata_ib_REG[54] ( .CK(clk), .CE(n37), .R(n1750), .D(n1699), .Q(tdata_ib[54]));
Q_FDP4EP \tdata_ib_REG[53] ( .CK(clk), .CE(n37), .R(n1750), .D(n1698), .Q(tdata_ib[53]));
Q_FDP4EP \tdata_ib_REG[52] ( .CK(clk), .CE(n37), .R(n1750), .D(n1697), .Q(tdata_ib[52]));
Q_FDP4EP \tdata_ib_REG[51] ( .CK(clk), .CE(n37), .R(n1750), .D(n1696), .Q(tdata_ib[51]));
Q_FDP4EP \tdata_ib_REG[50] ( .CK(clk), .CE(n37), .R(n1750), .D(n1695), .Q(tdata_ib[50]));
Q_FDP4EP \tdata_ib_REG[49] ( .CK(clk), .CE(n37), .R(n1750), .D(n1694), .Q(tdata_ib[49]));
Q_FDP4EP \tdata_ib_REG[48] ( .CK(clk), .CE(n37), .R(n1750), .D(n1693), .Q(tdata_ib[48]));
Q_FDP4EP \tdata_ib_REG[47] ( .CK(clk), .CE(n37), .R(n1750), .D(n1692), .Q(tdata_ib[47]));
Q_FDP4EP \tdata_ib_REG[46] ( .CK(clk), .CE(n37), .R(n1750), .D(n1691), .Q(tdata_ib[46]));
Q_FDP4EP \tdata_ib_REG[45] ( .CK(clk), .CE(n37), .R(n1750), .D(n1690), .Q(tdata_ib[45]));
Q_FDP4EP \tdata_ib_REG[44] ( .CK(clk), .CE(n37), .R(n1750), .D(n1689), .Q(tdata_ib[44]));
Q_FDP4EP \tdata_ib_REG[43] ( .CK(clk), .CE(n37), .R(n1750), .D(n1688), .Q(tdata_ib[43]));
Q_FDP4EP \tdata_ib_REG[42] ( .CK(clk), .CE(n37), .R(n1750), .D(n1687), .Q(tdata_ib[42]));
Q_FDP4EP \tdata_ib_REG[41] ( .CK(clk), .CE(n37), .R(n1750), .D(n1686), .Q(tdata_ib[41]));
Q_FDP4EP \tdata_ib_REG[40] ( .CK(clk), .CE(n37), .R(n1750), .D(n1685), .Q(tdata_ib[40]));
Q_FDP4EP \tdata_ib_REG[39] ( .CK(clk), .CE(n37), .R(n1750), .D(n1684), .Q(tdata_ib[39]));
Q_FDP4EP \tdata_ib_REG[38] ( .CK(clk), .CE(n37), .R(n1750), .D(n1683), .Q(tdata_ib[38]));
Q_FDP4EP \tdata_ib_REG[37] ( .CK(clk), .CE(n37), .R(n1750), .D(n1682), .Q(tdata_ib[37]));
Q_FDP4EP \tdata_ib_REG[36] ( .CK(clk), .CE(n37), .R(n1750), .D(n1681), .Q(tdata_ib[36]));
Q_FDP4EP \tdata_ib_REG[35] ( .CK(clk), .CE(n37), .R(n1750), .D(n1680), .Q(tdata_ib[35]));
Q_FDP4EP \tdata_ib_REG[34] ( .CK(clk), .CE(n37), .R(n1750), .D(n1679), .Q(tdata_ib[34]));
Q_FDP4EP \tdata_ib_REG[33] ( .CK(clk), .CE(n37), .R(n1750), .D(n1678), .Q(tdata_ib[33]));
Q_FDP4EP \tdata_ib_REG[32] ( .CK(clk), .CE(n37), .R(n1750), .D(n1677), .Q(tdata_ib[32]));
Q_FDP4EP \tdata_ib_REG[31] ( .CK(clk), .CE(n37), .R(n1750), .D(n1676), .Q(tdata_ib[31]));
Q_FDP4EP \tdata_ib_REG[30] ( .CK(clk), .CE(n37), .R(n1750), .D(n1675), .Q(tdata_ib[30]));
Q_FDP4EP \tdata_ib_REG[29] ( .CK(clk), .CE(n37), .R(n1750), .D(n1674), .Q(tdata_ib[29]));
Q_FDP4EP \tdata_ib_REG[28] ( .CK(clk), .CE(n37), .R(n1750), .D(n1673), .Q(tdata_ib[28]));
Q_FDP4EP \tdata_ib_REG[27] ( .CK(clk), .CE(n37), .R(n1750), .D(n1672), .Q(tdata_ib[27]));
Q_FDP4EP \tdata_ib_REG[26] ( .CK(clk), .CE(n37), .R(n1750), .D(n1671), .Q(tdata_ib[26]));
Q_FDP4EP \tdata_ib_REG[25] ( .CK(clk), .CE(n37), .R(n1750), .D(n1670), .Q(tdata_ib[25]));
Q_FDP4EP \tdata_ib_REG[24] ( .CK(clk), .CE(n37), .R(n1750), .D(n1669), .Q(tdata_ib[24]));
Q_FDP4EP \tdata_ib_REG[23] ( .CK(clk), .CE(n37), .R(n1750), .D(n1668), .Q(tdata_ib[23]));
Q_FDP4EP \tdata_ib_REG[22] ( .CK(clk), .CE(n37), .R(n1750), .D(n1667), .Q(tdata_ib[22]));
Q_FDP4EP \tdata_ib_REG[21] ( .CK(clk), .CE(n37), .R(n1750), .D(n1666), .Q(tdata_ib[21]));
Q_FDP4EP \tdata_ib_REG[20] ( .CK(clk), .CE(n37), .R(n1750), .D(n1665), .Q(tdata_ib[20]));
Q_FDP4EP \tdata_ib_REG[19] ( .CK(clk), .CE(n37), .R(n1750), .D(n1664), .Q(tdata_ib[19]));
Q_FDP4EP \tdata_ib_REG[18] ( .CK(clk), .CE(n37), .R(n1750), .D(n1663), .Q(tdata_ib[18]));
Q_FDP4EP \tdata_ib_REG[17] ( .CK(clk), .CE(n37), .R(n1750), .D(n1662), .Q(tdata_ib[17]));
Q_FDP4EP \tdata_ib_REG[16] ( .CK(clk), .CE(n37), .R(n1750), .D(n1661), .Q(tdata_ib[16]));
Q_FDP4EP \tdata_ib_REG[15] ( .CK(clk), .CE(n37), .R(n1750), .D(n1660), .Q(tdata_ib[15]));
Q_FDP4EP \tdata_ib_REG[14] ( .CK(clk), .CE(n37), .R(n1750), .D(n1659), .Q(tdata_ib[14]));
Q_FDP4EP \tdata_ib_REG[13] ( .CK(clk), .CE(n37), .R(n1750), .D(n1658), .Q(tdata_ib[13]));
Q_FDP4EP \tdata_ib_REG[12] ( .CK(clk), .CE(n37), .R(n1750), .D(n1657), .Q(tdata_ib[12]));
Q_FDP4EP \tdata_ib_REG[11] ( .CK(clk), .CE(n37), .R(n1750), .D(n1656), .Q(tdata_ib[11]));
Q_FDP4EP \tdata_ib_REG[10] ( .CK(clk), .CE(n37), .R(n1750), .D(n1655), .Q(tdata_ib[10]));
Q_FDP4EP \tdata_ib_REG[9] ( .CK(clk), .CE(n37), .R(n1750), .D(n1654), .Q(tdata_ib[9]));
Q_FDP4EP \tdata_ib_REG[8] ( .CK(clk), .CE(n37), .R(n1750), .D(n1653), .Q(tdata_ib[8]));
Q_FDP4EP \tdata_ib_REG[7] ( .CK(clk), .CE(n37), .R(n1750), .D(n1652), .Q(tdata_ib[7]));
Q_FDP4EP \tdata_ib_REG[6] ( .CK(clk), .CE(n37), .R(n1750), .D(n1651), .Q(tdata_ib[6]));
Q_FDP4EP \tdata_ib_REG[5] ( .CK(clk), .CE(n37), .R(n1750), .D(n1650), .Q(tdata_ib[5]));
Q_FDP4EP \tdata_ib_REG[4] ( .CK(clk), .CE(n37), .R(n1750), .D(n1649), .Q(tdata_ib[4]));
Q_FDP4EP \tdata_ib_REG[3] ( .CK(clk), .CE(n37), .R(n1750), .D(n1648), .Q(tdata_ib[3]));
Q_FDP4EP \tdata_ib_REG[2] ( .CK(clk), .CE(n37), .R(n1750), .D(n1647), .Q(tdata_ib[2]));
Q_FDP4EP \tdata_ib_REG[1] ( .CK(clk), .CE(n37), .R(n1750), .D(n1646), .Q(tdata_ib[1]));
Q_FDP4EP \tdata_ib_REG[0] ( .CK(clk), .CE(n37), .R(n1750), .D(n1645), .Q(tdata_ib[0]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[31] ( .CK(clk), .CE(n37), .R(n1750), .D(n1352), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [31]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[30] ( .CK(clk), .CE(n37), .R(n1750), .D(n1351), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [30]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[29] ( .CK(clk), .CE(n37), .R(n1750), .D(n1350), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [29]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[28] ( .CK(clk), .CE(n37), .R(n1750), .D(n1349), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [28]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[27] ( .CK(clk), .CE(n37), .R(n1750), .D(n1348), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [27]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[26] ( .CK(clk), .CE(n37), .R(n1750), .D(n1347), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [26]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[25] ( .CK(clk), .CE(n37), .R(n1750), .D(n1346), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [25]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[24] ( .CK(clk), .CE(n37), .R(n1750), .D(n1345), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [24]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[23] ( .CK(clk), .CE(n37), .R(n1750), .D(n1344), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [23]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[22] ( .CK(clk), .CE(n37), .R(n1750), .D(n1343), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [22]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[21] ( .CK(clk), .CE(n37), .R(n1750), .D(n1342), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [21]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[20] ( .CK(clk), .CE(n37), .R(n1750), .D(n1341), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [20]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[19] ( .CK(clk), .CE(n37), .R(n1750), .D(n1340), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [19]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[18] ( .CK(clk), .CE(n37), .R(n1750), .D(n1339), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [18]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[17] ( .CK(clk), .CE(n37), .R(n1750), .D(n1338), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [17]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[16] ( .CK(clk), .CE(n37), .R(n1750), .D(n1337), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [16]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[15] ( .CK(clk), .CE(n37), .R(n1750), .D(n1336), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [15]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[14] ( .CK(clk), .CE(n37), .R(n1750), .D(n1335), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [14]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[13] ( .CK(clk), .CE(n37), .R(n1750), .D(n1334), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [13]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[12] ( .CK(clk), .CE(n37), .R(n1750), .D(n1333), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [12]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[11] ( .CK(clk), .CE(n37), .R(n1750), .D(n1332), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [11]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[10] ( .CK(clk), .CE(n37), .R(n1750), .D(n1331), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [10]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[9] ( .CK(clk), .CE(n37), .R(n1750), .D(n1330), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [9]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[8] ( .CK(clk), .CE(n37), .R(n1750), .D(n1329), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [8]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[7] ( .CK(clk), .CE(n37), .R(n1750), .D(n1328), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [7]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[6] ( .CK(clk), .CE(n37), .R(n1750), .D(n1327), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [6]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[5] ( .CK(clk), .CE(n37), .R(n1750), .D(n1326), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [5]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[4] ( .CK(clk), .CE(n37), .R(n1750), .D(n1325), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [4]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[3] ( .CK(clk), .CE(n37), .R(n1750), .D(n1324), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [3]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[2] ( .CK(clk), .CE(n37), .R(n1750), .D(n1323), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [2]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[1] ( .CK(clk), .CE(n37), .R(n1750), .D(n1322), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [1]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6_REG[0] ( .CK(clk), .CE(n37), .R(n1750), .D(n1321), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytuser_string_L207_tfiV6 [0]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[31] ( .CK(clk), .CE(n37), .R(n1750), .D(n1414), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [31]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[30] ( .CK(clk), .CE(n37), .R(n1750), .D(n1413), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [30]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[29] ( .CK(clk), .CE(n37), .R(n1750), .D(n1412), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [29]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[28] ( .CK(clk), .CE(n37), .R(n1750), .D(n1411), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [28]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[27] ( .CK(clk), .CE(n37), .R(n1750), .D(n1410), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [27]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[26] ( .CK(clk), .CE(n37), .R(n1750), .D(n1409), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [26]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[25] ( .CK(clk), .CE(n37), .R(n1750), .D(n1408), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [25]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[24] ( .CK(clk), .CE(n37), .R(n1750), .D(n1407), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [24]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[23] ( .CK(clk), .CE(n37), .R(n1750), .D(n1406), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [23]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[22] ( .CK(clk), .CE(n37), .R(n1750), .D(n1405), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [22]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[21] ( .CK(clk), .CE(n37), .R(n1750), .D(n1404), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [21]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[20] ( .CK(clk), .CE(n37), .R(n1750), .D(n1403), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [20]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[19] ( .CK(clk), .CE(n37), .R(n1750), .D(n1402), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [19]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[18] ( .CK(clk), .CE(n37), .R(n1750), .D(n1401), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [18]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[17] ( .CK(clk), .CE(n37), .R(n1750), .D(n1400), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [17]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[16] ( .CK(clk), .CE(n37), .R(n1750), .D(n1399), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [16]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[15] ( .CK(clk), .CE(n37), .R(n1750), .D(n1398), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [15]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[14] ( .CK(clk), .CE(n37), .R(n1750), .D(n1397), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [14]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[13] ( .CK(clk), .CE(n37), .R(n1750), .D(n1396), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [13]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[12] ( .CK(clk), .CE(n37), .R(n1750), .D(n1395), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [12]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[11] ( .CK(clk), .CE(n37), .R(n1750), .D(n1394), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [11]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[10] ( .CK(clk), .CE(n37), .R(n1750), .D(n1393), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [10]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[9] ( .CK(clk), .CE(n37), .R(n1750), .D(n1392), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [9]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[8] ( .CK(clk), .CE(n37), .R(n1750), .D(n1391), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [8]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[7] ( .CK(clk), .CE(n37), .R(n1750), .D(n1390), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [7]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[6] ( .CK(clk), .CE(n37), .R(n1750), .D(n1389), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [6]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[5] ( .CK(clk), .CE(n37), .R(n1750), .D(n1388), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [5]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[4] ( .CK(clk), .CE(n37), .R(n1750), .D(n1387), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [4]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[3] ( .CK(clk), .CE(n37), .R(n1750), .D(n1386), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [3]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[2] ( .CK(clk), .CE(n37), .R(n1750), .D(n1385), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [2]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[1] ( .CK(clk), .CE(n37), .R(n1750), .D(n1384), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [1]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8_REG[0] ( .CK(clk), .CE(n37), .R(n1750), .D(n1383), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zystr_get_L207_tfiV8 [0]));
Q_FDP4EP \tuser_string_ib_REG[31] ( .CK(clk), .CE(n37), .R(n1750), .D(n1352), .Q(tuser_string_ib[31]));
Q_FDP4EP \tuser_string_ib_REG[30] ( .CK(clk), .CE(n37), .R(n1750), .D(n1351), .Q(tuser_string_ib[30]));
Q_FDP4EP \tuser_string_ib_REG[29] ( .CK(clk), .CE(n37), .R(n1750), .D(n1350), .Q(tuser_string_ib[29]));
Q_FDP4EP \tuser_string_ib_REG[28] ( .CK(clk), .CE(n37), .R(n1750), .D(n1349), .Q(tuser_string_ib[28]));
Q_FDP4EP \tuser_string_ib_REG[27] ( .CK(clk), .CE(n37), .R(n1750), .D(n1348), .Q(tuser_string_ib[27]));
Q_FDP4EP \tuser_string_ib_REG[26] ( .CK(clk), .CE(n37), .R(n1750), .D(n1347), .Q(tuser_string_ib[26]));
Q_FDP4EP \tuser_string_ib_REG[25] ( .CK(clk), .CE(n37), .R(n1750), .D(n1346), .Q(tuser_string_ib[25]));
Q_FDP4EP \tuser_string_ib_REG[24] ( .CK(clk), .CE(n37), .R(n1750), .D(n1345), .Q(tuser_string_ib[24]));
Q_FDP4EP \tuser_string_ib_REG[23] ( .CK(clk), .CE(n37), .R(n1750), .D(n1344), .Q(tuser_string_ib[23]));
Q_FDP4EP \tuser_string_ib_REG[22] ( .CK(clk), .CE(n37), .R(n1750), .D(n1343), .Q(tuser_string_ib[22]));
Q_FDP4EP \tuser_string_ib_REG[21] ( .CK(clk), .CE(n37), .R(n1750), .D(n1342), .Q(tuser_string_ib[21]));
Q_FDP4EP \tuser_string_ib_REG[20] ( .CK(clk), .CE(n37), .R(n1750), .D(n1341), .Q(tuser_string_ib[20]));
Q_FDP4EP \tuser_string_ib_REG[19] ( .CK(clk), .CE(n37), .R(n1750), .D(n1340), .Q(tuser_string_ib[19]));
Q_FDP4EP \tuser_string_ib_REG[18] ( .CK(clk), .CE(n37), .R(n1750), .D(n1339), .Q(tuser_string_ib[18]));
Q_FDP4EP \tuser_string_ib_REG[17] ( .CK(clk), .CE(n37), .R(n1750), .D(n1338), .Q(tuser_string_ib[17]));
Q_FDP4EP \tuser_string_ib_REG[16] ( .CK(clk), .CE(n37), .R(n1750), .D(n1337), .Q(tuser_string_ib[16]));
Q_FDP4EP \tuser_string_ib_REG[15] ( .CK(clk), .CE(n37), .R(n1750), .D(n1336), .Q(tuser_string_ib[15]));
Q_FDP4EP \tuser_string_ib_REG[14] ( .CK(clk), .CE(n37), .R(n1750), .D(n1335), .Q(tuser_string_ib[14]));
Q_FDP4EP \tuser_string_ib_REG[13] ( .CK(clk), .CE(n37), .R(n1750), .D(n1334), .Q(tuser_string_ib[13]));
Q_FDP4EP \tuser_string_ib_REG[12] ( .CK(clk), .CE(n37), .R(n1750), .D(n1333), .Q(tuser_string_ib[12]));
Q_FDP4EP \tuser_string_ib_REG[11] ( .CK(clk), .CE(n37), .R(n1750), .D(n1332), .Q(tuser_string_ib[11]));
Q_FDP4EP \tuser_string_ib_REG[10] ( .CK(clk), .CE(n37), .R(n1750), .D(n1331), .Q(tuser_string_ib[10]));
Q_FDP4EP \tuser_string_ib_REG[9] ( .CK(clk), .CE(n37), .R(n1750), .D(n1330), .Q(tuser_string_ib[9]));
Q_FDP4EP \tuser_string_ib_REG[8] ( .CK(clk), .CE(n37), .R(n1750), .D(n1329), .Q(tuser_string_ib[8]));
Q_FDP4EP \tuser_string_ib_REG[7] ( .CK(clk), .CE(n37), .R(n1750), .D(n1328), .Q(tuser_string_ib[7]));
Q_FDP4EP \tuser_string_ib_REG[6] ( .CK(clk), .CE(n37), .R(n1750), .D(n1327), .Q(tuser_string_ib[6]));
Q_FDP4EP \tuser_string_ib_REG[5] ( .CK(clk), .CE(n37), .R(n1750), .D(n1326), .Q(tuser_string_ib[5]));
Q_FDP4EP \tuser_string_ib_REG[4] ( .CK(clk), .CE(n37), .R(n1750), .D(n1325), .Q(tuser_string_ib[4]));
Q_FDP4EP \tuser_string_ib_REG[3] ( .CK(clk), .CE(n37), .R(n1750), .D(n1324), .Q(tuser_string_ib[3]));
Q_FDP4EP \tuser_string_ib_REG[2] ( .CK(clk), .CE(n37), .R(n1750), .D(n1323), .Q(tuser_string_ib[2]));
Q_FDP4EP \tuser_string_ib_REG[1] ( .CK(clk), .CE(n37), .R(n1750), .D(n1322), .Q(tuser_string_ib[1]));
Q_FDP4EP \tuser_string_ib_REG[0] ( .CK(clk), .CE(n37), .R(n1750), .D(n1321), .Q(tuser_string_ib[0]));
Q_FDP4EP \str_get_ib_REG[31] ( .CK(clk), .CE(n37), .R(n1750), .D(n1414), .Q(str_get_ib[31]));
Q_FDP4EP \str_get_ib_REG[30] ( .CK(clk), .CE(n37), .R(n1750), .D(n1413), .Q(str_get_ib[30]));
Q_FDP4EP \str_get_ib_REG[29] ( .CK(clk), .CE(n37), .R(n1750), .D(n1412), .Q(str_get_ib[29]));
Q_FDP4EP \str_get_ib_REG[28] ( .CK(clk), .CE(n37), .R(n1750), .D(n1411), .Q(str_get_ib[28]));
Q_FDP4EP \str_get_ib_REG[27] ( .CK(clk), .CE(n37), .R(n1750), .D(n1410), .Q(str_get_ib[27]));
Q_FDP4EP \str_get_ib_REG[26] ( .CK(clk), .CE(n37), .R(n1750), .D(n1409), .Q(str_get_ib[26]));
Q_FDP4EP \str_get_ib_REG[25] ( .CK(clk), .CE(n37), .R(n1750), .D(n1408), .Q(str_get_ib[25]));
Q_FDP4EP \str_get_ib_REG[24] ( .CK(clk), .CE(n37), .R(n1750), .D(n1407), .Q(str_get_ib[24]));
Q_FDP4EP \str_get_ib_REG[23] ( .CK(clk), .CE(n37), .R(n1750), .D(n1406), .Q(str_get_ib[23]));
Q_FDP4EP \str_get_ib_REG[22] ( .CK(clk), .CE(n37), .R(n1750), .D(n1405), .Q(str_get_ib[22]));
Q_FDP4EP \str_get_ib_REG[21] ( .CK(clk), .CE(n37), .R(n1750), .D(n1404), .Q(str_get_ib[21]));
Q_FDP4EP \str_get_ib_REG[20] ( .CK(clk), .CE(n37), .R(n1750), .D(n1403), .Q(str_get_ib[20]));
Q_FDP4EP \str_get_ib_REG[19] ( .CK(clk), .CE(n37), .R(n1750), .D(n1402), .Q(str_get_ib[19]));
Q_FDP4EP \str_get_ib_REG[18] ( .CK(clk), .CE(n37), .R(n1750), .D(n1401), .Q(str_get_ib[18]));
Q_FDP4EP \str_get_ib_REG[17] ( .CK(clk), .CE(n37), .R(n1750), .D(n1400), .Q(str_get_ib[17]));
Q_FDP4EP \str_get_ib_REG[16] ( .CK(clk), .CE(n37), .R(n1750), .D(n1399), .Q(str_get_ib[16]));
Q_FDP4EP \str_get_ib_REG[15] ( .CK(clk), .CE(n37), .R(n1750), .D(n1398), .Q(str_get_ib[15]));
Q_FDP4EP \str_get_ib_REG[14] ( .CK(clk), .CE(n37), .R(n1750), .D(n1397), .Q(str_get_ib[14]));
Q_FDP4EP \str_get_ib_REG[13] ( .CK(clk), .CE(n37), .R(n1750), .D(n1396), .Q(str_get_ib[13]));
Q_FDP4EP \str_get_ib_REG[12] ( .CK(clk), .CE(n37), .R(n1750), .D(n1395), .Q(str_get_ib[12]));
Q_FDP4EP \str_get_ib_REG[11] ( .CK(clk), .CE(n37), .R(n1750), .D(n1394), .Q(str_get_ib[11]));
Q_FDP4EP \str_get_ib_REG[10] ( .CK(clk), .CE(n37), .R(n1750), .D(n1393), .Q(str_get_ib[10]));
Q_FDP4EP \str_get_ib_REG[9] ( .CK(clk), .CE(n37), .R(n1750), .D(n1392), .Q(str_get_ib[9]));
Q_FDP4EP \str_get_ib_REG[8] ( .CK(clk), .CE(n37), .R(n1750), .D(n1391), .Q(str_get_ib[8]));
Q_FDP4EP \str_get_ib_REG[7] ( .CK(clk), .CE(n37), .R(n1750), .D(n1390), .Q(str_get_ib[7]));
Q_FDP4EP \str_get_ib_REG[6] ( .CK(clk), .CE(n37), .R(n1750), .D(n1389), .Q(str_get_ib[6]));
Q_FDP4EP \str_get_ib_REG[5] ( .CK(clk), .CE(n37), .R(n1750), .D(n1388), .Q(str_get_ib[5]));
Q_FDP4EP \str_get_ib_REG[4] ( .CK(clk), .CE(n37), .R(n1750), .D(n1387), .Q(str_get_ib[4]));
Q_FDP4EP \str_get_ib_REG[3] ( .CK(clk), .CE(n37), .R(n1750), .D(n1386), .Q(str_get_ib[3]));
Q_FDP4EP \str_get_ib_REG[2] ( .CK(clk), .CE(n37), .R(n1750), .D(n1385), .Q(str_get_ib[2]));
Q_FDP4EP \str_get_ib_REG[1] ( .CK(clk), .CE(n37), .R(n1750), .D(n1384), .Q(str_get_ib[1]));
Q_FDP4EP \str_get_ib_REG[0] ( .CK(clk), .CE(n37), .R(n1750), .D(n1383), .Q(str_get_ib[0]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytstrb_L207_tfiV7_REG[7] ( .CK(clk), .CE(n37), .R(n1750), .D(n1382), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytstrb_L207_tfiV7 [7]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytstrb_L207_tfiV7_REG[6] ( .CK(clk), .CE(n37), .R(n1750), .D(n1381), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytstrb_L207_tfiV7 [6]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytstrb_L207_tfiV7_REG[5] ( .CK(clk), .CE(n37), .R(n1750), .D(n1380), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytstrb_L207_tfiV7 [5]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytstrb_L207_tfiV7_REG[4] ( .CK(clk), .CE(n37), .R(n1750), .D(n1379), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytstrb_L207_tfiV7 [4]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytstrb_L207_tfiV7_REG[3] ( .CK(clk), .CE(n37), .R(n1750), .D(n1378), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytstrb_L207_tfiV7 [3]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytstrb_L207_tfiV7_REG[2] ( .CK(clk), .CE(n37), .R(n1750), .D(n1377), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytstrb_L207_tfiV7 [2]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytstrb_L207_tfiV7_REG[1] ( .CK(clk), .CE(n37), .R(n1750), .D(n1376), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytstrb_L207_tfiV7 [1]));
Q_FDP4EP \_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytstrb_L207_tfiV7_REG[0] ( .CK(clk), .CE(n37), .R(n1750), .D(n1375), .Q(\_zyL368_meSwitch4._zygfifotfiCscp1_L370_ib_service_data_isf_meScp5._zytstrb_L207_tfiV7 [0]));
Q_FDP4EP \tstrb_ib_REG[7] ( .CK(clk), .CE(n37), .R(n1750), .D(n1382), .Q(tstrb_ib[7]));
Q_FDP4EP \tstrb_ib_REG[6] ( .CK(clk), .CE(n37), .R(n1750), .D(n1381), .Q(tstrb_ib[6]));
Q_FDP4EP \tstrb_ib_REG[5] ( .CK(clk), .CE(n37), .R(n1750), .D(n1380), .Q(tstrb_ib[5]));
Q_FDP4EP \tstrb_ib_REG[4] ( .CK(clk), .CE(n37), .R(n1750), .D(n1379), .Q(tstrb_ib[4]));
Q_FDP4EP \tstrb_ib_REG[3] ( .CK(clk), .CE(n37), .R(n1750), .D(n1378), .Q(tstrb_ib[3]));
Q_FDP4EP \tstrb_ib_REG[2] ( .CK(clk), .CE(n37), .R(n1750), .D(n1377), .Q(tstrb_ib[2]));
Q_FDP4EP \tstrb_ib_REG[1] ( .CK(clk), .CE(n37), .R(n1750), .D(n1376), .Q(tstrb_ib[1]));
Q_FDP4EP \tstrb_ib_REG[0] ( .CK(clk), .CE(n37), .R(n1750), .D(n1375), .Q(tstrb_ib[0]));
Q_FDP4EP \_zygsfis_ib_service_data_rptr_REG[4] ( .CK(clk), .CE(n37), .R(n1750), .D(n1273), .Q(_zygsfis_ib_service_data_rptr[4]));
Q_FDP4EP \_zygsfis_ib_service_data_rptr_REG[3] ( .CK(clk), .CE(n37), .R(n1750), .D(n1272), .Q(_zygsfis_ib_service_data_rptr[3]));
Q_FDP4EP \_zygsfis_ib_service_data_rptr_REG[2] ( .CK(clk), .CE(n37), .R(n1750), .D(n1271), .Q(_zygsfis_ib_service_data_rptr[2]));
Q_FDP4EP \_zygsfis_ib_service_data_rptr_REG[1] ( .CK(clk), .CE(n37), .R(n1750), .D(n1270), .Q(_zygsfis_ib_service_data_rptr[1]));
Q_FDP4EP \_zygsfis_ib_service_data_rptr_REG[0] ( .CK(clk), .CE(n37), .R(n1750), .D(n1269), .Q(_zygsfis_ib_service_data_rptr[0]));
Q_FDP4EP \_zygsfis_ib_service_data_space_REG[4] ( .CK(clk), .CE(n37), .R(n1750), .D(n1465), .Q(_zygsfis_ib_service_data_space[4]));
Q_FDP4EP \_zygsfis_ib_service_data_space_REG[3] ( .CK(clk), .CE(n37), .R(n1750), .D(n1463), .Q(_zygsfis_ib_service_data_space[3]));
Q_FDP4EP \_zygsfis_ib_service_data_space_REG[2] ( .CK(clk), .CE(n37), .R(n1750), .D(n1461), .Q(_zygsfis_ib_service_data_space[2]));
Q_FDP4EP \_zygsfis_ib_service_data_space_REG[1] ( .CK(clk), .CE(n37), .R(n1750), .D(n1459), .Q(_zygsfis_ib_service_data_space[1]));
Q_FDP4EP \_zygsfis_ib_service_data_space_REG[0] ( .CK(clk), .CE(n37), .R(n1750), .D(n1457), .Q(_zygsfis_ib_service_data_space[0]));
Q_FDP4EP _zzM2L368_mdxP3_kme_ib_tlast_wr1_REG  ( .CK(clk), .CE(n1635), .R(n1750), .D(n1637), .Q(_zzM2L368_mdxP3_kme_ib_tlast_wr1));
Q_FDP4EP \_zyL372_tfiRv5_REG[24] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL372_tfiRv5[24]));
Q_FDP4EP \_zyL372_tfiRv5_REG[23] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL372_tfiRv5[23]));
Q_FDP4EP \_zyL372_tfiRv5_REG[22] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(_zyL372_tfiRv5[22]));
Q_FDP4EP \_zyL372_tfiRv5_REG[21] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL372_tfiRv5[21]));
Q_FDP4EP \_zyL372_tfiRv5_REG[20] ( .CK(clk), .CE(n37), .R(n1750), .D(n1632), .Q(_zyL372_tfiRv5[20]));
Q_FDP4EP \_zyL372_tfiRv5_REG[19] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL372_tfiRv5[19]));
Q_FDP4EP \_zyL372_tfiRv5_REG[18] ( .CK(clk), .CE(n37), .R(n1750), .D(n1631), .Q(_zyL372_tfiRv5[18]));
Q_FDP4EP \_zyL372_tfiRv5_REG[17] ( .CK(clk), .CE(n37), .R(n1750), .D(n1632), .Q(_zyL372_tfiRv5[17]));
Q_FDP4EP \_zyL372_tfiRv5_REG[16] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(_zyL372_tfiRv5[16]));
Q_FDP4EP \_zyL372_tfiRv5_REG[15] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL372_tfiRv5[15]));
Q_FDP4EP \_zyL372_tfiRv5_REG[14] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(_zyL372_tfiRv5[14]));
Q_FDP4EP \_zyL372_tfiRv5_REG[13] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(_zyL372_tfiRv5[13]));
Q_FDP4EP \_zyL372_tfiRv5_REG[12] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL372_tfiRv5[12]));
Q_FDP4EP \_zyL372_tfiRv5_REG[11] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(_zyL372_tfiRv5[11]));
Q_FDP4EP \_zyL372_tfiRv5_REG[10] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(_zyL372_tfiRv5[10]));
Q_FDP4EP \_zyL372_tfiRv5_REG[9] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(_zyL372_tfiRv5[9]));
Q_FDP4EP \_zyL372_tfiRv5_REG[8] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(_zyL372_tfiRv5[8]));
Q_FDP4EP \_zyL372_tfiRv5_REG[7] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL372_tfiRv5[7]));
Q_FDP4EP \_zyL372_tfiRv5_REG[6] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(_zyL372_tfiRv5[6]));
Q_FDP4EP \_zyL372_tfiRv5_REG[5] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL372_tfiRv5[5]));
Q_FDP4EP \_zyL372_tfiRv5_REG[4] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(_zyL372_tfiRv5[4]));
Q_FDP4EP \_zyL372_tfiRv5_REG[3] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL372_tfiRv5[3]));
Q_FDP4EP \_zyL372_tfiRv5_REG[2] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(_zyL372_tfiRv5[2]));
Q_FDP4EP \_zyL372_tfiRv5_REG[1] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL372_tfiRv5[1]));
Q_FDP4EP \_zyL372_tfiRv5_REG[0] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL372_tfiRv5[0]));
Q_FDP4EP \user_string_ib_REG[24] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(user_string_ib[24]));
Q_FDP4EP \user_string_ib_REG[23] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(user_string_ib[23]));
Q_FDP4EP \user_string_ib_REG[22] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(user_string_ib[22]));
Q_FDP4EP \user_string_ib_REG[21] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(user_string_ib[21]));
Q_FDP4EP \user_string_ib_REG[20] ( .CK(clk), .CE(n37), .R(n1750), .D(n1632), .Q(user_string_ib[20]));
Q_FDP4EP \user_string_ib_REG[19] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(user_string_ib[19]));
Q_FDP4EP \user_string_ib_REG[18] ( .CK(clk), .CE(n37), .R(n1750), .D(n1631), .Q(user_string_ib[18]));
Q_FDP4EP \user_string_ib_REG[17] ( .CK(clk), .CE(n37), .R(n1750), .D(n1632), .Q(user_string_ib[17]));
Q_FDP4EP \user_string_ib_REG[16] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(user_string_ib[16]));
Q_FDP4EP \user_string_ib_REG[15] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(user_string_ib[15]));
Q_FDP4EP \user_string_ib_REG[14] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(user_string_ib[14]));
Q_FDP4EP \user_string_ib_REG[13] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(user_string_ib[13]));
Q_FDP4EP \user_string_ib_REG[12] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(user_string_ib[12]));
Q_FDP4EP \user_string_ib_REG[11] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(user_string_ib[11]));
Q_FDP4EP \user_string_ib_REG[10] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(user_string_ib[10]));
Q_FDP4EP \user_string_ib_REG[9] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(user_string_ib[9]));
Q_FDP4EP \user_string_ib_REG[8] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(user_string_ib[8]));
Q_FDP4EP \user_string_ib_REG[7] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(user_string_ib[7]));
Q_FDP4EP \user_string_ib_REG[6] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(user_string_ib[6]));
Q_FDP4EP \user_string_ib_REG[5] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(user_string_ib[5]));
Q_FDP4EP \user_string_ib_REG[4] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(user_string_ib[4]));
Q_FDP4EP \user_string_ib_REG[3] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(user_string_ib[3]));
Q_FDP4EP \user_string_ib_REG[2] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(user_string_ib[2]));
Q_FDP4EP \user_string_ib_REG[1] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(user_string_ib[1]));
Q_FDP4EP \user_string_ib_REG[0] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(user_string_ib[0]));
Q_FDP4EP \_zyL406_tfiRv6_REG[7] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1750), .Q(_zyL406_tfiRv6[7]));
Q_FDP4EP \_zyL406_tfiRv6_REG[6] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1750), .Q(_zyL406_tfiRv6[6]));
Q_FDP4EP \_zyL406_tfiRv6_REG[5] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1750), .Q(_zyL406_tfiRv6[5]));
Q_FDP4EP \_zyL406_tfiRv6_REG[4] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1750), .Q(_zyL406_tfiRv6[4]));
Q_FDP4EP \_zyL406_tfiRv6_REG[3] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1750), .Q(_zyL406_tfiRv6[3]));
Q_FDP4EP \_zyL406_tfiRv6_REG[2] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1750), .Q(_zyL406_tfiRv6[2]));
Q_FDP4EP \_zyL406_tfiRv6_REG[1] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1358), .Q(_zyL406_tfiRv6[1]));
Q_FDP4EP \_zyL406_tfiRv6_REG[0] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1471), .Q(_zyL406_tfiRv6[0]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[31] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyGfifoF14_L373_data_0[31]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[30] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyGfifoF14_L373_data_0[30]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[29] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyGfifoF14_L373_data_0[29]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[28] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyGfifoF14_L373_data_0[28]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[27] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyGfifoF14_L373_data_0[27]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[26] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyGfifoF14_L373_data_0[26]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[25] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyGfifoF14_L373_data_0[25]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[24] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyGfifoF14_L373_data_0[24]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[23] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyGfifoF14_L373_data_0[23]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[22] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(_zyGfifoF14_L373_data_0[22]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[21] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyGfifoF14_L373_data_0[21]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[20] ( .CK(clk), .CE(n37), .R(n1750), .D(n1632), .Q(_zyGfifoF14_L373_data_0[20]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[19] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyGfifoF14_L373_data_0[19]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[18] ( .CK(clk), .CE(n37), .R(n1750), .D(n1631), .Q(_zyGfifoF14_L373_data_0[18]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[17] ( .CK(clk), .CE(n37), .R(n1750), .D(n1632), .Q(_zyGfifoF14_L373_data_0[17]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[16] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(_zyGfifoF14_L373_data_0[16]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[15] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyGfifoF14_L373_data_0[15]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[14] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(_zyGfifoF14_L373_data_0[14]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[13] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(_zyGfifoF14_L373_data_0[13]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[12] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyGfifoF14_L373_data_0[12]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[11] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(_zyGfifoF14_L373_data_0[11]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[10] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(_zyGfifoF14_L373_data_0[10]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[9] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(_zyGfifoF14_L373_data_0[9]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[8] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(_zyGfifoF14_L373_data_0[8]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[7] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyGfifoF14_L373_data_0[7]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[6] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(_zyGfifoF14_L373_data_0[6]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[5] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyGfifoF14_L373_data_0[5]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[4] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(_zyGfifoF14_L373_data_0[4]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[3] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyGfifoF14_L373_data_0[3]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[2] ( .CK(clk), .CE(n37), .R(n1750), .D(n1466), .Q(_zyGfifoF14_L373_data_0[2]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[1] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyGfifoF14_L373_data_0[1]));
Q_FDP4EP \_zyGfifoF14_L373_data_0_REG[0] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyGfifoF14_L373_data_0[0]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[31] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1750), .Q(_zyGfifoF18_L530_data_0[31]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[30] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1750), .Q(_zyGfifoF18_L530_data_0[30]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[29] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1750), .Q(_zyGfifoF18_L530_data_0[29]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[28] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1750), .Q(_zyGfifoF18_L530_data_0[28]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[27] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1750), .Q(_zyGfifoF18_L530_data_0[27]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[26] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1750), .Q(_zyGfifoF18_L530_data_0[26]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[25] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1750), .Q(_zyGfifoF18_L530_data_0[25]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[24] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1750), .Q(_zyGfifoF18_L530_data_0[24]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[23] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1750), .Q(_zyGfifoF18_L530_data_0[23]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[22] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1466), .Q(_zyGfifoF18_L530_data_0[22]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[21] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1750), .Q(_zyGfifoF18_L530_data_0[21]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[20] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1632), .Q(_zyGfifoF18_L530_data_0[20]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[19] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1750), .Q(_zyGfifoF18_L530_data_0[19]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[18] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1631), .Q(_zyGfifoF18_L530_data_0[18]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[17] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1632), .Q(_zyGfifoF18_L530_data_0[17]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[16] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1466), .Q(_zyGfifoF18_L530_data_0[16]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[15] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1750), .Q(_zyGfifoF18_L530_data_0[15]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[14] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1466), .Q(_zyGfifoF18_L530_data_0[14]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[13] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1466), .Q(_zyGfifoF18_L530_data_0[13]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[12] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1750), .Q(_zyGfifoF18_L530_data_0[12]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[11] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1466), .Q(_zyGfifoF18_L530_data_0[11]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[10] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1466), .Q(_zyGfifoF18_L530_data_0[10]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[9] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1466), .Q(_zyGfifoF18_L530_data_0[9]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[8] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1466), .Q(_zyGfifoF18_L530_data_0[8]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[7] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1750), .Q(_zyGfifoF18_L530_data_0[7]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[6] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1466), .Q(_zyGfifoF18_L530_data_0[6]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[5] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1750), .Q(_zyGfifoF18_L530_data_0[5]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[4] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1466), .Q(_zyGfifoF18_L530_data_0[4]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[3] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1750), .Q(_zyGfifoF18_L530_data_0[3]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[2] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1466), .Q(_zyGfifoF18_L530_data_0[2]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[1] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1750), .Q(_zyGfifoF18_L530_data_0[1]));
Q_FDP4EP \_zyGfifoF18_L530_data_0_REG[0] ( .CK(clk), .CE(n1640), .R(n1750), .D(n1750), .Q(_zyGfifoF18_L530_data_0[0]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tuser_wr4_REG[7] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1750), .Q(_zzM2L368_mdxP3_kme_ib_tuser_wr4[7]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tuser_wr4_REG[6] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1750), .Q(_zzM2L368_mdxP3_kme_ib_tuser_wr4[6]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tuser_wr4_REG[5] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1750), .Q(_zzM2L368_mdxP3_kme_ib_tuser_wr4[5]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tuser_wr4_REG[4] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1750), .Q(_zzM2L368_mdxP3_kme_ib_tuser_wr4[4]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tuser_wr4_REG[3] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1750), .Q(_zzM2L368_mdxP3_kme_ib_tuser_wr4[3]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tuser_wr4_REG[2] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1750), .Q(_zzM2L368_mdxP3_kme_ib_tuser_wr4[2]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tuser_wr4_REG[1] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1468), .Q(_zzM2L368_mdxP3_kme_ib_tuser_wr4[1]));
Q_FDP4EP \_zzM2L368_mdxP3_kme_ib_tuser_wr4_REG[0] ( .CK(clk), .CE(n1635), .R(n1750), .D(n1467), .Q(_zzM2L368_mdxP3_kme_ib_tuser_wr4[0]));
Q_FDP4EP \_zyL370_tfiRv18_REG[31] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[31]));
Q_FDP4EP \_zyL370_tfiRv18_REG[30] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[30]));
Q_FDP4EP \_zyL370_tfiRv18_REG[29] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[29]));
Q_FDP4EP \_zyL370_tfiRv18_REG[28] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[28]));
Q_FDP4EP \_zyL370_tfiRv18_REG[27] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[27]));
Q_FDP4EP \_zyL370_tfiRv18_REG[26] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[26]));
Q_FDP4EP \_zyL370_tfiRv18_REG[25] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[25]));
Q_FDP4EP \_zyL370_tfiRv18_REG[24] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[24]));
Q_FDP4EP \_zyL370_tfiRv18_REG[23] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[23]));
Q_FDP4EP \_zyL370_tfiRv18_REG[22] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[22]));
Q_FDP4EP \_zyL370_tfiRv18_REG[21] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[21]));
Q_FDP4EP \_zyL370_tfiRv18_REG[20] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[20]));
Q_FDP4EP \_zyL370_tfiRv18_REG[19] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[19]));
Q_FDP4EP \_zyL370_tfiRv18_REG[18] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[18]));
Q_FDP4EP \_zyL370_tfiRv18_REG[17] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[17]));
Q_FDP4EP \_zyL370_tfiRv18_REG[16] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[16]));
Q_FDP4EP \_zyL370_tfiRv18_REG[15] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[15]));
Q_FDP4EP \_zyL370_tfiRv18_REG[14] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[14]));
Q_FDP4EP \_zyL370_tfiRv18_REG[13] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[13]));
Q_FDP4EP \_zyL370_tfiRv18_REG[12] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[12]));
Q_FDP4EP \_zyL370_tfiRv18_REG[11] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[11]));
Q_FDP4EP \_zyL370_tfiRv18_REG[10] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[10]));
Q_FDP4EP \_zyL370_tfiRv18_REG[9] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[9]));
Q_FDP4EP \_zyL370_tfiRv18_REG[8] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[8]));
Q_FDP4EP \_zyL370_tfiRv18_REG[7] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[7]));
Q_FDP4EP \_zyL370_tfiRv18_REG[6] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[6]));
Q_FDP4EP \_zyL370_tfiRv18_REG[5] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[5]));
Q_FDP4EP \_zyL370_tfiRv18_REG[4] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[4]));
Q_FDP4EP \_zyL370_tfiRv18_REG[3] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[3]));
Q_FDP4EP \_zyL370_tfiRv18_REG[2] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(_zyL370_tfiRv18[2]));
Q_FDP4EP \_zyL370_tfiRv18_REG[1] ( .CK(clk), .CE(n37), .R(n1750), .D(n1639), .Q(_zyL370_tfiRv18[1]));
Q_FDP4EP \_zyL370_tfiRv18_REG[0] ( .CK(clk), .CE(n37), .R(n1750), .D(n1629), .Q(_zyL370_tfiRv18[0]));
Q_FDP4EP \retval_ib_REG[31] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[31]));
Q_FDP4EP \retval_ib_REG[30] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[30]));
Q_FDP4EP \retval_ib_REG[29] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[29]));
Q_FDP4EP \retval_ib_REG[28] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[28]));
Q_FDP4EP \retval_ib_REG[27] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[27]));
Q_FDP4EP \retval_ib_REG[26] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[26]));
Q_FDP4EP \retval_ib_REG[25] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[25]));
Q_FDP4EP \retval_ib_REG[24] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[24]));
Q_FDP4EP \retval_ib_REG[23] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[23]));
Q_FDP4EP \retval_ib_REG[22] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[22]));
Q_FDP4EP \retval_ib_REG[21] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[21]));
Q_FDP4EP \retval_ib_REG[20] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[20]));
Q_FDP4EP \retval_ib_REG[19] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[19]));
Q_FDP4EP \retval_ib_REG[18] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[18]));
Q_FDP4EP \retval_ib_REG[17] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[17]));
Q_FDP4EP \retval_ib_REG[16] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[16]));
Q_FDP4EP \retval_ib_REG[15] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[15]));
Q_FDP4EP \retval_ib_REG[14] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[14]));
Q_FDP4EP \retval_ib_REG[13] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[13]));
Q_FDP4EP \retval_ib_REG[12] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[12]));
Q_FDP4EP \retval_ib_REG[11] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[11]));
Q_FDP4EP \retval_ib_REG[10] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[10]));
Q_FDP4EP \retval_ib_REG[9] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[9]));
Q_FDP4EP \retval_ib_REG[8] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[8]));
Q_FDP4EP \retval_ib_REG[7] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[7]));
Q_FDP4EP \retval_ib_REG[6] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[6]));
Q_FDP4EP \retval_ib_REG[5] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[5]));
Q_FDP4EP \retval_ib_REG[4] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[4]));
Q_FDP4EP \retval_ib_REG[3] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[3]));
Q_FDP4EP \retval_ib_REG[2] ( .CK(clk), .CE(n37), .R(n1750), .D(n1750), .Q(retval_ib[2]));
Q_FDP4EP \retval_ib_REG[1] ( .CK(clk), .CE(n37), .R(n1750), .D(n1639), .Q(retval_ib[1]));
Q_FDP4EP \retval_ib_REG[0] ( .CK(clk), .CE(n37), .R(n1750), .D(n1629), .Q(retval_ib[0]));
Q_FDP4EP _zyictd_finish_L454_2_REG  ( .CK(clk), .CE(n3310), .R(n1750), .D(n5382), .Q(_zyictd_finish_L454_2));
Q_INV U7271 ( .A(n3390), .Z(n34));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[63] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[63]), .Q(_zyGfifoF25_L460_data_0[63]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[62] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[62]), .Q(_zyGfifoF25_L460_data_0[62]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[61] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[61]), .Q(_zyGfifoF25_L460_data_0[61]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[60] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[60]), .Q(_zyGfifoF25_L460_data_0[60]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[59] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[59]), .Q(_zyGfifoF25_L460_data_0[59]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[58] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[58]), .Q(_zyGfifoF25_L460_data_0[58]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[57] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[57]), .Q(_zyGfifoF25_L460_data_0[57]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[56] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[56]), .Q(_zyGfifoF25_L460_data_0[56]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[55] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[55]), .Q(_zyGfifoF25_L460_data_0[55]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[54] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[54]), .Q(_zyGfifoF25_L460_data_0[54]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[53] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[53]), .Q(_zyGfifoF25_L460_data_0[53]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[52] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[52]), .Q(_zyGfifoF25_L460_data_0[52]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[51] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[51]), .Q(_zyGfifoF25_L460_data_0[51]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[50] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[50]), .Q(_zyGfifoF25_L460_data_0[50]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[49] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[49]), .Q(_zyGfifoF25_L460_data_0[49]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[48] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[48]), .Q(_zyGfifoF25_L460_data_0[48]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[47] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[47]), .Q(_zyGfifoF25_L460_data_0[47]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[46] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[46]), .Q(_zyGfifoF25_L460_data_0[46]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[45] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[45]), .Q(_zyGfifoF25_L460_data_0[45]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[44] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[44]), .Q(_zyGfifoF25_L460_data_0[44]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[43] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[43]), .Q(_zyGfifoF25_L460_data_0[43]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[42] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[42]), .Q(_zyGfifoF25_L460_data_0[42]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[41] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[41]), .Q(_zyGfifoF25_L460_data_0[41]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[40] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[40]), .Q(_zyGfifoF25_L460_data_0[40]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[39] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[39]), .Q(_zyGfifoF25_L460_data_0[39]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[38] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[38]), .Q(_zyGfifoF25_L460_data_0[38]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[37] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[37]), .Q(_zyGfifoF25_L460_data_0[37]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[36] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[36]), .Q(_zyGfifoF25_L460_data_0[36]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[35] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[35]), .Q(_zyGfifoF25_L460_data_0[35]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[34] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[34]), .Q(_zyGfifoF25_L460_data_0[34]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[33] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[33]), .Q(_zyGfifoF25_L460_data_0[33]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[32] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[32]), .Q(_zyGfifoF25_L460_data_0[32]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[31] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[31]), .Q(_zyGfifoF25_L460_data_0[31]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[30] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[30]), .Q(_zyGfifoF25_L460_data_0[30]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[29] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[29]), .Q(_zyGfifoF25_L460_data_0[29]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[28] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[28]), .Q(_zyGfifoF25_L460_data_0[28]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[27] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[27]), .Q(_zyGfifoF25_L460_data_0[27]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[26] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[26]), .Q(_zyGfifoF25_L460_data_0[26]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[25] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[25]), .Q(_zyGfifoF25_L460_data_0[25]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[24] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[24]), .Q(_zyGfifoF25_L460_data_0[24]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[23] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[23]), .Q(_zyGfifoF25_L460_data_0[23]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[22] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[22]), .Q(_zyGfifoF25_L460_data_0[22]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[21] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[21]), .Q(_zyGfifoF25_L460_data_0[21]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[20] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[20]), .Q(_zyGfifoF25_L460_data_0[20]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[19] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[19]), .Q(_zyGfifoF25_L460_data_0[19]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[18] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[18]), .Q(_zyGfifoF25_L460_data_0[18]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[17] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[17]), .Q(_zyGfifoF25_L460_data_0[17]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[16] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[16]), .Q(_zyGfifoF25_L460_data_0[16]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[15] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[15]), .Q(_zyGfifoF25_L460_data_0[15]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[14] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[14]), .Q(_zyGfifoF25_L460_data_0[14]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[13] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[13]), .Q(_zyGfifoF25_L460_data_0[13]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[12] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[12]), .Q(_zyGfifoF25_L460_data_0[12]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[11] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[11]), .Q(_zyGfifoF25_L460_data_0[11]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[10] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[10]), .Q(_zyGfifoF25_L460_data_0[10]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[9] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[9]), .Q(_zyGfifoF25_L460_data_0[9]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[8] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[8]), .Q(_zyGfifoF25_L460_data_0[8]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[7] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[7]), .Q(_zyGfifoF25_L460_data_0[7]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[6] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[6]), .Q(_zyGfifoF25_L460_data_0[6]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[5] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[5]), .Q(_zyGfifoF25_L460_data_0[5]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[4] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[4]), .Q(_zyGfifoF25_L460_data_0[4]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[3] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[3]), .Q(_zyGfifoF25_L460_data_0[3]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[2] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[2]), .Q(_zyGfifoF25_L460_data_0[2]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[1] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[1]), .Q(_zyGfifoF25_L460_data_0[1]));
Q_FDP4EP \_zyGfifoF25_L460_data_0_REG[0] ( .CK(clk), .CE(n34), .R(n1750), .D(kme_ob_tdata[0]), .Q(_zyGfifoF25_L460_data_0[0]));
Q_INV U7336 ( .A(n3322), .Z(n33));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[127] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[63]), .Q(_zyGfifoF28_L482_data_0[127]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[126] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[62]), .Q(_zyGfifoF28_L482_data_0[126]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[125] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[61]), .Q(_zyGfifoF28_L482_data_0[125]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[124] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[60]), .Q(_zyGfifoF28_L482_data_0[124]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[123] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[59]), .Q(_zyGfifoF28_L482_data_0[123]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[122] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[58]), .Q(_zyGfifoF28_L482_data_0[122]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[121] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[57]), .Q(_zyGfifoF28_L482_data_0[121]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[120] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[56]), .Q(_zyGfifoF28_L482_data_0[120]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[119] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[55]), .Q(_zyGfifoF28_L482_data_0[119]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[118] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[54]), .Q(_zyGfifoF28_L482_data_0[118]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[117] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[53]), .Q(_zyGfifoF28_L482_data_0[117]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[116] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[52]), .Q(_zyGfifoF28_L482_data_0[116]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[115] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[51]), .Q(_zyGfifoF28_L482_data_0[115]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[114] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[50]), .Q(_zyGfifoF28_L482_data_0[114]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[113] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[49]), .Q(_zyGfifoF28_L482_data_0[113]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[112] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[48]), .Q(_zyGfifoF28_L482_data_0[112]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[111] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[47]), .Q(_zyGfifoF28_L482_data_0[111]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[110] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[46]), .Q(_zyGfifoF28_L482_data_0[110]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[109] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[45]), .Q(_zyGfifoF28_L482_data_0[109]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[108] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[44]), .Q(_zyGfifoF28_L482_data_0[108]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[107] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[43]), .Q(_zyGfifoF28_L482_data_0[107]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[106] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[42]), .Q(_zyGfifoF28_L482_data_0[106]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[105] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[41]), .Q(_zyGfifoF28_L482_data_0[105]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[104] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[40]), .Q(_zyGfifoF28_L482_data_0[104]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[103] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[39]), .Q(_zyGfifoF28_L482_data_0[103]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[102] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[38]), .Q(_zyGfifoF28_L482_data_0[102]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[101] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[37]), .Q(_zyGfifoF28_L482_data_0[101]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[100] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[36]), .Q(_zyGfifoF28_L482_data_0[100]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[99] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[35]), .Q(_zyGfifoF28_L482_data_0[99]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[98] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[34]), .Q(_zyGfifoF28_L482_data_0[98]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[97] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[33]), .Q(_zyGfifoF28_L482_data_0[97]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[96] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[32]), .Q(_zyGfifoF28_L482_data_0[96]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[95] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[31]), .Q(_zyGfifoF28_L482_data_0[95]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[94] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[30]), .Q(_zyGfifoF28_L482_data_0[94]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[93] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[29]), .Q(_zyGfifoF28_L482_data_0[93]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[92] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[28]), .Q(_zyGfifoF28_L482_data_0[92]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[91] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[27]), .Q(_zyGfifoF28_L482_data_0[91]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[90] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[26]), .Q(_zyGfifoF28_L482_data_0[90]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[89] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[25]), .Q(_zyGfifoF28_L482_data_0[89]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[88] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[24]), .Q(_zyGfifoF28_L482_data_0[88]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[87] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[23]), .Q(_zyGfifoF28_L482_data_0[87]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[86] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[22]), .Q(_zyGfifoF28_L482_data_0[86]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[85] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[21]), .Q(_zyGfifoF28_L482_data_0[85]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[84] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[20]), .Q(_zyGfifoF28_L482_data_0[84]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[83] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[19]), .Q(_zyGfifoF28_L482_data_0[83]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[82] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[18]), .Q(_zyGfifoF28_L482_data_0[82]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[81] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[17]), .Q(_zyGfifoF28_L482_data_0[81]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[80] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[16]), .Q(_zyGfifoF28_L482_data_0[80]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[79] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[15]), .Q(_zyGfifoF28_L482_data_0[79]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[78] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[14]), .Q(_zyGfifoF28_L482_data_0[78]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[77] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[13]), .Q(_zyGfifoF28_L482_data_0[77]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[76] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[12]), .Q(_zyGfifoF28_L482_data_0[76]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[75] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[11]), .Q(_zyGfifoF28_L482_data_0[75]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[74] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[10]), .Q(_zyGfifoF28_L482_data_0[74]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[73] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[9]), .Q(_zyGfifoF28_L482_data_0[73]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[72] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[8]), .Q(_zyGfifoF28_L482_data_0[72]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[71] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[7]), .Q(_zyGfifoF28_L482_data_0[71]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[70] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[6]), .Q(_zyGfifoF28_L482_data_0[70]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[69] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[5]), .Q(_zyGfifoF28_L482_data_0[69]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[68] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[4]), .Q(_zyGfifoF28_L482_data_0[68]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[67] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[3]), .Q(_zyGfifoF28_L482_data_0[67]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[66] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[2]), .Q(_zyGfifoF28_L482_data_0[66]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[65] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[1]), .Q(_zyGfifoF28_L482_data_0[65]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[64] ( .CK(clk), .CE(n33), .R(n1750), .D(kme_ob_tdata[0]), .Q(_zyGfifoF28_L482_data_0[64]));
Q_INV U7401 ( .A(n3338), .Z(n32));
Q_FDP4EP \_zyGfifoF29_L487_data_0_REG[15] ( .CK(clk), .CE(n32), .R(n1750), .D(kme_ob_tuser[7]), .Q(_zyGfifoF29_L487_data_0[15]));
Q_FDP4EP \_zyGfifoF29_L487_data_0_REG[14] ( .CK(clk), .CE(n32), .R(n1750), .D(kme_ob_tuser[6]), .Q(_zyGfifoF29_L487_data_0[14]));
Q_FDP4EP \_zyGfifoF29_L487_data_0_REG[13] ( .CK(clk), .CE(n32), .R(n1750), .D(kme_ob_tuser[5]), .Q(_zyGfifoF29_L487_data_0[13]));
Q_FDP4EP \_zyGfifoF29_L487_data_0_REG[12] ( .CK(clk), .CE(n32), .R(n1750), .D(kme_ob_tuser[4]), .Q(_zyGfifoF29_L487_data_0[12]));
Q_FDP4EP \_zyGfifoF29_L487_data_0_REG[11] ( .CK(clk), .CE(n32), .R(n1750), .D(kme_ob_tuser[3]), .Q(_zyGfifoF29_L487_data_0[11]));
Q_FDP4EP \_zyGfifoF29_L487_data_0_REG[10] ( .CK(clk), .CE(n32), .R(n1750), .D(kme_ob_tuser[2]), .Q(_zyGfifoF29_L487_data_0[10]));
Q_FDP4EP \_zyGfifoF29_L487_data_0_REG[9] ( .CK(clk), .CE(n32), .R(n1750), .D(kme_ob_tuser[1]), .Q(_zyGfifoF29_L487_data_0[9]));
Q_FDP4EP \_zyGfifoF29_L487_data_0_REG[8] ( .CK(clk), .CE(n32), .R(n1750), .D(kme_ob_tuser[0]), .Q(_zyGfifoF29_L487_data_0[8]));
Q_INV U7410 ( .A(n3343), .Z(n31));
Q_FDP4EP \_zyGfifoF30_L491_data_0_REG[15] ( .CK(clk), .CE(n31), .R(n1750), .D(kme_ob_tstrb[7]), .Q(_zyGfifoF30_L491_data_0[15]));
Q_FDP4EP \_zyGfifoF30_L491_data_0_REG[14] ( .CK(clk), .CE(n31), .R(n1750), .D(kme_ob_tstrb[6]), .Q(_zyGfifoF30_L491_data_0[14]));
Q_FDP4EP \_zyGfifoF30_L491_data_0_REG[13] ( .CK(clk), .CE(n31), .R(n1750), .D(kme_ob_tstrb[5]), .Q(_zyGfifoF30_L491_data_0[13]));
Q_FDP4EP \_zyGfifoF30_L491_data_0_REG[12] ( .CK(clk), .CE(n31), .R(n1750), .D(kme_ob_tstrb[4]), .Q(_zyGfifoF30_L491_data_0[12]));
Q_FDP4EP \_zyGfifoF30_L491_data_0_REG[11] ( .CK(clk), .CE(n31), .R(n1750), .D(kme_ob_tstrb[3]), .Q(_zyGfifoF30_L491_data_0[11]));
Q_FDP4EP \_zyGfifoF30_L491_data_0_REG[10] ( .CK(clk), .CE(n31), .R(n1750), .D(kme_ob_tstrb[2]), .Q(_zyGfifoF30_L491_data_0[10]));
Q_FDP4EP \_zyGfifoF30_L491_data_0_REG[9] ( .CK(clk), .CE(n31), .R(n1750), .D(kme_ob_tstrb[1]), .Q(_zyGfifoF30_L491_data_0[9]));
Q_FDP4EP \_zyGfifoF30_L491_data_0_REG[8] ( .CK(clk), .CE(n31), .R(n1750), .D(kme_ob_tstrb[0]), .Q(_zyGfifoF30_L491_data_0[8]));
Q_INV U7419 ( .A(n3348), .Z(n30));
Q_FDP4EP \_zyGfifoF31_L496_data_0_REG[8] ( .CK(clk), .CE(n30), .R(n1750), .D(kme_ob_tlast), .Q(_zyGfifoF31_L496_data_0[8]));
Q_FDP4EP _zzM2L439_mdxP4_En_REG  ( .CK(clk), .CE(n3551), .R(n1750), .D(_zzM2L439_mdxP4_EnNxt), .Q(_zzM2L439_mdxP4_En));
Q_INV U7422 ( .A(_zygsfis_ob_service_data_req[4]), .Z(n29));
Q_FDP4EP \_zygsfis_ob_service_data_req_REG[4] ( .CK(clk), .CE(n5877), .R(n1750), .D(n29), .Q(_zygsfis_ob_service_data_req[4]));
Q_FDP4EP \_zygsfis_ob_service_data_req_REG[3] ( .CK(clk), .CE(n3559), .R(n1750), .D(n2382), .Q(_zygsfis_ob_service_data_req[3]));
Q_FDP4EP \_zygsfis_ob_service_data_req_REG[2] ( .CK(clk), .CE(n3559), .R(n1750), .D(n2380), .Q(_zygsfis_ob_service_data_req[2]));
Q_FDP4EP \_zygsfis_ob_service_data_req_REG[1] ( .CK(clk), .CE(n3559), .R(n1750), .D(n2378), .Q(_zygsfis_ob_service_data_req[1]));
Q_INV U7427 ( .A(_zygsfis_ob_service_data_req[0]), .Z(n28));
Q_FDP4EP \_zygsfis_ob_service_data_req_REG[0] ( .CK(clk), .CE(n3559), .R(n1750), .D(n28), .Q(_zygsfis_ob_service_data_req[0]));
Q_FDP4EP _zyGfifoF20_L209_req_0_REG  ( .CK(clk), .CE(n3559), .R(n1750), .D(n1898), .Q(_zyGfifoF20_L209_req_0));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[31] ( .CK(clk), .CE(n3559), .R(n1750), .D(n1750), .Q(_zyGfifoF20_L209_data_0[31]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[30] ( .CK(clk), .CE(n3559), .R(n1750), .D(n1750), .Q(_zyGfifoF20_L209_data_0[30]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[29] ( .CK(clk), .CE(n3559), .R(n1750), .D(n1750), .Q(_zyGfifoF20_L209_data_0[29]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[28] ( .CK(clk), .CE(n3559), .R(n1750), .D(n1750), .Q(_zyGfifoF20_L209_data_0[28]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[27] ( .CK(clk), .CE(n3559), .R(n1750), .D(n1750), .Q(_zyGfifoF20_L209_data_0[27]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[26] ( .CK(clk), .CE(n3559), .R(n1750), .D(n1750), .Q(_zyGfifoF20_L209_data_0[26]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[25] ( .CK(clk), .CE(n3559), .R(n1750), .D(n1750), .Q(_zyGfifoF20_L209_data_0[25]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[24] ( .CK(clk), .CE(n3559), .R(n1750), .D(n1750), .Q(_zyGfifoF20_L209_data_0[24]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[23] ( .CK(clk), .CE(n3559), .R(n1750), .D(n1750), .Q(_zyGfifoF20_L209_data_0[23]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[22] ( .CK(clk), .CE(n3559), .R(n1750), .D(n1750), .Q(_zyGfifoF20_L209_data_0[22]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[21] ( .CK(clk), .CE(n3559), .R(n1750), .D(n1750), .Q(_zyGfifoF20_L209_data_0[21]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[20] ( .CK(clk), .CE(n3559), .R(n1750), .D(n1750), .Q(_zyGfifoF20_L209_data_0[20]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[19] ( .CK(clk), .CE(n3559), .R(n1750), .D(n1750), .Q(_zyGfifoF20_L209_data_0[19]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[18] ( .CK(clk), .CE(n3559), .R(n1750), .D(n1750), .Q(_zyGfifoF20_L209_data_0[18]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[17] ( .CK(clk), .CE(n3559), .R(n1750), .D(n1750), .Q(_zyGfifoF20_L209_data_0[17]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[16] ( .CK(clk), .CE(n3559), .R(n1750), .D(n1750), .Q(_zyGfifoF20_L209_data_0[16]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[15] ( .CK(clk), .CE(n3559), .R(n1750), .D(n1750), .Q(_zyGfifoF20_L209_data_0[15]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[14] ( .CK(clk), .CE(n3559), .R(n1750), .D(n1750), .Q(_zyGfifoF20_L209_data_0[14]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[13] ( .CK(clk), .CE(n3559), .R(n1750), .D(n1750), .Q(_zyGfifoF20_L209_data_0[13]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[12] ( .CK(clk), .CE(n3559), .R(n1750), .D(n1750), .Q(_zyGfifoF20_L209_data_0[12]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[11] ( .CK(clk), .CE(n3559), .R(n1750), .D(n1750), .Q(_zyGfifoF20_L209_data_0[11]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[10] ( .CK(clk), .CE(n3559), .R(n1750), .D(n1750), .Q(_zyGfifoF20_L209_data_0[10]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[9] ( .CK(clk), .CE(n3559), .R(n1750), .D(n1750), .Q(_zyGfifoF20_L209_data_0[9]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[8] ( .CK(clk), .CE(n3559), .R(n1750), .D(n1750), .Q(_zyGfifoF20_L209_data_0[8]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[7] ( .CK(clk), .CE(n3559), .R(n1750), .D(n1750), .Q(_zyGfifoF20_L209_data_0[7]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[6] ( .CK(clk), .CE(n3559), .R(n1750), .D(n1750), .Q(_zyGfifoF20_L209_data_0[6]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[5] ( .CK(clk), .CE(n3559), .R(n1750), .D(n1750), .Q(_zyGfifoF20_L209_data_0[5]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[4] ( .CK(clk), .CE(n3559), .R(n1750), .D(n2431), .Q(_zyGfifoF20_L209_data_0[4]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[3] ( .CK(clk), .CE(n3559), .R(n1750), .D(n2430), .Q(_zyGfifoF20_L209_data_0[3]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[2] ( .CK(clk), .CE(n3559), .R(n1750), .D(n2429), .Q(_zyGfifoF20_L209_data_0[2]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[1] ( .CK(clk), .CE(n3559), .R(n1750), .D(n2428), .Q(_zyGfifoF20_L209_data_0[1]));
Q_FDP4EP \_zyGfifoF20_L209_data_0_REG[0] ( .CK(clk), .CE(n3559), .R(n1750), .D(n2427), .Q(_zyGfifoF20_L209_data_0[0]));
Q_INV U7462 ( .A(n3316), .Z(n27));
Q_FDP4EP _zyGfifoF0_L439_s2_req_5_REG  ( .CK(clk), .CE(n27), .R(n1750), .D(n3093), .Q(_zyGfifoF0_L439_s2_req_5));
Q_FDP4EP \_zyGfifoF0_L439_s2_cbid_5_REG[19] ( .CK(clk), .CE(n27), .R(n1750), .D(n3092), .Q(_zyGfifoF0_L439_s2_cbid_5[19]));
Q_FDP4EP \_zyGfifoF0_L439_s2_cbid_5_REG[18] ( .CK(clk), .CE(n27), .R(n1750), .D(n3091), .Q(_zyGfifoF0_L439_s2_cbid_5[18]));
Q_FDP4EP \_zyGfifoF0_L439_s2_cbid_5_REG[17] ( .CK(clk), .CE(n27), .R(n1750), .D(n3090), .Q(_zyGfifoF0_L439_s2_cbid_5[17]));
Q_FDP4EP \_zyGfifoF0_L439_s2_cbid_5_REG[16] ( .CK(clk), .CE(n27), .R(n1750), .D(n3089), .Q(_zyGfifoF0_L439_s2_cbid_5[16]));
Q_FDP4EP \_zyGfifoF0_L439_s2_cbid_5_REG[15] ( .CK(clk), .CE(n27), .R(n1750), .D(n3088), .Q(_zyGfifoF0_L439_s2_cbid_5[15]));
Q_FDP4EP \_zyGfifoF0_L439_s2_cbid_5_REG[14] ( .CK(clk), .CE(n27), .R(n1750), .D(n3087), .Q(_zyGfifoF0_L439_s2_cbid_5[14]));
Q_FDP4EP \_zyGfifoF0_L439_s2_cbid_5_REG[13] ( .CK(clk), .CE(n27), .R(n1750), .D(n3086), .Q(_zyGfifoF0_L439_s2_cbid_5[13]));
Q_FDP4EP \_zyGfifoF0_L439_s2_cbid_5_REG[12] ( .CK(clk), .CE(n27), .R(n1750), .D(n3085), .Q(_zyGfifoF0_L439_s2_cbid_5[12]));
Q_FDP4EP \_zyGfifoF0_L439_s2_cbid_5_REG[11] ( .CK(clk), .CE(n27), .R(n1750), .D(n3084), .Q(_zyGfifoF0_L439_s2_cbid_5[11]));
Q_FDP4EP \_zyGfifoF0_L439_s2_cbid_5_REG[10] ( .CK(clk), .CE(n27), .R(n1750), .D(n3083), .Q(_zyGfifoF0_L439_s2_cbid_5[10]));
Q_FDP4EP \_zyGfifoF0_L439_s2_cbid_5_REG[9] ( .CK(clk), .CE(n27), .R(n1750), .D(n3082), .Q(_zyGfifoF0_L439_s2_cbid_5[9]));
Q_FDP4EP \_zyGfifoF0_L439_s2_cbid_5_REG[8] ( .CK(clk), .CE(n27), .R(n1750), .D(n3081), .Q(_zyGfifoF0_L439_s2_cbid_5[8]));
Q_FDP4EP \_zyGfifoF0_L439_s2_cbid_5_REG[7] ( .CK(clk), .CE(n27), .R(n1750), .D(n3080), .Q(_zyGfifoF0_L439_s2_cbid_5[7]));
Q_FDP4EP \_zyGfifoF0_L439_s2_cbid_5_REG[6] ( .CK(clk), .CE(n27), .R(n1750), .D(n3079), .Q(_zyGfifoF0_L439_s2_cbid_5[6]));
Q_FDP4EP \_zyGfifoF0_L439_s2_cbid_5_REG[5] ( .CK(clk), .CE(n27), .R(n1750), .D(n3078), .Q(_zyGfifoF0_L439_s2_cbid_5[5]));
Q_FDP4EP \_zyGfifoF0_L439_s2_cbid_5_REG[4] ( .CK(clk), .CE(n27), .R(n1750), .D(n3077), .Q(_zyGfifoF0_L439_s2_cbid_5[4]));
Q_FDP4EP \_zyGfifoF0_L439_s2_cbid_5_REG[3] ( .CK(clk), .CE(n27), .R(n1750), .D(n3076), .Q(_zyGfifoF0_L439_s2_cbid_5[3]));
Q_FDP4EP \_zyGfifoF0_L439_s2_cbid_5_REG[2] ( .CK(clk), .CE(n27), .R(n1750), .D(n3075), .Q(_zyGfifoF0_L439_s2_cbid_5[2]));
Q_FDP4EP \_zyGfifoF0_L439_s2_cbid_5_REG[1] ( .CK(clk), .CE(n27), .R(n1750), .D(n3074), .Q(_zyGfifoF0_L439_s2_cbid_5[1]));
Q_FDP4EP \_zyGfifoF0_L439_s2_cbid_5_REG[0] ( .CK(clk), .CE(n27), .R(n1750), .D(n3073), .Q(_zyGfifoF0_L439_s2_cbid_5[0]));
Q_INV U7484 ( .A(n3319), .Z(n26));
Q_FDP4EP _zyGfifoF23_L444_req_0_REG  ( .CK(clk), .CE(n26), .R(n1750), .D(n1900), .Q(_zyGfifoF23_L444_req_0));
Q_INV U7486 ( .A(n3320), .Z(n25));
Q_FDP4EP _zyGfifoF24_L446_req_0_REG  ( .CK(clk), .CE(n25), .R(n1750), .D(n1901), .Q(_zyGfifoF24_L446_req_0));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[135] ( .CK(clk), .CE(n25), .R(n1750), .D(n1972), .Q(_zyGfifoF24_L446_data_0[135]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[134] ( .CK(clk), .CE(n25), .R(n1750), .D(n1971), .Q(_zyGfifoF24_L446_data_0[134]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[133] ( .CK(clk), .CE(n25), .R(n1750), .D(n1970), .Q(_zyGfifoF24_L446_data_0[133]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[132] ( .CK(clk), .CE(n25), .R(n1750), .D(n1969), .Q(_zyGfifoF24_L446_data_0[132]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[131] ( .CK(clk), .CE(n25), .R(n1750), .D(n1968), .Q(_zyGfifoF24_L446_data_0[131]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[130] ( .CK(clk), .CE(n25), .R(n1750), .D(n1967), .Q(_zyGfifoF24_L446_data_0[130]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[129] ( .CK(clk), .CE(n25), .R(n1750), .D(n1966), .Q(_zyGfifoF24_L446_data_0[129]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[128] ( .CK(clk), .CE(n25), .R(n1750), .D(n1965), .Q(_zyGfifoF24_L446_data_0[128]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[127] ( .CK(clk), .CE(n25), .R(n1750), .D(n1964), .Q(_zyGfifoF24_L446_data_0[127]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[126] ( .CK(clk), .CE(n25), .R(n1750), .D(n1963), .Q(_zyGfifoF24_L446_data_0[126]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[125] ( .CK(clk), .CE(n25), .R(n1750), .D(n1962), .Q(_zyGfifoF24_L446_data_0[125]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[124] ( .CK(clk), .CE(n25), .R(n1750), .D(n1961), .Q(_zyGfifoF24_L446_data_0[124]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[123] ( .CK(clk), .CE(n25), .R(n1750), .D(n1960), .Q(_zyGfifoF24_L446_data_0[123]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[122] ( .CK(clk), .CE(n25), .R(n1750), .D(n1959), .Q(_zyGfifoF24_L446_data_0[122]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[121] ( .CK(clk), .CE(n25), .R(n1750), .D(n1958), .Q(_zyGfifoF24_L446_data_0[121]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[120] ( .CK(clk), .CE(n25), .R(n1750), .D(n1957), .Q(_zyGfifoF24_L446_data_0[120]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[119] ( .CK(clk), .CE(n25), .R(n1750), .D(n1956), .Q(_zyGfifoF24_L446_data_0[119]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[118] ( .CK(clk), .CE(n25), .R(n1750), .D(n1955), .Q(_zyGfifoF24_L446_data_0[118]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[117] ( .CK(clk), .CE(n25), .R(n1750), .D(n1954), .Q(_zyGfifoF24_L446_data_0[117]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[116] ( .CK(clk), .CE(n25), .R(n1750), .D(n1953), .Q(_zyGfifoF24_L446_data_0[116]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[115] ( .CK(clk), .CE(n25), .R(n1750), .D(n1952), .Q(_zyGfifoF24_L446_data_0[115]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[114] ( .CK(clk), .CE(n25), .R(n1750), .D(n1951), .Q(_zyGfifoF24_L446_data_0[114]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[113] ( .CK(clk), .CE(n25), .R(n1750), .D(n1950), .Q(_zyGfifoF24_L446_data_0[113]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[112] ( .CK(clk), .CE(n25), .R(n1750), .D(n1949), .Q(_zyGfifoF24_L446_data_0[112]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[111] ( .CK(clk), .CE(n25), .R(n1750), .D(n1948), .Q(_zyGfifoF24_L446_data_0[111]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[110] ( .CK(clk), .CE(n25), .R(n1750), .D(n1947), .Q(_zyGfifoF24_L446_data_0[110]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[109] ( .CK(clk), .CE(n25), .R(n1750), .D(n1946), .Q(_zyGfifoF24_L446_data_0[109]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[108] ( .CK(clk), .CE(n25), .R(n1750), .D(n1945), .Q(_zyGfifoF24_L446_data_0[108]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[107] ( .CK(clk), .CE(n25), .R(n1750), .D(n1944), .Q(_zyGfifoF24_L446_data_0[107]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[106] ( .CK(clk), .CE(n25), .R(n1750), .D(n1943), .Q(_zyGfifoF24_L446_data_0[106]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[105] ( .CK(clk), .CE(n25), .R(n1750), .D(n1942), .Q(_zyGfifoF24_L446_data_0[105]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[104] ( .CK(clk), .CE(n25), .R(n1750), .D(n1941), .Q(_zyGfifoF24_L446_data_0[104]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[103] ( .CK(clk), .CE(n25), .R(n1750), .D(n1940), .Q(_zyGfifoF24_L446_data_0[103]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[102] ( .CK(clk), .CE(n25), .R(n1750), .D(n1939), .Q(_zyGfifoF24_L446_data_0[102]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[101] ( .CK(clk), .CE(n25), .R(n1750), .D(n1938), .Q(_zyGfifoF24_L446_data_0[101]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[100] ( .CK(clk), .CE(n25), .R(n1750), .D(n1937), .Q(_zyGfifoF24_L446_data_0[100]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[99] ( .CK(clk), .CE(n25), .R(n1750), .D(n1936), .Q(_zyGfifoF24_L446_data_0[99]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[98] ( .CK(clk), .CE(n25), .R(n1750), .D(n1935), .Q(_zyGfifoF24_L446_data_0[98]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[97] ( .CK(clk), .CE(n25), .R(n1750), .D(n1934), .Q(_zyGfifoF24_L446_data_0[97]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[96] ( .CK(clk), .CE(n25), .R(n1750), .D(n1933), .Q(_zyGfifoF24_L446_data_0[96]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[95] ( .CK(clk), .CE(n25), .R(n1750), .D(n1932), .Q(_zyGfifoF24_L446_data_0[95]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[94] ( .CK(clk), .CE(n25), .R(n1750), .D(n1931), .Q(_zyGfifoF24_L446_data_0[94]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[93] ( .CK(clk), .CE(n25), .R(n1750), .D(n1930), .Q(_zyGfifoF24_L446_data_0[93]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[92] ( .CK(clk), .CE(n25), .R(n1750), .D(n1929), .Q(_zyGfifoF24_L446_data_0[92]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[91] ( .CK(clk), .CE(n25), .R(n1750), .D(n1928), .Q(_zyGfifoF24_L446_data_0[91]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[90] ( .CK(clk), .CE(n25), .R(n1750), .D(n1927), .Q(_zyGfifoF24_L446_data_0[90]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[89] ( .CK(clk), .CE(n25), .R(n1750), .D(n1926), .Q(_zyGfifoF24_L446_data_0[89]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[88] ( .CK(clk), .CE(n25), .R(n1750), .D(n1925), .Q(_zyGfifoF24_L446_data_0[88]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[87] ( .CK(clk), .CE(n25), .R(n1750), .D(n1924), .Q(_zyGfifoF24_L446_data_0[87]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[86] ( .CK(clk), .CE(n25), .R(n1750), .D(n1923), .Q(_zyGfifoF24_L446_data_0[86]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[85] ( .CK(clk), .CE(n25), .R(n1750), .D(n1922), .Q(_zyGfifoF24_L446_data_0[85]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[84] ( .CK(clk), .CE(n25), .R(n1750), .D(n1921), .Q(_zyGfifoF24_L446_data_0[84]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[83] ( .CK(clk), .CE(n25), .R(n1750), .D(n1920), .Q(_zyGfifoF24_L446_data_0[83]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[82] ( .CK(clk), .CE(n25), .R(n1750), .D(n1919), .Q(_zyGfifoF24_L446_data_0[82]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[81] ( .CK(clk), .CE(n25), .R(n1750), .D(n1918), .Q(_zyGfifoF24_L446_data_0[81]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[80] ( .CK(clk), .CE(n25), .R(n1750), .D(n1917), .Q(_zyGfifoF24_L446_data_0[80]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[79] ( .CK(clk), .CE(n25), .R(n1750), .D(n1916), .Q(_zyGfifoF24_L446_data_0[79]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[78] ( .CK(clk), .CE(n25), .R(n1750), .D(n1915), .Q(_zyGfifoF24_L446_data_0[78]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[77] ( .CK(clk), .CE(n25), .R(n1750), .D(n1914), .Q(_zyGfifoF24_L446_data_0[77]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[76] ( .CK(clk), .CE(n25), .R(n1750), .D(n1913), .Q(_zyGfifoF24_L446_data_0[76]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[75] ( .CK(clk), .CE(n25), .R(n1750), .D(n1912), .Q(_zyGfifoF24_L446_data_0[75]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[74] ( .CK(clk), .CE(n25), .R(n1750), .D(n1911), .Q(_zyGfifoF24_L446_data_0[74]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[73] ( .CK(clk), .CE(n25), .R(n1750), .D(n1910), .Q(_zyGfifoF24_L446_data_0[73]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[72] ( .CK(clk), .CE(n25), .R(n1750), .D(n1909), .Q(_zyGfifoF24_L446_data_0[72]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[71] ( .CK(clk), .CE(n25), .R(n1750), .D(n2108), .Q(_zyGfifoF24_L446_data_0[71]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[70] ( .CK(clk), .CE(n25), .R(n1750), .D(n2107), .Q(_zyGfifoF24_L446_data_0[70]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[69] ( .CK(clk), .CE(n25), .R(n1750), .D(n2106), .Q(_zyGfifoF24_L446_data_0[69]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[68] ( .CK(clk), .CE(n25), .R(n1750), .D(n2105), .Q(_zyGfifoF24_L446_data_0[68]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[67] ( .CK(clk), .CE(n25), .R(n1750), .D(n2104), .Q(_zyGfifoF24_L446_data_0[67]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[66] ( .CK(clk), .CE(n25), .R(n1750), .D(n2103), .Q(_zyGfifoF24_L446_data_0[66]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[65] ( .CK(clk), .CE(n25), .R(n1750), .D(n2102), .Q(_zyGfifoF24_L446_data_0[65]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[64] ( .CK(clk), .CE(n25), .R(n1750), .D(n2101), .Q(_zyGfifoF24_L446_data_0[64]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[63] ( .CK(clk), .CE(n25), .R(n1750), .D(n2100), .Q(_zyGfifoF24_L446_data_0[63]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[62] ( .CK(clk), .CE(n25), .R(n1750), .D(n2099), .Q(_zyGfifoF24_L446_data_0[62]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[61] ( .CK(clk), .CE(n25), .R(n1750), .D(n2098), .Q(_zyGfifoF24_L446_data_0[61]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[60] ( .CK(clk), .CE(n25), .R(n1750), .D(n2097), .Q(_zyGfifoF24_L446_data_0[60]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[59] ( .CK(clk), .CE(n25), .R(n1750), .D(n2096), .Q(_zyGfifoF24_L446_data_0[59]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[58] ( .CK(clk), .CE(n25), .R(n1750), .D(n2095), .Q(_zyGfifoF24_L446_data_0[58]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[57] ( .CK(clk), .CE(n25), .R(n1750), .D(n2094), .Q(_zyGfifoF24_L446_data_0[57]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[56] ( .CK(clk), .CE(n25), .R(n1750), .D(n2093), .Q(_zyGfifoF24_L446_data_0[56]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[55] ( .CK(clk), .CE(n25), .R(n1750), .D(n2092), .Q(_zyGfifoF24_L446_data_0[55]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[54] ( .CK(clk), .CE(n25), .R(n1750), .D(n2091), .Q(_zyGfifoF24_L446_data_0[54]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[53] ( .CK(clk), .CE(n25), .R(n1750), .D(n2090), .Q(_zyGfifoF24_L446_data_0[53]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[52] ( .CK(clk), .CE(n25), .R(n1750), .D(n2089), .Q(_zyGfifoF24_L446_data_0[52]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[51] ( .CK(clk), .CE(n25), .R(n1750), .D(n2088), .Q(_zyGfifoF24_L446_data_0[51]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[50] ( .CK(clk), .CE(n25), .R(n1750), .D(n2087), .Q(_zyGfifoF24_L446_data_0[50]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[49] ( .CK(clk), .CE(n25), .R(n1750), .D(n2086), .Q(_zyGfifoF24_L446_data_0[49]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[48] ( .CK(clk), .CE(n25), .R(n1750), .D(n2085), .Q(_zyGfifoF24_L446_data_0[48]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[47] ( .CK(clk), .CE(n25), .R(n1750), .D(n2084), .Q(_zyGfifoF24_L446_data_0[47]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[46] ( .CK(clk), .CE(n25), .R(n1750), .D(n2083), .Q(_zyGfifoF24_L446_data_0[46]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[45] ( .CK(clk), .CE(n25), .R(n1750), .D(n2082), .Q(_zyGfifoF24_L446_data_0[45]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[44] ( .CK(clk), .CE(n25), .R(n1750), .D(n2081), .Q(_zyGfifoF24_L446_data_0[44]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[43] ( .CK(clk), .CE(n25), .R(n1750), .D(n2080), .Q(_zyGfifoF24_L446_data_0[43]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[42] ( .CK(clk), .CE(n25), .R(n1750), .D(n2079), .Q(_zyGfifoF24_L446_data_0[42]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[41] ( .CK(clk), .CE(n25), .R(n1750), .D(n2078), .Q(_zyGfifoF24_L446_data_0[41]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[40] ( .CK(clk), .CE(n25), .R(n1750), .D(n2077), .Q(_zyGfifoF24_L446_data_0[40]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[39] ( .CK(clk), .CE(n25), .R(n1750), .D(n2138), .Q(_zyGfifoF24_L446_data_0[39]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[38] ( .CK(clk), .CE(n25), .R(n1750), .D(n2137), .Q(_zyGfifoF24_L446_data_0[38]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[37] ( .CK(clk), .CE(n25), .R(n1750), .D(n2136), .Q(_zyGfifoF24_L446_data_0[37]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[36] ( .CK(clk), .CE(n25), .R(n1750), .D(n2135), .Q(_zyGfifoF24_L446_data_0[36]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[35] ( .CK(clk), .CE(n25), .R(n1750), .D(n2134), .Q(_zyGfifoF24_L446_data_0[35]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[34] ( .CK(clk), .CE(n25), .R(n1750), .D(n2133), .Q(_zyGfifoF24_L446_data_0[34]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[33] ( .CK(clk), .CE(n25), .R(n1750), .D(n2132), .Q(_zyGfifoF24_L446_data_0[33]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[32] ( .CK(clk), .CE(n25), .R(n1750), .D(n2131), .Q(_zyGfifoF24_L446_data_0[32]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[31] ( .CK(clk), .CE(n25), .R(n1750), .D(n2182), .Q(_zyGfifoF24_L446_data_0[31]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[30] ( .CK(clk), .CE(n25), .R(n1750), .D(n2181), .Q(_zyGfifoF24_L446_data_0[30]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[29] ( .CK(clk), .CE(n25), .R(n1750), .D(n2180), .Q(_zyGfifoF24_L446_data_0[29]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[28] ( .CK(clk), .CE(n25), .R(n1750), .D(n2179), .Q(_zyGfifoF24_L446_data_0[28]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[27] ( .CK(clk), .CE(n25), .R(n1750), .D(n2178), .Q(_zyGfifoF24_L446_data_0[27]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[26] ( .CK(clk), .CE(n25), .R(n1750), .D(n2177), .Q(_zyGfifoF24_L446_data_0[26]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[25] ( .CK(clk), .CE(n25), .R(n1750), .D(n2176), .Q(_zyGfifoF24_L446_data_0[25]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[24] ( .CK(clk), .CE(n25), .R(n1750), .D(n2175), .Q(_zyGfifoF24_L446_data_0[24]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[23] ( .CK(clk), .CE(n25), .R(n1750), .D(n2174), .Q(_zyGfifoF24_L446_data_0[23]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[22] ( .CK(clk), .CE(n25), .R(n1750), .D(n2173), .Q(_zyGfifoF24_L446_data_0[22]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[21] ( .CK(clk), .CE(n25), .R(n1750), .D(n2172), .Q(_zyGfifoF24_L446_data_0[21]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[20] ( .CK(clk), .CE(n25), .R(n1750), .D(n2171), .Q(_zyGfifoF24_L446_data_0[20]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[19] ( .CK(clk), .CE(n25), .R(n1750), .D(n2170), .Q(_zyGfifoF24_L446_data_0[19]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[18] ( .CK(clk), .CE(n25), .R(n1750), .D(n2169), .Q(_zyGfifoF24_L446_data_0[18]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[17] ( .CK(clk), .CE(n25), .R(n1750), .D(n2168), .Q(_zyGfifoF24_L446_data_0[17]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[16] ( .CK(clk), .CE(n25), .R(n1750), .D(n2167), .Q(_zyGfifoF24_L446_data_0[16]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[15] ( .CK(clk), .CE(n25), .R(n1750), .D(n2166), .Q(_zyGfifoF24_L446_data_0[15]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[14] ( .CK(clk), .CE(n25), .R(n1750), .D(n2165), .Q(_zyGfifoF24_L446_data_0[14]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[13] ( .CK(clk), .CE(n25), .R(n1750), .D(n2164), .Q(_zyGfifoF24_L446_data_0[13]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[12] ( .CK(clk), .CE(n25), .R(n1750), .D(n2163), .Q(_zyGfifoF24_L446_data_0[12]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[11] ( .CK(clk), .CE(n25), .R(n1750), .D(n2162), .Q(_zyGfifoF24_L446_data_0[11]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[10] ( .CK(clk), .CE(n25), .R(n1750), .D(n2161), .Q(_zyGfifoF24_L446_data_0[10]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[9] ( .CK(clk), .CE(n25), .R(n1750), .D(n2160), .Q(_zyGfifoF24_L446_data_0[9]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[8] ( .CK(clk), .CE(n25), .R(n1750), .D(n2159), .Q(_zyGfifoF24_L446_data_0[8]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[7] ( .CK(clk), .CE(n25), .R(n1750), .D(n2158), .Q(_zyGfifoF24_L446_data_0[7]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[6] ( .CK(clk), .CE(n25), .R(n1750), .D(n2157), .Q(_zyGfifoF24_L446_data_0[6]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[5] ( .CK(clk), .CE(n25), .R(n1750), .D(n2156), .Q(_zyGfifoF24_L446_data_0[5]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[4] ( .CK(clk), .CE(n25), .R(n1750), .D(n2155), .Q(_zyGfifoF24_L446_data_0[4]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[3] ( .CK(clk), .CE(n25), .R(n1750), .D(n2154), .Q(_zyGfifoF24_L446_data_0[3]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[2] ( .CK(clk), .CE(n25), .R(n1750), .D(n2153), .Q(_zyGfifoF24_L446_data_0[2]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[1] ( .CK(clk), .CE(n25), .R(n1750), .D(n2152), .Q(_zyGfifoF24_L446_data_0[1]));
Q_FDP4EP \_zyGfifoF24_L446_data_0_REG[0] ( .CK(clk), .CE(n25), .R(n1750), .D(n2151), .Q(_zyGfifoF24_L446_data_0[0]));
Q_FDP4EP _zyGfifoF25_L460_req_0_REG  ( .CK(clk), .CE(n34), .R(n1750), .D(n1902), .Q(_zyGfifoF25_L460_req_0));
Q_FDP4EP _zyGfifoF26_L530_req_0_REG  ( .CK(clk), .CE(n3558), .R(n1750), .D(n1903), .Q(_zyGfifoF26_L530_req_0));
Q_FDP4EP _zyGfifoF27_L480_req_0_REG  ( .CK(clk), .CE(n34), .R(n1750), .D(n1904), .Q(_zyGfifoF27_L480_req_0));
Q_FDP4EP _zyGfifoF28_L482_req_0_REG  ( .CK(clk), .CE(n33), .R(n1750), .D(n1905), .Q(_zyGfifoF28_L482_req_0));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[63] ( .CK(clk), .CE(n33), .R(n1750), .D(n3072), .Q(_zyGfifoF28_L482_data_0[63]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[62] ( .CK(clk), .CE(n33), .R(n1750), .D(n3071), .Q(_zyGfifoF28_L482_data_0[62]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[61] ( .CK(clk), .CE(n33), .R(n1750), .D(n3070), .Q(_zyGfifoF28_L482_data_0[61]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[60] ( .CK(clk), .CE(n33), .R(n1750), .D(n3069), .Q(_zyGfifoF28_L482_data_0[60]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[59] ( .CK(clk), .CE(n33), .R(n1750), .D(n3068), .Q(_zyGfifoF28_L482_data_0[59]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[58] ( .CK(clk), .CE(n33), .R(n1750), .D(n3067), .Q(_zyGfifoF28_L482_data_0[58]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[57] ( .CK(clk), .CE(n33), .R(n1750), .D(n3066), .Q(_zyGfifoF28_L482_data_0[57]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[56] ( .CK(clk), .CE(n33), .R(n1750), .D(n3065), .Q(_zyGfifoF28_L482_data_0[56]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[55] ( .CK(clk), .CE(n33), .R(n1750), .D(n3064), .Q(_zyGfifoF28_L482_data_0[55]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[54] ( .CK(clk), .CE(n33), .R(n1750), .D(n3063), .Q(_zyGfifoF28_L482_data_0[54]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[53] ( .CK(clk), .CE(n33), .R(n1750), .D(n3062), .Q(_zyGfifoF28_L482_data_0[53]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[52] ( .CK(clk), .CE(n33), .R(n1750), .D(n3061), .Q(_zyGfifoF28_L482_data_0[52]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[51] ( .CK(clk), .CE(n33), .R(n1750), .D(n3060), .Q(_zyGfifoF28_L482_data_0[51]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[50] ( .CK(clk), .CE(n33), .R(n1750), .D(n3059), .Q(_zyGfifoF28_L482_data_0[50]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[49] ( .CK(clk), .CE(n33), .R(n1750), .D(n3058), .Q(_zyGfifoF28_L482_data_0[49]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[48] ( .CK(clk), .CE(n33), .R(n1750), .D(n3057), .Q(_zyGfifoF28_L482_data_0[48]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[47] ( .CK(clk), .CE(n33), .R(n1750), .D(n3056), .Q(_zyGfifoF28_L482_data_0[47]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[46] ( .CK(clk), .CE(n33), .R(n1750), .D(n3055), .Q(_zyGfifoF28_L482_data_0[46]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[45] ( .CK(clk), .CE(n33), .R(n1750), .D(n3054), .Q(_zyGfifoF28_L482_data_0[45]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[44] ( .CK(clk), .CE(n33), .R(n1750), .D(n3053), .Q(_zyGfifoF28_L482_data_0[44]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[43] ( .CK(clk), .CE(n33), .R(n1750), .D(n3052), .Q(_zyGfifoF28_L482_data_0[43]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[42] ( .CK(clk), .CE(n33), .R(n1750), .D(n3051), .Q(_zyGfifoF28_L482_data_0[42]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[41] ( .CK(clk), .CE(n33), .R(n1750), .D(n3050), .Q(_zyGfifoF28_L482_data_0[41]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[40] ( .CK(clk), .CE(n33), .R(n1750), .D(n3049), .Q(_zyGfifoF28_L482_data_0[40]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[39] ( .CK(clk), .CE(n33), .R(n1750), .D(n3048), .Q(_zyGfifoF28_L482_data_0[39]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[38] ( .CK(clk), .CE(n33), .R(n1750), .D(n3047), .Q(_zyGfifoF28_L482_data_0[38]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[37] ( .CK(clk), .CE(n33), .R(n1750), .D(n3046), .Q(_zyGfifoF28_L482_data_0[37]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[36] ( .CK(clk), .CE(n33), .R(n1750), .D(n3045), .Q(_zyGfifoF28_L482_data_0[36]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[35] ( .CK(clk), .CE(n33), .R(n1750), .D(n3044), .Q(_zyGfifoF28_L482_data_0[35]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[34] ( .CK(clk), .CE(n33), .R(n1750), .D(n3043), .Q(_zyGfifoF28_L482_data_0[34]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[33] ( .CK(clk), .CE(n33), .R(n1750), .D(n3042), .Q(_zyGfifoF28_L482_data_0[33]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[32] ( .CK(clk), .CE(n33), .R(n1750), .D(n3041), .Q(_zyGfifoF28_L482_data_0[32]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[31] ( .CK(clk), .CE(n33), .R(n1750), .D(n3040), .Q(_zyGfifoF28_L482_data_0[31]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[30] ( .CK(clk), .CE(n33), .R(n1750), .D(n3039), .Q(_zyGfifoF28_L482_data_0[30]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[29] ( .CK(clk), .CE(n33), .R(n1750), .D(n3038), .Q(_zyGfifoF28_L482_data_0[29]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[28] ( .CK(clk), .CE(n33), .R(n1750), .D(n3037), .Q(_zyGfifoF28_L482_data_0[28]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[27] ( .CK(clk), .CE(n33), .R(n1750), .D(n3036), .Q(_zyGfifoF28_L482_data_0[27]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[26] ( .CK(clk), .CE(n33), .R(n1750), .D(n3035), .Q(_zyGfifoF28_L482_data_0[26]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[25] ( .CK(clk), .CE(n33), .R(n1750), .D(n3034), .Q(_zyGfifoF28_L482_data_0[25]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[24] ( .CK(clk), .CE(n33), .R(n1750), .D(n3033), .Q(_zyGfifoF28_L482_data_0[24]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[23] ( .CK(clk), .CE(n33), .R(n1750), .D(n3032), .Q(_zyGfifoF28_L482_data_0[23]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[22] ( .CK(clk), .CE(n33), .R(n1750), .D(n3031), .Q(_zyGfifoF28_L482_data_0[22]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[21] ( .CK(clk), .CE(n33), .R(n1750), .D(n3030), .Q(_zyGfifoF28_L482_data_0[21]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[20] ( .CK(clk), .CE(n33), .R(n1750), .D(n3029), .Q(_zyGfifoF28_L482_data_0[20]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[19] ( .CK(clk), .CE(n33), .R(n1750), .D(n3028), .Q(_zyGfifoF28_L482_data_0[19]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[18] ( .CK(clk), .CE(n33), .R(n1750), .D(n3027), .Q(_zyGfifoF28_L482_data_0[18]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[17] ( .CK(clk), .CE(n33), .R(n1750), .D(n3026), .Q(_zyGfifoF28_L482_data_0[17]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[16] ( .CK(clk), .CE(n33), .R(n1750), .D(n3025), .Q(_zyGfifoF28_L482_data_0[16]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[15] ( .CK(clk), .CE(n33), .R(n1750), .D(n3024), .Q(_zyGfifoF28_L482_data_0[15]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[14] ( .CK(clk), .CE(n33), .R(n1750), .D(n3023), .Q(_zyGfifoF28_L482_data_0[14]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[13] ( .CK(clk), .CE(n33), .R(n1750), .D(n3022), .Q(_zyGfifoF28_L482_data_0[13]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[12] ( .CK(clk), .CE(n33), .R(n1750), .D(n3021), .Q(_zyGfifoF28_L482_data_0[12]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[11] ( .CK(clk), .CE(n33), .R(n1750), .D(n3020), .Q(_zyGfifoF28_L482_data_0[11]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[10] ( .CK(clk), .CE(n33), .R(n1750), .D(n3019), .Q(_zyGfifoF28_L482_data_0[10]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[9] ( .CK(clk), .CE(n33), .R(n1750), .D(n3018), .Q(_zyGfifoF28_L482_data_0[9]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[8] ( .CK(clk), .CE(n33), .R(n1750), .D(n3017), .Q(_zyGfifoF28_L482_data_0[8]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[7] ( .CK(clk), .CE(n33), .R(n1750), .D(n3016), .Q(_zyGfifoF28_L482_data_0[7]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[6] ( .CK(clk), .CE(n33), .R(n1750), .D(n3015), .Q(_zyGfifoF28_L482_data_0[6]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[5] ( .CK(clk), .CE(n33), .R(n1750), .D(n3014), .Q(_zyGfifoF28_L482_data_0[5]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[4] ( .CK(clk), .CE(n33), .R(n1750), .D(n3013), .Q(_zyGfifoF28_L482_data_0[4]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[3] ( .CK(clk), .CE(n33), .R(n1750), .D(n3012), .Q(_zyGfifoF28_L482_data_0[3]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[2] ( .CK(clk), .CE(n33), .R(n1750), .D(n3011), .Q(_zyGfifoF28_L482_data_0[2]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[1] ( .CK(clk), .CE(n33), .R(n1750), .D(n3010), .Q(_zyGfifoF28_L482_data_0[1]));
Q_FDP4EP \_zyGfifoF28_L482_data_0_REG[0] ( .CK(clk), .CE(n33), .R(n1750), .D(n3009), .Q(_zyGfifoF28_L482_data_0[0]));
Q_FDP4EP _zyGfifoF29_L487_req_0_REG  ( .CK(clk), .CE(n32), .R(n1750), .D(n1906), .Q(_zyGfifoF29_L487_req_0));
Q_FDP4EP _zyGfifoF30_L491_req_0_REG  ( .CK(clk), .CE(n31), .R(n1750), .D(n1907), .Q(_zyGfifoF30_L491_req_0));
Q_FDP4EP \_zyGfifoF30_L491_data_0_REG[7] ( .CK(clk), .CE(n31), .R(n1750), .D(n3008), .Q(_zyGfifoF30_L491_data_0[7]));
Q_FDP4EP \_zyGfifoF30_L491_data_0_REG[6] ( .CK(clk), .CE(n31), .R(n1750), .D(n3007), .Q(_zyGfifoF30_L491_data_0[6]));
Q_FDP4EP \_zyGfifoF30_L491_data_0_REG[5] ( .CK(clk), .CE(n31), .R(n1750), .D(n3006), .Q(_zyGfifoF30_L491_data_0[5]));
Q_FDP4EP \_zyGfifoF30_L491_data_0_REG[4] ( .CK(clk), .CE(n31), .R(n1750), .D(n3005), .Q(_zyGfifoF30_L491_data_0[4]));
Q_FDP4EP \_zyGfifoF30_L491_data_0_REG[3] ( .CK(clk), .CE(n31), .R(n1750), .D(n3004), .Q(_zyGfifoF30_L491_data_0[3]));
Q_FDP4EP \_zyGfifoF30_L491_data_0_REG[2] ( .CK(clk), .CE(n31), .R(n1750), .D(n3003), .Q(_zyGfifoF30_L491_data_0[2]));
Q_FDP4EP \_zyGfifoF30_L491_data_0_REG[1] ( .CK(clk), .CE(n31), .R(n1750), .D(n3002), .Q(_zyGfifoF30_L491_data_0[1]));
Q_FDP4EP \_zyGfifoF30_L491_data_0_REG[0] ( .CK(clk), .CE(n31), .R(n1750), .D(n3001), .Q(_zyGfifoF30_L491_data_0[0]));
Q_FDP4EP _zyGfifoF31_L496_req_0_REG  ( .CK(clk), .CE(n30), .R(n1750), .D(n1908), .Q(_zyGfifoF31_L496_req_0));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[63] ( .CK(clk), .CE(n26), .R(n1750), .D(n1972), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [63]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[62] ( .CK(clk), .CE(n26), .R(n1750), .D(n1971), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [62]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[61] ( .CK(clk), .CE(n26), .R(n1750), .D(n1970), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [61]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[60] ( .CK(clk), .CE(n26), .R(n1750), .D(n1969), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [60]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[59] ( .CK(clk), .CE(n26), .R(n1750), .D(n1968), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [59]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[58] ( .CK(clk), .CE(n26), .R(n1750), .D(n1967), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [58]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[57] ( .CK(clk), .CE(n26), .R(n1750), .D(n1966), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [57]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[56] ( .CK(clk), .CE(n26), .R(n1750), .D(n1965), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [56]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[55] ( .CK(clk), .CE(n26), .R(n1750), .D(n1964), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [55]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[54] ( .CK(clk), .CE(n26), .R(n1750), .D(n1963), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [54]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[53] ( .CK(clk), .CE(n26), .R(n1750), .D(n1962), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [53]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[52] ( .CK(clk), .CE(n26), .R(n1750), .D(n1961), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [52]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[51] ( .CK(clk), .CE(n26), .R(n1750), .D(n1960), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [51]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[50] ( .CK(clk), .CE(n26), .R(n1750), .D(n1959), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [50]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[49] ( .CK(clk), .CE(n26), .R(n1750), .D(n1958), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [49]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[48] ( .CK(clk), .CE(n26), .R(n1750), .D(n1957), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [48]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[47] ( .CK(clk), .CE(n26), .R(n1750), .D(n1956), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [47]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[46] ( .CK(clk), .CE(n26), .R(n1750), .D(n1955), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [46]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[45] ( .CK(clk), .CE(n26), .R(n1750), .D(n1954), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [45]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[44] ( .CK(clk), .CE(n26), .R(n1750), .D(n1953), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [44]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[43] ( .CK(clk), .CE(n26), .R(n1750), .D(n1952), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [43]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[42] ( .CK(clk), .CE(n26), .R(n1750), .D(n1951), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [42]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[41] ( .CK(clk), .CE(n26), .R(n1750), .D(n1950), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [41]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[40] ( .CK(clk), .CE(n26), .R(n1750), .D(n1949), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [40]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[39] ( .CK(clk), .CE(n26), .R(n1750), .D(n1948), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [39]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[38] ( .CK(clk), .CE(n26), .R(n1750), .D(n1947), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [38]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[37] ( .CK(clk), .CE(n26), .R(n1750), .D(n1946), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [37]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[36] ( .CK(clk), .CE(n26), .R(n1750), .D(n1945), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [36]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[35] ( .CK(clk), .CE(n26), .R(n1750), .D(n1944), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [35]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[34] ( .CK(clk), .CE(n26), .R(n1750), .D(n1943), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [34]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[33] ( .CK(clk), .CE(n26), .R(n1750), .D(n1942), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [33]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[32] ( .CK(clk), .CE(n26), .R(n1750), .D(n1941), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [32]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[31] ( .CK(clk), .CE(n26), .R(n1750), .D(n1940), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [31]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[30] ( .CK(clk), .CE(n26), .R(n1750), .D(n1939), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [30]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[29] ( .CK(clk), .CE(n26), .R(n1750), .D(n1938), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [29]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[28] ( .CK(clk), .CE(n26), .R(n1750), .D(n1937), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [28]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[27] ( .CK(clk), .CE(n26), .R(n1750), .D(n1936), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [27]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[26] ( .CK(clk), .CE(n26), .R(n1750), .D(n1935), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [26]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[25] ( .CK(clk), .CE(n26), .R(n1750), .D(n1934), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [25]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[24] ( .CK(clk), .CE(n26), .R(n1750), .D(n1933), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [24]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[23] ( .CK(clk), .CE(n26), .R(n1750), .D(n1932), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [23]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[22] ( .CK(clk), .CE(n26), .R(n1750), .D(n1931), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [22]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[21] ( .CK(clk), .CE(n26), .R(n1750), .D(n1930), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [21]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[20] ( .CK(clk), .CE(n26), .R(n1750), .D(n1929), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [20]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[19] ( .CK(clk), .CE(n26), .R(n1750), .D(n1928), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [19]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[18] ( .CK(clk), .CE(n26), .R(n1750), .D(n1927), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [18]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[17] ( .CK(clk), .CE(n26), .R(n1750), .D(n1926), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [17]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[16] ( .CK(clk), .CE(n26), .R(n1750), .D(n1925), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [16]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[15] ( .CK(clk), .CE(n26), .R(n1750), .D(n1924), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [15]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[14] ( .CK(clk), .CE(n26), .R(n1750), .D(n1923), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [14]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[13] ( .CK(clk), .CE(n26), .R(n1750), .D(n1922), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [13]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[12] ( .CK(clk), .CE(n26), .R(n1750), .D(n1921), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [12]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[11] ( .CK(clk), .CE(n26), .R(n1750), .D(n1920), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [11]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[10] ( .CK(clk), .CE(n26), .R(n1750), .D(n1919), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [10]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[9] ( .CK(clk), .CE(n26), .R(n1750), .D(n1918), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [9]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[8] ( .CK(clk), .CE(n26), .R(n1750), .D(n1917), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [8]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[7] ( .CK(clk), .CE(n26), .R(n1750), .D(n1916), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [7]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[6] ( .CK(clk), .CE(n26), .R(n1750), .D(n1915), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [6]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[5] ( .CK(clk), .CE(n26), .R(n1750), .D(n1914), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [5]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[4] ( .CK(clk), .CE(n26), .R(n1750), .D(n1913), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [4]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[3] ( .CK(clk), .CE(n26), .R(n1750), .D(n1912), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [3]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[2] ( .CK(clk), .CE(n26), .R(n1750), .D(n1911), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [2]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[1] ( .CK(clk), .CE(n26), .R(n1750), .D(n1910), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [1]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11_REG[0] ( .CK(clk), .CE(n26), .R(n1750), .D(n1909), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytdata_L209_tfiV11 [0]));
Q_FDP4EP \tdata_ob_REG[63] ( .CK(clk), .CE(n26), .R(n1750), .D(n1972), .Q(tdata_ob[63]));
Q_FDP4EP \tdata_ob_REG[62] ( .CK(clk), .CE(n26), .R(n1750), .D(n1971), .Q(tdata_ob[62]));
Q_FDP4EP \tdata_ob_REG[61] ( .CK(clk), .CE(n26), .R(n1750), .D(n1970), .Q(tdata_ob[61]));
Q_FDP4EP \tdata_ob_REG[60] ( .CK(clk), .CE(n26), .R(n1750), .D(n1969), .Q(tdata_ob[60]));
Q_FDP4EP \tdata_ob_REG[59] ( .CK(clk), .CE(n26), .R(n1750), .D(n1968), .Q(tdata_ob[59]));
Q_FDP4EP \tdata_ob_REG[58] ( .CK(clk), .CE(n26), .R(n1750), .D(n1967), .Q(tdata_ob[58]));
Q_FDP4EP \tdata_ob_REG[57] ( .CK(clk), .CE(n26), .R(n1750), .D(n1966), .Q(tdata_ob[57]));
Q_FDP4EP \tdata_ob_REG[56] ( .CK(clk), .CE(n26), .R(n1750), .D(n1965), .Q(tdata_ob[56]));
Q_FDP4EP \tdata_ob_REG[55] ( .CK(clk), .CE(n26), .R(n1750), .D(n1964), .Q(tdata_ob[55]));
Q_FDP4EP \tdata_ob_REG[54] ( .CK(clk), .CE(n26), .R(n1750), .D(n1963), .Q(tdata_ob[54]));
Q_FDP4EP \tdata_ob_REG[53] ( .CK(clk), .CE(n26), .R(n1750), .D(n1962), .Q(tdata_ob[53]));
Q_FDP4EP \tdata_ob_REG[52] ( .CK(clk), .CE(n26), .R(n1750), .D(n1961), .Q(tdata_ob[52]));
Q_FDP4EP \tdata_ob_REG[51] ( .CK(clk), .CE(n26), .R(n1750), .D(n1960), .Q(tdata_ob[51]));
Q_FDP4EP \tdata_ob_REG[50] ( .CK(clk), .CE(n26), .R(n1750), .D(n1959), .Q(tdata_ob[50]));
Q_FDP4EP \tdata_ob_REG[49] ( .CK(clk), .CE(n26), .R(n1750), .D(n1958), .Q(tdata_ob[49]));
Q_FDP4EP \tdata_ob_REG[48] ( .CK(clk), .CE(n26), .R(n1750), .D(n1957), .Q(tdata_ob[48]));
Q_FDP4EP \tdata_ob_REG[47] ( .CK(clk), .CE(n26), .R(n1750), .D(n1956), .Q(tdata_ob[47]));
Q_FDP4EP \tdata_ob_REG[46] ( .CK(clk), .CE(n26), .R(n1750), .D(n1955), .Q(tdata_ob[46]));
Q_FDP4EP \tdata_ob_REG[45] ( .CK(clk), .CE(n26), .R(n1750), .D(n1954), .Q(tdata_ob[45]));
Q_FDP4EP \tdata_ob_REG[44] ( .CK(clk), .CE(n26), .R(n1750), .D(n1953), .Q(tdata_ob[44]));
Q_FDP4EP \tdata_ob_REG[43] ( .CK(clk), .CE(n26), .R(n1750), .D(n1952), .Q(tdata_ob[43]));
Q_FDP4EP \tdata_ob_REG[42] ( .CK(clk), .CE(n26), .R(n1750), .D(n1951), .Q(tdata_ob[42]));
Q_FDP4EP \tdata_ob_REG[41] ( .CK(clk), .CE(n26), .R(n1750), .D(n1950), .Q(tdata_ob[41]));
Q_FDP4EP \tdata_ob_REG[40] ( .CK(clk), .CE(n26), .R(n1750), .D(n1949), .Q(tdata_ob[40]));
Q_FDP4EP \tdata_ob_REG[39] ( .CK(clk), .CE(n26), .R(n1750), .D(n1948), .Q(tdata_ob[39]));
Q_FDP4EP \tdata_ob_REG[38] ( .CK(clk), .CE(n26), .R(n1750), .D(n1947), .Q(tdata_ob[38]));
Q_FDP4EP \tdata_ob_REG[37] ( .CK(clk), .CE(n26), .R(n1750), .D(n1946), .Q(tdata_ob[37]));
Q_FDP4EP \tdata_ob_REG[36] ( .CK(clk), .CE(n26), .R(n1750), .D(n1945), .Q(tdata_ob[36]));
Q_FDP4EP \tdata_ob_REG[35] ( .CK(clk), .CE(n26), .R(n1750), .D(n1944), .Q(tdata_ob[35]));
Q_FDP4EP \tdata_ob_REG[34] ( .CK(clk), .CE(n26), .R(n1750), .D(n1943), .Q(tdata_ob[34]));
Q_FDP4EP \tdata_ob_REG[33] ( .CK(clk), .CE(n26), .R(n1750), .D(n1942), .Q(tdata_ob[33]));
Q_FDP4EP \tdata_ob_REG[32] ( .CK(clk), .CE(n26), .R(n1750), .D(n1941), .Q(tdata_ob[32]));
Q_FDP4EP \tdata_ob_REG[31] ( .CK(clk), .CE(n26), .R(n1750), .D(n1940), .Q(tdata_ob[31]));
Q_FDP4EP \tdata_ob_REG[30] ( .CK(clk), .CE(n26), .R(n1750), .D(n1939), .Q(tdata_ob[30]));
Q_FDP4EP \tdata_ob_REG[29] ( .CK(clk), .CE(n26), .R(n1750), .D(n1938), .Q(tdata_ob[29]));
Q_FDP4EP \tdata_ob_REG[28] ( .CK(clk), .CE(n26), .R(n1750), .D(n1937), .Q(tdata_ob[28]));
Q_FDP4EP \tdata_ob_REG[27] ( .CK(clk), .CE(n26), .R(n1750), .D(n1936), .Q(tdata_ob[27]));
Q_FDP4EP \tdata_ob_REG[26] ( .CK(clk), .CE(n26), .R(n1750), .D(n1935), .Q(tdata_ob[26]));
Q_FDP4EP \tdata_ob_REG[25] ( .CK(clk), .CE(n26), .R(n1750), .D(n1934), .Q(tdata_ob[25]));
Q_FDP4EP \tdata_ob_REG[24] ( .CK(clk), .CE(n26), .R(n1750), .D(n1933), .Q(tdata_ob[24]));
Q_FDP4EP \tdata_ob_REG[23] ( .CK(clk), .CE(n26), .R(n1750), .D(n1932), .Q(tdata_ob[23]));
Q_FDP4EP \tdata_ob_REG[22] ( .CK(clk), .CE(n26), .R(n1750), .D(n1931), .Q(tdata_ob[22]));
Q_FDP4EP \tdata_ob_REG[21] ( .CK(clk), .CE(n26), .R(n1750), .D(n1930), .Q(tdata_ob[21]));
Q_FDP4EP \tdata_ob_REG[20] ( .CK(clk), .CE(n26), .R(n1750), .D(n1929), .Q(tdata_ob[20]));
Q_FDP4EP \tdata_ob_REG[19] ( .CK(clk), .CE(n26), .R(n1750), .D(n1928), .Q(tdata_ob[19]));
Q_FDP4EP \tdata_ob_REG[18] ( .CK(clk), .CE(n26), .R(n1750), .D(n1927), .Q(tdata_ob[18]));
Q_FDP4EP \tdata_ob_REG[17] ( .CK(clk), .CE(n26), .R(n1750), .D(n1926), .Q(tdata_ob[17]));
Q_FDP4EP \tdata_ob_REG[16] ( .CK(clk), .CE(n26), .R(n1750), .D(n1925), .Q(tdata_ob[16]));
Q_FDP4EP \tdata_ob_REG[15] ( .CK(clk), .CE(n26), .R(n1750), .D(n1924), .Q(tdata_ob[15]));
Q_FDP4EP \tdata_ob_REG[14] ( .CK(clk), .CE(n26), .R(n1750), .D(n1923), .Q(tdata_ob[14]));
Q_FDP4EP \tdata_ob_REG[13] ( .CK(clk), .CE(n26), .R(n1750), .D(n1922), .Q(tdata_ob[13]));
Q_FDP4EP \tdata_ob_REG[12] ( .CK(clk), .CE(n26), .R(n1750), .D(n1921), .Q(tdata_ob[12]));
Q_FDP4EP \tdata_ob_REG[11] ( .CK(clk), .CE(n26), .R(n1750), .D(n1920), .Q(tdata_ob[11]));
Q_FDP4EP \tdata_ob_REG[10] ( .CK(clk), .CE(n26), .R(n1750), .D(n1919), .Q(tdata_ob[10]));
Q_FDP4EP \tdata_ob_REG[9] ( .CK(clk), .CE(n26), .R(n1750), .D(n1918), .Q(tdata_ob[9]));
Q_FDP4EP \tdata_ob_REG[8] ( .CK(clk), .CE(n26), .R(n1750), .D(n1917), .Q(tdata_ob[8]));
Q_FDP4EP \tdata_ob_REG[7] ( .CK(clk), .CE(n26), .R(n1750), .D(n1916), .Q(tdata_ob[7]));
Q_FDP4EP \tdata_ob_REG[6] ( .CK(clk), .CE(n26), .R(n1750), .D(n1915), .Q(tdata_ob[6]));
Q_FDP4EP \tdata_ob_REG[5] ( .CK(clk), .CE(n26), .R(n1750), .D(n1914), .Q(tdata_ob[5]));
Q_FDP4EP \tdata_ob_REG[4] ( .CK(clk), .CE(n26), .R(n1750), .D(n1913), .Q(tdata_ob[4]));
Q_FDP4EP \tdata_ob_REG[3] ( .CK(clk), .CE(n26), .R(n1750), .D(n1912), .Q(tdata_ob[3]));
Q_INV U7828 ( .A(tdata_ob[3]), .Z(n1776));
Q_FDP4EP \tdata_ob_REG[2] ( .CK(clk), .CE(n26), .R(n1750), .D(n1911), .Q(tdata_ob[2]));
Q_FDP4EP \tdata_ob_REG[1] ( .CK(clk), .CE(n26), .R(n1750), .D(n1910), .Q(tdata_ob[1]));
Q_FDP4EP \tdata_ob_REG[0] ( .CK(clk), .CE(n26), .R(n1750), .D(n1909), .Q(tdata_ob[0]));
Q_INV U7832 ( .A(tdata_ob[0]), .Z(n1775));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[31] ( .CK(clk), .CE(n26), .R(n1750), .D(n2108), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [31]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[30] ( .CK(clk), .CE(n26), .R(n1750), .D(n2107), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [30]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[29] ( .CK(clk), .CE(n26), .R(n1750), .D(n2106), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [29]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[28] ( .CK(clk), .CE(n26), .R(n1750), .D(n2105), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [28]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[27] ( .CK(clk), .CE(n26), .R(n1750), .D(n2104), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [27]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[26] ( .CK(clk), .CE(n26), .R(n1750), .D(n2103), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [26]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[25] ( .CK(clk), .CE(n26), .R(n1750), .D(n2102), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [25]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[24] ( .CK(clk), .CE(n26), .R(n1750), .D(n2101), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [24]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[23] ( .CK(clk), .CE(n26), .R(n1750), .D(n2100), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [23]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[22] ( .CK(clk), .CE(n26), .R(n1750), .D(n2099), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [22]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[21] ( .CK(clk), .CE(n26), .R(n1750), .D(n2098), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [21]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[20] ( .CK(clk), .CE(n26), .R(n1750), .D(n2097), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [20]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[19] ( .CK(clk), .CE(n26), .R(n1750), .D(n2096), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [19]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[18] ( .CK(clk), .CE(n26), .R(n1750), .D(n2095), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [18]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[17] ( .CK(clk), .CE(n26), .R(n1750), .D(n2094), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [17]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[16] ( .CK(clk), .CE(n26), .R(n1750), .D(n2093), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [16]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[15] ( .CK(clk), .CE(n26), .R(n1750), .D(n2092), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [15]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[14] ( .CK(clk), .CE(n26), .R(n1750), .D(n2091), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [14]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[13] ( .CK(clk), .CE(n26), .R(n1750), .D(n2090), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [13]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[12] ( .CK(clk), .CE(n26), .R(n1750), .D(n2089), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [12]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[11] ( .CK(clk), .CE(n26), .R(n1750), .D(n2088), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [11]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[10] ( .CK(clk), .CE(n26), .R(n1750), .D(n2087), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [10]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[9] ( .CK(clk), .CE(n26), .R(n1750), .D(n2086), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [9]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[8] ( .CK(clk), .CE(n26), .R(n1750), .D(n2085), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [8]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[7] ( .CK(clk), .CE(n26), .R(n1750), .D(n2084), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [7]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[6] ( .CK(clk), .CE(n26), .R(n1750), .D(n2083), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [6]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[5] ( .CK(clk), .CE(n26), .R(n1750), .D(n2082), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [5]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[4] ( .CK(clk), .CE(n26), .R(n1750), .D(n2081), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [4]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[3] ( .CK(clk), .CE(n26), .R(n1750), .D(n2080), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [3]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[2] ( .CK(clk), .CE(n26), .R(n1750), .D(n2079), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [2]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[1] ( .CK(clk), .CE(n26), .R(n1750), .D(n2078), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [1]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12_REG[0] ( .CK(clk), .CE(n26), .R(n1750), .D(n2077), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytuser_string_L209_tfiV12 [0]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[31] ( .CK(clk), .CE(n26), .R(n1750), .D(n2182), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [31]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[30] ( .CK(clk), .CE(n26), .R(n1750), .D(n2181), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [30]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[29] ( .CK(clk), .CE(n26), .R(n1750), .D(n2180), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [29]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[28] ( .CK(clk), .CE(n26), .R(n1750), .D(n2179), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [28]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[27] ( .CK(clk), .CE(n26), .R(n1750), .D(n2178), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [27]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[26] ( .CK(clk), .CE(n26), .R(n1750), .D(n2177), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [26]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[25] ( .CK(clk), .CE(n26), .R(n1750), .D(n2176), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [25]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[24] ( .CK(clk), .CE(n26), .R(n1750), .D(n2175), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [24]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[23] ( .CK(clk), .CE(n26), .R(n1750), .D(n2174), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [23]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[22] ( .CK(clk), .CE(n26), .R(n1750), .D(n2173), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [22]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[21] ( .CK(clk), .CE(n26), .R(n1750), .D(n2172), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [21]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[20] ( .CK(clk), .CE(n26), .R(n1750), .D(n2171), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [20]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[19] ( .CK(clk), .CE(n26), .R(n1750), .D(n2170), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [19]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[18] ( .CK(clk), .CE(n26), .R(n1750), .D(n2169), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [18]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[17] ( .CK(clk), .CE(n26), .R(n1750), .D(n2168), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [17]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[16] ( .CK(clk), .CE(n26), .R(n1750), .D(n2167), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [16]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[15] ( .CK(clk), .CE(n26), .R(n1750), .D(n2166), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [15]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[14] ( .CK(clk), .CE(n26), .R(n1750), .D(n2165), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [14]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[13] ( .CK(clk), .CE(n26), .R(n1750), .D(n2164), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [13]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[12] ( .CK(clk), .CE(n26), .R(n1750), .D(n2163), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [12]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[11] ( .CK(clk), .CE(n26), .R(n1750), .D(n2162), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [11]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[10] ( .CK(clk), .CE(n26), .R(n1750), .D(n2161), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [10]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[9] ( .CK(clk), .CE(n26), .R(n1750), .D(n2160), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [9]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[8] ( .CK(clk), .CE(n26), .R(n1750), .D(n2159), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [8]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[7] ( .CK(clk), .CE(n26), .R(n1750), .D(n2158), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [7]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[6] ( .CK(clk), .CE(n26), .R(n1750), .D(n2157), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [6]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[5] ( .CK(clk), .CE(n26), .R(n1750), .D(n2156), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [5]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[4] ( .CK(clk), .CE(n26), .R(n1750), .D(n2155), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [4]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[3] ( .CK(clk), .CE(n26), .R(n1750), .D(n2154), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [3]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[2] ( .CK(clk), .CE(n26), .R(n1750), .D(n2153), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [2]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[1] ( .CK(clk), .CE(n26), .R(n1750), .D(n2152), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [1]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14_REG[0] ( .CK(clk), .CE(n26), .R(n1750), .D(n2151), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zystr_get_L209_tfiV14 [0]));
Q_FDP4EP \tuser_string_ob_REG[31] ( .CK(clk), .CE(n26), .R(n1750), .D(n2108), .Q(tuser_string_ob[31]));
Q_FDP4EP \tuser_string_ob_REG[30] ( .CK(clk), .CE(n26), .R(n1750), .D(n2107), .Q(tuser_string_ob[30]));
Q_FDP4EP \tuser_string_ob_REG[29] ( .CK(clk), .CE(n26), .R(n1750), .D(n2106), .Q(tuser_string_ob[29]));
Q_FDP4EP \tuser_string_ob_REG[28] ( .CK(clk), .CE(n26), .R(n1750), .D(n2105), .Q(tuser_string_ob[28]));
Q_FDP4EP \tuser_string_ob_REG[27] ( .CK(clk), .CE(n26), .R(n1750), .D(n2104), .Q(tuser_string_ob[27]));
Q_FDP4EP \tuser_string_ob_REG[26] ( .CK(clk), .CE(n26), .R(n1750), .D(n2103), .Q(tuser_string_ob[26]));
Q_FDP4EP \tuser_string_ob_REG[25] ( .CK(clk), .CE(n26), .R(n1750), .D(n2102), .Q(tuser_string_ob[25]));
Q_FDP4EP \tuser_string_ob_REG[24] ( .CK(clk), .CE(n26), .R(n1750), .D(n2101), .Q(tuser_string_ob[24]));
Q_FDP4EP \tuser_string_ob_REG[23] ( .CK(clk), .CE(n26), .R(n1750), .D(n2100), .Q(tuser_string_ob[23]));
Q_FDP4EP \tuser_string_ob_REG[22] ( .CK(clk), .CE(n26), .R(n1750), .D(n2099), .Q(tuser_string_ob[22]));
Q_FDP4EP \tuser_string_ob_REG[21] ( .CK(clk), .CE(n26), .R(n1750), .D(n2098), .Q(tuser_string_ob[21]));
Q_FDP4EP \tuser_string_ob_REG[20] ( .CK(clk), .CE(n26), .R(n1750), .D(n2097), .Q(tuser_string_ob[20]));
Q_FDP4EP \tuser_string_ob_REG[19] ( .CK(clk), .CE(n26), .R(n1750), .D(n2096), .Q(tuser_string_ob[19]));
Q_FDP4EP \tuser_string_ob_REG[18] ( .CK(clk), .CE(n26), .R(n1750), .D(n2095), .Q(tuser_string_ob[18]));
Q_FDP4EP \tuser_string_ob_REG[17] ( .CK(clk), .CE(n26), .R(n1750), .D(n2094), .Q(tuser_string_ob[17]));
Q_FDP4EP \tuser_string_ob_REG[16] ( .CK(clk), .CE(n26), .R(n1750), .D(n2093), .Q(tuser_string_ob[16]));
Q_FDP4EP \tuser_string_ob_REG[15] ( .CK(clk), .CE(n26), .R(n1750), .D(n2092), .Q(tuser_string_ob[15]));
Q_FDP4EP \tuser_string_ob_REG[14] ( .CK(clk), .CE(n26), .R(n1750), .D(n2091), .Q(tuser_string_ob[14]));
Q_FDP4EP \tuser_string_ob_REG[13] ( .CK(clk), .CE(n26), .R(n1750), .D(n2090), .Q(tuser_string_ob[13]));
Q_FDP4EP \tuser_string_ob_REG[12] ( .CK(clk), .CE(n26), .R(n1750), .D(n2089), .Q(tuser_string_ob[12]));
Q_FDP4EP \tuser_string_ob_REG[11] ( .CK(clk), .CE(n26), .R(n1750), .D(n2088), .Q(tuser_string_ob[11]));
Q_FDP4EP \tuser_string_ob_REG[10] ( .CK(clk), .CE(n26), .R(n1750), .D(n2087), .Q(tuser_string_ob[10]));
Q_FDP4EP \tuser_string_ob_REG[9] ( .CK(clk), .CE(n26), .R(n1750), .D(n2086), .Q(tuser_string_ob[9]));
Q_FDP4EP \tuser_string_ob_REG[8] ( .CK(clk), .CE(n26), .R(n1750), .D(n2085), .Q(tuser_string_ob[8]));
Q_FDP4EP \tuser_string_ob_REG[7] ( .CK(clk), .CE(n26), .R(n1750), .D(n2084), .Q(tuser_string_ob[7]));
Q_FDP4EP \tuser_string_ob_REG[6] ( .CK(clk), .CE(n26), .R(n1750), .D(n2083), .Q(tuser_string_ob[6]));
Q_FDP4EP \tuser_string_ob_REG[5] ( .CK(clk), .CE(n26), .R(n1750), .D(n2082), .Q(tuser_string_ob[5]));
Q_FDP4EP \tuser_string_ob_REG[4] ( .CK(clk), .CE(n26), .R(n1750), .D(n2081), .Q(tuser_string_ob[4]));
Q_FDP4EP \tuser_string_ob_REG[3] ( .CK(clk), .CE(n26), .R(n1750), .D(n2080), .Q(tuser_string_ob[3]));
Q_FDP4EP \tuser_string_ob_REG[2] ( .CK(clk), .CE(n26), .R(n1750), .D(n2079), .Q(tuser_string_ob[2]));
Q_FDP4EP \tuser_string_ob_REG[1] ( .CK(clk), .CE(n26), .R(n1750), .D(n2078), .Q(tuser_string_ob[1]));
Q_FDP4EP \tuser_string_ob_REG[0] ( .CK(clk), .CE(n26), .R(n1750), .D(n2077), .Q(tuser_string_ob[0]));
Q_FDP4EP \str_get_ob_REG[31] ( .CK(clk), .CE(n26), .R(n1750), .D(n2182), .Q(str_get_ob[31]));
Q_FDP4EP \str_get_ob_REG[30] ( .CK(clk), .CE(n26), .R(n1750), .D(n2181), .Q(str_get_ob[30]));
Q_FDP4EP \str_get_ob_REG[29] ( .CK(clk), .CE(n26), .R(n1750), .D(n2180), .Q(str_get_ob[29]));
Q_FDP4EP \str_get_ob_REG[28] ( .CK(clk), .CE(n26), .R(n1750), .D(n2179), .Q(str_get_ob[28]));
Q_FDP4EP \str_get_ob_REG[27] ( .CK(clk), .CE(n26), .R(n1750), .D(n2178), .Q(str_get_ob[27]));
Q_FDP4EP \str_get_ob_REG[26] ( .CK(clk), .CE(n26), .R(n1750), .D(n2177), .Q(str_get_ob[26]));
Q_FDP4EP \str_get_ob_REG[25] ( .CK(clk), .CE(n26), .R(n1750), .D(n2176), .Q(str_get_ob[25]));
Q_FDP4EP \str_get_ob_REG[24] ( .CK(clk), .CE(n26), .R(n1750), .D(n2175), .Q(str_get_ob[24]));
Q_FDP4EP \str_get_ob_REG[23] ( .CK(clk), .CE(n26), .R(n1750), .D(n2174), .Q(str_get_ob[23]));
Q_FDP4EP \str_get_ob_REG[22] ( .CK(clk), .CE(n26), .R(n1750), .D(n2173), .Q(str_get_ob[22]));
Q_FDP4EP \str_get_ob_REG[21] ( .CK(clk), .CE(n26), .R(n1750), .D(n2172), .Q(str_get_ob[21]));
Q_FDP4EP \str_get_ob_REG[20] ( .CK(clk), .CE(n26), .R(n1750), .D(n2171), .Q(str_get_ob[20]));
Q_FDP4EP \str_get_ob_REG[19] ( .CK(clk), .CE(n26), .R(n1750), .D(n2170), .Q(str_get_ob[19]));
Q_FDP4EP \str_get_ob_REG[18] ( .CK(clk), .CE(n26), .R(n1750), .D(n2169), .Q(str_get_ob[18]));
Q_FDP4EP \str_get_ob_REG[17] ( .CK(clk), .CE(n26), .R(n1750), .D(n2168), .Q(str_get_ob[17]));
Q_FDP4EP \str_get_ob_REG[16] ( .CK(clk), .CE(n26), .R(n1750), .D(n2167), .Q(str_get_ob[16]));
Q_FDP4EP \str_get_ob_REG[15] ( .CK(clk), .CE(n26), .R(n1750), .D(n2166), .Q(str_get_ob[15]));
Q_FDP4EP \str_get_ob_REG[14] ( .CK(clk), .CE(n26), .R(n1750), .D(n2165), .Q(str_get_ob[14]));
Q_FDP4EP \str_get_ob_REG[13] ( .CK(clk), .CE(n26), .R(n1750), .D(n2164), .Q(str_get_ob[13]));
Q_FDP4EP \str_get_ob_REG[12] ( .CK(clk), .CE(n26), .R(n1750), .D(n2163), .Q(str_get_ob[12]));
Q_FDP4EP \str_get_ob_REG[11] ( .CK(clk), .CE(n26), .R(n1750), .D(n2162), .Q(str_get_ob[11]));
Q_FDP4EP \str_get_ob_REG[10] ( .CK(clk), .CE(n26), .R(n1750), .D(n2161), .Q(str_get_ob[10]));
Q_FDP4EP \str_get_ob_REG[9] ( .CK(clk), .CE(n26), .R(n1750), .D(n2160), .Q(str_get_ob[9]));
Q_FDP4EP \str_get_ob_REG[8] ( .CK(clk), .CE(n26), .R(n1750), .D(n2159), .Q(str_get_ob[8]));
Q_FDP4EP \str_get_ob_REG[7] ( .CK(clk), .CE(n26), .R(n1750), .D(n2158), .Q(str_get_ob[7]));
Q_FDP4EP \str_get_ob_REG[6] ( .CK(clk), .CE(n26), .R(n1750), .D(n2157), .Q(str_get_ob[6]));
Q_FDP4EP \str_get_ob_REG[5] ( .CK(clk), .CE(n26), .R(n1750), .D(n2156), .Q(str_get_ob[5]));
Q_FDP4EP \str_get_ob_REG[4] ( .CK(clk), .CE(n26), .R(n1750), .D(n2155), .Q(str_get_ob[4]));
Q_FDP4EP \str_get_ob_REG[3] ( .CK(clk), .CE(n26), .R(n1750), .D(n2154), .Q(str_get_ob[3]));
Q_FDP4EP \str_get_ob_REG[2] ( .CK(clk), .CE(n26), .R(n1750), .D(n2153), .Q(str_get_ob[2]));
Q_FDP4EP \str_get_ob_REG[1] ( .CK(clk), .CE(n26), .R(n1750), .D(n2152), .Q(str_get_ob[1]));
Q_INV U7960 ( .A(str_get_ob[1]), .Z(n1758));
Q_FDP4EP \str_get_ob_REG[0] ( .CK(clk), .CE(n26), .R(n1750), .D(n2151), .Q(str_get_ob[0]));
Q_INV U7962 ( .A(str_get_ob[0]), .Z(n1757));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytstrb_L209_tfiV13_REG[7] ( .CK(clk), .CE(n26), .R(n1750), .D(n2138), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytstrb_L209_tfiV13 [7]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytstrb_L209_tfiV13_REG[6] ( .CK(clk), .CE(n26), .R(n1750), .D(n2137), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytstrb_L209_tfiV13 [6]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytstrb_L209_tfiV13_REG[5] ( .CK(clk), .CE(n26), .R(n1750), .D(n2136), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytstrb_L209_tfiV13 [5]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytstrb_L209_tfiV13_REG[4] ( .CK(clk), .CE(n26), .R(n1750), .D(n2135), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytstrb_L209_tfiV13 [4]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytstrb_L209_tfiV13_REG[3] ( .CK(clk), .CE(n26), .R(n1750), .D(n2134), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytstrb_L209_tfiV13 [3]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytstrb_L209_tfiV13_REG[2] ( .CK(clk), .CE(n26), .R(n1750), .D(n2133), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytstrb_L209_tfiV13 [2]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytstrb_L209_tfiV13_REG[1] ( .CK(clk), .CE(n26), .R(n1750), .D(n2132), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytstrb_L209_tfiV13 [1]));
Q_FDP4EP \_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytstrb_L209_tfiV13_REG[0] ( .CK(clk), .CE(n26), .R(n1750), .D(n2131), .Q(\_zyL439_meSwitch8._zygfifotfiCscp2_L441_ob_service_data_isf_meScp9._zytstrb_L209_tfiV13 [0]));
Q_FDP4EP \tstrb_ob_REG[7] ( .CK(clk), .CE(n26), .R(n1750), .D(n2138), .Q(tstrb_ob[7]));
Q_FDP4EP \tstrb_ob_REG[6] ( .CK(clk), .CE(n26), .R(n1750), .D(n2137), .Q(tstrb_ob[6]));
Q_FDP4EP \tstrb_ob_REG[5] ( .CK(clk), .CE(n26), .R(n1750), .D(n2136), .Q(tstrb_ob[5]));
Q_FDP4EP \tstrb_ob_REG[4] ( .CK(clk), .CE(n26), .R(n1750), .D(n2135), .Q(tstrb_ob[4]));
Q_FDP4EP \tstrb_ob_REG[3] ( .CK(clk), .CE(n26), .R(n1750), .D(n2134), .Q(tstrb_ob[3]));
Q_FDP4EP \tstrb_ob_REG[2] ( .CK(clk), .CE(n26), .R(n1750), .D(n2133), .Q(tstrb_ob[2]));
Q_FDP4EP \tstrb_ob_REG[1] ( .CK(clk), .CE(n26), .R(n1750), .D(n2132), .Q(tstrb_ob[1]));
Q_FDP4EP \tstrb_ob_REG[0] ( .CK(clk), .CE(n26), .R(n1750), .D(n2131), .Q(tstrb_ob[0]));
Q_FDP4EP \_zygsfis_ob_service_data_rptr_REG[4] ( .CK(clk), .CE(n26), .R(n1750), .D(n2405), .Q(_zygsfis_ob_service_data_rptr[4]));
Q_FDP4EP \_zygsfis_ob_service_data_rptr_REG[3] ( .CK(clk), .CE(n26), .R(n1750), .D(n2404), .Q(_zygsfis_ob_service_data_rptr[3]));
Q_FDP4EP \_zygsfis_ob_service_data_rptr_REG[2] ( .CK(clk), .CE(n26), .R(n1750), .D(n2403), .Q(_zygsfis_ob_service_data_rptr[2]));
Q_FDP4EP \_zygsfis_ob_service_data_rptr_REG[1] ( .CK(clk), .CE(n26), .R(n1750), .D(n2402), .Q(_zygsfis_ob_service_data_rptr[1]));
Q_FDP4EP \_zygsfis_ob_service_data_rptr_REG[0] ( .CK(clk), .CE(n26), .R(n1750), .D(n2401), .Q(_zygsfis_ob_service_data_rptr[0]));
Q_FDP4EP \_zygsfis_ob_service_data_space_REG[4] ( .CK(clk), .CE(n26), .R(n1750), .D(n3200), .Q(_zygsfis_ob_service_data_space[4]));
Q_FDP4EP \_zygsfis_ob_service_data_space_REG[3] ( .CK(clk), .CE(n26), .R(n1750), .D(n3198), .Q(_zygsfis_ob_service_data_space[3]));
Q_FDP4EP \_zygsfis_ob_service_data_space_REG[2] ( .CK(clk), .CE(n26), .R(n1750), .D(n3196), .Q(_zygsfis_ob_service_data_space[2]));
Q_FDP4EP \_zygsfis_ob_service_data_space_REG[1] ( .CK(clk), .CE(n26), .R(n1750), .D(n3194), .Q(_zygsfis_ob_service_data_space[1]));
Q_FDP4EP \_zygsfis_ob_service_data_space_REG[0] ( .CK(clk), .CE(n26), .R(n1750), .D(n3192), .Q(_zygsfis_ob_service_data_space[0]));
Q_INV U7989 ( .A(n3352), .Z(n24));
Q_FDP4EP \_zyL439_meState8_REG[1] ( .CK(clk), .CE(n24), .R(n1750), .D(n3273), .Q(_zyL439_meState8[1]));
Q_INV U7991 ( .A(_zyL439_meState8[1]), .Z(n3272));
Q_FDP4EP \_zyL439_meState8_REG[0] ( .CK(clk), .CE(n24), .R(n1750), .D(n3552), .Q(_zyL439_meState8[0]));
Q_INV U7993 ( .A(_zyL439_meState8[0]), .Z(n2465));
Q_FDP4EP \_zyL443_tfiRv7_REG[24] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL443_tfiRv7[24]));
Q_FDP4EP \_zyL443_tfiRv7_REG[23] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL443_tfiRv7[23]));
Q_FDP4EP \_zyL443_tfiRv7_REG[22] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(_zyL443_tfiRv7[22]));
Q_FDP4EP \_zyL443_tfiRv7_REG[21] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL443_tfiRv7[21]));
Q_FDP4EP \_zyL443_tfiRv7_REG[20] ( .CK(clk), .CE(n26), .R(n1750), .D(n3537), .Q(_zyL443_tfiRv7[20]));
Q_FDP4EP \_zyL443_tfiRv7_REG[19] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL443_tfiRv7[19]));
Q_FDP4EP \_zyL443_tfiRv7_REG[18] ( .CK(clk), .CE(n26), .R(n1750), .D(n3536), .Q(_zyL443_tfiRv7[18]));
Q_FDP4EP \_zyL443_tfiRv7_REG[17] ( .CK(clk), .CE(n26), .R(n1750), .D(n3537), .Q(_zyL443_tfiRv7[17]));
Q_FDP4EP \_zyL443_tfiRv7_REG[16] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(_zyL443_tfiRv7[16]));
Q_FDP4EP \_zyL443_tfiRv7_REG[15] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL443_tfiRv7[15]));
Q_FDP4EP \_zyL443_tfiRv7_REG[14] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(_zyL443_tfiRv7[14]));
Q_FDP4EP \_zyL443_tfiRv7_REG[13] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(_zyL443_tfiRv7[13]));
Q_FDP4EP \_zyL443_tfiRv7_REG[12] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL443_tfiRv7[12]));
Q_FDP4EP \_zyL443_tfiRv7_REG[11] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(_zyL443_tfiRv7[11]));
Q_FDP4EP \_zyL443_tfiRv7_REG[10] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(_zyL443_tfiRv7[10]));
Q_FDP4EP \_zyL443_tfiRv7_REG[9] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(_zyL443_tfiRv7[9]));
Q_FDP4EP \_zyL443_tfiRv7_REG[8] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(_zyL443_tfiRv7[8]));
Q_FDP4EP \_zyL443_tfiRv7_REG[7] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL443_tfiRv7[7]));
Q_FDP4EP \_zyL443_tfiRv7_REG[6] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(_zyL443_tfiRv7[6]));
Q_FDP4EP \_zyL443_tfiRv7_REG[5] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL443_tfiRv7[5]));
Q_FDP4EP \_zyL443_tfiRv7_REG[4] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(_zyL443_tfiRv7[4]));
Q_FDP4EP \_zyL443_tfiRv7_REG[3] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL443_tfiRv7[3]));
Q_FDP4EP \_zyL443_tfiRv7_REG[2] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(_zyL443_tfiRv7[2]));
Q_FDP4EP \_zyL443_tfiRv7_REG[1] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL443_tfiRv7[1]));
Q_FDP4EP \_zyL443_tfiRv7_REG[0] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL443_tfiRv7[0]));
Q_FDP4EP \user_string_ob_REG[24] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(user_string_ob[24]));
Q_FDP4EP \user_string_ob_REG[23] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(user_string_ob[23]));
Q_FDP4EP \user_string_ob_REG[22] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(user_string_ob[22]));
Q_INV U8022 ( .A(user_string_ob[22]), .Z(n3335));
Q_FDP4EP \user_string_ob_REG[21] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(user_string_ob[21]));
Q_FDP4EP \user_string_ob_REG[20] ( .CK(clk), .CE(n26), .R(n1750), .D(n3537), .Q(user_string_ob[20]));
Q_FDP4EP \user_string_ob_REG[19] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(user_string_ob[19]));
Q_FDP4EP \user_string_ob_REG[18] ( .CK(clk), .CE(n26), .R(n1750), .D(n3536), .Q(user_string_ob[18]));
Q_INV U8027 ( .A(user_string_ob[18]), .Z(n3263));
Q_FDP4EP \user_string_ob_REG[17] ( .CK(clk), .CE(n26), .R(n1750), .D(n3537), .Q(user_string_ob[17]));
Q_FDP4EP \user_string_ob_REG[16] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(user_string_ob[16]));
Q_INV U8030 ( .A(user_string_ob[16]), .Z(n3258));
Q_FDP4EP \user_string_ob_REG[15] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(user_string_ob[15]));
Q_FDP4EP \user_string_ob_REG[14] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(user_string_ob[14]));
Q_INV U8033 ( .A(user_string_ob[14]), .Z(n3389));
Q_FDP4EP \user_string_ob_REG[13] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(user_string_ob[13]));
Q_FDP4EP \user_string_ob_REG[12] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(user_string_ob[12]));
Q_FDP4EP \user_string_ob_REG[11] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(user_string_ob[11]));
Q_FDP4EP \user_string_ob_REG[10] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(user_string_ob[10]));
Q_INV U8038 ( .A(user_string_ob[10]), .Z(n3259));
Q_FDP4EP \user_string_ob_REG[9] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(user_string_ob[9]));
Q_INV U8040 ( .A(user_string_ob[9]), .Z(n3388));
Q_FDP4EP \user_string_ob_REG[8] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(user_string_ob[8]));
Q_INV U8042 ( .A(user_string_ob[8]), .Z(n3332));
Q_FDP4EP \user_string_ob_REG[7] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(user_string_ob[7]));
Q_FDP4EP \user_string_ob_REG[6] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(user_string_ob[6]));
Q_FDP4EP \user_string_ob_REG[5] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(user_string_ob[5]));
Q_FDP4EP \user_string_ob_REG[4] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(user_string_ob[4]));
Q_FDP4EP \user_string_ob_REG[3] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(user_string_ob[3]));
Q_FDP4EP \user_string_ob_REG[2] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(user_string_ob[2]));
Q_INV U8049 ( .A(user_string_ob[2]), .Z(n3336));
Q_FDP4EP \user_string_ob_REG[1] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(user_string_ob[1]));
Q_FDP4EP \user_string_ob_REG[0] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(user_string_ob[0]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[31] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyGfifoF23_L444_data_0[31]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[30] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyGfifoF23_L444_data_0[30]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[29] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyGfifoF23_L444_data_0[29]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[28] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyGfifoF23_L444_data_0[28]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[27] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyGfifoF23_L444_data_0[27]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[26] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyGfifoF23_L444_data_0[26]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[25] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyGfifoF23_L444_data_0[25]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[24] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyGfifoF23_L444_data_0[24]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[23] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyGfifoF23_L444_data_0[23]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[22] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(_zyGfifoF23_L444_data_0[22]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[21] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyGfifoF23_L444_data_0[21]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[20] ( .CK(clk), .CE(n26), .R(n1750), .D(n3537), .Q(_zyGfifoF23_L444_data_0[20]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[19] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyGfifoF23_L444_data_0[19]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[18] ( .CK(clk), .CE(n26), .R(n1750), .D(n3536), .Q(_zyGfifoF23_L444_data_0[18]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[17] ( .CK(clk), .CE(n26), .R(n1750), .D(n3537), .Q(_zyGfifoF23_L444_data_0[17]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[16] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(_zyGfifoF23_L444_data_0[16]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[15] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyGfifoF23_L444_data_0[15]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[14] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(_zyGfifoF23_L444_data_0[14]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[13] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(_zyGfifoF23_L444_data_0[13]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[12] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyGfifoF23_L444_data_0[12]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[11] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(_zyGfifoF23_L444_data_0[11]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[10] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(_zyGfifoF23_L444_data_0[10]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[9] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(_zyGfifoF23_L444_data_0[9]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[8] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(_zyGfifoF23_L444_data_0[8]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[7] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyGfifoF23_L444_data_0[7]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[6] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(_zyGfifoF23_L444_data_0[6]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[5] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyGfifoF23_L444_data_0[5]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[4] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(_zyGfifoF23_L444_data_0[4]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[3] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyGfifoF23_L444_data_0[3]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[2] ( .CK(clk), .CE(n26), .R(n1750), .D(n3201), .Q(_zyGfifoF23_L444_data_0[2]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[1] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyGfifoF23_L444_data_0[1]));
Q_FDP4EP \_zyGfifoF23_L444_data_0_REG[0] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyGfifoF23_L444_data_0[0]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[31] ( .CK(clk), .CE(n3558), .R(n1750), .D(n1750), .Q(_zyGfifoF26_L530_data_0[31]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[30] ( .CK(clk), .CE(n3558), .R(n1750), .D(n1750), .Q(_zyGfifoF26_L530_data_0[30]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[29] ( .CK(clk), .CE(n3558), .R(n1750), .D(n1750), .Q(_zyGfifoF26_L530_data_0[29]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[28] ( .CK(clk), .CE(n3558), .R(n1750), .D(n1750), .Q(_zyGfifoF26_L530_data_0[28]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[27] ( .CK(clk), .CE(n3558), .R(n1750), .D(n1750), .Q(_zyGfifoF26_L530_data_0[27]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[26] ( .CK(clk), .CE(n3558), .R(n1750), .D(n1750), .Q(_zyGfifoF26_L530_data_0[26]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[25] ( .CK(clk), .CE(n3558), .R(n1750), .D(n1750), .Q(_zyGfifoF26_L530_data_0[25]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[24] ( .CK(clk), .CE(n3558), .R(n1750), .D(n3243), .Q(_zyGfifoF26_L530_data_0[24]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[23] ( .CK(clk), .CE(n3558), .R(n1750), .D(n3242), .Q(_zyGfifoF26_L530_data_0[23]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[22] ( .CK(clk), .CE(n3558), .R(n1750), .D(n3241), .Q(_zyGfifoF26_L530_data_0[22]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[21] ( .CK(clk), .CE(n3558), .R(n1750), .D(n3240), .Q(_zyGfifoF26_L530_data_0[21]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[20] ( .CK(clk), .CE(n3558), .R(n1750), .D(n3239), .Q(_zyGfifoF26_L530_data_0[20]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[19] ( .CK(clk), .CE(n3558), .R(n1750), .D(n3238), .Q(_zyGfifoF26_L530_data_0[19]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[18] ( .CK(clk), .CE(n3558), .R(n1750), .D(n3237), .Q(_zyGfifoF26_L530_data_0[18]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[17] ( .CK(clk), .CE(n3558), .R(n1750), .D(n3236), .Q(_zyGfifoF26_L530_data_0[17]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[16] ( .CK(clk), .CE(n3558), .R(n1750), .D(n3235), .Q(_zyGfifoF26_L530_data_0[16]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[15] ( .CK(clk), .CE(n3558), .R(n1750), .D(n3234), .Q(_zyGfifoF26_L530_data_0[15]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[14] ( .CK(clk), .CE(n3558), .R(n1750), .D(n3233), .Q(_zyGfifoF26_L530_data_0[14]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[13] ( .CK(clk), .CE(n3558), .R(n1750), .D(n3232), .Q(_zyGfifoF26_L530_data_0[13]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[12] ( .CK(clk), .CE(n3558), .R(n1750), .D(n3231), .Q(_zyGfifoF26_L530_data_0[12]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[11] ( .CK(clk), .CE(n3558), .R(n1750), .D(n3230), .Q(_zyGfifoF26_L530_data_0[11]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[10] ( .CK(clk), .CE(n3558), .R(n1750), .D(n3229), .Q(_zyGfifoF26_L530_data_0[10]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[9] ( .CK(clk), .CE(n3558), .R(n1750), .D(n3228), .Q(_zyGfifoF26_L530_data_0[9]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[8] ( .CK(clk), .CE(n3558), .R(n1750), .D(n3227), .Q(_zyGfifoF26_L530_data_0[8]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[7] ( .CK(clk), .CE(n3558), .R(n1750), .D(n3226), .Q(_zyGfifoF26_L530_data_0[7]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[6] ( .CK(clk), .CE(n3558), .R(n1750), .D(n3225), .Q(_zyGfifoF26_L530_data_0[6]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[5] ( .CK(clk), .CE(n3558), .R(n1750), .D(n3224), .Q(_zyGfifoF26_L530_data_0[5]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[4] ( .CK(clk), .CE(n3558), .R(n1750), .D(n3223), .Q(_zyGfifoF26_L530_data_0[4]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[3] ( .CK(clk), .CE(n3558), .R(n1750), .D(n3222), .Q(_zyGfifoF26_L530_data_0[3]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[2] ( .CK(clk), .CE(n3558), .R(n1750), .D(n3221), .Q(_zyGfifoF26_L530_data_0[2]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[1] ( .CK(clk), .CE(n3558), .R(n1750), .D(n3220), .Q(_zyGfifoF26_L530_data_0[1]));
Q_FDP4EP \_zyGfifoF26_L530_data_0_REG[0] ( .CK(clk), .CE(n3558), .R(n1750), .D(n3219), .Q(_zyGfifoF26_L530_data_0[0]));
Q_FDP4EP \_zyGfifoF27_L480_data_0_REG[7] ( .CK(clk), .CE(n34), .R(n1750), .D(n1750), .Q(_zyGfifoF27_L480_data_0[7]));
Q_FDP4EP \_zyGfifoF27_L480_data_0_REG[6] ( .CK(clk), .CE(n34), .R(n1750), .D(n1750), .Q(_zyGfifoF27_L480_data_0[6]));
Q_FDP4EP \_zyGfifoF27_L480_data_0_REG[5] ( .CK(clk), .CE(n34), .R(n1750), .D(n1750), .Q(_zyGfifoF27_L480_data_0[5]));
Q_FDP4EP \_zyGfifoF27_L480_data_0_REG[4] ( .CK(clk), .CE(n34), .R(n1750), .D(n1750), .Q(_zyGfifoF27_L480_data_0[4]));
Q_FDP4EP \_zyGfifoF27_L480_data_0_REG[3] ( .CK(clk), .CE(n34), .R(n1750), .D(n1750), .Q(_zyGfifoF27_L480_data_0[3]));
Q_FDP4EP \_zyGfifoF27_L480_data_0_REG[2] ( .CK(clk), .CE(n34), .R(n1750), .D(n1750), .Q(_zyGfifoF27_L480_data_0[2]));
Q_FDP4EP \_zyGfifoF27_L480_data_0_REG[1] ( .CK(clk), .CE(n34), .R(n1750), .D(n3245), .Q(_zyGfifoF27_L480_data_0[1]));
Q_FDP4EP \_zyGfifoF27_L480_data_0_REG[0] ( .CK(clk), .CE(n34), .R(n1750), .D(n3244), .Q(_zyGfifoF27_L480_data_0[0]));
Q_FDP4EP \_zyGfifoF29_L487_data_0_REG[7] ( .CK(clk), .CE(n32), .R(n1750), .D(n1750), .Q(_zyGfifoF29_L487_data_0[7]));
Q_FDP4EP \_zyGfifoF29_L487_data_0_REG[6] ( .CK(clk), .CE(n32), .R(n1750), .D(n1750), .Q(_zyGfifoF29_L487_data_0[6]));
Q_FDP4EP \_zyGfifoF29_L487_data_0_REG[5] ( .CK(clk), .CE(n32), .R(n1750), .D(n1750), .Q(_zyGfifoF29_L487_data_0[5]));
Q_FDP4EP \_zyGfifoF29_L487_data_0_REG[4] ( .CK(clk), .CE(n32), .R(n1750), .D(n1750), .Q(_zyGfifoF29_L487_data_0[4]));
Q_FDP4EP \_zyGfifoF29_L487_data_0_REG[3] ( .CK(clk), .CE(n32), .R(n1750), .D(n1750), .Q(_zyGfifoF29_L487_data_0[3]));
Q_FDP4EP \_zyGfifoF29_L487_data_0_REG[2] ( .CK(clk), .CE(n32), .R(n1750), .D(n1750), .Q(_zyGfifoF29_L487_data_0[2]));
Q_FDP4EP \_zyGfifoF29_L487_data_0_REG[1] ( .CK(clk), .CE(n32), .R(n1750), .D(n3245), .Q(_zyGfifoF29_L487_data_0[1]));
Q_FDP4EP \_zyGfifoF29_L487_data_0_REG[0] ( .CK(clk), .CE(n32), .R(n1750), .D(n3244), .Q(_zyGfifoF29_L487_data_0[0]));
Q_FDP4EP \_zyGfifoF31_L496_data_0_REG[0] ( .CK(clk), .CE(n30), .R(n1750), .D(n3218), .Q(_zyGfifoF31_L496_data_0[0]));
Q_FDP4EP tlast_REG  ( .CK(clk), .CE(n34), .R(n1750), .D(n3218), .Q(tlast));
Q_FDP4EP ignore_compare_result_REG  ( .CK(clk), .CE(n34), .R(n1750), .D(n3217), .Q(ignore_compare_result));
Q_FDP4EP \_zyL441_tfiRv19_REG[31] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[31]));
Q_FDP4EP \_zyL441_tfiRv19_REG[30] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[30]));
Q_FDP4EP \_zyL441_tfiRv19_REG[29] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[29]));
Q_FDP4EP \_zyL441_tfiRv19_REG[28] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[28]));
Q_FDP4EP \_zyL441_tfiRv19_REG[27] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[27]));
Q_FDP4EP \_zyL441_tfiRv19_REG[26] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[26]));
Q_FDP4EP \_zyL441_tfiRv19_REG[25] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[25]));
Q_FDP4EP \_zyL441_tfiRv19_REG[24] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[24]));
Q_FDP4EP \_zyL441_tfiRv19_REG[23] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[23]));
Q_FDP4EP \_zyL441_tfiRv19_REG[22] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[22]));
Q_FDP4EP \_zyL441_tfiRv19_REG[21] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[21]));
Q_FDP4EP \_zyL441_tfiRv19_REG[20] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[20]));
Q_FDP4EP \_zyL441_tfiRv19_REG[19] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[19]));
Q_FDP4EP \_zyL441_tfiRv19_REG[18] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[18]));
Q_FDP4EP \_zyL441_tfiRv19_REG[17] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[17]));
Q_FDP4EP \_zyL441_tfiRv19_REG[16] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[16]));
Q_FDP4EP \_zyL441_tfiRv19_REG[15] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[15]));
Q_FDP4EP \_zyL441_tfiRv19_REG[14] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[14]));
Q_FDP4EP \_zyL441_tfiRv19_REG[13] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[13]));
Q_FDP4EP \_zyL441_tfiRv19_REG[12] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[12]));
Q_FDP4EP \_zyL441_tfiRv19_REG[11] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[11]));
Q_FDP4EP \_zyL441_tfiRv19_REG[10] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[10]));
Q_FDP4EP \_zyL441_tfiRv19_REG[9] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[9]));
Q_FDP4EP \_zyL441_tfiRv19_REG[8] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[8]));
Q_FDP4EP \_zyL441_tfiRv19_REG[7] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[7]));
Q_FDP4EP \_zyL441_tfiRv19_REG[6] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[6]));
Q_FDP4EP \_zyL441_tfiRv19_REG[5] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[5]));
Q_FDP4EP \_zyL441_tfiRv19_REG[4] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[4]));
Q_FDP4EP \_zyL441_tfiRv19_REG[3] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[3]));
Q_FDP4EP \_zyL441_tfiRv19_REG[2] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(_zyL441_tfiRv19[2]));
Q_FDP4EP \_zyL441_tfiRv19_REG[1] ( .CK(clk), .CE(n26), .R(n1750), .D(n3557), .Q(_zyL441_tfiRv19[1]));
Q_FDP4EP \_zyL441_tfiRv19_REG[0] ( .CK(clk), .CE(n26), .R(n1750), .D(n3534), .Q(_zyL441_tfiRv19[0]));
Q_FDP4EP \retval_ob_REG[31] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[31]));
Q_FDP4EP \retval_ob_REG[30] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[30]));
Q_FDP4EP \retval_ob_REG[29] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[29]));
Q_FDP4EP \retval_ob_REG[28] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[28]));
Q_FDP4EP \retval_ob_REG[27] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[27]));
Q_FDP4EP \retval_ob_REG[26] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[26]));
Q_FDP4EP \retval_ob_REG[25] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[25]));
Q_FDP4EP \retval_ob_REG[24] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[24]));
Q_FDP4EP \retval_ob_REG[23] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[23]));
Q_FDP4EP \retval_ob_REG[22] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[22]));
Q_FDP4EP \retval_ob_REG[21] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[21]));
Q_FDP4EP \retval_ob_REG[20] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[20]));
Q_FDP4EP \retval_ob_REG[19] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[19]));
Q_FDP4EP \retval_ob_REG[18] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[18]));
Q_FDP4EP \retval_ob_REG[17] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[17]));
Q_FDP4EP \retval_ob_REG[16] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[16]));
Q_FDP4EP \retval_ob_REG[15] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[15]));
Q_FDP4EP \retval_ob_REG[14] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[14]));
Q_FDP4EP \retval_ob_REG[13] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[13]));
Q_FDP4EP \retval_ob_REG[12] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[12]));
Q_FDP4EP \retval_ob_REG[11] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[11]));
Q_FDP4EP \retval_ob_REG[10] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[10]));
Q_FDP4EP \retval_ob_REG[9] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[9]));
Q_FDP4EP \retval_ob_REG[8] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[8]));
Q_FDP4EP \retval_ob_REG[7] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[7]));
Q_FDP4EP \retval_ob_REG[6] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[6]));
Q_FDP4EP \retval_ob_REG[5] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[5]));
Q_FDP4EP \retval_ob_REG[4] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[4]));
Q_FDP4EP \retval_ob_REG[3] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[3]));
Q_FDP4EP \retval_ob_REG[2] ( .CK(clk), .CE(n26), .R(n1750), .D(n1750), .Q(retval_ob[2]));
Q_FDP4EP \retval_ob_REG[1] ( .CK(clk), .CE(n26), .R(n1750), .D(n3557), .Q(retval_ob[1]));
Q_FDP4EP \retval_ob_REG[0] ( .CK(clk), .CE(n26), .R(n1750), .D(n3534), .Q(retval_ob[0]));
Q_FDP4EP \_zyL462_tfiRv8_REG[7] ( .CK(clk), .CE(n3558), .R(n1750), .D(n1750), .Q(_zyL462_tfiRv8[7]));
Q_FDP4EP \_zyL462_tfiRv8_REG[6] ( .CK(clk), .CE(n3558), .R(n1750), .D(n1750), .Q(_zyL462_tfiRv8[6]));
Q_FDP4EP \_zyL462_tfiRv8_REG[5] ( .CK(clk), .CE(n3558), .R(n1750), .D(n1750), .Q(_zyL462_tfiRv8[5]));
Q_FDP4EP \_zyL462_tfiRv8_REG[4] ( .CK(clk), .CE(n3558), .R(n1750), .D(n1750), .Q(_zyL462_tfiRv8[4]));
Q_FDP4EP \_zyL462_tfiRv8_REG[3] ( .CK(clk), .CE(n3558), .R(n1750), .D(n1750), .Q(_zyL462_tfiRv8[3]));
Q_FDP4EP \_zyL462_tfiRv8_REG[2] ( .CK(clk), .CE(n3558), .R(n1750), .D(n1750), .Q(_zyL462_tfiRv8[2]));
Q_FDP4EP \_zyL462_tfiRv8_REG[1] ( .CK(clk), .CE(n3558), .R(n1750), .D(n3247), .Q(_zyL462_tfiRv8[1]));
Q_FDP4EP \_zyL462_tfiRv8_REG[0] ( .CK(clk), .CE(n3558), .R(n1750), .D(n3246), .Q(_zyL462_tfiRv8[0]));
Q_FDP4EP \tuser_REG[7] ( .CK(clk), .CE(n34), .R(n1750), .D(n1750), .Q(tuser[7]));
Q_FDP4EP \tuser_REG[6] ( .CK(clk), .CE(n34), .R(n1750), .D(n1750), .Q(tuser[6]));
Q_FDP4EP \tuser_REG[5] ( .CK(clk), .CE(n34), .R(n1750), .D(n1750), .Q(tuser[5]));
Q_FDP4EP \tuser_REG[4] ( .CK(clk), .CE(n34), .R(n1750), .D(n1750), .Q(tuser[4]));
Q_FDP4EP \tuser_REG[3] ( .CK(clk), .CE(n34), .R(n1750), .D(n1750), .Q(tuser[3]));
Q_FDP4EP \tuser_REG[2] ( .CK(clk), .CE(n34), .R(n1750), .D(n1750), .Q(tuser[2]));
Q_FDP4EP \tuser_REG[1] ( .CK(clk), .CE(n34), .R(n1750), .D(n3245), .Q(tuser[1]));
Q_FDP4EP \tuser_REG[0] ( .CK(clk), .CE(n34), .R(n1750), .D(n3244), .Q(tuser[0]));
Q_FDP4EP \kme_ib_tid_REG[0] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(kme_ib_tid[0]));
Q_FDP4EP kme_ob_tready_REG  ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n5382), .Q(kme_ob_tready));
Q_FDP4EP config_done_REG  ( .CK(_zyM2L253_pbcMevClk12), .CE(n5334), .R(n1750), .D(n5382), .Q(config_done));
Q_FDP4EP config_ready_REG  ( .CK(_zyM2L253_pbcMevClk12), .CE(n5335), .R(n1750), .D(n5382), .Q(config_ready));
Q_INV U8219 ( .A(config_ready), .Z(n1024));
Q_INV U8220 ( .A(n5295), .Z(n23));
Q_FDP4EP \_zz_58_258_2_REG[31] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[31]), .Q(_zz_58_258_2[31]));
Q_FDP4EP \_zz_58_258_2_REG[30] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[30]), .Q(_zz_58_258_2[30]));
Q_FDP4EP \_zz_58_258_2_REG[29] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[29]), .Q(_zz_58_258_2[29]));
Q_FDP4EP \_zz_58_258_2_REG[28] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[28]), .Q(_zz_58_258_2[28]));
Q_FDP4EP \_zz_58_258_2_REG[27] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[27]), .Q(_zz_58_258_2[27]));
Q_FDP4EP \_zz_58_258_2_REG[26] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[26]), .Q(_zz_58_258_2[26]));
Q_FDP4EP \_zz_58_258_2_REG[25] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[25]), .Q(_zz_58_258_2[25]));
Q_FDP4EP \_zz_58_258_2_REG[24] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[24]), .Q(_zz_58_258_2[24]));
Q_FDP4EP \_zz_58_258_2_REG[23] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[23]), .Q(_zz_58_258_2[23]));
Q_FDP4EP \_zz_58_258_2_REG[22] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[22]), .Q(_zz_58_258_2[22]));
Q_FDP4EP \_zz_58_258_2_REG[21] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[21]), .Q(_zz_58_258_2[21]));
Q_FDP4EP \_zz_58_258_2_REG[20] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[20]), .Q(_zz_58_258_2[20]));
Q_FDP4EP \_zz_58_258_2_REG[19] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[19]), .Q(_zz_58_258_2[19]));
Q_FDP4EP \_zz_58_258_2_REG[18] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[18]), .Q(_zz_58_258_2[18]));
Q_FDP4EP \_zz_58_258_2_REG[17] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[17]), .Q(_zz_58_258_2[17]));
Q_FDP4EP \_zz_58_258_2_REG[16] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[16]), .Q(_zz_58_258_2[16]));
Q_FDP4EP \_zz_58_258_2_REG[15] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[15]), .Q(_zz_58_258_2[15]));
Q_FDP4EP \_zz_58_258_2_REG[14] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[14]), .Q(_zz_58_258_2[14]));
Q_FDP4EP \_zz_58_258_2_REG[13] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[13]), .Q(_zz_58_258_2[13]));
Q_FDP4EP \_zz_58_258_2_REG[12] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[12]), .Q(_zz_58_258_2[12]));
Q_FDP4EP \_zz_58_258_2_REG[11] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[11]), .Q(_zz_58_258_2[11]));
Q_FDP4EP \_zz_58_258_2_REG[10] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[10]), .Q(_zz_58_258_2[10]));
Q_FDP4EP \_zz_58_258_2_REG[9] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[9]), .Q(_zz_58_258_2[9]));
Q_FDP4EP \_zz_58_258_2_REG[8] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[8]), .Q(_zz_58_258_2[8]));
Q_FDP4EP \_zz_58_258_2_REG[7] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[7]), .Q(_zz_58_258_2[7]));
Q_FDP4EP \_zz_58_258_2_REG[6] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[6]), .Q(_zz_58_258_2[6]));
Q_FDP4EP \_zz_58_258_2_REG[5] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[5]), .Q(_zz_58_258_2[5]));
Q_FDP4EP \_zz_58_258_2_REG[4] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[4]), .Q(_zz_58_258_2[4]));
Q_FDP4EP \_zz_58_258_2_REG[3] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[3]), .Q(_zz_58_258_2[3]));
Q_FDP4EP \_zz_58_258_2_REG[2] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[2]), .Q(_zz_58_258_2[2]));
Q_FDP4EP \_zz_58_258_2_REG[1] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[1]), .Q(_zz_58_258_2[1]));
Q_FDP4EP \_zz_58_258_2_REG[0] ( .CK(_zyM2L253_pbcMevClk12), .CE(n23), .R(n1750), .D(_zyictd_sysfunc_36_L258_1[0]), .Q(_zz_58_258_2[0]));
Q_INV U8253 ( .A(n5297), .Z(n22));
Q_FDP4EP \_zz_58_264_3_REG[31] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[31]), .Q(_zz_58_264_3[31]));
Q_FDP4EP \_zz_58_264_3_REG[30] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[30]), .Q(_zz_58_264_3[30]));
Q_FDP4EP \_zz_58_264_3_REG[29] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[29]), .Q(_zz_58_264_3[29]));
Q_FDP4EP \_zz_58_264_3_REG[28] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[28]), .Q(_zz_58_264_3[28]));
Q_FDP4EP \_zz_58_264_3_REG[27] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[27]), .Q(_zz_58_264_3[27]));
Q_FDP4EP \_zz_58_264_3_REG[26] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[26]), .Q(_zz_58_264_3[26]));
Q_FDP4EP \_zz_58_264_3_REG[25] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[25]), .Q(_zz_58_264_3[25]));
Q_FDP4EP \_zz_58_264_3_REG[24] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[24]), .Q(_zz_58_264_3[24]));
Q_FDP4EP \_zz_58_264_3_REG[23] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[23]), .Q(_zz_58_264_3[23]));
Q_FDP4EP \_zz_58_264_3_REG[22] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[22]), .Q(_zz_58_264_3[22]));
Q_FDP4EP \_zz_58_264_3_REG[21] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[21]), .Q(_zz_58_264_3[21]));
Q_FDP4EP \_zz_58_264_3_REG[20] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[20]), .Q(_zz_58_264_3[20]));
Q_FDP4EP \_zz_58_264_3_REG[19] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[19]), .Q(_zz_58_264_3[19]));
Q_FDP4EP \_zz_58_264_3_REG[18] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[18]), .Q(_zz_58_264_3[18]));
Q_FDP4EP \_zz_58_264_3_REG[17] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[17]), .Q(_zz_58_264_3[17]));
Q_FDP4EP \_zz_58_264_3_REG[16] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[16]), .Q(_zz_58_264_3[16]));
Q_FDP4EP \_zz_58_264_3_REG[15] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[15]), .Q(_zz_58_264_3[15]));
Q_FDP4EP \_zz_58_264_3_REG[14] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[14]), .Q(_zz_58_264_3[14]));
Q_FDP4EP \_zz_58_264_3_REG[13] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[13]), .Q(_zz_58_264_3[13]));
Q_FDP4EP \_zz_58_264_3_REG[12] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[12]), .Q(_zz_58_264_3[12]));
Q_FDP4EP \_zz_58_264_3_REG[11] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[11]), .Q(_zz_58_264_3[11]));
Q_FDP4EP \_zz_58_264_3_REG[10] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[10]), .Q(_zz_58_264_3[10]));
Q_FDP4EP \_zz_58_264_3_REG[9] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[9]), .Q(_zz_58_264_3[9]));
Q_FDP4EP \_zz_58_264_3_REG[8] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[8]), .Q(_zz_58_264_3[8]));
Q_FDP4EP \_zz_58_264_3_REG[7] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[7]), .Q(_zz_58_264_3[7]));
Q_FDP4EP \_zz_58_264_3_REG[6] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[6]), .Q(_zz_58_264_3[6]));
Q_FDP4EP \_zz_58_264_3_REG[5] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[5]), .Q(_zz_58_264_3[5]));
Q_FDP4EP \_zz_58_264_3_REG[4] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[4]), .Q(_zz_58_264_3[4]));
Q_FDP4EP \_zz_58_264_3_REG[3] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[3]), .Q(_zz_58_264_3[3]));
Q_FDP4EP \_zz_58_264_3_REG[2] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[2]), .Q(_zz_58_264_3[2]));
Q_FDP4EP \_zz_58_264_3_REG[1] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[1]), .Q(_zz_58_264_3[1]));
Q_FDP4EP \_zz_58_264_3_REG[0] ( .CK(_zyM2L253_pbcMevClk12), .CE(n22), .R(n1750), .D(_zyictd_sysfunc_36_L264_4[0]), .Q(_zz_58_264_3[0]));
Q_INV U8286 ( .A(n5300), .Z(n21));
Q_FDP4EP _zzM2L253_mdxP5_En_REG  ( .CK(_zyM2L253_pbcMevClk12), .CE(n21), .R(n1750), .D(_zzM2L253_mdxP5_EnNxt), .Q(_zzM2L253_mdxP5_En));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[31] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[31]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[30] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[30]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[29] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[29]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[28] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[28]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[27] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[27]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[26] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[26]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[25] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[25]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[24] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[24]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[23] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[23]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[22] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[22]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[21] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[21]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[20] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[20]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[19] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[19]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[18] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[18]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[17] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[17]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[16] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[16]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[15] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[15]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[14] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[14]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[13] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[13]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[12] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[12]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[11] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[11]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[10] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[10]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[9] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[9]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[8] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[8]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[7] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[7]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[6] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[6]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[5] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[5]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[4] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[4]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[3] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[3]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[2] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[2]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[1] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[1]));
Q_FDP4EP \_zzM2L253_mdxP5_error_cntr_wr0_REG[0] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_error_cntr_wr0[0]));
Q_FDP4EP _zzM2L253_mdxP5_kme_ib_tvalid_wr1_REG  ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tvalid_wr1));
Q_FDP4EP _zzM2L253_mdxP5_kme_ib_tlast_wr2_REG  ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tlast_wr2));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[63] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[63]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[62] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[62]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[61] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[61]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[60] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[60]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[59] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[59]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[58] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[58]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[57] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[57]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[56] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[56]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[55] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[55]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[54] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[54]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[53] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[53]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[52] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[52]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[51] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[51]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[50] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[50]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[49] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[49]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[48] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[48]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[47] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[47]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[46] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[46]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[45] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[45]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[44] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[44]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[43] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[43]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[42] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[42]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[41] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[41]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[40] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[40]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[39] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[39]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[38] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[38]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[37] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[37]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[36] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[36]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[35] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[35]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[34] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[34]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[33] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[33]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[32] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[32]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[31] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[31]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[30] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[30]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[29] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[29]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[28] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[28]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[27] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[27]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[26] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[26]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[25] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[25]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[24] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[24]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[23] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[23]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[22] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[22]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[21] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[21]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[20] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[20]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[19] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[19]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[18] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[18]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[17] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[17]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[16] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[16]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[15] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[15]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[14] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[14]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[13] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[13]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[12] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[12]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[11] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[11]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[10] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[10]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[9] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[9]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[8] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[8]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[7] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[7]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[6] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[6]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[5] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[5]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[4] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[4]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[3] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[3]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[2] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[2]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[1] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[1]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tdata_wr3_REG[0] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tdata_wr3[0]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tstrb_wr4_REG[7] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tstrb_wr4[7]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tstrb_wr4_REG[6] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tstrb_wr4[6]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tstrb_wr4_REG[5] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tstrb_wr4[5]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tstrb_wr4_REG[4] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tstrb_wr4[4]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tstrb_wr4_REG[3] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tstrb_wr4[3]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tstrb_wr4_REG[2] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tstrb_wr4[2]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tstrb_wr4_REG[1] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tstrb_wr4[1]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tstrb_wr4_REG[0] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tstrb_wr4[0]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tuser_wr5_REG[7] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tuser_wr5[7]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tuser_wr5_REG[6] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tuser_wr5[6]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tuser_wr5_REG[5] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tuser_wr5[5]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tuser_wr5_REG[4] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tuser_wr5[4]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tuser_wr5_REG[3] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tuser_wr5[3]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tuser_wr5_REG[2] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tuser_wr5[2]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tuser_wr5_REG[1] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tuser_wr5[1]));
Q_FDP4EP \_zzM2L253_mdxP5_kme_ib_tuser_wr5_REG[0] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5320), .R(n1750), .D(n1750), .Q(_zzM2L253_mdxP5_kme_ib_tuser_wr5[0]));
Q_INV U8402 ( .A(_zyixc_port_0_0_ack), .Z(n20));
Q_FDP4EP _zyixc_port_0_0_ack_REG  ( .CK(_zyM2L253_pbcMevClk12), .CE(n5336), .R(n1750), .D(n20), .Q(_zyixc_port_0_0_ack));
Q_INV U8404 ( .A(n5299), .Z(n19));
Q_FDP4EP _zyGfifoF0_L253_s4_req_6_REG  ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4850), .Q(_zyGfifoF0_L253_s4_req_6));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[559] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4849), .Q(_zyGfifoF0_L253_s4_data_6[559]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[558] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4848), .Q(_zyGfifoF0_L253_s4_data_6[558]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[557] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4847), .Q(_zyGfifoF0_L253_s4_data_6[557]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[556] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4846), .Q(_zyGfifoF0_L253_s4_data_6[556]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[555] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4845), .Q(_zyGfifoF0_L253_s4_data_6[555]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[554] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4844), .Q(_zyGfifoF0_L253_s4_data_6[554]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[553] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4843), .Q(_zyGfifoF0_L253_s4_data_6[553]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[552] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4842), .Q(_zyGfifoF0_L253_s4_data_6[552]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[551] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4841), .Q(_zyGfifoF0_L253_s4_data_6[551]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[550] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4840), .Q(_zyGfifoF0_L253_s4_data_6[550]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[549] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4839), .Q(_zyGfifoF0_L253_s4_data_6[549]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[548] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4838), .Q(_zyGfifoF0_L253_s4_data_6[548]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[547] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4837), .Q(_zyGfifoF0_L253_s4_data_6[547]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[546] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4836), .Q(_zyGfifoF0_L253_s4_data_6[546]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[545] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4835), .Q(_zyGfifoF0_L253_s4_data_6[545]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[544] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4834), .Q(_zyGfifoF0_L253_s4_data_6[544]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[543] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4833), .Q(_zyGfifoF0_L253_s4_data_6[543]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[542] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4832), .Q(_zyGfifoF0_L253_s4_data_6[542]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[541] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4831), .Q(_zyGfifoF0_L253_s4_data_6[541]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[540] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4830), .Q(_zyGfifoF0_L253_s4_data_6[540]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[539] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4829), .Q(_zyGfifoF0_L253_s4_data_6[539]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[538] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4828), .Q(_zyGfifoF0_L253_s4_data_6[538]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[537] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4827), .Q(_zyGfifoF0_L253_s4_data_6[537]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[536] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4826), .Q(_zyGfifoF0_L253_s4_data_6[536]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[535] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4825), .Q(_zyGfifoF0_L253_s4_data_6[535]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[534] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4824), .Q(_zyGfifoF0_L253_s4_data_6[534]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[533] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4823), .Q(_zyGfifoF0_L253_s4_data_6[533]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[532] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4822), .Q(_zyGfifoF0_L253_s4_data_6[532]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[531] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4821), .Q(_zyGfifoF0_L253_s4_data_6[531]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[530] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4820), .Q(_zyGfifoF0_L253_s4_data_6[530]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[529] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4819), .Q(_zyGfifoF0_L253_s4_data_6[529]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[528] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4818), .Q(_zyGfifoF0_L253_s4_data_6[528]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[527] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4817), .Q(_zyGfifoF0_L253_s4_data_6[527]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[526] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4816), .Q(_zyGfifoF0_L253_s4_data_6[526]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[525] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4815), .Q(_zyGfifoF0_L253_s4_data_6[525]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[524] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4814), .Q(_zyGfifoF0_L253_s4_data_6[524]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[523] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4813), .Q(_zyGfifoF0_L253_s4_data_6[523]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[522] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4812), .Q(_zyGfifoF0_L253_s4_data_6[522]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[521] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4811), .Q(_zyGfifoF0_L253_s4_data_6[521]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[520] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4810), .Q(_zyGfifoF0_L253_s4_data_6[520]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[519] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4809), .Q(_zyGfifoF0_L253_s4_data_6[519]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[518] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4808), .Q(_zyGfifoF0_L253_s4_data_6[518]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[517] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4807), .Q(_zyGfifoF0_L253_s4_data_6[517]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[516] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4806), .Q(_zyGfifoF0_L253_s4_data_6[516]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[515] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4805), .Q(_zyGfifoF0_L253_s4_data_6[515]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[514] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4804), .Q(_zyGfifoF0_L253_s4_data_6[514]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[513] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4803), .Q(_zyGfifoF0_L253_s4_data_6[513]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[512] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4802), .Q(_zyGfifoF0_L253_s4_data_6[512]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[511] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4801), .Q(_zyGfifoF0_L253_s4_data_6[511]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[510] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4800), .Q(_zyGfifoF0_L253_s4_data_6[510]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[509] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4799), .Q(_zyGfifoF0_L253_s4_data_6[509]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[508] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4798), .Q(_zyGfifoF0_L253_s4_data_6[508]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[507] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4797), .Q(_zyGfifoF0_L253_s4_data_6[507]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[506] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4796), .Q(_zyGfifoF0_L253_s4_data_6[506]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[505] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4795), .Q(_zyGfifoF0_L253_s4_data_6[505]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[504] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4794), .Q(_zyGfifoF0_L253_s4_data_6[504]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[503] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4793), .Q(_zyGfifoF0_L253_s4_data_6[503]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[502] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4792), .Q(_zyGfifoF0_L253_s4_data_6[502]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[501] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4791), .Q(_zyGfifoF0_L253_s4_data_6[501]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[500] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4790), .Q(_zyGfifoF0_L253_s4_data_6[500]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[499] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4789), .Q(_zyGfifoF0_L253_s4_data_6[499]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[498] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4788), .Q(_zyGfifoF0_L253_s4_data_6[498]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[497] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4787), .Q(_zyGfifoF0_L253_s4_data_6[497]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[496] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4786), .Q(_zyGfifoF0_L253_s4_data_6[496]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[495] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4785), .Q(_zyGfifoF0_L253_s4_data_6[495]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[494] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4784), .Q(_zyGfifoF0_L253_s4_data_6[494]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[493] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4783), .Q(_zyGfifoF0_L253_s4_data_6[493]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[492] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4782), .Q(_zyGfifoF0_L253_s4_data_6[492]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[491] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4781), .Q(_zyGfifoF0_L253_s4_data_6[491]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[490] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4780), .Q(_zyGfifoF0_L253_s4_data_6[490]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[489] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4779), .Q(_zyGfifoF0_L253_s4_data_6[489]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[488] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4778), .Q(_zyGfifoF0_L253_s4_data_6[488]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[487] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4777), .Q(_zyGfifoF0_L253_s4_data_6[487]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[486] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4776), .Q(_zyGfifoF0_L253_s4_data_6[486]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[485] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4775), .Q(_zyGfifoF0_L253_s4_data_6[485]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[484] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4774), .Q(_zyGfifoF0_L253_s4_data_6[484]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[483] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4773), .Q(_zyGfifoF0_L253_s4_data_6[483]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[482] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4772), .Q(_zyGfifoF0_L253_s4_data_6[482]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[481] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4771), .Q(_zyGfifoF0_L253_s4_data_6[481]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[480] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4770), .Q(_zyGfifoF0_L253_s4_data_6[480]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[479] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4769), .Q(_zyGfifoF0_L253_s4_data_6[479]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[478] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4768), .Q(_zyGfifoF0_L253_s4_data_6[478]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[477] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4767), .Q(_zyGfifoF0_L253_s4_data_6[477]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[476] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4766), .Q(_zyGfifoF0_L253_s4_data_6[476]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[475] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4765), .Q(_zyGfifoF0_L253_s4_data_6[475]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[474] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4764), .Q(_zyGfifoF0_L253_s4_data_6[474]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[473] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4763), .Q(_zyGfifoF0_L253_s4_data_6[473]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[472] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4762), .Q(_zyGfifoF0_L253_s4_data_6[472]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[471] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4761), .Q(_zyGfifoF0_L253_s4_data_6[471]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[470] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4760), .Q(_zyGfifoF0_L253_s4_data_6[470]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[469] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4759), .Q(_zyGfifoF0_L253_s4_data_6[469]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[468] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4758), .Q(_zyGfifoF0_L253_s4_data_6[468]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[467] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4757), .Q(_zyGfifoF0_L253_s4_data_6[467]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[466] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4756), .Q(_zyGfifoF0_L253_s4_data_6[466]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[465] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4755), .Q(_zyGfifoF0_L253_s4_data_6[465]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[464] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4754), .Q(_zyGfifoF0_L253_s4_data_6[464]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[463] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4753), .Q(_zyGfifoF0_L253_s4_data_6[463]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[462] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4752), .Q(_zyGfifoF0_L253_s4_data_6[462]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[461] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4751), .Q(_zyGfifoF0_L253_s4_data_6[461]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[460] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4750), .Q(_zyGfifoF0_L253_s4_data_6[460]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[459] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4749), .Q(_zyGfifoF0_L253_s4_data_6[459]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[458] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4748), .Q(_zyGfifoF0_L253_s4_data_6[458]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[457] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4747), .Q(_zyGfifoF0_L253_s4_data_6[457]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[456] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4746), .Q(_zyGfifoF0_L253_s4_data_6[456]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[455] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4745), .Q(_zyGfifoF0_L253_s4_data_6[455]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[454] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4744), .Q(_zyGfifoF0_L253_s4_data_6[454]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[453] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4743), .Q(_zyGfifoF0_L253_s4_data_6[453]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[452] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4742), .Q(_zyGfifoF0_L253_s4_data_6[452]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[451] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4741), .Q(_zyGfifoF0_L253_s4_data_6[451]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[450] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4740), .Q(_zyGfifoF0_L253_s4_data_6[450]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[449] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4739), .Q(_zyGfifoF0_L253_s4_data_6[449]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[448] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4738), .Q(_zyGfifoF0_L253_s4_data_6[448]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[447] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4737), .Q(_zyGfifoF0_L253_s4_data_6[447]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[446] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4736), .Q(_zyGfifoF0_L253_s4_data_6[446]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[445] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4735), .Q(_zyGfifoF0_L253_s4_data_6[445]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[444] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4734), .Q(_zyGfifoF0_L253_s4_data_6[444]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[443] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4733), .Q(_zyGfifoF0_L253_s4_data_6[443]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[442] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4732), .Q(_zyGfifoF0_L253_s4_data_6[442]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[441] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4731), .Q(_zyGfifoF0_L253_s4_data_6[441]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[440] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4730), .Q(_zyGfifoF0_L253_s4_data_6[440]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[439] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4729), .Q(_zyGfifoF0_L253_s4_data_6[439]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[438] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4728), .Q(_zyGfifoF0_L253_s4_data_6[438]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[437] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4727), .Q(_zyGfifoF0_L253_s4_data_6[437]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[436] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4726), .Q(_zyGfifoF0_L253_s4_data_6[436]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[435] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4725), .Q(_zyGfifoF0_L253_s4_data_6[435]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[434] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4724), .Q(_zyGfifoF0_L253_s4_data_6[434]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[433] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4723), .Q(_zyGfifoF0_L253_s4_data_6[433]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[432] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4722), .Q(_zyGfifoF0_L253_s4_data_6[432]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[431] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4721), .Q(_zyGfifoF0_L253_s4_data_6[431]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[430] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4720), .Q(_zyGfifoF0_L253_s4_data_6[430]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[429] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4719), .Q(_zyGfifoF0_L253_s4_data_6[429]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[428] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4718), .Q(_zyGfifoF0_L253_s4_data_6[428]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[427] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4717), .Q(_zyGfifoF0_L253_s4_data_6[427]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[426] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4716), .Q(_zyGfifoF0_L253_s4_data_6[426]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[425] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4715), .Q(_zyGfifoF0_L253_s4_data_6[425]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[424] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4714), .Q(_zyGfifoF0_L253_s4_data_6[424]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[423] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4713), .Q(_zyGfifoF0_L253_s4_data_6[423]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[422] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4712), .Q(_zyGfifoF0_L253_s4_data_6[422]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[421] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4711), .Q(_zyGfifoF0_L253_s4_data_6[421]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[420] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4710), .Q(_zyGfifoF0_L253_s4_data_6[420]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[419] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4709), .Q(_zyGfifoF0_L253_s4_data_6[419]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[418] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4708), .Q(_zyGfifoF0_L253_s4_data_6[418]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[417] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4707), .Q(_zyGfifoF0_L253_s4_data_6[417]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[416] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4706), .Q(_zyGfifoF0_L253_s4_data_6[416]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[415] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4705), .Q(_zyGfifoF0_L253_s4_data_6[415]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[414] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4704), .Q(_zyGfifoF0_L253_s4_data_6[414]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[413] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4703), .Q(_zyGfifoF0_L253_s4_data_6[413]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[412] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4702), .Q(_zyGfifoF0_L253_s4_data_6[412]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[411] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4701), .Q(_zyGfifoF0_L253_s4_data_6[411]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[410] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4700), .Q(_zyGfifoF0_L253_s4_data_6[410]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[409] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4699), .Q(_zyGfifoF0_L253_s4_data_6[409]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[408] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4698), .Q(_zyGfifoF0_L253_s4_data_6[408]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[407] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4697), .Q(_zyGfifoF0_L253_s4_data_6[407]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[406] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4696), .Q(_zyGfifoF0_L253_s4_data_6[406]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[405] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4695), .Q(_zyGfifoF0_L253_s4_data_6[405]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[404] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4694), .Q(_zyGfifoF0_L253_s4_data_6[404]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[403] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4693), .Q(_zyGfifoF0_L253_s4_data_6[403]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[402] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4692), .Q(_zyGfifoF0_L253_s4_data_6[402]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[401] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4691), .Q(_zyGfifoF0_L253_s4_data_6[401]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[400] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4690), .Q(_zyGfifoF0_L253_s4_data_6[400]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[399] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4689), .Q(_zyGfifoF0_L253_s4_data_6[399]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[398] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4688), .Q(_zyGfifoF0_L253_s4_data_6[398]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[397] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4687), .Q(_zyGfifoF0_L253_s4_data_6[397]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[396] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4686), .Q(_zyGfifoF0_L253_s4_data_6[396]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[395] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4685), .Q(_zyGfifoF0_L253_s4_data_6[395]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[394] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4684), .Q(_zyGfifoF0_L253_s4_data_6[394]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[393] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4683), .Q(_zyGfifoF0_L253_s4_data_6[393]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[392] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4682), .Q(_zyGfifoF0_L253_s4_data_6[392]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[391] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4681), .Q(_zyGfifoF0_L253_s4_data_6[391]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[390] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4680), .Q(_zyGfifoF0_L253_s4_data_6[390]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[389] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4679), .Q(_zyGfifoF0_L253_s4_data_6[389]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[388] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4678), .Q(_zyGfifoF0_L253_s4_data_6[388]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[387] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4677), .Q(_zyGfifoF0_L253_s4_data_6[387]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[386] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4676), .Q(_zyGfifoF0_L253_s4_data_6[386]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[385] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4675), .Q(_zyGfifoF0_L253_s4_data_6[385]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[384] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4674), .Q(_zyGfifoF0_L253_s4_data_6[384]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[383] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4673), .Q(_zyGfifoF0_L253_s4_data_6[383]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[382] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4672), .Q(_zyGfifoF0_L253_s4_data_6[382]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[381] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4671), .Q(_zyGfifoF0_L253_s4_data_6[381]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[380] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4670), .Q(_zyGfifoF0_L253_s4_data_6[380]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[379] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4669), .Q(_zyGfifoF0_L253_s4_data_6[379]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[378] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4668), .Q(_zyGfifoF0_L253_s4_data_6[378]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[377] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4667), .Q(_zyGfifoF0_L253_s4_data_6[377]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[376] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4666), .Q(_zyGfifoF0_L253_s4_data_6[376]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[375] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4665), .Q(_zyGfifoF0_L253_s4_data_6[375]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[374] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4664), .Q(_zyGfifoF0_L253_s4_data_6[374]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[373] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4663), .Q(_zyGfifoF0_L253_s4_data_6[373]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[372] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4662), .Q(_zyGfifoF0_L253_s4_data_6[372]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[371] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4661), .Q(_zyGfifoF0_L253_s4_data_6[371]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[370] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4660), .Q(_zyGfifoF0_L253_s4_data_6[370]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[369] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4659), .Q(_zyGfifoF0_L253_s4_data_6[369]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[368] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4658), .Q(_zyGfifoF0_L253_s4_data_6[368]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[367] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4657), .Q(_zyGfifoF0_L253_s4_data_6[367]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[366] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4656), .Q(_zyGfifoF0_L253_s4_data_6[366]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[365] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4655), .Q(_zyGfifoF0_L253_s4_data_6[365]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[364] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4654), .Q(_zyGfifoF0_L253_s4_data_6[364]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[363] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4653), .Q(_zyGfifoF0_L253_s4_data_6[363]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[362] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4652), .Q(_zyGfifoF0_L253_s4_data_6[362]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[361] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4651), .Q(_zyGfifoF0_L253_s4_data_6[361]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[360] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4650), .Q(_zyGfifoF0_L253_s4_data_6[360]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[359] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4649), .Q(_zyGfifoF0_L253_s4_data_6[359]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[358] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4648), .Q(_zyGfifoF0_L253_s4_data_6[358]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[357] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4647), .Q(_zyGfifoF0_L253_s4_data_6[357]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[356] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4646), .Q(_zyGfifoF0_L253_s4_data_6[356]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[355] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4645), .Q(_zyGfifoF0_L253_s4_data_6[355]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[354] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4644), .Q(_zyGfifoF0_L253_s4_data_6[354]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[353] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4643), .Q(_zyGfifoF0_L253_s4_data_6[353]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[352] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4642), .Q(_zyGfifoF0_L253_s4_data_6[352]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[351] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4641), .Q(_zyGfifoF0_L253_s4_data_6[351]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[350] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4640), .Q(_zyGfifoF0_L253_s4_data_6[350]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[349] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4639), .Q(_zyGfifoF0_L253_s4_data_6[349]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[348] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4638), .Q(_zyGfifoF0_L253_s4_data_6[348]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[347] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4637), .Q(_zyGfifoF0_L253_s4_data_6[347]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[346] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4636), .Q(_zyGfifoF0_L253_s4_data_6[346]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[345] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4635), .Q(_zyGfifoF0_L253_s4_data_6[345]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[344] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4634), .Q(_zyGfifoF0_L253_s4_data_6[344]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[343] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4633), .Q(_zyGfifoF0_L253_s4_data_6[343]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[342] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4632), .Q(_zyGfifoF0_L253_s4_data_6[342]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[341] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4631), .Q(_zyGfifoF0_L253_s4_data_6[341]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[340] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4630), .Q(_zyGfifoF0_L253_s4_data_6[340]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[339] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4629), .Q(_zyGfifoF0_L253_s4_data_6[339]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[338] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4628), .Q(_zyGfifoF0_L253_s4_data_6[338]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[337] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4627), .Q(_zyGfifoF0_L253_s4_data_6[337]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[336] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4626), .Q(_zyGfifoF0_L253_s4_data_6[336]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[335] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4625), .Q(_zyGfifoF0_L253_s4_data_6[335]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[334] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4624), .Q(_zyGfifoF0_L253_s4_data_6[334]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[333] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4623), .Q(_zyGfifoF0_L253_s4_data_6[333]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[332] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4622), .Q(_zyGfifoF0_L253_s4_data_6[332]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[331] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4621), .Q(_zyGfifoF0_L253_s4_data_6[331]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[330] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4620), .Q(_zyGfifoF0_L253_s4_data_6[330]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[329] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4619), .Q(_zyGfifoF0_L253_s4_data_6[329]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[328] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4618), .Q(_zyGfifoF0_L253_s4_data_6[328]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[327] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4617), .Q(_zyGfifoF0_L253_s4_data_6[327]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[326] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4616), .Q(_zyGfifoF0_L253_s4_data_6[326]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[325] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4615), .Q(_zyGfifoF0_L253_s4_data_6[325]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[324] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4614), .Q(_zyGfifoF0_L253_s4_data_6[324]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[323] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4613), .Q(_zyGfifoF0_L253_s4_data_6[323]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[322] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4612), .Q(_zyGfifoF0_L253_s4_data_6[322]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[321] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4611), .Q(_zyGfifoF0_L253_s4_data_6[321]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[320] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4610), .Q(_zyGfifoF0_L253_s4_data_6[320]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[319] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4609), .Q(_zyGfifoF0_L253_s4_data_6[319]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[318] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4608), .Q(_zyGfifoF0_L253_s4_data_6[318]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[317] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4607), .Q(_zyGfifoF0_L253_s4_data_6[317]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[316] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4606), .Q(_zyGfifoF0_L253_s4_data_6[316]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[315] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4605), .Q(_zyGfifoF0_L253_s4_data_6[315]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[314] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4604), .Q(_zyGfifoF0_L253_s4_data_6[314]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[313] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4603), .Q(_zyGfifoF0_L253_s4_data_6[313]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[312] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4602), .Q(_zyGfifoF0_L253_s4_data_6[312]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[311] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4601), .Q(_zyGfifoF0_L253_s4_data_6[311]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[310] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4600), .Q(_zyGfifoF0_L253_s4_data_6[310]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[309] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4599), .Q(_zyGfifoF0_L253_s4_data_6[309]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[308] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4598), .Q(_zyGfifoF0_L253_s4_data_6[308]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[307] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4597), .Q(_zyGfifoF0_L253_s4_data_6[307]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[306] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4596), .Q(_zyGfifoF0_L253_s4_data_6[306]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[305] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4595), .Q(_zyGfifoF0_L253_s4_data_6[305]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[304] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4594), .Q(_zyGfifoF0_L253_s4_data_6[304]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[303] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4593), .Q(_zyGfifoF0_L253_s4_data_6[303]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[302] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4592), .Q(_zyGfifoF0_L253_s4_data_6[302]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[301] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4591), .Q(_zyGfifoF0_L253_s4_data_6[301]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[300] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4590), .Q(_zyGfifoF0_L253_s4_data_6[300]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[299] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4589), .Q(_zyGfifoF0_L253_s4_data_6[299]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[298] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4588), .Q(_zyGfifoF0_L253_s4_data_6[298]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[297] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4587), .Q(_zyGfifoF0_L253_s4_data_6[297]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[296] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4586), .Q(_zyGfifoF0_L253_s4_data_6[296]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[295] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4585), .Q(_zyGfifoF0_L253_s4_data_6[295]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[294] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4584), .Q(_zyGfifoF0_L253_s4_data_6[294]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[293] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4583), .Q(_zyGfifoF0_L253_s4_data_6[293]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[292] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4582), .Q(_zyGfifoF0_L253_s4_data_6[292]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[291] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4581), .Q(_zyGfifoF0_L253_s4_data_6[291]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[290] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4580), .Q(_zyGfifoF0_L253_s4_data_6[290]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[289] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4579), .Q(_zyGfifoF0_L253_s4_data_6[289]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[288] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4578), .Q(_zyGfifoF0_L253_s4_data_6[288]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[287] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4577), .Q(_zyGfifoF0_L253_s4_data_6[287]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[286] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4576), .Q(_zyGfifoF0_L253_s4_data_6[286]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[285] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4575), .Q(_zyGfifoF0_L253_s4_data_6[285]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[284] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4574), .Q(_zyGfifoF0_L253_s4_data_6[284]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[283] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4573), .Q(_zyGfifoF0_L253_s4_data_6[283]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[282] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4572), .Q(_zyGfifoF0_L253_s4_data_6[282]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[281] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4571), .Q(_zyGfifoF0_L253_s4_data_6[281]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[280] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4570), .Q(_zyGfifoF0_L253_s4_data_6[280]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[279] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4569), .Q(_zyGfifoF0_L253_s4_data_6[279]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[278] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4568), .Q(_zyGfifoF0_L253_s4_data_6[278]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[277] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4567), .Q(_zyGfifoF0_L253_s4_data_6[277]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[276] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4566), .Q(_zyGfifoF0_L253_s4_data_6[276]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[275] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4565), .Q(_zyGfifoF0_L253_s4_data_6[275]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[274] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4564), .Q(_zyGfifoF0_L253_s4_data_6[274]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[273] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4563), .Q(_zyGfifoF0_L253_s4_data_6[273]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[272] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4562), .Q(_zyGfifoF0_L253_s4_data_6[272]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[271] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4561), .Q(_zyGfifoF0_L253_s4_data_6[271]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[270] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4560), .Q(_zyGfifoF0_L253_s4_data_6[270]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[269] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4559), .Q(_zyGfifoF0_L253_s4_data_6[269]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[268] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4558), .Q(_zyGfifoF0_L253_s4_data_6[268]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[267] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4557), .Q(_zyGfifoF0_L253_s4_data_6[267]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[266] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4556), .Q(_zyGfifoF0_L253_s4_data_6[266]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[265] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4555), .Q(_zyGfifoF0_L253_s4_data_6[265]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[264] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4554), .Q(_zyGfifoF0_L253_s4_data_6[264]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[263] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4553), .Q(_zyGfifoF0_L253_s4_data_6[263]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[262] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4552), .Q(_zyGfifoF0_L253_s4_data_6[262]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[261] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4551), .Q(_zyGfifoF0_L253_s4_data_6[261]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[260] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4550), .Q(_zyGfifoF0_L253_s4_data_6[260]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[259] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4549), .Q(_zyGfifoF0_L253_s4_data_6[259]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[258] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4548), .Q(_zyGfifoF0_L253_s4_data_6[258]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[257] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4547), .Q(_zyGfifoF0_L253_s4_data_6[257]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[256] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4546), .Q(_zyGfifoF0_L253_s4_data_6[256]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[255] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4545), .Q(_zyGfifoF0_L253_s4_data_6[255]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[254] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4544), .Q(_zyGfifoF0_L253_s4_data_6[254]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[253] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4543), .Q(_zyGfifoF0_L253_s4_data_6[253]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[252] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4542), .Q(_zyGfifoF0_L253_s4_data_6[252]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[251] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4541), .Q(_zyGfifoF0_L253_s4_data_6[251]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[250] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4540), .Q(_zyGfifoF0_L253_s4_data_6[250]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[249] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4539), .Q(_zyGfifoF0_L253_s4_data_6[249]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[248] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4538), .Q(_zyGfifoF0_L253_s4_data_6[248]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[247] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4537), .Q(_zyGfifoF0_L253_s4_data_6[247]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[246] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4536), .Q(_zyGfifoF0_L253_s4_data_6[246]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[245] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4535), .Q(_zyGfifoF0_L253_s4_data_6[245]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[244] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4534), .Q(_zyGfifoF0_L253_s4_data_6[244]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[243] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4533), .Q(_zyGfifoF0_L253_s4_data_6[243]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[242] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4532), .Q(_zyGfifoF0_L253_s4_data_6[242]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[241] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4531), .Q(_zyGfifoF0_L253_s4_data_6[241]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[240] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4530), .Q(_zyGfifoF0_L253_s4_data_6[240]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[239] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4529), .Q(_zyGfifoF0_L253_s4_data_6[239]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[238] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4528), .Q(_zyGfifoF0_L253_s4_data_6[238]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[237] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4527), .Q(_zyGfifoF0_L253_s4_data_6[237]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[236] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4526), .Q(_zyGfifoF0_L253_s4_data_6[236]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[235] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4525), .Q(_zyGfifoF0_L253_s4_data_6[235]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[234] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4524), .Q(_zyGfifoF0_L253_s4_data_6[234]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[233] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4523), .Q(_zyGfifoF0_L253_s4_data_6[233]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[232] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4522), .Q(_zyGfifoF0_L253_s4_data_6[232]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[231] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4521), .Q(_zyGfifoF0_L253_s4_data_6[231]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[230] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4520), .Q(_zyGfifoF0_L253_s4_data_6[230]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[229] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4519), .Q(_zyGfifoF0_L253_s4_data_6[229]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[228] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4518), .Q(_zyGfifoF0_L253_s4_data_6[228]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[227] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4517), .Q(_zyGfifoF0_L253_s4_data_6[227]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[226] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4516), .Q(_zyGfifoF0_L253_s4_data_6[226]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[225] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4515), .Q(_zyGfifoF0_L253_s4_data_6[225]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[224] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4514), .Q(_zyGfifoF0_L253_s4_data_6[224]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[223] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4513), .Q(_zyGfifoF0_L253_s4_data_6[223]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[222] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4512), .Q(_zyGfifoF0_L253_s4_data_6[222]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[221] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4511), .Q(_zyGfifoF0_L253_s4_data_6[221]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[220] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4510), .Q(_zyGfifoF0_L253_s4_data_6[220]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[219] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4509), .Q(_zyGfifoF0_L253_s4_data_6[219]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[218] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4508), .Q(_zyGfifoF0_L253_s4_data_6[218]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[217] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4507), .Q(_zyGfifoF0_L253_s4_data_6[217]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[216] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4506), .Q(_zyGfifoF0_L253_s4_data_6[216]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[215] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4505), .Q(_zyGfifoF0_L253_s4_data_6[215]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[214] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4504), .Q(_zyGfifoF0_L253_s4_data_6[214]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[213] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4503), .Q(_zyGfifoF0_L253_s4_data_6[213]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[212] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4502), .Q(_zyGfifoF0_L253_s4_data_6[212]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[211] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4501), .Q(_zyGfifoF0_L253_s4_data_6[211]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[210] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4500), .Q(_zyGfifoF0_L253_s4_data_6[210]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[209] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4499), .Q(_zyGfifoF0_L253_s4_data_6[209]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[208] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4498), .Q(_zyGfifoF0_L253_s4_data_6[208]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[207] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4497), .Q(_zyGfifoF0_L253_s4_data_6[207]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[206] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4496), .Q(_zyGfifoF0_L253_s4_data_6[206]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[205] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4495), .Q(_zyGfifoF0_L253_s4_data_6[205]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[204] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4494), .Q(_zyGfifoF0_L253_s4_data_6[204]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[203] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4493), .Q(_zyGfifoF0_L253_s4_data_6[203]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[202] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4492), .Q(_zyGfifoF0_L253_s4_data_6[202]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[201] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4491), .Q(_zyGfifoF0_L253_s4_data_6[201]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[200] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4490), .Q(_zyGfifoF0_L253_s4_data_6[200]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[199] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4489), .Q(_zyGfifoF0_L253_s4_data_6[199]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[198] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4488), .Q(_zyGfifoF0_L253_s4_data_6[198]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[197] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4487), .Q(_zyGfifoF0_L253_s4_data_6[197]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[196] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4486), .Q(_zyGfifoF0_L253_s4_data_6[196]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[195] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4485), .Q(_zyGfifoF0_L253_s4_data_6[195]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[194] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4484), .Q(_zyGfifoF0_L253_s4_data_6[194]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[193] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4483), .Q(_zyGfifoF0_L253_s4_data_6[193]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[192] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4482), .Q(_zyGfifoF0_L253_s4_data_6[192]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[191] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4481), .Q(_zyGfifoF0_L253_s4_data_6[191]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[190] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4480), .Q(_zyGfifoF0_L253_s4_data_6[190]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[189] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4479), .Q(_zyGfifoF0_L253_s4_data_6[189]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[188] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4478), .Q(_zyGfifoF0_L253_s4_data_6[188]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[187] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4477), .Q(_zyGfifoF0_L253_s4_data_6[187]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[186] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4476), .Q(_zyGfifoF0_L253_s4_data_6[186]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[185] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4475), .Q(_zyGfifoF0_L253_s4_data_6[185]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[184] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4474), .Q(_zyGfifoF0_L253_s4_data_6[184]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[183] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4473), .Q(_zyGfifoF0_L253_s4_data_6[183]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[182] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4472), .Q(_zyGfifoF0_L253_s4_data_6[182]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[181] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4471), .Q(_zyGfifoF0_L253_s4_data_6[181]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[180] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4470), .Q(_zyGfifoF0_L253_s4_data_6[180]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[179] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4469), .Q(_zyGfifoF0_L253_s4_data_6[179]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[178] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4468), .Q(_zyGfifoF0_L253_s4_data_6[178]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[177] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4467), .Q(_zyGfifoF0_L253_s4_data_6[177]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[176] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4466), .Q(_zyGfifoF0_L253_s4_data_6[176]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[175] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4465), .Q(_zyGfifoF0_L253_s4_data_6[175]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[174] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4464), .Q(_zyGfifoF0_L253_s4_data_6[174]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[173] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4463), .Q(_zyGfifoF0_L253_s4_data_6[173]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[172] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4462), .Q(_zyGfifoF0_L253_s4_data_6[172]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[171] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4461), .Q(_zyGfifoF0_L253_s4_data_6[171]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[170] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4460), .Q(_zyGfifoF0_L253_s4_data_6[170]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[169] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4459), .Q(_zyGfifoF0_L253_s4_data_6[169]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[168] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4458), .Q(_zyGfifoF0_L253_s4_data_6[168]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[167] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4457), .Q(_zyGfifoF0_L253_s4_data_6[167]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[166] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4456), .Q(_zyGfifoF0_L253_s4_data_6[166]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[165] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4455), .Q(_zyGfifoF0_L253_s4_data_6[165]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[164] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4454), .Q(_zyGfifoF0_L253_s4_data_6[164]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[163] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4453), .Q(_zyGfifoF0_L253_s4_data_6[163]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[162] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4452), .Q(_zyGfifoF0_L253_s4_data_6[162]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[161] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4451), .Q(_zyGfifoF0_L253_s4_data_6[161]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[160] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4450), .Q(_zyGfifoF0_L253_s4_data_6[160]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[159] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4449), .Q(_zyGfifoF0_L253_s4_data_6[159]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[158] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4448), .Q(_zyGfifoF0_L253_s4_data_6[158]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[157] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4447), .Q(_zyGfifoF0_L253_s4_data_6[157]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[156] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4446), .Q(_zyGfifoF0_L253_s4_data_6[156]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[155] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4445), .Q(_zyGfifoF0_L253_s4_data_6[155]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[154] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4444), .Q(_zyGfifoF0_L253_s4_data_6[154]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[153] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4443), .Q(_zyGfifoF0_L253_s4_data_6[153]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[152] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4442), .Q(_zyGfifoF0_L253_s4_data_6[152]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[151] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4441), .Q(_zyGfifoF0_L253_s4_data_6[151]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[150] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4440), .Q(_zyGfifoF0_L253_s4_data_6[150]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[149] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4439), .Q(_zyGfifoF0_L253_s4_data_6[149]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[148] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4438), .Q(_zyGfifoF0_L253_s4_data_6[148]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[147] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4437), .Q(_zyGfifoF0_L253_s4_data_6[147]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[146] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4436), .Q(_zyGfifoF0_L253_s4_data_6[146]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[145] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4435), .Q(_zyGfifoF0_L253_s4_data_6[145]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[144] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4434), .Q(_zyGfifoF0_L253_s4_data_6[144]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[143] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4433), .Q(_zyGfifoF0_L253_s4_data_6[143]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[142] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4432), .Q(_zyGfifoF0_L253_s4_data_6[142]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[141] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4431), .Q(_zyGfifoF0_L253_s4_data_6[141]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[140] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4430), .Q(_zyGfifoF0_L253_s4_data_6[140]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[139] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4429), .Q(_zyGfifoF0_L253_s4_data_6[139]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[138] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4428), .Q(_zyGfifoF0_L253_s4_data_6[138]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[137] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4427), .Q(_zyGfifoF0_L253_s4_data_6[137]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[136] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4426), .Q(_zyGfifoF0_L253_s4_data_6[136]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[135] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4425), .Q(_zyGfifoF0_L253_s4_data_6[135]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[134] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4424), .Q(_zyGfifoF0_L253_s4_data_6[134]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[133] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4423), .Q(_zyGfifoF0_L253_s4_data_6[133]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[132] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4422), .Q(_zyGfifoF0_L253_s4_data_6[132]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[131] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4421), .Q(_zyGfifoF0_L253_s4_data_6[131]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[130] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4420), .Q(_zyGfifoF0_L253_s4_data_6[130]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[129] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4419), .Q(_zyGfifoF0_L253_s4_data_6[129]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[128] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4418), .Q(_zyGfifoF0_L253_s4_data_6[128]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[127] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4417), .Q(_zyGfifoF0_L253_s4_data_6[127]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[126] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4416), .Q(_zyGfifoF0_L253_s4_data_6[126]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[125] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4415), .Q(_zyGfifoF0_L253_s4_data_6[125]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[124] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4414), .Q(_zyGfifoF0_L253_s4_data_6[124]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[123] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4413), .Q(_zyGfifoF0_L253_s4_data_6[123]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[122] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4412), .Q(_zyGfifoF0_L253_s4_data_6[122]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[121] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4411), .Q(_zyGfifoF0_L253_s4_data_6[121]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[120] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4410), .Q(_zyGfifoF0_L253_s4_data_6[120]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[119] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4409), .Q(_zyGfifoF0_L253_s4_data_6[119]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[118] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4408), .Q(_zyGfifoF0_L253_s4_data_6[118]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[117] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4407), .Q(_zyGfifoF0_L253_s4_data_6[117]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[116] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4406), .Q(_zyGfifoF0_L253_s4_data_6[116]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[115] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4405), .Q(_zyGfifoF0_L253_s4_data_6[115]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[114] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4404), .Q(_zyGfifoF0_L253_s4_data_6[114]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[113] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4403), .Q(_zyGfifoF0_L253_s4_data_6[113]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[112] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4402), .Q(_zyGfifoF0_L253_s4_data_6[112]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[111] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4401), .Q(_zyGfifoF0_L253_s4_data_6[111]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[110] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4400), .Q(_zyGfifoF0_L253_s4_data_6[110]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[109] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4399), .Q(_zyGfifoF0_L253_s4_data_6[109]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[108] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4398), .Q(_zyGfifoF0_L253_s4_data_6[108]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[107] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4397), .Q(_zyGfifoF0_L253_s4_data_6[107]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[106] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4396), .Q(_zyGfifoF0_L253_s4_data_6[106]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[105] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4395), .Q(_zyGfifoF0_L253_s4_data_6[105]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[104] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4394), .Q(_zyGfifoF0_L253_s4_data_6[104]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[103] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4393), .Q(_zyGfifoF0_L253_s4_data_6[103]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[102] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4392), .Q(_zyGfifoF0_L253_s4_data_6[102]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[101] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4391), .Q(_zyGfifoF0_L253_s4_data_6[101]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[100] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4390), .Q(_zyGfifoF0_L253_s4_data_6[100]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[99] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4389), .Q(_zyGfifoF0_L253_s4_data_6[99]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[98] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4388), .Q(_zyGfifoF0_L253_s4_data_6[98]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[97] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4387), .Q(_zyGfifoF0_L253_s4_data_6[97]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[96] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4386), .Q(_zyGfifoF0_L253_s4_data_6[96]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[95] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4385), .Q(_zyGfifoF0_L253_s4_data_6[95]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[94] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4384), .Q(_zyGfifoF0_L253_s4_data_6[94]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[93] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4383), .Q(_zyGfifoF0_L253_s4_data_6[93]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[92] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4382), .Q(_zyGfifoF0_L253_s4_data_6[92]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[91] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4381), .Q(_zyGfifoF0_L253_s4_data_6[91]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[90] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4380), .Q(_zyGfifoF0_L253_s4_data_6[90]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[89] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4379), .Q(_zyGfifoF0_L253_s4_data_6[89]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[88] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4378), .Q(_zyGfifoF0_L253_s4_data_6[88]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[87] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4377), .Q(_zyGfifoF0_L253_s4_data_6[87]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[86] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4376), .Q(_zyGfifoF0_L253_s4_data_6[86]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[85] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4375), .Q(_zyGfifoF0_L253_s4_data_6[85]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[84] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4374), .Q(_zyGfifoF0_L253_s4_data_6[84]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[83] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4373), .Q(_zyGfifoF0_L253_s4_data_6[83]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[82] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4372), .Q(_zyGfifoF0_L253_s4_data_6[82]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[81] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4371), .Q(_zyGfifoF0_L253_s4_data_6[81]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[80] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4370), .Q(_zyGfifoF0_L253_s4_data_6[80]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[79] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4369), .Q(_zyGfifoF0_L253_s4_data_6[79]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[78] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4368), .Q(_zyGfifoF0_L253_s4_data_6[78]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[77] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4367), .Q(_zyGfifoF0_L253_s4_data_6[77]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[76] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4366), .Q(_zyGfifoF0_L253_s4_data_6[76]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[75] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4365), .Q(_zyGfifoF0_L253_s4_data_6[75]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[74] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4364), .Q(_zyGfifoF0_L253_s4_data_6[74]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[73] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4363), .Q(_zyGfifoF0_L253_s4_data_6[73]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[72] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4362), .Q(_zyGfifoF0_L253_s4_data_6[72]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[71] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4361), .Q(_zyGfifoF0_L253_s4_data_6[71]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[70] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4360), .Q(_zyGfifoF0_L253_s4_data_6[70]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[69] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4359), .Q(_zyGfifoF0_L253_s4_data_6[69]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[68] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4358), .Q(_zyGfifoF0_L253_s4_data_6[68]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[67] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4357), .Q(_zyGfifoF0_L253_s4_data_6[67]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[66] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4356), .Q(_zyGfifoF0_L253_s4_data_6[66]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[65] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4355), .Q(_zyGfifoF0_L253_s4_data_6[65]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[64] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4354), .Q(_zyGfifoF0_L253_s4_data_6[64]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[63] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4353), .Q(_zyGfifoF0_L253_s4_data_6[63]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[62] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4352), .Q(_zyGfifoF0_L253_s4_data_6[62]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[61] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4351), .Q(_zyGfifoF0_L253_s4_data_6[61]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[60] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4350), .Q(_zyGfifoF0_L253_s4_data_6[60]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[59] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4349), .Q(_zyGfifoF0_L253_s4_data_6[59]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[58] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4348), .Q(_zyGfifoF0_L253_s4_data_6[58]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[57] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4347), .Q(_zyGfifoF0_L253_s4_data_6[57]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[56] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4346), .Q(_zyGfifoF0_L253_s4_data_6[56]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[55] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4345), .Q(_zyGfifoF0_L253_s4_data_6[55]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[54] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4344), .Q(_zyGfifoF0_L253_s4_data_6[54]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[53] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4343), .Q(_zyGfifoF0_L253_s4_data_6[53]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[52] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4342), .Q(_zyGfifoF0_L253_s4_data_6[52]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[51] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4341), .Q(_zyGfifoF0_L253_s4_data_6[51]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[50] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4340), .Q(_zyGfifoF0_L253_s4_data_6[50]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[49] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4339), .Q(_zyGfifoF0_L253_s4_data_6[49]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[48] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4338), .Q(_zyGfifoF0_L253_s4_data_6[48]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[47] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4337), .Q(_zyGfifoF0_L253_s4_data_6[47]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[46] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4336), .Q(_zyGfifoF0_L253_s4_data_6[46]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[45] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4335), .Q(_zyGfifoF0_L253_s4_data_6[45]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[44] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4334), .Q(_zyGfifoF0_L253_s4_data_6[44]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[43] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4333), .Q(_zyGfifoF0_L253_s4_data_6[43]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[42] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4332), .Q(_zyGfifoF0_L253_s4_data_6[42]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[41] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4331), .Q(_zyGfifoF0_L253_s4_data_6[41]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[40] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4330), .Q(_zyGfifoF0_L253_s4_data_6[40]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[39] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4329), .Q(_zyGfifoF0_L253_s4_data_6[39]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[38] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4328), .Q(_zyGfifoF0_L253_s4_data_6[38]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[37] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4327), .Q(_zyGfifoF0_L253_s4_data_6[37]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[36] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4326), .Q(_zyGfifoF0_L253_s4_data_6[36]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[35] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4325), .Q(_zyGfifoF0_L253_s4_data_6[35]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[34] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4324), .Q(_zyGfifoF0_L253_s4_data_6[34]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[33] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4323), .Q(_zyGfifoF0_L253_s4_data_6[33]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[32] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4322), .Q(_zyGfifoF0_L253_s4_data_6[32]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[31] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4321), .Q(_zyGfifoF0_L253_s4_data_6[31]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[30] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4320), .Q(_zyGfifoF0_L253_s4_data_6[30]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[29] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4319), .Q(_zyGfifoF0_L253_s4_data_6[29]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[28] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4318), .Q(_zyGfifoF0_L253_s4_data_6[28]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[27] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4317), .Q(_zyGfifoF0_L253_s4_data_6[27]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[26] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4316), .Q(_zyGfifoF0_L253_s4_data_6[26]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[25] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4315), .Q(_zyGfifoF0_L253_s4_data_6[25]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[24] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4314), .Q(_zyGfifoF0_L253_s4_data_6[24]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[23] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4313), .Q(_zyGfifoF0_L253_s4_data_6[23]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[22] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4312), .Q(_zyGfifoF0_L253_s4_data_6[22]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[21] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4311), .Q(_zyGfifoF0_L253_s4_data_6[21]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[20] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4310), .Q(_zyGfifoF0_L253_s4_data_6[20]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[19] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4309), .Q(_zyGfifoF0_L253_s4_data_6[19]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[18] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4308), .Q(_zyGfifoF0_L253_s4_data_6[18]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[17] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4307), .Q(_zyGfifoF0_L253_s4_data_6[17]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[16] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4306), .Q(_zyGfifoF0_L253_s4_data_6[16]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[15] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4305), .Q(_zyGfifoF0_L253_s4_data_6[15]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[14] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4304), .Q(_zyGfifoF0_L253_s4_data_6[14]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[13] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4303), .Q(_zyGfifoF0_L253_s4_data_6[13]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[12] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4302), .Q(_zyGfifoF0_L253_s4_data_6[12]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[11] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4301), .Q(_zyGfifoF0_L253_s4_data_6[11]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[10] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4300), .Q(_zyGfifoF0_L253_s4_data_6[10]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[9] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4299), .Q(_zyGfifoF0_L253_s4_data_6[9]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[8] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4298), .Q(_zyGfifoF0_L253_s4_data_6[8]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[7] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4297), .Q(_zyGfifoF0_L253_s4_data_6[7]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[6] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4296), .Q(_zyGfifoF0_L253_s4_data_6[6]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[5] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4295), .Q(_zyGfifoF0_L253_s4_data_6[5]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[4] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4294), .Q(_zyGfifoF0_L253_s4_data_6[4]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[3] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4293), .Q(_zyGfifoF0_L253_s4_data_6[3]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[2] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4292), .Q(_zyGfifoF0_L253_s4_data_6[2]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[1] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4291), .Q(_zyGfifoF0_L253_s4_data_6[1]));
Q_FDP4EP \_zyGfifoF0_L253_s4_data_6_REG[0] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4290), .Q(_zyGfifoF0_L253_s4_data_6[0]));
Q_FDP4EP \_zyGfifoF0_L253_s4_cbid_6_REG[19] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4289), .Q(_zyGfifoF0_L253_s4_cbid_6[19]));
Q_FDP4EP \_zyGfifoF0_L253_s4_cbid_6_REG[18] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4288), .Q(_zyGfifoF0_L253_s4_cbid_6[18]));
Q_FDP4EP \_zyGfifoF0_L253_s4_cbid_6_REG[17] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4287), .Q(_zyGfifoF0_L253_s4_cbid_6[17]));
Q_FDP4EP \_zyGfifoF0_L253_s4_cbid_6_REG[16] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4286), .Q(_zyGfifoF0_L253_s4_cbid_6[16]));
Q_FDP4EP \_zyGfifoF0_L253_s4_cbid_6_REG[15] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4285), .Q(_zyGfifoF0_L253_s4_cbid_6[15]));
Q_FDP4EP \_zyGfifoF0_L253_s4_cbid_6_REG[14] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4284), .Q(_zyGfifoF0_L253_s4_cbid_6[14]));
Q_FDP4EP \_zyGfifoF0_L253_s4_cbid_6_REG[13] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4283), .Q(_zyGfifoF0_L253_s4_cbid_6[13]));
Q_FDP4EP \_zyGfifoF0_L253_s4_cbid_6_REG[12] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4282), .Q(_zyGfifoF0_L253_s4_cbid_6[12]));
Q_FDP4EP \_zyGfifoF0_L253_s4_cbid_6_REG[11] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4281), .Q(_zyGfifoF0_L253_s4_cbid_6[11]));
Q_FDP4EP \_zyGfifoF0_L253_s4_cbid_6_REG[10] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4280), .Q(_zyGfifoF0_L253_s4_cbid_6[10]));
Q_FDP4EP \_zyGfifoF0_L253_s4_cbid_6_REG[9] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4279), .Q(_zyGfifoF0_L253_s4_cbid_6[9]));
Q_FDP4EP \_zyGfifoF0_L253_s4_cbid_6_REG[8] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4278), .Q(_zyGfifoF0_L253_s4_cbid_6[8]));
Q_FDP4EP \_zyGfifoF0_L253_s4_cbid_6_REG[7] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4277), .Q(_zyGfifoF0_L253_s4_cbid_6[7]));
Q_FDP4EP \_zyGfifoF0_L253_s4_cbid_6_REG[6] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4276), .Q(_zyGfifoF0_L253_s4_cbid_6[6]));
Q_FDP4EP \_zyGfifoF0_L253_s4_cbid_6_REG[5] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4275), .Q(_zyGfifoF0_L253_s4_cbid_6[5]));
Q_FDP4EP \_zyGfifoF0_L253_s4_cbid_6_REG[4] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4274), .Q(_zyGfifoF0_L253_s4_cbid_6[4]));
Q_FDP4EP \_zyGfifoF0_L253_s4_cbid_6_REG[3] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4273), .Q(_zyGfifoF0_L253_s4_cbid_6[3]));
Q_FDP4EP \_zyGfifoF0_L253_s4_cbid_6_REG[2] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4272), .Q(_zyGfifoF0_L253_s4_cbid_6[2]));
Q_FDP4EP \_zyGfifoF0_L253_s4_cbid_6_REG[1] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4271), .Q(_zyGfifoF0_L253_s4_cbid_6[1]));
Q_FDP4EP \_zyGfifoF0_L253_s4_cbid_6_REG[0] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n4270), .Q(_zyGfifoF0_L253_s4_cbid_6[0]));
Q_INV U8986 ( .A(n5302), .Z(n18));
Q_FDP4EP _zyGfifoF1_L253_s2_req_7_REG  ( .CK(_zyM2L253_pbcMevClk12), .CE(n18), .R(n1750), .D(n4269), .Q(_zyGfifoF1_L253_s2_req_7));
Q_FDP4EP \_zyGfifoF1_L253_s2_cbid_7_REG[19] ( .CK(_zyM2L253_pbcMevClk12), .CE(n18), .R(n1750), .D(n4268), .Q(_zyGfifoF1_L253_s2_cbid_7[19]));
Q_FDP4EP \_zyGfifoF1_L253_s2_cbid_7_REG[18] ( .CK(_zyM2L253_pbcMevClk12), .CE(n18), .R(n1750), .D(n4267), .Q(_zyGfifoF1_L253_s2_cbid_7[18]));
Q_FDP4EP \_zyGfifoF1_L253_s2_cbid_7_REG[17] ( .CK(_zyM2L253_pbcMevClk12), .CE(n18), .R(n1750), .D(n4266), .Q(_zyGfifoF1_L253_s2_cbid_7[17]));
Q_FDP4EP \_zyGfifoF1_L253_s2_cbid_7_REG[16] ( .CK(_zyM2L253_pbcMevClk12), .CE(n18), .R(n1750), .D(n4265), .Q(_zyGfifoF1_L253_s2_cbid_7[16]));
Q_FDP4EP \_zyGfifoF1_L253_s2_cbid_7_REG[15] ( .CK(_zyM2L253_pbcMevClk12), .CE(n18), .R(n1750), .D(n4264), .Q(_zyGfifoF1_L253_s2_cbid_7[15]));
Q_FDP4EP \_zyGfifoF1_L253_s2_cbid_7_REG[14] ( .CK(_zyM2L253_pbcMevClk12), .CE(n18), .R(n1750), .D(n4263), .Q(_zyGfifoF1_L253_s2_cbid_7[14]));
Q_FDP4EP \_zyGfifoF1_L253_s2_cbid_7_REG[13] ( .CK(_zyM2L253_pbcMevClk12), .CE(n18), .R(n1750), .D(n4262), .Q(_zyGfifoF1_L253_s2_cbid_7[13]));
Q_FDP4EP \_zyGfifoF1_L253_s2_cbid_7_REG[12] ( .CK(_zyM2L253_pbcMevClk12), .CE(n18), .R(n1750), .D(n4261), .Q(_zyGfifoF1_L253_s2_cbid_7[12]));
Q_FDP4EP \_zyGfifoF1_L253_s2_cbid_7_REG[11] ( .CK(_zyM2L253_pbcMevClk12), .CE(n18), .R(n1750), .D(n4260), .Q(_zyGfifoF1_L253_s2_cbid_7[11]));
Q_FDP4EP \_zyGfifoF1_L253_s2_cbid_7_REG[10] ( .CK(_zyM2L253_pbcMevClk12), .CE(n18), .R(n1750), .D(n4259), .Q(_zyGfifoF1_L253_s2_cbid_7[10]));
Q_FDP4EP \_zyGfifoF1_L253_s2_cbid_7_REG[9] ( .CK(_zyM2L253_pbcMevClk12), .CE(n18), .R(n1750), .D(n4258), .Q(_zyGfifoF1_L253_s2_cbid_7[9]));
Q_FDP4EP \_zyGfifoF1_L253_s2_cbid_7_REG[8] ( .CK(_zyM2L253_pbcMevClk12), .CE(n18), .R(n1750), .D(n4257), .Q(_zyGfifoF1_L253_s2_cbid_7[8]));
Q_FDP4EP \_zyGfifoF1_L253_s2_cbid_7_REG[7] ( .CK(_zyM2L253_pbcMevClk12), .CE(n18), .R(n1750), .D(n4256), .Q(_zyGfifoF1_L253_s2_cbid_7[7]));
Q_FDP4EP \_zyGfifoF1_L253_s2_cbid_7_REG[6] ( .CK(_zyM2L253_pbcMevClk12), .CE(n18), .R(n1750), .D(n4255), .Q(_zyGfifoF1_L253_s2_cbid_7[6]));
Q_FDP4EP \_zyGfifoF1_L253_s2_cbid_7_REG[5] ( .CK(_zyM2L253_pbcMevClk12), .CE(n18), .R(n1750), .D(n4254), .Q(_zyGfifoF1_L253_s2_cbid_7[5]));
Q_FDP4EP \_zyGfifoF1_L253_s2_cbid_7_REG[4] ( .CK(_zyM2L253_pbcMevClk12), .CE(n18), .R(n1750), .D(n4253), .Q(_zyGfifoF1_L253_s2_cbid_7[4]));
Q_FDP4EP \_zyGfifoF1_L253_s2_cbid_7_REG[3] ( .CK(_zyM2L253_pbcMevClk12), .CE(n18), .R(n1750), .D(n4252), .Q(_zyGfifoF1_L253_s2_cbid_7[3]));
Q_FDP4EP \_zyGfifoF1_L253_s2_cbid_7_REG[2] ( .CK(_zyM2L253_pbcMevClk12), .CE(n18), .R(n1750), .D(n4251), .Q(_zyGfifoF1_L253_s2_cbid_7[2]));
Q_FDP4EP \_zyGfifoF1_L253_s2_cbid_7_REG[1] ( .CK(_zyM2L253_pbcMevClk12), .CE(n18), .R(n1750), .D(n4250), .Q(_zyGfifoF1_L253_s2_cbid_7[1]));
Q_FDP4EP \_zyGfifoF1_L253_s2_cbid_7_REG[0] ( .CK(_zyM2L253_pbcMevClk12), .CE(n18), .R(n1750), .D(n4249), .Q(_zyGfifoF1_L253_s2_cbid_7[0]));
Q_FDP4EP \seed_REG[279] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4248), .Q(seed[279]));
Q_FDP4EP \seed_REG[278] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4247), .Q(seed[278]));
Q_FDP4EP \seed_REG[277] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4246), .Q(seed[277]));
Q_FDP4EP \seed_REG[276] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4245), .Q(seed[276]));
Q_FDP4EP \seed_REG[275] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4244), .Q(seed[275]));
Q_FDP4EP \seed_REG[274] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4243), .Q(seed[274]));
Q_FDP4EP \seed_REG[273] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4242), .Q(seed[273]));
Q_FDP4EP \seed_REG[272] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4241), .Q(seed[272]));
Q_FDP4EP \seed_REG[271] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4240), .Q(seed[271]));
Q_FDP4EP \seed_REG[270] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4239), .Q(seed[270]));
Q_FDP4EP \seed_REG[269] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4238), .Q(seed[269]));
Q_FDP4EP \seed_REG[268] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4237), .Q(seed[268]));
Q_FDP4EP \seed_REG[267] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4236), .Q(seed[267]));
Q_FDP4EP \seed_REG[266] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4235), .Q(seed[266]));
Q_FDP4EP \seed_REG[265] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4234), .Q(seed[265]));
Q_FDP4EP \seed_REG[264] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4233), .Q(seed[264]));
Q_FDP4EP \seed_REG[263] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4232), .Q(seed[263]));
Q_FDP4EP \seed_REG[262] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4231), .Q(seed[262]));
Q_FDP4EP \seed_REG[261] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4230), .Q(seed[261]));
Q_FDP4EP \seed_REG[260] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4229), .Q(seed[260]));
Q_FDP4EP \seed_REG[259] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4228), .Q(seed[259]));
Q_FDP4EP \seed_REG[258] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4227), .Q(seed[258]));
Q_FDP4EP \seed_REG[257] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4226), .Q(seed[257]));
Q_FDP4EP \seed_REG[256] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4225), .Q(seed[256]));
Q_FDP4EP \seed_REG[255] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4224), .Q(seed[255]));
Q_FDP4EP \seed_REG[254] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4223), .Q(seed[254]));
Q_FDP4EP \seed_REG[253] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4222), .Q(seed[253]));
Q_FDP4EP \seed_REG[252] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4221), .Q(seed[252]));
Q_FDP4EP \seed_REG[251] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4220), .Q(seed[251]));
Q_FDP4EP \seed_REG[250] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4219), .Q(seed[250]));
Q_FDP4EP \seed_REG[249] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4218), .Q(seed[249]));
Q_FDP4EP \seed_REG[248] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4217), .Q(seed[248]));
Q_FDP4EP \seed_REG[247] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4216), .Q(seed[247]));
Q_FDP4EP \seed_REG[246] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4215), .Q(seed[246]));
Q_FDP4EP \seed_REG[245] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4214), .Q(seed[245]));
Q_FDP4EP \seed_REG[244] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4213), .Q(seed[244]));
Q_FDP4EP \seed_REG[243] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4212), .Q(seed[243]));
Q_FDP4EP \seed_REG[242] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4211), .Q(seed[242]));
Q_FDP4EP \seed_REG[241] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4210), .Q(seed[241]));
Q_FDP4EP \seed_REG[240] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4209), .Q(seed[240]));
Q_FDP4EP \seed_REG[239] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4208), .Q(seed[239]));
Q_FDP4EP \seed_REG[238] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4207), .Q(seed[238]));
Q_FDP4EP \seed_REG[237] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4206), .Q(seed[237]));
Q_FDP4EP \seed_REG[236] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4205), .Q(seed[236]));
Q_FDP4EP \seed_REG[235] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4204), .Q(seed[235]));
Q_FDP4EP \seed_REG[234] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4203), .Q(seed[234]));
Q_FDP4EP \seed_REG[233] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4202), .Q(seed[233]));
Q_FDP4EP \seed_REG[232] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4201), .Q(seed[232]));
Q_FDP4EP \seed_REG[231] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4200), .Q(seed[231]));
Q_FDP4EP \seed_REG[230] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4199), .Q(seed[230]));
Q_FDP4EP \seed_REG[229] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4198), .Q(seed[229]));
Q_FDP4EP \seed_REG[228] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4197), .Q(seed[228]));
Q_FDP4EP \seed_REG[227] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4196), .Q(seed[227]));
Q_FDP4EP \seed_REG[226] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4195), .Q(seed[226]));
Q_FDP4EP \seed_REG[225] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4194), .Q(seed[225]));
Q_FDP4EP \seed_REG[224] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4193), .Q(seed[224]));
Q_FDP4EP \seed_REG[223] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4192), .Q(seed[223]));
Q_FDP4EP \seed_REG[222] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4191), .Q(seed[222]));
Q_FDP4EP \seed_REG[221] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4190), .Q(seed[221]));
Q_FDP4EP \seed_REG[220] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4189), .Q(seed[220]));
Q_FDP4EP \seed_REG[219] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4188), .Q(seed[219]));
Q_FDP4EP \seed_REG[218] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4187), .Q(seed[218]));
Q_FDP4EP \seed_REG[217] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4186), .Q(seed[217]));
Q_FDP4EP \seed_REG[216] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4185), .Q(seed[216]));
Q_FDP4EP \seed_REG[215] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4184), .Q(seed[215]));
Q_FDP4EP \seed_REG[214] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4183), .Q(seed[214]));
Q_FDP4EP \seed_REG[213] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4182), .Q(seed[213]));
Q_FDP4EP \seed_REG[212] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4181), .Q(seed[212]));
Q_FDP4EP \seed_REG[211] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4180), .Q(seed[211]));
Q_FDP4EP \seed_REG[210] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4179), .Q(seed[210]));
Q_FDP4EP \seed_REG[209] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4178), .Q(seed[209]));
Q_FDP4EP \seed_REG[208] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4177), .Q(seed[208]));
Q_FDP4EP \seed_REG[207] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4176), .Q(seed[207]));
Q_FDP4EP \seed_REG[206] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4175), .Q(seed[206]));
Q_FDP4EP \seed_REG[205] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4174), .Q(seed[205]));
Q_FDP4EP \seed_REG[204] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4173), .Q(seed[204]));
Q_FDP4EP \seed_REG[203] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4172), .Q(seed[203]));
Q_FDP4EP \seed_REG[202] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4171), .Q(seed[202]));
Q_FDP4EP \seed_REG[201] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4170), .Q(seed[201]));
Q_FDP4EP \seed_REG[200] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4169), .Q(seed[200]));
Q_FDP4EP \seed_REG[199] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4168), .Q(seed[199]));
Q_FDP4EP \seed_REG[198] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4167), .Q(seed[198]));
Q_FDP4EP \seed_REG[197] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4166), .Q(seed[197]));
Q_FDP4EP \seed_REG[196] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4165), .Q(seed[196]));
Q_FDP4EP \seed_REG[195] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4164), .Q(seed[195]));
Q_FDP4EP \seed_REG[194] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4163), .Q(seed[194]));
Q_FDP4EP \seed_REG[193] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4162), .Q(seed[193]));
Q_FDP4EP \seed_REG[192] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4161), .Q(seed[192]));
Q_FDP4EP \seed_REG[191] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4160), .Q(seed[191]));
Q_FDP4EP \seed_REG[190] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4159), .Q(seed[190]));
Q_FDP4EP \seed_REG[189] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4158), .Q(seed[189]));
Q_FDP4EP \seed_REG[188] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4157), .Q(seed[188]));
Q_FDP4EP \seed_REG[187] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4156), .Q(seed[187]));
Q_FDP4EP \seed_REG[186] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4155), .Q(seed[186]));
Q_FDP4EP \seed_REG[185] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4154), .Q(seed[185]));
Q_FDP4EP \seed_REG[184] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4153), .Q(seed[184]));
Q_FDP4EP \seed_REG[183] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4152), .Q(seed[183]));
Q_FDP4EP \seed_REG[182] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4151), .Q(seed[182]));
Q_FDP4EP \seed_REG[181] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4150), .Q(seed[181]));
Q_FDP4EP \seed_REG[180] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4149), .Q(seed[180]));
Q_FDP4EP \seed_REG[179] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4148), .Q(seed[179]));
Q_FDP4EP \seed_REG[178] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4147), .Q(seed[178]));
Q_FDP4EP \seed_REG[177] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4146), .Q(seed[177]));
Q_FDP4EP \seed_REG[176] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4145), .Q(seed[176]));
Q_FDP4EP \seed_REG[175] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4144), .Q(seed[175]));
Q_FDP4EP \seed_REG[174] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4143), .Q(seed[174]));
Q_FDP4EP \seed_REG[173] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4142), .Q(seed[173]));
Q_FDP4EP \seed_REG[172] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4141), .Q(seed[172]));
Q_FDP4EP \seed_REG[171] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4140), .Q(seed[171]));
Q_FDP4EP \seed_REG[170] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4139), .Q(seed[170]));
Q_FDP4EP \seed_REG[169] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4138), .Q(seed[169]));
Q_FDP4EP \seed_REG[168] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4137), .Q(seed[168]));
Q_FDP4EP \seed_REG[167] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4136), .Q(seed[167]));
Q_FDP4EP \seed_REG[166] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4135), .Q(seed[166]));
Q_FDP4EP \seed_REG[165] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4134), .Q(seed[165]));
Q_FDP4EP \seed_REG[164] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4133), .Q(seed[164]));
Q_FDP4EP \seed_REG[163] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4132), .Q(seed[163]));
Q_FDP4EP \seed_REG[162] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4131), .Q(seed[162]));
Q_FDP4EP \seed_REG[161] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4130), .Q(seed[161]));
Q_FDP4EP \seed_REG[160] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4129), .Q(seed[160]));
Q_FDP4EP \seed_REG[159] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4128), .Q(seed[159]));
Q_FDP4EP \seed_REG[158] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4127), .Q(seed[158]));
Q_FDP4EP \seed_REG[157] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4126), .Q(seed[157]));
Q_FDP4EP \seed_REG[156] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4125), .Q(seed[156]));
Q_FDP4EP \seed_REG[155] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4124), .Q(seed[155]));
Q_FDP4EP \seed_REG[154] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4123), .Q(seed[154]));
Q_FDP4EP \seed_REG[153] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4122), .Q(seed[153]));
Q_FDP4EP \seed_REG[152] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4121), .Q(seed[152]));
Q_FDP4EP \seed_REG[151] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4120), .Q(seed[151]));
Q_FDP4EP \seed_REG[150] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4119), .Q(seed[150]));
Q_FDP4EP \seed_REG[149] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4118), .Q(seed[149]));
Q_FDP4EP \seed_REG[148] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4117), .Q(seed[148]));
Q_FDP4EP \seed_REG[147] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4116), .Q(seed[147]));
Q_FDP4EP \seed_REG[146] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4115), .Q(seed[146]));
Q_FDP4EP \seed_REG[145] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4114), .Q(seed[145]));
Q_FDP4EP \seed_REG[144] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4113), .Q(seed[144]));
Q_FDP4EP \seed_REG[143] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4112), .Q(seed[143]));
Q_FDP4EP \seed_REG[142] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4111), .Q(seed[142]));
Q_FDP4EP \seed_REG[141] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4110), .Q(seed[141]));
Q_FDP4EP \seed_REG[140] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4109), .Q(seed[140]));
Q_FDP4EP \seed_REG[139] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4108), .Q(seed[139]));
Q_FDP4EP \seed_REG[138] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4107), .Q(seed[138]));
Q_FDP4EP \seed_REG[137] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4106), .Q(seed[137]));
Q_FDP4EP \seed_REG[136] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4105), .Q(seed[136]));
Q_FDP4EP \seed_REG[135] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4104), .Q(seed[135]));
Q_FDP4EP \seed_REG[134] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4103), .Q(seed[134]));
Q_FDP4EP \seed_REG[133] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4102), .Q(seed[133]));
Q_FDP4EP \seed_REG[132] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4101), .Q(seed[132]));
Q_FDP4EP \seed_REG[131] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4100), .Q(seed[131]));
Q_FDP4EP \seed_REG[130] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4099), .Q(seed[130]));
Q_FDP4EP \seed_REG[129] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4098), .Q(seed[129]));
Q_FDP4EP \seed_REG[128] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4097), .Q(seed[128]));
Q_FDP4EP \seed_REG[127] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4096), .Q(seed[127]));
Q_FDP4EP \seed_REG[126] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4095), .Q(seed[126]));
Q_FDP4EP \seed_REG[125] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4094), .Q(seed[125]));
Q_FDP4EP \seed_REG[124] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4093), .Q(seed[124]));
Q_FDP4EP \seed_REG[123] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4092), .Q(seed[123]));
Q_FDP4EP \seed_REG[122] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4091), .Q(seed[122]));
Q_FDP4EP \seed_REG[121] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4090), .Q(seed[121]));
Q_FDP4EP \seed_REG[120] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4089), .Q(seed[120]));
Q_FDP4EP \seed_REG[119] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4088), .Q(seed[119]));
Q_FDP4EP \seed_REG[118] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4087), .Q(seed[118]));
Q_FDP4EP \seed_REG[117] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4086), .Q(seed[117]));
Q_FDP4EP \seed_REG[116] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4085), .Q(seed[116]));
Q_FDP4EP \seed_REG[115] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4084), .Q(seed[115]));
Q_FDP4EP \seed_REG[114] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4083), .Q(seed[114]));
Q_FDP4EP \seed_REG[113] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4082), .Q(seed[113]));
Q_FDP4EP \seed_REG[112] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4081), .Q(seed[112]));
Q_FDP4EP \seed_REG[111] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4080), .Q(seed[111]));
Q_FDP4EP \seed_REG[110] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4079), .Q(seed[110]));
Q_FDP4EP \seed_REG[109] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4078), .Q(seed[109]));
Q_FDP4EP \seed_REG[108] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4077), .Q(seed[108]));
Q_FDP4EP \seed_REG[107] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4076), .Q(seed[107]));
Q_FDP4EP \seed_REG[106] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4075), .Q(seed[106]));
Q_FDP4EP \seed_REG[105] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4074), .Q(seed[105]));
Q_FDP4EP \seed_REG[104] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4073), .Q(seed[104]));
Q_FDP4EP \seed_REG[103] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4072), .Q(seed[103]));
Q_FDP4EP \seed_REG[102] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4071), .Q(seed[102]));
Q_FDP4EP \seed_REG[101] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4070), .Q(seed[101]));
Q_FDP4EP \seed_REG[100] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4069), .Q(seed[100]));
Q_FDP4EP \seed_REG[99] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4068), .Q(seed[99]));
Q_FDP4EP \seed_REG[98] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4067), .Q(seed[98]));
Q_FDP4EP \seed_REG[97] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4066), .Q(seed[97]));
Q_FDP4EP \seed_REG[96] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4065), .Q(seed[96]));
Q_FDP4EP \seed_REG[95] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4064), .Q(seed[95]));
Q_FDP4EP \seed_REG[94] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4063), .Q(seed[94]));
Q_FDP4EP \seed_REG[93] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4062), .Q(seed[93]));
Q_FDP4EP \seed_REG[92] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4061), .Q(seed[92]));
Q_FDP4EP \seed_REG[91] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4060), .Q(seed[91]));
Q_FDP4EP \seed_REG[90] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4059), .Q(seed[90]));
Q_FDP4EP \seed_REG[89] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4058), .Q(seed[89]));
Q_FDP4EP \seed_REG[88] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4057), .Q(seed[88]));
Q_FDP4EP \seed_REG[87] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4056), .Q(seed[87]));
Q_FDP4EP \seed_REG[86] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4055), .Q(seed[86]));
Q_FDP4EP \seed_REG[85] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4054), .Q(seed[85]));
Q_FDP4EP \seed_REG[84] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4053), .Q(seed[84]));
Q_FDP4EP \seed_REG[83] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4052), .Q(seed[83]));
Q_FDP4EP \seed_REG[82] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4051), .Q(seed[82]));
Q_FDP4EP \seed_REG[81] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4050), .Q(seed[81]));
Q_FDP4EP \seed_REG[80] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4049), .Q(seed[80]));
Q_FDP4EP \seed_REG[79] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4048), .Q(seed[79]));
Q_FDP4EP \seed_REG[78] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4047), .Q(seed[78]));
Q_FDP4EP \seed_REG[77] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4046), .Q(seed[77]));
Q_FDP4EP \seed_REG[76] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4045), .Q(seed[76]));
Q_FDP4EP \seed_REG[75] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4044), .Q(seed[75]));
Q_FDP4EP \seed_REG[74] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4043), .Q(seed[74]));
Q_FDP4EP \seed_REG[73] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4042), .Q(seed[73]));
Q_FDP4EP \seed_REG[72] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4041), .Q(seed[72]));
Q_FDP4EP \seed_REG[71] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4040), .Q(seed[71]));
Q_FDP4EP \seed_REG[70] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4039), .Q(seed[70]));
Q_FDP4EP \seed_REG[69] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4038), .Q(seed[69]));
Q_FDP4EP \seed_REG[68] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4037), .Q(seed[68]));
Q_FDP4EP \seed_REG[67] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4036), .Q(seed[67]));
Q_FDP4EP \seed_REG[66] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4035), .Q(seed[66]));
Q_FDP4EP \seed_REG[65] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4034), .Q(seed[65]));
Q_FDP4EP \seed_REG[64] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4033), .Q(seed[64]));
Q_FDP4EP \seed_REG[63] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4032), .Q(seed[63]));
Q_FDP4EP \seed_REG[62] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4031), .Q(seed[62]));
Q_FDP4EP \seed_REG[61] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4030), .Q(seed[61]));
Q_FDP4EP \seed_REG[60] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4029), .Q(seed[60]));
Q_FDP4EP \seed_REG[59] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4028), .Q(seed[59]));
Q_FDP4EP \seed_REG[58] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4027), .Q(seed[58]));
Q_FDP4EP \seed_REG[57] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4026), .Q(seed[57]));
Q_FDP4EP \seed_REG[56] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4025), .Q(seed[56]));
Q_FDP4EP \seed_REG[55] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4024), .Q(seed[55]));
Q_FDP4EP \seed_REG[54] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4023), .Q(seed[54]));
Q_FDP4EP \seed_REG[53] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4022), .Q(seed[53]));
Q_FDP4EP \seed_REG[52] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4021), .Q(seed[52]));
Q_FDP4EP \seed_REG[51] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4020), .Q(seed[51]));
Q_FDP4EP \seed_REG[50] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4019), .Q(seed[50]));
Q_FDP4EP \seed_REG[49] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4018), .Q(seed[49]));
Q_FDP4EP \seed_REG[48] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4017), .Q(seed[48]));
Q_FDP4EP \seed_REG[47] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4016), .Q(seed[47]));
Q_FDP4EP \seed_REG[46] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4015), .Q(seed[46]));
Q_FDP4EP \seed_REG[45] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4014), .Q(seed[45]));
Q_FDP4EP \seed_REG[44] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4013), .Q(seed[44]));
Q_FDP4EP \seed_REG[43] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4012), .Q(seed[43]));
Q_FDP4EP \seed_REG[42] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4011), .Q(seed[42]));
Q_FDP4EP \seed_REG[41] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4010), .Q(seed[41]));
Q_FDP4EP \seed_REG[40] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4009), .Q(seed[40]));
Q_FDP4EP \seed_REG[39] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4008), .Q(seed[39]));
Q_FDP4EP \seed_REG[38] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4007), .Q(seed[38]));
Q_FDP4EP \seed_REG[37] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4006), .Q(seed[37]));
Q_FDP4EP \seed_REG[36] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4005), .Q(seed[36]));
Q_FDP4EP \seed_REG[35] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4004), .Q(seed[35]));
Q_FDP4EP \seed_REG[34] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4003), .Q(seed[34]));
Q_FDP4EP \seed_REG[33] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4002), .Q(seed[33]));
Q_FDP4EP \seed_REG[32] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4001), .Q(seed[32]));
Q_FDP4EP \seed_REG[31] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4000), .Q(seed[31]));
Q_FDP4EP \seed_REG[30] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3999), .Q(seed[30]));
Q_FDP4EP \seed_REG[29] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3998), .Q(seed[29]));
Q_FDP4EP \seed_REG[28] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3997), .Q(seed[28]));
Q_FDP4EP \seed_REG[27] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3996), .Q(seed[27]));
Q_FDP4EP \seed_REG[26] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3995), .Q(seed[26]));
Q_FDP4EP \seed_REG[25] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3994), .Q(seed[25]));
Q_FDP4EP \seed_REG[24] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3993), .Q(seed[24]));
Q_FDP4EP \seed_REG[23] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3992), .Q(seed[23]));
Q_FDP4EP \seed_REG[22] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3991), .Q(seed[22]));
Q_FDP4EP \seed_REG[21] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3990), .Q(seed[21]));
Q_FDP4EP \seed_REG[20] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3989), .Q(seed[20]));
Q_FDP4EP \seed_REG[19] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3988), .Q(seed[19]));
Q_FDP4EP \seed_REG[18] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3987), .Q(seed[18]));
Q_FDP4EP \seed_REG[17] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3986), .Q(seed[17]));
Q_FDP4EP \seed_REG[16] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3985), .Q(seed[16]));
Q_FDP4EP \seed_REG[15] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3984), .Q(seed[15]));
Q_FDP4EP \seed_REG[14] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3983), .Q(seed[14]));
Q_FDP4EP \seed_REG[13] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3982), .Q(seed[13]));
Q_FDP4EP \seed_REG[12] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3981), .Q(seed[12]));
Q_FDP4EP \seed_REG[11] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3980), .Q(seed[11]));
Q_FDP4EP \seed_REG[10] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3979), .Q(seed[10]));
Q_FDP4EP \seed_REG[9] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3978), .Q(seed[9]));
Q_FDP4EP \seed_REG[8] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3977), .Q(seed[8]));
Q_FDP4EP \seed_REG[7] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3976), .Q(seed[7]));
Q_FDP4EP \seed_REG[6] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3975), .Q(seed[6]));
Q_FDP4EP \seed_REG[5] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3974), .Q(seed[5]));
Q_FDP4EP \seed_REG[4] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3973), .Q(seed[4]));
Q_FDP4EP \seed_REG[3] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3972), .Q(seed[3]));
Q_FDP4EP \seed_REG[2] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3971), .Q(seed[2]));
Q_FDP4EP \seed_REG[1] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3970), .Q(seed[1]));
Q_FDP4EP \seed_REG[0] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n3969), .Q(seed[0]));
Q_FDP4EP \testname_REG[279] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5130), .Q(testname[279]));
Q_FDP4EP \testname_REG[278] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5129), .Q(testname[278]));
Q_FDP4EP \testname_REG[277] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5128), .Q(testname[277]));
Q_FDP4EP \testname_REG[276] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5127), .Q(testname[276]));
Q_FDP4EP \testname_REG[275] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5126), .Q(testname[275]));
Q_FDP4EP \testname_REG[274] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5125), .Q(testname[274]));
Q_FDP4EP \testname_REG[273] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5124), .Q(testname[273]));
Q_FDP4EP \testname_REG[272] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5123), .Q(testname[272]));
Q_FDP4EP \testname_REG[271] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5122), .Q(testname[271]));
Q_FDP4EP \testname_REG[270] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5121), .Q(testname[270]));
Q_FDP4EP \testname_REG[269] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5120), .Q(testname[269]));
Q_FDP4EP \testname_REG[268] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5119), .Q(testname[268]));
Q_FDP4EP \testname_REG[267] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5118), .Q(testname[267]));
Q_FDP4EP \testname_REG[266] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5117), .Q(testname[266]));
Q_FDP4EP \testname_REG[265] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5116), .Q(testname[265]));
Q_FDP4EP \testname_REG[264] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5115), .Q(testname[264]));
Q_FDP4EP \testname_REG[263] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5114), .Q(testname[263]));
Q_FDP4EP \testname_REG[262] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5113), .Q(testname[262]));
Q_FDP4EP \testname_REG[261] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5112), .Q(testname[261]));
Q_FDP4EP \testname_REG[260] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5111), .Q(testname[260]));
Q_FDP4EP \testname_REG[259] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5110), .Q(testname[259]));
Q_FDP4EP \testname_REG[258] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5109), .Q(testname[258]));
Q_FDP4EP \testname_REG[257] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5108), .Q(testname[257]));
Q_FDP4EP \testname_REG[256] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5107), .Q(testname[256]));
Q_FDP4EP \testname_REG[255] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5106), .Q(testname[255]));
Q_FDP4EP \testname_REG[254] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5105), .Q(testname[254]));
Q_FDP4EP \testname_REG[253] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5104), .Q(testname[253]));
Q_FDP4EP \testname_REG[252] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5103), .Q(testname[252]));
Q_FDP4EP \testname_REG[251] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5102), .Q(testname[251]));
Q_FDP4EP \testname_REG[250] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5101), .Q(testname[250]));
Q_FDP4EP \testname_REG[249] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5100), .Q(testname[249]));
Q_FDP4EP \testname_REG[248] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5099), .Q(testname[248]));
Q_FDP4EP \testname_REG[247] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5098), .Q(testname[247]));
Q_FDP4EP \testname_REG[246] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5097), .Q(testname[246]));
Q_FDP4EP \testname_REG[245] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5096), .Q(testname[245]));
Q_FDP4EP \testname_REG[244] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5095), .Q(testname[244]));
Q_FDP4EP \testname_REG[243] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5094), .Q(testname[243]));
Q_FDP4EP \testname_REG[242] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5093), .Q(testname[242]));
Q_FDP4EP \testname_REG[241] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5092), .Q(testname[241]));
Q_FDP4EP \testname_REG[240] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5091), .Q(testname[240]));
Q_FDP4EP \testname_REG[239] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5090), .Q(testname[239]));
Q_FDP4EP \testname_REG[238] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5089), .Q(testname[238]));
Q_FDP4EP \testname_REG[237] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5088), .Q(testname[237]));
Q_FDP4EP \testname_REG[236] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5087), .Q(testname[236]));
Q_FDP4EP \testname_REG[235] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5086), .Q(testname[235]));
Q_FDP4EP \testname_REG[234] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5085), .Q(testname[234]));
Q_FDP4EP \testname_REG[233] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5084), .Q(testname[233]));
Q_FDP4EP \testname_REG[232] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5083), .Q(testname[232]));
Q_FDP4EP \testname_REG[231] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5082), .Q(testname[231]));
Q_FDP4EP \testname_REG[230] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5081), .Q(testname[230]));
Q_FDP4EP \testname_REG[229] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5080), .Q(testname[229]));
Q_FDP4EP \testname_REG[228] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5079), .Q(testname[228]));
Q_FDP4EP \testname_REG[227] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5078), .Q(testname[227]));
Q_FDP4EP \testname_REG[226] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5077), .Q(testname[226]));
Q_FDP4EP \testname_REG[225] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5076), .Q(testname[225]));
Q_FDP4EP \testname_REG[224] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5075), .Q(testname[224]));
Q_FDP4EP \testname_REG[223] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5074), .Q(testname[223]));
Q_FDP4EP \testname_REG[222] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5073), .Q(testname[222]));
Q_FDP4EP \testname_REG[221] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5072), .Q(testname[221]));
Q_FDP4EP \testname_REG[220] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5071), .Q(testname[220]));
Q_FDP4EP \testname_REG[219] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5070), .Q(testname[219]));
Q_FDP4EP \testname_REG[218] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5069), .Q(testname[218]));
Q_FDP4EP \testname_REG[217] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5068), .Q(testname[217]));
Q_FDP4EP \testname_REG[216] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5067), .Q(testname[216]));
Q_FDP4EP \testname_REG[215] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5066), .Q(testname[215]));
Q_FDP4EP \testname_REG[214] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5065), .Q(testname[214]));
Q_FDP4EP \testname_REG[213] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5064), .Q(testname[213]));
Q_FDP4EP \testname_REG[212] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5063), .Q(testname[212]));
Q_FDP4EP \testname_REG[211] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5062), .Q(testname[211]));
Q_FDP4EP \testname_REG[210] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5061), .Q(testname[210]));
Q_FDP4EP \testname_REG[209] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5060), .Q(testname[209]));
Q_FDP4EP \testname_REG[208] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5059), .Q(testname[208]));
Q_FDP4EP \testname_REG[207] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5058), .Q(testname[207]));
Q_FDP4EP \testname_REG[206] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5057), .Q(testname[206]));
Q_FDP4EP \testname_REG[205] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5056), .Q(testname[205]));
Q_FDP4EP \testname_REG[204] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5055), .Q(testname[204]));
Q_FDP4EP \testname_REG[203] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5054), .Q(testname[203]));
Q_FDP4EP \testname_REG[202] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5053), .Q(testname[202]));
Q_FDP4EP \testname_REG[201] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5052), .Q(testname[201]));
Q_FDP4EP \testname_REG[200] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5051), .Q(testname[200]));
Q_FDP4EP \testname_REG[199] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5050), .Q(testname[199]));
Q_FDP4EP \testname_REG[198] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5049), .Q(testname[198]));
Q_FDP4EP \testname_REG[197] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5048), .Q(testname[197]));
Q_FDP4EP \testname_REG[196] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5047), .Q(testname[196]));
Q_FDP4EP \testname_REG[195] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5046), .Q(testname[195]));
Q_FDP4EP \testname_REG[194] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5045), .Q(testname[194]));
Q_FDP4EP \testname_REG[193] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5044), .Q(testname[193]));
Q_FDP4EP \testname_REG[192] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5043), .Q(testname[192]));
Q_FDP4EP \testname_REG[191] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5042), .Q(testname[191]));
Q_FDP4EP \testname_REG[190] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5041), .Q(testname[190]));
Q_FDP4EP \testname_REG[189] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5040), .Q(testname[189]));
Q_FDP4EP \testname_REG[188] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5039), .Q(testname[188]));
Q_FDP4EP \testname_REG[187] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5038), .Q(testname[187]));
Q_FDP4EP \testname_REG[186] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5037), .Q(testname[186]));
Q_FDP4EP \testname_REG[185] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5036), .Q(testname[185]));
Q_FDP4EP \testname_REG[184] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5035), .Q(testname[184]));
Q_FDP4EP \testname_REG[183] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5034), .Q(testname[183]));
Q_FDP4EP \testname_REG[182] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5033), .Q(testname[182]));
Q_FDP4EP \testname_REG[181] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5032), .Q(testname[181]));
Q_FDP4EP \testname_REG[180] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5031), .Q(testname[180]));
Q_FDP4EP \testname_REG[179] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5030), .Q(testname[179]));
Q_FDP4EP \testname_REG[178] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5029), .Q(testname[178]));
Q_FDP4EP \testname_REG[177] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5028), .Q(testname[177]));
Q_FDP4EP \testname_REG[176] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5027), .Q(testname[176]));
Q_FDP4EP \testname_REG[175] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5026), .Q(testname[175]));
Q_FDP4EP \testname_REG[174] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5025), .Q(testname[174]));
Q_FDP4EP \testname_REG[173] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5024), .Q(testname[173]));
Q_FDP4EP \testname_REG[172] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5023), .Q(testname[172]));
Q_FDP4EP \testname_REG[171] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5022), .Q(testname[171]));
Q_FDP4EP \testname_REG[170] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5021), .Q(testname[170]));
Q_FDP4EP \testname_REG[169] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5020), .Q(testname[169]));
Q_FDP4EP \testname_REG[168] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5019), .Q(testname[168]));
Q_FDP4EP \testname_REG[167] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5018), .Q(testname[167]));
Q_FDP4EP \testname_REG[166] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5017), .Q(testname[166]));
Q_FDP4EP \testname_REG[165] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5016), .Q(testname[165]));
Q_FDP4EP \testname_REG[164] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5015), .Q(testname[164]));
Q_FDP4EP \testname_REG[163] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5014), .Q(testname[163]));
Q_FDP4EP \testname_REG[162] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5013), .Q(testname[162]));
Q_FDP4EP \testname_REG[161] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5012), .Q(testname[161]));
Q_FDP4EP \testname_REG[160] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5011), .Q(testname[160]));
Q_FDP4EP \testname_REG[159] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5010), .Q(testname[159]));
Q_FDP4EP \testname_REG[158] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5009), .Q(testname[158]));
Q_FDP4EP \testname_REG[157] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5008), .Q(testname[157]));
Q_FDP4EP \testname_REG[156] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5007), .Q(testname[156]));
Q_FDP4EP \testname_REG[155] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5006), .Q(testname[155]));
Q_FDP4EP \testname_REG[154] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5005), .Q(testname[154]));
Q_FDP4EP \testname_REG[153] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5004), .Q(testname[153]));
Q_FDP4EP \testname_REG[152] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5003), .Q(testname[152]));
Q_FDP4EP \testname_REG[151] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5002), .Q(testname[151]));
Q_FDP4EP \testname_REG[150] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5001), .Q(testname[150]));
Q_FDP4EP \testname_REG[149] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n5000), .Q(testname[149]));
Q_FDP4EP \testname_REG[148] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4999), .Q(testname[148]));
Q_FDP4EP \testname_REG[147] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4998), .Q(testname[147]));
Q_FDP4EP \testname_REG[146] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4997), .Q(testname[146]));
Q_FDP4EP \testname_REG[145] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4996), .Q(testname[145]));
Q_FDP4EP \testname_REG[144] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4995), .Q(testname[144]));
Q_FDP4EP \testname_REG[143] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4994), .Q(testname[143]));
Q_FDP4EP \testname_REG[142] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4993), .Q(testname[142]));
Q_FDP4EP \testname_REG[141] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4992), .Q(testname[141]));
Q_FDP4EP \testname_REG[140] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4991), .Q(testname[140]));
Q_FDP4EP \testname_REG[139] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4990), .Q(testname[139]));
Q_FDP4EP \testname_REG[138] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4989), .Q(testname[138]));
Q_FDP4EP \testname_REG[137] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4988), .Q(testname[137]));
Q_FDP4EP \testname_REG[136] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4987), .Q(testname[136]));
Q_FDP4EP \testname_REG[135] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4986), .Q(testname[135]));
Q_FDP4EP \testname_REG[134] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4985), .Q(testname[134]));
Q_FDP4EP \testname_REG[133] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4984), .Q(testname[133]));
Q_FDP4EP \testname_REG[132] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4983), .Q(testname[132]));
Q_FDP4EP \testname_REG[131] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4982), .Q(testname[131]));
Q_FDP4EP \testname_REG[130] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4981), .Q(testname[130]));
Q_FDP4EP \testname_REG[129] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4980), .Q(testname[129]));
Q_FDP4EP \testname_REG[128] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4979), .Q(testname[128]));
Q_FDP4EP \testname_REG[127] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4978), .Q(testname[127]));
Q_FDP4EP \testname_REG[126] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4977), .Q(testname[126]));
Q_FDP4EP \testname_REG[125] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4976), .Q(testname[125]));
Q_FDP4EP \testname_REG[124] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4975), .Q(testname[124]));
Q_FDP4EP \testname_REG[123] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4974), .Q(testname[123]));
Q_FDP4EP \testname_REG[122] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4973), .Q(testname[122]));
Q_FDP4EP \testname_REG[121] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4972), .Q(testname[121]));
Q_FDP4EP \testname_REG[120] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4971), .Q(testname[120]));
Q_FDP4EP \testname_REG[119] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4970), .Q(testname[119]));
Q_FDP4EP \testname_REG[118] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4969), .Q(testname[118]));
Q_FDP4EP \testname_REG[117] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4968), .Q(testname[117]));
Q_FDP4EP \testname_REG[116] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4967), .Q(testname[116]));
Q_FDP4EP \testname_REG[115] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4966), .Q(testname[115]));
Q_FDP4EP \testname_REG[114] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4965), .Q(testname[114]));
Q_FDP4EP \testname_REG[113] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4964), .Q(testname[113]));
Q_FDP4EP \testname_REG[112] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4963), .Q(testname[112]));
Q_FDP4EP \testname_REG[111] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4962), .Q(testname[111]));
Q_FDP4EP \testname_REG[110] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4961), .Q(testname[110]));
Q_FDP4EP \testname_REG[109] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4960), .Q(testname[109]));
Q_FDP4EP \testname_REG[108] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4959), .Q(testname[108]));
Q_FDP4EP \testname_REG[107] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4958), .Q(testname[107]));
Q_FDP4EP \testname_REG[106] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4957), .Q(testname[106]));
Q_FDP4EP \testname_REG[105] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4956), .Q(testname[105]));
Q_FDP4EP \testname_REG[104] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4955), .Q(testname[104]));
Q_FDP4EP \testname_REG[103] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4954), .Q(testname[103]));
Q_FDP4EP \testname_REG[102] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4953), .Q(testname[102]));
Q_FDP4EP \testname_REG[101] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4952), .Q(testname[101]));
Q_FDP4EP \testname_REG[100] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4951), .Q(testname[100]));
Q_FDP4EP \testname_REG[99] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4950), .Q(testname[99]));
Q_FDP4EP \testname_REG[98] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4949), .Q(testname[98]));
Q_FDP4EP \testname_REG[97] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4948), .Q(testname[97]));
Q_FDP4EP \testname_REG[96] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4947), .Q(testname[96]));
Q_FDP4EP \testname_REG[95] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4946), .Q(testname[95]));
Q_FDP4EP \testname_REG[94] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4945), .Q(testname[94]));
Q_FDP4EP \testname_REG[93] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4944), .Q(testname[93]));
Q_FDP4EP \testname_REG[92] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4943), .Q(testname[92]));
Q_FDP4EP \testname_REG[91] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4942), .Q(testname[91]));
Q_FDP4EP \testname_REG[90] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4941), .Q(testname[90]));
Q_FDP4EP \testname_REG[89] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4940), .Q(testname[89]));
Q_FDP4EP \testname_REG[88] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4939), .Q(testname[88]));
Q_FDP4EP \testname_REG[87] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4938), .Q(testname[87]));
Q_FDP4EP \testname_REG[86] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4937), .Q(testname[86]));
Q_FDP4EP \testname_REG[85] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4936), .Q(testname[85]));
Q_FDP4EP \testname_REG[84] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4935), .Q(testname[84]));
Q_FDP4EP \testname_REG[83] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4934), .Q(testname[83]));
Q_FDP4EP \testname_REG[82] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4933), .Q(testname[82]));
Q_FDP4EP \testname_REG[81] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4932), .Q(testname[81]));
Q_FDP4EP \testname_REG[80] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4931), .Q(testname[80]));
Q_FDP4EP \testname_REG[79] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4930), .Q(testname[79]));
Q_FDP4EP \testname_REG[78] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4929), .Q(testname[78]));
Q_FDP4EP \testname_REG[77] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4928), .Q(testname[77]));
Q_FDP4EP \testname_REG[76] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4927), .Q(testname[76]));
Q_FDP4EP \testname_REG[75] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4926), .Q(testname[75]));
Q_FDP4EP \testname_REG[74] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4925), .Q(testname[74]));
Q_FDP4EP \testname_REG[73] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4924), .Q(testname[73]));
Q_FDP4EP \testname_REG[72] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4923), .Q(testname[72]));
Q_FDP4EP \testname_REG[71] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4922), .Q(testname[71]));
Q_FDP4EP \testname_REG[70] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4921), .Q(testname[70]));
Q_FDP4EP \testname_REG[69] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4920), .Q(testname[69]));
Q_FDP4EP \testname_REG[68] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4919), .Q(testname[68]));
Q_FDP4EP \testname_REG[67] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4918), .Q(testname[67]));
Q_FDP4EP \testname_REG[66] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4917), .Q(testname[66]));
Q_FDP4EP \testname_REG[65] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4916), .Q(testname[65]));
Q_FDP4EP \testname_REG[64] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4915), .Q(testname[64]));
Q_FDP4EP \testname_REG[63] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4914), .Q(testname[63]));
Q_FDP4EP \testname_REG[62] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4913), .Q(testname[62]));
Q_FDP4EP \testname_REG[61] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4912), .Q(testname[61]));
Q_FDP4EP \testname_REG[60] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4911), .Q(testname[60]));
Q_FDP4EP \testname_REG[59] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4910), .Q(testname[59]));
Q_FDP4EP \testname_REG[58] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4909), .Q(testname[58]));
Q_FDP4EP \testname_REG[57] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4908), .Q(testname[57]));
Q_FDP4EP \testname_REG[56] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4907), .Q(testname[56]));
Q_FDP4EP \testname_REG[55] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4906), .Q(testname[55]));
Q_FDP4EP \testname_REG[54] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4905), .Q(testname[54]));
Q_FDP4EP \testname_REG[53] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4904), .Q(testname[53]));
Q_FDP4EP \testname_REG[52] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4903), .Q(testname[52]));
Q_FDP4EP \testname_REG[51] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4902), .Q(testname[51]));
Q_FDP4EP \testname_REG[50] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4901), .Q(testname[50]));
Q_FDP4EP \testname_REG[49] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4900), .Q(testname[49]));
Q_FDP4EP \testname_REG[48] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4899), .Q(testname[48]));
Q_FDP4EP \testname_REG[47] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4898), .Q(testname[47]));
Q_FDP4EP \testname_REG[46] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4897), .Q(testname[46]));
Q_FDP4EP \testname_REG[45] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4896), .Q(testname[45]));
Q_FDP4EP \testname_REG[44] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4895), .Q(testname[44]));
Q_FDP4EP \testname_REG[43] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4894), .Q(testname[43]));
Q_FDP4EP \testname_REG[42] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4893), .Q(testname[42]));
Q_FDP4EP \testname_REG[41] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4892), .Q(testname[41]));
Q_FDP4EP \testname_REG[40] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4891), .Q(testname[40]));
Q_FDP4EP \testname_REG[39] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4890), .Q(testname[39]));
Q_FDP4EP \testname_REG[38] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4889), .Q(testname[38]));
Q_FDP4EP \testname_REG[37] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4888), .Q(testname[37]));
Q_FDP4EP \testname_REG[36] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4887), .Q(testname[36]));
Q_FDP4EP \testname_REG[35] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4886), .Q(testname[35]));
Q_FDP4EP \testname_REG[34] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4885), .Q(testname[34]));
Q_FDP4EP \testname_REG[33] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4884), .Q(testname[33]));
Q_FDP4EP \testname_REG[32] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4883), .Q(testname[32]));
Q_FDP4EP \testname_REG[31] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4882), .Q(testname[31]));
Q_FDP4EP \testname_REG[30] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4881), .Q(testname[30]));
Q_FDP4EP \testname_REG[29] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4880), .Q(testname[29]));
Q_FDP4EP \testname_REG[28] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4879), .Q(testname[28]));
Q_FDP4EP \testname_REG[27] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4878), .Q(testname[27]));
Q_FDP4EP \testname_REG[26] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4877), .Q(testname[26]));
Q_FDP4EP \testname_REG[25] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4876), .Q(testname[25]));
Q_FDP4EP \testname_REG[24] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4875), .Q(testname[24]));
Q_FDP4EP \testname_REG[23] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4874), .Q(testname[23]));
Q_FDP4EP \testname_REG[22] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4873), .Q(testname[22]));
Q_FDP4EP \testname_REG[21] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4872), .Q(testname[21]));
Q_FDP4EP \testname_REG[20] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4871), .Q(testname[20]));
Q_FDP4EP \testname_REG[19] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4870), .Q(testname[19]));
Q_FDP4EP \testname_REG[18] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4869), .Q(testname[18]));
Q_FDP4EP \testname_REG[17] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4868), .Q(testname[17]));
Q_FDP4EP \testname_REG[16] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4867), .Q(testname[16]));
Q_FDP4EP \testname_REG[15] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4866), .Q(testname[15]));
Q_FDP4EP \testname_REG[14] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4865), .Q(testname[14]));
Q_FDP4EP \testname_REG[13] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4864), .Q(testname[13]));
Q_FDP4EP \testname_REG[12] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4863), .Q(testname[12]));
Q_FDP4EP \testname_REG[11] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4862), .Q(testname[11]));
Q_FDP4EP \testname_REG[10] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4861), .Q(testname[10]));
Q_FDP4EP \testname_REG[9] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4860), .Q(testname[9]));
Q_FDP4EP \testname_REG[8] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4859), .Q(testname[8]));
Q_FDP4EP \testname_REG[7] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4858), .Q(testname[7]));
Q_FDP4EP \testname_REG[6] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4857), .Q(testname[6]));
Q_FDP4EP \testname_REG[5] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4856), .Q(testname[5]));
Q_FDP4EP \testname_REG[4] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4855), .Q(testname[4]));
Q_FDP4EP \testname_REG[3] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4854), .Q(testname[3]));
Q_FDP4EP \testname_REG[2] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4853), .Q(testname[2]));
Q_FDP4EP \testname_REG[1] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4852), .Q(testname[1]));
Q_FDP4EP \testname_REG[0] ( .CK(_zyM2L253_pbcMevClk12), .CE(n5321), .R(n1750), .D(n4851), .Q(testname[0]));
Q_INV U9568 ( .A(n5296), .Z(n17));
Q_FDP4EP \_zyM2L273_pbcT0_REG[31] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5260), .Q(_zyM2L273_pbcT0[31]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[30] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5259), .Q(_zyM2L273_pbcT0[30]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[29] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5258), .Q(_zyM2L273_pbcT0[29]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[28] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5257), .Q(_zyM2L273_pbcT0[28]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[27] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5256), .Q(_zyM2L273_pbcT0[27]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[26] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5255), .Q(_zyM2L273_pbcT0[26]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[25] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5254), .Q(_zyM2L273_pbcT0[25]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[24] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5253), .Q(_zyM2L273_pbcT0[24]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[23] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5252), .Q(_zyM2L273_pbcT0[23]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[22] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5251), .Q(_zyM2L273_pbcT0[22]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[21] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5250), .Q(_zyM2L273_pbcT0[21]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[20] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5249), .Q(_zyM2L273_pbcT0[20]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[19] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5248), .Q(_zyM2L273_pbcT0[19]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[18] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5247), .Q(_zyM2L273_pbcT0[18]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[17] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5246), .Q(_zyM2L273_pbcT0[17]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[16] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5245), .Q(_zyM2L273_pbcT0[16]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[15] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5244), .Q(_zyM2L273_pbcT0[15]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[14] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5243), .Q(_zyM2L273_pbcT0[14]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[13] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5242), .Q(_zyM2L273_pbcT0[13]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[12] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5241), .Q(_zyM2L273_pbcT0[12]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[11] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5240), .Q(_zyM2L273_pbcT0[11]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[10] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5239), .Q(_zyM2L273_pbcT0[10]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[9] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5238), .Q(_zyM2L273_pbcT0[9]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[8] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5237), .Q(_zyM2L273_pbcT0[8]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[7] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5236), .Q(_zyM2L273_pbcT0[7]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[6] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5235), .Q(_zyM2L273_pbcT0[6]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[5] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5234), .Q(_zyM2L273_pbcT0[5]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[4] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5233), .Q(_zyM2L273_pbcT0[4]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[3] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5232), .Q(_zyM2L273_pbcT0[3]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[2] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5231), .Q(_zyM2L273_pbcT0[2]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[1] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5230), .Q(_zyM2L273_pbcT0[1]));
Q_FDP4EP \_zyM2L273_pbcT0_REG[0] ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5229), .Q(_zyM2L273_pbcT0[0]));
Q_INV U9601 ( .A(_zyM2L273_pbcT0[0]), .Z(n3886));
Q_INV U9602 ( .A(n5306), .Z(n16));
Q_FDP4EP \_zyM2L286_pbcT1_REG[31] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5227), .Q(_zyM2L286_pbcT1[31]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[30] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5226), .Q(_zyM2L286_pbcT1[30]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[29] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5225), .Q(_zyM2L286_pbcT1[29]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[28] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5224), .Q(_zyM2L286_pbcT1[28]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[27] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5223), .Q(_zyM2L286_pbcT1[27]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[26] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5222), .Q(_zyM2L286_pbcT1[26]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[25] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5221), .Q(_zyM2L286_pbcT1[25]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[24] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5220), .Q(_zyM2L286_pbcT1[24]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[23] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5219), .Q(_zyM2L286_pbcT1[23]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[22] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5218), .Q(_zyM2L286_pbcT1[22]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[21] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5217), .Q(_zyM2L286_pbcT1[21]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[20] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5216), .Q(_zyM2L286_pbcT1[20]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[19] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5215), .Q(_zyM2L286_pbcT1[19]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[18] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5214), .Q(_zyM2L286_pbcT1[18]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[17] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5213), .Q(_zyM2L286_pbcT1[17]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[16] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5212), .Q(_zyM2L286_pbcT1[16]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[15] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5211), .Q(_zyM2L286_pbcT1[15]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[14] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5210), .Q(_zyM2L286_pbcT1[14]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[13] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5209), .Q(_zyM2L286_pbcT1[13]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[12] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5208), .Q(_zyM2L286_pbcT1[12]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[11] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5207), .Q(_zyM2L286_pbcT1[11]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[10] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5206), .Q(_zyM2L286_pbcT1[10]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[9] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5205), .Q(_zyM2L286_pbcT1[9]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[8] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5204), .Q(_zyM2L286_pbcT1[8]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[7] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5203), .Q(_zyM2L286_pbcT1[7]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[6] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5202), .Q(_zyM2L286_pbcT1[6]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[5] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5201), .Q(_zyM2L286_pbcT1[5]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[4] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5200), .Q(_zyM2L286_pbcT1[4]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[3] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5199), .Q(_zyM2L286_pbcT1[3]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[2] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5198), .Q(_zyM2L286_pbcT1[2]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[1] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5197), .Q(_zyM2L286_pbcT1[1]));
Q_FDP4EP \_zyM2L286_pbcT1_REG[0] ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5196), .Q(_zyM2L286_pbcT1[0]));
Q_INV U9635 ( .A(_zyM2L286_pbcT1[0]), .Z(n3804));
Q_INV U9636 ( .A(n5308), .Z(n15));
Q_FDP4EP \_zyM2L292_pbcT2_REG[31] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5195), .Q(_zyM2L292_pbcT2[31]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[30] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5194), .Q(_zyM2L292_pbcT2[30]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[29] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5193), .Q(_zyM2L292_pbcT2[29]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[28] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5192), .Q(_zyM2L292_pbcT2[28]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[27] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5191), .Q(_zyM2L292_pbcT2[27]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[26] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5190), .Q(_zyM2L292_pbcT2[26]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[25] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5189), .Q(_zyM2L292_pbcT2[25]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[24] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5188), .Q(_zyM2L292_pbcT2[24]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[23] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5187), .Q(_zyM2L292_pbcT2[23]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[22] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5186), .Q(_zyM2L292_pbcT2[22]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[21] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5185), .Q(_zyM2L292_pbcT2[21]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[20] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5184), .Q(_zyM2L292_pbcT2[20]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[19] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5183), .Q(_zyM2L292_pbcT2[19]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[18] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5182), .Q(_zyM2L292_pbcT2[18]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[17] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5181), .Q(_zyM2L292_pbcT2[17]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[16] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5180), .Q(_zyM2L292_pbcT2[16]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[15] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5179), .Q(_zyM2L292_pbcT2[15]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[14] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5178), .Q(_zyM2L292_pbcT2[14]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[13] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5177), .Q(_zyM2L292_pbcT2[13]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[12] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5176), .Q(_zyM2L292_pbcT2[12]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[11] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5175), .Q(_zyM2L292_pbcT2[11]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[10] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5174), .Q(_zyM2L292_pbcT2[10]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[9] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5173), .Q(_zyM2L292_pbcT2[9]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[8] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5172), .Q(_zyM2L292_pbcT2[8]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[7] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5171), .Q(_zyM2L292_pbcT2[7]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[6] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5170), .Q(_zyM2L292_pbcT2[6]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[5] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5169), .Q(_zyM2L292_pbcT2[5]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[4] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5168), .Q(_zyM2L292_pbcT2[4]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[3] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5167), .Q(_zyM2L292_pbcT2[3]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[2] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5166), .Q(_zyM2L292_pbcT2[2]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[1] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5165), .Q(_zyM2L292_pbcT2[1]));
Q_FDP4EP \_zyM2L292_pbcT2_REG[0] ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5164), .Q(_zyM2L292_pbcT2[0]));
Q_INV U9669 ( .A(_zyM2L292_pbcT2[0]), .Z(n3722));
Q_INV U9670 ( .A(n5283), .Z(n14));
Q_FDP4EP \_zyM2L299_pbcT3_REG[31] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5162), .Q(_zyM2L299_pbcT3[31]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[30] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5161), .Q(_zyM2L299_pbcT3[30]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[29] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5160), .Q(_zyM2L299_pbcT3[29]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[28] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5159), .Q(_zyM2L299_pbcT3[28]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[27] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5158), .Q(_zyM2L299_pbcT3[27]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[26] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5157), .Q(_zyM2L299_pbcT3[26]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[25] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5156), .Q(_zyM2L299_pbcT3[25]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[24] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5155), .Q(_zyM2L299_pbcT3[24]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[23] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5154), .Q(_zyM2L299_pbcT3[23]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[22] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5153), .Q(_zyM2L299_pbcT3[22]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[21] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5152), .Q(_zyM2L299_pbcT3[21]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[20] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5151), .Q(_zyM2L299_pbcT3[20]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[19] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5150), .Q(_zyM2L299_pbcT3[19]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[18] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5149), .Q(_zyM2L299_pbcT3[18]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[17] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5148), .Q(_zyM2L299_pbcT3[17]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[16] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5147), .Q(_zyM2L299_pbcT3[16]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[15] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5146), .Q(_zyM2L299_pbcT3[15]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[14] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5145), .Q(_zyM2L299_pbcT3[14]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[13] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5144), .Q(_zyM2L299_pbcT3[13]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[12] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5143), .Q(_zyM2L299_pbcT3[12]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[11] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5142), .Q(_zyM2L299_pbcT3[11]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[10] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5141), .Q(_zyM2L299_pbcT3[10]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[9] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5140), .Q(_zyM2L299_pbcT3[9]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[8] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5139), .Q(_zyM2L299_pbcT3[8]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[7] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5138), .Q(_zyM2L299_pbcT3[7]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[6] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5137), .Q(_zyM2L299_pbcT3[6]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[5] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5136), .Q(_zyM2L299_pbcT3[5]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[4] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5135), .Q(_zyM2L299_pbcT3[4]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[3] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5134), .Q(_zyM2L299_pbcT3[3]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[2] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5133), .Q(_zyM2L299_pbcT3[2]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[1] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5132), .Q(_zyM2L299_pbcT3[1]));
Q_FDP4EP \_zyM2L299_pbcT3_REG[0] ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5131), .Q(_zyM2L299_pbcT3[0]));
Q_INV U9703 ( .A(_zyM2L299_pbcT3[0]), .Z(n3640));
Q_FDP4EP rst_n_REG  ( .CK(_zyM2L253_pbcMevClk12), .CE(n18), .R(n1750), .D(_zyM2L253_pbcFsm2_s[1]), .Q(rst_n));
Q_FDP4EP \_zyGfifoF0_L253_s4_len_6_REG[11] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n1750), .Q(_zyGfifoF0_L253_s4_len_6[11]));
Q_FDP4EP \_zyGfifoF0_L253_s4_len_6_REG[10] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n1750), .Q(_zyGfifoF0_L253_s4_len_6[10]));
Q_FDP4EP \_zyGfifoF0_L253_s4_len_6_REG[9] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n1750), .Q(_zyGfifoF0_L253_s4_len_6[9]));
Q_FDP4EP \_zyGfifoF0_L253_s4_len_6_REG[8] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n1750), .Q(_zyGfifoF0_L253_s4_len_6[8]));
Q_FDP4EP \_zyGfifoF0_L253_s4_len_6_REG[7] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n1750), .Q(_zyGfifoF0_L253_s4_len_6[7]));
Q_FDP4EP \_zyGfifoF0_L253_s4_len_6_REG[6] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n1750), .Q(_zyGfifoF0_L253_s4_len_6[6]));
Q_FDP4EP \_zyGfifoF0_L253_s4_len_6_REG[5] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n1750), .Q(_zyGfifoF0_L253_s4_len_6[5]));
Q_FDP4EP \_zyGfifoF0_L253_s4_len_6_REG[4] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n5326), .Q(_zyGfifoF0_L253_s4_len_6[4]));
Q_FDP4EP \_zyGfifoF0_L253_s4_len_6_REG[3] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n1750), .Q(_zyGfifoF0_L253_s4_len_6[3]));
Q_FDP4EP \_zyGfifoF0_L253_s4_len_6_REG[2] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n1750), .Q(_zyGfifoF0_L253_s4_len_6[2]));
Q_FDP4EP \_zyGfifoF0_L253_s4_len_6_REG[1] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n5326), .Q(_zyGfifoF0_L253_s4_len_6[1]));
Q_FDP4EP \_zyGfifoF0_L253_s4_len_6_REG[0] ( .CK(_zyM2L253_pbcMevClk12), .CE(n19), .R(n1750), .D(n1750), .Q(_zyGfifoF0_L253_s4_len_6[0]));
Q_INV U9717 ( .A(n5304), .Z(n13));
Q_FDP4EP _zyM2L253_pbcCapEn5_REG  ( .CK(_zyM2L253_pbcMevClk12), .CE(n13), .R(n1750), .D(_zyM2L253_pbcFsm2_s[1]), .Q(_zyM2L253_pbcCapEn5));
Q_FDP4EP _zyM2L274_pbcCapEn6_REG  ( .CK(_zyM2L253_pbcMevClk12), .CE(n17), .R(n1750), .D(n5329), .Q(_zyM2L274_pbcCapEn6));
Q_FDP4EP _zyM2L287_pbcCapEn7_REG  ( .CK(_zyM2L253_pbcMevClk12), .CE(n16), .R(n1750), .D(n5328), .Q(_zyM2L287_pbcCapEn7));
Q_FDP4EP _zyM2L293_pbcCapEn8_REG  ( .CK(_zyM2L253_pbcMevClk12), .CE(n15), .R(n1750), .D(n5327), .Q(_zyM2L293_pbcCapEn8));
Q_INV U9722 ( .A(n5312), .Z(n12));
Q_FDP4EP _zyM2L295_pbcCapEn9_REG  ( .CK(_zyM2L253_pbcMevClk12), .CE(n12), .R(n1750), .D(_zyM2L253_pbcFsm2_s[0]), .Q(_zyM2L295_pbcCapEn9));
Q_INV U9724 ( .A(n5313), .Z(n11));
Q_FDP4EP _zyM2L364_pbcCapEn10_REG  ( .CK(_zyM2L253_pbcMevClk12), .CE(n11), .R(n1750), .D(n5326), .Q(_zyM2L364_pbcCapEn10));
Q_FDP4EP _zyM2L300_pbcCapEn11_REG  ( .CK(_zyM2L253_pbcMevClk12), .CE(n14), .R(n1750), .D(n5325), .Q(_zyM2L300_pbcCapEn11));
Q_INV U9727 ( .A(n5314), .Z(n10));
Q_FDP4EP \_zyM2L253_pbcFsm2_s_REG[2] ( .CK(_zyM2L253_pbcMevClk12), .CE(n10), .R(n1750), .D(n5267), .Q(_zyM2L253_pbcFsm2_s[2]));
Q_INV U9729 ( .A(_zyM2L253_pbcFsm2_s[2]), .Z(n5276));
Q_FDP4EP \_zyM2L253_pbcFsm2_s_REG[1] ( .CK(_zyM2L253_pbcMevClk12), .CE(n10), .R(n1750), .D(n5263), .Q(_zyM2L253_pbcFsm2_s[1]));
Q_INV U9731 ( .A(_zyM2L253_pbcFsm2_s[1]), .Z(n5330));
Q_FDP4EP \_zyM2L253_pbcFsm2_s_REG[0] ( .CK(_zyM2L253_pbcMevClk12), .CE(n10), .R(n1750), .D(n5262), .Q(_zyM2L253_pbcFsm2_s[0]));
Q_INV U9733 ( .A(_zyM2L253_pbcFsm2_s[0]), .Z(n5163));
Q_INV U9734 ( .A(n5316), .Z(n9));
Q_FDP4EP _zyM2L253_pbcEn14_REG  ( .CK(_zyM2L253_pbcMevClk12), .CE(n9), .R(n1750), .D(n5271), .Q(_zyM2L253_pbcEn14));
Q_INV U9736 ( .A(_zygsfis_get_config_data_ack[4]), .Z(n8));
Q_FDP4EP \_zygsfis_get_config_data_ack_REG[4] ( .CK(_zySfifoF0_call), .CE(n5340), .R(n1750), .D(n8), .Q(_zygsfis_get_config_data_ack[4]));
Q_INV U9738 ( .A(_zygsfis_get_config_data_wptr[4]), .Z(n7));
Q_FDP4EP \_zygsfis_get_config_data_wptr_REG[4] ( .CK(_zySfifoF1_call), .CE(n5347), .R(n1750), .D(n7), .Q(_zygsfis_get_config_data_wptr[4]));
Q_INV U9740 ( .A(_zygsfis_ib_service_data_ack[4]), .Z(n6));
Q_FDP4EP \_zygsfis_ib_service_data_ack_REG[4] ( .CK(_zySfifoF2_call), .CE(n5354), .R(n1750), .D(n6), .Q(_zygsfis_ib_service_data_ack[4]));
Q_INV U9742 ( .A(_zygsfis_ib_service_data_wptr[4]), .Z(n5));
Q_FDP4EP \_zygsfis_ib_service_data_wptr_REG[4] ( .CK(_zySfifoF3_call), .CE(n5361), .R(n1750), .D(n5), .Q(_zygsfis_ib_service_data_wptr[4]));
Q_INV U9744 ( .A(_zygsfis_ob_service_data_ack[4]), .Z(n4));
Q_FDP4EP \_zygsfis_ob_service_data_ack_REG[4] ( .CK(_zySfifoF4_call), .CE(n5368), .R(n1750), .D(n4), .Q(_zygsfis_ob_service_data_ack[4]));
Q_INV U9746 ( .A(_zygsfis_ob_service_data_wptr[4]), .Z(n3));
Q_FDP4EP \_zygsfis_ob_service_data_wptr_REG[4] ( .CK(_zySfifoF5_call), .CE(n5375), .R(n1750), .D(n3), .Q(_zygsfis_ob_service_data_wptr[4]));
Q_FDP4EP \_zzM2_bcBehEval_REG[31] ( .CK(_zzM2_bcBehEvalClk), .CE(n5456), .R(n1750), .D(_zzM2_bcBehHalt), .Q(_zzM2_bcBehEval[31]));
Q_INV U9749 ( .A(_zzM2_bcBehEval[30]), .Z(n2));
Q_FDP4EP \_zzM2_bcBehEval_REG[30] ( .CK(_zzM2_bcBehEvalClk), .CE(n5876), .R(n1750), .D(n2), .Q(_zzM2_bcBehEval[30]));
Q_FDP4EP \_zzM2_bcBehEval_REG[29] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n5454), .Q(_zzM2_bcBehEval[29]));
Q_FDP4EP \_zzM2_bcBehEval_REG[28] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n5452), .Q(_zzM2_bcBehEval[28]));
Q_FDP4EP \_zzM2_bcBehEval_REG[27] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n5450), .Q(_zzM2_bcBehEval[27]));
Q_FDP4EP \_zzM2_bcBehEval_REG[26] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n5448), .Q(_zzM2_bcBehEval[26]));
Q_FDP4EP \_zzM2_bcBehEval_REG[25] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n5446), .Q(_zzM2_bcBehEval[25]));
Q_FDP4EP \_zzM2_bcBehEval_REG[24] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n5444), .Q(_zzM2_bcBehEval[24]));
Q_FDP4EP \_zzM2_bcBehEval_REG[23] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n5442), .Q(_zzM2_bcBehEval[23]));
Q_FDP4EP \_zzM2_bcBehEval_REG[22] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n5440), .Q(_zzM2_bcBehEval[22]));
Q_FDP4EP \_zzM2_bcBehEval_REG[21] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n5438), .Q(_zzM2_bcBehEval[21]));
Q_FDP4EP \_zzM2_bcBehEval_REG[20] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n5436), .Q(_zzM2_bcBehEval[20]));
Q_FDP4EP \_zzM2_bcBehEval_REG[19] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n5434), .Q(_zzM2_bcBehEval[19]));
Q_FDP4EP \_zzM2_bcBehEval_REG[18] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n5432), .Q(_zzM2_bcBehEval[18]));
Q_FDP4EP \_zzM2_bcBehEval_REG[17] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n5430), .Q(_zzM2_bcBehEval[17]));
Q_FDP4EP \_zzM2_bcBehEval_REG[16] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n5428), .Q(_zzM2_bcBehEval[16]));
Q_FDP4EP \_zzM2_bcBehEval_REG[15] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n5426), .Q(_zzM2_bcBehEval[15]));
Q_FDP4EP \_zzM2_bcBehEval_REG[14] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n5424), .Q(_zzM2_bcBehEval[14]));
Q_FDP4EP \_zzM2_bcBehEval_REG[13] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n5422), .Q(_zzM2_bcBehEval[13]));
Q_FDP4EP \_zzM2_bcBehEval_REG[12] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n5420), .Q(_zzM2_bcBehEval[12]));
Q_FDP4EP \_zzM2_bcBehEval_REG[11] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n5418), .Q(_zzM2_bcBehEval[11]));
Q_FDP4EP \_zzM2_bcBehEval_REG[10] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n5416), .Q(_zzM2_bcBehEval[10]));
Q_FDP4EP \_zzM2_bcBehEval_REG[9] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n5414), .Q(_zzM2_bcBehEval[9]));
Q_FDP4EP \_zzM2_bcBehEval_REG[8] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n5412), .Q(_zzM2_bcBehEval[8]));
Q_FDP4EP \_zzM2_bcBehEval_REG[7] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n5410), .Q(_zzM2_bcBehEval[7]));
Q_FDP4EP \_zzM2_bcBehEval_REG[6] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n5408), .Q(_zzM2_bcBehEval[6]));
Q_FDP4EP \_zzM2_bcBehEval_REG[5] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n5406), .Q(_zzM2_bcBehEval[5]));
Q_FDP4EP \_zzM2_bcBehEval_REG[4] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n5404), .Q(_zzM2_bcBehEval[4]));
Q_FDP4EP \_zzM2_bcBehEval_REG[3] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n5402), .Q(_zzM2_bcBehEval[3]));
Q_FDP4EP \_zzM2_bcBehEval_REG[2] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n5400), .Q(_zzM2_bcBehEval[2]));
Q_FDP4EP \_zzM2_bcBehEval_REG[1] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n5398), .Q(_zzM2_bcBehEval[1]));
Q_INV U9780 ( .A(_zzM2_bcBehEval[0]), .Z(n1));
Q_FDP4EP \_zzM2_bcBehEval_REG[0] ( .CK(_zzM2_bcBehEvalClk), .CE(n5457), .R(n1750), .D(n1), .Q(_zzM2_bcBehEval[0]));
`ifdef CBV

reg [71:0] _zygsfis_get_config_data_fifo [0:31];
initial begin: U9782
  integer i;
  for (i=0; i<=31; i=i+1) _zygsfis_get_config_data_fifo[i] =
`ifdef CBV_MEM_INIT1
  {72{1'b1}};
`else
  72'b0;
`endif
end
reg [71:0] n5887;
assign {n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122} = n5887; 
always @(n5512 or n5511 or n5510 or n5509 or n5508
 or n5584 or n5583 or n5582 or n5581 or n5580 or n5579 or n5578 or n5577
 or n5576 or n5575 or n5574 or n5573 or n5572 or n5571 or n5570 or n5569
 or n5568 or n5567 or n5566 or n5565 or n5564 or n5563 or n5562 or n5561
 or n5560 or n5559 or n5558 or n5557 or n5556 or n5555 or n5554 or n5553
 or n5552 or n5551 or n5550 or n5549 or n5548 or n5547 or n5546 or n5545
 or n5544 or n5543 or n5542 or n5541 or n5540 or n5539 or n5538 or n5537
 or n5536 or n5535 or n5534 or n5533 or n5532 or n5531 or n5530 or n5529
 or n5528 or n5527 or n5526 or n5525 or n5524 or n5523 or n5522 or n5521
 or n5520 or n5519 or n5518 or n5517 or n5516 or n5515 or n5514 or n5513
 or n5507 or _zygsfis_get_config_data_rptr[4] or _zygsfis_get_config_data_rptr[3] or _zygsfis_get_config_data_rptr[2] or _zygsfis_get_config_data_rptr[1] or _zygsfis_get_config_data_rptr[0])
#0 begin
if (n5507)
_zygsfis_get_config_data_fifo[{n5512, n5511, n5510, n5509, n5508}] =
{n5584, n5583, n5582, n5581, n5580,
 n5579, n5578, n5577, n5576, n5575, n5574, n5573, n5572,
 n5571, n5570, n5569, n5568, n5567, n5566, n5565, n5564,
 n5563, n5562, n5561, n5560, n5559, n5558, n5557, n5556,
 n5555, n5554, n5553, n5552, n5551, n5550, n5549, n5548,
 n5547, n5546, n5545, n5544, n5543, n5542, n5541, n5540,
 n5539, n5538, n5537, n5536, n5535, n5534, n5533, n5532,
 n5531, n5530, n5529, n5528, n5527, n5526, n5525, n5524,
 n5523, n5522, n5521, n5520, n5519, n5518, n5517, n5516,
 n5515, n5514, n5513};
n5887 = _zygsfis_get_config_data_fifo[{_zygsfis_get_config_data_rptr[4], _zygsfis_get_config_data_rptr[3], _zygsfis_get_config_data_rptr[2], _zygsfis_get_config_data_rptr[1], _zygsfis_get_config_data_rptr[0]}];
end
`else

MPW32X72 _zygsfis_get_config_data_fifo ( .A4(n5512), .A3(n5511), .A2(n5510), .A1(n5509), .A0(n5508), .DI71(n5584),
 .DI70(n5583), .DI69(n5582), .DI68(n5581), .DI67(n5580), .DI66(n5579), .DI65(n5578), .DI64(n5577), .DI63(n5576),
 .DI62(n5575), .DI61(n5574), .DI60(n5573), .DI59(n5572), .DI58(n5571), .DI57(n5570), .DI56(n5569), .DI55(n5568),
 .DI54(n5567), .DI53(n5566), .DI52(n5565), .DI51(n5564), .DI50(n5563), .DI49(n5562), .DI48(n5561), .DI47(n5560),
 .DI46(n5559), .DI45(n5558), .DI44(n5557), .DI43(n5556), .DI42(n5555), .DI41(n5554), .DI40(n5553), .DI39(n5552),
 .DI38(n5551), .DI37(n5550), .DI36(n5549), .DI35(n5548), .DI34(n5547), .DI33(n5546), .DI32(n5545), .DI31(n5544),
 .DI30(n5543), .DI29(n5542), .DI28(n5541), .DI27(n5540), .DI26(n5539), .DI25(n5538), .DI24(n5537), .DI23(n5536),
 .DI22(n5535), .DI21(n5534), .DI20(n5533), .DI19(n5532), .DI18(n5531), .DI17(n5530), .DI16(n5529), .DI15(n5528),
 .DI14(n5527), .DI13(n5526), .DI12(n5525), .DI11(n5524), .DI10(n5523), .DI9(n5522), .DI8(n5521), .DI7(n5520),
 .DI6(n5519), .DI5(n5518), .DI4(n5517), .DI3(n5516), .DI2(n5515), .DI1(n5514), .DI0(n5513), .WE(n5507),
 .SYNC_IN(n1750), .SYNC_OUT(n5887));
// pragma CVASTRPROP INSTANCE "_zygsfis_get_config_data_fifo" HDL_MEMORY_DECL "1 71 0 0 31"
MPR32X72 U9783 ( .A4(_zygsfis_get_config_data_rptr[4]), .A3(_zygsfis_get_config_data_rptr[3]), .A2(_zygsfis_get_config_data_rptr[2]), .A1(_zygsfis_get_config_data_rptr[1]), .A0(_zygsfis_get_config_data_rptr[0]), .SYNC_IN(n5887),
 .DO71(n1051), .DO70(n1052), .DO69(n1053), .DO68(n1054), .DO67(n1055), .DO66(n1056), .DO65(n1057), .DO64(n1058),
 .DO63(n1059), .DO62(n1060), .DO61(n1061), .DO60(n1062), .DO59(n1063), .DO58(n1064), .DO57(n1065), .DO56(n1066),
 .DO55(n1067), .DO54(n1068), .DO53(n1069), .DO52(n1070), .DO51(n1071), .DO50(n1072), .DO49(n1073), .DO48(n1074),
 .DO47(n1075), .DO46(n1076), .DO45(n1077), .DO44(n1078), .DO43(n1079), .DO42(n1080), .DO41(n1081), .DO40(n1082),
 .DO39(n1083), .DO38(n1084), .DO37(n1085), .DO36(n1086), .DO35(n1087), .DO34(n1088), .DO33(n1089), .DO32(n1090),
 .DO31(n1091), .DO30(n1092), .DO29(n1093), .DO28(n1094), .DO27(n1095), .DO26(n1096), .DO25(n1097), .DO24(n1098),
 .DO23(n1099), .DO22(n1100), .DO21(n1101), .DO20(n1102), .DO19(n1103), .DO18(n1104), .DO17(n1105), .DO16(n1106),
 .DO15(n1107), .DO14(n1108), .DO13(n1109), .DO12(n1110), .DO11(n1111), .DO10(n1112), .DO9(n1113), .DO8(n1114),
 .DO7(n1115), .DO6(n1116), .DO5(n1117), .DO4(n1118), .DO3(n1119), .DO2(n1120), .DO1(n1121), .DO0(n1122),
 .SYNC_OUT( ));
`endif
`ifdef CBV

reg [135:0] _zygsfis_ib_service_data_fifo [0:31];
initial begin: U9784
  integer i;
  for (i=0; i<=31; i=i+1) _zygsfis_ib_service_data_fifo[i] =
`ifdef CBV_MEM_INIT1
  {136{1'b1}};
`else
  136'b0;
`endif
end
reg [135:0] n5888;
assign {n1493, n1494, n1495, n1496, n1497, n1498, n1499,
n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
n1628} = n5888; 
always @(n5593 or n5592 or n5591 or n5590 or n5589
 or n5729 or n5728 or n5727 or n5726 or n5725 or n5724 or n5723 or n5722
 or n5721 or n5720 or n5719 or n5718 or n5717 or n5716 or n5715 or n5714
 or n5713 or n5712 or n5711 or n5710 or n5709 or n5708 or n5707 or n5706
 or n5705 or n5704 or n5703 or n5702 or n5701 or n5700 or n5699 or n5698
 or n5697 or n5696 or n5695 or n5694 or n5693 or n5692 or n5691 or n5690
 or n5689 or n5688 or n5687 or n5686 or n5685 or n5684 or n5683 or n5682
 or n5681 or n5680 or n5679 or n5678 or n5677 or n5676 or n5675 or n5674
 or n5673 or n5672 or n5671 or n5670 or n5669 or n5668 or n5667 or n5666
 or n5665 or n5664 or n5663 or n5662 or n5661 or n5660 or n5659 or n5658
 or n5657 or n5656 or n5655 or n5654 or n5653 or n5652 or n5651 or n5650
 or n5649 or n5648 or n5647 or n5646 or n5645 or n5644 or n5643 or n5642
 or n5641 or n5640 or n5639 or n5638 or n5637 or n5636 or n5635 or n5634
 or n5633 or n5632 or n5631 or n5630 or n5629 or n5628 or n5627 or n5626
 or n5625 or n5624 or n5623 or n5622 or n5621 or n5620 or n5619 or n5618
 or n5617 or n5616 or n5615 or n5614 or n5613 or n5612 or n5611 or n5610
 or n5609 or n5608 or n5607 or n5606 or n5605 or n5604 or n5603 or n5602
 or n5601 or n5600 or n5599 or n5598 or n5597 or n5596 or n5595 or n5594
 or n5588 or _zygsfis_ib_service_data_rptr[4] or _zygsfis_ib_service_data_rptr[3] or _zygsfis_ib_service_data_rptr[2] or _zygsfis_ib_service_data_rptr[1] or _zygsfis_ib_service_data_rptr[0])
#0 begin
if (n5588)
_zygsfis_ib_service_data_fifo[{n5593, n5592, n5591, n5590, n5589}] =
{n5729, n5728, n5727, n5726, n5725,
 n5724, n5723, n5722, n5721, n5720, n5719, n5718, n5717,
 n5716, n5715, n5714, n5713, n5712, n5711, n5710, n5709,
 n5708, n5707, n5706, n5705, n5704, n5703, n5702, n5701,
 n5700, n5699, n5698, n5697, n5696, n5695, n5694, n5693,
 n5692, n5691, n5690, n5689, n5688, n5687, n5686, n5685,
 n5684, n5683, n5682, n5681, n5680, n5679, n5678, n5677,
 n5676, n5675, n5674, n5673, n5672, n5671, n5670, n5669,
 n5668, n5667, n5666, n5665, n5664, n5663, n5662, n5661,
 n5660, n5659, n5658, n5657, n5656, n5655, n5654, n5653,
 n5652, n5651, n5650, n5649, n5648, n5647, n5646, n5645,
 n5644, n5643, n5642, n5641, n5640, n5639, n5638, n5637,
 n5636, n5635, n5634, n5633, n5632, n5631, n5630, n5629,
 n5628, n5627, n5626, n5625, n5624, n5623, n5622, n5621,
 n5620, n5619, n5618, n5617, n5616, n5615, n5614, n5613,
 n5612, n5611, n5610, n5609, n5608, n5607, n5606, n5605,
 n5604, n5603, n5602, n5601, n5600, n5599, n5598, n5597,
 n5596, n5595, n5594};
n5888 = _zygsfis_ib_service_data_fifo[{_zygsfis_ib_service_data_rptr[4], _zygsfis_ib_service_data_rptr[3], _zygsfis_ib_service_data_rptr[2], _zygsfis_ib_service_data_rptr[1], _zygsfis_ib_service_data_rptr[0]}];
end
`else

MPW32X136 _zygsfis_ib_service_data_fifo ( .A4(n5593), .A3(n5592), .A2(n5591), .A1(n5590), .A0(n5589), .DI135(n5729),
 .DI134(n5728), .DI133(n5727), .DI132(n5726), .DI131(n5725), .DI130(n5724), .DI129(n5723), .DI128(n5722), .DI127(n5721),
 .DI126(n5720), .DI125(n5719), .DI124(n5718), .DI123(n5717), .DI122(n5716), .DI121(n5715), .DI120(n5714), .DI119(n5713),
 .DI118(n5712), .DI117(n5711), .DI116(n5710), .DI115(n5709), .DI114(n5708), .DI113(n5707), .DI112(n5706), .DI111(n5705),
 .DI110(n5704), .DI109(n5703), .DI108(n5702), .DI107(n5701), .DI106(n5700), .DI105(n5699), .DI104(n5698), .DI103(n5697),
 .DI102(n5696), .DI101(n5695), .DI100(n5694), .DI99(n5693), .DI98(n5692), .DI97(n5691), .DI96(n5690), .DI95(n5689),
 .DI94(n5688), .DI93(n5687), .DI92(n5686), .DI91(n5685), .DI90(n5684), .DI89(n5683), .DI88(n5682), .DI87(n5681),
 .DI86(n5680), .DI85(n5679), .DI84(n5678), .DI83(n5677), .DI82(n5676), .DI81(n5675), .DI80(n5674), .DI79(n5673),
 .DI78(n5672), .DI77(n5671), .DI76(n5670), .DI75(n5669), .DI74(n5668), .DI73(n5667), .DI72(n5666), .DI71(n5665),
 .DI70(n5664), .DI69(n5663), .DI68(n5662), .DI67(n5661), .DI66(n5660), .DI65(n5659), .DI64(n5658), .DI63(n5657),
 .DI62(n5656), .DI61(n5655), .DI60(n5654), .DI59(n5653), .DI58(n5652), .DI57(n5651), .DI56(n5650), .DI55(n5649),
 .DI54(n5648), .DI53(n5647), .DI52(n5646), .DI51(n5645), .DI50(n5644), .DI49(n5643), .DI48(n5642), .DI47(n5641),
 .DI46(n5640), .DI45(n5639), .DI44(n5638), .DI43(n5637), .DI42(n5636), .DI41(n5635), .DI40(n5634), .DI39(n5633),
 .DI38(n5632), .DI37(n5631), .DI36(n5630), .DI35(n5629), .DI34(n5628), .DI33(n5627), .DI32(n5626), .DI31(n5625),
 .DI30(n5624), .DI29(n5623), .DI28(n5622), .DI27(n5621), .DI26(n5620), .DI25(n5619), .DI24(n5618), .DI23(n5617),
 .DI22(n5616), .DI21(n5615), .DI20(n5614), .DI19(n5613), .DI18(n5612), .DI17(n5611), .DI16(n5610), .DI15(n5609),
 .DI14(n5608), .DI13(n5607), .DI12(n5606), .DI11(n5605), .DI10(n5604), .DI9(n5603), .DI8(n5602), .DI7(n5601),
 .DI6(n5600), .DI5(n5599), .DI4(n5598), .DI3(n5597), .DI2(n5596), .DI1(n5595), .DI0(n5594), .WE(n5588),
 .SYNC_IN(n1750), .SYNC_OUT(n5888));
// pragma CVASTRPROP INSTANCE "_zygsfis_ib_service_data_fifo" HDL_MEMORY_DECL "1 135 0 0 31"
MPR32X136 U9785 ( .A4(_zygsfis_ib_service_data_rptr[4]), .A3(_zygsfis_ib_service_data_rptr[3]), .A2(_zygsfis_ib_service_data_rptr[2]), .A1(_zygsfis_ib_service_data_rptr[1]), .A0(_zygsfis_ib_service_data_rptr[0]), .SYNC_IN(n5888),
 .DO135(n1493), .DO134(n1494), .DO133(n1495), .DO132(n1496), .DO131(n1497), .DO130(n1498), .DO129(n1499), .DO128(n1500),
 .DO127(n1501), .DO126(n1502), .DO125(n1503), .DO124(n1504), .DO123(n1505), .DO122(n1506), .DO121(n1507), .DO120(n1508),
 .DO119(n1509), .DO118(n1510), .DO117(n1511), .DO116(n1512), .DO115(n1513), .DO114(n1514), .DO113(n1515), .DO112(n1516),
 .DO111(n1517), .DO110(n1518), .DO109(n1519), .DO108(n1520), .DO107(n1521), .DO106(n1522), .DO105(n1523), .DO104(n1524),
 .DO103(n1525), .DO102(n1526), .DO101(n1527), .DO100(n1528), .DO99(n1529), .DO98(n1530), .DO97(n1531), .DO96(n1532),
 .DO95(n1533), .DO94(n1534), .DO93(n1535), .DO92(n1536), .DO91(n1537), .DO90(n1538), .DO89(n1539), .DO88(n1540),
 .DO87(n1541), .DO86(n1542), .DO85(n1543), .DO84(n1544), .DO83(n1545), .DO82(n1546), .DO81(n1547), .DO80(n1548),
 .DO79(n1549), .DO78(n1550), .DO77(n1551), .DO76(n1552), .DO75(n1553), .DO74(n1554), .DO73(n1555), .DO72(n1556),
 .DO71(n1557), .DO70(n1558), .DO69(n1559), .DO68(n1560), .DO67(n1561), .DO66(n1562), .DO65(n1563), .DO64(n1564),
 .DO63(n1565), .DO62(n1566), .DO61(n1567), .DO60(n1568), .DO59(n1569), .DO58(n1570), .DO57(n1571), .DO56(n1572),
 .DO55(n1573), .DO54(n1574), .DO53(n1575), .DO52(n1576), .DO51(n1577), .DO50(n1578), .DO49(n1579), .DO48(n1580),
 .DO47(n1581), .DO46(n1582), .DO45(n1583), .DO44(n1584), .DO43(n1585), .DO42(n1586), .DO41(n1587), .DO40(n1588),
 .DO39(n1589), .DO38(n1590), .DO37(n1591), .DO36(n1592), .DO35(n1593), .DO34(n1594), .DO33(n1595), .DO32(n1596),
 .DO31(n1597), .DO30(n1598), .DO29(n1599), .DO28(n1600), .DO27(n1601), .DO26(n1602), .DO25(n1603), .DO24(n1604),
 .DO23(n1605), .DO22(n1606), .DO21(n1607), .DO20(n1608), .DO19(n1609), .DO18(n1610), .DO17(n1611), .DO16(n1612),
 .DO15(n1613), .DO14(n1614), .DO13(n1615), .DO12(n1616), .DO11(n1617), .DO10(n1618), .DO9(n1619), .DO8(n1620),
 .DO7(n1621), .DO6(n1622), .DO5(n1623), .DO4(n1624), .DO3(n1625), .DO2(n1626), .DO1(n1627), .DO0(n1628),
 .SYNC_OUT( ));
`endif
`ifdef CBV

reg [135:0] _zygsfis_ob_service_data_fifo [0:31];
initial begin: U9786
  integer i;
  for (i=0; i<=31; i=i+1) _zygsfis_ob_service_data_fifo[i] =
`ifdef CBV_MEM_INIT1
  {136{1'b1}};
`else
  136'b0;
`endif
end
reg [135:0] n5889;
assign {n3398, n3399, n3400, n3401, n3402, n3403, n3404,
n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
n3533} = n5889; 
always @(n5738 or n5737 or n5736 or n5735 or n5734
 or n5874 or n5873 or n5872 or n5871 or n5870 or n5869 or n5868 or n5867
 or n5866 or n5865 or n5864 or n5863 or n5862 or n5861 or n5860 or n5859
 or n5858 or n5857 or n5856 or n5855 or n5854 or n5853 or n5852 or n5851
 or n5850 or n5849 or n5848 or n5847 or n5846 or n5845 or n5844 or n5843
 or n5842 or n5841 or n5840 or n5839 or n5838 or n5837 or n5836 or n5835
 or n5834 or n5833 or n5832 or n5831 or n5830 or n5829 or n5828 or n5827
 or n5826 or n5825 or n5824 or n5823 or n5822 or n5821 or n5820 or n5819
 or n5818 or n5817 or n5816 or n5815 or n5814 or n5813 or n5812 or n5811
 or n5810 or n5809 or n5808 or n5807 or n5806 or n5805 or n5804 or n5803
 or n5802 or n5801 or n5800 or n5799 or n5798 or n5797 or n5796 or n5795
 or n5794 or n5793 or n5792 or n5791 or n5790 or n5789 or n5788 or n5787
 or n5786 or n5785 or n5784 or n5783 or n5782 or n5781 or n5780 or n5779
 or n5778 or n5777 or n5776 or n5775 or n5774 or n5773 or n5772 or n5771
 or n5770 or n5769 or n5768 or n5767 or n5766 or n5765 or n5764 or n5763
 or n5762 or n5761 or n5760 or n5759 or n5758 or n5757 or n5756 or n5755
 or n5754 or n5753 or n5752 or n5751 or n5750 or n5749 or n5748 or n5747
 or n5746 or n5745 or n5744 or n5743 or n5742 or n5741 or n5740 or n5739
 or n5733 or _zygsfis_ob_service_data_rptr[4] or _zygsfis_ob_service_data_rptr[3] or _zygsfis_ob_service_data_rptr[2] or _zygsfis_ob_service_data_rptr[1] or _zygsfis_ob_service_data_rptr[0])
#0 begin
if (n5733)
_zygsfis_ob_service_data_fifo[{n5738, n5737, n5736, n5735, n5734}] =
{n5874, n5873, n5872, n5871, n5870,
 n5869, n5868, n5867, n5866, n5865, n5864, n5863, n5862,
 n5861, n5860, n5859, n5858, n5857, n5856, n5855, n5854,
 n5853, n5852, n5851, n5850, n5849, n5848, n5847, n5846,
 n5845, n5844, n5843, n5842, n5841, n5840, n5839, n5838,
 n5837, n5836, n5835, n5834, n5833, n5832, n5831, n5830,
 n5829, n5828, n5827, n5826, n5825, n5824, n5823, n5822,
 n5821, n5820, n5819, n5818, n5817, n5816, n5815, n5814,
 n5813, n5812, n5811, n5810, n5809, n5808, n5807, n5806,
 n5805, n5804, n5803, n5802, n5801, n5800, n5799, n5798,
 n5797, n5796, n5795, n5794, n5793, n5792, n5791, n5790,
 n5789, n5788, n5787, n5786, n5785, n5784, n5783, n5782,
 n5781, n5780, n5779, n5778, n5777, n5776, n5775, n5774,
 n5773, n5772, n5771, n5770, n5769, n5768, n5767, n5766,
 n5765, n5764, n5763, n5762, n5761, n5760, n5759, n5758,
 n5757, n5756, n5755, n5754, n5753, n5752, n5751, n5750,
 n5749, n5748, n5747, n5746, n5745, n5744, n5743, n5742,
 n5741, n5740, n5739};
n5889 = _zygsfis_ob_service_data_fifo[{_zygsfis_ob_service_data_rptr[4], _zygsfis_ob_service_data_rptr[3], _zygsfis_ob_service_data_rptr[2], _zygsfis_ob_service_data_rptr[1], _zygsfis_ob_service_data_rptr[0]}];
end
`else

MPW32X136 _zygsfis_ob_service_data_fifo ( .A4(n5738), .A3(n5737), .A2(n5736), .A1(n5735), .A0(n5734), .DI135(n5874),
 .DI134(n5873), .DI133(n5872), .DI132(n5871), .DI131(n5870), .DI130(n5869), .DI129(n5868), .DI128(n5867), .DI127(n5866),
 .DI126(n5865), .DI125(n5864), .DI124(n5863), .DI123(n5862), .DI122(n5861), .DI121(n5860), .DI120(n5859), .DI119(n5858),
 .DI118(n5857), .DI117(n5856), .DI116(n5855), .DI115(n5854), .DI114(n5853), .DI113(n5852), .DI112(n5851), .DI111(n5850),
 .DI110(n5849), .DI109(n5848), .DI108(n5847), .DI107(n5846), .DI106(n5845), .DI105(n5844), .DI104(n5843), .DI103(n5842),
 .DI102(n5841), .DI101(n5840), .DI100(n5839), .DI99(n5838), .DI98(n5837), .DI97(n5836), .DI96(n5835), .DI95(n5834),
 .DI94(n5833), .DI93(n5832), .DI92(n5831), .DI91(n5830), .DI90(n5829), .DI89(n5828), .DI88(n5827), .DI87(n5826),
 .DI86(n5825), .DI85(n5824), .DI84(n5823), .DI83(n5822), .DI82(n5821), .DI81(n5820), .DI80(n5819), .DI79(n5818),
 .DI78(n5817), .DI77(n5816), .DI76(n5815), .DI75(n5814), .DI74(n5813), .DI73(n5812), .DI72(n5811), .DI71(n5810),
 .DI70(n5809), .DI69(n5808), .DI68(n5807), .DI67(n5806), .DI66(n5805), .DI65(n5804), .DI64(n5803), .DI63(n5802),
 .DI62(n5801), .DI61(n5800), .DI60(n5799), .DI59(n5798), .DI58(n5797), .DI57(n5796), .DI56(n5795), .DI55(n5794),
 .DI54(n5793), .DI53(n5792), .DI52(n5791), .DI51(n5790), .DI50(n5789), .DI49(n5788), .DI48(n5787), .DI47(n5786),
 .DI46(n5785), .DI45(n5784), .DI44(n5783), .DI43(n5782), .DI42(n5781), .DI41(n5780), .DI40(n5779), .DI39(n5778),
 .DI38(n5777), .DI37(n5776), .DI36(n5775), .DI35(n5774), .DI34(n5773), .DI33(n5772), .DI32(n5771), .DI31(n5770),
 .DI30(n5769), .DI29(n5768), .DI28(n5767), .DI27(n5766), .DI26(n5765), .DI25(n5764), .DI24(n5763), .DI23(n5762),
 .DI22(n5761), .DI21(n5760), .DI20(n5759), .DI19(n5758), .DI18(n5757), .DI17(n5756), .DI16(n5755), .DI15(n5754),
 .DI14(n5753), .DI13(n5752), .DI12(n5751), .DI11(n5750), .DI10(n5749), .DI9(n5748), .DI8(n5747), .DI7(n5746),
 .DI6(n5745), .DI5(n5744), .DI4(n5743), .DI3(n5742), .DI2(n5741), .DI1(n5740), .DI0(n5739), .WE(n5733),
 .SYNC_IN(n1750), .SYNC_OUT(n5889));
// pragma CVASTRPROP INSTANCE "_zygsfis_ob_service_data_fifo" HDL_MEMORY_DECL "1 135 0 0 31"
MPR32X136 U9787 ( .A4(_zygsfis_ob_service_data_rptr[4]), .A3(_zygsfis_ob_service_data_rptr[3]), .A2(_zygsfis_ob_service_data_rptr[2]), .A1(_zygsfis_ob_service_data_rptr[1]), .A0(_zygsfis_ob_service_data_rptr[0]), .SYNC_IN(n5889),
 .DO135(n3398), .DO134(n3399), .DO133(n3400), .DO132(n3401), .DO131(n3402), .DO130(n3403), .DO129(n3404), .DO128(n3405),
 .DO127(n3406), .DO126(n3407), .DO125(n3408), .DO124(n3409), .DO123(n3410), .DO122(n3411), .DO121(n3412), .DO120(n3413),
 .DO119(n3414), .DO118(n3415), .DO117(n3416), .DO116(n3417), .DO115(n3418), .DO114(n3419), .DO113(n3420), .DO112(n3421),
 .DO111(n3422), .DO110(n3423), .DO109(n3424), .DO108(n3425), .DO107(n3426), .DO106(n3427), .DO105(n3428), .DO104(n3429),
 .DO103(n3430), .DO102(n3431), .DO101(n3432), .DO100(n3433), .DO99(n3434), .DO98(n3435), .DO97(n3436), .DO96(n3437),
 .DO95(n3438), .DO94(n3439), .DO93(n3440), .DO92(n3441), .DO91(n3442), .DO90(n3443), .DO89(n3444), .DO88(n3445),
 .DO87(n3446), .DO86(n3447), .DO85(n3448), .DO84(n3449), .DO83(n3450), .DO82(n3451), .DO81(n3452), .DO80(n3453),
 .DO79(n3454), .DO78(n3455), .DO77(n3456), .DO76(n3457), .DO75(n3458), .DO74(n3459), .DO73(n3460), .DO72(n3461),
 .DO71(n3462), .DO70(n3463), .DO69(n3464), .DO68(n3465), .DO67(n3466), .DO66(n3467), .DO65(n3468), .DO64(n3469),
 .DO63(n3470), .DO62(n3471), .DO61(n3472), .DO60(n3473), .DO59(n3474), .DO58(n3475), .DO57(n3476), .DO56(n3477),
 .DO55(n3478), .DO54(n3479), .DO53(n3480), .DO52(n3481), .DO51(n3482), .DO50(n3483), .DO49(n3484), .DO48(n3485),
 .DO47(n3486), .DO46(n3487), .DO45(n3488), .DO44(n3489), .DO43(n3490), .DO42(n3491), .DO41(n3492), .DO40(n3493),
 .DO39(n3494), .DO38(n3495), .DO37(n3496), .DO36(n3497), .DO35(n3498), .DO34(n3499), .DO33(n3500), .DO32(n3501),
 .DO31(n3502), .DO30(n3503), .DO29(n3504), .DO28(n3505), .DO27(n3506), .DO26(n3507), .DO25(n3508), .DO24(n3509),
 .DO23(n3510), .DO22(n3511), .DO21(n3512), .DO20(n3513), .DO19(n3514), .DO18(n3515), .DO17(n3516), .DO16(n3517),
 .DO15(n3518), .DO14(n3519), .DO13(n3520), .DO12(n3521), .DO11(n3522), .DO10(n3523), .DO9(n3524), .DO8(n3525),
 .DO7(n3526), .DO6(n3527), .DO5(n3528), .DO4(n3529), .DO3(n3530), .DO2(n3531), .DO1(n3532), .DO0(n3533),
 .SYNC_OUT( ));
`endif
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "_zygsfis_get_config_data_fifo 1 71 0 0 31"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m2 "_zygsfis_ib_service_data_fifo 1 135 0 0 31"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m3 "_zygsfis_ob_service_data_fifo 1 135 0 0 31"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "3"
// pragma CVASTRPROP MODULE HDLICE PROP_RANOFF TRUE
endmodule
`ifdef CBV
`else
`ifdef MPW32X136_MPR32X136
`else
module MPW32X136( A4, A3, A2, A1, A0, DI135, DI134,
 DI133, DI132, DI131, DI130, DI129, DI128, DI127, DI126,
 DI125, DI124, DI123, DI122, DI121, DI120, DI119, DI118,
 DI117, DI116, DI115, DI114, DI113, DI112, DI111, DI110,
 DI109, DI108, DI107, DI106, DI105, DI104, DI103, DI102,
 DI101, DI100, DI99, DI98, DI97, DI96, DI95, DI94,
 DI93, DI92, DI91, DI90, DI89, DI88, DI87, DI86,
 DI85, DI84, DI83, DI82, DI81, DI80, DI79, DI78,
 DI77, DI76, DI75, DI74, DI73, DI72, DI71, DI70,
 DI69, DI68, DI67, DI66, DI65, DI64, DI63, DI62,
 DI61, DI60, DI59, DI58, DI57, DI56, DI55, DI54,
 DI53, DI52, DI51, DI50, DI49, DI48, DI47, DI46,
 DI45, DI44, DI43, DI42, DI41, DI40, DI39, DI38,
 DI37, DI36, DI35, DI34, DI33, DI32, DI31, DI30,
 DI29, DI28, DI27, DI26, DI25, DI24, DI23, DI22,
 DI21, DI20, DI19, DI18, DI17, DI16, DI15, DI14,
 DI13, DI12, DI11, DI10, DI9, DI8, DI7, DI6,
 DI5, DI4, DI3, DI2, DI1, DI0, WE, SYNC_IN,
 SYNC_OUT);
input  A4, A3, A2, A1, A0, DI135, DI134, DI133,
 DI132, DI131, DI130, DI129, DI128, DI127, DI126, DI125, DI124, DI123,
 DI122, DI121, DI120, DI119, DI118, DI117, DI116, DI115, DI114, DI113,
 DI112, DI111, DI110, DI109, DI108, DI107, DI106, DI105, DI104, DI103,
 DI102, DI101, DI100, DI99, DI98, DI97, DI96, DI95, DI94, DI93,
 DI92, DI91, DI90, DI89, DI88, DI87, DI86, DI85, DI84, DI83,
 DI82, DI81, DI80, DI79, DI78, DI77, DI76, DI75, DI74, DI73,
 DI72, DI71, DI70, DI69, DI68, DI67, DI66, DI65, DI64, DI63,
 DI62, DI61, DI60, DI59, DI58, DI57, DI56, DI55, DI54, DI53,
 DI52, DI51, DI50, DI49, DI48, DI47, DI46, DI45, DI44, DI43,
 DI42, DI41, DI40, DI39, DI38, DI37, DI36, DI35, DI34, DI33,
 DI32, DI31, DI30, DI29, DI28, DI27, DI26, DI25, DI24, DI23,
 DI22, DI21, DI20, DI19, DI18, DI17, DI16, DI15, DI14, DI13,
 DI12, DI11, DI10, DI9, DI8, DI7, DI6, DI5, DI4, DI3,
 DI2, DI1, DI0, WE, SYNC_IN;
output  SYNC_OUT;
endmodule
`ifdef _MPR32X136_
`else
module MPR32X136( A4, A3, A2, A1, A0, SYNC_IN, DO135,
 DO134, DO133, DO132, DO131, DO130, DO129, DO128, DO127,
 DO126, DO125, DO124, DO123, DO122, DO121, DO120, DO119,
 DO118, DO117, DO116, DO115, DO114, DO113, DO112, DO111,
 DO110, DO109, DO108, DO107, DO106, DO105, DO104, DO103,
 DO102, DO101, DO100, DO99, DO98, DO97, DO96, DO95,
 DO94, DO93, DO92, DO91, DO90, DO89, DO88, DO87,
 DO86, DO85, DO84, DO83, DO82, DO81, DO80, DO79,
 DO78, DO77, DO76, DO75, DO74, DO73, DO72, DO71,
 DO70, DO69, DO68, DO67, DO66, DO65, DO64, DO63,
 DO62, DO61, DO60, DO59, DO58, DO57, DO56, DO55,
 DO54, DO53, DO52, DO51, DO50, DO49, DO48, DO47,
 DO46, DO45, DO44, DO43, DO42, DO41, DO40, DO39,
 DO38, DO37, DO36, DO35, DO34, DO33, DO32, DO31,
 DO30, DO29, DO28, DO27, DO26, DO25, DO24, DO23,
 DO22, DO21, DO20, DO19, DO18, DO17, DO16, DO15,
 DO14, DO13, DO12, DO11, DO10, DO9, DO8, DO7,
 DO6, DO5, DO4, DO3, DO2, DO1, DO0, SYNC_OUT);
input  A4, A3, A2, A1, A0, SYNC_IN;
output  DO135, DO134, DO133, DO132, DO131, DO130, DO129, DO128,
 DO127, DO126, DO125, DO124, DO123, DO122, DO121, DO120, DO119, DO118,
 DO117, DO116, DO115, DO114, DO113, DO112, DO111, DO110, DO109, DO108,
 DO107, DO106, DO105, DO104, DO103, DO102, DO101, DO100, DO99, DO98,
 DO97, DO96, DO95, DO94, DO93, DO92, DO91, DO90, DO89, DO88,
 DO87, DO86, DO85, DO84, DO83, DO82, DO81, DO80, DO79, DO78,
 DO77, DO76, DO75, DO74, DO73, DO72, DO71, DO70, DO69, DO68,
 DO67, DO66, DO65, DO64, DO63, DO62, DO61, DO60, DO59, DO58,
 DO57, DO56, DO55, DO54, DO53, DO52, DO51, DO50, DO49, DO48,
 DO47, DO46, DO45, DO44, DO43, DO42, DO41, DO40, DO39, DO38,
 DO37, DO36, DO35, DO34, DO33, DO32, DO31, DO30, DO29, DO28,
 DO27, DO26, DO25, DO24, DO23, DO22, DO21, DO20, DO19, DO18,
 DO17, DO16, DO15, DO14, DO13, DO12, DO11, DO10, DO9, DO8,
 DO7, DO6, DO5, DO4, DO3, DO2, DO1, DO0, SYNC_OUT;
endmodule
`define _MPR32X136_
`endif
`define MPW32X136_MPR32X136
`endif
`ifdef MPW32X72_MPR32X72
`else
module MPW32X72( A4, A3, A2, A1, A0, DI71, DI70,
 DI69, DI68, DI67, DI66, DI65, DI64, DI63, DI62,
 DI61, DI60, DI59, DI58, DI57, DI56, DI55, DI54,
 DI53, DI52, DI51, DI50, DI49, DI48, DI47, DI46,
 DI45, DI44, DI43, DI42, DI41, DI40, DI39, DI38,
 DI37, DI36, DI35, DI34, DI33, DI32, DI31, DI30,
 DI29, DI28, DI27, DI26, DI25, DI24, DI23, DI22,
 DI21, DI20, DI19, DI18, DI17, DI16, DI15, DI14,
 DI13, DI12, DI11, DI10, DI9, DI8, DI7, DI6,
 DI5, DI4, DI3, DI2, DI1, DI0, WE, SYNC_IN,
 SYNC_OUT);
input  A4, A3, A2, A1, A0, DI71, DI70, DI69,
 DI68, DI67, DI66, DI65, DI64, DI63, DI62, DI61, DI60, DI59,
 DI58, DI57, DI56, DI55, DI54, DI53, DI52, DI51, DI50, DI49,
 DI48, DI47, DI46, DI45, DI44, DI43, DI42, DI41, DI40, DI39,
 DI38, DI37, DI36, DI35, DI34, DI33, DI32, DI31, DI30, DI29,
 DI28, DI27, DI26, DI25, DI24, DI23, DI22, DI21, DI20, DI19,
 DI18, DI17, DI16, DI15, DI14, DI13, DI12, DI11, DI10, DI9,
 DI8, DI7, DI6, DI5, DI4, DI3, DI2, DI1, DI0, WE,
 SYNC_IN;
output  SYNC_OUT;
endmodule
`ifdef _MPR32X72_
`else
module MPR32X72( A4, A3, A2, A1, A0, SYNC_IN, DO71,
 DO70, DO69, DO68, DO67, DO66, DO65, DO64, DO63,
 DO62, DO61, DO60, DO59, DO58, DO57, DO56, DO55,
 DO54, DO53, DO52, DO51, DO50, DO49, DO48, DO47,
 DO46, DO45, DO44, DO43, DO42, DO41, DO40, DO39,
 DO38, DO37, DO36, DO35, DO34, DO33, DO32, DO31,
 DO30, DO29, DO28, DO27, DO26, DO25, DO24, DO23,
 DO22, DO21, DO20, DO19, DO18, DO17, DO16, DO15,
 DO14, DO13, DO12, DO11, DO10, DO9, DO8, DO7,
 DO6, DO5, DO4, DO3, DO2, DO1, DO0, SYNC_OUT);
input  A4, A3, A2, A1, A0, SYNC_IN;
output  DO71, DO70, DO69, DO68, DO67, DO66, DO65, DO64,
 DO63, DO62, DO61, DO60, DO59, DO58, DO57, DO56, DO55, DO54,
 DO53, DO52, DO51, DO50, DO49, DO48, DO47, DO46, DO45, DO44,
 DO43, DO42, DO41, DO40, DO39, DO38, DO37, DO36, DO35, DO34,
 DO33, DO32, DO31, DO30, DO29, DO28, DO27, DO26, DO25, DO24,
 DO23, DO22, DO21, DO20, DO19, DO18, DO17, DO16, DO15, DO14,
 DO13, DO12, DO11, DO10, DO9, DO8, DO7, DO6, DO5, DO4,
 DO3, DO2, DO1, DO0, SYNC_OUT;
endmodule
`define _MPR32X72_
`endif
`define MPW32X72_MPR32X72
`endif
`endif
