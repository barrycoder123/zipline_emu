architecture module of ixc_sfifo_bind_1_2 is

begin
end module;
