library ieee, quickturn ;
use ieee.std_logic_1164.all ;
use quickturn.verilog.all ;
entity cr_kme_regs is
  generic (
    IDLE : std_logic_vector := std_logic_vector'("000");
    WR_PREP : std_logic_vector := std_logic_vector'("001");
    WR_REG : std_logic_vector := std_logic_vector'("011");
    DUMMY0 : std_logic_vector := std_logic_vector'("100");
    RD_PREP : std_logic_vector := std_logic_vector'("101");
    RD_REG : std_logic_vector := std_logic_vector'("111")
  ) ;
  port (
    clk : in std_logic ;
    i_reset_ : in std_logic ;
    i_sw_init : in std_logic ;
    i_addr : in std_logic_vector(10 downto 0) ;
    i_wr_strb : in std_logic ;
    i_wr_data : in std_logic_vector(31 downto 0) ;
    i_rd_strb : in std_logic ;
    o_rd_data : out std_logic_vector(31 downto 0) ;
    o_ack : out std_logic ;
    o_err_ack : out std_logic ;
    o_spare_config : out std_logic_vector(31 downto 0) ;
    o_cceip0_out_ia_wdata_part0 : out std_logic_vector(31 downto 0) ;
    o_cceip0_out_ia_wdata_part1 : out std_logic_vector(31 downto 0) ;
    o_cceip0_out_ia_wdata_part2 : out std_logic_vector(31 downto 0) ;
    o_cceip0_out_ia_config : out std_logic_vector(12 downto 0) ;
    o_cceip0_out_im_config : out std_logic_vector(11 downto 0) ;
    o_cceip0_out_im_read_done : out std_logic_vector(1 downto 0) ;
    o_cceip1_out_ia_wdata_part0 : out std_logic_vector(31 downto 0) ;
    o_cceip1_out_ia_wdata_part1 : out std_logic_vector(31 downto 0) ;
    o_cceip1_out_ia_wdata_part2 : out std_logic_vector(31 downto 0) ;
    o_cceip1_out_ia_config : out std_logic_vector(12 downto 0) ;
    o_cceip1_out_im_config : out std_logic_vector(11 downto 0) ;
    o_cceip1_out_im_read_done : out std_logic_vector(1 downto 0) ;
    o_cceip2_out_ia_wdata_part0 : out std_logic_vector(31 downto 0) ;
    o_cceip2_out_ia_wdata_part1 : out std_logic_vector(31 downto 0) ;
    o_cceip2_out_ia_wdata_part2 : out std_logic_vector(31 downto 0) ;
    o_cceip2_out_ia_config : out std_logic_vector(12 downto 0) ;
    o_cceip2_out_im_config : out std_logic_vector(11 downto 0) ;
    o_cceip2_out_im_read_done : out std_logic_vector(1 downto 0) ;
    o_cceip3_out_ia_wdata_part0 : out std_logic_vector(31 downto 0) ;
    o_cceip3_out_ia_wdata_part1 : out std_logic_vector(31 downto 0) ;
    o_cceip3_out_ia_wdata_part2 : out std_logic_vector(31 downto 0) ;
    o_cceip3_out_ia_config : out std_logic_vector(12 downto 0) ;
    o_cceip3_out_im_config : out std_logic_vector(11 downto 0) ;
    o_cceip3_out_im_read_done : out std_logic_vector(1 downto 0) ;
    o_cddip0_out_ia_wdata_part0 : out std_logic_vector(31 downto 0) ;
    o_cddip0_out_ia_wdata_part1 : out std_logic_vector(31 downto 0) ;
    o_cddip0_out_ia_wdata_part2 : out std_logic_vector(31 downto 0) ;
    o_cddip0_out_ia_config : out std_logic_vector(12 downto 0) ;
    o_cddip0_out_im_config : out std_logic_vector(11 downto 0) ;
    o_cddip0_out_im_read_done : out std_logic_vector(1 downto 0) ;
    o_cddip1_out_ia_wdata_part0 : out std_logic_vector(31 downto 0) ;
    o_cddip1_out_ia_wdata_part1 : out std_logic_vector(31 downto 0) ;
    o_cddip1_out_ia_wdata_part2 : out std_logic_vector(31 downto 0) ;
    o_cddip1_out_ia_config : out std_logic_vector(12 downto 0) ;
    o_cddip1_out_im_config : out std_logic_vector(11 downto 0) ;
    o_cddip1_out_im_read_done : out std_logic_vector(1 downto 0) ;
    o_cddip2_out_ia_wdata_part0 : out std_logic_vector(31 downto 0) ;
    o_cddip2_out_ia_wdata_part1 : out std_logic_vector(31 downto 0) ;
    o_cddip2_out_ia_wdata_part2 : out std_logic_vector(31 downto 0) ;
    o_cddip2_out_ia_config : out std_logic_vector(12 downto 0) ;
    o_cddip2_out_im_config : out std_logic_vector(11 downto 0) ;
    o_cddip2_out_im_read_done : out std_logic_vector(1 downto 0) ;
    o_cddip3_out_ia_wdata_part0 : out std_logic_vector(31 downto 0) ;
    o_cddip3_out_ia_wdata_part1 : out std_logic_vector(31 downto 0) ;
    o_cddip3_out_ia_wdata_part2 : out std_logic_vector(31 downto 0) ;
    o_cddip3_out_ia_config : out std_logic_vector(12 downto 0) ;
    o_cddip3_out_im_config : out std_logic_vector(11 downto 0) ;
    o_cddip3_out_im_read_done : out std_logic_vector(1 downto 0) ;
    o_ckv_ia_wdata_part0 : out std_logic_vector(31 downto 0) ;
    o_ckv_ia_wdata_part1 : out std_logic_vector(31 downto 0) ;
    o_ckv_ia_config : out std_logic_vector(18 downto 0) ;
    o_kim_ia_wdata_part0 : out std_logic_vector(20 downto 0) ;
    o_kim_ia_wdata_part1 : out std_logic_vector(16 downto 0) ;
    o_kim_ia_config : out std_logic_vector(17 downto 0) ;
    o_label0_config : out std_logic_vector(15 downto 0) ;
    o_label0_data7 : out std_logic_vector(31 downto 0) ;
    o_label0_data6 : out std_logic_vector(31 downto 0) ;
    o_label0_data5 : out std_logic_vector(31 downto 0) ;
    o_label0_data4 : out std_logic_vector(31 downto 0) ;
    o_label0_data3 : out std_logic_vector(31 downto 0) ;
    o_label0_data2 : out std_logic_vector(31 downto 0) ;
    o_label0_data1 : out std_logic_vector(31 downto 0) ;
    o_label0_data0 : out std_logic_vector(31 downto 0) ;
    o_label1_config : out std_logic_vector(15 downto 0) ;
    o_label1_data7 : out std_logic_vector(31 downto 0) ;
    o_label1_data6 : out std_logic_vector(31 downto 0) ;
    o_label1_data5 : out std_logic_vector(31 downto 0) ;
    o_label1_data4 : out std_logic_vector(31 downto 0) ;
    o_label1_data3 : out std_logic_vector(31 downto 0) ;
    o_label1_data2 : out std_logic_vector(31 downto 0) ;
    o_label1_data1 : out std_logic_vector(31 downto 0) ;
    o_label1_data0 : out std_logic_vector(31 downto 0) ;
    o_label2_config : out std_logic_vector(15 downto 0) ;
    o_label2_data7 : out std_logic_vector(31 downto 0) ;
    o_label2_data6 : out std_logic_vector(31 downto 0) ;
    o_label2_data5 : out std_logic_vector(31 downto 0) ;
    o_label2_data4 : out std_logic_vector(31 downto 0) ;
    o_label2_data3 : out std_logic_vector(31 downto 0) ;
    o_label2_data2 : out std_logic_vector(31 downto 0) ;
    o_label2_data1 : out std_logic_vector(31 downto 0) ;
    o_label2_data0 : out std_logic_vector(31 downto 0) ;
    o_label3_config : out std_logic_vector(15 downto 0) ;
    o_label3_data7 : out std_logic_vector(31 downto 0) ;
    o_label3_data6 : out std_logic_vector(31 downto 0) ;
    o_label3_data5 : out std_logic_vector(31 downto 0) ;
    o_label3_data4 : out std_logic_vector(31 downto 0) ;
    o_label3_data3 : out std_logic_vector(31 downto 0) ;
    o_label3_data2 : out std_logic_vector(31 downto 0) ;
    o_label3_data1 : out std_logic_vector(31 downto 0) ;
    o_label3_data0 : out std_logic_vector(31 downto 0) ;
    o_label4_config : out std_logic_vector(15 downto 0) ;
    o_label4_data7 : out std_logic_vector(31 downto 0) ;
    o_label4_data6 : out std_logic_vector(31 downto 0) ;
    o_label4_data5 : out std_logic_vector(31 downto 0) ;
    o_label4_data4 : out std_logic_vector(31 downto 0) ;
    o_label4_data3 : out std_logic_vector(31 downto 0) ;
    o_label4_data2 : out std_logic_vector(31 downto 0) ;
    o_label4_data1 : out std_logic_vector(31 downto 0) ;
    o_label4_data0 : out std_logic_vector(31 downto 0) ;
    o_label5_config : out std_logic_vector(15 downto 0) ;
    o_label5_data7 : out std_logic_vector(31 downto 0) ;
    o_label5_data6 : out std_logic_vector(31 downto 0) ;
    o_label5_data5 : out std_logic_vector(31 downto 0) ;
    o_label5_data4 : out std_logic_vector(31 downto 0) ;
    o_label5_data3 : out std_logic_vector(31 downto 0) ;
    o_label5_data2 : out std_logic_vector(31 downto 0) ;
    o_label5_data1 : out std_logic_vector(31 downto 0) ;
    o_label5_data0 : out std_logic_vector(31 downto 0) ;
    o_label6_config : out std_logic_vector(15 downto 0) ;
    o_label6_data7 : out std_logic_vector(31 downto 0) ;
    o_label6_data6 : out std_logic_vector(31 downto 0) ;
    o_label6_data5 : out std_logic_vector(31 downto 0) ;
    o_label6_data4 : out std_logic_vector(31 downto 0) ;
    o_label6_data3 : out std_logic_vector(31 downto 0) ;
    o_label6_data2 : out std_logic_vector(31 downto 0) ;
    o_label6_data1 : out std_logic_vector(31 downto 0) ;
    o_label6_data0 : out std_logic_vector(31 downto 0) ;
    o_label7_config : out std_logic_vector(15 downto 0) ;
    o_label7_data7 : out std_logic_vector(31 downto 0) ;
    o_label7_data6 : out std_logic_vector(31 downto 0) ;
    o_label7_data5 : out std_logic_vector(31 downto 0) ;
    o_label7_data4 : out std_logic_vector(31 downto 0) ;
    o_label7_data3 : out std_logic_vector(31 downto 0) ;
    o_label7_data2 : out std_logic_vector(31 downto 0) ;
    o_label7_data1 : out std_logic_vector(31 downto 0) ;
    o_label7_data0 : out std_logic_vector(31 downto 0) ;
    o_kdf_drbg_ctrl : out std_logic_vector(1 downto 0) ;
    o_kdf_drbg_seed_0_state_key_31_0 : out std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_0_state_key_63_32 : out std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_0_state_key_95_64 : out std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_0_state_key_127_96 : out std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_0_state_key_159_128 : out std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_0_state_key_191_160 : out std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_0_state_key_223_192 : out std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_0_state_key_255_224 : out std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_0_state_value_31_0 : out std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_0_state_value_63_32 : out std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_0_state_value_95_64 : out std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_0_state_value_127_96 : out std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_0_reseed_interval_0 : out std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_0_reseed_interval_1 : out std_logic_vector(15 downto 0) ;
    o_kdf_drbg_seed_1_state_key_31_0 : out std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_1_state_key_63_32 : out std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_1_state_key_95_64 : out std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_1_state_key_127_96 : out std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_1_state_key_159_128 : out std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_1_state_key_191_160 : out std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_1_state_key_223_192 : out std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_1_state_key_255_224 : out std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_1_state_value_31_0 : out std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_1_state_value_63_32 : out std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_1_state_value_95_64 : out std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_1_state_value_127_96 : out std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_1_reseed_interval_0 : out std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_1_reseed_interval_1 : out std_logic_vector(15 downto 0) ;
    o_interrupt_status : out std_logic_vector(4 downto 0) ;
    o_interrupt_mask : out std_logic_vector(4 downto 0) ;
    o_engine_sticky_status : out std_logic_vector(7 downto 0) ;
    o_bimc_monitor_mask : out std_logic_vector(6 downto 0) ;
    o_bimc_ecc_uncorrectable_error_cnt : out std_logic_vector(31 downto 0) ;
    o_bimc_ecc_correctable_error_cnt : out std_logic_vector(31 downto 0) ;
    o_bimc_parity_error_cnt : out std_logic_vector(31 downto 0) ;
    o_bimc_global_config : out std_logic_vector(31 downto 0) ;
    o_bimc_eccpar_debug : out std_logic_vector(28 downto 0) ;
    o_bimc_cmd2 : out std_logic_vector(10 downto 0) ;
    o_bimc_cmd1 : out std_logic_vector(31 downto 0) ;
    o_bimc_cmd0 : out std_logic_vector(31 downto 0) ;
    o_bimc_rxcmd2 : out std_logic_vector(9 downto 0) ;
    o_bimc_rxrsp2 : out std_logic_vector(9 downto 0) ;
    o_bimc_pollrsp2 : out std_logic_vector(9 downto 0) ;
    o_bimc_dbgcmd2 : out std_logic_vector(9 downto 0) ;
    o_im_consumed : out std_logic_vector(15 downto 0) ;
    o_tready_override : out std_logic_vector(8 downto 0) ;
    o_regs_sa_ctrl : out std_logic_vector(31 downto 0) ;
    o_sa_snapshot_ia_wdata_part0 : out std_logic_vector(31 downto 0) ;
    o_sa_snapshot_ia_wdata_part1 : out std_logic_vector(31 downto 0) ;
    o_sa_snapshot_ia_config : out std_logic_vector(8 downto 0) ;
    o_sa_count_ia_wdata_part0 : out std_logic_vector(31 downto 0) ;
    o_sa_count_ia_wdata_part1 : out std_logic_vector(31 downto 0) ;
    o_sa_count_ia_config : out std_logic_vector(8 downto 0) ;
    o_cceip_encrypt_kop_fifo_override : out std_logic_vector(6 downto 0) ;
    o_cceip_validate_kop_fifo_override : out std_logic_vector(6 downto 0) ;
    o_cddip_decrypt_kop_fifo_override : out std_logic_vector(6 downto 0) ;
    o_sa_global_ctrl : out std_logic_vector(31 downto 0) ;
    o_sa_ctrl_ia_wdata_part0 : out std_logic_vector(31 downto 0) ;
    o_sa_ctrl_ia_config : out std_logic_vector(8 downto 0) ;
    o_kdf_test_key_size_config : out std_logic_vector(31 downto 0) ;
    i_blkid_revid_config : in std_logic_vector(31 downto 0) ;
    i_revision_config : in std_logic_vector(7 downto 0) ;
    i_spare_config : in std_logic_vector(31 downto 0) ;
    i_cceip0_out_ia_capability : in std_logic_vector(19 downto 0) ;
    i_cceip0_out_ia_status : in std_logic_vector(16 downto 0) ;
    i_cceip0_out_ia_rdata_part0 : in std_logic_vector(31 downto 0) ;
    i_cceip0_out_ia_rdata_part1 : in std_logic_vector(31 downto 0) ;
    i_cceip0_out_ia_rdata_part2 : in std_logic_vector(31 downto 0) ;
    i_cceip0_out_im_status : in std_logic_vector(11 downto 0) ;
    i_cceip0_out_im_read_done : in std_logic_vector(1 downto 0) ;
    i_cceip1_out_ia_capability : in std_logic_vector(19 downto 0) ;
    i_cceip1_out_ia_status : in std_logic_vector(16 downto 0) ;
    i_cceip1_out_ia_rdata_part0 : in std_logic_vector(31 downto 0) ;
    i_cceip1_out_ia_rdata_part1 : in std_logic_vector(31 downto 0) ;
    i_cceip1_out_ia_rdata_part2 : in std_logic_vector(31 downto 0) ;
    i_cceip1_out_im_status : in std_logic_vector(11 downto 0) ;
    i_cceip1_out_im_read_done : in std_logic_vector(1 downto 0) ;
    i_cceip2_out_ia_capability : in std_logic_vector(19 downto 0) ;
    i_cceip2_out_ia_status : in std_logic_vector(16 downto 0) ;
    i_cceip2_out_ia_rdata_part0 : in std_logic_vector(31 downto 0) ;
    i_cceip2_out_ia_rdata_part1 : in std_logic_vector(31 downto 0) ;
    i_cceip2_out_ia_rdata_part2 : in std_logic_vector(31 downto 0) ;
    i_cceip2_out_im_status : in std_logic_vector(11 downto 0) ;
    i_cceip2_out_im_read_done : in std_logic_vector(1 downto 0) ;
    i_cceip3_out_ia_capability : in std_logic_vector(19 downto 0) ;
    i_cceip3_out_ia_status : in std_logic_vector(16 downto 0) ;
    i_cceip3_out_ia_rdata_part0 : in std_logic_vector(31 downto 0) ;
    i_cceip3_out_ia_rdata_part1 : in std_logic_vector(31 downto 0) ;
    i_cceip3_out_ia_rdata_part2 : in std_logic_vector(31 downto 0) ;
    i_cceip3_out_im_status : in std_logic_vector(11 downto 0) ;
    i_cceip3_out_im_read_done : in std_logic_vector(1 downto 0) ;
    i_cddip0_out_ia_capability : in std_logic_vector(19 downto 0) ;
    i_cddip0_out_ia_status : in std_logic_vector(16 downto 0) ;
    i_cddip0_out_ia_rdata_part0 : in std_logic_vector(31 downto 0) ;
    i_cddip0_out_ia_rdata_part1 : in std_logic_vector(31 downto 0) ;
    i_cddip0_out_ia_rdata_part2 : in std_logic_vector(31 downto 0) ;
    i_cddip0_out_im_status : in std_logic_vector(11 downto 0) ;
    i_cddip0_out_im_read_done : in std_logic_vector(1 downto 0) ;
    i_cddip1_out_ia_capability : in std_logic_vector(19 downto 0) ;
    i_cddip1_out_ia_status : in std_logic_vector(16 downto 0) ;
    i_cddip1_out_ia_rdata_part0 : in std_logic_vector(31 downto 0) ;
    i_cddip1_out_ia_rdata_part1 : in std_logic_vector(31 downto 0) ;
    i_cddip1_out_ia_rdata_part2 : in std_logic_vector(31 downto 0) ;
    i_cddip1_out_im_status : in std_logic_vector(11 downto 0) ;
    i_cddip1_out_im_read_done : in std_logic_vector(1 downto 0) ;
    i_cddip2_out_ia_capability : in std_logic_vector(19 downto 0) ;
    i_cddip2_out_ia_status : in std_logic_vector(16 downto 0) ;
    i_cddip2_out_ia_rdata_part0 : in std_logic_vector(31 downto 0) ;
    i_cddip2_out_ia_rdata_part1 : in std_logic_vector(31 downto 0) ;
    i_cddip2_out_ia_rdata_part2 : in std_logic_vector(31 downto 0) ;
    i_cddip2_out_im_status : in std_logic_vector(11 downto 0) ;
    i_cddip2_out_im_read_done : in std_logic_vector(1 downto 0) ;
    i_cddip3_out_ia_capability : in std_logic_vector(19 downto 0) ;
    i_cddip3_out_ia_status : in std_logic_vector(16 downto 0) ;
    i_cddip3_out_ia_rdata_part0 : in std_logic_vector(31 downto 0) ;
    i_cddip3_out_ia_rdata_part1 : in std_logic_vector(31 downto 0) ;
    i_cddip3_out_ia_rdata_part2 : in std_logic_vector(31 downto 0) ;
    i_cddip3_out_im_status : in std_logic_vector(11 downto 0) ;
    i_cddip3_out_im_read_done : in std_logic_vector(1 downto 0) ;
    i_ckv_ia_capability : in std_logic_vector(19 downto 0) ;
    i_ckv_ia_status : in std_logic_vector(22 downto 0) ;
    i_ckv_ia_rdata_part0 : in std_logic_vector(31 downto 0) ;
    i_ckv_ia_rdata_part1 : in std_logic_vector(31 downto 0) ;
    i_kim_ia_capability : in std_logic_vector(19 downto 0) ;
    i_kim_ia_status : in std_logic_vector(21 downto 0) ;
    i_kim_ia_rdata_part0 : in std_logic_vector(20 downto 0) ;
    i_kim_ia_rdata_part1 : in std_logic_vector(16 downto 0) ;
    i_kdf_drbg_ctrl : in std_logic_vector(1 downto 0) ;
    i_interrupt_status : in std_logic_vector(4 downto 0) ;
    i_engine_sticky_status : in std_logic_vector(7 downto 0) ;
    i_bimc_monitor : in std_logic_vector(6 downto 0) ;
    i_bimc_ecc_uncorrectable_error_cnt : in std_logic_vector(31 downto 0) ;
    i_bimc_ecc_correctable_error_cnt : in std_logic_vector(31 downto 0) ;
    i_bimc_parity_error_cnt : in std_logic_vector(31 downto 0) ;
    i_bimc_global_config : in std_logic_vector(31 downto 0) ;
    i_bimc_memid : in std_logic_vector(11 downto 0) ;
    i_bimc_eccpar_debug : in std_logic_vector(28 downto 0) ;
    i_bimc_cmd2 : in std_logic_vector(10 downto 0) ;
    i_bimc_rxcmd2 : in std_logic_vector(9 downto 0) ;
    i_bimc_rxcmd1 : in std_logic_vector(31 downto 0) ;
    i_bimc_rxcmd0 : in std_logic_vector(31 downto 0) ;
    i_bimc_rxrsp2 : in std_logic_vector(9 downto 0) ;
    i_bimc_rxrsp1 : in std_logic_vector(31 downto 0) ;
    i_bimc_rxrsp0 : in std_logic_vector(31 downto 0) ;
    i_bimc_pollrsp2 : in std_logic_vector(9 downto 0) ;
    i_bimc_pollrsp1 : in std_logic_vector(31 downto 0) ;
    i_bimc_pollrsp0 : in std_logic_vector(31 downto 0) ;
    i_bimc_dbgcmd2 : in std_logic_vector(9 downto 0) ;
    i_bimc_dbgcmd1 : in std_logic_vector(31 downto 0) ;
    i_bimc_dbgcmd0 : in std_logic_vector(31 downto 0) ;
    i_im_available : in std_logic_vector(15 downto 0) ;
    i_im_consumed : in std_logic_vector(15 downto 0) ;
    i_tready_override : in std_logic_vector(8 downto 0) ;
    i_regs_sa_ctrl : in std_logic_vector(31 downto 0) ;
    i_sa_snapshot_ia_capability : in std_logic_vector(19 downto 0) ;
    i_sa_snapshot_ia_status : in std_logic_vector(12 downto 0) ;
    i_sa_snapshot_ia_rdata_part0 : in std_logic_vector(31 downto 0) ;
    i_sa_snapshot_ia_rdata_part1 : in std_logic_vector(31 downto 0) ;
    i_sa_count_ia_capability : in std_logic_vector(19 downto 0) ;
    i_sa_count_ia_status : in std_logic_vector(12 downto 0) ;
    i_sa_count_ia_rdata_part0 : in std_logic_vector(31 downto 0) ;
    i_sa_count_ia_rdata_part1 : in std_logic_vector(31 downto 0) ;
    i_idle_components : in std_logic_vector(31 downto 0) ;
    i_sa_global_ctrl : in std_logic_vector(31 downto 0) ;
    i_sa_ctrl_ia_capability : in std_logic_vector(19 downto 0) ;
    i_sa_ctrl_ia_status : in std_logic_vector(12 downto 0) ;
    i_sa_ctrl_ia_rdata_part0 : in std_logic_vector(31 downto 0) ;
    o_reg_written : out std_logic ;
    o_reg_read : out std_logic ;
    o_reg_wr_data : out std_logic_vector(31 downto 0) ;
  o_reg_addr : out std_logic_vector(10 downto 0) ) ;
  attribute _2_state_: integer;
end cr_kme_regs ;
