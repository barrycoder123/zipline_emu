
module xcva_top ;
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
kme_tb kme_tb ();
my_clks my_clks ();
IXC_GFIFO IXC_GFIFO ();
ixc_time ixc_time ();
_ixc_isc _ixc_isc ();
xc_top_1 xc_top ();
ASSERTION ASSERTION ();
// pragma CVASTRPROP MODULE HDLICE PROP_IXCOM_MOD TRUE
endmodule
