
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
`_2_ (* upf_always_on = 1 *) 
module ixc_gfifo_port_560_3 ( tkout, tkin, ireq, cbid, len, idata, CGFtsReq, 
	CGFcbid, CGFlen, CGFidata, CGFfull, CLBreq, CLBrd, CLBwr, CLBfull, 
	Rtkin);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output tkout;
input tkin;
input ireq;
input [19:0] cbid;
input [11:0] len;
input [559:0] idata;
output CGFtsReq;
output [19:0] CGFcbid;
output [11:0] CGFlen;
output [511:0] CGFidata;
input CGFfull;
output CLBreq;
input [3:0] CLBrd;
input [3:0] CLBwr;
input CLBfull;
input Rtkin;
wire fclk;
wire enq;
wire CLBreqWhileFull;
`_2_ wire en;
`_2_ wire ack;
`_2_ wire [559:0] odata;
`_2_ wire oreq;
`_2_ wire [19:0] ocbid;
`_2_ wire [19:0] xcbid;
`_2_ wire [11:0] olen;
`_2_ wire [11:0] xlen;
`_2_ wire [1:0] sel;
`_2_ wire [511:0] xdata;
wire [31:0] i;
`_2_ wire ireqR;
wire State_Var;
supply1 n6;
Q_AN02 U0 ( .A0(n169), .A1(n113), .Z(n1));
Q_NOT_TOUCH _zzqnthw ( .sig());
Q_EV_WOR_START qi ( .A(CLBreqWhileFull));
Q_INV U3 ( .A(n5), .Z(tkout));
Q_XNR2 U4 ( .A0(oreq), .A1(ack), .Z(n5));
Q_CCLKCHK cchk ( .sig(ireq));
Q_AN02 U6 ( .A0(enq), .A1(CLBfull), .Z(CLBreqWhileFull));
Q_AN02 U7 ( .A0(n3), .A1(n4), .Z(enq));
Q_INV U8 ( .A(xc_top.GFLock2), .Z(n4));
Q_XOR2 U9 ( .A0(ireq), .A1(ireqR), .Z(n3));
Q_BUFZP U10 ( .OE(CLBreqWhileFull), .A(n6), .Z(xc_top.GFLBfull));
Q_BUFZP U11 ( .OE(en), .A(xcbid[0]), .Z(CGFcbid[0]));
Q_BUFZP U12 ( .OE(en), .A(xcbid[1]), .Z(CGFcbid[1]));
Q_BUFZP U13 ( .OE(en), .A(xcbid[2]), .Z(CGFcbid[2]));
Q_BUFZP U14 ( .OE(en), .A(xcbid[3]), .Z(CGFcbid[3]));
Q_BUFZP U15 ( .OE(en), .A(xcbid[4]), .Z(CGFcbid[4]));
Q_BUFZP U16 ( .OE(en), .A(xcbid[5]), .Z(CGFcbid[5]));
Q_BUFZP U17 ( .OE(en), .A(xcbid[6]), .Z(CGFcbid[6]));
Q_BUFZP U18 ( .OE(en), .A(xcbid[7]), .Z(CGFcbid[7]));
Q_BUFZP U19 ( .OE(en), .A(xcbid[8]), .Z(CGFcbid[8]));
Q_BUFZP U20 ( .OE(en), .A(xcbid[9]), .Z(CGFcbid[9]));
Q_BUFZP U21 ( .OE(en), .A(xcbid[10]), .Z(CGFcbid[10]));
Q_BUFZP U22 ( .OE(en), .A(xcbid[11]), .Z(CGFcbid[11]));
Q_BUFZP U23 ( .OE(en), .A(xcbid[12]), .Z(CGFcbid[12]));
Q_BUFZP U24 ( .OE(en), .A(xcbid[13]), .Z(CGFcbid[13]));
Q_BUFZP U25 ( .OE(en), .A(xcbid[14]), .Z(CGFcbid[14]));
Q_BUFZP U26 ( .OE(en), .A(xcbid[15]), .Z(CGFcbid[15]));
Q_BUFZP U27 ( .OE(en), .A(xcbid[16]), .Z(CGFcbid[16]));
Q_BUFZP U28 ( .OE(en), .A(xcbid[17]), .Z(CGFcbid[17]));
Q_BUFZP U29 ( .OE(en), .A(xcbid[18]), .Z(CGFcbid[18]));
Q_BUFZP U30 ( .OE(en), .A(xcbid[19]), .Z(CGFcbid[19]));
Q_BUFZP U31 ( .OE(en), .A(xlen[0]), .Z(CGFlen[0]));
Q_BUFZP U32 ( .OE(en), .A(xlen[1]), .Z(CGFlen[1]));
Q_BUFZP U33 ( .OE(en), .A(xlen[2]), .Z(CGFlen[2]));
Q_BUFZP U34 ( .OE(en), .A(xlen[3]), .Z(CGFlen[3]));
Q_BUFZP U35 ( .OE(en), .A(xlen[4]), .Z(CGFlen[4]));
Q_BUFZP U36 ( .OE(en), .A(xlen[5]), .Z(CGFlen[5]));
Q_BUFZP U37 ( .OE(en), .A(xlen[6]), .Z(CGFlen[6]));
Q_BUFZP U38 ( .OE(en), .A(xlen[7]), .Z(CGFlen[7]));
Q_BUFZP U39 ( .OE(en), .A(xlen[8]), .Z(CGFlen[8]));
Q_BUFZP U40 ( .OE(en), .A(xlen[9]), .Z(CGFlen[9]));
Q_BUFZP U41 ( .OE(en), .A(xlen[10]), .Z(CGFlen[10]));
Q_BUFZP U42 ( .OE(en), .A(xlen[11]), .Z(CGFlen[11]));
Q_BUFZP U43 ( .OE(en), .A(xdata[0]), .Z(CGFidata[0]));
Q_BUFZP U44 ( .OE(en), .A(xdata[1]), .Z(CGFidata[1]));
Q_BUFZP U45 ( .OE(en), .A(xdata[2]), .Z(CGFidata[2]));
Q_BUFZP U46 ( .OE(en), .A(xdata[3]), .Z(CGFidata[3]));
Q_BUFZP U47 ( .OE(en), .A(xdata[4]), .Z(CGFidata[4]));
Q_BUFZP U48 ( .OE(en), .A(xdata[5]), .Z(CGFidata[5]));
Q_BUFZP U49 ( .OE(en), .A(xdata[6]), .Z(CGFidata[6]));
Q_BUFZP U50 ( .OE(en), .A(xdata[7]), .Z(CGFidata[7]));
Q_BUFZP U51 ( .OE(en), .A(xdata[8]), .Z(CGFidata[8]));
Q_BUFZP U52 ( .OE(en), .A(xdata[9]), .Z(CGFidata[9]));
Q_BUFZP U53 ( .OE(en), .A(xdata[10]), .Z(CGFidata[10]));
Q_BUFZP U54 ( .OE(en), .A(xdata[11]), .Z(CGFidata[11]));
Q_BUFZP U55 ( .OE(en), .A(xdata[12]), .Z(CGFidata[12]));
Q_BUFZP U56 ( .OE(en), .A(xdata[13]), .Z(CGFidata[13]));
Q_BUFZP U57 ( .OE(en), .A(xdata[14]), .Z(CGFidata[14]));
Q_BUFZP U58 ( .OE(en), .A(xdata[15]), .Z(CGFidata[15]));
Q_BUFZP U59 ( .OE(en), .A(xdata[16]), .Z(CGFidata[16]));
Q_BUFZP U60 ( .OE(en), .A(xdata[17]), .Z(CGFidata[17]));
Q_BUFZP U61 ( .OE(en), .A(xdata[18]), .Z(CGFidata[18]));
Q_BUFZP U62 ( .OE(en), .A(xdata[19]), .Z(CGFidata[19]));
Q_BUFZP U63 ( .OE(en), .A(xdata[20]), .Z(CGFidata[20]));
Q_BUFZP U64 ( .OE(en), .A(xdata[21]), .Z(CGFidata[21]));
Q_BUFZP U65 ( .OE(en), .A(xdata[22]), .Z(CGFidata[22]));
Q_BUFZP U66 ( .OE(en), .A(xdata[23]), .Z(CGFidata[23]));
Q_BUFZP U67 ( .OE(en), .A(xdata[24]), .Z(CGFidata[24]));
Q_BUFZP U68 ( .OE(en), .A(xdata[25]), .Z(CGFidata[25]));
Q_BUFZP U69 ( .OE(en), .A(xdata[26]), .Z(CGFidata[26]));
Q_BUFZP U70 ( .OE(en), .A(xdata[27]), .Z(CGFidata[27]));
Q_BUFZP U71 ( .OE(en), .A(xdata[28]), .Z(CGFidata[28]));
Q_BUFZP U72 ( .OE(en), .A(xdata[29]), .Z(CGFidata[29]));
Q_BUFZP U73 ( .OE(en), .A(xdata[30]), .Z(CGFidata[30]));
Q_BUFZP U74 ( .OE(en), .A(xdata[31]), .Z(CGFidata[31]));
Q_BUFZP U75 ( .OE(en), .A(xdata[32]), .Z(CGFidata[32]));
Q_BUFZP U76 ( .OE(en), .A(xdata[33]), .Z(CGFidata[33]));
Q_BUFZP U77 ( .OE(en), .A(xdata[34]), .Z(CGFidata[34]));
Q_BUFZP U78 ( .OE(en), .A(xdata[35]), .Z(CGFidata[35]));
Q_BUFZP U79 ( .OE(en), .A(xdata[36]), .Z(CGFidata[36]));
Q_BUFZP U80 ( .OE(en), .A(xdata[37]), .Z(CGFidata[37]));
Q_BUFZP U81 ( .OE(en), .A(xdata[38]), .Z(CGFidata[38]));
Q_BUFZP U82 ( .OE(en), .A(xdata[39]), .Z(CGFidata[39]));
Q_BUFZP U83 ( .OE(en), .A(xdata[40]), .Z(CGFidata[40]));
Q_BUFZP U84 ( .OE(en), .A(xdata[41]), .Z(CGFidata[41]));
Q_BUFZP U85 ( .OE(en), .A(xdata[42]), .Z(CGFidata[42]));
Q_BUFZP U86 ( .OE(en), .A(xdata[43]), .Z(CGFidata[43]));
Q_BUFZP U87 ( .OE(en), .A(xdata[44]), .Z(CGFidata[44]));
Q_BUFZP U88 ( .OE(en), .A(xdata[45]), .Z(CGFidata[45]));
Q_BUFZP U89 ( .OE(en), .A(xdata[46]), .Z(CGFidata[46]));
Q_BUFZP U90 ( .OE(en), .A(xdata[47]), .Z(CGFidata[47]));
Q_BUFZP U91 ( .OE(en), .A(xdata[48]), .Z(CGFidata[48]));
Q_BUFZP U92 ( .OE(en), .A(xdata[49]), .Z(CGFidata[49]));
Q_BUFZP U93 ( .OE(en), .A(xdata[50]), .Z(CGFidata[50]));
Q_BUFZP U94 ( .OE(en), .A(xdata[51]), .Z(CGFidata[51]));
Q_BUFZP U95 ( .OE(en), .A(xdata[52]), .Z(CGFidata[52]));
Q_BUFZP U96 ( .OE(en), .A(xdata[53]), .Z(CGFidata[53]));
Q_BUFZP U97 ( .OE(en), .A(xdata[54]), .Z(CGFidata[54]));
Q_BUFZP U98 ( .OE(en), .A(xdata[55]), .Z(CGFidata[55]));
Q_BUFZP U99 ( .OE(en), .A(xdata[56]), .Z(CGFidata[56]));
Q_BUFZP U100 ( .OE(en), .A(xdata[57]), .Z(CGFidata[57]));
Q_BUFZP U101 ( .OE(en), .A(xdata[58]), .Z(CGFidata[58]));
Q_BUFZP U102 ( .OE(en), .A(xdata[59]), .Z(CGFidata[59]));
Q_BUFZP U103 ( .OE(en), .A(xdata[60]), .Z(CGFidata[60]));
Q_BUFZP U104 ( .OE(en), .A(xdata[61]), .Z(CGFidata[61]));
Q_BUFZP U105 ( .OE(en), .A(xdata[62]), .Z(CGFidata[62]));
Q_BUFZP U106 ( .OE(en), .A(xdata[63]), .Z(CGFidata[63]));
Q_BUFZP U107 ( .OE(en), .A(xdata[64]), .Z(CGFidata[64]));
Q_BUFZP U108 ( .OE(en), .A(xdata[65]), .Z(CGFidata[65]));
Q_BUFZP U109 ( .OE(en), .A(xdata[66]), .Z(CGFidata[66]));
Q_BUFZP U110 ( .OE(en), .A(xdata[67]), .Z(CGFidata[67]));
Q_BUFZP U111 ( .OE(en), .A(xdata[68]), .Z(CGFidata[68]));
Q_BUFZP U112 ( .OE(en), .A(xdata[69]), .Z(CGFidata[69]));
Q_BUFZP U113 ( .OE(en), .A(xdata[70]), .Z(CGFidata[70]));
Q_BUFZP U114 ( .OE(en), .A(xdata[71]), .Z(CGFidata[71]));
Q_BUFZP U115 ( .OE(en), .A(xdata[72]), .Z(CGFidata[72]));
Q_BUFZP U116 ( .OE(en), .A(xdata[73]), .Z(CGFidata[73]));
Q_BUFZP U117 ( .OE(en), .A(xdata[74]), .Z(CGFidata[74]));
Q_BUFZP U118 ( .OE(en), .A(xdata[75]), .Z(CGFidata[75]));
Q_BUFZP U119 ( .OE(en), .A(xdata[76]), .Z(CGFidata[76]));
Q_BUFZP U120 ( .OE(en), .A(xdata[77]), .Z(CGFidata[77]));
Q_BUFZP U121 ( .OE(en), .A(xdata[78]), .Z(CGFidata[78]));
Q_BUFZP U122 ( .OE(en), .A(xdata[79]), .Z(CGFidata[79]));
Q_BUFZP U123 ( .OE(en), .A(xdata[80]), .Z(CGFidata[80]));
Q_BUFZP U124 ( .OE(en), .A(xdata[81]), .Z(CGFidata[81]));
Q_BUFZP U125 ( .OE(en), .A(xdata[82]), .Z(CGFidata[82]));
Q_BUFZP U126 ( .OE(en), .A(xdata[83]), .Z(CGFidata[83]));
Q_BUFZP U127 ( .OE(en), .A(xdata[84]), .Z(CGFidata[84]));
Q_BUFZP U128 ( .OE(en), .A(xdata[85]), .Z(CGFidata[85]));
Q_BUFZP U129 ( .OE(en), .A(xdata[86]), .Z(CGFidata[86]));
Q_BUFZP U130 ( .OE(en), .A(xdata[87]), .Z(CGFidata[87]));
Q_BUFZP U131 ( .OE(en), .A(xdata[88]), .Z(CGFidata[88]));
Q_BUFZP U132 ( .OE(en), .A(xdata[89]), .Z(CGFidata[89]));
Q_BUFZP U133 ( .OE(en), .A(xdata[90]), .Z(CGFidata[90]));
Q_BUFZP U134 ( .OE(en), .A(xdata[91]), .Z(CGFidata[91]));
Q_BUFZP U135 ( .OE(en), .A(xdata[92]), .Z(CGFidata[92]));
Q_BUFZP U136 ( .OE(en), .A(xdata[93]), .Z(CGFidata[93]));
Q_BUFZP U137 ( .OE(en), .A(xdata[94]), .Z(CGFidata[94]));
Q_BUFZP U138 ( .OE(en), .A(xdata[95]), .Z(CGFidata[95]));
Q_BUFZP U139 ( .OE(en), .A(xdata[96]), .Z(CGFidata[96]));
Q_BUFZP U140 ( .OE(en), .A(xdata[97]), .Z(CGFidata[97]));
Q_BUFZP U141 ( .OE(en), .A(xdata[98]), .Z(CGFidata[98]));
Q_BUFZP U142 ( .OE(en), .A(xdata[99]), .Z(CGFidata[99]));
Q_BUFZP U143 ( .OE(en), .A(xdata[100]), .Z(CGFidata[100]));
Q_BUFZP U144 ( .OE(en), .A(xdata[101]), .Z(CGFidata[101]));
Q_BUFZP U145 ( .OE(en), .A(xdata[102]), .Z(CGFidata[102]));
Q_BUFZP U146 ( .OE(en), .A(xdata[103]), .Z(CGFidata[103]));
Q_BUFZP U147 ( .OE(en), .A(xdata[104]), .Z(CGFidata[104]));
Q_BUFZP U148 ( .OE(en), .A(xdata[105]), .Z(CGFidata[105]));
Q_BUFZP U149 ( .OE(en), .A(xdata[106]), .Z(CGFidata[106]));
Q_BUFZP U150 ( .OE(en), .A(xdata[107]), .Z(CGFidata[107]));
Q_BUFZP U151 ( .OE(en), .A(xdata[108]), .Z(CGFidata[108]));
Q_BUFZP U152 ( .OE(en), .A(xdata[109]), .Z(CGFidata[109]));
Q_BUFZP U153 ( .OE(en), .A(xdata[110]), .Z(CGFidata[110]));
Q_BUFZP U154 ( .OE(en), .A(xdata[111]), .Z(CGFidata[111]));
Q_BUFZP U155 ( .OE(en), .A(xdata[112]), .Z(CGFidata[112]));
Q_BUFZP U156 ( .OE(en), .A(xdata[113]), .Z(CGFidata[113]));
Q_BUFZP U157 ( .OE(en), .A(xdata[114]), .Z(CGFidata[114]));
Q_BUFZP U158 ( .OE(en), .A(xdata[115]), .Z(CGFidata[115]));
Q_BUFZP U159 ( .OE(en), .A(xdata[116]), .Z(CGFidata[116]));
Q_BUFZP U160 ( .OE(en), .A(xdata[117]), .Z(CGFidata[117]));
Q_BUFZP U161 ( .OE(en), .A(xdata[118]), .Z(CGFidata[118]));
Q_BUFZP U162 ( .OE(en), .A(xdata[119]), .Z(CGFidata[119]));
Q_BUFZP U163 ( .OE(en), .A(xdata[120]), .Z(CGFidata[120]));
Q_BUFZP U164 ( .OE(en), .A(xdata[121]), .Z(CGFidata[121]));
Q_BUFZP U165 ( .OE(en), .A(xdata[122]), .Z(CGFidata[122]));
Q_BUFZP U166 ( .OE(en), .A(xdata[123]), .Z(CGFidata[123]));
Q_BUFZP U167 ( .OE(en), .A(xdata[124]), .Z(CGFidata[124]));
Q_BUFZP U168 ( .OE(en), .A(xdata[125]), .Z(CGFidata[125]));
Q_BUFZP U169 ( .OE(en), .A(xdata[126]), .Z(CGFidata[126]));
Q_BUFZP U170 ( .OE(en), .A(xdata[127]), .Z(CGFidata[127]));
Q_BUFZP U171 ( .OE(en), .A(xdata[128]), .Z(CGFidata[128]));
Q_BUFZP U172 ( .OE(en), .A(xdata[129]), .Z(CGFidata[129]));
Q_BUFZP U173 ( .OE(en), .A(xdata[130]), .Z(CGFidata[130]));
Q_BUFZP U174 ( .OE(en), .A(xdata[131]), .Z(CGFidata[131]));
Q_BUFZP U175 ( .OE(en), .A(xdata[132]), .Z(CGFidata[132]));
Q_BUFZP U176 ( .OE(en), .A(xdata[133]), .Z(CGFidata[133]));
Q_BUFZP U177 ( .OE(en), .A(xdata[134]), .Z(CGFidata[134]));
Q_BUFZP U178 ( .OE(en), .A(xdata[135]), .Z(CGFidata[135]));
Q_BUFZP U179 ( .OE(en), .A(xdata[136]), .Z(CGFidata[136]));
Q_BUFZP U180 ( .OE(en), .A(xdata[137]), .Z(CGFidata[137]));
Q_BUFZP U181 ( .OE(en), .A(xdata[138]), .Z(CGFidata[138]));
Q_BUFZP U182 ( .OE(en), .A(xdata[139]), .Z(CGFidata[139]));
Q_BUFZP U183 ( .OE(en), .A(xdata[140]), .Z(CGFidata[140]));
Q_BUFZP U184 ( .OE(en), .A(xdata[141]), .Z(CGFidata[141]));
Q_BUFZP U185 ( .OE(en), .A(xdata[142]), .Z(CGFidata[142]));
Q_BUFZP U186 ( .OE(en), .A(xdata[143]), .Z(CGFidata[143]));
Q_BUFZP U187 ( .OE(en), .A(xdata[144]), .Z(CGFidata[144]));
Q_BUFZP U188 ( .OE(en), .A(xdata[145]), .Z(CGFidata[145]));
Q_BUFZP U189 ( .OE(en), .A(xdata[146]), .Z(CGFidata[146]));
Q_BUFZP U190 ( .OE(en), .A(xdata[147]), .Z(CGFidata[147]));
Q_BUFZP U191 ( .OE(en), .A(xdata[148]), .Z(CGFidata[148]));
Q_BUFZP U192 ( .OE(en), .A(xdata[149]), .Z(CGFidata[149]));
Q_BUFZP U193 ( .OE(en), .A(xdata[150]), .Z(CGFidata[150]));
Q_BUFZP U194 ( .OE(en), .A(xdata[151]), .Z(CGFidata[151]));
Q_BUFZP U195 ( .OE(en), .A(xdata[152]), .Z(CGFidata[152]));
Q_BUFZP U196 ( .OE(en), .A(xdata[153]), .Z(CGFidata[153]));
Q_BUFZP U197 ( .OE(en), .A(xdata[154]), .Z(CGFidata[154]));
Q_BUFZP U198 ( .OE(en), .A(xdata[155]), .Z(CGFidata[155]));
Q_BUFZP U199 ( .OE(en), .A(xdata[156]), .Z(CGFidata[156]));
Q_BUFZP U200 ( .OE(en), .A(xdata[157]), .Z(CGFidata[157]));
Q_BUFZP U201 ( .OE(en), .A(xdata[158]), .Z(CGFidata[158]));
Q_BUFZP U202 ( .OE(en), .A(xdata[159]), .Z(CGFidata[159]));
Q_BUFZP U203 ( .OE(en), .A(xdata[160]), .Z(CGFidata[160]));
Q_BUFZP U204 ( .OE(en), .A(xdata[161]), .Z(CGFidata[161]));
Q_BUFZP U205 ( .OE(en), .A(xdata[162]), .Z(CGFidata[162]));
Q_BUFZP U206 ( .OE(en), .A(xdata[163]), .Z(CGFidata[163]));
Q_BUFZP U207 ( .OE(en), .A(xdata[164]), .Z(CGFidata[164]));
Q_BUFZP U208 ( .OE(en), .A(xdata[165]), .Z(CGFidata[165]));
Q_BUFZP U209 ( .OE(en), .A(xdata[166]), .Z(CGFidata[166]));
Q_BUFZP U210 ( .OE(en), .A(xdata[167]), .Z(CGFidata[167]));
Q_BUFZP U211 ( .OE(en), .A(xdata[168]), .Z(CGFidata[168]));
Q_BUFZP U212 ( .OE(en), .A(xdata[169]), .Z(CGFidata[169]));
Q_BUFZP U213 ( .OE(en), .A(xdata[170]), .Z(CGFidata[170]));
Q_BUFZP U214 ( .OE(en), .A(xdata[171]), .Z(CGFidata[171]));
Q_BUFZP U215 ( .OE(en), .A(xdata[172]), .Z(CGFidata[172]));
Q_BUFZP U216 ( .OE(en), .A(xdata[173]), .Z(CGFidata[173]));
Q_BUFZP U217 ( .OE(en), .A(xdata[174]), .Z(CGFidata[174]));
Q_BUFZP U218 ( .OE(en), .A(xdata[175]), .Z(CGFidata[175]));
Q_BUFZP U219 ( .OE(en), .A(xdata[176]), .Z(CGFidata[176]));
Q_BUFZP U220 ( .OE(en), .A(xdata[177]), .Z(CGFidata[177]));
Q_BUFZP U221 ( .OE(en), .A(xdata[178]), .Z(CGFidata[178]));
Q_BUFZP U222 ( .OE(en), .A(xdata[179]), .Z(CGFidata[179]));
Q_BUFZP U223 ( .OE(en), .A(xdata[180]), .Z(CGFidata[180]));
Q_BUFZP U224 ( .OE(en), .A(xdata[181]), .Z(CGFidata[181]));
Q_BUFZP U225 ( .OE(en), .A(xdata[182]), .Z(CGFidata[182]));
Q_BUFZP U226 ( .OE(en), .A(xdata[183]), .Z(CGFidata[183]));
Q_BUFZP U227 ( .OE(en), .A(xdata[184]), .Z(CGFidata[184]));
Q_BUFZP U228 ( .OE(en), .A(xdata[185]), .Z(CGFidata[185]));
Q_BUFZP U229 ( .OE(en), .A(xdata[186]), .Z(CGFidata[186]));
Q_BUFZP U230 ( .OE(en), .A(xdata[187]), .Z(CGFidata[187]));
Q_BUFZP U231 ( .OE(en), .A(xdata[188]), .Z(CGFidata[188]));
Q_BUFZP U232 ( .OE(en), .A(xdata[189]), .Z(CGFidata[189]));
Q_BUFZP U233 ( .OE(en), .A(xdata[190]), .Z(CGFidata[190]));
Q_BUFZP U234 ( .OE(en), .A(xdata[191]), .Z(CGFidata[191]));
Q_BUFZP U235 ( .OE(en), .A(xdata[192]), .Z(CGFidata[192]));
Q_BUFZP U236 ( .OE(en), .A(xdata[193]), .Z(CGFidata[193]));
Q_BUFZP U237 ( .OE(en), .A(xdata[194]), .Z(CGFidata[194]));
Q_BUFZP U238 ( .OE(en), .A(xdata[195]), .Z(CGFidata[195]));
Q_BUFZP U239 ( .OE(en), .A(xdata[196]), .Z(CGFidata[196]));
Q_BUFZP U240 ( .OE(en), .A(xdata[197]), .Z(CGFidata[197]));
Q_BUFZP U241 ( .OE(en), .A(xdata[198]), .Z(CGFidata[198]));
Q_BUFZP U242 ( .OE(en), .A(xdata[199]), .Z(CGFidata[199]));
Q_BUFZP U243 ( .OE(en), .A(xdata[200]), .Z(CGFidata[200]));
Q_BUFZP U244 ( .OE(en), .A(xdata[201]), .Z(CGFidata[201]));
Q_BUFZP U245 ( .OE(en), .A(xdata[202]), .Z(CGFidata[202]));
Q_BUFZP U246 ( .OE(en), .A(xdata[203]), .Z(CGFidata[203]));
Q_BUFZP U247 ( .OE(en), .A(xdata[204]), .Z(CGFidata[204]));
Q_BUFZP U248 ( .OE(en), .A(xdata[205]), .Z(CGFidata[205]));
Q_BUFZP U249 ( .OE(en), .A(xdata[206]), .Z(CGFidata[206]));
Q_BUFZP U250 ( .OE(en), .A(xdata[207]), .Z(CGFidata[207]));
Q_BUFZP U251 ( .OE(en), .A(xdata[208]), .Z(CGFidata[208]));
Q_BUFZP U252 ( .OE(en), .A(xdata[209]), .Z(CGFidata[209]));
Q_BUFZP U253 ( .OE(en), .A(xdata[210]), .Z(CGFidata[210]));
Q_BUFZP U254 ( .OE(en), .A(xdata[211]), .Z(CGFidata[211]));
Q_BUFZP U255 ( .OE(en), .A(xdata[212]), .Z(CGFidata[212]));
Q_BUFZP U256 ( .OE(en), .A(xdata[213]), .Z(CGFidata[213]));
Q_BUFZP U257 ( .OE(en), .A(xdata[214]), .Z(CGFidata[214]));
Q_BUFZP U258 ( .OE(en), .A(xdata[215]), .Z(CGFidata[215]));
Q_BUFZP U259 ( .OE(en), .A(xdata[216]), .Z(CGFidata[216]));
Q_BUFZP U260 ( .OE(en), .A(xdata[217]), .Z(CGFidata[217]));
Q_BUFZP U261 ( .OE(en), .A(xdata[218]), .Z(CGFidata[218]));
Q_BUFZP U262 ( .OE(en), .A(xdata[219]), .Z(CGFidata[219]));
Q_BUFZP U263 ( .OE(en), .A(xdata[220]), .Z(CGFidata[220]));
Q_BUFZP U264 ( .OE(en), .A(xdata[221]), .Z(CGFidata[221]));
Q_BUFZP U265 ( .OE(en), .A(xdata[222]), .Z(CGFidata[222]));
Q_BUFZP U266 ( .OE(en), .A(xdata[223]), .Z(CGFidata[223]));
Q_BUFZP U267 ( .OE(en), .A(xdata[224]), .Z(CGFidata[224]));
Q_BUFZP U268 ( .OE(en), .A(xdata[225]), .Z(CGFidata[225]));
Q_BUFZP U269 ( .OE(en), .A(xdata[226]), .Z(CGFidata[226]));
Q_BUFZP U270 ( .OE(en), .A(xdata[227]), .Z(CGFidata[227]));
Q_BUFZP U271 ( .OE(en), .A(xdata[228]), .Z(CGFidata[228]));
Q_BUFZP U272 ( .OE(en), .A(xdata[229]), .Z(CGFidata[229]));
Q_BUFZP U273 ( .OE(en), .A(xdata[230]), .Z(CGFidata[230]));
Q_BUFZP U274 ( .OE(en), .A(xdata[231]), .Z(CGFidata[231]));
Q_BUFZP U275 ( .OE(en), .A(xdata[232]), .Z(CGFidata[232]));
Q_BUFZP U276 ( .OE(en), .A(xdata[233]), .Z(CGFidata[233]));
Q_BUFZP U277 ( .OE(en), .A(xdata[234]), .Z(CGFidata[234]));
Q_BUFZP U278 ( .OE(en), .A(xdata[235]), .Z(CGFidata[235]));
Q_BUFZP U279 ( .OE(en), .A(xdata[236]), .Z(CGFidata[236]));
Q_BUFZP U280 ( .OE(en), .A(xdata[237]), .Z(CGFidata[237]));
Q_BUFZP U281 ( .OE(en), .A(xdata[238]), .Z(CGFidata[238]));
Q_BUFZP U282 ( .OE(en), .A(xdata[239]), .Z(CGFidata[239]));
Q_BUFZP U283 ( .OE(en), .A(xdata[240]), .Z(CGFidata[240]));
Q_BUFZP U284 ( .OE(en), .A(xdata[241]), .Z(CGFidata[241]));
Q_BUFZP U285 ( .OE(en), .A(xdata[242]), .Z(CGFidata[242]));
Q_BUFZP U286 ( .OE(en), .A(xdata[243]), .Z(CGFidata[243]));
Q_BUFZP U287 ( .OE(en), .A(xdata[244]), .Z(CGFidata[244]));
Q_BUFZP U288 ( .OE(en), .A(xdata[245]), .Z(CGFidata[245]));
Q_BUFZP U289 ( .OE(en), .A(xdata[246]), .Z(CGFidata[246]));
Q_BUFZP U290 ( .OE(en), .A(xdata[247]), .Z(CGFidata[247]));
Q_BUFZP U291 ( .OE(en), .A(xdata[248]), .Z(CGFidata[248]));
Q_BUFZP U292 ( .OE(en), .A(xdata[249]), .Z(CGFidata[249]));
Q_BUFZP U293 ( .OE(en), .A(xdata[250]), .Z(CGFidata[250]));
Q_BUFZP U294 ( .OE(en), .A(xdata[251]), .Z(CGFidata[251]));
Q_BUFZP U295 ( .OE(en), .A(xdata[252]), .Z(CGFidata[252]));
Q_BUFZP U296 ( .OE(en), .A(xdata[253]), .Z(CGFidata[253]));
Q_BUFZP U297 ( .OE(en), .A(xdata[254]), .Z(CGFidata[254]));
Q_BUFZP U298 ( .OE(en), .A(xdata[255]), .Z(CGFidata[255]));
Q_BUFZP U299 ( .OE(en), .A(xdata[256]), .Z(CGFidata[256]));
Q_BUFZP U300 ( .OE(en), .A(xdata[257]), .Z(CGFidata[257]));
Q_BUFZP U301 ( .OE(en), .A(xdata[258]), .Z(CGFidata[258]));
Q_BUFZP U302 ( .OE(en), .A(xdata[259]), .Z(CGFidata[259]));
Q_BUFZP U303 ( .OE(en), .A(xdata[260]), .Z(CGFidata[260]));
Q_BUFZP U304 ( .OE(en), .A(xdata[261]), .Z(CGFidata[261]));
Q_BUFZP U305 ( .OE(en), .A(xdata[262]), .Z(CGFidata[262]));
Q_BUFZP U306 ( .OE(en), .A(xdata[263]), .Z(CGFidata[263]));
Q_BUFZP U307 ( .OE(en), .A(xdata[264]), .Z(CGFidata[264]));
Q_BUFZP U308 ( .OE(en), .A(xdata[265]), .Z(CGFidata[265]));
Q_BUFZP U309 ( .OE(en), .A(xdata[266]), .Z(CGFidata[266]));
Q_BUFZP U310 ( .OE(en), .A(xdata[267]), .Z(CGFidata[267]));
Q_BUFZP U311 ( .OE(en), .A(xdata[268]), .Z(CGFidata[268]));
Q_BUFZP U312 ( .OE(en), .A(xdata[269]), .Z(CGFidata[269]));
Q_BUFZP U313 ( .OE(en), .A(xdata[270]), .Z(CGFidata[270]));
Q_BUFZP U314 ( .OE(en), .A(xdata[271]), .Z(CGFidata[271]));
Q_BUFZP U315 ( .OE(en), .A(xdata[272]), .Z(CGFidata[272]));
Q_BUFZP U316 ( .OE(en), .A(xdata[273]), .Z(CGFidata[273]));
Q_BUFZP U317 ( .OE(en), .A(xdata[274]), .Z(CGFidata[274]));
Q_BUFZP U318 ( .OE(en), .A(xdata[275]), .Z(CGFidata[275]));
Q_BUFZP U319 ( .OE(en), .A(xdata[276]), .Z(CGFidata[276]));
Q_BUFZP U320 ( .OE(en), .A(xdata[277]), .Z(CGFidata[277]));
Q_BUFZP U321 ( .OE(en), .A(xdata[278]), .Z(CGFidata[278]));
Q_BUFZP U322 ( .OE(en), .A(xdata[279]), .Z(CGFidata[279]));
Q_BUFZP U323 ( .OE(en), .A(xdata[280]), .Z(CGFidata[280]));
Q_BUFZP U324 ( .OE(en), .A(xdata[281]), .Z(CGFidata[281]));
Q_BUFZP U325 ( .OE(en), .A(xdata[282]), .Z(CGFidata[282]));
Q_BUFZP U326 ( .OE(en), .A(xdata[283]), .Z(CGFidata[283]));
Q_BUFZP U327 ( .OE(en), .A(xdata[284]), .Z(CGFidata[284]));
Q_BUFZP U328 ( .OE(en), .A(xdata[285]), .Z(CGFidata[285]));
Q_BUFZP U329 ( .OE(en), .A(xdata[286]), .Z(CGFidata[286]));
Q_BUFZP U330 ( .OE(en), .A(xdata[287]), .Z(CGFidata[287]));
Q_BUFZP U331 ( .OE(en), .A(xdata[288]), .Z(CGFidata[288]));
Q_BUFZP U332 ( .OE(en), .A(xdata[289]), .Z(CGFidata[289]));
Q_BUFZP U333 ( .OE(en), .A(xdata[290]), .Z(CGFidata[290]));
Q_BUFZP U334 ( .OE(en), .A(xdata[291]), .Z(CGFidata[291]));
Q_BUFZP U335 ( .OE(en), .A(xdata[292]), .Z(CGFidata[292]));
Q_BUFZP U336 ( .OE(en), .A(xdata[293]), .Z(CGFidata[293]));
Q_BUFZP U337 ( .OE(en), .A(xdata[294]), .Z(CGFidata[294]));
Q_BUFZP U338 ( .OE(en), .A(xdata[295]), .Z(CGFidata[295]));
Q_BUFZP U339 ( .OE(en), .A(xdata[296]), .Z(CGFidata[296]));
Q_BUFZP U340 ( .OE(en), .A(xdata[297]), .Z(CGFidata[297]));
Q_BUFZP U341 ( .OE(en), .A(xdata[298]), .Z(CGFidata[298]));
Q_BUFZP U342 ( .OE(en), .A(xdata[299]), .Z(CGFidata[299]));
Q_BUFZP U343 ( .OE(en), .A(xdata[300]), .Z(CGFidata[300]));
Q_BUFZP U344 ( .OE(en), .A(xdata[301]), .Z(CGFidata[301]));
Q_BUFZP U345 ( .OE(en), .A(xdata[302]), .Z(CGFidata[302]));
Q_BUFZP U346 ( .OE(en), .A(xdata[303]), .Z(CGFidata[303]));
Q_BUFZP U347 ( .OE(en), .A(xdata[304]), .Z(CGFidata[304]));
Q_BUFZP U348 ( .OE(en), .A(xdata[305]), .Z(CGFidata[305]));
Q_BUFZP U349 ( .OE(en), .A(xdata[306]), .Z(CGFidata[306]));
Q_BUFZP U350 ( .OE(en), .A(xdata[307]), .Z(CGFidata[307]));
Q_BUFZP U351 ( .OE(en), .A(xdata[308]), .Z(CGFidata[308]));
Q_BUFZP U352 ( .OE(en), .A(xdata[309]), .Z(CGFidata[309]));
Q_BUFZP U353 ( .OE(en), .A(xdata[310]), .Z(CGFidata[310]));
Q_BUFZP U354 ( .OE(en), .A(xdata[311]), .Z(CGFidata[311]));
Q_BUFZP U355 ( .OE(en), .A(xdata[312]), .Z(CGFidata[312]));
Q_BUFZP U356 ( .OE(en), .A(xdata[313]), .Z(CGFidata[313]));
Q_BUFZP U357 ( .OE(en), .A(xdata[314]), .Z(CGFidata[314]));
Q_BUFZP U358 ( .OE(en), .A(xdata[315]), .Z(CGFidata[315]));
Q_BUFZP U359 ( .OE(en), .A(xdata[316]), .Z(CGFidata[316]));
Q_BUFZP U360 ( .OE(en), .A(xdata[317]), .Z(CGFidata[317]));
Q_BUFZP U361 ( .OE(en), .A(xdata[318]), .Z(CGFidata[318]));
Q_BUFZP U362 ( .OE(en), .A(xdata[319]), .Z(CGFidata[319]));
Q_BUFZP U363 ( .OE(en), .A(xdata[320]), .Z(CGFidata[320]));
Q_BUFZP U364 ( .OE(en), .A(xdata[321]), .Z(CGFidata[321]));
Q_BUFZP U365 ( .OE(en), .A(xdata[322]), .Z(CGFidata[322]));
Q_BUFZP U366 ( .OE(en), .A(xdata[323]), .Z(CGFidata[323]));
Q_BUFZP U367 ( .OE(en), .A(xdata[324]), .Z(CGFidata[324]));
Q_BUFZP U368 ( .OE(en), .A(xdata[325]), .Z(CGFidata[325]));
Q_BUFZP U369 ( .OE(en), .A(xdata[326]), .Z(CGFidata[326]));
Q_BUFZP U370 ( .OE(en), .A(xdata[327]), .Z(CGFidata[327]));
Q_BUFZP U371 ( .OE(en), .A(xdata[328]), .Z(CGFidata[328]));
Q_BUFZP U372 ( .OE(en), .A(xdata[329]), .Z(CGFidata[329]));
Q_BUFZP U373 ( .OE(en), .A(xdata[330]), .Z(CGFidata[330]));
Q_BUFZP U374 ( .OE(en), .A(xdata[331]), .Z(CGFidata[331]));
Q_BUFZP U375 ( .OE(en), .A(xdata[332]), .Z(CGFidata[332]));
Q_BUFZP U376 ( .OE(en), .A(xdata[333]), .Z(CGFidata[333]));
Q_BUFZP U377 ( .OE(en), .A(xdata[334]), .Z(CGFidata[334]));
Q_BUFZP U378 ( .OE(en), .A(xdata[335]), .Z(CGFidata[335]));
Q_BUFZP U379 ( .OE(en), .A(xdata[336]), .Z(CGFidata[336]));
Q_BUFZP U380 ( .OE(en), .A(xdata[337]), .Z(CGFidata[337]));
Q_BUFZP U381 ( .OE(en), .A(xdata[338]), .Z(CGFidata[338]));
Q_BUFZP U382 ( .OE(en), .A(xdata[339]), .Z(CGFidata[339]));
Q_BUFZP U383 ( .OE(en), .A(xdata[340]), .Z(CGFidata[340]));
Q_BUFZP U384 ( .OE(en), .A(xdata[341]), .Z(CGFidata[341]));
Q_BUFZP U385 ( .OE(en), .A(xdata[342]), .Z(CGFidata[342]));
Q_BUFZP U386 ( .OE(en), .A(xdata[343]), .Z(CGFidata[343]));
Q_BUFZP U387 ( .OE(en), .A(xdata[344]), .Z(CGFidata[344]));
Q_BUFZP U388 ( .OE(en), .A(xdata[345]), .Z(CGFidata[345]));
Q_BUFZP U389 ( .OE(en), .A(xdata[346]), .Z(CGFidata[346]));
Q_BUFZP U390 ( .OE(en), .A(xdata[347]), .Z(CGFidata[347]));
Q_BUFZP U391 ( .OE(en), .A(xdata[348]), .Z(CGFidata[348]));
Q_BUFZP U392 ( .OE(en), .A(xdata[349]), .Z(CGFidata[349]));
Q_BUFZP U393 ( .OE(en), .A(xdata[350]), .Z(CGFidata[350]));
Q_BUFZP U394 ( .OE(en), .A(xdata[351]), .Z(CGFidata[351]));
Q_BUFZP U395 ( .OE(en), .A(xdata[352]), .Z(CGFidata[352]));
Q_BUFZP U396 ( .OE(en), .A(xdata[353]), .Z(CGFidata[353]));
Q_BUFZP U397 ( .OE(en), .A(xdata[354]), .Z(CGFidata[354]));
Q_BUFZP U398 ( .OE(en), .A(xdata[355]), .Z(CGFidata[355]));
Q_BUFZP U399 ( .OE(en), .A(xdata[356]), .Z(CGFidata[356]));
Q_BUFZP U400 ( .OE(en), .A(xdata[357]), .Z(CGFidata[357]));
Q_BUFZP U401 ( .OE(en), .A(xdata[358]), .Z(CGFidata[358]));
Q_BUFZP U402 ( .OE(en), .A(xdata[359]), .Z(CGFidata[359]));
Q_BUFZP U403 ( .OE(en), .A(xdata[360]), .Z(CGFidata[360]));
Q_BUFZP U404 ( .OE(en), .A(xdata[361]), .Z(CGFidata[361]));
Q_BUFZP U405 ( .OE(en), .A(xdata[362]), .Z(CGFidata[362]));
Q_BUFZP U406 ( .OE(en), .A(xdata[363]), .Z(CGFidata[363]));
Q_BUFZP U407 ( .OE(en), .A(xdata[364]), .Z(CGFidata[364]));
Q_BUFZP U408 ( .OE(en), .A(xdata[365]), .Z(CGFidata[365]));
Q_BUFZP U409 ( .OE(en), .A(xdata[366]), .Z(CGFidata[366]));
Q_BUFZP U410 ( .OE(en), .A(xdata[367]), .Z(CGFidata[367]));
Q_BUFZP U411 ( .OE(en), .A(xdata[368]), .Z(CGFidata[368]));
Q_BUFZP U412 ( .OE(en), .A(xdata[369]), .Z(CGFidata[369]));
Q_BUFZP U413 ( .OE(en), .A(xdata[370]), .Z(CGFidata[370]));
Q_BUFZP U414 ( .OE(en), .A(xdata[371]), .Z(CGFidata[371]));
Q_BUFZP U415 ( .OE(en), .A(xdata[372]), .Z(CGFidata[372]));
Q_BUFZP U416 ( .OE(en), .A(xdata[373]), .Z(CGFidata[373]));
Q_BUFZP U417 ( .OE(en), .A(xdata[374]), .Z(CGFidata[374]));
Q_BUFZP U418 ( .OE(en), .A(xdata[375]), .Z(CGFidata[375]));
Q_BUFZP U419 ( .OE(en), .A(xdata[376]), .Z(CGFidata[376]));
Q_BUFZP U420 ( .OE(en), .A(xdata[377]), .Z(CGFidata[377]));
Q_BUFZP U421 ( .OE(en), .A(xdata[378]), .Z(CGFidata[378]));
Q_BUFZP U422 ( .OE(en), .A(xdata[379]), .Z(CGFidata[379]));
Q_BUFZP U423 ( .OE(en), .A(xdata[380]), .Z(CGFidata[380]));
Q_BUFZP U424 ( .OE(en), .A(xdata[381]), .Z(CGFidata[381]));
Q_BUFZP U425 ( .OE(en), .A(xdata[382]), .Z(CGFidata[382]));
Q_BUFZP U426 ( .OE(en), .A(xdata[383]), .Z(CGFidata[383]));
Q_BUFZP U427 ( .OE(en), .A(xdata[384]), .Z(CGFidata[384]));
Q_BUFZP U428 ( .OE(en), .A(xdata[385]), .Z(CGFidata[385]));
Q_BUFZP U429 ( .OE(en), .A(xdata[386]), .Z(CGFidata[386]));
Q_BUFZP U430 ( .OE(en), .A(xdata[387]), .Z(CGFidata[387]));
Q_BUFZP U431 ( .OE(en), .A(xdata[388]), .Z(CGFidata[388]));
Q_BUFZP U432 ( .OE(en), .A(xdata[389]), .Z(CGFidata[389]));
Q_BUFZP U433 ( .OE(en), .A(xdata[390]), .Z(CGFidata[390]));
Q_BUFZP U434 ( .OE(en), .A(xdata[391]), .Z(CGFidata[391]));
Q_BUFZP U435 ( .OE(en), .A(xdata[392]), .Z(CGFidata[392]));
Q_BUFZP U436 ( .OE(en), .A(xdata[393]), .Z(CGFidata[393]));
Q_BUFZP U437 ( .OE(en), .A(xdata[394]), .Z(CGFidata[394]));
Q_BUFZP U438 ( .OE(en), .A(xdata[395]), .Z(CGFidata[395]));
Q_BUFZP U439 ( .OE(en), .A(xdata[396]), .Z(CGFidata[396]));
Q_BUFZP U440 ( .OE(en), .A(xdata[397]), .Z(CGFidata[397]));
Q_BUFZP U441 ( .OE(en), .A(xdata[398]), .Z(CGFidata[398]));
Q_BUFZP U442 ( .OE(en), .A(xdata[399]), .Z(CGFidata[399]));
Q_BUFZP U443 ( .OE(en), .A(xdata[400]), .Z(CGFidata[400]));
Q_BUFZP U444 ( .OE(en), .A(xdata[401]), .Z(CGFidata[401]));
Q_BUFZP U445 ( .OE(en), .A(xdata[402]), .Z(CGFidata[402]));
Q_BUFZP U446 ( .OE(en), .A(xdata[403]), .Z(CGFidata[403]));
Q_BUFZP U447 ( .OE(en), .A(xdata[404]), .Z(CGFidata[404]));
Q_BUFZP U448 ( .OE(en), .A(xdata[405]), .Z(CGFidata[405]));
Q_BUFZP U449 ( .OE(en), .A(xdata[406]), .Z(CGFidata[406]));
Q_BUFZP U450 ( .OE(en), .A(xdata[407]), .Z(CGFidata[407]));
Q_BUFZP U451 ( .OE(en), .A(xdata[408]), .Z(CGFidata[408]));
Q_BUFZP U452 ( .OE(en), .A(xdata[409]), .Z(CGFidata[409]));
Q_BUFZP U453 ( .OE(en), .A(xdata[410]), .Z(CGFidata[410]));
Q_BUFZP U454 ( .OE(en), .A(xdata[411]), .Z(CGFidata[411]));
Q_BUFZP U455 ( .OE(en), .A(xdata[412]), .Z(CGFidata[412]));
Q_BUFZP U456 ( .OE(en), .A(xdata[413]), .Z(CGFidata[413]));
Q_BUFZP U457 ( .OE(en), .A(xdata[414]), .Z(CGFidata[414]));
Q_BUFZP U458 ( .OE(en), .A(xdata[415]), .Z(CGFidata[415]));
Q_BUFZP U459 ( .OE(en), .A(xdata[416]), .Z(CGFidata[416]));
Q_BUFZP U460 ( .OE(en), .A(xdata[417]), .Z(CGFidata[417]));
Q_BUFZP U461 ( .OE(en), .A(xdata[418]), .Z(CGFidata[418]));
Q_BUFZP U462 ( .OE(en), .A(xdata[419]), .Z(CGFidata[419]));
Q_BUFZP U463 ( .OE(en), .A(xdata[420]), .Z(CGFidata[420]));
Q_BUFZP U464 ( .OE(en), .A(xdata[421]), .Z(CGFidata[421]));
Q_BUFZP U465 ( .OE(en), .A(xdata[422]), .Z(CGFidata[422]));
Q_BUFZP U466 ( .OE(en), .A(xdata[423]), .Z(CGFidata[423]));
Q_BUFZP U467 ( .OE(en), .A(xdata[424]), .Z(CGFidata[424]));
Q_BUFZP U468 ( .OE(en), .A(xdata[425]), .Z(CGFidata[425]));
Q_BUFZP U469 ( .OE(en), .A(xdata[426]), .Z(CGFidata[426]));
Q_BUFZP U470 ( .OE(en), .A(xdata[427]), .Z(CGFidata[427]));
Q_BUFZP U471 ( .OE(en), .A(xdata[428]), .Z(CGFidata[428]));
Q_BUFZP U472 ( .OE(en), .A(xdata[429]), .Z(CGFidata[429]));
Q_BUFZP U473 ( .OE(en), .A(xdata[430]), .Z(CGFidata[430]));
Q_BUFZP U474 ( .OE(en), .A(xdata[431]), .Z(CGFidata[431]));
Q_BUFZP U475 ( .OE(en), .A(xdata[432]), .Z(CGFidata[432]));
Q_BUFZP U476 ( .OE(en), .A(xdata[433]), .Z(CGFidata[433]));
Q_BUFZP U477 ( .OE(en), .A(xdata[434]), .Z(CGFidata[434]));
Q_BUFZP U478 ( .OE(en), .A(xdata[435]), .Z(CGFidata[435]));
Q_BUFZP U479 ( .OE(en), .A(xdata[436]), .Z(CGFidata[436]));
Q_BUFZP U480 ( .OE(en), .A(xdata[437]), .Z(CGFidata[437]));
Q_BUFZP U481 ( .OE(en), .A(xdata[438]), .Z(CGFidata[438]));
Q_BUFZP U482 ( .OE(en), .A(xdata[439]), .Z(CGFidata[439]));
Q_BUFZP U483 ( .OE(en), .A(xdata[440]), .Z(CGFidata[440]));
Q_BUFZP U484 ( .OE(en), .A(xdata[441]), .Z(CGFidata[441]));
Q_BUFZP U485 ( .OE(en), .A(xdata[442]), .Z(CGFidata[442]));
Q_BUFZP U486 ( .OE(en), .A(xdata[443]), .Z(CGFidata[443]));
Q_BUFZP U487 ( .OE(en), .A(xdata[444]), .Z(CGFidata[444]));
Q_BUFZP U488 ( .OE(en), .A(xdata[445]), .Z(CGFidata[445]));
Q_BUFZP U489 ( .OE(en), .A(xdata[446]), .Z(CGFidata[446]));
Q_BUFZP U490 ( .OE(en), .A(xdata[447]), .Z(CGFidata[447]));
Q_BUFZP U491 ( .OE(en), .A(xdata[448]), .Z(CGFidata[448]));
Q_BUFZP U492 ( .OE(en), .A(xdata[449]), .Z(CGFidata[449]));
Q_BUFZP U493 ( .OE(en), .A(xdata[450]), .Z(CGFidata[450]));
Q_BUFZP U494 ( .OE(en), .A(xdata[451]), .Z(CGFidata[451]));
Q_BUFZP U495 ( .OE(en), .A(xdata[452]), .Z(CGFidata[452]));
Q_BUFZP U496 ( .OE(en), .A(xdata[453]), .Z(CGFidata[453]));
Q_BUFZP U497 ( .OE(en), .A(xdata[454]), .Z(CGFidata[454]));
Q_BUFZP U498 ( .OE(en), .A(xdata[455]), .Z(CGFidata[455]));
Q_BUFZP U499 ( .OE(en), .A(xdata[456]), .Z(CGFidata[456]));
Q_BUFZP U500 ( .OE(en), .A(xdata[457]), .Z(CGFidata[457]));
Q_BUFZP U501 ( .OE(en), .A(xdata[458]), .Z(CGFidata[458]));
Q_BUFZP U502 ( .OE(en), .A(xdata[459]), .Z(CGFidata[459]));
Q_BUFZP U503 ( .OE(en), .A(xdata[460]), .Z(CGFidata[460]));
Q_BUFZP U504 ( .OE(en), .A(xdata[461]), .Z(CGFidata[461]));
Q_BUFZP U505 ( .OE(en), .A(xdata[462]), .Z(CGFidata[462]));
Q_BUFZP U506 ( .OE(en), .A(xdata[463]), .Z(CGFidata[463]));
Q_BUFZP U507 ( .OE(en), .A(xdata[464]), .Z(CGFidata[464]));
Q_BUFZP U508 ( .OE(en), .A(xdata[465]), .Z(CGFidata[465]));
Q_BUFZP U509 ( .OE(en), .A(xdata[466]), .Z(CGFidata[466]));
Q_BUFZP U510 ( .OE(en), .A(xdata[467]), .Z(CGFidata[467]));
Q_BUFZP U511 ( .OE(en), .A(xdata[468]), .Z(CGFidata[468]));
Q_BUFZP U512 ( .OE(en), .A(xdata[469]), .Z(CGFidata[469]));
Q_BUFZP U513 ( .OE(en), .A(xdata[470]), .Z(CGFidata[470]));
Q_BUFZP U514 ( .OE(en), .A(xdata[471]), .Z(CGFidata[471]));
Q_BUFZP U515 ( .OE(en), .A(xdata[472]), .Z(CGFidata[472]));
Q_BUFZP U516 ( .OE(en), .A(xdata[473]), .Z(CGFidata[473]));
Q_BUFZP U517 ( .OE(en), .A(xdata[474]), .Z(CGFidata[474]));
Q_BUFZP U518 ( .OE(en), .A(xdata[475]), .Z(CGFidata[475]));
Q_BUFZP U519 ( .OE(en), .A(xdata[476]), .Z(CGFidata[476]));
Q_BUFZP U520 ( .OE(en), .A(xdata[477]), .Z(CGFidata[477]));
Q_BUFZP U521 ( .OE(en), .A(xdata[478]), .Z(CGFidata[478]));
Q_BUFZP U522 ( .OE(en), .A(xdata[479]), .Z(CGFidata[479]));
Q_BUFZP U523 ( .OE(en), .A(xdata[480]), .Z(CGFidata[480]));
Q_BUFZP U524 ( .OE(en), .A(xdata[481]), .Z(CGFidata[481]));
Q_BUFZP U525 ( .OE(en), .A(xdata[482]), .Z(CGFidata[482]));
Q_BUFZP U526 ( .OE(en), .A(xdata[483]), .Z(CGFidata[483]));
Q_BUFZP U527 ( .OE(en), .A(xdata[484]), .Z(CGFidata[484]));
Q_BUFZP U528 ( .OE(en), .A(xdata[485]), .Z(CGFidata[485]));
Q_BUFZP U529 ( .OE(en), .A(xdata[486]), .Z(CGFidata[486]));
Q_BUFZP U530 ( .OE(en), .A(xdata[487]), .Z(CGFidata[487]));
Q_BUFZP U531 ( .OE(en), .A(xdata[488]), .Z(CGFidata[488]));
Q_BUFZP U532 ( .OE(en), .A(xdata[489]), .Z(CGFidata[489]));
Q_BUFZP U533 ( .OE(en), .A(xdata[490]), .Z(CGFidata[490]));
Q_BUFZP U534 ( .OE(en), .A(xdata[491]), .Z(CGFidata[491]));
Q_BUFZP U535 ( .OE(en), .A(xdata[492]), .Z(CGFidata[492]));
Q_BUFZP U536 ( .OE(en), .A(xdata[493]), .Z(CGFidata[493]));
Q_BUFZP U537 ( .OE(en), .A(xdata[494]), .Z(CGFidata[494]));
Q_BUFZP U538 ( .OE(en), .A(xdata[495]), .Z(CGFidata[495]));
Q_BUFZP U539 ( .OE(en), .A(xdata[496]), .Z(CGFidata[496]));
Q_BUFZP U540 ( .OE(en), .A(xdata[497]), .Z(CGFidata[497]));
Q_BUFZP U541 ( .OE(en), .A(xdata[498]), .Z(CGFidata[498]));
Q_BUFZP U542 ( .OE(en), .A(xdata[499]), .Z(CGFidata[499]));
Q_BUFZP U543 ( .OE(en), .A(xdata[500]), .Z(CGFidata[500]));
Q_BUFZP U544 ( .OE(en), .A(xdata[501]), .Z(CGFidata[501]));
Q_BUFZP U545 ( .OE(en), .A(xdata[502]), .Z(CGFidata[502]));
Q_BUFZP U546 ( .OE(en), .A(xdata[503]), .Z(CGFidata[503]));
Q_BUFZP U547 ( .OE(en), .A(xdata[504]), .Z(CGFidata[504]));
Q_BUFZP U548 ( .OE(en), .A(xdata[505]), .Z(CGFidata[505]));
Q_BUFZP U549 ( .OE(en), .A(xdata[506]), .Z(CGFidata[506]));
Q_BUFZP U550 ( .OE(en), .A(xdata[507]), .Z(CGFidata[507]));
Q_BUFZP U551 ( .OE(en), .A(xdata[508]), .Z(CGFidata[508]));
Q_BUFZP U552 ( .OE(en), .A(xdata[509]), .Z(CGFidata[509]));
Q_BUFZP U553 ( .OE(en), .A(xdata[510]), .Z(CGFidata[510]));
Q_BUFZP U554 ( .OE(en), .A(xdata[511]), .Z(CGFidata[511]));
Q_AO21 U555 ( .A0(sel[0]), .A1(odata[0]), .B0(n7), .Z(xdata[0]));
Q_AO21 U556 ( .A0(sel[0]), .A1(odata[1]), .B0(n8), .Z(xdata[1]));
Q_AO21 U557 ( .A0(sel[0]), .A1(odata[2]), .B0(n9), .Z(xdata[2]));
Q_AO21 U558 ( .A0(sel[0]), .A1(odata[3]), .B0(n10), .Z(xdata[3]));
Q_AO21 U559 ( .A0(sel[0]), .A1(odata[4]), .B0(n11), .Z(xdata[4]));
Q_AO21 U560 ( .A0(sel[0]), .A1(odata[5]), .B0(n12), .Z(xdata[5]));
Q_AO21 U561 ( .A0(sel[0]), .A1(odata[6]), .B0(n13), .Z(xdata[6]));
Q_AO21 U562 ( .A0(sel[0]), .A1(odata[7]), .B0(n14), .Z(xdata[7]));
Q_AO21 U563 ( .A0(sel[0]), .A1(odata[8]), .B0(n15), .Z(xdata[8]));
Q_AO21 U564 ( .A0(sel[0]), .A1(odata[9]), .B0(n16), .Z(xdata[9]));
Q_AO21 U565 ( .A0(sel[0]), .A1(odata[10]), .B0(n17), .Z(xdata[10]));
Q_AO21 U566 ( .A0(sel[0]), .A1(odata[11]), .B0(n18), .Z(xdata[11]));
Q_AO21 U567 ( .A0(sel[0]), .A1(odata[12]), .B0(n19), .Z(xdata[12]));
Q_AO21 U568 ( .A0(sel[0]), .A1(odata[13]), .B0(n20), .Z(xdata[13]));
Q_AO21 U569 ( .A0(sel[0]), .A1(odata[14]), .B0(n21), .Z(xdata[14]));
Q_AO21 U570 ( .A0(sel[0]), .A1(odata[15]), .B0(n22), .Z(xdata[15]));
Q_AO21 U571 ( .A0(sel[0]), .A1(odata[16]), .B0(n23), .Z(xdata[16]));
Q_AO21 U572 ( .A0(sel[0]), .A1(odata[17]), .B0(n24), .Z(xdata[17]));
Q_AO21 U573 ( .A0(sel[0]), .A1(odata[18]), .B0(n25), .Z(xdata[18]));
Q_AO21 U574 ( .A0(sel[0]), .A1(odata[19]), .B0(n26), .Z(xdata[19]));
Q_AO21 U575 ( .A0(sel[0]), .A1(odata[20]), .B0(n27), .Z(xdata[20]));
Q_AO21 U576 ( .A0(sel[0]), .A1(odata[21]), .B0(n28), .Z(xdata[21]));
Q_AO21 U577 ( .A0(sel[0]), .A1(odata[22]), .B0(n29), .Z(xdata[22]));
Q_AO21 U578 ( .A0(sel[0]), .A1(odata[23]), .B0(n30), .Z(xdata[23]));
Q_AO21 U579 ( .A0(sel[0]), .A1(odata[24]), .B0(n31), .Z(xdata[24]));
Q_AO21 U580 ( .A0(sel[0]), .A1(odata[25]), .B0(n32), .Z(xdata[25]));
Q_AO21 U581 ( .A0(sel[0]), .A1(odata[26]), .B0(n33), .Z(xdata[26]));
Q_AO21 U582 ( .A0(sel[0]), .A1(odata[27]), .B0(n34), .Z(xdata[27]));
Q_AO21 U583 ( .A0(sel[0]), .A1(odata[28]), .B0(n35), .Z(xdata[28]));
Q_AO21 U584 ( .A0(sel[0]), .A1(odata[29]), .B0(n36), .Z(xdata[29]));
Q_AO21 U585 ( .A0(sel[0]), .A1(odata[30]), .B0(n37), .Z(xdata[30]));
Q_AO21 U586 ( .A0(sel[0]), .A1(odata[31]), .B0(n38), .Z(xdata[31]));
Q_AO21 U587 ( .A0(sel[0]), .A1(odata[32]), .B0(n39), .Z(xdata[32]));
Q_AO21 U588 ( .A0(sel[0]), .A1(odata[33]), .B0(n40), .Z(xdata[33]));
Q_AO21 U589 ( .A0(sel[0]), .A1(odata[34]), .B0(n41), .Z(xdata[34]));
Q_AO21 U590 ( .A0(sel[0]), .A1(odata[35]), .B0(n42), .Z(xdata[35]));
Q_AO21 U591 ( .A0(sel[0]), .A1(odata[36]), .B0(n43), .Z(xdata[36]));
Q_AO21 U592 ( .A0(sel[0]), .A1(odata[37]), .B0(n44), .Z(xdata[37]));
Q_AO21 U593 ( .A0(sel[0]), .A1(odata[38]), .B0(n45), .Z(xdata[38]));
Q_AO21 U594 ( .A0(sel[0]), .A1(odata[39]), .B0(n46), .Z(xdata[39]));
Q_AO21 U595 ( .A0(sel[0]), .A1(odata[40]), .B0(n47), .Z(xdata[40]));
Q_AO21 U596 ( .A0(sel[0]), .A1(odata[41]), .B0(n48), .Z(xdata[41]));
Q_AO21 U597 ( .A0(sel[0]), .A1(odata[42]), .B0(n49), .Z(xdata[42]));
Q_AO21 U598 ( .A0(sel[0]), .A1(odata[43]), .B0(n50), .Z(xdata[43]));
Q_AO21 U599 ( .A0(sel[0]), .A1(odata[44]), .B0(n51), .Z(xdata[44]));
Q_AO21 U600 ( .A0(sel[0]), .A1(odata[45]), .B0(n52), .Z(xdata[45]));
Q_AO21 U601 ( .A0(sel[0]), .A1(odata[46]), .B0(n53), .Z(xdata[46]));
Q_AO21 U602 ( .A0(sel[0]), .A1(odata[47]), .B0(n54), .Z(xdata[47]));
Q_AN02 U603 ( .A0(sel[0]), .A1(odata[48]), .Z(xdata[48]));
Q_AN02 U604 ( .A0(sel[0]), .A1(odata[49]), .Z(xdata[49]));
Q_AN02 U605 ( .A0(sel[0]), .A1(odata[50]), .Z(xdata[50]));
Q_AN02 U606 ( .A0(sel[0]), .A1(odata[51]), .Z(xdata[51]));
Q_AN02 U607 ( .A0(sel[0]), .A1(odata[52]), .Z(xdata[52]));
Q_AN02 U608 ( .A0(sel[0]), .A1(odata[53]), .Z(xdata[53]));
Q_AN02 U609 ( .A0(sel[0]), .A1(odata[54]), .Z(xdata[54]));
Q_AN02 U610 ( .A0(sel[0]), .A1(odata[55]), .Z(xdata[55]));
Q_AN02 U611 ( .A0(sel[0]), .A1(odata[56]), .Z(xdata[56]));
Q_AN02 U612 ( .A0(sel[0]), .A1(odata[57]), .Z(xdata[57]));
Q_AN02 U613 ( .A0(sel[0]), .A1(odata[58]), .Z(xdata[58]));
Q_AN02 U614 ( .A0(sel[0]), .A1(odata[59]), .Z(xdata[59]));
Q_AN02 U615 ( .A0(sel[0]), .A1(odata[60]), .Z(xdata[60]));
Q_AN02 U616 ( .A0(sel[0]), .A1(odata[61]), .Z(xdata[61]));
Q_AN02 U617 ( .A0(sel[0]), .A1(odata[62]), .Z(xdata[62]));
Q_AN02 U618 ( .A0(sel[0]), .A1(odata[63]), .Z(xdata[63]));
Q_AN02 U619 ( .A0(sel[0]), .A1(odata[64]), .Z(xdata[64]));
Q_AN02 U620 ( .A0(sel[0]), .A1(odata[65]), .Z(xdata[65]));
Q_AN02 U621 ( .A0(sel[0]), .A1(odata[66]), .Z(xdata[66]));
Q_AN02 U622 ( .A0(sel[0]), .A1(odata[67]), .Z(xdata[67]));
Q_AN02 U623 ( .A0(sel[0]), .A1(odata[68]), .Z(xdata[68]));
Q_AN02 U624 ( .A0(sel[0]), .A1(odata[69]), .Z(xdata[69]));
Q_AN02 U625 ( .A0(sel[0]), .A1(odata[70]), .Z(xdata[70]));
Q_AN02 U626 ( .A0(sel[0]), .A1(odata[71]), .Z(xdata[71]));
Q_AN02 U627 ( .A0(sel[0]), .A1(odata[72]), .Z(xdata[72]));
Q_AN02 U628 ( .A0(sel[0]), .A1(odata[73]), .Z(xdata[73]));
Q_AN02 U629 ( .A0(sel[0]), .A1(odata[74]), .Z(xdata[74]));
Q_AN02 U630 ( .A0(sel[0]), .A1(odata[75]), .Z(xdata[75]));
Q_AN02 U631 ( .A0(sel[0]), .A1(odata[76]), .Z(xdata[76]));
Q_AN02 U632 ( .A0(sel[0]), .A1(odata[77]), .Z(xdata[77]));
Q_AN02 U633 ( .A0(sel[0]), .A1(odata[78]), .Z(xdata[78]));
Q_AN02 U634 ( .A0(sel[0]), .A1(odata[79]), .Z(xdata[79]));
Q_AN02 U635 ( .A0(sel[0]), .A1(odata[80]), .Z(xdata[80]));
Q_AN02 U636 ( .A0(sel[0]), .A1(odata[81]), .Z(xdata[81]));
Q_AN02 U637 ( .A0(sel[0]), .A1(odata[82]), .Z(xdata[82]));
Q_AN02 U638 ( .A0(sel[0]), .A1(odata[83]), .Z(xdata[83]));
Q_AN02 U639 ( .A0(sel[0]), .A1(odata[84]), .Z(xdata[84]));
Q_AN02 U640 ( .A0(sel[0]), .A1(odata[85]), .Z(xdata[85]));
Q_AN02 U641 ( .A0(sel[0]), .A1(odata[86]), .Z(xdata[86]));
Q_AN02 U642 ( .A0(sel[0]), .A1(odata[87]), .Z(xdata[87]));
Q_AN02 U643 ( .A0(sel[0]), .A1(odata[88]), .Z(xdata[88]));
Q_AN02 U644 ( .A0(sel[0]), .A1(odata[89]), .Z(xdata[89]));
Q_AN02 U645 ( .A0(sel[0]), .A1(odata[90]), .Z(xdata[90]));
Q_AN02 U646 ( .A0(sel[0]), .A1(odata[91]), .Z(xdata[91]));
Q_AN02 U647 ( .A0(sel[0]), .A1(odata[92]), .Z(xdata[92]));
Q_AN02 U648 ( .A0(sel[0]), .A1(odata[93]), .Z(xdata[93]));
Q_AN02 U649 ( .A0(sel[0]), .A1(odata[94]), .Z(xdata[94]));
Q_AN02 U650 ( .A0(sel[0]), .A1(odata[95]), .Z(xdata[95]));
Q_AN02 U651 ( .A0(sel[0]), .A1(odata[96]), .Z(xdata[96]));
Q_AN02 U652 ( .A0(sel[0]), .A1(odata[97]), .Z(xdata[97]));
Q_AN02 U653 ( .A0(sel[0]), .A1(odata[98]), .Z(xdata[98]));
Q_AN02 U654 ( .A0(sel[0]), .A1(odata[99]), .Z(xdata[99]));
Q_AN02 U655 ( .A0(sel[0]), .A1(odata[100]), .Z(xdata[100]));
Q_AN02 U656 ( .A0(sel[0]), .A1(odata[101]), .Z(xdata[101]));
Q_AN02 U657 ( .A0(sel[0]), .A1(odata[102]), .Z(xdata[102]));
Q_AN02 U658 ( .A0(sel[0]), .A1(odata[103]), .Z(xdata[103]));
Q_AN02 U659 ( .A0(sel[0]), .A1(odata[104]), .Z(xdata[104]));
Q_AN02 U660 ( .A0(sel[0]), .A1(odata[105]), .Z(xdata[105]));
Q_AN02 U661 ( .A0(sel[0]), .A1(odata[106]), .Z(xdata[106]));
Q_AN02 U662 ( .A0(sel[0]), .A1(odata[107]), .Z(xdata[107]));
Q_AN02 U663 ( .A0(sel[0]), .A1(odata[108]), .Z(xdata[108]));
Q_AN02 U664 ( .A0(sel[0]), .A1(odata[109]), .Z(xdata[109]));
Q_AN02 U665 ( .A0(sel[0]), .A1(odata[110]), .Z(xdata[110]));
Q_AN02 U666 ( .A0(sel[0]), .A1(odata[111]), .Z(xdata[111]));
Q_AN02 U667 ( .A0(sel[0]), .A1(odata[112]), .Z(xdata[112]));
Q_AN02 U668 ( .A0(sel[0]), .A1(odata[113]), .Z(xdata[113]));
Q_AN02 U669 ( .A0(sel[0]), .A1(odata[114]), .Z(xdata[114]));
Q_AN02 U670 ( .A0(sel[0]), .A1(odata[115]), .Z(xdata[115]));
Q_AN02 U671 ( .A0(sel[0]), .A1(odata[116]), .Z(xdata[116]));
Q_AN02 U672 ( .A0(sel[0]), .A1(odata[117]), .Z(xdata[117]));
Q_AN02 U673 ( .A0(sel[0]), .A1(odata[118]), .Z(xdata[118]));
Q_AN02 U674 ( .A0(sel[0]), .A1(odata[119]), .Z(xdata[119]));
Q_AN02 U675 ( .A0(sel[0]), .A1(odata[120]), .Z(xdata[120]));
Q_AN02 U676 ( .A0(sel[0]), .A1(odata[121]), .Z(xdata[121]));
Q_AN02 U677 ( .A0(sel[0]), .A1(odata[122]), .Z(xdata[122]));
Q_AN02 U678 ( .A0(sel[0]), .A1(odata[123]), .Z(xdata[123]));
Q_AN02 U679 ( .A0(sel[0]), .A1(odata[124]), .Z(xdata[124]));
Q_AN02 U680 ( .A0(sel[0]), .A1(odata[125]), .Z(xdata[125]));
Q_AN02 U681 ( .A0(sel[0]), .A1(odata[126]), .Z(xdata[126]));
Q_AN02 U682 ( .A0(sel[0]), .A1(odata[127]), .Z(xdata[127]));
Q_AN02 U683 ( .A0(sel[0]), .A1(odata[128]), .Z(xdata[128]));
Q_AN02 U684 ( .A0(sel[0]), .A1(odata[129]), .Z(xdata[129]));
Q_AN02 U685 ( .A0(sel[0]), .A1(odata[130]), .Z(xdata[130]));
Q_AN02 U686 ( .A0(sel[0]), .A1(odata[131]), .Z(xdata[131]));
Q_AN02 U687 ( .A0(sel[0]), .A1(odata[132]), .Z(xdata[132]));
Q_AN02 U688 ( .A0(sel[0]), .A1(odata[133]), .Z(xdata[133]));
Q_AN02 U689 ( .A0(sel[0]), .A1(odata[134]), .Z(xdata[134]));
Q_AN02 U690 ( .A0(sel[0]), .A1(odata[135]), .Z(xdata[135]));
Q_AN02 U691 ( .A0(sel[0]), .A1(odata[136]), .Z(xdata[136]));
Q_AN02 U692 ( .A0(sel[0]), .A1(odata[137]), .Z(xdata[137]));
Q_AN02 U693 ( .A0(sel[0]), .A1(odata[138]), .Z(xdata[138]));
Q_AN02 U694 ( .A0(sel[0]), .A1(odata[139]), .Z(xdata[139]));
Q_AN02 U695 ( .A0(sel[0]), .A1(odata[140]), .Z(xdata[140]));
Q_AN02 U696 ( .A0(sel[0]), .A1(odata[141]), .Z(xdata[141]));
Q_AN02 U697 ( .A0(sel[0]), .A1(odata[142]), .Z(xdata[142]));
Q_AN02 U698 ( .A0(sel[0]), .A1(odata[143]), .Z(xdata[143]));
Q_AN02 U699 ( .A0(sel[0]), .A1(odata[144]), .Z(xdata[144]));
Q_AN02 U700 ( .A0(sel[0]), .A1(odata[145]), .Z(xdata[145]));
Q_AN02 U701 ( .A0(sel[0]), .A1(odata[146]), .Z(xdata[146]));
Q_AN02 U702 ( .A0(sel[0]), .A1(odata[147]), .Z(xdata[147]));
Q_AN02 U703 ( .A0(sel[0]), .A1(odata[148]), .Z(xdata[148]));
Q_AN02 U704 ( .A0(sel[0]), .A1(odata[149]), .Z(xdata[149]));
Q_AN02 U705 ( .A0(sel[0]), .A1(odata[150]), .Z(xdata[150]));
Q_AN02 U706 ( .A0(sel[0]), .A1(odata[151]), .Z(xdata[151]));
Q_AN02 U707 ( .A0(sel[0]), .A1(odata[152]), .Z(xdata[152]));
Q_AN02 U708 ( .A0(sel[0]), .A1(odata[153]), .Z(xdata[153]));
Q_AN02 U709 ( .A0(sel[0]), .A1(odata[154]), .Z(xdata[154]));
Q_AN02 U710 ( .A0(sel[0]), .A1(odata[155]), .Z(xdata[155]));
Q_AN02 U711 ( .A0(sel[0]), .A1(odata[156]), .Z(xdata[156]));
Q_AN02 U712 ( .A0(sel[0]), .A1(odata[157]), .Z(xdata[157]));
Q_AN02 U713 ( .A0(sel[0]), .A1(odata[158]), .Z(xdata[158]));
Q_AN02 U714 ( .A0(sel[0]), .A1(odata[159]), .Z(xdata[159]));
Q_AN02 U715 ( .A0(sel[0]), .A1(odata[160]), .Z(xdata[160]));
Q_AN02 U716 ( .A0(sel[0]), .A1(odata[161]), .Z(xdata[161]));
Q_AN02 U717 ( .A0(sel[0]), .A1(odata[162]), .Z(xdata[162]));
Q_AN02 U718 ( .A0(sel[0]), .A1(odata[163]), .Z(xdata[163]));
Q_AN02 U719 ( .A0(sel[0]), .A1(odata[164]), .Z(xdata[164]));
Q_AN02 U720 ( .A0(sel[0]), .A1(odata[165]), .Z(xdata[165]));
Q_AN02 U721 ( .A0(sel[0]), .A1(odata[166]), .Z(xdata[166]));
Q_AN02 U722 ( .A0(sel[0]), .A1(odata[167]), .Z(xdata[167]));
Q_AN02 U723 ( .A0(sel[0]), .A1(odata[168]), .Z(xdata[168]));
Q_AN02 U724 ( .A0(sel[0]), .A1(odata[169]), .Z(xdata[169]));
Q_AN02 U725 ( .A0(sel[0]), .A1(odata[170]), .Z(xdata[170]));
Q_AN02 U726 ( .A0(sel[0]), .A1(odata[171]), .Z(xdata[171]));
Q_AN02 U727 ( .A0(sel[0]), .A1(odata[172]), .Z(xdata[172]));
Q_AN02 U728 ( .A0(sel[0]), .A1(odata[173]), .Z(xdata[173]));
Q_AN02 U729 ( .A0(sel[0]), .A1(odata[174]), .Z(xdata[174]));
Q_AN02 U730 ( .A0(sel[0]), .A1(odata[175]), .Z(xdata[175]));
Q_AN02 U731 ( .A0(sel[0]), .A1(odata[176]), .Z(xdata[176]));
Q_AN02 U732 ( .A0(sel[0]), .A1(odata[177]), .Z(xdata[177]));
Q_AN02 U733 ( .A0(sel[0]), .A1(odata[178]), .Z(xdata[178]));
Q_AN02 U734 ( .A0(sel[0]), .A1(odata[179]), .Z(xdata[179]));
Q_AN02 U735 ( .A0(sel[0]), .A1(odata[180]), .Z(xdata[180]));
Q_AN02 U736 ( .A0(sel[0]), .A1(odata[181]), .Z(xdata[181]));
Q_AN02 U737 ( .A0(sel[0]), .A1(odata[182]), .Z(xdata[182]));
Q_AN02 U738 ( .A0(sel[0]), .A1(odata[183]), .Z(xdata[183]));
Q_AN02 U739 ( .A0(sel[0]), .A1(odata[184]), .Z(xdata[184]));
Q_AN02 U740 ( .A0(sel[0]), .A1(odata[185]), .Z(xdata[185]));
Q_AN02 U741 ( .A0(sel[0]), .A1(odata[186]), .Z(xdata[186]));
Q_AN02 U742 ( .A0(sel[0]), .A1(odata[187]), .Z(xdata[187]));
Q_AN02 U743 ( .A0(sel[0]), .A1(odata[188]), .Z(xdata[188]));
Q_AN02 U744 ( .A0(sel[0]), .A1(odata[189]), .Z(xdata[189]));
Q_AN02 U745 ( .A0(sel[0]), .A1(odata[190]), .Z(xdata[190]));
Q_AN02 U746 ( .A0(sel[0]), .A1(odata[191]), .Z(xdata[191]));
Q_AN02 U747 ( .A0(sel[0]), .A1(odata[192]), .Z(xdata[192]));
Q_AN02 U748 ( .A0(sel[0]), .A1(odata[193]), .Z(xdata[193]));
Q_AN02 U749 ( .A0(sel[0]), .A1(odata[194]), .Z(xdata[194]));
Q_AN02 U750 ( .A0(sel[0]), .A1(odata[195]), .Z(xdata[195]));
Q_AN02 U751 ( .A0(sel[0]), .A1(odata[196]), .Z(xdata[196]));
Q_AN02 U752 ( .A0(sel[0]), .A1(odata[197]), .Z(xdata[197]));
Q_AN02 U753 ( .A0(sel[0]), .A1(odata[198]), .Z(xdata[198]));
Q_AN02 U754 ( .A0(sel[0]), .A1(odata[199]), .Z(xdata[199]));
Q_AN02 U755 ( .A0(sel[0]), .A1(odata[200]), .Z(xdata[200]));
Q_AN02 U756 ( .A0(sel[0]), .A1(odata[201]), .Z(xdata[201]));
Q_AN02 U757 ( .A0(sel[0]), .A1(odata[202]), .Z(xdata[202]));
Q_AN02 U758 ( .A0(sel[0]), .A1(odata[203]), .Z(xdata[203]));
Q_AN02 U759 ( .A0(sel[0]), .A1(odata[204]), .Z(xdata[204]));
Q_AN02 U760 ( .A0(sel[0]), .A1(odata[205]), .Z(xdata[205]));
Q_AN02 U761 ( .A0(sel[0]), .A1(odata[206]), .Z(xdata[206]));
Q_AN02 U762 ( .A0(sel[0]), .A1(odata[207]), .Z(xdata[207]));
Q_AN02 U763 ( .A0(sel[0]), .A1(odata[208]), .Z(xdata[208]));
Q_AN02 U764 ( .A0(sel[0]), .A1(odata[209]), .Z(xdata[209]));
Q_AN02 U765 ( .A0(sel[0]), .A1(odata[210]), .Z(xdata[210]));
Q_AN02 U766 ( .A0(sel[0]), .A1(odata[211]), .Z(xdata[211]));
Q_AN02 U767 ( .A0(sel[0]), .A1(odata[212]), .Z(xdata[212]));
Q_AN02 U768 ( .A0(sel[0]), .A1(odata[213]), .Z(xdata[213]));
Q_AN02 U769 ( .A0(sel[0]), .A1(odata[214]), .Z(xdata[214]));
Q_AN02 U770 ( .A0(sel[0]), .A1(odata[215]), .Z(xdata[215]));
Q_AN02 U771 ( .A0(sel[0]), .A1(odata[216]), .Z(xdata[216]));
Q_AN02 U772 ( .A0(sel[0]), .A1(odata[217]), .Z(xdata[217]));
Q_AN02 U773 ( .A0(sel[0]), .A1(odata[218]), .Z(xdata[218]));
Q_AN02 U774 ( .A0(sel[0]), .A1(odata[219]), .Z(xdata[219]));
Q_AN02 U775 ( .A0(sel[0]), .A1(odata[220]), .Z(xdata[220]));
Q_AN02 U776 ( .A0(sel[0]), .A1(odata[221]), .Z(xdata[221]));
Q_AN02 U777 ( .A0(sel[0]), .A1(odata[222]), .Z(xdata[222]));
Q_AN02 U778 ( .A0(sel[0]), .A1(odata[223]), .Z(xdata[223]));
Q_AN02 U779 ( .A0(sel[0]), .A1(odata[224]), .Z(xdata[224]));
Q_AN02 U780 ( .A0(sel[0]), .A1(odata[225]), .Z(xdata[225]));
Q_AN02 U781 ( .A0(sel[0]), .A1(odata[226]), .Z(xdata[226]));
Q_AN02 U782 ( .A0(sel[0]), .A1(odata[227]), .Z(xdata[227]));
Q_AN02 U783 ( .A0(sel[0]), .A1(odata[228]), .Z(xdata[228]));
Q_AN02 U784 ( .A0(sel[0]), .A1(odata[229]), .Z(xdata[229]));
Q_AN02 U785 ( .A0(sel[0]), .A1(odata[230]), .Z(xdata[230]));
Q_AN02 U786 ( .A0(sel[0]), .A1(odata[231]), .Z(xdata[231]));
Q_AN02 U787 ( .A0(sel[0]), .A1(odata[232]), .Z(xdata[232]));
Q_AN02 U788 ( .A0(sel[0]), .A1(odata[233]), .Z(xdata[233]));
Q_AN02 U789 ( .A0(sel[0]), .A1(odata[234]), .Z(xdata[234]));
Q_AN02 U790 ( .A0(sel[0]), .A1(odata[235]), .Z(xdata[235]));
Q_AN02 U791 ( .A0(sel[0]), .A1(odata[236]), .Z(xdata[236]));
Q_AN02 U792 ( .A0(sel[0]), .A1(odata[237]), .Z(xdata[237]));
Q_AN02 U793 ( .A0(sel[0]), .A1(odata[238]), .Z(xdata[238]));
Q_AN02 U794 ( .A0(sel[0]), .A1(odata[239]), .Z(xdata[239]));
Q_AN02 U795 ( .A0(sel[0]), .A1(odata[240]), .Z(xdata[240]));
Q_AN02 U796 ( .A0(sel[0]), .A1(odata[241]), .Z(xdata[241]));
Q_AN02 U797 ( .A0(sel[0]), .A1(odata[242]), .Z(xdata[242]));
Q_AN02 U798 ( .A0(sel[0]), .A1(odata[243]), .Z(xdata[243]));
Q_AN02 U799 ( .A0(sel[0]), .A1(odata[244]), .Z(xdata[244]));
Q_AN02 U800 ( .A0(sel[0]), .A1(odata[245]), .Z(xdata[245]));
Q_AN02 U801 ( .A0(sel[0]), .A1(odata[246]), .Z(xdata[246]));
Q_AN02 U802 ( .A0(sel[0]), .A1(odata[247]), .Z(xdata[247]));
Q_AN02 U803 ( .A0(sel[0]), .A1(odata[248]), .Z(xdata[248]));
Q_AN02 U804 ( .A0(sel[0]), .A1(odata[249]), .Z(xdata[249]));
Q_AN02 U805 ( .A0(sel[0]), .A1(odata[250]), .Z(xdata[250]));
Q_AN02 U806 ( .A0(sel[0]), .A1(odata[251]), .Z(xdata[251]));
Q_AN02 U807 ( .A0(sel[0]), .A1(odata[252]), .Z(xdata[252]));
Q_AN02 U808 ( .A0(sel[0]), .A1(odata[253]), .Z(xdata[253]));
Q_AN02 U809 ( .A0(sel[0]), .A1(odata[254]), .Z(xdata[254]));
Q_AN02 U810 ( .A0(sel[0]), .A1(odata[255]), .Z(xdata[255]));
Q_AN02 U811 ( .A0(sel[0]), .A1(odata[256]), .Z(xdata[256]));
Q_AN02 U812 ( .A0(sel[0]), .A1(odata[257]), .Z(xdata[257]));
Q_AN02 U813 ( .A0(sel[0]), .A1(odata[258]), .Z(xdata[258]));
Q_AN02 U814 ( .A0(sel[0]), .A1(odata[259]), .Z(xdata[259]));
Q_AN02 U815 ( .A0(sel[0]), .A1(odata[260]), .Z(xdata[260]));
Q_AN02 U816 ( .A0(sel[0]), .A1(odata[261]), .Z(xdata[261]));
Q_AN02 U817 ( .A0(sel[0]), .A1(odata[262]), .Z(xdata[262]));
Q_AN02 U818 ( .A0(sel[0]), .A1(odata[263]), .Z(xdata[263]));
Q_AN02 U819 ( .A0(sel[0]), .A1(odata[264]), .Z(xdata[264]));
Q_AN02 U820 ( .A0(sel[0]), .A1(odata[265]), .Z(xdata[265]));
Q_AN02 U821 ( .A0(sel[0]), .A1(odata[266]), .Z(xdata[266]));
Q_AN02 U822 ( .A0(sel[0]), .A1(odata[267]), .Z(xdata[267]));
Q_AN02 U823 ( .A0(sel[0]), .A1(odata[268]), .Z(xdata[268]));
Q_AN02 U824 ( .A0(sel[0]), .A1(odata[269]), .Z(xdata[269]));
Q_AN02 U825 ( .A0(sel[0]), .A1(odata[270]), .Z(xdata[270]));
Q_AN02 U826 ( .A0(sel[0]), .A1(odata[271]), .Z(xdata[271]));
Q_AN02 U827 ( .A0(sel[0]), .A1(odata[272]), .Z(xdata[272]));
Q_AN02 U828 ( .A0(sel[0]), .A1(odata[273]), .Z(xdata[273]));
Q_AN02 U829 ( .A0(sel[0]), .A1(odata[274]), .Z(xdata[274]));
Q_AN02 U830 ( .A0(sel[0]), .A1(odata[275]), .Z(xdata[275]));
Q_AN02 U831 ( .A0(sel[0]), .A1(odata[276]), .Z(xdata[276]));
Q_AN02 U832 ( .A0(sel[0]), .A1(odata[277]), .Z(xdata[277]));
Q_AN02 U833 ( .A0(sel[0]), .A1(odata[278]), .Z(xdata[278]));
Q_AN02 U834 ( .A0(sel[0]), .A1(odata[279]), .Z(xdata[279]));
Q_AN02 U835 ( .A0(sel[0]), .A1(odata[280]), .Z(xdata[280]));
Q_AN02 U836 ( .A0(sel[0]), .A1(odata[281]), .Z(xdata[281]));
Q_AN02 U837 ( .A0(sel[0]), .A1(odata[282]), .Z(xdata[282]));
Q_AN02 U838 ( .A0(sel[0]), .A1(odata[283]), .Z(xdata[283]));
Q_AN02 U839 ( .A0(sel[0]), .A1(odata[284]), .Z(xdata[284]));
Q_AN02 U840 ( .A0(sel[0]), .A1(odata[285]), .Z(xdata[285]));
Q_AN02 U841 ( .A0(sel[0]), .A1(odata[286]), .Z(xdata[286]));
Q_AN02 U842 ( .A0(sel[0]), .A1(odata[287]), .Z(xdata[287]));
Q_AN02 U843 ( .A0(sel[0]), .A1(odata[288]), .Z(xdata[288]));
Q_AN02 U844 ( .A0(sel[0]), .A1(odata[289]), .Z(xdata[289]));
Q_AN02 U845 ( .A0(sel[0]), .A1(odata[290]), .Z(xdata[290]));
Q_AN02 U846 ( .A0(sel[0]), .A1(odata[291]), .Z(xdata[291]));
Q_AN02 U847 ( .A0(sel[0]), .A1(odata[292]), .Z(xdata[292]));
Q_AN02 U848 ( .A0(sel[0]), .A1(odata[293]), .Z(xdata[293]));
Q_AN02 U849 ( .A0(sel[0]), .A1(odata[294]), .Z(xdata[294]));
Q_AN02 U850 ( .A0(sel[0]), .A1(odata[295]), .Z(xdata[295]));
Q_AN02 U851 ( .A0(sel[0]), .A1(odata[296]), .Z(xdata[296]));
Q_AN02 U852 ( .A0(sel[0]), .A1(odata[297]), .Z(xdata[297]));
Q_AN02 U853 ( .A0(sel[0]), .A1(odata[298]), .Z(xdata[298]));
Q_AN02 U854 ( .A0(sel[0]), .A1(odata[299]), .Z(xdata[299]));
Q_AN02 U855 ( .A0(sel[0]), .A1(odata[300]), .Z(xdata[300]));
Q_AN02 U856 ( .A0(sel[0]), .A1(odata[301]), .Z(xdata[301]));
Q_AN02 U857 ( .A0(sel[0]), .A1(odata[302]), .Z(xdata[302]));
Q_AN02 U858 ( .A0(sel[0]), .A1(odata[303]), .Z(xdata[303]));
Q_AN02 U859 ( .A0(sel[0]), .A1(odata[304]), .Z(xdata[304]));
Q_AN02 U860 ( .A0(sel[0]), .A1(odata[305]), .Z(xdata[305]));
Q_AN02 U861 ( .A0(sel[0]), .A1(odata[306]), .Z(xdata[306]));
Q_AN02 U862 ( .A0(sel[0]), .A1(odata[307]), .Z(xdata[307]));
Q_AN02 U863 ( .A0(sel[0]), .A1(odata[308]), .Z(xdata[308]));
Q_AN02 U864 ( .A0(sel[0]), .A1(odata[309]), .Z(xdata[309]));
Q_AN02 U865 ( .A0(sel[0]), .A1(odata[310]), .Z(xdata[310]));
Q_AN02 U866 ( .A0(sel[0]), .A1(odata[311]), .Z(xdata[311]));
Q_AN02 U867 ( .A0(sel[0]), .A1(odata[312]), .Z(xdata[312]));
Q_AN02 U868 ( .A0(sel[0]), .A1(odata[313]), .Z(xdata[313]));
Q_AN02 U869 ( .A0(sel[0]), .A1(odata[314]), .Z(xdata[314]));
Q_AN02 U870 ( .A0(sel[0]), .A1(odata[315]), .Z(xdata[315]));
Q_AN02 U871 ( .A0(sel[0]), .A1(odata[316]), .Z(xdata[316]));
Q_AN02 U872 ( .A0(sel[0]), .A1(odata[317]), .Z(xdata[317]));
Q_AN02 U873 ( .A0(sel[0]), .A1(odata[318]), .Z(xdata[318]));
Q_AN02 U874 ( .A0(sel[0]), .A1(odata[319]), .Z(xdata[319]));
Q_AN02 U875 ( .A0(sel[0]), .A1(odata[320]), .Z(xdata[320]));
Q_AN02 U876 ( .A0(sel[0]), .A1(odata[321]), .Z(xdata[321]));
Q_AN02 U877 ( .A0(sel[0]), .A1(odata[322]), .Z(xdata[322]));
Q_AN02 U878 ( .A0(sel[0]), .A1(odata[323]), .Z(xdata[323]));
Q_AN02 U879 ( .A0(sel[0]), .A1(odata[324]), .Z(xdata[324]));
Q_AN02 U880 ( .A0(sel[0]), .A1(odata[325]), .Z(xdata[325]));
Q_AN02 U881 ( .A0(sel[0]), .A1(odata[326]), .Z(xdata[326]));
Q_AN02 U882 ( .A0(sel[0]), .A1(odata[327]), .Z(xdata[327]));
Q_AN02 U883 ( .A0(sel[0]), .A1(odata[328]), .Z(xdata[328]));
Q_AN02 U884 ( .A0(sel[0]), .A1(odata[329]), .Z(xdata[329]));
Q_AN02 U885 ( .A0(sel[0]), .A1(odata[330]), .Z(xdata[330]));
Q_AN02 U886 ( .A0(sel[0]), .A1(odata[331]), .Z(xdata[331]));
Q_AN02 U887 ( .A0(sel[0]), .A1(odata[332]), .Z(xdata[332]));
Q_AN02 U888 ( .A0(sel[0]), .A1(odata[333]), .Z(xdata[333]));
Q_AN02 U889 ( .A0(sel[0]), .A1(odata[334]), .Z(xdata[334]));
Q_AN02 U890 ( .A0(sel[0]), .A1(odata[335]), .Z(xdata[335]));
Q_AN02 U891 ( .A0(sel[0]), .A1(odata[336]), .Z(xdata[336]));
Q_AN02 U892 ( .A0(sel[0]), .A1(odata[337]), .Z(xdata[337]));
Q_AN02 U893 ( .A0(sel[0]), .A1(odata[338]), .Z(xdata[338]));
Q_AN02 U894 ( .A0(sel[0]), .A1(odata[339]), .Z(xdata[339]));
Q_AN02 U895 ( .A0(sel[0]), .A1(odata[340]), .Z(xdata[340]));
Q_AN02 U896 ( .A0(sel[0]), .A1(odata[341]), .Z(xdata[341]));
Q_AN02 U897 ( .A0(sel[0]), .A1(odata[342]), .Z(xdata[342]));
Q_AN02 U898 ( .A0(sel[0]), .A1(odata[343]), .Z(xdata[343]));
Q_AN02 U899 ( .A0(sel[0]), .A1(odata[344]), .Z(xdata[344]));
Q_AN02 U900 ( .A0(sel[0]), .A1(odata[345]), .Z(xdata[345]));
Q_AN02 U901 ( .A0(sel[0]), .A1(odata[346]), .Z(xdata[346]));
Q_AN02 U902 ( .A0(sel[0]), .A1(odata[347]), .Z(xdata[347]));
Q_AN02 U903 ( .A0(sel[0]), .A1(odata[348]), .Z(xdata[348]));
Q_AN02 U904 ( .A0(sel[0]), .A1(odata[349]), .Z(xdata[349]));
Q_AN02 U905 ( .A0(sel[0]), .A1(odata[350]), .Z(xdata[350]));
Q_AN02 U906 ( .A0(sel[0]), .A1(odata[351]), .Z(xdata[351]));
Q_AN02 U907 ( .A0(sel[0]), .A1(odata[352]), .Z(xdata[352]));
Q_AN02 U908 ( .A0(sel[0]), .A1(odata[353]), .Z(xdata[353]));
Q_AN02 U909 ( .A0(sel[0]), .A1(odata[354]), .Z(xdata[354]));
Q_AN02 U910 ( .A0(sel[0]), .A1(odata[355]), .Z(xdata[355]));
Q_AN02 U911 ( .A0(sel[0]), .A1(odata[356]), .Z(xdata[356]));
Q_AN02 U912 ( .A0(sel[0]), .A1(odata[357]), .Z(xdata[357]));
Q_AN02 U913 ( .A0(sel[0]), .A1(odata[358]), .Z(xdata[358]));
Q_AN02 U914 ( .A0(sel[0]), .A1(odata[359]), .Z(xdata[359]));
Q_AN02 U915 ( .A0(sel[0]), .A1(odata[360]), .Z(xdata[360]));
Q_AN02 U916 ( .A0(sel[0]), .A1(odata[361]), .Z(xdata[361]));
Q_AN02 U917 ( .A0(sel[0]), .A1(odata[362]), .Z(xdata[362]));
Q_AN02 U918 ( .A0(sel[0]), .A1(odata[363]), .Z(xdata[363]));
Q_AN02 U919 ( .A0(sel[0]), .A1(odata[364]), .Z(xdata[364]));
Q_AN02 U920 ( .A0(sel[0]), .A1(odata[365]), .Z(xdata[365]));
Q_AN02 U921 ( .A0(sel[0]), .A1(odata[366]), .Z(xdata[366]));
Q_AN02 U922 ( .A0(sel[0]), .A1(odata[367]), .Z(xdata[367]));
Q_AN02 U923 ( .A0(sel[0]), .A1(odata[368]), .Z(xdata[368]));
Q_AN02 U924 ( .A0(sel[0]), .A1(odata[369]), .Z(xdata[369]));
Q_AN02 U925 ( .A0(sel[0]), .A1(odata[370]), .Z(xdata[370]));
Q_AN02 U926 ( .A0(sel[0]), .A1(odata[371]), .Z(xdata[371]));
Q_AN02 U927 ( .A0(sel[0]), .A1(odata[372]), .Z(xdata[372]));
Q_AN02 U928 ( .A0(sel[0]), .A1(odata[373]), .Z(xdata[373]));
Q_AN02 U929 ( .A0(sel[0]), .A1(odata[374]), .Z(xdata[374]));
Q_AN02 U930 ( .A0(sel[0]), .A1(odata[375]), .Z(xdata[375]));
Q_AN02 U931 ( .A0(sel[0]), .A1(odata[376]), .Z(xdata[376]));
Q_AN02 U932 ( .A0(sel[0]), .A1(odata[377]), .Z(xdata[377]));
Q_AN02 U933 ( .A0(sel[0]), .A1(odata[378]), .Z(xdata[378]));
Q_AN02 U934 ( .A0(sel[0]), .A1(odata[379]), .Z(xdata[379]));
Q_AN02 U935 ( .A0(sel[0]), .A1(odata[380]), .Z(xdata[380]));
Q_AN02 U936 ( .A0(sel[0]), .A1(odata[381]), .Z(xdata[381]));
Q_AN02 U937 ( .A0(sel[0]), .A1(odata[382]), .Z(xdata[382]));
Q_AN02 U938 ( .A0(sel[0]), .A1(odata[383]), .Z(xdata[383]));
Q_AN02 U939 ( .A0(sel[0]), .A1(odata[384]), .Z(xdata[384]));
Q_AN02 U940 ( .A0(sel[0]), .A1(odata[385]), .Z(xdata[385]));
Q_AN02 U941 ( .A0(sel[0]), .A1(odata[386]), .Z(xdata[386]));
Q_AN02 U942 ( .A0(sel[0]), .A1(odata[387]), .Z(xdata[387]));
Q_AN02 U943 ( .A0(sel[0]), .A1(odata[388]), .Z(xdata[388]));
Q_AN02 U944 ( .A0(sel[0]), .A1(odata[389]), .Z(xdata[389]));
Q_AN02 U945 ( .A0(sel[0]), .A1(odata[390]), .Z(xdata[390]));
Q_AN02 U946 ( .A0(sel[0]), .A1(odata[391]), .Z(xdata[391]));
Q_AN02 U947 ( .A0(sel[0]), .A1(odata[392]), .Z(xdata[392]));
Q_AN02 U948 ( .A0(sel[0]), .A1(odata[393]), .Z(xdata[393]));
Q_AN02 U949 ( .A0(sel[0]), .A1(odata[394]), .Z(xdata[394]));
Q_AN02 U950 ( .A0(sel[0]), .A1(odata[395]), .Z(xdata[395]));
Q_AN02 U951 ( .A0(sel[0]), .A1(odata[396]), .Z(xdata[396]));
Q_AN02 U952 ( .A0(sel[0]), .A1(odata[397]), .Z(xdata[397]));
Q_AN02 U953 ( .A0(sel[0]), .A1(odata[398]), .Z(xdata[398]));
Q_AN02 U954 ( .A0(sel[0]), .A1(odata[399]), .Z(xdata[399]));
Q_AN02 U955 ( .A0(sel[0]), .A1(odata[400]), .Z(xdata[400]));
Q_AN02 U956 ( .A0(sel[0]), .A1(odata[401]), .Z(xdata[401]));
Q_AN02 U957 ( .A0(sel[0]), .A1(odata[402]), .Z(xdata[402]));
Q_AN02 U958 ( .A0(sel[0]), .A1(odata[403]), .Z(xdata[403]));
Q_AN02 U959 ( .A0(sel[0]), .A1(odata[404]), .Z(xdata[404]));
Q_AN02 U960 ( .A0(sel[0]), .A1(odata[405]), .Z(xdata[405]));
Q_AN02 U961 ( .A0(sel[0]), .A1(odata[406]), .Z(xdata[406]));
Q_AN02 U962 ( .A0(sel[0]), .A1(odata[407]), .Z(xdata[407]));
Q_AN02 U963 ( .A0(sel[0]), .A1(odata[408]), .Z(xdata[408]));
Q_AN02 U964 ( .A0(sel[0]), .A1(odata[409]), .Z(xdata[409]));
Q_AN02 U965 ( .A0(sel[0]), .A1(odata[410]), .Z(xdata[410]));
Q_AN02 U966 ( .A0(sel[0]), .A1(odata[411]), .Z(xdata[411]));
Q_AN02 U967 ( .A0(sel[0]), .A1(odata[412]), .Z(xdata[412]));
Q_AN02 U968 ( .A0(sel[0]), .A1(odata[413]), .Z(xdata[413]));
Q_AN02 U969 ( .A0(sel[0]), .A1(odata[414]), .Z(xdata[414]));
Q_AN02 U970 ( .A0(sel[0]), .A1(odata[415]), .Z(xdata[415]));
Q_AN02 U971 ( .A0(sel[0]), .A1(odata[416]), .Z(xdata[416]));
Q_AN02 U972 ( .A0(sel[0]), .A1(odata[417]), .Z(xdata[417]));
Q_AN02 U973 ( .A0(sel[0]), .A1(odata[418]), .Z(xdata[418]));
Q_AN02 U974 ( .A0(sel[0]), .A1(odata[419]), .Z(xdata[419]));
Q_AN02 U975 ( .A0(sel[0]), .A1(odata[420]), .Z(xdata[420]));
Q_AN02 U976 ( .A0(sel[0]), .A1(odata[421]), .Z(xdata[421]));
Q_AN02 U977 ( .A0(sel[0]), .A1(odata[422]), .Z(xdata[422]));
Q_AN02 U978 ( .A0(sel[0]), .A1(odata[423]), .Z(xdata[423]));
Q_AN02 U979 ( .A0(sel[0]), .A1(odata[424]), .Z(xdata[424]));
Q_AN02 U980 ( .A0(sel[0]), .A1(odata[425]), .Z(xdata[425]));
Q_AN02 U981 ( .A0(sel[0]), .A1(odata[426]), .Z(xdata[426]));
Q_AN02 U982 ( .A0(sel[0]), .A1(odata[427]), .Z(xdata[427]));
Q_AN02 U983 ( .A0(sel[0]), .A1(odata[428]), .Z(xdata[428]));
Q_AN02 U984 ( .A0(sel[0]), .A1(odata[429]), .Z(xdata[429]));
Q_AN02 U985 ( .A0(sel[0]), .A1(odata[430]), .Z(xdata[430]));
Q_AN02 U986 ( .A0(sel[0]), .A1(odata[431]), .Z(xdata[431]));
Q_AN02 U987 ( .A0(sel[0]), .A1(odata[432]), .Z(xdata[432]));
Q_AN02 U988 ( .A0(sel[0]), .A1(odata[433]), .Z(xdata[433]));
Q_AN02 U989 ( .A0(sel[0]), .A1(odata[434]), .Z(xdata[434]));
Q_AN02 U990 ( .A0(sel[0]), .A1(odata[435]), .Z(xdata[435]));
Q_AN02 U991 ( .A0(sel[0]), .A1(odata[436]), .Z(xdata[436]));
Q_AN02 U992 ( .A0(sel[0]), .A1(odata[437]), .Z(xdata[437]));
Q_AN02 U993 ( .A0(sel[0]), .A1(odata[438]), .Z(xdata[438]));
Q_AN02 U994 ( .A0(sel[0]), .A1(odata[439]), .Z(xdata[439]));
Q_AN02 U995 ( .A0(sel[0]), .A1(odata[440]), .Z(xdata[440]));
Q_AN02 U996 ( .A0(sel[0]), .A1(odata[441]), .Z(xdata[441]));
Q_AN02 U997 ( .A0(sel[0]), .A1(odata[442]), .Z(xdata[442]));
Q_AN02 U998 ( .A0(sel[0]), .A1(odata[443]), .Z(xdata[443]));
Q_AN02 U999 ( .A0(sel[0]), .A1(odata[444]), .Z(xdata[444]));
Q_AN02 U1000 ( .A0(sel[0]), .A1(odata[445]), .Z(xdata[445]));
Q_AN02 U1001 ( .A0(sel[0]), .A1(odata[446]), .Z(xdata[446]));
Q_AN02 U1002 ( .A0(sel[0]), .A1(odata[447]), .Z(xdata[447]));
Q_AN02 U1003 ( .A0(sel[0]), .A1(odata[448]), .Z(xdata[448]));
Q_AN02 U1004 ( .A0(sel[0]), .A1(odata[449]), .Z(xdata[449]));
Q_AN02 U1005 ( .A0(sel[0]), .A1(odata[450]), .Z(xdata[450]));
Q_AN02 U1006 ( .A0(sel[0]), .A1(odata[451]), .Z(xdata[451]));
Q_AN02 U1007 ( .A0(sel[0]), .A1(odata[452]), .Z(xdata[452]));
Q_AN02 U1008 ( .A0(sel[0]), .A1(odata[453]), .Z(xdata[453]));
Q_AN02 U1009 ( .A0(sel[0]), .A1(odata[454]), .Z(xdata[454]));
Q_AN02 U1010 ( .A0(sel[0]), .A1(odata[455]), .Z(xdata[455]));
Q_AN02 U1011 ( .A0(sel[0]), .A1(odata[456]), .Z(xdata[456]));
Q_AN02 U1012 ( .A0(sel[0]), .A1(odata[457]), .Z(xdata[457]));
Q_AN02 U1013 ( .A0(sel[0]), .A1(odata[458]), .Z(xdata[458]));
Q_AN02 U1014 ( .A0(sel[0]), .A1(odata[459]), .Z(xdata[459]));
Q_AN02 U1015 ( .A0(sel[0]), .A1(odata[460]), .Z(xdata[460]));
Q_AN02 U1016 ( .A0(sel[0]), .A1(odata[461]), .Z(xdata[461]));
Q_AN02 U1017 ( .A0(sel[0]), .A1(odata[462]), .Z(xdata[462]));
Q_AN02 U1018 ( .A0(sel[0]), .A1(odata[463]), .Z(xdata[463]));
Q_AN02 U1019 ( .A0(sel[0]), .A1(odata[464]), .Z(xdata[464]));
Q_AN02 U1020 ( .A0(sel[0]), .A1(odata[465]), .Z(xdata[465]));
Q_AN02 U1021 ( .A0(sel[0]), .A1(odata[466]), .Z(xdata[466]));
Q_AN02 U1022 ( .A0(sel[0]), .A1(odata[467]), .Z(xdata[467]));
Q_AN02 U1023 ( .A0(sel[0]), .A1(odata[468]), .Z(xdata[468]));
Q_AN02 U1024 ( .A0(sel[0]), .A1(odata[469]), .Z(xdata[469]));
Q_AN02 U1025 ( .A0(sel[0]), .A1(odata[470]), .Z(xdata[470]));
Q_AN02 U1026 ( .A0(sel[0]), .A1(odata[471]), .Z(xdata[471]));
Q_AN02 U1027 ( .A0(sel[0]), .A1(odata[472]), .Z(xdata[472]));
Q_AN02 U1028 ( .A0(sel[0]), .A1(odata[473]), .Z(xdata[473]));
Q_AN02 U1029 ( .A0(sel[0]), .A1(odata[474]), .Z(xdata[474]));
Q_AN02 U1030 ( .A0(sel[0]), .A1(odata[475]), .Z(xdata[475]));
Q_AN02 U1031 ( .A0(sel[0]), .A1(odata[476]), .Z(xdata[476]));
Q_AN02 U1032 ( .A0(sel[0]), .A1(odata[477]), .Z(xdata[477]));
Q_AN02 U1033 ( .A0(sel[0]), .A1(odata[478]), .Z(xdata[478]));
Q_AN02 U1034 ( .A0(sel[0]), .A1(odata[479]), .Z(xdata[479]));
Q_AN02 U1035 ( .A0(sel[0]), .A1(odata[480]), .Z(xdata[480]));
Q_AN02 U1036 ( .A0(sel[0]), .A1(odata[481]), .Z(xdata[481]));
Q_AN02 U1037 ( .A0(sel[0]), .A1(odata[482]), .Z(xdata[482]));
Q_AN02 U1038 ( .A0(sel[0]), .A1(odata[483]), .Z(xdata[483]));
Q_AN02 U1039 ( .A0(sel[0]), .A1(odata[484]), .Z(xdata[484]));
Q_AN02 U1040 ( .A0(sel[0]), .A1(odata[485]), .Z(xdata[485]));
Q_AN02 U1041 ( .A0(sel[0]), .A1(odata[486]), .Z(xdata[486]));
Q_AN02 U1042 ( .A0(sel[0]), .A1(odata[487]), .Z(xdata[487]));
Q_AN02 U1043 ( .A0(sel[0]), .A1(odata[488]), .Z(xdata[488]));
Q_AN02 U1044 ( .A0(sel[0]), .A1(odata[489]), .Z(xdata[489]));
Q_AN02 U1045 ( .A0(sel[0]), .A1(odata[490]), .Z(xdata[490]));
Q_AN02 U1046 ( .A0(sel[0]), .A1(odata[491]), .Z(xdata[491]));
Q_AN02 U1047 ( .A0(sel[0]), .A1(odata[492]), .Z(xdata[492]));
Q_AN02 U1048 ( .A0(sel[0]), .A1(odata[493]), .Z(xdata[493]));
Q_AN02 U1049 ( .A0(sel[0]), .A1(odata[494]), .Z(xdata[494]));
Q_AN02 U1050 ( .A0(sel[0]), .A1(odata[495]), .Z(xdata[495]));
Q_AN02 U1051 ( .A0(sel[0]), .A1(odata[496]), .Z(xdata[496]));
Q_AN02 U1052 ( .A0(sel[0]), .A1(odata[497]), .Z(xdata[497]));
Q_AN02 U1053 ( .A0(sel[0]), .A1(odata[498]), .Z(xdata[498]));
Q_AN02 U1054 ( .A0(sel[0]), .A1(odata[499]), .Z(xdata[499]));
Q_AN02 U1055 ( .A0(sel[0]), .A1(odata[500]), .Z(xdata[500]));
Q_AN02 U1056 ( .A0(sel[0]), .A1(odata[501]), .Z(xdata[501]));
Q_AN02 U1057 ( .A0(sel[0]), .A1(odata[502]), .Z(xdata[502]));
Q_AN02 U1058 ( .A0(sel[0]), .A1(odata[503]), .Z(xdata[503]));
Q_AN02 U1059 ( .A0(sel[0]), .A1(odata[504]), .Z(xdata[504]));
Q_AN02 U1060 ( .A0(sel[0]), .A1(odata[505]), .Z(xdata[505]));
Q_AN02 U1061 ( .A0(sel[0]), .A1(odata[506]), .Z(xdata[506]));
Q_AN02 U1062 ( .A0(sel[0]), .A1(odata[507]), .Z(xdata[507]));
Q_AN02 U1063 ( .A0(sel[0]), .A1(odata[508]), .Z(xdata[508]));
Q_AN02 U1064 ( .A0(sel[0]), .A1(odata[509]), .Z(xdata[509]));
Q_AN02 U1065 ( .A0(sel[0]), .A1(odata[510]), .Z(xdata[510]));
Q_AN02 U1066 ( .A0(sel[0]), .A1(odata[511]), .Z(xdata[511]));
Q_AN02 U1067 ( .A0(sel[1]), .A1(odata[512]), .Z(n7));
Q_AN02 U1068 ( .A0(sel[1]), .A1(odata[513]), .Z(n8));
Q_AN02 U1069 ( .A0(sel[1]), .A1(odata[514]), .Z(n9));
Q_AN02 U1070 ( .A0(sel[1]), .A1(odata[515]), .Z(n10));
Q_AN02 U1071 ( .A0(sel[1]), .A1(odata[516]), .Z(n11));
Q_AN02 U1072 ( .A0(sel[1]), .A1(odata[517]), .Z(n12));
Q_AN02 U1073 ( .A0(sel[1]), .A1(odata[518]), .Z(n13));
Q_AN02 U1074 ( .A0(sel[1]), .A1(odata[519]), .Z(n14));
Q_AN02 U1075 ( .A0(sel[1]), .A1(odata[520]), .Z(n15));
Q_AN02 U1076 ( .A0(sel[1]), .A1(odata[521]), .Z(n16));
Q_AN02 U1077 ( .A0(sel[1]), .A1(odata[522]), .Z(n17));
Q_AN02 U1078 ( .A0(sel[1]), .A1(odata[523]), .Z(n18));
Q_AN02 U1079 ( .A0(sel[1]), .A1(odata[524]), .Z(n19));
Q_AN02 U1080 ( .A0(sel[1]), .A1(odata[525]), .Z(n20));
Q_AN02 U1081 ( .A0(sel[1]), .A1(odata[526]), .Z(n21));
Q_AN02 U1082 ( .A0(sel[1]), .A1(odata[527]), .Z(n22));
Q_AN02 U1083 ( .A0(sel[1]), .A1(odata[528]), .Z(n23));
Q_AN02 U1084 ( .A0(sel[1]), .A1(odata[529]), .Z(n24));
Q_AN02 U1085 ( .A0(sel[1]), .A1(odata[530]), .Z(n25));
Q_AN02 U1086 ( .A0(sel[1]), .A1(odata[531]), .Z(n26));
Q_AN02 U1087 ( .A0(sel[1]), .A1(odata[532]), .Z(n27));
Q_AN02 U1088 ( .A0(sel[1]), .A1(odata[533]), .Z(n28));
Q_AN02 U1089 ( .A0(sel[1]), .A1(odata[534]), .Z(n29));
Q_AN02 U1090 ( .A0(sel[1]), .A1(odata[535]), .Z(n30));
Q_AN02 U1091 ( .A0(sel[1]), .A1(odata[536]), .Z(n31));
Q_AN02 U1092 ( .A0(sel[1]), .A1(odata[537]), .Z(n32));
Q_AN02 U1093 ( .A0(sel[1]), .A1(odata[538]), .Z(n33));
Q_AN02 U1094 ( .A0(sel[1]), .A1(odata[539]), .Z(n34));
Q_AN02 U1095 ( .A0(sel[1]), .A1(odata[540]), .Z(n35));
Q_AN02 U1096 ( .A0(sel[1]), .A1(odata[541]), .Z(n36));
Q_AN02 U1097 ( .A0(sel[1]), .A1(odata[542]), .Z(n37));
Q_AN02 U1098 ( .A0(sel[1]), .A1(odata[543]), .Z(n38));
Q_AN02 U1099 ( .A0(sel[1]), .A1(odata[544]), .Z(n39));
Q_AN02 U1100 ( .A0(sel[1]), .A1(odata[545]), .Z(n40));
Q_AN02 U1101 ( .A0(sel[1]), .A1(odata[546]), .Z(n41));
Q_AN02 U1102 ( .A0(sel[1]), .A1(odata[547]), .Z(n42));
Q_AN02 U1103 ( .A0(sel[1]), .A1(odata[548]), .Z(n43));
Q_AN02 U1104 ( .A0(sel[1]), .A1(odata[549]), .Z(n44));
Q_AN02 U1105 ( .A0(sel[1]), .A1(odata[550]), .Z(n45));
Q_AN02 U1106 ( .A0(sel[1]), .A1(odata[551]), .Z(n46));
Q_AN02 U1107 ( .A0(sel[1]), .A1(odata[552]), .Z(n47));
Q_AN02 U1108 ( .A0(sel[1]), .A1(odata[553]), .Z(n48));
Q_AN02 U1109 ( .A0(sel[1]), .A1(odata[554]), .Z(n49));
Q_AN02 U1110 ( .A0(sel[1]), .A1(odata[555]), .Z(n50));
Q_AN02 U1111 ( .A0(sel[1]), .A1(odata[556]), .Z(n51));
Q_AN02 U1112 ( .A0(sel[1]), .A1(odata[557]), .Z(n52));
Q_AN02 U1113 ( .A0(sel[1]), .A1(odata[558]), .Z(n53));
Q_AN02 U1114 ( .A0(sel[1]), .A1(odata[559]), .Z(n54));
Q_BUFZP U1115 ( .OE(enq), .A(n6), .Z(CLBreq));
Q_BUFZP U1116 ( .OE(enq), .A(n6), .Z(CGFtsReq));
Q_INV U1117 ( .A(CLBwr[2]), .Z(n55));
ixc_bind \genblk3.b5 ( CLBfull, IXC_GFIFO.O.O.LBfull);
ixc_bind_4 \genblk3.b4 ( CLBwr[3:0], IXC_GFIFO.O.O.LBwr[3:0]);
ixc_bind_4 \genblk3.b3 ( CLBrd[3:0], IXC_GFIFO.O.O.LBrd[3:0]);
ixc_bind \genblk3.b2 ( CLBreq, IXC_GFIFO.O.O.LBreq);
ixc_bind \genblk3.b1 ( CGFfull, IXC_GFIFO.O.O.GFfull);
ixc_bind \genblk3.b0 ( CGFtsReq, IXC_GFIFO.O.O.GFtsReq);
Q_OR03 U1124 ( .A0(olen[9]), .A1(olen[8]), .A2(n57), .Z(n58));
Q_OR02 U1125 ( .A0(olen[11]), .A1(olen[10]), .Z(n57));
Q_OR03 U1126 ( .A0(olen[7]), .A1(olen[6]), .A2(olen[5]), .Z(n59));
Q_OR03 U1127 ( .A0(olen[1]), .A1(olen[0]), .A2(n60), .Z(n61));
Q_OR02 U1128 ( .A0(olen[3]), .A1(olen[2]), .Z(n60));
Q_AN02 U1129 ( .A0(olen[4]), .A1(n61), .Z(n62));
Q_OR03 U1130 ( .A0(n58), .A1(n59), .A2(n62), .Z(n171));
Q_XNR2 U1131 ( .A0(xlen[4]), .A1(CGFfull), .Z(n63));
Q_OR02 U1132 ( .A0(xlen[4]), .A1(CGFfull), .Z(n64));
Q_XNR2 U1133 ( .A0(xlen[5]), .A1(n64), .Z(n65));
Q_OR02 U1134 ( .A0(xlen[5]), .A1(n64), .Z(n66));
Q_XNR2 U1135 ( .A0(xlen[6]), .A1(n66), .Z(n67));
Q_OR02 U1136 ( .A0(xlen[6]), .A1(n66), .Z(n68));
Q_XNR2 U1137 ( .A0(xlen[7]), .A1(n68), .Z(n69));
Q_OR02 U1138 ( .A0(xlen[7]), .A1(n68), .Z(n70));
Q_XNR2 U1139 ( .A0(xlen[8]), .A1(n70), .Z(n71));
Q_OR02 U1140 ( .A0(xlen[8]), .A1(n70), .Z(n72));
Q_XNR2 U1141 ( .A0(xlen[9]), .A1(n72), .Z(n73));
Q_OR02 U1142 ( .A0(xlen[9]), .A1(n72), .Z(n74));
Q_XNR2 U1143 ( .A0(xlen[10]), .A1(n74), .Z(n75));
Q_OR02 U1144 ( .A0(xlen[10]), .A1(n74), .Z(n76));
Q_XNR2 U1145 ( .A0(xlen[11]), .A1(n76), .Z(n77));
Q_OR03 U1146 ( .A0(n73), .A1(n71), .A2(n78), .Z(n79));
Q_OR02 U1147 ( .A0(n77), .A1(n75), .Z(n78));
Q_OR03 U1148 ( .A0(n69), .A1(n67), .A2(n65), .Z(n80));
Q_OR03 U1149 ( .A0(xlen[1]), .A1(xlen[0]), .A2(n81), .Z(n82));
Q_OR02 U1150 ( .A0(xlen[3]), .A1(xlen[2]), .Z(n81));
Q_AN02 U1151 ( .A0(n63), .A1(n82), .Z(n83));
Q_OR03 U1152 ( .A0(n79), .A1(n80), .A2(n83), .Z(n172));
Q_OR02 U1153 ( .A0(State_Var), .A1(ocbid[0]), .Z(n84));
Q_OR02 U1154 ( .A0(State_Var), .A1(ocbid[1]), .Z(n85));
Q_OR02 U1155 ( .A0(State_Var), .A1(ocbid[2]), .Z(n86));
Q_OR02 U1156 ( .A0(State_Var), .A1(ocbid[3]), .Z(n87));
Q_OR02 U1157 ( .A0(State_Var), .A1(ocbid[4]), .Z(n88));
Q_OR02 U1158 ( .A0(State_Var), .A1(ocbid[5]), .Z(n89));
Q_OR02 U1159 ( .A0(State_Var), .A1(ocbid[6]), .Z(n90));
Q_OR02 U1160 ( .A0(State_Var), .A1(ocbid[7]), .Z(n91));
Q_OR02 U1161 ( .A0(State_Var), .A1(ocbid[8]), .Z(n92));
Q_OR02 U1162 ( .A0(State_Var), .A1(ocbid[9]), .Z(n93));
Q_OR02 U1163 ( .A0(State_Var), .A1(ocbid[10]), .Z(n94));
Q_OR02 U1164 ( .A0(State_Var), .A1(ocbid[11]), .Z(n95));
Q_OR02 U1165 ( .A0(State_Var), .A1(ocbid[12]), .Z(n96));
Q_OR02 U1166 ( .A0(State_Var), .A1(ocbid[13]), .Z(n97));
Q_OR02 U1167 ( .A0(State_Var), .A1(ocbid[14]), .Z(n98));
Q_OR02 U1168 ( .A0(State_Var), .A1(ocbid[15]), .Z(n99));
Q_OR02 U1169 ( .A0(State_Var), .A1(ocbid[16]), .Z(n100));
Q_OR02 U1170 ( .A0(State_Var), .A1(ocbid[17]), .Z(n101));
Q_OR02 U1171 ( .A0(State_Var), .A1(ocbid[18]), .Z(n102));
Q_OR02 U1172 ( .A0(State_Var), .A1(ocbid[19]), .Z(n103));
Q_MX02 U1173 ( .S(n157), .A0(ireq), .A1(oreq), .Z(n104));
Q_MX02 U1174 ( .S(State_Var), .A0(olen[4]), .A1(n63), .Z(n105));
Q_MX02 U1175 ( .S(State_Var), .A0(olen[5]), .A1(n65), .Z(n106));
Q_MX02 U1176 ( .S(State_Var), .A0(olen[6]), .A1(n67), .Z(n107));
Q_MX02 U1177 ( .S(State_Var), .A0(olen[7]), .A1(n69), .Z(n108));
Q_MX02 U1178 ( .S(State_Var), .A0(olen[8]), .A1(n71), .Z(n109));
Q_MX02 U1179 ( .S(State_Var), .A0(olen[9]), .A1(n73), .Z(n110));
Q_MX02 U1180 ( .S(State_Var), .A0(olen[10]), .A1(n75), .Z(n111));
Q_MX02 U1181 ( .S(State_Var), .A0(olen[11]), .A1(n77), .Z(n112));
Q_INV U1182 ( .A(State_Var), .Z(n113));
Q_AN02 U1183 ( .A0(State_Var), .A1(sel[0]), .Z(n114));
Q_FDP0UA U1184 ( .D(n115), .QTFCLK( ), .Q(ack));
Q_MX02 U1185 ( .S(n170), .A0(ack), .A1(n104), .Z(n115));
Q_FDP0UA U1186 ( .D(n116), .QTFCLK( ), .Q(xcbid[19]));
Q_MX02 U1187 ( .S(n168), .A0(xcbid[19]), .A1(n103), .Z(n116));
Q_FDP0UA U1188 ( .D(n117), .QTFCLK( ), .Q(xcbid[18]));
Q_MX02 U1189 ( .S(n168), .A0(xcbid[18]), .A1(n102), .Z(n117));
Q_FDP0UA U1190 ( .D(n118), .QTFCLK( ), .Q(xcbid[17]));
Q_MX02 U1191 ( .S(n168), .A0(xcbid[17]), .A1(n101), .Z(n118));
Q_FDP0UA U1192 ( .D(n119), .QTFCLK( ), .Q(xcbid[16]));
Q_MX02 U1193 ( .S(n168), .A0(xcbid[16]), .A1(n100), .Z(n119));
Q_FDP0UA U1194 ( .D(n120), .QTFCLK( ), .Q(xcbid[15]));
Q_MX02 U1195 ( .S(n168), .A0(xcbid[15]), .A1(n99), .Z(n120));
Q_FDP0UA U1196 ( .D(n121), .QTFCLK( ), .Q(xcbid[14]));
Q_MX02 U1197 ( .S(n168), .A0(xcbid[14]), .A1(n98), .Z(n121));
Q_FDP0UA U1198 ( .D(n122), .QTFCLK( ), .Q(xcbid[13]));
Q_MX02 U1199 ( .S(n168), .A0(xcbid[13]), .A1(n97), .Z(n122));
Q_FDP0UA U1200 ( .D(n123), .QTFCLK( ), .Q(xcbid[12]));
Q_MX02 U1201 ( .S(n168), .A0(xcbid[12]), .A1(n96), .Z(n123));
Q_FDP0UA U1202 ( .D(n124), .QTFCLK( ), .Q(xcbid[11]));
Q_MX02 U1203 ( .S(n168), .A0(xcbid[11]), .A1(n95), .Z(n124));
Q_FDP0UA U1204 ( .D(n125), .QTFCLK( ), .Q(xcbid[10]));
Q_MX02 U1205 ( .S(n168), .A0(xcbid[10]), .A1(n94), .Z(n125));
Q_FDP0UA U1206 ( .D(n126), .QTFCLK( ), .Q(xcbid[9]));
Q_MX02 U1207 ( .S(n168), .A0(xcbid[9]), .A1(n93), .Z(n126));
Q_FDP0UA U1208 ( .D(n127), .QTFCLK( ), .Q(xcbid[8]));
Q_MX02 U1209 ( .S(n168), .A0(xcbid[8]), .A1(n92), .Z(n127));
Q_FDP0UA U1210 ( .D(n128), .QTFCLK( ), .Q(xcbid[7]));
Q_MX02 U1211 ( .S(n168), .A0(xcbid[7]), .A1(n91), .Z(n128));
Q_FDP0UA U1212 ( .D(n129), .QTFCLK( ), .Q(xcbid[6]));
Q_MX02 U1213 ( .S(n168), .A0(xcbid[6]), .A1(n90), .Z(n129));
Q_FDP0UA U1214 ( .D(n130), .QTFCLK( ), .Q(xcbid[5]));
Q_MX02 U1215 ( .S(n168), .A0(xcbid[5]), .A1(n89), .Z(n130));
Q_FDP0UA U1216 ( .D(n131), .QTFCLK( ), .Q(xcbid[4]));
Q_MX02 U1217 ( .S(n168), .A0(xcbid[4]), .A1(n88), .Z(n131));
Q_FDP0UA U1218 ( .D(n132), .QTFCLK( ), .Q(xcbid[3]));
Q_MX02 U1219 ( .S(n168), .A0(xcbid[3]), .A1(n87), .Z(n132));
Q_FDP0UA U1220 ( .D(n133), .QTFCLK( ), .Q(xcbid[2]));
Q_MX02 U1221 ( .S(n168), .A0(xcbid[2]), .A1(n86), .Z(n133));
Q_FDP0UA U1222 ( .D(n134), .QTFCLK( ), .Q(xcbid[1]));
Q_MX02 U1223 ( .S(n168), .A0(xcbid[1]), .A1(n85), .Z(n134));
Q_FDP0UA U1224 ( .D(n135), .QTFCLK( ), .Q(xcbid[0]));
Q_MX02 U1225 ( .S(n168), .A0(xcbid[0]), .A1(n84), .Z(n135));
Q_FDP0UA U1226 ( .D(n136), .QTFCLK( ), .Q(xlen[11]));
Q_MX02 U1227 ( .S(n169), .A0(xlen[11]), .A1(n112), .Z(n136));
Q_FDP0UA U1228 ( .D(n137), .QTFCLK( ), .Q(xlen[10]));
Q_MX02 U1229 ( .S(n169), .A0(xlen[10]), .A1(n111), .Z(n137));
Q_FDP0UA U1230 ( .D(n138), .QTFCLK( ), .Q(xlen[9]));
Q_MX02 U1231 ( .S(n169), .A0(xlen[9]), .A1(n110), .Z(n138));
Q_FDP0UA U1232 ( .D(n139), .QTFCLK( ), .Q(xlen[8]));
Q_MX02 U1233 ( .S(n169), .A0(xlen[8]), .A1(n109), .Z(n139));
Q_FDP0UA U1234 ( .D(n140), .QTFCLK( ), .Q(xlen[7]));
Q_MX02 U1235 ( .S(n169), .A0(xlen[7]), .A1(n108), .Z(n140));
Q_FDP0UA U1236 ( .D(n141), .QTFCLK( ), .Q(xlen[6]));
Q_MX02 U1237 ( .S(n169), .A0(xlen[6]), .A1(n107), .Z(n141));
Q_FDP0UA U1238 ( .D(n142), .QTFCLK( ), .Q(xlen[5]));
Q_MX02 U1239 ( .S(n169), .A0(xlen[5]), .A1(n106), .Z(n142));
Q_FDP0UA U1240 ( .D(n143), .QTFCLK( ), .Q(xlen[4]));
Q_MX02 U1241 ( .S(n169), .A0(xlen[4]), .A1(n105), .Z(n143));
Q_FDP0UA U1242 ( .D(n144), .QTFCLK( ), .Q(xlen[3]));
Q_MX02 U1243 ( .S(n1), .A0(xlen[3]), .A1(olen[3]), .Z(n144));
Q_FDP0UA U1244 ( .D(n145), .QTFCLK( ), .Q(xlen[2]));
Q_MX02 U1245 ( .S(n1), .A0(xlen[2]), .A1(olen[2]), .Z(n145));
Q_FDP0UA U1246 ( .D(n146), .QTFCLK( ), .Q(xlen[1]));
Q_MX02 U1247 ( .S(n1), .A0(xlen[1]), .A1(olen[1]), .Z(n146));
Q_FDP0UA U1248 ( .D(n147), .QTFCLK( ), .Q(xlen[0]));
Q_MX02 U1249 ( .S(n1), .A0(xlen[0]), .A1(olen[0]), .Z(n147));
Q_FDP0UA U1250 ( .D(n148), .QTFCLK( ), .Q(sel[1]));
Q_MX02 U1251 ( .S(n168), .A0(sel[1]), .A1(n114), .Z(n148));
Q_FDP0UA U1252 ( .D(n149), .QTFCLK( ), .Q(sel[0]));
Q_MX02 U1253 ( .S(n168), .A0(sel[0]), .A1(n113), .Z(n149));
Q_FDP0UA U1254 ( .D(n150), .QTFCLK( ), .Q(en));
Q_MX02 U1255 ( .S(State_Var), .A0(n167), .A1(en), .Z(n150));
Q_FDP0UA U1256 ( .D(n166), .QTFCLK( ), .Q(State_Var));
Q_AN02 U1257 ( .A0(State_Var), .A1(n172), .Z(n151));
Q_AO21 U1258 ( .A0(n152), .A1(n153), .B0(n151), .Z(n166));
Q_AN02 U1259 ( .A0(n154), .A1(n171), .Z(n153));
Q_AN02 U1260 ( .A0(n155), .A1(n156), .Z(n152));
Q_NR02 U1261 ( .A0(State_Var), .A1(xc_top.GFLock2), .Z(n155));
Q_ND02 U1262 ( .A0(n113), .A1(xc_top.GFLock2), .Z(n157));
Q_OR02 U1263 ( .A0(n167), .A1(State_Var), .Z(n169));
Q_AN02 U1264 ( .A0(n158), .A1(n154), .Z(n167));
Q_MX02 U1265 ( .S(State_Var), .A0(n160), .A1(n159), .Z(n170));
Q_INV U1266 ( .A(n172), .Z(n159));
Q_AO21 U1267 ( .A0(n154), .A1(n161), .B0(xc_top.GFLock2), .Z(n160));
Q_AN02 U1268 ( .A0(n156), .A1(n162), .Z(n161));
Q_INV U1269 ( .A(n171), .Z(n162));
Q_AN02 U1270 ( .A0(n163), .A1(n164), .Z(n154));
Q_INV U1271 ( .A(CGFfull), .Z(n164));
Q_OA21 U1272 ( .A0(State_Var), .A1(n165), .B0(n164), .Z(n168));
Q_AN02 U1273 ( .A0(n158), .A1(n163), .Z(n165));
Q_INV U1274 ( .A(Rtkin), .Z(n163));
Q_AN02 U1275 ( .A0(n4), .A1(n156), .Z(n158));
Q_NR02 U1276 ( .A0(n5), .A1(tkin), .Z(n156));
Q_MX02 U1277 ( .S(CLBfull), .A0(ireq), .A1(ireqR), .Z(n173));
Q_FDP0UA U1278 ( .D(n173), .QTFCLK( ), .Q(ireqR));
Q_AN02 U1279 ( .A0(CLBwr[0]), .A1(n55), .Z(n174));
Q_AN02 U1280 ( .A0(CLBwr[1]), .A1(n55), .Z(n175));
Q_INV U1281 ( .A(n174), .Z(n176));
Q_INV U1282 ( .A(n175), .Z(n177));
Q_NR02 U1283 ( .A0(n175), .A1(n174), .Z(n178));
Q_AN02 U1284 ( .A0(n177), .A1(n174), .Z(n179));
Q_AN02 U1285 ( .A0(n175), .A1(n176), .Z(n180));
Q_AN02 U1286 ( .A0(n175), .A1(n174), .Z(n181));
Q_AN02 U1287 ( .A0(n178), .A1(n55), .Z(n182));
Q_LDP0 \_zzLB_REG[0][0] ( .G(n182), .D(len[0]), .Q(\_zzLB[0][0] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][1] ( .G(n182), .D(len[1]), .Q(\_zzLB[0][1] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][2] ( .G(n182), .D(len[2]), .Q(\_zzLB[0][2] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][3] ( .G(n182), .D(len[3]), .Q(\_zzLB[0][3] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][4] ( .G(n182), .D(len[4]), .Q(\_zzLB[0][4] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][5] ( .G(n182), .D(len[5]), .Q(\_zzLB[0][5] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][6] ( .G(n182), .D(len[6]), .Q(\_zzLB[0][6] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][7] ( .G(n182), .D(len[7]), .Q(\_zzLB[0][7] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][8] ( .G(n182), .D(len[8]), .Q(\_zzLB[0][8] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][9] ( .G(n182), .D(len[9]), .Q(\_zzLB[0][9] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][10] ( .G(n182), .D(len[10]), .Q(\_zzLB[0][10] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][11] ( .G(n182), .D(len[11]), .Q(\_zzLB[0][11] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][12] ( .G(n182), .D(cbid[0]), .Q(\_zzLB[0][12] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][13] ( .G(n182), .D(cbid[1]), .Q(\_zzLB[0][13] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][14] ( .G(n182), .D(cbid[2]), .Q(\_zzLB[0][14] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][15] ( .G(n182), .D(cbid[3]), .Q(\_zzLB[0][15] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][16] ( .G(n182), .D(cbid[4]), .Q(\_zzLB[0][16] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][17] ( .G(n182), .D(cbid[5]), .Q(\_zzLB[0][17] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][18] ( .G(n182), .D(cbid[6]), .Q(\_zzLB[0][18] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][19] ( .G(n182), .D(cbid[7]), .Q(\_zzLB[0][19] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][20] ( .G(n182), .D(cbid[8]), .Q(\_zzLB[0][20] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][21] ( .G(n182), .D(cbid[9]), .Q(\_zzLB[0][21] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][22] ( .G(n182), .D(cbid[10]), .Q(\_zzLB[0][22] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][23] ( .G(n182), .D(cbid[11]), .Q(\_zzLB[0][23] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][24] ( .G(n182), .D(cbid[12]), .Q(\_zzLB[0][24] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][25] ( .G(n182), .D(cbid[13]), .Q(\_zzLB[0][25] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][26] ( .G(n182), .D(cbid[14]), .Q(\_zzLB[0][26] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][27] ( .G(n182), .D(cbid[15]), .Q(\_zzLB[0][27] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][28] ( .G(n182), .D(cbid[16]), .Q(\_zzLB[0][28] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][29] ( .G(n182), .D(cbid[17]), .Q(\_zzLB[0][29] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][30] ( .G(n182), .D(cbid[18]), .Q(\_zzLB[0][30] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][31] ( .G(n182), .D(cbid[19]), .Q(\_zzLB[0][31] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][32] ( .G(n182), .D(idata[0]), .Q(\_zzLB[0][32] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][33] ( .G(n182), .D(idata[1]), .Q(\_zzLB[0][33] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][34] ( .G(n182), .D(idata[2]), .Q(\_zzLB[0][34] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][35] ( .G(n182), .D(idata[3]), .Q(\_zzLB[0][35] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][36] ( .G(n182), .D(idata[4]), .Q(\_zzLB[0][36] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][37] ( .G(n182), .D(idata[5]), .Q(\_zzLB[0][37] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][38] ( .G(n182), .D(idata[6]), .Q(\_zzLB[0][38] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][39] ( .G(n182), .D(idata[7]), .Q(\_zzLB[0][39] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][40] ( .G(n182), .D(idata[8]), .Q(\_zzLB[0][40] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][41] ( .G(n182), .D(idata[9]), .Q(\_zzLB[0][41] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][42] ( .G(n182), .D(idata[10]), .Q(\_zzLB[0][42] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][43] ( .G(n182), .D(idata[11]), .Q(\_zzLB[0][43] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][44] ( .G(n182), .D(idata[12]), .Q(\_zzLB[0][44] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][45] ( .G(n182), .D(idata[13]), .Q(\_zzLB[0][45] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][46] ( .G(n182), .D(idata[14]), .Q(\_zzLB[0][46] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][47] ( .G(n182), .D(idata[15]), .Q(\_zzLB[0][47] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][48] ( .G(n182), .D(idata[16]), .Q(\_zzLB[0][48] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][49] ( .G(n182), .D(idata[17]), .Q(\_zzLB[0][49] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][50] ( .G(n182), .D(idata[18]), .Q(\_zzLB[0][50] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][51] ( .G(n182), .D(idata[19]), .Q(\_zzLB[0][51] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][52] ( .G(n182), .D(idata[20]), .Q(\_zzLB[0][52] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][53] ( .G(n182), .D(idata[21]), .Q(\_zzLB[0][53] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][54] ( .G(n182), .D(idata[22]), .Q(\_zzLB[0][54] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][55] ( .G(n182), .D(idata[23]), .Q(\_zzLB[0][55] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][56] ( .G(n182), .D(idata[24]), .Q(\_zzLB[0][56] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][57] ( .G(n182), .D(idata[25]), .Q(\_zzLB[0][57] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][58] ( .G(n182), .D(idata[26]), .Q(\_zzLB[0][58] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][59] ( .G(n182), .D(idata[27]), .Q(\_zzLB[0][59] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][60] ( .G(n182), .D(idata[28]), .Q(\_zzLB[0][60] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][61] ( .G(n182), .D(idata[29]), .Q(\_zzLB[0][61] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][62] ( .G(n182), .D(idata[30]), .Q(\_zzLB[0][62] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][63] ( .G(n182), .D(idata[31]), .Q(\_zzLB[0][63] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][64] ( .G(n182), .D(idata[32]), .Q(\_zzLB[0][64] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][65] ( .G(n182), .D(idata[33]), .Q(\_zzLB[0][65] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][66] ( .G(n182), .D(idata[34]), .Q(\_zzLB[0][66] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][67] ( .G(n182), .D(idata[35]), .Q(\_zzLB[0][67] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][68] ( .G(n182), .D(idata[36]), .Q(\_zzLB[0][68] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][69] ( .G(n182), .D(idata[37]), .Q(\_zzLB[0][69] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][70] ( .G(n182), .D(idata[38]), .Q(\_zzLB[0][70] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][71] ( .G(n182), .D(idata[39]), .Q(\_zzLB[0][71] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][72] ( .G(n182), .D(idata[40]), .Q(\_zzLB[0][72] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][73] ( .G(n182), .D(idata[41]), .Q(\_zzLB[0][73] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][74] ( .G(n182), .D(idata[42]), .Q(\_zzLB[0][74] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][75] ( .G(n182), .D(idata[43]), .Q(\_zzLB[0][75] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][76] ( .G(n182), .D(idata[44]), .Q(\_zzLB[0][76] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][77] ( .G(n182), .D(idata[45]), .Q(\_zzLB[0][77] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][78] ( .G(n182), .D(idata[46]), .Q(\_zzLB[0][78] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][79] ( .G(n182), .D(idata[47]), .Q(\_zzLB[0][79] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][80] ( .G(n182), .D(idata[48]), .Q(\_zzLB[0][80] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][81] ( .G(n182), .D(idata[49]), .Q(\_zzLB[0][81] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][82] ( .G(n182), .D(idata[50]), .Q(\_zzLB[0][82] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][83] ( .G(n182), .D(idata[51]), .Q(\_zzLB[0][83] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][84] ( .G(n182), .D(idata[52]), .Q(\_zzLB[0][84] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][85] ( .G(n182), .D(idata[53]), .Q(\_zzLB[0][85] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][86] ( .G(n182), .D(idata[54]), .Q(\_zzLB[0][86] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][87] ( .G(n182), .D(idata[55]), .Q(\_zzLB[0][87] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][88] ( .G(n182), .D(idata[56]), .Q(\_zzLB[0][88] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][89] ( .G(n182), .D(idata[57]), .Q(\_zzLB[0][89] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][90] ( .G(n182), .D(idata[58]), .Q(\_zzLB[0][90] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][91] ( .G(n182), .D(idata[59]), .Q(\_zzLB[0][91] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][92] ( .G(n182), .D(idata[60]), .Q(\_zzLB[0][92] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][93] ( .G(n182), .D(idata[61]), .Q(\_zzLB[0][93] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][94] ( .G(n182), .D(idata[62]), .Q(\_zzLB[0][94] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][95] ( .G(n182), .D(idata[63]), .Q(\_zzLB[0][95] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][96] ( .G(n182), .D(idata[64]), .Q(\_zzLB[0][96] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][97] ( .G(n182), .D(idata[65]), .Q(\_zzLB[0][97] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][98] ( .G(n182), .D(idata[66]), .Q(\_zzLB[0][98] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][99] ( .G(n182), .D(idata[67]), .Q(\_zzLB[0][99] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][100] ( .G(n182), .D(idata[68]), .Q(\_zzLB[0][100] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][101] ( .G(n182), .D(idata[69]), .Q(\_zzLB[0][101] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][102] ( .G(n182), .D(idata[70]), .Q(\_zzLB[0][102] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][103] ( .G(n182), .D(idata[71]), .Q(\_zzLB[0][103] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][104] ( .G(n182), .D(idata[72]), .Q(\_zzLB[0][104] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][105] ( .G(n182), .D(idata[73]), .Q(\_zzLB[0][105] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][106] ( .G(n182), .D(idata[74]), .Q(\_zzLB[0][106] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][107] ( .G(n182), .D(idata[75]), .Q(\_zzLB[0][107] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][108] ( .G(n182), .D(idata[76]), .Q(\_zzLB[0][108] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][109] ( .G(n182), .D(idata[77]), .Q(\_zzLB[0][109] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][110] ( .G(n182), .D(idata[78]), .Q(\_zzLB[0][110] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][111] ( .G(n182), .D(idata[79]), .Q(\_zzLB[0][111] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][112] ( .G(n182), .D(idata[80]), .Q(\_zzLB[0][112] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][113] ( .G(n182), .D(idata[81]), .Q(\_zzLB[0][113] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][114] ( .G(n182), .D(idata[82]), .Q(\_zzLB[0][114] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][115] ( .G(n182), .D(idata[83]), .Q(\_zzLB[0][115] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][116] ( .G(n182), .D(idata[84]), .Q(\_zzLB[0][116] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][117] ( .G(n182), .D(idata[85]), .Q(\_zzLB[0][117] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][118] ( .G(n182), .D(idata[86]), .Q(\_zzLB[0][118] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][119] ( .G(n182), .D(idata[87]), .Q(\_zzLB[0][119] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][120] ( .G(n182), .D(idata[88]), .Q(\_zzLB[0][120] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][121] ( .G(n182), .D(idata[89]), .Q(\_zzLB[0][121] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][122] ( .G(n182), .D(idata[90]), .Q(\_zzLB[0][122] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][123] ( .G(n182), .D(idata[91]), .Q(\_zzLB[0][123] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][124] ( .G(n182), .D(idata[92]), .Q(\_zzLB[0][124] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][125] ( .G(n182), .D(idata[93]), .Q(\_zzLB[0][125] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][126] ( .G(n182), .D(idata[94]), .Q(\_zzLB[0][126] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][127] ( .G(n182), .D(idata[95]), .Q(\_zzLB[0][127] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][128] ( .G(n182), .D(idata[96]), .Q(\_zzLB[0][128] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][129] ( .G(n182), .D(idata[97]), .Q(\_zzLB[0][129] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][130] ( .G(n182), .D(idata[98]), .Q(\_zzLB[0][130] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][131] ( .G(n182), .D(idata[99]), .Q(\_zzLB[0][131] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][132] ( .G(n182), .D(idata[100]), .Q(\_zzLB[0][132] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][133] ( .G(n182), .D(idata[101]), .Q(\_zzLB[0][133] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][134] ( .G(n182), .D(idata[102]), .Q(\_zzLB[0][134] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][135] ( .G(n182), .D(idata[103]), .Q(\_zzLB[0][135] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][136] ( .G(n182), .D(idata[104]), .Q(\_zzLB[0][136] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][137] ( .G(n182), .D(idata[105]), .Q(\_zzLB[0][137] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][138] ( .G(n182), .D(idata[106]), .Q(\_zzLB[0][138] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][139] ( .G(n182), .D(idata[107]), .Q(\_zzLB[0][139] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][140] ( .G(n182), .D(idata[108]), .Q(\_zzLB[0][140] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][141] ( .G(n182), .D(idata[109]), .Q(\_zzLB[0][141] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][142] ( .G(n182), .D(idata[110]), .Q(\_zzLB[0][142] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][143] ( .G(n182), .D(idata[111]), .Q(\_zzLB[0][143] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][144] ( .G(n182), .D(idata[112]), .Q(\_zzLB[0][144] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][145] ( .G(n182), .D(idata[113]), .Q(\_zzLB[0][145] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][146] ( .G(n182), .D(idata[114]), .Q(\_zzLB[0][146] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][147] ( .G(n182), .D(idata[115]), .Q(\_zzLB[0][147] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][148] ( .G(n182), .D(idata[116]), .Q(\_zzLB[0][148] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][149] ( .G(n182), .D(idata[117]), .Q(\_zzLB[0][149] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][150] ( .G(n182), .D(idata[118]), .Q(\_zzLB[0][150] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][151] ( .G(n182), .D(idata[119]), .Q(\_zzLB[0][151] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][152] ( .G(n182), .D(idata[120]), .Q(\_zzLB[0][152] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][153] ( .G(n182), .D(idata[121]), .Q(\_zzLB[0][153] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][154] ( .G(n182), .D(idata[122]), .Q(\_zzLB[0][154] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][155] ( .G(n182), .D(idata[123]), .Q(\_zzLB[0][155] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][156] ( .G(n182), .D(idata[124]), .Q(\_zzLB[0][156] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][157] ( .G(n182), .D(idata[125]), .Q(\_zzLB[0][157] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][158] ( .G(n182), .D(idata[126]), .Q(\_zzLB[0][158] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][159] ( .G(n182), .D(idata[127]), .Q(\_zzLB[0][159] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][160] ( .G(n182), .D(idata[128]), .Q(\_zzLB[0][160] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][161] ( .G(n182), .D(idata[129]), .Q(\_zzLB[0][161] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][162] ( .G(n182), .D(idata[130]), .Q(\_zzLB[0][162] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][163] ( .G(n182), .D(idata[131]), .Q(\_zzLB[0][163] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][164] ( .G(n182), .D(idata[132]), .Q(\_zzLB[0][164] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][165] ( .G(n182), .D(idata[133]), .Q(\_zzLB[0][165] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][166] ( .G(n182), .D(idata[134]), .Q(\_zzLB[0][166] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][167] ( .G(n182), .D(idata[135]), .Q(\_zzLB[0][167] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][168] ( .G(n182), .D(idata[136]), .Q(\_zzLB[0][168] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][169] ( .G(n182), .D(idata[137]), .Q(\_zzLB[0][169] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][170] ( .G(n182), .D(idata[138]), .Q(\_zzLB[0][170] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][171] ( .G(n182), .D(idata[139]), .Q(\_zzLB[0][171] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][172] ( .G(n182), .D(idata[140]), .Q(\_zzLB[0][172] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][173] ( .G(n182), .D(idata[141]), .Q(\_zzLB[0][173] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][174] ( .G(n182), .D(idata[142]), .Q(\_zzLB[0][174] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][175] ( .G(n182), .D(idata[143]), .Q(\_zzLB[0][175] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][176] ( .G(n182), .D(idata[144]), .Q(\_zzLB[0][176] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][177] ( .G(n182), .D(idata[145]), .Q(\_zzLB[0][177] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][178] ( .G(n182), .D(idata[146]), .Q(\_zzLB[0][178] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][179] ( .G(n182), .D(idata[147]), .Q(\_zzLB[0][179] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][180] ( .G(n182), .D(idata[148]), .Q(\_zzLB[0][180] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][181] ( .G(n182), .D(idata[149]), .Q(\_zzLB[0][181] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][182] ( .G(n182), .D(idata[150]), .Q(\_zzLB[0][182] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][183] ( .G(n182), .D(idata[151]), .Q(\_zzLB[0][183] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][184] ( .G(n182), .D(idata[152]), .Q(\_zzLB[0][184] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][185] ( .G(n182), .D(idata[153]), .Q(\_zzLB[0][185] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][186] ( .G(n182), .D(idata[154]), .Q(\_zzLB[0][186] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][187] ( .G(n182), .D(idata[155]), .Q(\_zzLB[0][187] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][188] ( .G(n182), .D(idata[156]), .Q(\_zzLB[0][188] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][189] ( .G(n182), .D(idata[157]), .Q(\_zzLB[0][189] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][190] ( .G(n182), .D(idata[158]), .Q(\_zzLB[0][190] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][191] ( .G(n182), .D(idata[159]), .Q(\_zzLB[0][191] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][192] ( .G(n182), .D(idata[160]), .Q(\_zzLB[0][192] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][193] ( .G(n182), .D(idata[161]), .Q(\_zzLB[0][193] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][194] ( .G(n182), .D(idata[162]), .Q(\_zzLB[0][194] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][195] ( .G(n182), .D(idata[163]), .Q(\_zzLB[0][195] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][196] ( .G(n182), .D(idata[164]), .Q(\_zzLB[0][196] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][197] ( .G(n182), .D(idata[165]), .Q(\_zzLB[0][197] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][198] ( .G(n182), .D(idata[166]), .Q(\_zzLB[0][198] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][199] ( .G(n182), .D(idata[167]), .Q(\_zzLB[0][199] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][200] ( .G(n182), .D(idata[168]), .Q(\_zzLB[0][200] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][201] ( .G(n182), .D(idata[169]), .Q(\_zzLB[0][201] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][202] ( .G(n182), .D(idata[170]), .Q(\_zzLB[0][202] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][203] ( .G(n182), .D(idata[171]), .Q(\_zzLB[0][203] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][204] ( .G(n182), .D(idata[172]), .Q(\_zzLB[0][204] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][205] ( .G(n182), .D(idata[173]), .Q(\_zzLB[0][205] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][206] ( .G(n182), .D(idata[174]), .Q(\_zzLB[0][206] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][207] ( .G(n182), .D(idata[175]), .Q(\_zzLB[0][207] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][208] ( .G(n182), .D(idata[176]), .Q(\_zzLB[0][208] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][209] ( .G(n182), .D(idata[177]), .Q(\_zzLB[0][209] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][210] ( .G(n182), .D(idata[178]), .Q(\_zzLB[0][210] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][211] ( .G(n182), .D(idata[179]), .Q(\_zzLB[0][211] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][212] ( .G(n182), .D(idata[180]), .Q(\_zzLB[0][212] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][213] ( .G(n182), .D(idata[181]), .Q(\_zzLB[0][213] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][214] ( .G(n182), .D(idata[182]), .Q(\_zzLB[0][214] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][215] ( .G(n182), .D(idata[183]), .Q(\_zzLB[0][215] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][216] ( .G(n182), .D(idata[184]), .Q(\_zzLB[0][216] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][217] ( .G(n182), .D(idata[185]), .Q(\_zzLB[0][217] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][218] ( .G(n182), .D(idata[186]), .Q(\_zzLB[0][218] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][219] ( .G(n182), .D(idata[187]), .Q(\_zzLB[0][219] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][220] ( .G(n182), .D(idata[188]), .Q(\_zzLB[0][220] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][221] ( .G(n182), .D(idata[189]), .Q(\_zzLB[0][221] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][222] ( .G(n182), .D(idata[190]), .Q(\_zzLB[0][222] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][223] ( .G(n182), .D(idata[191]), .Q(\_zzLB[0][223] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][224] ( .G(n182), .D(idata[192]), .Q(\_zzLB[0][224] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][225] ( .G(n182), .D(idata[193]), .Q(\_zzLB[0][225] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][226] ( .G(n182), .D(idata[194]), .Q(\_zzLB[0][226] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][227] ( .G(n182), .D(idata[195]), .Q(\_zzLB[0][227] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][228] ( .G(n182), .D(idata[196]), .Q(\_zzLB[0][228] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][229] ( .G(n182), .D(idata[197]), .Q(\_zzLB[0][229] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][230] ( .G(n182), .D(idata[198]), .Q(\_zzLB[0][230] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][231] ( .G(n182), .D(idata[199]), .Q(\_zzLB[0][231] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][232] ( .G(n182), .D(idata[200]), .Q(\_zzLB[0][232] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][233] ( .G(n182), .D(idata[201]), .Q(\_zzLB[0][233] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][234] ( .G(n182), .D(idata[202]), .Q(\_zzLB[0][234] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][235] ( .G(n182), .D(idata[203]), .Q(\_zzLB[0][235] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][236] ( .G(n182), .D(idata[204]), .Q(\_zzLB[0][236] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][237] ( .G(n182), .D(idata[205]), .Q(\_zzLB[0][237] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][238] ( .G(n182), .D(idata[206]), .Q(\_zzLB[0][238] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][239] ( .G(n182), .D(idata[207]), .Q(\_zzLB[0][239] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][240] ( .G(n182), .D(idata[208]), .Q(\_zzLB[0][240] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][241] ( .G(n182), .D(idata[209]), .Q(\_zzLB[0][241] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][242] ( .G(n182), .D(idata[210]), .Q(\_zzLB[0][242] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][243] ( .G(n182), .D(idata[211]), .Q(\_zzLB[0][243] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][244] ( .G(n182), .D(idata[212]), .Q(\_zzLB[0][244] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][245] ( .G(n182), .D(idata[213]), .Q(\_zzLB[0][245] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][246] ( .G(n182), .D(idata[214]), .Q(\_zzLB[0][246] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][247] ( .G(n182), .D(idata[215]), .Q(\_zzLB[0][247] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][248] ( .G(n182), .D(idata[216]), .Q(\_zzLB[0][248] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][249] ( .G(n182), .D(idata[217]), .Q(\_zzLB[0][249] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][250] ( .G(n182), .D(idata[218]), .Q(\_zzLB[0][250] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][251] ( .G(n182), .D(idata[219]), .Q(\_zzLB[0][251] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][252] ( .G(n182), .D(idata[220]), .Q(\_zzLB[0][252] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][253] ( .G(n182), .D(idata[221]), .Q(\_zzLB[0][253] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][254] ( .G(n182), .D(idata[222]), .Q(\_zzLB[0][254] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][255] ( .G(n182), .D(idata[223]), .Q(\_zzLB[0][255] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][256] ( .G(n182), .D(idata[224]), .Q(\_zzLB[0][256] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][257] ( .G(n182), .D(idata[225]), .Q(\_zzLB[0][257] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][258] ( .G(n182), .D(idata[226]), .Q(\_zzLB[0][258] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][259] ( .G(n182), .D(idata[227]), .Q(\_zzLB[0][259] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][260] ( .G(n182), .D(idata[228]), .Q(\_zzLB[0][260] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][261] ( .G(n182), .D(idata[229]), .Q(\_zzLB[0][261] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][262] ( .G(n182), .D(idata[230]), .Q(\_zzLB[0][262] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][263] ( .G(n182), .D(idata[231]), .Q(\_zzLB[0][263] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][264] ( .G(n182), .D(idata[232]), .Q(\_zzLB[0][264] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][265] ( .G(n182), .D(idata[233]), .Q(\_zzLB[0][265] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][266] ( .G(n182), .D(idata[234]), .Q(\_zzLB[0][266] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][267] ( .G(n182), .D(idata[235]), .Q(\_zzLB[0][267] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][268] ( .G(n182), .D(idata[236]), .Q(\_zzLB[0][268] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][269] ( .G(n182), .D(idata[237]), .Q(\_zzLB[0][269] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][270] ( .G(n182), .D(idata[238]), .Q(\_zzLB[0][270] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][271] ( .G(n182), .D(idata[239]), .Q(\_zzLB[0][271] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][272] ( .G(n182), .D(idata[240]), .Q(\_zzLB[0][272] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][273] ( .G(n182), .D(idata[241]), .Q(\_zzLB[0][273] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][274] ( .G(n182), .D(idata[242]), .Q(\_zzLB[0][274] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][275] ( .G(n182), .D(idata[243]), .Q(\_zzLB[0][275] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][276] ( .G(n182), .D(idata[244]), .Q(\_zzLB[0][276] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][277] ( .G(n182), .D(idata[245]), .Q(\_zzLB[0][277] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][278] ( .G(n182), .D(idata[246]), .Q(\_zzLB[0][278] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][279] ( .G(n182), .D(idata[247]), .Q(\_zzLB[0][279] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][280] ( .G(n182), .D(idata[248]), .Q(\_zzLB[0][280] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][281] ( .G(n182), .D(idata[249]), .Q(\_zzLB[0][281] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][282] ( .G(n182), .D(idata[250]), .Q(\_zzLB[0][282] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][283] ( .G(n182), .D(idata[251]), .Q(\_zzLB[0][283] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][284] ( .G(n182), .D(idata[252]), .Q(\_zzLB[0][284] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][285] ( .G(n182), .D(idata[253]), .Q(\_zzLB[0][285] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][286] ( .G(n182), .D(idata[254]), .Q(\_zzLB[0][286] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][287] ( .G(n182), .D(idata[255]), .Q(\_zzLB[0][287] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][288] ( .G(n182), .D(idata[256]), .Q(\_zzLB[0][288] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][289] ( .G(n182), .D(idata[257]), .Q(\_zzLB[0][289] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][290] ( .G(n182), .D(idata[258]), .Q(\_zzLB[0][290] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][291] ( .G(n182), .D(idata[259]), .Q(\_zzLB[0][291] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][292] ( .G(n182), .D(idata[260]), .Q(\_zzLB[0][292] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][293] ( .G(n182), .D(idata[261]), .Q(\_zzLB[0][293] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][294] ( .G(n182), .D(idata[262]), .Q(\_zzLB[0][294] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][295] ( .G(n182), .D(idata[263]), .Q(\_zzLB[0][295] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][296] ( .G(n182), .D(idata[264]), .Q(\_zzLB[0][296] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][297] ( .G(n182), .D(idata[265]), .Q(\_zzLB[0][297] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][298] ( .G(n182), .D(idata[266]), .Q(\_zzLB[0][298] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][299] ( .G(n182), .D(idata[267]), .Q(\_zzLB[0][299] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][300] ( .G(n182), .D(idata[268]), .Q(\_zzLB[0][300] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][301] ( .G(n182), .D(idata[269]), .Q(\_zzLB[0][301] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][302] ( .G(n182), .D(idata[270]), .Q(\_zzLB[0][302] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][303] ( .G(n182), .D(idata[271]), .Q(\_zzLB[0][303] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][304] ( .G(n182), .D(idata[272]), .Q(\_zzLB[0][304] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][305] ( .G(n182), .D(idata[273]), .Q(\_zzLB[0][305] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][306] ( .G(n182), .D(idata[274]), .Q(\_zzLB[0][306] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][307] ( .G(n182), .D(idata[275]), .Q(\_zzLB[0][307] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][308] ( .G(n182), .D(idata[276]), .Q(\_zzLB[0][308] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][309] ( .G(n182), .D(idata[277]), .Q(\_zzLB[0][309] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][310] ( .G(n182), .D(idata[278]), .Q(\_zzLB[0][310] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][311] ( .G(n182), .D(idata[279]), .Q(\_zzLB[0][311] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][312] ( .G(n182), .D(idata[280]), .Q(\_zzLB[0][312] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][313] ( .G(n182), .D(idata[281]), .Q(\_zzLB[0][313] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][314] ( .G(n182), .D(idata[282]), .Q(\_zzLB[0][314] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][315] ( .G(n182), .D(idata[283]), .Q(\_zzLB[0][315] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][316] ( .G(n182), .D(idata[284]), .Q(\_zzLB[0][316] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][317] ( .G(n182), .D(idata[285]), .Q(\_zzLB[0][317] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][318] ( .G(n182), .D(idata[286]), .Q(\_zzLB[0][318] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][319] ( .G(n182), .D(idata[287]), .Q(\_zzLB[0][319] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][320] ( .G(n182), .D(idata[288]), .Q(\_zzLB[0][320] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][321] ( .G(n182), .D(idata[289]), .Q(\_zzLB[0][321] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][322] ( .G(n182), .D(idata[290]), .Q(\_zzLB[0][322] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][323] ( .G(n182), .D(idata[291]), .Q(\_zzLB[0][323] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][324] ( .G(n182), .D(idata[292]), .Q(\_zzLB[0][324] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][325] ( .G(n182), .D(idata[293]), .Q(\_zzLB[0][325] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][326] ( .G(n182), .D(idata[294]), .Q(\_zzLB[0][326] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][327] ( .G(n182), .D(idata[295]), .Q(\_zzLB[0][327] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][328] ( .G(n182), .D(idata[296]), .Q(\_zzLB[0][328] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][329] ( .G(n182), .D(idata[297]), .Q(\_zzLB[0][329] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][330] ( .G(n182), .D(idata[298]), .Q(\_zzLB[0][330] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][331] ( .G(n182), .D(idata[299]), .Q(\_zzLB[0][331] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][332] ( .G(n182), .D(idata[300]), .Q(\_zzLB[0][332] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][333] ( .G(n182), .D(idata[301]), .Q(\_zzLB[0][333] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][334] ( .G(n182), .D(idata[302]), .Q(\_zzLB[0][334] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][335] ( .G(n182), .D(idata[303]), .Q(\_zzLB[0][335] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][336] ( .G(n182), .D(idata[304]), .Q(\_zzLB[0][336] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][337] ( .G(n182), .D(idata[305]), .Q(\_zzLB[0][337] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][338] ( .G(n182), .D(idata[306]), .Q(\_zzLB[0][338] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][339] ( .G(n182), .D(idata[307]), .Q(\_zzLB[0][339] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][340] ( .G(n182), .D(idata[308]), .Q(\_zzLB[0][340] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][341] ( .G(n182), .D(idata[309]), .Q(\_zzLB[0][341] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][342] ( .G(n182), .D(idata[310]), .Q(\_zzLB[0][342] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][343] ( .G(n182), .D(idata[311]), .Q(\_zzLB[0][343] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][344] ( .G(n182), .D(idata[312]), .Q(\_zzLB[0][344] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][345] ( .G(n182), .D(idata[313]), .Q(\_zzLB[0][345] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][346] ( .G(n182), .D(idata[314]), .Q(\_zzLB[0][346] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][347] ( .G(n182), .D(idata[315]), .Q(\_zzLB[0][347] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][348] ( .G(n182), .D(idata[316]), .Q(\_zzLB[0][348] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][349] ( .G(n182), .D(idata[317]), .Q(\_zzLB[0][349] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][350] ( .G(n182), .D(idata[318]), .Q(\_zzLB[0][350] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][351] ( .G(n182), .D(idata[319]), .Q(\_zzLB[0][351] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][352] ( .G(n182), .D(idata[320]), .Q(\_zzLB[0][352] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][353] ( .G(n182), .D(idata[321]), .Q(\_zzLB[0][353] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][354] ( .G(n182), .D(idata[322]), .Q(\_zzLB[0][354] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][355] ( .G(n182), .D(idata[323]), .Q(\_zzLB[0][355] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][356] ( .G(n182), .D(idata[324]), .Q(\_zzLB[0][356] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][357] ( .G(n182), .D(idata[325]), .Q(\_zzLB[0][357] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][358] ( .G(n182), .D(idata[326]), .Q(\_zzLB[0][358] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][359] ( .G(n182), .D(idata[327]), .Q(\_zzLB[0][359] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][360] ( .G(n182), .D(idata[328]), .Q(\_zzLB[0][360] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][361] ( .G(n182), .D(idata[329]), .Q(\_zzLB[0][361] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][362] ( .G(n182), .D(idata[330]), .Q(\_zzLB[0][362] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][363] ( .G(n182), .D(idata[331]), .Q(\_zzLB[0][363] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][364] ( .G(n182), .D(idata[332]), .Q(\_zzLB[0][364] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][365] ( .G(n182), .D(idata[333]), .Q(\_zzLB[0][365] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][366] ( .G(n182), .D(idata[334]), .Q(\_zzLB[0][366] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][367] ( .G(n182), .D(idata[335]), .Q(\_zzLB[0][367] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][368] ( .G(n182), .D(idata[336]), .Q(\_zzLB[0][368] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][369] ( .G(n182), .D(idata[337]), .Q(\_zzLB[0][369] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][370] ( .G(n182), .D(idata[338]), .Q(\_zzLB[0][370] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][371] ( .G(n182), .D(idata[339]), .Q(\_zzLB[0][371] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][372] ( .G(n182), .D(idata[340]), .Q(\_zzLB[0][372] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][373] ( .G(n182), .D(idata[341]), .Q(\_zzLB[0][373] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][374] ( .G(n182), .D(idata[342]), .Q(\_zzLB[0][374] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][375] ( .G(n182), .D(idata[343]), .Q(\_zzLB[0][375] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][376] ( .G(n182), .D(idata[344]), .Q(\_zzLB[0][376] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][377] ( .G(n182), .D(idata[345]), .Q(\_zzLB[0][377] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][378] ( .G(n182), .D(idata[346]), .Q(\_zzLB[0][378] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][379] ( .G(n182), .D(idata[347]), .Q(\_zzLB[0][379] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][380] ( .G(n182), .D(idata[348]), .Q(\_zzLB[0][380] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][381] ( .G(n182), .D(idata[349]), .Q(\_zzLB[0][381] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][382] ( .G(n182), .D(idata[350]), .Q(\_zzLB[0][382] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][383] ( .G(n182), .D(idata[351]), .Q(\_zzLB[0][383] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][384] ( .G(n182), .D(idata[352]), .Q(\_zzLB[0][384] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][385] ( .G(n182), .D(idata[353]), .Q(\_zzLB[0][385] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][386] ( .G(n182), .D(idata[354]), .Q(\_zzLB[0][386] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][387] ( .G(n182), .D(idata[355]), .Q(\_zzLB[0][387] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][388] ( .G(n182), .D(idata[356]), .Q(\_zzLB[0][388] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][389] ( .G(n182), .D(idata[357]), .Q(\_zzLB[0][389] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][390] ( .G(n182), .D(idata[358]), .Q(\_zzLB[0][390] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][391] ( .G(n182), .D(idata[359]), .Q(\_zzLB[0][391] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][392] ( .G(n182), .D(idata[360]), .Q(\_zzLB[0][392] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][393] ( .G(n182), .D(idata[361]), .Q(\_zzLB[0][393] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][394] ( .G(n182), .D(idata[362]), .Q(\_zzLB[0][394] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][395] ( .G(n182), .D(idata[363]), .Q(\_zzLB[0][395] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][396] ( .G(n182), .D(idata[364]), .Q(\_zzLB[0][396] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][397] ( .G(n182), .D(idata[365]), .Q(\_zzLB[0][397] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][398] ( .G(n182), .D(idata[366]), .Q(\_zzLB[0][398] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][399] ( .G(n182), .D(idata[367]), .Q(\_zzLB[0][399] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][400] ( .G(n182), .D(idata[368]), .Q(\_zzLB[0][400] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][401] ( .G(n182), .D(idata[369]), .Q(\_zzLB[0][401] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][402] ( .G(n182), .D(idata[370]), .Q(\_zzLB[0][402] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][403] ( .G(n182), .D(idata[371]), .Q(\_zzLB[0][403] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][404] ( .G(n182), .D(idata[372]), .Q(\_zzLB[0][404] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][405] ( .G(n182), .D(idata[373]), .Q(\_zzLB[0][405] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][406] ( .G(n182), .D(idata[374]), .Q(\_zzLB[0][406] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][407] ( .G(n182), .D(idata[375]), .Q(\_zzLB[0][407] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][408] ( .G(n182), .D(idata[376]), .Q(\_zzLB[0][408] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][409] ( .G(n182), .D(idata[377]), .Q(\_zzLB[0][409] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][410] ( .G(n182), .D(idata[378]), .Q(\_zzLB[0][410] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][411] ( .G(n182), .D(idata[379]), .Q(\_zzLB[0][411] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][412] ( .G(n182), .D(idata[380]), .Q(\_zzLB[0][412] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][413] ( .G(n182), .D(idata[381]), .Q(\_zzLB[0][413] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][414] ( .G(n182), .D(idata[382]), .Q(\_zzLB[0][414] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][415] ( .G(n182), .D(idata[383]), .Q(\_zzLB[0][415] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][416] ( .G(n182), .D(idata[384]), .Q(\_zzLB[0][416] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][417] ( .G(n182), .D(idata[385]), .Q(\_zzLB[0][417] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][418] ( .G(n182), .D(idata[386]), .Q(\_zzLB[0][418] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][419] ( .G(n182), .D(idata[387]), .Q(\_zzLB[0][419] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][420] ( .G(n182), .D(idata[388]), .Q(\_zzLB[0][420] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][421] ( .G(n182), .D(idata[389]), .Q(\_zzLB[0][421] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][422] ( .G(n182), .D(idata[390]), .Q(\_zzLB[0][422] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][423] ( .G(n182), .D(idata[391]), .Q(\_zzLB[0][423] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][424] ( .G(n182), .D(idata[392]), .Q(\_zzLB[0][424] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][425] ( .G(n182), .D(idata[393]), .Q(\_zzLB[0][425] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][426] ( .G(n182), .D(idata[394]), .Q(\_zzLB[0][426] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][427] ( .G(n182), .D(idata[395]), .Q(\_zzLB[0][427] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][428] ( .G(n182), .D(idata[396]), .Q(\_zzLB[0][428] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][429] ( .G(n182), .D(idata[397]), .Q(\_zzLB[0][429] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][430] ( .G(n182), .D(idata[398]), .Q(\_zzLB[0][430] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][431] ( .G(n182), .D(idata[399]), .Q(\_zzLB[0][431] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][432] ( .G(n182), .D(idata[400]), .Q(\_zzLB[0][432] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][433] ( .G(n182), .D(idata[401]), .Q(\_zzLB[0][433] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][434] ( .G(n182), .D(idata[402]), .Q(\_zzLB[0][434] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][435] ( .G(n182), .D(idata[403]), .Q(\_zzLB[0][435] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][436] ( .G(n182), .D(idata[404]), .Q(\_zzLB[0][436] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][437] ( .G(n182), .D(idata[405]), .Q(\_zzLB[0][437] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][438] ( .G(n182), .D(idata[406]), .Q(\_zzLB[0][438] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][439] ( .G(n182), .D(idata[407]), .Q(\_zzLB[0][439] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][440] ( .G(n182), .D(idata[408]), .Q(\_zzLB[0][440] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][441] ( .G(n182), .D(idata[409]), .Q(\_zzLB[0][441] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][442] ( .G(n182), .D(idata[410]), .Q(\_zzLB[0][442] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][443] ( .G(n182), .D(idata[411]), .Q(\_zzLB[0][443] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][444] ( .G(n182), .D(idata[412]), .Q(\_zzLB[0][444] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][445] ( .G(n182), .D(idata[413]), .Q(\_zzLB[0][445] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][446] ( .G(n182), .D(idata[414]), .Q(\_zzLB[0][446] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][447] ( .G(n182), .D(idata[415]), .Q(\_zzLB[0][447] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][448] ( .G(n182), .D(idata[416]), .Q(\_zzLB[0][448] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][449] ( .G(n182), .D(idata[417]), .Q(\_zzLB[0][449] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][450] ( .G(n182), .D(idata[418]), .Q(\_zzLB[0][450] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][451] ( .G(n182), .D(idata[419]), .Q(\_zzLB[0][451] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][452] ( .G(n182), .D(idata[420]), .Q(\_zzLB[0][452] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][453] ( .G(n182), .D(idata[421]), .Q(\_zzLB[0][453] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][454] ( .G(n182), .D(idata[422]), .Q(\_zzLB[0][454] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][455] ( .G(n182), .D(idata[423]), .Q(\_zzLB[0][455] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][456] ( .G(n182), .D(idata[424]), .Q(\_zzLB[0][456] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][457] ( .G(n182), .D(idata[425]), .Q(\_zzLB[0][457] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][458] ( .G(n182), .D(idata[426]), .Q(\_zzLB[0][458] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][459] ( .G(n182), .D(idata[427]), .Q(\_zzLB[0][459] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][460] ( .G(n182), .D(idata[428]), .Q(\_zzLB[0][460] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][461] ( .G(n182), .D(idata[429]), .Q(\_zzLB[0][461] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][462] ( .G(n182), .D(idata[430]), .Q(\_zzLB[0][462] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][463] ( .G(n182), .D(idata[431]), .Q(\_zzLB[0][463] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][464] ( .G(n182), .D(idata[432]), .Q(\_zzLB[0][464] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][465] ( .G(n182), .D(idata[433]), .Q(\_zzLB[0][465] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][466] ( .G(n182), .D(idata[434]), .Q(\_zzLB[0][466] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][467] ( .G(n182), .D(idata[435]), .Q(\_zzLB[0][467] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][468] ( .G(n182), .D(idata[436]), .Q(\_zzLB[0][468] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][469] ( .G(n182), .D(idata[437]), .Q(\_zzLB[0][469] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][470] ( .G(n182), .D(idata[438]), .Q(\_zzLB[0][470] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][471] ( .G(n182), .D(idata[439]), .Q(\_zzLB[0][471] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][472] ( .G(n182), .D(idata[440]), .Q(\_zzLB[0][472] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][473] ( .G(n182), .D(idata[441]), .Q(\_zzLB[0][473] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][474] ( .G(n182), .D(idata[442]), .Q(\_zzLB[0][474] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][475] ( .G(n182), .D(idata[443]), .Q(\_zzLB[0][475] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][476] ( .G(n182), .D(idata[444]), .Q(\_zzLB[0][476] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][477] ( .G(n182), .D(idata[445]), .Q(\_zzLB[0][477] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][478] ( .G(n182), .D(idata[446]), .Q(\_zzLB[0][478] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][479] ( .G(n182), .D(idata[447]), .Q(\_zzLB[0][479] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][480] ( .G(n182), .D(idata[448]), .Q(\_zzLB[0][480] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][481] ( .G(n182), .D(idata[449]), .Q(\_zzLB[0][481] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][482] ( .G(n182), .D(idata[450]), .Q(\_zzLB[0][482] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][483] ( .G(n182), .D(idata[451]), .Q(\_zzLB[0][483] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][484] ( .G(n182), .D(idata[452]), .Q(\_zzLB[0][484] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][485] ( .G(n182), .D(idata[453]), .Q(\_zzLB[0][485] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][486] ( .G(n182), .D(idata[454]), .Q(\_zzLB[0][486] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][487] ( .G(n182), .D(idata[455]), .Q(\_zzLB[0][487] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][488] ( .G(n182), .D(idata[456]), .Q(\_zzLB[0][488] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][489] ( .G(n182), .D(idata[457]), .Q(\_zzLB[0][489] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][490] ( .G(n182), .D(idata[458]), .Q(\_zzLB[0][490] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][491] ( .G(n182), .D(idata[459]), .Q(\_zzLB[0][491] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][492] ( .G(n182), .D(idata[460]), .Q(\_zzLB[0][492] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][493] ( .G(n182), .D(idata[461]), .Q(\_zzLB[0][493] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][494] ( .G(n182), .D(idata[462]), .Q(\_zzLB[0][494] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][495] ( .G(n182), .D(idata[463]), .Q(\_zzLB[0][495] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][496] ( .G(n182), .D(idata[464]), .Q(\_zzLB[0][496] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][497] ( .G(n182), .D(idata[465]), .Q(\_zzLB[0][497] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][498] ( .G(n182), .D(idata[466]), .Q(\_zzLB[0][498] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][499] ( .G(n182), .D(idata[467]), .Q(\_zzLB[0][499] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][500] ( .G(n182), .D(idata[468]), .Q(\_zzLB[0][500] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][501] ( .G(n182), .D(idata[469]), .Q(\_zzLB[0][501] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][502] ( .G(n182), .D(idata[470]), .Q(\_zzLB[0][502] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][503] ( .G(n182), .D(idata[471]), .Q(\_zzLB[0][503] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][504] ( .G(n182), .D(idata[472]), .Q(\_zzLB[0][504] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][505] ( .G(n182), .D(idata[473]), .Q(\_zzLB[0][505] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][506] ( .G(n182), .D(idata[474]), .Q(\_zzLB[0][506] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][507] ( .G(n182), .D(idata[475]), .Q(\_zzLB[0][507] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][508] ( .G(n182), .D(idata[476]), .Q(\_zzLB[0][508] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][509] ( .G(n182), .D(idata[477]), .Q(\_zzLB[0][509] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][510] ( .G(n182), .D(idata[478]), .Q(\_zzLB[0][510] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][511] ( .G(n182), .D(idata[479]), .Q(\_zzLB[0][511] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][512] ( .G(n182), .D(idata[480]), .Q(\_zzLB[0][512] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][513] ( .G(n182), .D(idata[481]), .Q(\_zzLB[0][513] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][514] ( .G(n182), .D(idata[482]), .Q(\_zzLB[0][514] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][515] ( .G(n182), .D(idata[483]), .Q(\_zzLB[0][515] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][516] ( .G(n182), .D(idata[484]), .Q(\_zzLB[0][516] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][517] ( .G(n182), .D(idata[485]), .Q(\_zzLB[0][517] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][518] ( .G(n182), .D(idata[486]), .Q(\_zzLB[0][518] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][519] ( .G(n182), .D(idata[487]), .Q(\_zzLB[0][519] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][520] ( .G(n182), .D(idata[488]), .Q(\_zzLB[0][520] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][521] ( .G(n182), .D(idata[489]), .Q(\_zzLB[0][521] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][522] ( .G(n182), .D(idata[490]), .Q(\_zzLB[0][522] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][523] ( .G(n182), .D(idata[491]), .Q(\_zzLB[0][523] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][524] ( .G(n182), .D(idata[492]), .Q(\_zzLB[0][524] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][525] ( .G(n182), .D(idata[493]), .Q(\_zzLB[0][525] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][526] ( .G(n182), .D(idata[494]), .Q(\_zzLB[0][526] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][527] ( .G(n182), .D(idata[495]), .Q(\_zzLB[0][527] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][528] ( .G(n182), .D(idata[496]), .Q(\_zzLB[0][528] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][529] ( .G(n182), .D(idata[497]), .Q(\_zzLB[0][529] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][530] ( .G(n182), .D(idata[498]), .Q(\_zzLB[0][530] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][531] ( .G(n182), .D(idata[499]), .Q(\_zzLB[0][531] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][532] ( .G(n182), .D(idata[500]), .Q(\_zzLB[0][532] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][533] ( .G(n182), .D(idata[501]), .Q(\_zzLB[0][533] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][534] ( .G(n182), .D(idata[502]), .Q(\_zzLB[0][534] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][535] ( .G(n182), .D(idata[503]), .Q(\_zzLB[0][535] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][536] ( .G(n182), .D(idata[504]), .Q(\_zzLB[0][536] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][537] ( .G(n182), .D(idata[505]), .Q(\_zzLB[0][537] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][538] ( .G(n182), .D(idata[506]), .Q(\_zzLB[0][538] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][539] ( .G(n182), .D(idata[507]), .Q(\_zzLB[0][539] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][540] ( .G(n182), .D(idata[508]), .Q(\_zzLB[0][540] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][541] ( .G(n182), .D(idata[509]), .Q(\_zzLB[0][541] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][542] ( .G(n182), .D(idata[510]), .Q(\_zzLB[0][542] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][543] ( .G(n182), .D(idata[511]), .Q(\_zzLB[0][543] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][544] ( .G(n182), .D(idata[512]), .Q(\_zzLB[0][544] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][545] ( .G(n182), .D(idata[513]), .Q(\_zzLB[0][545] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][546] ( .G(n182), .D(idata[514]), .Q(\_zzLB[0][546] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][547] ( .G(n182), .D(idata[515]), .Q(\_zzLB[0][547] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][548] ( .G(n182), .D(idata[516]), .Q(\_zzLB[0][548] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][549] ( .G(n182), .D(idata[517]), .Q(\_zzLB[0][549] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][550] ( .G(n182), .D(idata[518]), .Q(\_zzLB[0][550] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][551] ( .G(n182), .D(idata[519]), .Q(\_zzLB[0][551] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][552] ( .G(n182), .D(idata[520]), .Q(\_zzLB[0][552] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][553] ( .G(n182), .D(idata[521]), .Q(\_zzLB[0][553] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][554] ( .G(n182), .D(idata[522]), .Q(\_zzLB[0][554] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][555] ( .G(n182), .D(idata[523]), .Q(\_zzLB[0][555] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][556] ( .G(n182), .D(idata[524]), .Q(\_zzLB[0][556] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][557] ( .G(n182), .D(idata[525]), .Q(\_zzLB[0][557] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][558] ( .G(n182), .D(idata[526]), .Q(\_zzLB[0][558] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][559] ( .G(n182), .D(idata[527]), .Q(\_zzLB[0][559] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][560] ( .G(n182), .D(idata[528]), .Q(\_zzLB[0][560] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][561] ( .G(n182), .D(idata[529]), .Q(\_zzLB[0][561] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][562] ( .G(n182), .D(idata[530]), .Q(\_zzLB[0][562] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][563] ( .G(n182), .D(idata[531]), .Q(\_zzLB[0][563] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][564] ( .G(n182), .D(idata[532]), .Q(\_zzLB[0][564] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][565] ( .G(n182), .D(idata[533]), .Q(\_zzLB[0][565] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][566] ( .G(n182), .D(idata[534]), .Q(\_zzLB[0][566] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][567] ( .G(n182), .D(idata[535]), .Q(\_zzLB[0][567] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][568] ( .G(n182), .D(idata[536]), .Q(\_zzLB[0][568] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][569] ( .G(n182), .D(idata[537]), .Q(\_zzLB[0][569] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][570] ( .G(n182), .D(idata[538]), .Q(\_zzLB[0][570] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][571] ( .G(n182), .D(idata[539]), .Q(\_zzLB[0][571] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][572] ( .G(n182), .D(idata[540]), .Q(\_zzLB[0][572] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][573] ( .G(n182), .D(idata[541]), .Q(\_zzLB[0][573] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][574] ( .G(n182), .D(idata[542]), .Q(\_zzLB[0][574] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][575] ( .G(n182), .D(idata[543]), .Q(\_zzLB[0][575] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][576] ( .G(n182), .D(idata[544]), .Q(\_zzLB[0][576] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][577] ( .G(n182), .D(idata[545]), .Q(\_zzLB[0][577] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][578] ( .G(n182), .D(idata[546]), .Q(\_zzLB[0][578] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][579] ( .G(n182), .D(idata[547]), .Q(\_zzLB[0][579] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][580] ( .G(n182), .D(idata[548]), .Q(\_zzLB[0][580] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][581] ( .G(n182), .D(idata[549]), .Q(\_zzLB[0][581] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][582] ( .G(n182), .D(idata[550]), .Q(\_zzLB[0][582] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][583] ( .G(n182), .D(idata[551]), .Q(\_zzLB[0][583] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][584] ( .G(n182), .D(idata[552]), .Q(\_zzLB[0][584] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][585] ( .G(n182), .D(idata[553]), .Q(\_zzLB[0][585] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][586] ( .G(n182), .D(idata[554]), .Q(\_zzLB[0][586] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][587] ( .G(n182), .D(idata[555]), .Q(\_zzLB[0][587] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][588] ( .G(n182), .D(idata[556]), .Q(\_zzLB[0][588] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][589] ( .G(n182), .D(idata[557]), .Q(\_zzLB[0][589] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][590] ( .G(n182), .D(idata[558]), .Q(\_zzLB[0][590] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][591] ( .G(n182), .D(idata[559]), .Q(\_zzLB[0][591] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][592] ( .G(n182), .D(ireq), .Q(\_zzLB[0][592] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][0] ( .G(n179), .D(len[0]), .Q(\_zzLB[1][0] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][1] ( .G(n179), .D(len[1]), .Q(\_zzLB[1][1] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][2] ( .G(n179), .D(len[2]), .Q(\_zzLB[1][2] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][3] ( .G(n179), .D(len[3]), .Q(\_zzLB[1][3] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][4] ( .G(n179), .D(len[4]), .Q(\_zzLB[1][4] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][5] ( .G(n179), .D(len[5]), .Q(\_zzLB[1][5] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][6] ( .G(n179), .D(len[6]), .Q(\_zzLB[1][6] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][7] ( .G(n179), .D(len[7]), .Q(\_zzLB[1][7] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][8] ( .G(n179), .D(len[8]), .Q(\_zzLB[1][8] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][9] ( .G(n179), .D(len[9]), .Q(\_zzLB[1][9] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][10] ( .G(n179), .D(len[10]), .Q(\_zzLB[1][10] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][11] ( .G(n179), .D(len[11]), .Q(\_zzLB[1][11] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][12] ( .G(n179), .D(cbid[0]), .Q(\_zzLB[1][12] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][13] ( .G(n179), .D(cbid[1]), .Q(\_zzLB[1][13] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][14] ( .G(n179), .D(cbid[2]), .Q(\_zzLB[1][14] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][15] ( .G(n179), .D(cbid[3]), .Q(\_zzLB[1][15] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][16] ( .G(n179), .D(cbid[4]), .Q(\_zzLB[1][16] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][17] ( .G(n179), .D(cbid[5]), .Q(\_zzLB[1][17] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][18] ( .G(n179), .D(cbid[6]), .Q(\_zzLB[1][18] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][19] ( .G(n179), .D(cbid[7]), .Q(\_zzLB[1][19] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][20] ( .G(n179), .D(cbid[8]), .Q(\_zzLB[1][20] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][21] ( .G(n179), .D(cbid[9]), .Q(\_zzLB[1][21] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][22] ( .G(n179), .D(cbid[10]), .Q(\_zzLB[1][22] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][23] ( .G(n179), .D(cbid[11]), .Q(\_zzLB[1][23] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][24] ( .G(n179), .D(cbid[12]), .Q(\_zzLB[1][24] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][25] ( .G(n179), .D(cbid[13]), .Q(\_zzLB[1][25] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][26] ( .G(n179), .D(cbid[14]), .Q(\_zzLB[1][26] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][27] ( .G(n179), .D(cbid[15]), .Q(\_zzLB[1][27] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][28] ( .G(n179), .D(cbid[16]), .Q(\_zzLB[1][28] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][29] ( .G(n179), .D(cbid[17]), .Q(\_zzLB[1][29] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][30] ( .G(n179), .D(cbid[18]), .Q(\_zzLB[1][30] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][31] ( .G(n179), .D(cbid[19]), .Q(\_zzLB[1][31] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][32] ( .G(n179), .D(idata[0]), .Q(\_zzLB[1][32] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][33] ( .G(n179), .D(idata[1]), .Q(\_zzLB[1][33] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][34] ( .G(n179), .D(idata[2]), .Q(\_zzLB[1][34] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][35] ( .G(n179), .D(idata[3]), .Q(\_zzLB[1][35] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][36] ( .G(n179), .D(idata[4]), .Q(\_zzLB[1][36] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][37] ( .G(n179), .D(idata[5]), .Q(\_zzLB[1][37] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][38] ( .G(n179), .D(idata[6]), .Q(\_zzLB[1][38] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][39] ( .G(n179), .D(idata[7]), .Q(\_zzLB[1][39] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][40] ( .G(n179), .D(idata[8]), .Q(\_zzLB[1][40] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][41] ( .G(n179), .D(idata[9]), .Q(\_zzLB[1][41] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][42] ( .G(n179), .D(idata[10]), .Q(\_zzLB[1][42] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][43] ( .G(n179), .D(idata[11]), .Q(\_zzLB[1][43] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][44] ( .G(n179), .D(idata[12]), .Q(\_zzLB[1][44] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][45] ( .G(n179), .D(idata[13]), .Q(\_zzLB[1][45] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][46] ( .G(n179), .D(idata[14]), .Q(\_zzLB[1][46] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][47] ( .G(n179), .D(idata[15]), .Q(\_zzLB[1][47] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][48] ( .G(n179), .D(idata[16]), .Q(\_zzLB[1][48] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][49] ( .G(n179), .D(idata[17]), .Q(\_zzLB[1][49] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][50] ( .G(n179), .D(idata[18]), .Q(\_zzLB[1][50] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][51] ( .G(n179), .D(idata[19]), .Q(\_zzLB[1][51] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][52] ( .G(n179), .D(idata[20]), .Q(\_zzLB[1][52] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][53] ( .G(n179), .D(idata[21]), .Q(\_zzLB[1][53] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][54] ( .G(n179), .D(idata[22]), .Q(\_zzLB[1][54] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][55] ( .G(n179), .D(idata[23]), .Q(\_zzLB[1][55] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][56] ( .G(n179), .D(idata[24]), .Q(\_zzLB[1][56] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][57] ( .G(n179), .D(idata[25]), .Q(\_zzLB[1][57] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][58] ( .G(n179), .D(idata[26]), .Q(\_zzLB[1][58] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][59] ( .G(n179), .D(idata[27]), .Q(\_zzLB[1][59] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][60] ( .G(n179), .D(idata[28]), .Q(\_zzLB[1][60] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][61] ( .G(n179), .D(idata[29]), .Q(\_zzLB[1][61] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][62] ( .G(n179), .D(idata[30]), .Q(\_zzLB[1][62] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][63] ( .G(n179), .D(idata[31]), .Q(\_zzLB[1][63] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][64] ( .G(n179), .D(idata[32]), .Q(\_zzLB[1][64] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][65] ( .G(n179), .D(idata[33]), .Q(\_zzLB[1][65] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][66] ( .G(n179), .D(idata[34]), .Q(\_zzLB[1][66] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][67] ( .G(n179), .D(idata[35]), .Q(\_zzLB[1][67] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][68] ( .G(n179), .D(idata[36]), .Q(\_zzLB[1][68] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][69] ( .G(n179), .D(idata[37]), .Q(\_zzLB[1][69] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][70] ( .G(n179), .D(idata[38]), .Q(\_zzLB[1][70] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][71] ( .G(n179), .D(idata[39]), .Q(\_zzLB[1][71] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][72] ( .G(n179), .D(idata[40]), .Q(\_zzLB[1][72] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][73] ( .G(n179), .D(idata[41]), .Q(\_zzLB[1][73] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][74] ( .G(n179), .D(idata[42]), .Q(\_zzLB[1][74] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][75] ( .G(n179), .D(idata[43]), .Q(\_zzLB[1][75] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][76] ( .G(n179), .D(idata[44]), .Q(\_zzLB[1][76] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][77] ( .G(n179), .D(idata[45]), .Q(\_zzLB[1][77] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][78] ( .G(n179), .D(idata[46]), .Q(\_zzLB[1][78] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][79] ( .G(n179), .D(idata[47]), .Q(\_zzLB[1][79] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][80] ( .G(n179), .D(idata[48]), .Q(\_zzLB[1][80] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][81] ( .G(n179), .D(idata[49]), .Q(\_zzLB[1][81] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][82] ( .G(n179), .D(idata[50]), .Q(\_zzLB[1][82] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][83] ( .G(n179), .D(idata[51]), .Q(\_zzLB[1][83] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][84] ( .G(n179), .D(idata[52]), .Q(\_zzLB[1][84] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][85] ( .G(n179), .D(idata[53]), .Q(\_zzLB[1][85] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][86] ( .G(n179), .D(idata[54]), .Q(\_zzLB[1][86] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][87] ( .G(n179), .D(idata[55]), .Q(\_zzLB[1][87] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][88] ( .G(n179), .D(idata[56]), .Q(\_zzLB[1][88] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][89] ( .G(n179), .D(idata[57]), .Q(\_zzLB[1][89] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][90] ( .G(n179), .D(idata[58]), .Q(\_zzLB[1][90] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][91] ( .G(n179), .D(idata[59]), .Q(\_zzLB[1][91] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][92] ( .G(n179), .D(idata[60]), .Q(\_zzLB[1][92] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][93] ( .G(n179), .D(idata[61]), .Q(\_zzLB[1][93] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][94] ( .G(n179), .D(idata[62]), .Q(\_zzLB[1][94] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][95] ( .G(n179), .D(idata[63]), .Q(\_zzLB[1][95] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][96] ( .G(n179), .D(idata[64]), .Q(\_zzLB[1][96] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][97] ( .G(n179), .D(idata[65]), .Q(\_zzLB[1][97] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][98] ( .G(n179), .D(idata[66]), .Q(\_zzLB[1][98] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][99] ( .G(n179), .D(idata[67]), .Q(\_zzLB[1][99] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][100] ( .G(n179), .D(idata[68]), .Q(\_zzLB[1][100] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][101] ( .G(n179), .D(idata[69]), .Q(\_zzLB[1][101] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][102] ( .G(n179), .D(idata[70]), .Q(\_zzLB[1][102] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][103] ( .G(n179), .D(idata[71]), .Q(\_zzLB[1][103] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][104] ( .G(n179), .D(idata[72]), .Q(\_zzLB[1][104] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][105] ( .G(n179), .D(idata[73]), .Q(\_zzLB[1][105] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][106] ( .G(n179), .D(idata[74]), .Q(\_zzLB[1][106] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][107] ( .G(n179), .D(idata[75]), .Q(\_zzLB[1][107] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][108] ( .G(n179), .D(idata[76]), .Q(\_zzLB[1][108] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][109] ( .G(n179), .D(idata[77]), .Q(\_zzLB[1][109] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][110] ( .G(n179), .D(idata[78]), .Q(\_zzLB[1][110] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][111] ( .G(n179), .D(idata[79]), .Q(\_zzLB[1][111] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][112] ( .G(n179), .D(idata[80]), .Q(\_zzLB[1][112] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][113] ( .G(n179), .D(idata[81]), .Q(\_zzLB[1][113] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][114] ( .G(n179), .D(idata[82]), .Q(\_zzLB[1][114] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][115] ( .G(n179), .D(idata[83]), .Q(\_zzLB[1][115] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][116] ( .G(n179), .D(idata[84]), .Q(\_zzLB[1][116] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][117] ( .G(n179), .D(idata[85]), .Q(\_zzLB[1][117] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][118] ( .G(n179), .D(idata[86]), .Q(\_zzLB[1][118] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][119] ( .G(n179), .D(idata[87]), .Q(\_zzLB[1][119] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][120] ( .G(n179), .D(idata[88]), .Q(\_zzLB[1][120] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][121] ( .G(n179), .D(idata[89]), .Q(\_zzLB[1][121] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][122] ( .G(n179), .D(idata[90]), .Q(\_zzLB[1][122] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][123] ( .G(n179), .D(idata[91]), .Q(\_zzLB[1][123] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][124] ( .G(n179), .D(idata[92]), .Q(\_zzLB[1][124] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][125] ( .G(n179), .D(idata[93]), .Q(\_zzLB[1][125] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][126] ( .G(n179), .D(idata[94]), .Q(\_zzLB[1][126] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][127] ( .G(n179), .D(idata[95]), .Q(\_zzLB[1][127] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][128] ( .G(n179), .D(idata[96]), .Q(\_zzLB[1][128] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][129] ( .G(n179), .D(idata[97]), .Q(\_zzLB[1][129] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][130] ( .G(n179), .D(idata[98]), .Q(\_zzLB[1][130] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][131] ( .G(n179), .D(idata[99]), .Q(\_zzLB[1][131] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][132] ( .G(n179), .D(idata[100]), .Q(\_zzLB[1][132] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][133] ( .G(n179), .D(idata[101]), .Q(\_zzLB[1][133] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][134] ( .G(n179), .D(idata[102]), .Q(\_zzLB[1][134] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][135] ( .G(n179), .D(idata[103]), .Q(\_zzLB[1][135] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][136] ( .G(n179), .D(idata[104]), .Q(\_zzLB[1][136] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][137] ( .G(n179), .D(idata[105]), .Q(\_zzLB[1][137] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][138] ( .G(n179), .D(idata[106]), .Q(\_zzLB[1][138] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][139] ( .G(n179), .D(idata[107]), .Q(\_zzLB[1][139] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][140] ( .G(n179), .D(idata[108]), .Q(\_zzLB[1][140] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][141] ( .G(n179), .D(idata[109]), .Q(\_zzLB[1][141] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][142] ( .G(n179), .D(idata[110]), .Q(\_zzLB[1][142] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][143] ( .G(n179), .D(idata[111]), .Q(\_zzLB[1][143] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][144] ( .G(n179), .D(idata[112]), .Q(\_zzLB[1][144] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][145] ( .G(n179), .D(idata[113]), .Q(\_zzLB[1][145] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][146] ( .G(n179), .D(idata[114]), .Q(\_zzLB[1][146] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][147] ( .G(n179), .D(idata[115]), .Q(\_zzLB[1][147] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][148] ( .G(n179), .D(idata[116]), .Q(\_zzLB[1][148] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][149] ( .G(n179), .D(idata[117]), .Q(\_zzLB[1][149] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][150] ( .G(n179), .D(idata[118]), .Q(\_zzLB[1][150] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][151] ( .G(n179), .D(idata[119]), .Q(\_zzLB[1][151] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][152] ( .G(n179), .D(idata[120]), .Q(\_zzLB[1][152] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][153] ( .G(n179), .D(idata[121]), .Q(\_zzLB[1][153] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][154] ( .G(n179), .D(idata[122]), .Q(\_zzLB[1][154] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][155] ( .G(n179), .D(idata[123]), .Q(\_zzLB[1][155] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][156] ( .G(n179), .D(idata[124]), .Q(\_zzLB[1][156] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][157] ( .G(n179), .D(idata[125]), .Q(\_zzLB[1][157] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][158] ( .G(n179), .D(idata[126]), .Q(\_zzLB[1][158] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][159] ( .G(n179), .D(idata[127]), .Q(\_zzLB[1][159] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][160] ( .G(n179), .D(idata[128]), .Q(\_zzLB[1][160] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][161] ( .G(n179), .D(idata[129]), .Q(\_zzLB[1][161] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][162] ( .G(n179), .D(idata[130]), .Q(\_zzLB[1][162] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][163] ( .G(n179), .D(idata[131]), .Q(\_zzLB[1][163] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][164] ( .G(n179), .D(idata[132]), .Q(\_zzLB[1][164] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][165] ( .G(n179), .D(idata[133]), .Q(\_zzLB[1][165] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][166] ( .G(n179), .D(idata[134]), .Q(\_zzLB[1][166] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][167] ( .G(n179), .D(idata[135]), .Q(\_zzLB[1][167] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][168] ( .G(n179), .D(idata[136]), .Q(\_zzLB[1][168] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][169] ( .G(n179), .D(idata[137]), .Q(\_zzLB[1][169] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][170] ( .G(n179), .D(idata[138]), .Q(\_zzLB[1][170] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][171] ( .G(n179), .D(idata[139]), .Q(\_zzLB[1][171] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][172] ( .G(n179), .D(idata[140]), .Q(\_zzLB[1][172] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][173] ( .G(n179), .D(idata[141]), .Q(\_zzLB[1][173] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][174] ( .G(n179), .D(idata[142]), .Q(\_zzLB[1][174] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][175] ( .G(n179), .D(idata[143]), .Q(\_zzLB[1][175] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][176] ( .G(n179), .D(idata[144]), .Q(\_zzLB[1][176] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][177] ( .G(n179), .D(idata[145]), .Q(\_zzLB[1][177] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][178] ( .G(n179), .D(idata[146]), .Q(\_zzLB[1][178] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][179] ( .G(n179), .D(idata[147]), .Q(\_zzLB[1][179] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][180] ( .G(n179), .D(idata[148]), .Q(\_zzLB[1][180] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][181] ( .G(n179), .D(idata[149]), .Q(\_zzLB[1][181] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][182] ( .G(n179), .D(idata[150]), .Q(\_zzLB[1][182] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][183] ( .G(n179), .D(idata[151]), .Q(\_zzLB[1][183] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][184] ( .G(n179), .D(idata[152]), .Q(\_zzLB[1][184] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][185] ( .G(n179), .D(idata[153]), .Q(\_zzLB[1][185] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][186] ( .G(n179), .D(idata[154]), .Q(\_zzLB[1][186] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][187] ( .G(n179), .D(idata[155]), .Q(\_zzLB[1][187] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][188] ( .G(n179), .D(idata[156]), .Q(\_zzLB[1][188] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][189] ( .G(n179), .D(idata[157]), .Q(\_zzLB[1][189] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][190] ( .G(n179), .D(idata[158]), .Q(\_zzLB[1][190] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][191] ( .G(n179), .D(idata[159]), .Q(\_zzLB[1][191] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][192] ( .G(n179), .D(idata[160]), .Q(\_zzLB[1][192] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][193] ( .G(n179), .D(idata[161]), .Q(\_zzLB[1][193] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][194] ( .G(n179), .D(idata[162]), .Q(\_zzLB[1][194] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][195] ( .G(n179), .D(idata[163]), .Q(\_zzLB[1][195] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][196] ( .G(n179), .D(idata[164]), .Q(\_zzLB[1][196] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][197] ( .G(n179), .D(idata[165]), .Q(\_zzLB[1][197] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][198] ( .G(n179), .D(idata[166]), .Q(\_zzLB[1][198] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][199] ( .G(n179), .D(idata[167]), .Q(\_zzLB[1][199] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][200] ( .G(n179), .D(idata[168]), .Q(\_zzLB[1][200] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][201] ( .G(n179), .D(idata[169]), .Q(\_zzLB[1][201] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][202] ( .G(n179), .D(idata[170]), .Q(\_zzLB[1][202] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][203] ( .G(n179), .D(idata[171]), .Q(\_zzLB[1][203] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][204] ( .G(n179), .D(idata[172]), .Q(\_zzLB[1][204] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][205] ( .G(n179), .D(idata[173]), .Q(\_zzLB[1][205] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][206] ( .G(n179), .D(idata[174]), .Q(\_zzLB[1][206] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][207] ( .G(n179), .D(idata[175]), .Q(\_zzLB[1][207] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][208] ( .G(n179), .D(idata[176]), .Q(\_zzLB[1][208] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][209] ( .G(n179), .D(idata[177]), .Q(\_zzLB[1][209] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][210] ( .G(n179), .D(idata[178]), .Q(\_zzLB[1][210] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][211] ( .G(n179), .D(idata[179]), .Q(\_zzLB[1][211] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][212] ( .G(n179), .D(idata[180]), .Q(\_zzLB[1][212] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][213] ( .G(n179), .D(idata[181]), .Q(\_zzLB[1][213] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][214] ( .G(n179), .D(idata[182]), .Q(\_zzLB[1][214] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][215] ( .G(n179), .D(idata[183]), .Q(\_zzLB[1][215] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][216] ( .G(n179), .D(idata[184]), .Q(\_zzLB[1][216] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][217] ( .G(n179), .D(idata[185]), .Q(\_zzLB[1][217] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][218] ( .G(n179), .D(idata[186]), .Q(\_zzLB[1][218] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][219] ( .G(n179), .D(idata[187]), .Q(\_zzLB[1][219] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][220] ( .G(n179), .D(idata[188]), .Q(\_zzLB[1][220] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][221] ( .G(n179), .D(idata[189]), .Q(\_zzLB[1][221] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][222] ( .G(n179), .D(idata[190]), .Q(\_zzLB[1][222] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][223] ( .G(n179), .D(idata[191]), .Q(\_zzLB[1][223] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][224] ( .G(n179), .D(idata[192]), .Q(\_zzLB[1][224] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][225] ( .G(n179), .D(idata[193]), .Q(\_zzLB[1][225] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][226] ( .G(n179), .D(idata[194]), .Q(\_zzLB[1][226] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][227] ( .G(n179), .D(idata[195]), .Q(\_zzLB[1][227] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][228] ( .G(n179), .D(idata[196]), .Q(\_zzLB[1][228] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][229] ( .G(n179), .D(idata[197]), .Q(\_zzLB[1][229] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][230] ( .G(n179), .D(idata[198]), .Q(\_zzLB[1][230] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][231] ( .G(n179), .D(idata[199]), .Q(\_zzLB[1][231] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][232] ( .G(n179), .D(idata[200]), .Q(\_zzLB[1][232] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][233] ( .G(n179), .D(idata[201]), .Q(\_zzLB[1][233] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][234] ( .G(n179), .D(idata[202]), .Q(\_zzLB[1][234] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][235] ( .G(n179), .D(idata[203]), .Q(\_zzLB[1][235] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][236] ( .G(n179), .D(idata[204]), .Q(\_zzLB[1][236] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][237] ( .G(n179), .D(idata[205]), .Q(\_zzLB[1][237] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][238] ( .G(n179), .D(idata[206]), .Q(\_zzLB[1][238] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][239] ( .G(n179), .D(idata[207]), .Q(\_zzLB[1][239] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][240] ( .G(n179), .D(idata[208]), .Q(\_zzLB[1][240] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][241] ( .G(n179), .D(idata[209]), .Q(\_zzLB[1][241] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][242] ( .G(n179), .D(idata[210]), .Q(\_zzLB[1][242] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][243] ( .G(n179), .D(idata[211]), .Q(\_zzLB[1][243] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][244] ( .G(n179), .D(idata[212]), .Q(\_zzLB[1][244] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][245] ( .G(n179), .D(idata[213]), .Q(\_zzLB[1][245] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][246] ( .G(n179), .D(idata[214]), .Q(\_zzLB[1][246] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][247] ( .G(n179), .D(idata[215]), .Q(\_zzLB[1][247] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][248] ( .G(n179), .D(idata[216]), .Q(\_zzLB[1][248] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][249] ( .G(n179), .D(idata[217]), .Q(\_zzLB[1][249] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][250] ( .G(n179), .D(idata[218]), .Q(\_zzLB[1][250] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][251] ( .G(n179), .D(idata[219]), .Q(\_zzLB[1][251] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][252] ( .G(n179), .D(idata[220]), .Q(\_zzLB[1][252] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][253] ( .G(n179), .D(idata[221]), .Q(\_zzLB[1][253] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][254] ( .G(n179), .D(idata[222]), .Q(\_zzLB[1][254] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][255] ( .G(n179), .D(idata[223]), .Q(\_zzLB[1][255] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][256] ( .G(n179), .D(idata[224]), .Q(\_zzLB[1][256] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][257] ( .G(n179), .D(idata[225]), .Q(\_zzLB[1][257] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][258] ( .G(n179), .D(idata[226]), .Q(\_zzLB[1][258] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][259] ( .G(n179), .D(idata[227]), .Q(\_zzLB[1][259] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][260] ( .G(n179), .D(idata[228]), .Q(\_zzLB[1][260] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][261] ( .G(n179), .D(idata[229]), .Q(\_zzLB[1][261] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][262] ( .G(n179), .D(idata[230]), .Q(\_zzLB[1][262] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][263] ( .G(n179), .D(idata[231]), .Q(\_zzLB[1][263] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][264] ( .G(n179), .D(idata[232]), .Q(\_zzLB[1][264] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][265] ( .G(n179), .D(idata[233]), .Q(\_zzLB[1][265] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][266] ( .G(n179), .D(idata[234]), .Q(\_zzLB[1][266] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][267] ( .G(n179), .D(idata[235]), .Q(\_zzLB[1][267] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][268] ( .G(n179), .D(idata[236]), .Q(\_zzLB[1][268] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][269] ( .G(n179), .D(idata[237]), .Q(\_zzLB[1][269] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][270] ( .G(n179), .D(idata[238]), .Q(\_zzLB[1][270] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][271] ( .G(n179), .D(idata[239]), .Q(\_zzLB[1][271] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][272] ( .G(n179), .D(idata[240]), .Q(\_zzLB[1][272] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][273] ( .G(n179), .D(idata[241]), .Q(\_zzLB[1][273] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][274] ( .G(n179), .D(idata[242]), .Q(\_zzLB[1][274] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][275] ( .G(n179), .D(idata[243]), .Q(\_zzLB[1][275] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][276] ( .G(n179), .D(idata[244]), .Q(\_zzLB[1][276] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][277] ( .G(n179), .D(idata[245]), .Q(\_zzLB[1][277] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][278] ( .G(n179), .D(idata[246]), .Q(\_zzLB[1][278] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][279] ( .G(n179), .D(idata[247]), .Q(\_zzLB[1][279] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][280] ( .G(n179), .D(idata[248]), .Q(\_zzLB[1][280] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][281] ( .G(n179), .D(idata[249]), .Q(\_zzLB[1][281] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][282] ( .G(n179), .D(idata[250]), .Q(\_zzLB[1][282] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][283] ( .G(n179), .D(idata[251]), .Q(\_zzLB[1][283] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][284] ( .G(n179), .D(idata[252]), .Q(\_zzLB[1][284] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][285] ( .G(n179), .D(idata[253]), .Q(\_zzLB[1][285] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][286] ( .G(n179), .D(idata[254]), .Q(\_zzLB[1][286] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][287] ( .G(n179), .D(idata[255]), .Q(\_zzLB[1][287] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][288] ( .G(n179), .D(idata[256]), .Q(\_zzLB[1][288] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][289] ( .G(n179), .D(idata[257]), .Q(\_zzLB[1][289] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][290] ( .G(n179), .D(idata[258]), .Q(\_zzLB[1][290] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][291] ( .G(n179), .D(idata[259]), .Q(\_zzLB[1][291] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][292] ( .G(n179), .D(idata[260]), .Q(\_zzLB[1][292] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][293] ( .G(n179), .D(idata[261]), .Q(\_zzLB[1][293] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][294] ( .G(n179), .D(idata[262]), .Q(\_zzLB[1][294] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][295] ( .G(n179), .D(idata[263]), .Q(\_zzLB[1][295] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][296] ( .G(n179), .D(idata[264]), .Q(\_zzLB[1][296] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][297] ( .G(n179), .D(idata[265]), .Q(\_zzLB[1][297] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][298] ( .G(n179), .D(idata[266]), .Q(\_zzLB[1][298] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][299] ( .G(n179), .D(idata[267]), .Q(\_zzLB[1][299] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][300] ( .G(n179), .D(idata[268]), .Q(\_zzLB[1][300] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][301] ( .G(n179), .D(idata[269]), .Q(\_zzLB[1][301] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][302] ( .G(n179), .D(idata[270]), .Q(\_zzLB[1][302] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][303] ( .G(n179), .D(idata[271]), .Q(\_zzLB[1][303] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][304] ( .G(n179), .D(idata[272]), .Q(\_zzLB[1][304] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][305] ( .G(n179), .D(idata[273]), .Q(\_zzLB[1][305] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][306] ( .G(n179), .D(idata[274]), .Q(\_zzLB[1][306] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][307] ( .G(n179), .D(idata[275]), .Q(\_zzLB[1][307] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][308] ( .G(n179), .D(idata[276]), .Q(\_zzLB[1][308] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][309] ( .G(n179), .D(idata[277]), .Q(\_zzLB[1][309] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][310] ( .G(n179), .D(idata[278]), .Q(\_zzLB[1][310] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][311] ( .G(n179), .D(idata[279]), .Q(\_zzLB[1][311] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][312] ( .G(n179), .D(idata[280]), .Q(\_zzLB[1][312] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][313] ( .G(n179), .D(idata[281]), .Q(\_zzLB[1][313] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][314] ( .G(n179), .D(idata[282]), .Q(\_zzLB[1][314] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][315] ( .G(n179), .D(idata[283]), .Q(\_zzLB[1][315] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][316] ( .G(n179), .D(idata[284]), .Q(\_zzLB[1][316] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][317] ( .G(n179), .D(idata[285]), .Q(\_zzLB[1][317] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][318] ( .G(n179), .D(idata[286]), .Q(\_zzLB[1][318] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][319] ( .G(n179), .D(idata[287]), .Q(\_zzLB[1][319] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][320] ( .G(n179), .D(idata[288]), .Q(\_zzLB[1][320] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][321] ( .G(n179), .D(idata[289]), .Q(\_zzLB[1][321] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][322] ( .G(n179), .D(idata[290]), .Q(\_zzLB[1][322] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][323] ( .G(n179), .D(idata[291]), .Q(\_zzLB[1][323] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][324] ( .G(n179), .D(idata[292]), .Q(\_zzLB[1][324] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][325] ( .G(n179), .D(idata[293]), .Q(\_zzLB[1][325] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][326] ( .G(n179), .D(idata[294]), .Q(\_zzLB[1][326] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][327] ( .G(n179), .D(idata[295]), .Q(\_zzLB[1][327] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][328] ( .G(n179), .D(idata[296]), .Q(\_zzLB[1][328] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][329] ( .G(n179), .D(idata[297]), .Q(\_zzLB[1][329] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][330] ( .G(n179), .D(idata[298]), .Q(\_zzLB[1][330] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][331] ( .G(n179), .D(idata[299]), .Q(\_zzLB[1][331] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][332] ( .G(n179), .D(idata[300]), .Q(\_zzLB[1][332] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][333] ( .G(n179), .D(idata[301]), .Q(\_zzLB[1][333] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][334] ( .G(n179), .D(idata[302]), .Q(\_zzLB[1][334] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][335] ( .G(n179), .D(idata[303]), .Q(\_zzLB[1][335] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][336] ( .G(n179), .D(idata[304]), .Q(\_zzLB[1][336] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][337] ( .G(n179), .D(idata[305]), .Q(\_zzLB[1][337] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][338] ( .G(n179), .D(idata[306]), .Q(\_zzLB[1][338] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][339] ( .G(n179), .D(idata[307]), .Q(\_zzLB[1][339] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][340] ( .G(n179), .D(idata[308]), .Q(\_zzLB[1][340] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][341] ( .G(n179), .D(idata[309]), .Q(\_zzLB[1][341] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][342] ( .G(n179), .D(idata[310]), .Q(\_zzLB[1][342] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][343] ( .G(n179), .D(idata[311]), .Q(\_zzLB[1][343] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][344] ( .G(n179), .D(idata[312]), .Q(\_zzLB[1][344] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][345] ( .G(n179), .D(idata[313]), .Q(\_zzLB[1][345] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][346] ( .G(n179), .D(idata[314]), .Q(\_zzLB[1][346] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][347] ( .G(n179), .D(idata[315]), .Q(\_zzLB[1][347] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][348] ( .G(n179), .D(idata[316]), .Q(\_zzLB[1][348] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][349] ( .G(n179), .D(idata[317]), .Q(\_zzLB[1][349] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][350] ( .G(n179), .D(idata[318]), .Q(\_zzLB[1][350] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][351] ( .G(n179), .D(idata[319]), .Q(\_zzLB[1][351] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][352] ( .G(n179), .D(idata[320]), .Q(\_zzLB[1][352] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][353] ( .G(n179), .D(idata[321]), .Q(\_zzLB[1][353] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][354] ( .G(n179), .D(idata[322]), .Q(\_zzLB[1][354] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][355] ( .G(n179), .D(idata[323]), .Q(\_zzLB[1][355] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][356] ( .G(n179), .D(idata[324]), .Q(\_zzLB[1][356] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][357] ( .G(n179), .D(idata[325]), .Q(\_zzLB[1][357] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][358] ( .G(n179), .D(idata[326]), .Q(\_zzLB[1][358] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][359] ( .G(n179), .D(idata[327]), .Q(\_zzLB[1][359] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][360] ( .G(n179), .D(idata[328]), .Q(\_zzLB[1][360] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][361] ( .G(n179), .D(idata[329]), .Q(\_zzLB[1][361] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][362] ( .G(n179), .D(idata[330]), .Q(\_zzLB[1][362] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][363] ( .G(n179), .D(idata[331]), .Q(\_zzLB[1][363] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][364] ( .G(n179), .D(idata[332]), .Q(\_zzLB[1][364] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][365] ( .G(n179), .D(idata[333]), .Q(\_zzLB[1][365] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][366] ( .G(n179), .D(idata[334]), .Q(\_zzLB[1][366] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][367] ( .G(n179), .D(idata[335]), .Q(\_zzLB[1][367] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][368] ( .G(n179), .D(idata[336]), .Q(\_zzLB[1][368] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][369] ( .G(n179), .D(idata[337]), .Q(\_zzLB[1][369] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][370] ( .G(n179), .D(idata[338]), .Q(\_zzLB[1][370] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][371] ( .G(n179), .D(idata[339]), .Q(\_zzLB[1][371] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][372] ( .G(n179), .D(idata[340]), .Q(\_zzLB[1][372] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][373] ( .G(n179), .D(idata[341]), .Q(\_zzLB[1][373] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][374] ( .G(n179), .D(idata[342]), .Q(\_zzLB[1][374] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][375] ( .G(n179), .D(idata[343]), .Q(\_zzLB[1][375] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][376] ( .G(n179), .D(idata[344]), .Q(\_zzLB[1][376] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][377] ( .G(n179), .D(idata[345]), .Q(\_zzLB[1][377] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][378] ( .G(n179), .D(idata[346]), .Q(\_zzLB[1][378] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][379] ( .G(n179), .D(idata[347]), .Q(\_zzLB[1][379] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][380] ( .G(n179), .D(idata[348]), .Q(\_zzLB[1][380] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][381] ( .G(n179), .D(idata[349]), .Q(\_zzLB[1][381] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][382] ( .G(n179), .D(idata[350]), .Q(\_zzLB[1][382] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][383] ( .G(n179), .D(idata[351]), .Q(\_zzLB[1][383] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][384] ( .G(n179), .D(idata[352]), .Q(\_zzLB[1][384] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][385] ( .G(n179), .D(idata[353]), .Q(\_zzLB[1][385] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][386] ( .G(n179), .D(idata[354]), .Q(\_zzLB[1][386] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][387] ( .G(n179), .D(idata[355]), .Q(\_zzLB[1][387] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][388] ( .G(n179), .D(idata[356]), .Q(\_zzLB[1][388] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][389] ( .G(n179), .D(idata[357]), .Q(\_zzLB[1][389] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][390] ( .G(n179), .D(idata[358]), .Q(\_zzLB[1][390] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][391] ( .G(n179), .D(idata[359]), .Q(\_zzLB[1][391] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][392] ( .G(n179), .D(idata[360]), .Q(\_zzLB[1][392] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][393] ( .G(n179), .D(idata[361]), .Q(\_zzLB[1][393] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][394] ( .G(n179), .D(idata[362]), .Q(\_zzLB[1][394] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][395] ( .G(n179), .D(idata[363]), .Q(\_zzLB[1][395] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][396] ( .G(n179), .D(idata[364]), .Q(\_zzLB[1][396] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][397] ( .G(n179), .D(idata[365]), .Q(\_zzLB[1][397] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][398] ( .G(n179), .D(idata[366]), .Q(\_zzLB[1][398] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][399] ( .G(n179), .D(idata[367]), .Q(\_zzLB[1][399] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][400] ( .G(n179), .D(idata[368]), .Q(\_zzLB[1][400] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][401] ( .G(n179), .D(idata[369]), .Q(\_zzLB[1][401] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][402] ( .G(n179), .D(idata[370]), .Q(\_zzLB[1][402] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][403] ( .G(n179), .D(idata[371]), .Q(\_zzLB[1][403] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][404] ( .G(n179), .D(idata[372]), .Q(\_zzLB[1][404] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][405] ( .G(n179), .D(idata[373]), .Q(\_zzLB[1][405] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][406] ( .G(n179), .D(idata[374]), .Q(\_zzLB[1][406] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][407] ( .G(n179), .D(idata[375]), .Q(\_zzLB[1][407] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][408] ( .G(n179), .D(idata[376]), .Q(\_zzLB[1][408] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][409] ( .G(n179), .D(idata[377]), .Q(\_zzLB[1][409] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][410] ( .G(n179), .D(idata[378]), .Q(\_zzLB[1][410] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][411] ( .G(n179), .D(idata[379]), .Q(\_zzLB[1][411] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][412] ( .G(n179), .D(idata[380]), .Q(\_zzLB[1][412] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][413] ( .G(n179), .D(idata[381]), .Q(\_zzLB[1][413] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][414] ( .G(n179), .D(idata[382]), .Q(\_zzLB[1][414] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][415] ( .G(n179), .D(idata[383]), .Q(\_zzLB[1][415] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][416] ( .G(n179), .D(idata[384]), .Q(\_zzLB[1][416] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][417] ( .G(n179), .D(idata[385]), .Q(\_zzLB[1][417] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][418] ( .G(n179), .D(idata[386]), .Q(\_zzLB[1][418] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][419] ( .G(n179), .D(idata[387]), .Q(\_zzLB[1][419] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][420] ( .G(n179), .D(idata[388]), .Q(\_zzLB[1][420] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][421] ( .G(n179), .D(idata[389]), .Q(\_zzLB[1][421] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][422] ( .G(n179), .D(idata[390]), .Q(\_zzLB[1][422] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][423] ( .G(n179), .D(idata[391]), .Q(\_zzLB[1][423] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][424] ( .G(n179), .D(idata[392]), .Q(\_zzLB[1][424] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][425] ( .G(n179), .D(idata[393]), .Q(\_zzLB[1][425] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][426] ( .G(n179), .D(idata[394]), .Q(\_zzLB[1][426] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][427] ( .G(n179), .D(idata[395]), .Q(\_zzLB[1][427] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][428] ( .G(n179), .D(idata[396]), .Q(\_zzLB[1][428] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][429] ( .G(n179), .D(idata[397]), .Q(\_zzLB[1][429] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][430] ( .G(n179), .D(idata[398]), .Q(\_zzLB[1][430] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][431] ( .G(n179), .D(idata[399]), .Q(\_zzLB[1][431] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][432] ( .G(n179), .D(idata[400]), .Q(\_zzLB[1][432] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][433] ( .G(n179), .D(idata[401]), .Q(\_zzLB[1][433] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][434] ( .G(n179), .D(idata[402]), .Q(\_zzLB[1][434] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][435] ( .G(n179), .D(idata[403]), .Q(\_zzLB[1][435] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][436] ( .G(n179), .D(idata[404]), .Q(\_zzLB[1][436] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][437] ( .G(n179), .D(idata[405]), .Q(\_zzLB[1][437] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][438] ( .G(n179), .D(idata[406]), .Q(\_zzLB[1][438] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][439] ( .G(n179), .D(idata[407]), .Q(\_zzLB[1][439] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][440] ( .G(n179), .D(idata[408]), .Q(\_zzLB[1][440] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][441] ( .G(n179), .D(idata[409]), .Q(\_zzLB[1][441] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][442] ( .G(n179), .D(idata[410]), .Q(\_zzLB[1][442] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][443] ( .G(n179), .D(idata[411]), .Q(\_zzLB[1][443] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][444] ( .G(n179), .D(idata[412]), .Q(\_zzLB[1][444] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][445] ( .G(n179), .D(idata[413]), .Q(\_zzLB[1][445] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][446] ( .G(n179), .D(idata[414]), .Q(\_zzLB[1][446] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][447] ( .G(n179), .D(idata[415]), .Q(\_zzLB[1][447] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][448] ( .G(n179), .D(idata[416]), .Q(\_zzLB[1][448] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][449] ( .G(n179), .D(idata[417]), .Q(\_zzLB[1][449] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][450] ( .G(n179), .D(idata[418]), .Q(\_zzLB[1][450] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][451] ( .G(n179), .D(idata[419]), .Q(\_zzLB[1][451] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][452] ( .G(n179), .D(idata[420]), .Q(\_zzLB[1][452] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][453] ( .G(n179), .D(idata[421]), .Q(\_zzLB[1][453] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][454] ( .G(n179), .D(idata[422]), .Q(\_zzLB[1][454] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][455] ( .G(n179), .D(idata[423]), .Q(\_zzLB[1][455] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][456] ( .G(n179), .D(idata[424]), .Q(\_zzLB[1][456] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][457] ( .G(n179), .D(idata[425]), .Q(\_zzLB[1][457] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][458] ( .G(n179), .D(idata[426]), .Q(\_zzLB[1][458] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][459] ( .G(n179), .D(idata[427]), .Q(\_zzLB[1][459] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][460] ( .G(n179), .D(idata[428]), .Q(\_zzLB[1][460] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][461] ( .G(n179), .D(idata[429]), .Q(\_zzLB[1][461] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][462] ( .G(n179), .D(idata[430]), .Q(\_zzLB[1][462] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][463] ( .G(n179), .D(idata[431]), .Q(\_zzLB[1][463] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][464] ( .G(n179), .D(idata[432]), .Q(\_zzLB[1][464] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][465] ( .G(n179), .D(idata[433]), .Q(\_zzLB[1][465] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][466] ( .G(n179), .D(idata[434]), .Q(\_zzLB[1][466] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][467] ( .G(n179), .D(idata[435]), .Q(\_zzLB[1][467] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][468] ( .G(n179), .D(idata[436]), .Q(\_zzLB[1][468] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][469] ( .G(n179), .D(idata[437]), .Q(\_zzLB[1][469] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][470] ( .G(n179), .D(idata[438]), .Q(\_zzLB[1][470] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][471] ( .G(n179), .D(idata[439]), .Q(\_zzLB[1][471] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][472] ( .G(n179), .D(idata[440]), .Q(\_zzLB[1][472] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][473] ( .G(n179), .D(idata[441]), .Q(\_zzLB[1][473] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][474] ( .G(n179), .D(idata[442]), .Q(\_zzLB[1][474] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][475] ( .G(n179), .D(idata[443]), .Q(\_zzLB[1][475] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][476] ( .G(n179), .D(idata[444]), .Q(\_zzLB[1][476] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][477] ( .G(n179), .D(idata[445]), .Q(\_zzLB[1][477] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][478] ( .G(n179), .D(idata[446]), .Q(\_zzLB[1][478] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][479] ( .G(n179), .D(idata[447]), .Q(\_zzLB[1][479] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][480] ( .G(n179), .D(idata[448]), .Q(\_zzLB[1][480] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][481] ( .G(n179), .D(idata[449]), .Q(\_zzLB[1][481] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][482] ( .G(n179), .D(idata[450]), .Q(\_zzLB[1][482] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][483] ( .G(n179), .D(idata[451]), .Q(\_zzLB[1][483] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][484] ( .G(n179), .D(idata[452]), .Q(\_zzLB[1][484] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][485] ( .G(n179), .D(idata[453]), .Q(\_zzLB[1][485] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][486] ( .G(n179), .D(idata[454]), .Q(\_zzLB[1][486] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][487] ( .G(n179), .D(idata[455]), .Q(\_zzLB[1][487] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][488] ( .G(n179), .D(idata[456]), .Q(\_zzLB[1][488] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][489] ( .G(n179), .D(idata[457]), .Q(\_zzLB[1][489] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][490] ( .G(n179), .D(idata[458]), .Q(\_zzLB[1][490] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][491] ( .G(n179), .D(idata[459]), .Q(\_zzLB[1][491] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][492] ( .G(n179), .D(idata[460]), .Q(\_zzLB[1][492] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][493] ( .G(n179), .D(idata[461]), .Q(\_zzLB[1][493] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][494] ( .G(n179), .D(idata[462]), .Q(\_zzLB[1][494] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][495] ( .G(n179), .D(idata[463]), .Q(\_zzLB[1][495] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][496] ( .G(n179), .D(idata[464]), .Q(\_zzLB[1][496] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][497] ( .G(n179), .D(idata[465]), .Q(\_zzLB[1][497] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][498] ( .G(n179), .D(idata[466]), .Q(\_zzLB[1][498] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][499] ( .G(n179), .D(idata[467]), .Q(\_zzLB[1][499] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][500] ( .G(n179), .D(idata[468]), .Q(\_zzLB[1][500] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][501] ( .G(n179), .D(idata[469]), .Q(\_zzLB[1][501] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][502] ( .G(n179), .D(idata[470]), .Q(\_zzLB[1][502] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][503] ( .G(n179), .D(idata[471]), .Q(\_zzLB[1][503] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][504] ( .G(n179), .D(idata[472]), .Q(\_zzLB[1][504] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][505] ( .G(n179), .D(idata[473]), .Q(\_zzLB[1][505] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][506] ( .G(n179), .D(idata[474]), .Q(\_zzLB[1][506] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][507] ( .G(n179), .D(idata[475]), .Q(\_zzLB[1][507] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][508] ( .G(n179), .D(idata[476]), .Q(\_zzLB[1][508] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][509] ( .G(n179), .D(idata[477]), .Q(\_zzLB[1][509] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][510] ( .G(n179), .D(idata[478]), .Q(\_zzLB[1][510] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][511] ( .G(n179), .D(idata[479]), .Q(\_zzLB[1][511] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][512] ( .G(n179), .D(idata[480]), .Q(\_zzLB[1][512] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][513] ( .G(n179), .D(idata[481]), .Q(\_zzLB[1][513] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][514] ( .G(n179), .D(idata[482]), .Q(\_zzLB[1][514] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][515] ( .G(n179), .D(idata[483]), .Q(\_zzLB[1][515] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][516] ( .G(n179), .D(idata[484]), .Q(\_zzLB[1][516] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][517] ( .G(n179), .D(idata[485]), .Q(\_zzLB[1][517] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][518] ( .G(n179), .D(idata[486]), .Q(\_zzLB[1][518] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][519] ( .G(n179), .D(idata[487]), .Q(\_zzLB[1][519] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][520] ( .G(n179), .D(idata[488]), .Q(\_zzLB[1][520] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][521] ( .G(n179), .D(idata[489]), .Q(\_zzLB[1][521] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][522] ( .G(n179), .D(idata[490]), .Q(\_zzLB[1][522] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][523] ( .G(n179), .D(idata[491]), .Q(\_zzLB[1][523] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][524] ( .G(n179), .D(idata[492]), .Q(\_zzLB[1][524] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][525] ( .G(n179), .D(idata[493]), .Q(\_zzLB[1][525] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][526] ( .G(n179), .D(idata[494]), .Q(\_zzLB[1][526] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][527] ( .G(n179), .D(idata[495]), .Q(\_zzLB[1][527] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][528] ( .G(n179), .D(idata[496]), .Q(\_zzLB[1][528] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][529] ( .G(n179), .D(idata[497]), .Q(\_zzLB[1][529] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][530] ( .G(n179), .D(idata[498]), .Q(\_zzLB[1][530] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][531] ( .G(n179), .D(idata[499]), .Q(\_zzLB[1][531] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][532] ( .G(n179), .D(idata[500]), .Q(\_zzLB[1][532] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][533] ( .G(n179), .D(idata[501]), .Q(\_zzLB[1][533] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][534] ( .G(n179), .D(idata[502]), .Q(\_zzLB[1][534] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][535] ( .G(n179), .D(idata[503]), .Q(\_zzLB[1][535] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][536] ( .G(n179), .D(idata[504]), .Q(\_zzLB[1][536] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][537] ( .G(n179), .D(idata[505]), .Q(\_zzLB[1][537] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][538] ( .G(n179), .D(idata[506]), .Q(\_zzLB[1][538] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][539] ( .G(n179), .D(idata[507]), .Q(\_zzLB[1][539] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][540] ( .G(n179), .D(idata[508]), .Q(\_zzLB[1][540] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][541] ( .G(n179), .D(idata[509]), .Q(\_zzLB[1][541] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][542] ( .G(n179), .D(idata[510]), .Q(\_zzLB[1][542] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][543] ( .G(n179), .D(idata[511]), .Q(\_zzLB[1][543] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][544] ( .G(n179), .D(idata[512]), .Q(\_zzLB[1][544] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][545] ( .G(n179), .D(idata[513]), .Q(\_zzLB[1][545] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][546] ( .G(n179), .D(idata[514]), .Q(\_zzLB[1][546] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][547] ( .G(n179), .D(idata[515]), .Q(\_zzLB[1][547] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][548] ( .G(n179), .D(idata[516]), .Q(\_zzLB[1][548] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][549] ( .G(n179), .D(idata[517]), .Q(\_zzLB[1][549] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][550] ( .G(n179), .D(idata[518]), .Q(\_zzLB[1][550] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][551] ( .G(n179), .D(idata[519]), .Q(\_zzLB[1][551] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][552] ( .G(n179), .D(idata[520]), .Q(\_zzLB[1][552] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][553] ( .G(n179), .D(idata[521]), .Q(\_zzLB[1][553] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][554] ( .G(n179), .D(idata[522]), .Q(\_zzLB[1][554] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][555] ( .G(n179), .D(idata[523]), .Q(\_zzLB[1][555] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][556] ( .G(n179), .D(idata[524]), .Q(\_zzLB[1][556] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][557] ( .G(n179), .D(idata[525]), .Q(\_zzLB[1][557] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][558] ( .G(n179), .D(idata[526]), .Q(\_zzLB[1][558] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][559] ( .G(n179), .D(idata[527]), .Q(\_zzLB[1][559] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][560] ( .G(n179), .D(idata[528]), .Q(\_zzLB[1][560] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][561] ( .G(n179), .D(idata[529]), .Q(\_zzLB[1][561] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][562] ( .G(n179), .D(idata[530]), .Q(\_zzLB[1][562] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][563] ( .G(n179), .D(idata[531]), .Q(\_zzLB[1][563] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][564] ( .G(n179), .D(idata[532]), .Q(\_zzLB[1][564] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][565] ( .G(n179), .D(idata[533]), .Q(\_zzLB[1][565] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][566] ( .G(n179), .D(idata[534]), .Q(\_zzLB[1][566] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][567] ( .G(n179), .D(idata[535]), .Q(\_zzLB[1][567] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][568] ( .G(n179), .D(idata[536]), .Q(\_zzLB[1][568] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][569] ( .G(n179), .D(idata[537]), .Q(\_zzLB[1][569] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][570] ( .G(n179), .D(idata[538]), .Q(\_zzLB[1][570] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][571] ( .G(n179), .D(idata[539]), .Q(\_zzLB[1][571] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][572] ( .G(n179), .D(idata[540]), .Q(\_zzLB[1][572] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][573] ( .G(n179), .D(idata[541]), .Q(\_zzLB[1][573] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][574] ( .G(n179), .D(idata[542]), .Q(\_zzLB[1][574] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][575] ( .G(n179), .D(idata[543]), .Q(\_zzLB[1][575] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][576] ( .G(n179), .D(idata[544]), .Q(\_zzLB[1][576] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][577] ( .G(n179), .D(idata[545]), .Q(\_zzLB[1][577] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][578] ( .G(n179), .D(idata[546]), .Q(\_zzLB[1][578] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][579] ( .G(n179), .D(idata[547]), .Q(\_zzLB[1][579] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][580] ( .G(n179), .D(idata[548]), .Q(\_zzLB[1][580] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][581] ( .G(n179), .D(idata[549]), .Q(\_zzLB[1][581] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][582] ( .G(n179), .D(idata[550]), .Q(\_zzLB[1][582] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][583] ( .G(n179), .D(idata[551]), .Q(\_zzLB[1][583] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][584] ( .G(n179), .D(idata[552]), .Q(\_zzLB[1][584] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][585] ( .G(n179), .D(idata[553]), .Q(\_zzLB[1][585] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][586] ( .G(n179), .D(idata[554]), .Q(\_zzLB[1][586] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][587] ( .G(n179), .D(idata[555]), .Q(\_zzLB[1][587] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][588] ( .G(n179), .D(idata[556]), .Q(\_zzLB[1][588] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][589] ( .G(n179), .D(idata[557]), .Q(\_zzLB[1][589] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][590] ( .G(n179), .D(idata[558]), .Q(\_zzLB[1][590] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][591] ( .G(n179), .D(idata[559]), .Q(\_zzLB[1][591] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][592] ( .G(n179), .D(ireq), .Q(\_zzLB[1][592] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][0] ( .G(n180), .D(len[0]), .Q(\_zzLB[2][0] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][1] ( .G(n180), .D(len[1]), .Q(\_zzLB[2][1] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][2] ( .G(n180), .D(len[2]), .Q(\_zzLB[2][2] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][3] ( .G(n180), .D(len[3]), .Q(\_zzLB[2][3] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][4] ( .G(n180), .D(len[4]), .Q(\_zzLB[2][4] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][5] ( .G(n180), .D(len[5]), .Q(\_zzLB[2][5] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][6] ( .G(n180), .D(len[6]), .Q(\_zzLB[2][6] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][7] ( .G(n180), .D(len[7]), .Q(\_zzLB[2][7] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][8] ( .G(n180), .D(len[8]), .Q(\_zzLB[2][8] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][9] ( .G(n180), .D(len[9]), .Q(\_zzLB[2][9] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][10] ( .G(n180), .D(len[10]), .Q(\_zzLB[2][10] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][11] ( .G(n180), .D(len[11]), .Q(\_zzLB[2][11] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][12] ( .G(n180), .D(cbid[0]), .Q(\_zzLB[2][12] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][13] ( .G(n180), .D(cbid[1]), .Q(\_zzLB[2][13] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][14] ( .G(n180), .D(cbid[2]), .Q(\_zzLB[2][14] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][15] ( .G(n180), .D(cbid[3]), .Q(\_zzLB[2][15] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][16] ( .G(n180), .D(cbid[4]), .Q(\_zzLB[2][16] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][17] ( .G(n180), .D(cbid[5]), .Q(\_zzLB[2][17] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][18] ( .G(n180), .D(cbid[6]), .Q(\_zzLB[2][18] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][19] ( .G(n180), .D(cbid[7]), .Q(\_zzLB[2][19] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][20] ( .G(n180), .D(cbid[8]), .Q(\_zzLB[2][20] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][21] ( .G(n180), .D(cbid[9]), .Q(\_zzLB[2][21] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][22] ( .G(n180), .D(cbid[10]), .Q(\_zzLB[2][22] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][23] ( .G(n180), .D(cbid[11]), .Q(\_zzLB[2][23] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][24] ( .G(n180), .D(cbid[12]), .Q(\_zzLB[2][24] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][25] ( .G(n180), .D(cbid[13]), .Q(\_zzLB[2][25] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][26] ( .G(n180), .D(cbid[14]), .Q(\_zzLB[2][26] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][27] ( .G(n180), .D(cbid[15]), .Q(\_zzLB[2][27] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][28] ( .G(n180), .D(cbid[16]), .Q(\_zzLB[2][28] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][29] ( .G(n180), .D(cbid[17]), .Q(\_zzLB[2][29] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][30] ( .G(n180), .D(cbid[18]), .Q(\_zzLB[2][30] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][31] ( .G(n180), .D(cbid[19]), .Q(\_zzLB[2][31] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][32] ( .G(n180), .D(idata[0]), .Q(\_zzLB[2][32] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][33] ( .G(n180), .D(idata[1]), .Q(\_zzLB[2][33] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][34] ( .G(n180), .D(idata[2]), .Q(\_zzLB[2][34] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][35] ( .G(n180), .D(idata[3]), .Q(\_zzLB[2][35] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][36] ( .G(n180), .D(idata[4]), .Q(\_zzLB[2][36] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][37] ( .G(n180), .D(idata[5]), .Q(\_zzLB[2][37] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][38] ( .G(n180), .D(idata[6]), .Q(\_zzLB[2][38] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][39] ( .G(n180), .D(idata[7]), .Q(\_zzLB[2][39] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][40] ( .G(n180), .D(idata[8]), .Q(\_zzLB[2][40] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][41] ( .G(n180), .D(idata[9]), .Q(\_zzLB[2][41] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][42] ( .G(n180), .D(idata[10]), .Q(\_zzLB[2][42] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][43] ( .G(n180), .D(idata[11]), .Q(\_zzLB[2][43] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][44] ( .G(n180), .D(idata[12]), .Q(\_zzLB[2][44] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][45] ( .G(n180), .D(idata[13]), .Q(\_zzLB[2][45] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][46] ( .G(n180), .D(idata[14]), .Q(\_zzLB[2][46] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][47] ( .G(n180), .D(idata[15]), .Q(\_zzLB[2][47] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][48] ( .G(n180), .D(idata[16]), .Q(\_zzLB[2][48] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][49] ( .G(n180), .D(idata[17]), .Q(\_zzLB[2][49] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][50] ( .G(n180), .D(idata[18]), .Q(\_zzLB[2][50] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][51] ( .G(n180), .D(idata[19]), .Q(\_zzLB[2][51] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][52] ( .G(n180), .D(idata[20]), .Q(\_zzLB[2][52] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][53] ( .G(n180), .D(idata[21]), .Q(\_zzLB[2][53] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][54] ( .G(n180), .D(idata[22]), .Q(\_zzLB[2][54] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][55] ( .G(n180), .D(idata[23]), .Q(\_zzLB[2][55] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][56] ( .G(n180), .D(idata[24]), .Q(\_zzLB[2][56] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][57] ( .G(n180), .D(idata[25]), .Q(\_zzLB[2][57] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][58] ( .G(n180), .D(idata[26]), .Q(\_zzLB[2][58] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][59] ( .G(n180), .D(idata[27]), .Q(\_zzLB[2][59] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][60] ( .G(n180), .D(idata[28]), .Q(\_zzLB[2][60] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][61] ( .G(n180), .D(idata[29]), .Q(\_zzLB[2][61] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][62] ( .G(n180), .D(idata[30]), .Q(\_zzLB[2][62] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][63] ( .G(n180), .D(idata[31]), .Q(\_zzLB[2][63] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][64] ( .G(n180), .D(idata[32]), .Q(\_zzLB[2][64] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][65] ( .G(n180), .D(idata[33]), .Q(\_zzLB[2][65] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][66] ( .G(n180), .D(idata[34]), .Q(\_zzLB[2][66] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][67] ( .G(n180), .D(idata[35]), .Q(\_zzLB[2][67] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][68] ( .G(n180), .D(idata[36]), .Q(\_zzLB[2][68] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][69] ( .G(n180), .D(idata[37]), .Q(\_zzLB[2][69] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][70] ( .G(n180), .D(idata[38]), .Q(\_zzLB[2][70] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][71] ( .G(n180), .D(idata[39]), .Q(\_zzLB[2][71] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][72] ( .G(n180), .D(idata[40]), .Q(\_zzLB[2][72] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][73] ( .G(n180), .D(idata[41]), .Q(\_zzLB[2][73] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][74] ( .G(n180), .D(idata[42]), .Q(\_zzLB[2][74] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][75] ( .G(n180), .D(idata[43]), .Q(\_zzLB[2][75] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][76] ( .G(n180), .D(idata[44]), .Q(\_zzLB[2][76] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][77] ( .G(n180), .D(idata[45]), .Q(\_zzLB[2][77] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][78] ( .G(n180), .D(idata[46]), .Q(\_zzLB[2][78] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][79] ( .G(n180), .D(idata[47]), .Q(\_zzLB[2][79] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][80] ( .G(n180), .D(idata[48]), .Q(\_zzLB[2][80] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][81] ( .G(n180), .D(idata[49]), .Q(\_zzLB[2][81] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][82] ( .G(n180), .D(idata[50]), .Q(\_zzLB[2][82] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][83] ( .G(n180), .D(idata[51]), .Q(\_zzLB[2][83] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][84] ( .G(n180), .D(idata[52]), .Q(\_zzLB[2][84] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][85] ( .G(n180), .D(idata[53]), .Q(\_zzLB[2][85] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][86] ( .G(n180), .D(idata[54]), .Q(\_zzLB[2][86] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][87] ( .G(n180), .D(idata[55]), .Q(\_zzLB[2][87] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][88] ( .G(n180), .D(idata[56]), .Q(\_zzLB[2][88] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][89] ( .G(n180), .D(idata[57]), .Q(\_zzLB[2][89] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][90] ( .G(n180), .D(idata[58]), .Q(\_zzLB[2][90] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][91] ( .G(n180), .D(idata[59]), .Q(\_zzLB[2][91] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][92] ( .G(n180), .D(idata[60]), .Q(\_zzLB[2][92] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][93] ( .G(n180), .D(idata[61]), .Q(\_zzLB[2][93] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][94] ( .G(n180), .D(idata[62]), .Q(\_zzLB[2][94] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][95] ( .G(n180), .D(idata[63]), .Q(\_zzLB[2][95] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][96] ( .G(n180), .D(idata[64]), .Q(\_zzLB[2][96] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][97] ( .G(n180), .D(idata[65]), .Q(\_zzLB[2][97] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][98] ( .G(n180), .D(idata[66]), .Q(\_zzLB[2][98] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][99] ( .G(n180), .D(idata[67]), .Q(\_zzLB[2][99] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][100] ( .G(n180), .D(idata[68]), .Q(\_zzLB[2][100] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][101] ( .G(n180), .D(idata[69]), .Q(\_zzLB[2][101] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][102] ( .G(n180), .D(idata[70]), .Q(\_zzLB[2][102] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][103] ( .G(n180), .D(idata[71]), .Q(\_zzLB[2][103] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][104] ( .G(n180), .D(idata[72]), .Q(\_zzLB[2][104] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][105] ( .G(n180), .D(idata[73]), .Q(\_zzLB[2][105] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][106] ( .G(n180), .D(idata[74]), .Q(\_zzLB[2][106] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][107] ( .G(n180), .D(idata[75]), .Q(\_zzLB[2][107] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][108] ( .G(n180), .D(idata[76]), .Q(\_zzLB[2][108] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][109] ( .G(n180), .D(idata[77]), .Q(\_zzLB[2][109] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][110] ( .G(n180), .D(idata[78]), .Q(\_zzLB[2][110] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][111] ( .G(n180), .D(idata[79]), .Q(\_zzLB[2][111] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][112] ( .G(n180), .D(idata[80]), .Q(\_zzLB[2][112] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][113] ( .G(n180), .D(idata[81]), .Q(\_zzLB[2][113] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][114] ( .G(n180), .D(idata[82]), .Q(\_zzLB[2][114] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][115] ( .G(n180), .D(idata[83]), .Q(\_zzLB[2][115] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][116] ( .G(n180), .D(idata[84]), .Q(\_zzLB[2][116] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][117] ( .G(n180), .D(idata[85]), .Q(\_zzLB[2][117] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][118] ( .G(n180), .D(idata[86]), .Q(\_zzLB[2][118] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][119] ( .G(n180), .D(idata[87]), .Q(\_zzLB[2][119] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][120] ( .G(n180), .D(idata[88]), .Q(\_zzLB[2][120] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][121] ( .G(n180), .D(idata[89]), .Q(\_zzLB[2][121] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][122] ( .G(n180), .D(idata[90]), .Q(\_zzLB[2][122] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][123] ( .G(n180), .D(idata[91]), .Q(\_zzLB[2][123] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][124] ( .G(n180), .D(idata[92]), .Q(\_zzLB[2][124] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][125] ( .G(n180), .D(idata[93]), .Q(\_zzLB[2][125] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][126] ( .G(n180), .D(idata[94]), .Q(\_zzLB[2][126] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][127] ( .G(n180), .D(idata[95]), .Q(\_zzLB[2][127] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][128] ( .G(n180), .D(idata[96]), .Q(\_zzLB[2][128] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][129] ( .G(n180), .D(idata[97]), .Q(\_zzLB[2][129] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][130] ( .G(n180), .D(idata[98]), .Q(\_zzLB[2][130] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][131] ( .G(n180), .D(idata[99]), .Q(\_zzLB[2][131] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][132] ( .G(n180), .D(idata[100]), .Q(\_zzLB[2][132] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][133] ( .G(n180), .D(idata[101]), .Q(\_zzLB[2][133] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][134] ( .G(n180), .D(idata[102]), .Q(\_zzLB[2][134] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][135] ( .G(n180), .D(idata[103]), .Q(\_zzLB[2][135] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][136] ( .G(n180), .D(idata[104]), .Q(\_zzLB[2][136] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][137] ( .G(n180), .D(idata[105]), .Q(\_zzLB[2][137] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][138] ( .G(n180), .D(idata[106]), .Q(\_zzLB[2][138] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][139] ( .G(n180), .D(idata[107]), .Q(\_zzLB[2][139] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][140] ( .G(n180), .D(idata[108]), .Q(\_zzLB[2][140] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][141] ( .G(n180), .D(idata[109]), .Q(\_zzLB[2][141] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][142] ( .G(n180), .D(idata[110]), .Q(\_zzLB[2][142] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][143] ( .G(n180), .D(idata[111]), .Q(\_zzLB[2][143] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][144] ( .G(n180), .D(idata[112]), .Q(\_zzLB[2][144] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][145] ( .G(n180), .D(idata[113]), .Q(\_zzLB[2][145] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][146] ( .G(n180), .D(idata[114]), .Q(\_zzLB[2][146] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][147] ( .G(n180), .D(idata[115]), .Q(\_zzLB[2][147] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][148] ( .G(n180), .D(idata[116]), .Q(\_zzLB[2][148] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][149] ( .G(n180), .D(idata[117]), .Q(\_zzLB[2][149] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][150] ( .G(n180), .D(idata[118]), .Q(\_zzLB[2][150] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][151] ( .G(n180), .D(idata[119]), .Q(\_zzLB[2][151] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][152] ( .G(n180), .D(idata[120]), .Q(\_zzLB[2][152] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][153] ( .G(n180), .D(idata[121]), .Q(\_zzLB[2][153] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][154] ( .G(n180), .D(idata[122]), .Q(\_zzLB[2][154] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][155] ( .G(n180), .D(idata[123]), .Q(\_zzLB[2][155] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][156] ( .G(n180), .D(idata[124]), .Q(\_zzLB[2][156] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][157] ( .G(n180), .D(idata[125]), .Q(\_zzLB[2][157] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][158] ( .G(n180), .D(idata[126]), .Q(\_zzLB[2][158] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][159] ( .G(n180), .D(idata[127]), .Q(\_zzLB[2][159] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][160] ( .G(n180), .D(idata[128]), .Q(\_zzLB[2][160] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][161] ( .G(n180), .D(idata[129]), .Q(\_zzLB[2][161] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][162] ( .G(n180), .D(idata[130]), .Q(\_zzLB[2][162] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][163] ( .G(n180), .D(idata[131]), .Q(\_zzLB[2][163] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][164] ( .G(n180), .D(idata[132]), .Q(\_zzLB[2][164] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][165] ( .G(n180), .D(idata[133]), .Q(\_zzLB[2][165] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][166] ( .G(n180), .D(idata[134]), .Q(\_zzLB[2][166] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][167] ( .G(n180), .D(idata[135]), .Q(\_zzLB[2][167] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][168] ( .G(n180), .D(idata[136]), .Q(\_zzLB[2][168] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][169] ( .G(n180), .D(idata[137]), .Q(\_zzLB[2][169] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][170] ( .G(n180), .D(idata[138]), .Q(\_zzLB[2][170] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][171] ( .G(n180), .D(idata[139]), .Q(\_zzLB[2][171] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][172] ( .G(n180), .D(idata[140]), .Q(\_zzLB[2][172] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][173] ( .G(n180), .D(idata[141]), .Q(\_zzLB[2][173] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][174] ( .G(n180), .D(idata[142]), .Q(\_zzLB[2][174] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][175] ( .G(n180), .D(idata[143]), .Q(\_zzLB[2][175] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][176] ( .G(n180), .D(idata[144]), .Q(\_zzLB[2][176] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][177] ( .G(n180), .D(idata[145]), .Q(\_zzLB[2][177] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][178] ( .G(n180), .D(idata[146]), .Q(\_zzLB[2][178] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][179] ( .G(n180), .D(idata[147]), .Q(\_zzLB[2][179] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][180] ( .G(n180), .D(idata[148]), .Q(\_zzLB[2][180] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][181] ( .G(n180), .D(idata[149]), .Q(\_zzLB[2][181] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][182] ( .G(n180), .D(idata[150]), .Q(\_zzLB[2][182] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][183] ( .G(n180), .D(idata[151]), .Q(\_zzLB[2][183] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][184] ( .G(n180), .D(idata[152]), .Q(\_zzLB[2][184] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][185] ( .G(n180), .D(idata[153]), .Q(\_zzLB[2][185] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][186] ( .G(n180), .D(idata[154]), .Q(\_zzLB[2][186] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][187] ( .G(n180), .D(idata[155]), .Q(\_zzLB[2][187] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][188] ( .G(n180), .D(idata[156]), .Q(\_zzLB[2][188] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][189] ( .G(n180), .D(idata[157]), .Q(\_zzLB[2][189] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][190] ( .G(n180), .D(idata[158]), .Q(\_zzLB[2][190] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][191] ( .G(n180), .D(idata[159]), .Q(\_zzLB[2][191] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][192] ( .G(n180), .D(idata[160]), .Q(\_zzLB[2][192] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][193] ( .G(n180), .D(idata[161]), .Q(\_zzLB[2][193] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][194] ( .G(n180), .D(idata[162]), .Q(\_zzLB[2][194] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][195] ( .G(n180), .D(idata[163]), .Q(\_zzLB[2][195] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][196] ( .G(n180), .D(idata[164]), .Q(\_zzLB[2][196] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][197] ( .G(n180), .D(idata[165]), .Q(\_zzLB[2][197] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][198] ( .G(n180), .D(idata[166]), .Q(\_zzLB[2][198] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][199] ( .G(n180), .D(idata[167]), .Q(\_zzLB[2][199] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][200] ( .G(n180), .D(idata[168]), .Q(\_zzLB[2][200] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][201] ( .G(n180), .D(idata[169]), .Q(\_zzLB[2][201] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][202] ( .G(n180), .D(idata[170]), .Q(\_zzLB[2][202] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][203] ( .G(n180), .D(idata[171]), .Q(\_zzLB[2][203] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][204] ( .G(n180), .D(idata[172]), .Q(\_zzLB[2][204] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][205] ( .G(n180), .D(idata[173]), .Q(\_zzLB[2][205] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][206] ( .G(n180), .D(idata[174]), .Q(\_zzLB[2][206] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][207] ( .G(n180), .D(idata[175]), .Q(\_zzLB[2][207] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][208] ( .G(n180), .D(idata[176]), .Q(\_zzLB[2][208] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][209] ( .G(n180), .D(idata[177]), .Q(\_zzLB[2][209] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][210] ( .G(n180), .D(idata[178]), .Q(\_zzLB[2][210] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][211] ( .G(n180), .D(idata[179]), .Q(\_zzLB[2][211] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][212] ( .G(n180), .D(idata[180]), .Q(\_zzLB[2][212] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][213] ( .G(n180), .D(idata[181]), .Q(\_zzLB[2][213] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][214] ( .G(n180), .D(idata[182]), .Q(\_zzLB[2][214] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][215] ( .G(n180), .D(idata[183]), .Q(\_zzLB[2][215] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][216] ( .G(n180), .D(idata[184]), .Q(\_zzLB[2][216] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][217] ( .G(n180), .D(idata[185]), .Q(\_zzLB[2][217] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][218] ( .G(n180), .D(idata[186]), .Q(\_zzLB[2][218] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][219] ( .G(n180), .D(idata[187]), .Q(\_zzLB[2][219] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][220] ( .G(n180), .D(idata[188]), .Q(\_zzLB[2][220] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][221] ( .G(n180), .D(idata[189]), .Q(\_zzLB[2][221] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][222] ( .G(n180), .D(idata[190]), .Q(\_zzLB[2][222] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][223] ( .G(n180), .D(idata[191]), .Q(\_zzLB[2][223] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][224] ( .G(n180), .D(idata[192]), .Q(\_zzLB[2][224] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][225] ( .G(n180), .D(idata[193]), .Q(\_zzLB[2][225] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][226] ( .G(n180), .D(idata[194]), .Q(\_zzLB[2][226] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][227] ( .G(n180), .D(idata[195]), .Q(\_zzLB[2][227] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][228] ( .G(n180), .D(idata[196]), .Q(\_zzLB[2][228] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][229] ( .G(n180), .D(idata[197]), .Q(\_zzLB[2][229] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][230] ( .G(n180), .D(idata[198]), .Q(\_zzLB[2][230] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][231] ( .G(n180), .D(idata[199]), .Q(\_zzLB[2][231] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][232] ( .G(n180), .D(idata[200]), .Q(\_zzLB[2][232] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][233] ( .G(n180), .D(idata[201]), .Q(\_zzLB[2][233] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][234] ( .G(n180), .D(idata[202]), .Q(\_zzLB[2][234] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][235] ( .G(n180), .D(idata[203]), .Q(\_zzLB[2][235] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][236] ( .G(n180), .D(idata[204]), .Q(\_zzLB[2][236] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][237] ( .G(n180), .D(idata[205]), .Q(\_zzLB[2][237] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][238] ( .G(n180), .D(idata[206]), .Q(\_zzLB[2][238] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][239] ( .G(n180), .D(idata[207]), .Q(\_zzLB[2][239] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][240] ( .G(n180), .D(idata[208]), .Q(\_zzLB[2][240] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][241] ( .G(n180), .D(idata[209]), .Q(\_zzLB[2][241] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][242] ( .G(n180), .D(idata[210]), .Q(\_zzLB[2][242] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][243] ( .G(n180), .D(idata[211]), .Q(\_zzLB[2][243] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][244] ( .G(n180), .D(idata[212]), .Q(\_zzLB[2][244] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][245] ( .G(n180), .D(idata[213]), .Q(\_zzLB[2][245] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][246] ( .G(n180), .D(idata[214]), .Q(\_zzLB[2][246] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][247] ( .G(n180), .D(idata[215]), .Q(\_zzLB[2][247] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][248] ( .G(n180), .D(idata[216]), .Q(\_zzLB[2][248] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][249] ( .G(n180), .D(idata[217]), .Q(\_zzLB[2][249] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][250] ( .G(n180), .D(idata[218]), .Q(\_zzLB[2][250] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][251] ( .G(n180), .D(idata[219]), .Q(\_zzLB[2][251] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][252] ( .G(n180), .D(idata[220]), .Q(\_zzLB[2][252] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][253] ( .G(n180), .D(idata[221]), .Q(\_zzLB[2][253] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][254] ( .G(n180), .D(idata[222]), .Q(\_zzLB[2][254] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][255] ( .G(n180), .D(idata[223]), .Q(\_zzLB[2][255] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][256] ( .G(n180), .D(idata[224]), .Q(\_zzLB[2][256] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][257] ( .G(n180), .D(idata[225]), .Q(\_zzLB[2][257] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][258] ( .G(n180), .D(idata[226]), .Q(\_zzLB[2][258] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][259] ( .G(n180), .D(idata[227]), .Q(\_zzLB[2][259] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][260] ( .G(n180), .D(idata[228]), .Q(\_zzLB[2][260] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][261] ( .G(n180), .D(idata[229]), .Q(\_zzLB[2][261] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][262] ( .G(n180), .D(idata[230]), .Q(\_zzLB[2][262] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][263] ( .G(n180), .D(idata[231]), .Q(\_zzLB[2][263] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][264] ( .G(n180), .D(idata[232]), .Q(\_zzLB[2][264] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][265] ( .G(n180), .D(idata[233]), .Q(\_zzLB[2][265] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][266] ( .G(n180), .D(idata[234]), .Q(\_zzLB[2][266] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][267] ( .G(n180), .D(idata[235]), .Q(\_zzLB[2][267] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][268] ( .G(n180), .D(idata[236]), .Q(\_zzLB[2][268] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][269] ( .G(n180), .D(idata[237]), .Q(\_zzLB[2][269] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][270] ( .G(n180), .D(idata[238]), .Q(\_zzLB[2][270] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][271] ( .G(n180), .D(idata[239]), .Q(\_zzLB[2][271] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][272] ( .G(n180), .D(idata[240]), .Q(\_zzLB[2][272] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][273] ( .G(n180), .D(idata[241]), .Q(\_zzLB[2][273] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][274] ( .G(n180), .D(idata[242]), .Q(\_zzLB[2][274] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][275] ( .G(n180), .D(idata[243]), .Q(\_zzLB[2][275] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][276] ( .G(n180), .D(idata[244]), .Q(\_zzLB[2][276] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][277] ( .G(n180), .D(idata[245]), .Q(\_zzLB[2][277] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][278] ( .G(n180), .D(idata[246]), .Q(\_zzLB[2][278] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][279] ( .G(n180), .D(idata[247]), .Q(\_zzLB[2][279] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][280] ( .G(n180), .D(idata[248]), .Q(\_zzLB[2][280] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][281] ( .G(n180), .D(idata[249]), .Q(\_zzLB[2][281] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][282] ( .G(n180), .D(idata[250]), .Q(\_zzLB[2][282] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][283] ( .G(n180), .D(idata[251]), .Q(\_zzLB[2][283] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][284] ( .G(n180), .D(idata[252]), .Q(\_zzLB[2][284] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][285] ( .G(n180), .D(idata[253]), .Q(\_zzLB[2][285] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][286] ( .G(n180), .D(idata[254]), .Q(\_zzLB[2][286] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][287] ( .G(n180), .D(idata[255]), .Q(\_zzLB[2][287] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][288] ( .G(n180), .D(idata[256]), .Q(\_zzLB[2][288] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][289] ( .G(n180), .D(idata[257]), .Q(\_zzLB[2][289] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][290] ( .G(n180), .D(idata[258]), .Q(\_zzLB[2][290] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][291] ( .G(n180), .D(idata[259]), .Q(\_zzLB[2][291] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][292] ( .G(n180), .D(idata[260]), .Q(\_zzLB[2][292] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][293] ( .G(n180), .D(idata[261]), .Q(\_zzLB[2][293] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][294] ( .G(n180), .D(idata[262]), .Q(\_zzLB[2][294] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][295] ( .G(n180), .D(idata[263]), .Q(\_zzLB[2][295] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][296] ( .G(n180), .D(idata[264]), .Q(\_zzLB[2][296] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][297] ( .G(n180), .D(idata[265]), .Q(\_zzLB[2][297] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][298] ( .G(n180), .D(idata[266]), .Q(\_zzLB[2][298] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][299] ( .G(n180), .D(idata[267]), .Q(\_zzLB[2][299] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][300] ( .G(n180), .D(idata[268]), .Q(\_zzLB[2][300] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][301] ( .G(n180), .D(idata[269]), .Q(\_zzLB[2][301] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][302] ( .G(n180), .D(idata[270]), .Q(\_zzLB[2][302] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][303] ( .G(n180), .D(idata[271]), .Q(\_zzLB[2][303] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][304] ( .G(n180), .D(idata[272]), .Q(\_zzLB[2][304] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][305] ( .G(n180), .D(idata[273]), .Q(\_zzLB[2][305] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][306] ( .G(n180), .D(idata[274]), .Q(\_zzLB[2][306] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][307] ( .G(n180), .D(idata[275]), .Q(\_zzLB[2][307] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][308] ( .G(n180), .D(idata[276]), .Q(\_zzLB[2][308] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][309] ( .G(n180), .D(idata[277]), .Q(\_zzLB[2][309] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][310] ( .G(n180), .D(idata[278]), .Q(\_zzLB[2][310] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][311] ( .G(n180), .D(idata[279]), .Q(\_zzLB[2][311] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][312] ( .G(n180), .D(idata[280]), .Q(\_zzLB[2][312] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][313] ( .G(n180), .D(idata[281]), .Q(\_zzLB[2][313] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][314] ( .G(n180), .D(idata[282]), .Q(\_zzLB[2][314] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][315] ( .G(n180), .D(idata[283]), .Q(\_zzLB[2][315] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][316] ( .G(n180), .D(idata[284]), .Q(\_zzLB[2][316] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][317] ( .G(n180), .D(idata[285]), .Q(\_zzLB[2][317] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][318] ( .G(n180), .D(idata[286]), .Q(\_zzLB[2][318] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][319] ( .G(n180), .D(idata[287]), .Q(\_zzLB[2][319] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][320] ( .G(n180), .D(idata[288]), .Q(\_zzLB[2][320] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][321] ( .G(n180), .D(idata[289]), .Q(\_zzLB[2][321] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][322] ( .G(n180), .D(idata[290]), .Q(\_zzLB[2][322] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][323] ( .G(n180), .D(idata[291]), .Q(\_zzLB[2][323] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][324] ( .G(n180), .D(idata[292]), .Q(\_zzLB[2][324] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][325] ( .G(n180), .D(idata[293]), .Q(\_zzLB[2][325] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][326] ( .G(n180), .D(idata[294]), .Q(\_zzLB[2][326] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][327] ( .G(n180), .D(idata[295]), .Q(\_zzLB[2][327] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][328] ( .G(n180), .D(idata[296]), .Q(\_zzLB[2][328] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][329] ( .G(n180), .D(idata[297]), .Q(\_zzLB[2][329] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][330] ( .G(n180), .D(idata[298]), .Q(\_zzLB[2][330] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][331] ( .G(n180), .D(idata[299]), .Q(\_zzLB[2][331] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][332] ( .G(n180), .D(idata[300]), .Q(\_zzLB[2][332] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][333] ( .G(n180), .D(idata[301]), .Q(\_zzLB[2][333] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][334] ( .G(n180), .D(idata[302]), .Q(\_zzLB[2][334] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][335] ( .G(n180), .D(idata[303]), .Q(\_zzLB[2][335] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][336] ( .G(n180), .D(idata[304]), .Q(\_zzLB[2][336] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][337] ( .G(n180), .D(idata[305]), .Q(\_zzLB[2][337] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][338] ( .G(n180), .D(idata[306]), .Q(\_zzLB[2][338] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][339] ( .G(n180), .D(idata[307]), .Q(\_zzLB[2][339] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][340] ( .G(n180), .D(idata[308]), .Q(\_zzLB[2][340] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][341] ( .G(n180), .D(idata[309]), .Q(\_zzLB[2][341] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][342] ( .G(n180), .D(idata[310]), .Q(\_zzLB[2][342] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][343] ( .G(n180), .D(idata[311]), .Q(\_zzLB[2][343] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][344] ( .G(n180), .D(idata[312]), .Q(\_zzLB[2][344] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][345] ( .G(n180), .D(idata[313]), .Q(\_zzLB[2][345] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][346] ( .G(n180), .D(idata[314]), .Q(\_zzLB[2][346] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][347] ( .G(n180), .D(idata[315]), .Q(\_zzLB[2][347] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][348] ( .G(n180), .D(idata[316]), .Q(\_zzLB[2][348] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][349] ( .G(n180), .D(idata[317]), .Q(\_zzLB[2][349] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][350] ( .G(n180), .D(idata[318]), .Q(\_zzLB[2][350] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][351] ( .G(n180), .D(idata[319]), .Q(\_zzLB[2][351] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][352] ( .G(n180), .D(idata[320]), .Q(\_zzLB[2][352] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][353] ( .G(n180), .D(idata[321]), .Q(\_zzLB[2][353] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][354] ( .G(n180), .D(idata[322]), .Q(\_zzLB[2][354] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][355] ( .G(n180), .D(idata[323]), .Q(\_zzLB[2][355] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][356] ( .G(n180), .D(idata[324]), .Q(\_zzLB[2][356] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][357] ( .G(n180), .D(idata[325]), .Q(\_zzLB[2][357] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][358] ( .G(n180), .D(idata[326]), .Q(\_zzLB[2][358] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][359] ( .G(n180), .D(idata[327]), .Q(\_zzLB[2][359] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][360] ( .G(n180), .D(idata[328]), .Q(\_zzLB[2][360] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][361] ( .G(n180), .D(idata[329]), .Q(\_zzLB[2][361] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][362] ( .G(n180), .D(idata[330]), .Q(\_zzLB[2][362] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][363] ( .G(n180), .D(idata[331]), .Q(\_zzLB[2][363] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][364] ( .G(n180), .D(idata[332]), .Q(\_zzLB[2][364] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][365] ( .G(n180), .D(idata[333]), .Q(\_zzLB[2][365] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][366] ( .G(n180), .D(idata[334]), .Q(\_zzLB[2][366] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][367] ( .G(n180), .D(idata[335]), .Q(\_zzLB[2][367] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][368] ( .G(n180), .D(idata[336]), .Q(\_zzLB[2][368] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][369] ( .G(n180), .D(idata[337]), .Q(\_zzLB[2][369] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][370] ( .G(n180), .D(idata[338]), .Q(\_zzLB[2][370] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][371] ( .G(n180), .D(idata[339]), .Q(\_zzLB[2][371] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][372] ( .G(n180), .D(idata[340]), .Q(\_zzLB[2][372] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][373] ( .G(n180), .D(idata[341]), .Q(\_zzLB[2][373] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][374] ( .G(n180), .D(idata[342]), .Q(\_zzLB[2][374] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][375] ( .G(n180), .D(idata[343]), .Q(\_zzLB[2][375] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][376] ( .G(n180), .D(idata[344]), .Q(\_zzLB[2][376] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][377] ( .G(n180), .D(idata[345]), .Q(\_zzLB[2][377] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][378] ( .G(n180), .D(idata[346]), .Q(\_zzLB[2][378] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][379] ( .G(n180), .D(idata[347]), .Q(\_zzLB[2][379] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][380] ( .G(n180), .D(idata[348]), .Q(\_zzLB[2][380] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][381] ( .G(n180), .D(idata[349]), .Q(\_zzLB[2][381] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][382] ( .G(n180), .D(idata[350]), .Q(\_zzLB[2][382] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][383] ( .G(n180), .D(idata[351]), .Q(\_zzLB[2][383] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][384] ( .G(n180), .D(idata[352]), .Q(\_zzLB[2][384] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][385] ( .G(n180), .D(idata[353]), .Q(\_zzLB[2][385] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][386] ( .G(n180), .D(idata[354]), .Q(\_zzLB[2][386] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][387] ( .G(n180), .D(idata[355]), .Q(\_zzLB[2][387] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][388] ( .G(n180), .D(idata[356]), .Q(\_zzLB[2][388] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][389] ( .G(n180), .D(idata[357]), .Q(\_zzLB[2][389] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][390] ( .G(n180), .D(idata[358]), .Q(\_zzLB[2][390] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][391] ( .G(n180), .D(idata[359]), .Q(\_zzLB[2][391] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][392] ( .G(n180), .D(idata[360]), .Q(\_zzLB[2][392] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][393] ( .G(n180), .D(idata[361]), .Q(\_zzLB[2][393] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][394] ( .G(n180), .D(idata[362]), .Q(\_zzLB[2][394] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][395] ( .G(n180), .D(idata[363]), .Q(\_zzLB[2][395] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][396] ( .G(n180), .D(idata[364]), .Q(\_zzLB[2][396] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][397] ( .G(n180), .D(idata[365]), .Q(\_zzLB[2][397] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][398] ( .G(n180), .D(idata[366]), .Q(\_zzLB[2][398] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][399] ( .G(n180), .D(idata[367]), .Q(\_zzLB[2][399] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][400] ( .G(n180), .D(idata[368]), .Q(\_zzLB[2][400] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][401] ( .G(n180), .D(idata[369]), .Q(\_zzLB[2][401] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][402] ( .G(n180), .D(idata[370]), .Q(\_zzLB[2][402] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][403] ( .G(n180), .D(idata[371]), .Q(\_zzLB[2][403] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][404] ( .G(n180), .D(idata[372]), .Q(\_zzLB[2][404] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][405] ( .G(n180), .D(idata[373]), .Q(\_zzLB[2][405] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][406] ( .G(n180), .D(idata[374]), .Q(\_zzLB[2][406] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][407] ( .G(n180), .D(idata[375]), .Q(\_zzLB[2][407] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][408] ( .G(n180), .D(idata[376]), .Q(\_zzLB[2][408] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][409] ( .G(n180), .D(idata[377]), .Q(\_zzLB[2][409] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][410] ( .G(n180), .D(idata[378]), .Q(\_zzLB[2][410] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][411] ( .G(n180), .D(idata[379]), .Q(\_zzLB[2][411] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][412] ( .G(n180), .D(idata[380]), .Q(\_zzLB[2][412] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][413] ( .G(n180), .D(idata[381]), .Q(\_zzLB[2][413] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][414] ( .G(n180), .D(idata[382]), .Q(\_zzLB[2][414] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][415] ( .G(n180), .D(idata[383]), .Q(\_zzLB[2][415] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][416] ( .G(n180), .D(idata[384]), .Q(\_zzLB[2][416] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][417] ( .G(n180), .D(idata[385]), .Q(\_zzLB[2][417] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][418] ( .G(n180), .D(idata[386]), .Q(\_zzLB[2][418] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][419] ( .G(n180), .D(idata[387]), .Q(\_zzLB[2][419] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][420] ( .G(n180), .D(idata[388]), .Q(\_zzLB[2][420] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][421] ( .G(n180), .D(idata[389]), .Q(\_zzLB[2][421] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][422] ( .G(n180), .D(idata[390]), .Q(\_zzLB[2][422] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][423] ( .G(n180), .D(idata[391]), .Q(\_zzLB[2][423] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][424] ( .G(n180), .D(idata[392]), .Q(\_zzLB[2][424] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][425] ( .G(n180), .D(idata[393]), .Q(\_zzLB[2][425] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][426] ( .G(n180), .D(idata[394]), .Q(\_zzLB[2][426] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][427] ( .G(n180), .D(idata[395]), .Q(\_zzLB[2][427] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][428] ( .G(n180), .D(idata[396]), .Q(\_zzLB[2][428] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][429] ( .G(n180), .D(idata[397]), .Q(\_zzLB[2][429] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][430] ( .G(n180), .D(idata[398]), .Q(\_zzLB[2][430] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][431] ( .G(n180), .D(idata[399]), .Q(\_zzLB[2][431] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][432] ( .G(n180), .D(idata[400]), .Q(\_zzLB[2][432] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][433] ( .G(n180), .D(idata[401]), .Q(\_zzLB[2][433] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][434] ( .G(n180), .D(idata[402]), .Q(\_zzLB[2][434] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][435] ( .G(n180), .D(idata[403]), .Q(\_zzLB[2][435] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][436] ( .G(n180), .D(idata[404]), .Q(\_zzLB[2][436] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][437] ( .G(n180), .D(idata[405]), .Q(\_zzLB[2][437] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][438] ( .G(n180), .D(idata[406]), .Q(\_zzLB[2][438] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][439] ( .G(n180), .D(idata[407]), .Q(\_zzLB[2][439] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][440] ( .G(n180), .D(idata[408]), .Q(\_zzLB[2][440] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][441] ( .G(n180), .D(idata[409]), .Q(\_zzLB[2][441] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][442] ( .G(n180), .D(idata[410]), .Q(\_zzLB[2][442] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][443] ( .G(n180), .D(idata[411]), .Q(\_zzLB[2][443] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][444] ( .G(n180), .D(idata[412]), .Q(\_zzLB[2][444] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][445] ( .G(n180), .D(idata[413]), .Q(\_zzLB[2][445] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][446] ( .G(n180), .D(idata[414]), .Q(\_zzLB[2][446] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][447] ( .G(n180), .D(idata[415]), .Q(\_zzLB[2][447] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][448] ( .G(n180), .D(idata[416]), .Q(\_zzLB[2][448] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][449] ( .G(n180), .D(idata[417]), .Q(\_zzLB[2][449] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][450] ( .G(n180), .D(idata[418]), .Q(\_zzLB[2][450] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][451] ( .G(n180), .D(idata[419]), .Q(\_zzLB[2][451] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][452] ( .G(n180), .D(idata[420]), .Q(\_zzLB[2][452] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][453] ( .G(n180), .D(idata[421]), .Q(\_zzLB[2][453] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][454] ( .G(n180), .D(idata[422]), .Q(\_zzLB[2][454] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][455] ( .G(n180), .D(idata[423]), .Q(\_zzLB[2][455] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][456] ( .G(n180), .D(idata[424]), .Q(\_zzLB[2][456] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][457] ( .G(n180), .D(idata[425]), .Q(\_zzLB[2][457] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][458] ( .G(n180), .D(idata[426]), .Q(\_zzLB[2][458] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][459] ( .G(n180), .D(idata[427]), .Q(\_zzLB[2][459] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][460] ( .G(n180), .D(idata[428]), .Q(\_zzLB[2][460] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][461] ( .G(n180), .D(idata[429]), .Q(\_zzLB[2][461] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][462] ( .G(n180), .D(idata[430]), .Q(\_zzLB[2][462] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][463] ( .G(n180), .D(idata[431]), .Q(\_zzLB[2][463] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][464] ( .G(n180), .D(idata[432]), .Q(\_zzLB[2][464] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][465] ( .G(n180), .D(idata[433]), .Q(\_zzLB[2][465] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][466] ( .G(n180), .D(idata[434]), .Q(\_zzLB[2][466] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][467] ( .G(n180), .D(idata[435]), .Q(\_zzLB[2][467] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][468] ( .G(n180), .D(idata[436]), .Q(\_zzLB[2][468] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][469] ( .G(n180), .D(idata[437]), .Q(\_zzLB[2][469] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][470] ( .G(n180), .D(idata[438]), .Q(\_zzLB[2][470] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][471] ( .G(n180), .D(idata[439]), .Q(\_zzLB[2][471] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][472] ( .G(n180), .D(idata[440]), .Q(\_zzLB[2][472] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][473] ( .G(n180), .D(idata[441]), .Q(\_zzLB[2][473] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][474] ( .G(n180), .D(idata[442]), .Q(\_zzLB[2][474] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][475] ( .G(n180), .D(idata[443]), .Q(\_zzLB[2][475] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][476] ( .G(n180), .D(idata[444]), .Q(\_zzLB[2][476] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][477] ( .G(n180), .D(idata[445]), .Q(\_zzLB[2][477] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][478] ( .G(n180), .D(idata[446]), .Q(\_zzLB[2][478] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][479] ( .G(n180), .D(idata[447]), .Q(\_zzLB[2][479] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][480] ( .G(n180), .D(idata[448]), .Q(\_zzLB[2][480] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][481] ( .G(n180), .D(idata[449]), .Q(\_zzLB[2][481] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][482] ( .G(n180), .D(idata[450]), .Q(\_zzLB[2][482] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][483] ( .G(n180), .D(idata[451]), .Q(\_zzLB[2][483] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][484] ( .G(n180), .D(idata[452]), .Q(\_zzLB[2][484] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][485] ( .G(n180), .D(idata[453]), .Q(\_zzLB[2][485] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][486] ( .G(n180), .D(idata[454]), .Q(\_zzLB[2][486] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][487] ( .G(n180), .D(idata[455]), .Q(\_zzLB[2][487] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][488] ( .G(n180), .D(idata[456]), .Q(\_zzLB[2][488] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][489] ( .G(n180), .D(idata[457]), .Q(\_zzLB[2][489] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][490] ( .G(n180), .D(idata[458]), .Q(\_zzLB[2][490] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][491] ( .G(n180), .D(idata[459]), .Q(\_zzLB[2][491] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][492] ( .G(n180), .D(idata[460]), .Q(\_zzLB[2][492] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][493] ( .G(n180), .D(idata[461]), .Q(\_zzLB[2][493] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][494] ( .G(n180), .D(idata[462]), .Q(\_zzLB[2][494] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][495] ( .G(n180), .D(idata[463]), .Q(\_zzLB[2][495] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][496] ( .G(n180), .D(idata[464]), .Q(\_zzLB[2][496] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][497] ( .G(n180), .D(idata[465]), .Q(\_zzLB[2][497] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][498] ( .G(n180), .D(idata[466]), .Q(\_zzLB[2][498] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][499] ( .G(n180), .D(idata[467]), .Q(\_zzLB[2][499] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][500] ( .G(n180), .D(idata[468]), .Q(\_zzLB[2][500] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][501] ( .G(n180), .D(idata[469]), .Q(\_zzLB[2][501] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][502] ( .G(n180), .D(idata[470]), .Q(\_zzLB[2][502] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][503] ( .G(n180), .D(idata[471]), .Q(\_zzLB[2][503] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][504] ( .G(n180), .D(idata[472]), .Q(\_zzLB[2][504] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][505] ( .G(n180), .D(idata[473]), .Q(\_zzLB[2][505] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][506] ( .G(n180), .D(idata[474]), .Q(\_zzLB[2][506] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][507] ( .G(n180), .D(idata[475]), .Q(\_zzLB[2][507] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][508] ( .G(n180), .D(idata[476]), .Q(\_zzLB[2][508] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][509] ( .G(n180), .D(idata[477]), .Q(\_zzLB[2][509] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][510] ( .G(n180), .D(idata[478]), .Q(\_zzLB[2][510] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][511] ( .G(n180), .D(idata[479]), .Q(\_zzLB[2][511] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][512] ( .G(n180), .D(idata[480]), .Q(\_zzLB[2][512] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][513] ( .G(n180), .D(idata[481]), .Q(\_zzLB[2][513] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][514] ( .G(n180), .D(idata[482]), .Q(\_zzLB[2][514] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][515] ( .G(n180), .D(idata[483]), .Q(\_zzLB[2][515] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][516] ( .G(n180), .D(idata[484]), .Q(\_zzLB[2][516] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][517] ( .G(n180), .D(idata[485]), .Q(\_zzLB[2][517] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][518] ( .G(n180), .D(idata[486]), .Q(\_zzLB[2][518] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][519] ( .G(n180), .D(idata[487]), .Q(\_zzLB[2][519] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][520] ( .G(n180), .D(idata[488]), .Q(\_zzLB[2][520] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][521] ( .G(n180), .D(idata[489]), .Q(\_zzLB[2][521] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][522] ( .G(n180), .D(idata[490]), .Q(\_zzLB[2][522] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][523] ( .G(n180), .D(idata[491]), .Q(\_zzLB[2][523] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][524] ( .G(n180), .D(idata[492]), .Q(\_zzLB[2][524] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][525] ( .G(n180), .D(idata[493]), .Q(\_zzLB[2][525] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][526] ( .G(n180), .D(idata[494]), .Q(\_zzLB[2][526] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][527] ( .G(n180), .D(idata[495]), .Q(\_zzLB[2][527] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][528] ( .G(n180), .D(idata[496]), .Q(\_zzLB[2][528] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][529] ( .G(n180), .D(idata[497]), .Q(\_zzLB[2][529] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][530] ( .G(n180), .D(idata[498]), .Q(\_zzLB[2][530] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][531] ( .G(n180), .D(idata[499]), .Q(\_zzLB[2][531] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][532] ( .G(n180), .D(idata[500]), .Q(\_zzLB[2][532] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][533] ( .G(n180), .D(idata[501]), .Q(\_zzLB[2][533] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][534] ( .G(n180), .D(idata[502]), .Q(\_zzLB[2][534] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][535] ( .G(n180), .D(idata[503]), .Q(\_zzLB[2][535] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][536] ( .G(n180), .D(idata[504]), .Q(\_zzLB[2][536] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][537] ( .G(n180), .D(idata[505]), .Q(\_zzLB[2][537] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][538] ( .G(n180), .D(idata[506]), .Q(\_zzLB[2][538] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][539] ( .G(n180), .D(idata[507]), .Q(\_zzLB[2][539] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][540] ( .G(n180), .D(idata[508]), .Q(\_zzLB[2][540] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][541] ( .G(n180), .D(idata[509]), .Q(\_zzLB[2][541] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][542] ( .G(n180), .D(idata[510]), .Q(\_zzLB[2][542] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][543] ( .G(n180), .D(idata[511]), .Q(\_zzLB[2][543] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][544] ( .G(n180), .D(idata[512]), .Q(\_zzLB[2][544] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][545] ( .G(n180), .D(idata[513]), .Q(\_zzLB[2][545] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][546] ( .G(n180), .D(idata[514]), .Q(\_zzLB[2][546] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][547] ( .G(n180), .D(idata[515]), .Q(\_zzLB[2][547] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][548] ( .G(n180), .D(idata[516]), .Q(\_zzLB[2][548] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][549] ( .G(n180), .D(idata[517]), .Q(\_zzLB[2][549] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][550] ( .G(n180), .D(idata[518]), .Q(\_zzLB[2][550] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][551] ( .G(n180), .D(idata[519]), .Q(\_zzLB[2][551] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][552] ( .G(n180), .D(idata[520]), .Q(\_zzLB[2][552] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][553] ( .G(n180), .D(idata[521]), .Q(\_zzLB[2][553] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][554] ( .G(n180), .D(idata[522]), .Q(\_zzLB[2][554] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][555] ( .G(n180), .D(idata[523]), .Q(\_zzLB[2][555] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][556] ( .G(n180), .D(idata[524]), .Q(\_zzLB[2][556] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][557] ( .G(n180), .D(idata[525]), .Q(\_zzLB[2][557] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][558] ( .G(n180), .D(idata[526]), .Q(\_zzLB[2][558] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][559] ( .G(n180), .D(idata[527]), .Q(\_zzLB[2][559] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][560] ( .G(n180), .D(idata[528]), .Q(\_zzLB[2][560] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][561] ( .G(n180), .D(idata[529]), .Q(\_zzLB[2][561] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][562] ( .G(n180), .D(idata[530]), .Q(\_zzLB[2][562] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][563] ( .G(n180), .D(idata[531]), .Q(\_zzLB[2][563] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][564] ( .G(n180), .D(idata[532]), .Q(\_zzLB[2][564] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][565] ( .G(n180), .D(idata[533]), .Q(\_zzLB[2][565] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][566] ( .G(n180), .D(idata[534]), .Q(\_zzLB[2][566] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][567] ( .G(n180), .D(idata[535]), .Q(\_zzLB[2][567] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][568] ( .G(n180), .D(idata[536]), .Q(\_zzLB[2][568] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][569] ( .G(n180), .D(idata[537]), .Q(\_zzLB[2][569] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][570] ( .G(n180), .D(idata[538]), .Q(\_zzLB[2][570] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][571] ( .G(n180), .D(idata[539]), .Q(\_zzLB[2][571] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][572] ( .G(n180), .D(idata[540]), .Q(\_zzLB[2][572] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][573] ( .G(n180), .D(idata[541]), .Q(\_zzLB[2][573] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][574] ( .G(n180), .D(idata[542]), .Q(\_zzLB[2][574] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][575] ( .G(n180), .D(idata[543]), .Q(\_zzLB[2][575] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][576] ( .G(n180), .D(idata[544]), .Q(\_zzLB[2][576] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][577] ( .G(n180), .D(idata[545]), .Q(\_zzLB[2][577] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][578] ( .G(n180), .D(idata[546]), .Q(\_zzLB[2][578] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][579] ( .G(n180), .D(idata[547]), .Q(\_zzLB[2][579] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][580] ( .G(n180), .D(idata[548]), .Q(\_zzLB[2][580] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][581] ( .G(n180), .D(idata[549]), .Q(\_zzLB[2][581] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][582] ( .G(n180), .D(idata[550]), .Q(\_zzLB[2][582] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][583] ( .G(n180), .D(idata[551]), .Q(\_zzLB[2][583] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][584] ( .G(n180), .D(idata[552]), .Q(\_zzLB[2][584] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][585] ( .G(n180), .D(idata[553]), .Q(\_zzLB[2][585] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][586] ( .G(n180), .D(idata[554]), .Q(\_zzLB[2][586] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][587] ( .G(n180), .D(idata[555]), .Q(\_zzLB[2][587] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][588] ( .G(n180), .D(idata[556]), .Q(\_zzLB[2][588] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][589] ( .G(n180), .D(idata[557]), .Q(\_zzLB[2][589] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][590] ( .G(n180), .D(idata[558]), .Q(\_zzLB[2][590] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][591] ( .G(n180), .D(idata[559]), .Q(\_zzLB[2][591] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][592] ( .G(n180), .D(ireq), .Q(\_zzLB[2][592] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][0] ( .G(n181), .D(len[0]), .Q(\_zzLB[3][0] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][1] ( .G(n181), .D(len[1]), .Q(\_zzLB[3][1] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][2] ( .G(n181), .D(len[2]), .Q(\_zzLB[3][2] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][3] ( .G(n181), .D(len[3]), .Q(\_zzLB[3][3] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][4] ( .G(n181), .D(len[4]), .Q(\_zzLB[3][4] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][5] ( .G(n181), .D(len[5]), .Q(\_zzLB[3][5] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][6] ( .G(n181), .D(len[6]), .Q(\_zzLB[3][6] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][7] ( .G(n181), .D(len[7]), .Q(\_zzLB[3][7] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][8] ( .G(n181), .D(len[8]), .Q(\_zzLB[3][8] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][9] ( .G(n181), .D(len[9]), .Q(\_zzLB[3][9] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][10] ( .G(n181), .D(len[10]), .Q(\_zzLB[3][10] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][11] ( .G(n181), .D(len[11]), .Q(\_zzLB[3][11] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][12] ( .G(n181), .D(cbid[0]), .Q(\_zzLB[3][12] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][13] ( .G(n181), .D(cbid[1]), .Q(\_zzLB[3][13] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][14] ( .G(n181), .D(cbid[2]), .Q(\_zzLB[3][14] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][15] ( .G(n181), .D(cbid[3]), .Q(\_zzLB[3][15] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][16] ( .G(n181), .D(cbid[4]), .Q(\_zzLB[3][16] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][17] ( .G(n181), .D(cbid[5]), .Q(\_zzLB[3][17] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][18] ( .G(n181), .D(cbid[6]), .Q(\_zzLB[3][18] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][19] ( .G(n181), .D(cbid[7]), .Q(\_zzLB[3][19] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][20] ( .G(n181), .D(cbid[8]), .Q(\_zzLB[3][20] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][21] ( .G(n181), .D(cbid[9]), .Q(\_zzLB[3][21] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][22] ( .G(n181), .D(cbid[10]), .Q(\_zzLB[3][22] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][23] ( .G(n181), .D(cbid[11]), .Q(\_zzLB[3][23] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][24] ( .G(n181), .D(cbid[12]), .Q(\_zzLB[3][24] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][25] ( .G(n181), .D(cbid[13]), .Q(\_zzLB[3][25] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][26] ( .G(n181), .D(cbid[14]), .Q(\_zzLB[3][26] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][27] ( .G(n181), .D(cbid[15]), .Q(\_zzLB[3][27] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][28] ( .G(n181), .D(cbid[16]), .Q(\_zzLB[3][28] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][29] ( .G(n181), .D(cbid[17]), .Q(\_zzLB[3][29] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][30] ( .G(n181), .D(cbid[18]), .Q(\_zzLB[3][30] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][31] ( .G(n181), .D(cbid[19]), .Q(\_zzLB[3][31] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][32] ( .G(n181), .D(idata[0]), .Q(\_zzLB[3][32] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][33] ( .G(n181), .D(idata[1]), .Q(\_zzLB[3][33] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][34] ( .G(n181), .D(idata[2]), .Q(\_zzLB[3][34] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][35] ( .G(n181), .D(idata[3]), .Q(\_zzLB[3][35] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][36] ( .G(n181), .D(idata[4]), .Q(\_zzLB[3][36] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][37] ( .G(n181), .D(idata[5]), .Q(\_zzLB[3][37] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][38] ( .G(n181), .D(idata[6]), .Q(\_zzLB[3][38] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][39] ( .G(n181), .D(idata[7]), .Q(\_zzLB[3][39] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][40] ( .G(n181), .D(idata[8]), .Q(\_zzLB[3][40] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][41] ( .G(n181), .D(idata[9]), .Q(\_zzLB[3][41] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][42] ( .G(n181), .D(idata[10]), .Q(\_zzLB[3][42] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][43] ( .G(n181), .D(idata[11]), .Q(\_zzLB[3][43] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][44] ( .G(n181), .D(idata[12]), .Q(\_zzLB[3][44] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][45] ( .G(n181), .D(idata[13]), .Q(\_zzLB[3][45] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][46] ( .G(n181), .D(idata[14]), .Q(\_zzLB[3][46] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][47] ( .G(n181), .D(idata[15]), .Q(\_zzLB[3][47] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][48] ( .G(n181), .D(idata[16]), .Q(\_zzLB[3][48] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][49] ( .G(n181), .D(idata[17]), .Q(\_zzLB[3][49] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][50] ( .G(n181), .D(idata[18]), .Q(\_zzLB[3][50] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][51] ( .G(n181), .D(idata[19]), .Q(\_zzLB[3][51] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][52] ( .G(n181), .D(idata[20]), .Q(\_zzLB[3][52] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][53] ( .G(n181), .D(idata[21]), .Q(\_zzLB[3][53] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][54] ( .G(n181), .D(idata[22]), .Q(\_zzLB[3][54] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][55] ( .G(n181), .D(idata[23]), .Q(\_zzLB[3][55] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][56] ( .G(n181), .D(idata[24]), .Q(\_zzLB[3][56] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][57] ( .G(n181), .D(idata[25]), .Q(\_zzLB[3][57] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][58] ( .G(n181), .D(idata[26]), .Q(\_zzLB[3][58] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][59] ( .G(n181), .D(idata[27]), .Q(\_zzLB[3][59] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][60] ( .G(n181), .D(idata[28]), .Q(\_zzLB[3][60] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][61] ( .G(n181), .D(idata[29]), .Q(\_zzLB[3][61] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][62] ( .G(n181), .D(idata[30]), .Q(\_zzLB[3][62] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][63] ( .G(n181), .D(idata[31]), .Q(\_zzLB[3][63] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][64] ( .G(n181), .D(idata[32]), .Q(\_zzLB[3][64] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][65] ( .G(n181), .D(idata[33]), .Q(\_zzLB[3][65] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][66] ( .G(n181), .D(idata[34]), .Q(\_zzLB[3][66] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][67] ( .G(n181), .D(idata[35]), .Q(\_zzLB[3][67] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][68] ( .G(n181), .D(idata[36]), .Q(\_zzLB[3][68] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][69] ( .G(n181), .D(idata[37]), .Q(\_zzLB[3][69] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][70] ( .G(n181), .D(idata[38]), .Q(\_zzLB[3][70] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][71] ( .G(n181), .D(idata[39]), .Q(\_zzLB[3][71] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][72] ( .G(n181), .D(idata[40]), .Q(\_zzLB[3][72] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][73] ( .G(n181), .D(idata[41]), .Q(\_zzLB[3][73] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][74] ( .G(n181), .D(idata[42]), .Q(\_zzLB[3][74] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][75] ( .G(n181), .D(idata[43]), .Q(\_zzLB[3][75] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][76] ( .G(n181), .D(idata[44]), .Q(\_zzLB[3][76] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][77] ( .G(n181), .D(idata[45]), .Q(\_zzLB[3][77] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][78] ( .G(n181), .D(idata[46]), .Q(\_zzLB[3][78] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][79] ( .G(n181), .D(idata[47]), .Q(\_zzLB[3][79] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][80] ( .G(n181), .D(idata[48]), .Q(\_zzLB[3][80] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][81] ( .G(n181), .D(idata[49]), .Q(\_zzLB[3][81] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][82] ( .G(n181), .D(idata[50]), .Q(\_zzLB[3][82] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][83] ( .G(n181), .D(idata[51]), .Q(\_zzLB[3][83] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][84] ( .G(n181), .D(idata[52]), .Q(\_zzLB[3][84] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][85] ( .G(n181), .D(idata[53]), .Q(\_zzLB[3][85] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][86] ( .G(n181), .D(idata[54]), .Q(\_zzLB[3][86] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][87] ( .G(n181), .D(idata[55]), .Q(\_zzLB[3][87] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][88] ( .G(n181), .D(idata[56]), .Q(\_zzLB[3][88] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][89] ( .G(n181), .D(idata[57]), .Q(\_zzLB[3][89] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][90] ( .G(n181), .D(idata[58]), .Q(\_zzLB[3][90] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][91] ( .G(n181), .D(idata[59]), .Q(\_zzLB[3][91] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][92] ( .G(n181), .D(idata[60]), .Q(\_zzLB[3][92] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][93] ( .G(n181), .D(idata[61]), .Q(\_zzLB[3][93] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][94] ( .G(n181), .D(idata[62]), .Q(\_zzLB[3][94] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][95] ( .G(n181), .D(idata[63]), .Q(\_zzLB[3][95] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][96] ( .G(n181), .D(idata[64]), .Q(\_zzLB[3][96] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][97] ( .G(n181), .D(idata[65]), .Q(\_zzLB[3][97] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][98] ( .G(n181), .D(idata[66]), .Q(\_zzLB[3][98] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][99] ( .G(n181), .D(idata[67]), .Q(\_zzLB[3][99] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][100] ( .G(n181), .D(idata[68]), .Q(\_zzLB[3][100] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][101] ( .G(n181), .D(idata[69]), .Q(\_zzLB[3][101] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][102] ( .G(n181), .D(idata[70]), .Q(\_zzLB[3][102] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][103] ( .G(n181), .D(idata[71]), .Q(\_zzLB[3][103] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][104] ( .G(n181), .D(idata[72]), .Q(\_zzLB[3][104] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][105] ( .G(n181), .D(idata[73]), .Q(\_zzLB[3][105] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][106] ( .G(n181), .D(idata[74]), .Q(\_zzLB[3][106] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][107] ( .G(n181), .D(idata[75]), .Q(\_zzLB[3][107] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][108] ( .G(n181), .D(idata[76]), .Q(\_zzLB[3][108] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][109] ( .G(n181), .D(idata[77]), .Q(\_zzLB[3][109] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][110] ( .G(n181), .D(idata[78]), .Q(\_zzLB[3][110] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][111] ( .G(n181), .D(idata[79]), .Q(\_zzLB[3][111] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][112] ( .G(n181), .D(idata[80]), .Q(\_zzLB[3][112] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][113] ( .G(n181), .D(idata[81]), .Q(\_zzLB[3][113] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][114] ( .G(n181), .D(idata[82]), .Q(\_zzLB[3][114] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][115] ( .G(n181), .D(idata[83]), .Q(\_zzLB[3][115] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][116] ( .G(n181), .D(idata[84]), .Q(\_zzLB[3][116] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][117] ( .G(n181), .D(idata[85]), .Q(\_zzLB[3][117] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][118] ( .G(n181), .D(idata[86]), .Q(\_zzLB[3][118] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][119] ( .G(n181), .D(idata[87]), .Q(\_zzLB[3][119] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][120] ( .G(n181), .D(idata[88]), .Q(\_zzLB[3][120] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][121] ( .G(n181), .D(idata[89]), .Q(\_zzLB[3][121] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][122] ( .G(n181), .D(idata[90]), .Q(\_zzLB[3][122] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][123] ( .G(n181), .D(idata[91]), .Q(\_zzLB[3][123] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][124] ( .G(n181), .D(idata[92]), .Q(\_zzLB[3][124] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][125] ( .G(n181), .D(idata[93]), .Q(\_zzLB[3][125] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][126] ( .G(n181), .D(idata[94]), .Q(\_zzLB[3][126] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][127] ( .G(n181), .D(idata[95]), .Q(\_zzLB[3][127] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][128] ( .G(n181), .D(idata[96]), .Q(\_zzLB[3][128] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][129] ( .G(n181), .D(idata[97]), .Q(\_zzLB[3][129] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][130] ( .G(n181), .D(idata[98]), .Q(\_zzLB[3][130] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][131] ( .G(n181), .D(idata[99]), .Q(\_zzLB[3][131] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][132] ( .G(n181), .D(idata[100]), .Q(\_zzLB[3][132] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][133] ( .G(n181), .D(idata[101]), .Q(\_zzLB[3][133] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][134] ( .G(n181), .D(idata[102]), .Q(\_zzLB[3][134] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][135] ( .G(n181), .D(idata[103]), .Q(\_zzLB[3][135] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][136] ( .G(n181), .D(idata[104]), .Q(\_zzLB[3][136] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][137] ( .G(n181), .D(idata[105]), .Q(\_zzLB[3][137] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][138] ( .G(n181), .D(idata[106]), .Q(\_zzLB[3][138] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][139] ( .G(n181), .D(idata[107]), .Q(\_zzLB[3][139] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][140] ( .G(n181), .D(idata[108]), .Q(\_zzLB[3][140] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][141] ( .G(n181), .D(idata[109]), .Q(\_zzLB[3][141] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][142] ( .G(n181), .D(idata[110]), .Q(\_zzLB[3][142] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][143] ( .G(n181), .D(idata[111]), .Q(\_zzLB[3][143] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][144] ( .G(n181), .D(idata[112]), .Q(\_zzLB[3][144] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][145] ( .G(n181), .D(idata[113]), .Q(\_zzLB[3][145] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][146] ( .G(n181), .D(idata[114]), .Q(\_zzLB[3][146] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][147] ( .G(n181), .D(idata[115]), .Q(\_zzLB[3][147] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][148] ( .G(n181), .D(idata[116]), .Q(\_zzLB[3][148] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][149] ( .G(n181), .D(idata[117]), .Q(\_zzLB[3][149] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][150] ( .G(n181), .D(idata[118]), .Q(\_zzLB[3][150] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][151] ( .G(n181), .D(idata[119]), .Q(\_zzLB[3][151] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][152] ( .G(n181), .D(idata[120]), .Q(\_zzLB[3][152] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][153] ( .G(n181), .D(idata[121]), .Q(\_zzLB[3][153] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][154] ( .G(n181), .D(idata[122]), .Q(\_zzLB[3][154] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][155] ( .G(n181), .D(idata[123]), .Q(\_zzLB[3][155] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][156] ( .G(n181), .D(idata[124]), .Q(\_zzLB[3][156] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][157] ( .G(n181), .D(idata[125]), .Q(\_zzLB[3][157] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][158] ( .G(n181), .D(idata[126]), .Q(\_zzLB[3][158] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][159] ( .G(n181), .D(idata[127]), .Q(\_zzLB[3][159] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][160] ( .G(n181), .D(idata[128]), .Q(\_zzLB[3][160] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][161] ( .G(n181), .D(idata[129]), .Q(\_zzLB[3][161] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][162] ( .G(n181), .D(idata[130]), .Q(\_zzLB[3][162] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][163] ( .G(n181), .D(idata[131]), .Q(\_zzLB[3][163] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][164] ( .G(n181), .D(idata[132]), .Q(\_zzLB[3][164] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][165] ( .G(n181), .D(idata[133]), .Q(\_zzLB[3][165] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][166] ( .G(n181), .D(idata[134]), .Q(\_zzLB[3][166] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][167] ( .G(n181), .D(idata[135]), .Q(\_zzLB[3][167] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][168] ( .G(n181), .D(idata[136]), .Q(\_zzLB[3][168] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][169] ( .G(n181), .D(idata[137]), .Q(\_zzLB[3][169] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][170] ( .G(n181), .D(idata[138]), .Q(\_zzLB[3][170] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][171] ( .G(n181), .D(idata[139]), .Q(\_zzLB[3][171] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][172] ( .G(n181), .D(idata[140]), .Q(\_zzLB[3][172] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][173] ( .G(n181), .D(idata[141]), .Q(\_zzLB[3][173] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][174] ( .G(n181), .D(idata[142]), .Q(\_zzLB[3][174] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][175] ( .G(n181), .D(idata[143]), .Q(\_zzLB[3][175] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][176] ( .G(n181), .D(idata[144]), .Q(\_zzLB[3][176] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][177] ( .G(n181), .D(idata[145]), .Q(\_zzLB[3][177] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][178] ( .G(n181), .D(idata[146]), .Q(\_zzLB[3][178] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][179] ( .G(n181), .D(idata[147]), .Q(\_zzLB[3][179] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][180] ( .G(n181), .D(idata[148]), .Q(\_zzLB[3][180] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][181] ( .G(n181), .D(idata[149]), .Q(\_zzLB[3][181] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][182] ( .G(n181), .D(idata[150]), .Q(\_zzLB[3][182] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][183] ( .G(n181), .D(idata[151]), .Q(\_zzLB[3][183] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][184] ( .G(n181), .D(idata[152]), .Q(\_zzLB[3][184] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][185] ( .G(n181), .D(idata[153]), .Q(\_zzLB[3][185] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][186] ( .G(n181), .D(idata[154]), .Q(\_zzLB[3][186] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][187] ( .G(n181), .D(idata[155]), .Q(\_zzLB[3][187] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][188] ( .G(n181), .D(idata[156]), .Q(\_zzLB[3][188] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][189] ( .G(n181), .D(idata[157]), .Q(\_zzLB[3][189] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][190] ( .G(n181), .D(idata[158]), .Q(\_zzLB[3][190] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][191] ( .G(n181), .D(idata[159]), .Q(\_zzLB[3][191] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][192] ( .G(n181), .D(idata[160]), .Q(\_zzLB[3][192] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][193] ( .G(n181), .D(idata[161]), .Q(\_zzLB[3][193] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][194] ( .G(n181), .D(idata[162]), .Q(\_zzLB[3][194] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][195] ( .G(n181), .D(idata[163]), .Q(\_zzLB[3][195] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][196] ( .G(n181), .D(idata[164]), .Q(\_zzLB[3][196] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][197] ( .G(n181), .D(idata[165]), .Q(\_zzLB[3][197] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][198] ( .G(n181), .D(idata[166]), .Q(\_zzLB[3][198] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][199] ( .G(n181), .D(idata[167]), .Q(\_zzLB[3][199] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][200] ( .G(n181), .D(idata[168]), .Q(\_zzLB[3][200] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][201] ( .G(n181), .D(idata[169]), .Q(\_zzLB[3][201] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][202] ( .G(n181), .D(idata[170]), .Q(\_zzLB[3][202] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][203] ( .G(n181), .D(idata[171]), .Q(\_zzLB[3][203] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][204] ( .G(n181), .D(idata[172]), .Q(\_zzLB[3][204] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][205] ( .G(n181), .D(idata[173]), .Q(\_zzLB[3][205] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][206] ( .G(n181), .D(idata[174]), .Q(\_zzLB[3][206] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][207] ( .G(n181), .D(idata[175]), .Q(\_zzLB[3][207] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][208] ( .G(n181), .D(idata[176]), .Q(\_zzLB[3][208] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][209] ( .G(n181), .D(idata[177]), .Q(\_zzLB[3][209] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][210] ( .G(n181), .D(idata[178]), .Q(\_zzLB[3][210] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][211] ( .G(n181), .D(idata[179]), .Q(\_zzLB[3][211] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][212] ( .G(n181), .D(idata[180]), .Q(\_zzLB[3][212] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][213] ( .G(n181), .D(idata[181]), .Q(\_zzLB[3][213] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][214] ( .G(n181), .D(idata[182]), .Q(\_zzLB[3][214] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][215] ( .G(n181), .D(idata[183]), .Q(\_zzLB[3][215] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][216] ( .G(n181), .D(idata[184]), .Q(\_zzLB[3][216] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][217] ( .G(n181), .D(idata[185]), .Q(\_zzLB[3][217] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][218] ( .G(n181), .D(idata[186]), .Q(\_zzLB[3][218] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][219] ( .G(n181), .D(idata[187]), .Q(\_zzLB[3][219] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][220] ( .G(n181), .D(idata[188]), .Q(\_zzLB[3][220] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][221] ( .G(n181), .D(idata[189]), .Q(\_zzLB[3][221] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][222] ( .G(n181), .D(idata[190]), .Q(\_zzLB[3][222] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][223] ( .G(n181), .D(idata[191]), .Q(\_zzLB[3][223] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][224] ( .G(n181), .D(idata[192]), .Q(\_zzLB[3][224] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][225] ( .G(n181), .D(idata[193]), .Q(\_zzLB[3][225] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][226] ( .G(n181), .D(idata[194]), .Q(\_zzLB[3][226] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][227] ( .G(n181), .D(idata[195]), .Q(\_zzLB[3][227] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][228] ( .G(n181), .D(idata[196]), .Q(\_zzLB[3][228] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][229] ( .G(n181), .D(idata[197]), .Q(\_zzLB[3][229] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][230] ( .G(n181), .D(idata[198]), .Q(\_zzLB[3][230] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][231] ( .G(n181), .D(idata[199]), .Q(\_zzLB[3][231] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][232] ( .G(n181), .D(idata[200]), .Q(\_zzLB[3][232] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][233] ( .G(n181), .D(idata[201]), .Q(\_zzLB[3][233] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][234] ( .G(n181), .D(idata[202]), .Q(\_zzLB[3][234] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][235] ( .G(n181), .D(idata[203]), .Q(\_zzLB[3][235] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][236] ( .G(n181), .D(idata[204]), .Q(\_zzLB[3][236] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][237] ( .G(n181), .D(idata[205]), .Q(\_zzLB[3][237] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][238] ( .G(n181), .D(idata[206]), .Q(\_zzLB[3][238] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][239] ( .G(n181), .D(idata[207]), .Q(\_zzLB[3][239] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][240] ( .G(n181), .D(idata[208]), .Q(\_zzLB[3][240] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][241] ( .G(n181), .D(idata[209]), .Q(\_zzLB[3][241] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][242] ( .G(n181), .D(idata[210]), .Q(\_zzLB[3][242] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][243] ( .G(n181), .D(idata[211]), .Q(\_zzLB[3][243] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][244] ( .G(n181), .D(idata[212]), .Q(\_zzLB[3][244] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][245] ( .G(n181), .D(idata[213]), .Q(\_zzLB[3][245] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][246] ( .G(n181), .D(idata[214]), .Q(\_zzLB[3][246] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][247] ( .G(n181), .D(idata[215]), .Q(\_zzLB[3][247] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][248] ( .G(n181), .D(idata[216]), .Q(\_zzLB[3][248] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][249] ( .G(n181), .D(idata[217]), .Q(\_zzLB[3][249] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][250] ( .G(n181), .D(idata[218]), .Q(\_zzLB[3][250] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][251] ( .G(n181), .D(idata[219]), .Q(\_zzLB[3][251] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][252] ( .G(n181), .D(idata[220]), .Q(\_zzLB[3][252] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][253] ( .G(n181), .D(idata[221]), .Q(\_zzLB[3][253] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][254] ( .G(n181), .D(idata[222]), .Q(\_zzLB[3][254] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][255] ( .G(n181), .D(idata[223]), .Q(\_zzLB[3][255] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][256] ( .G(n181), .D(idata[224]), .Q(\_zzLB[3][256] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][257] ( .G(n181), .D(idata[225]), .Q(\_zzLB[3][257] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][258] ( .G(n181), .D(idata[226]), .Q(\_zzLB[3][258] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][259] ( .G(n181), .D(idata[227]), .Q(\_zzLB[3][259] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][260] ( .G(n181), .D(idata[228]), .Q(\_zzLB[3][260] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][261] ( .G(n181), .D(idata[229]), .Q(\_zzLB[3][261] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][262] ( .G(n181), .D(idata[230]), .Q(\_zzLB[3][262] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][263] ( .G(n181), .D(idata[231]), .Q(\_zzLB[3][263] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][264] ( .G(n181), .D(idata[232]), .Q(\_zzLB[3][264] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][265] ( .G(n181), .D(idata[233]), .Q(\_zzLB[3][265] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][266] ( .G(n181), .D(idata[234]), .Q(\_zzLB[3][266] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][267] ( .G(n181), .D(idata[235]), .Q(\_zzLB[3][267] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][268] ( .G(n181), .D(idata[236]), .Q(\_zzLB[3][268] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][269] ( .G(n181), .D(idata[237]), .Q(\_zzLB[3][269] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][270] ( .G(n181), .D(idata[238]), .Q(\_zzLB[3][270] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][271] ( .G(n181), .D(idata[239]), .Q(\_zzLB[3][271] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][272] ( .G(n181), .D(idata[240]), .Q(\_zzLB[3][272] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][273] ( .G(n181), .D(idata[241]), .Q(\_zzLB[3][273] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][274] ( .G(n181), .D(idata[242]), .Q(\_zzLB[3][274] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][275] ( .G(n181), .D(idata[243]), .Q(\_zzLB[3][275] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][276] ( .G(n181), .D(idata[244]), .Q(\_zzLB[3][276] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][277] ( .G(n181), .D(idata[245]), .Q(\_zzLB[3][277] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][278] ( .G(n181), .D(idata[246]), .Q(\_zzLB[3][278] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][279] ( .G(n181), .D(idata[247]), .Q(\_zzLB[3][279] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][280] ( .G(n181), .D(idata[248]), .Q(\_zzLB[3][280] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][281] ( .G(n181), .D(idata[249]), .Q(\_zzLB[3][281] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][282] ( .G(n181), .D(idata[250]), .Q(\_zzLB[3][282] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][283] ( .G(n181), .D(idata[251]), .Q(\_zzLB[3][283] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][284] ( .G(n181), .D(idata[252]), .Q(\_zzLB[3][284] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][285] ( .G(n181), .D(idata[253]), .Q(\_zzLB[3][285] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][286] ( .G(n181), .D(idata[254]), .Q(\_zzLB[3][286] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][287] ( .G(n181), .D(idata[255]), .Q(\_zzLB[3][287] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][288] ( .G(n181), .D(idata[256]), .Q(\_zzLB[3][288] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][289] ( .G(n181), .D(idata[257]), .Q(\_zzLB[3][289] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][290] ( .G(n181), .D(idata[258]), .Q(\_zzLB[3][290] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][291] ( .G(n181), .D(idata[259]), .Q(\_zzLB[3][291] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][292] ( .G(n181), .D(idata[260]), .Q(\_zzLB[3][292] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][293] ( .G(n181), .D(idata[261]), .Q(\_zzLB[3][293] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][294] ( .G(n181), .D(idata[262]), .Q(\_zzLB[3][294] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][295] ( .G(n181), .D(idata[263]), .Q(\_zzLB[3][295] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][296] ( .G(n181), .D(idata[264]), .Q(\_zzLB[3][296] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][297] ( .G(n181), .D(idata[265]), .Q(\_zzLB[3][297] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][298] ( .G(n181), .D(idata[266]), .Q(\_zzLB[3][298] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][299] ( .G(n181), .D(idata[267]), .Q(\_zzLB[3][299] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][300] ( .G(n181), .D(idata[268]), .Q(\_zzLB[3][300] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][301] ( .G(n181), .D(idata[269]), .Q(\_zzLB[3][301] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][302] ( .G(n181), .D(idata[270]), .Q(\_zzLB[3][302] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][303] ( .G(n181), .D(idata[271]), .Q(\_zzLB[3][303] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][304] ( .G(n181), .D(idata[272]), .Q(\_zzLB[3][304] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][305] ( .G(n181), .D(idata[273]), .Q(\_zzLB[3][305] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][306] ( .G(n181), .D(idata[274]), .Q(\_zzLB[3][306] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][307] ( .G(n181), .D(idata[275]), .Q(\_zzLB[3][307] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][308] ( .G(n181), .D(idata[276]), .Q(\_zzLB[3][308] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][309] ( .G(n181), .D(idata[277]), .Q(\_zzLB[3][309] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][310] ( .G(n181), .D(idata[278]), .Q(\_zzLB[3][310] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][311] ( .G(n181), .D(idata[279]), .Q(\_zzLB[3][311] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][312] ( .G(n181), .D(idata[280]), .Q(\_zzLB[3][312] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][313] ( .G(n181), .D(idata[281]), .Q(\_zzLB[3][313] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][314] ( .G(n181), .D(idata[282]), .Q(\_zzLB[3][314] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][315] ( .G(n181), .D(idata[283]), .Q(\_zzLB[3][315] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][316] ( .G(n181), .D(idata[284]), .Q(\_zzLB[3][316] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][317] ( .G(n181), .D(idata[285]), .Q(\_zzLB[3][317] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][318] ( .G(n181), .D(idata[286]), .Q(\_zzLB[3][318] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][319] ( .G(n181), .D(idata[287]), .Q(\_zzLB[3][319] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][320] ( .G(n181), .D(idata[288]), .Q(\_zzLB[3][320] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][321] ( .G(n181), .D(idata[289]), .Q(\_zzLB[3][321] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][322] ( .G(n181), .D(idata[290]), .Q(\_zzLB[3][322] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][323] ( .G(n181), .D(idata[291]), .Q(\_zzLB[3][323] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][324] ( .G(n181), .D(idata[292]), .Q(\_zzLB[3][324] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][325] ( .G(n181), .D(idata[293]), .Q(\_zzLB[3][325] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][326] ( .G(n181), .D(idata[294]), .Q(\_zzLB[3][326] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][327] ( .G(n181), .D(idata[295]), .Q(\_zzLB[3][327] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][328] ( .G(n181), .D(idata[296]), .Q(\_zzLB[3][328] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][329] ( .G(n181), .D(idata[297]), .Q(\_zzLB[3][329] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][330] ( .G(n181), .D(idata[298]), .Q(\_zzLB[3][330] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][331] ( .G(n181), .D(idata[299]), .Q(\_zzLB[3][331] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][332] ( .G(n181), .D(idata[300]), .Q(\_zzLB[3][332] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][333] ( .G(n181), .D(idata[301]), .Q(\_zzLB[3][333] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][334] ( .G(n181), .D(idata[302]), .Q(\_zzLB[3][334] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][335] ( .G(n181), .D(idata[303]), .Q(\_zzLB[3][335] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][336] ( .G(n181), .D(idata[304]), .Q(\_zzLB[3][336] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][337] ( .G(n181), .D(idata[305]), .Q(\_zzLB[3][337] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][338] ( .G(n181), .D(idata[306]), .Q(\_zzLB[3][338] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][339] ( .G(n181), .D(idata[307]), .Q(\_zzLB[3][339] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][340] ( .G(n181), .D(idata[308]), .Q(\_zzLB[3][340] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][341] ( .G(n181), .D(idata[309]), .Q(\_zzLB[3][341] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][342] ( .G(n181), .D(idata[310]), .Q(\_zzLB[3][342] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][343] ( .G(n181), .D(idata[311]), .Q(\_zzLB[3][343] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][344] ( .G(n181), .D(idata[312]), .Q(\_zzLB[3][344] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][345] ( .G(n181), .D(idata[313]), .Q(\_zzLB[3][345] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][346] ( .G(n181), .D(idata[314]), .Q(\_zzLB[3][346] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][347] ( .G(n181), .D(idata[315]), .Q(\_zzLB[3][347] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][348] ( .G(n181), .D(idata[316]), .Q(\_zzLB[3][348] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][349] ( .G(n181), .D(idata[317]), .Q(\_zzLB[3][349] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][350] ( .G(n181), .D(idata[318]), .Q(\_zzLB[3][350] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][351] ( .G(n181), .D(idata[319]), .Q(\_zzLB[3][351] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][352] ( .G(n181), .D(idata[320]), .Q(\_zzLB[3][352] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][353] ( .G(n181), .D(idata[321]), .Q(\_zzLB[3][353] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][354] ( .G(n181), .D(idata[322]), .Q(\_zzLB[3][354] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][355] ( .G(n181), .D(idata[323]), .Q(\_zzLB[3][355] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][356] ( .G(n181), .D(idata[324]), .Q(\_zzLB[3][356] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][357] ( .G(n181), .D(idata[325]), .Q(\_zzLB[3][357] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][358] ( .G(n181), .D(idata[326]), .Q(\_zzLB[3][358] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][359] ( .G(n181), .D(idata[327]), .Q(\_zzLB[3][359] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][360] ( .G(n181), .D(idata[328]), .Q(\_zzLB[3][360] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][361] ( .G(n181), .D(idata[329]), .Q(\_zzLB[3][361] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][362] ( .G(n181), .D(idata[330]), .Q(\_zzLB[3][362] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][363] ( .G(n181), .D(idata[331]), .Q(\_zzLB[3][363] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][364] ( .G(n181), .D(idata[332]), .Q(\_zzLB[3][364] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][365] ( .G(n181), .D(idata[333]), .Q(\_zzLB[3][365] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][366] ( .G(n181), .D(idata[334]), .Q(\_zzLB[3][366] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][367] ( .G(n181), .D(idata[335]), .Q(\_zzLB[3][367] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][368] ( .G(n181), .D(idata[336]), .Q(\_zzLB[3][368] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][369] ( .G(n181), .D(idata[337]), .Q(\_zzLB[3][369] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][370] ( .G(n181), .D(idata[338]), .Q(\_zzLB[3][370] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][371] ( .G(n181), .D(idata[339]), .Q(\_zzLB[3][371] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][372] ( .G(n181), .D(idata[340]), .Q(\_zzLB[3][372] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][373] ( .G(n181), .D(idata[341]), .Q(\_zzLB[3][373] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][374] ( .G(n181), .D(idata[342]), .Q(\_zzLB[3][374] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][375] ( .G(n181), .D(idata[343]), .Q(\_zzLB[3][375] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][376] ( .G(n181), .D(idata[344]), .Q(\_zzLB[3][376] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][377] ( .G(n181), .D(idata[345]), .Q(\_zzLB[3][377] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][378] ( .G(n181), .D(idata[346]), .Q(\_zzLB[3][378] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][379] ( .G(n181), .D(idata[347]), .Q(\_zzLB[3][379] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][380] ( .G(n181), .D(idata[348]), .Q(\_zzLB[3][380] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][381] ( .G(n181), .D(idata[349]), .Q(\_zzLB[3][381] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][382] ( .G(n181), .D(idata[350]), .Q(\_zzLB[3][382] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][383] ( .G(n181), .D(idata[351]), .Q(\_zzLB[3][383] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][384] ( .G(n181), .D(idata[352]), .Q(\_zzLB[3][384] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][385] ( .G(n181), .D(idata[353]), .Q(\_zzLB[3][385] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][386] ( .G(n181), .D(idata[354]), .Q(\_zzLB[3][386] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][387] ( .G(n181), .D(idata[355]), .Q(\_zzLB[3][387] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][388] ( .G(n181), .D(idata[356]), .Q(\_zzLB[3][388] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][389] ( .G(n181), .D(idata[357]), .Q(\_zzLB[3][389] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][390] ( .G(n181), .D(idata[358]), .Q(\_zzLB[3][390] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][391] ( .G(n181), .D(idata[359]), .Q(\_zzLB[3][391] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][392] ( .G(n181), .D(idata[360]), .Q(\_zzLB[3][392] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][393] ( .G(n181), .D(idata[361]), .Q(\_zzLB[3][393] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][394] ( .G(n181), .D(idata[362]), .Q(\_zzLB[3][394] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][395] ( .G(n181), .D(idata[363]), .Q(\_zzLB[3][395] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][396] ( .G(n181), .D(idata[364]), .Q(\_zzLB[3][396] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][397] ( .G(n181), .D(idata[365]), .Q(\_zzLB[3][397] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][398] ( .G(n181), .D(idata[366]), .Q(\_zzLB[3][398] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][399] ( .G(n181), .D(idata[367]), .Q(\_zzLB[3][399] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][400] ( .G(n181), .D(idata[368]), .Q(\_zzLB[3][400] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][401] ( .G(n181), .D(idata[369]), .Q(\_zzLB[3][401] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][402] ( .G(n181), .D(idata[370]), .Q(\_zzLB[3][402] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][403] ( .G(n181), .D(idata[371]), .Q(\_zzLB[3][403] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][404] ( .G(n181), .D(idata[372]), .Q(\_zzLB[3][404] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][405] ( .G(n181), .D(idata[373]), .Q(\_zzLB[3][405] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][406] ( .G(n181), .D(idata[374]), .Q(\_zzLB[3][406] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][407] ( .G(n181), .D(idata[375]), .Q(\_zzLB[3][407] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][408] ( .G(n181), .D(idata[376]), .Q(\_zzLB[3][408] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][409] ( .G(n181), .D(idata[377]), .Q(\_zzLB[3][409] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][410] ( .G(n181), .D(idata[378]), .Q(\_zzLB[3][410] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][411] ( .G(n181), .D(idata[379]), .Q(\_zzLB[3][411] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][412] ( .G(n181), .D(idata[380]), .Q(\_zzLB[3][412] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][413] ( .G(n181), .D(idata[381]), .Q(\_zzLB[3][413] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][414] ( .G(n181), .D(idata[382]), .Q(\_zzLB[3][414] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][415] ( .G(n181), .D(idata[383]), .Q(\_zzLB[3][415] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][416] ( .G(n181), .D(idata[384]), .Q(\_zzLB[3][416] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][417] ( .G(n181), .D(idata[385]), .Q(\_zzLB[3][417] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][418] ( .G(n181), .D(idata[386]), .Q(\_zzLB[3][418] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][419] ( .G(n181), .D(idata[387]), .Q(\_zzLB[3][419] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][420] ( .G(n181), .D(idata[388]), .Q(\_zzLB[3][420] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][421] ( .G(n181), .D(idata[389]), .Q(\_zzLB[3][421] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][422] ( .G(n181), .D(idata[390]), .Q(\_zzLB[3][422] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][423] ( .G(n181), .D(idata[391]), .Q(\_zzLB[3][423] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][424] ( .G(n181), .D(idata[392]), .Q(\_zzLB[3][424] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][425] ( .G(n181), .D(idata[393]), .Q(\_zzLB[3][425] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][426] ( .G(n181), .D(idata[394]), .Q(\_zzLB[3][426] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][427] ( .G(n181), .D(idata[395]), .Q(\_zzLB[3][427] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][428] ( .G(n181), .D(idata[396]), .Q(\_zzLB[3][428] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][429] ( .G(n181), .D(idata[397]), .Q(\_zzLB[3][429] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][430] ( .G(n181), .D(idata[398]), .Q(\_zzLB[3][430] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][431] ( .G(n181), .D(idata[399]), .Q(\_zzLB[3][431] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][432] ( .G(n181), .D(idata[400]), .Q(\_zzLB[3][432] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][433] ( .G(n181), .D(idata[401]), .Q(\_zzLB[3][433] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][434] ( .G(n181), .D(idata[402]), .Q(\_zzLB[3][434] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][435] ( .G(n181), .D(idata[403]), .Q(\_zzLB[3][435] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][436] ( .G(n181), .D(idata[404]), .Q(\_zzLB[3][436] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][437] ( .G(n181), .D(idata[405]), .Q(\_zzLB[3][437] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][438] ( .G(n181), .D(idata[406]), .Q(\_zzLB[3][438] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][439] ( .G(n181), .D(idata[407]), .Q(\_zzLB[3][439] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][440] ( .G(n181), .D(idata[408]), .Q(\_zzLB[3][440] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][441] ( .G(n181), .D(idata[409]), .Q(\_zzLB[3][441] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][442] ( .G(n181), .D(idata[410]), .Q(\_zzLB[3][442] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][443] ( .G(n181), .D(idata[411]), .Q(\_zzLB[3][443] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][444] ( .G(n181), .D(idata[412]), .Q(\_zzLB[3][444] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][445] ( .G(n181), .D(idata[413]), .Q(\_zzLB[3][445] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][446] ( .G(n181), .D(idata[414]), .Q(\_zzLB[3][446] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][447] ( .G(n181), .D(idata[415]), .Q(\_zzLB[3][447] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][448] ( .G(n181), .D(idata[416]), .Q(\_zzLB[3][448] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][449] ( .G(n181), .D(idata[417]), .Q(\_zzLB[3][449] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][450] ( .G(n181), .D(idata[418]), .Q(\_zzLB[3][450] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][451] ( .G(n181), .D(idata[419]), .Q(\_zzLB[3][451] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][452] ( .G(n181), .D(idata[420]), .Q(\_zzLB[3][452] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][453] ( .G(n181), .D(idata[421]), .Q(\_zzLB[3][453] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][454] ( .G(n181), .D(idata[422]), .Q(\_zzLB[3][454] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][455] ( .G(n181), .D(idata[423]), .Q(\_zzLB[3][455] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][456] ( .G(n181), .D(idata[424]), .Q(\_zzLB[3][456] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][457] ( .G(n181), .D(idata[425]), .Q(\_zzLB[3][457] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][458] ( .G(n181), .D(idata[426]), .Q(\_zzLB[3][458] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][459] ( .G(n181), .D(idata[427]), .Q(\_zzLB[3][459] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][460] ( .G(n181), .D(idata[428]), .Q(\_zzLB[3][460] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][461] ( .G(n181), .D(idata[429]), .Q(\_zzLB[3][461] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][462] ( .G(n181), .D(idata[430]), .Q(\_zzLB[3][462] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][463] ( .G(n181), .D(idata[431]), .Q(\_zzLB[3][463] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][464] ( .G(n181), .D(idata[432]), .Q(\_zzLB[3][464] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][465] ( .G(n181), .D(idata[433]), .Q(\_zzLB[3][465] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][466] ( .G(n181), .D(idata[434]), .Q(\_zzLB[3][466] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][467] ( .G(n181), .D(idata[435]), .Q(\_zzLB[3][467] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][468] ( .G(n181), .D(idata[436]), .Q(\_zzLB[3][468] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][469] ( .G(n181), .D(idata[437]), .Q(\_zzLB[3][469] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][470] ( .G(n181), .D(idata[438]), .Q(\_zzLB[3][470] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][471] ( .G(n181), .D(idata[439]), .Q(\_zzLB[3][471] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][472] ( .G(n181), .D(idata[440]), .Q(\_zzLB[3][472] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][473] ( .G(n181), .D(idata[441]), .Q(\_zzLB[3][473] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][474] ( .G(n181), .D(idata[442]), .Q(\_zzLB[3][474] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][475] ( .G(n181), .D(idata[443]), .Q(\_zzLB[3][475] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][476] ( .G(n181), .D(idata[444]), .Q(\_zzLB[3][476] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][477] ( .G(n181), .D(idata[445]), .Q(\_zzLB[3][477] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][478] ( .G(n181), .D(idata[446]), .Q(\_zzLB[3][478] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][479] ( .G(n181), .D(idata[447]), .Q(\_zzLB[3][479] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][480] ( .G(n181), .D(idata[448]), .Q(\_zzLB[3][480] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][481] ( .G(n181), .D(idata[449]), .Q(\_zzLB[3][481] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][482] ( .G(n181), .D(idata[450]), .Q(\_zzLB[3][482] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][483] ( .G(n181), .D(idata[451]), .Q(\_zzLB[3][483] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][484] ( .G(n181), .D(idata[452]), .Q(\_zzLB[3][484] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][485] ( .G(n181), .D(idata[453]), .Q(\_zzLB[3][485] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][486] ( .G(n181), .D(idata[454]), .Q(\_zzLB[3][486] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][487] ( .G(n181), .D(idata[455]), .Q(\_zzLB[3][487] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][488] ( .G(n181), .D(idata[456]), .Q(\_zzLB[3][488] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][489] ( .G(n181), .D(idata[457]), .Q(\_zzLB[3][489] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][490] ( .G(n181), .D(idata[458]), .Q(\_zzLB[3][490] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][491] ( .G(n181), .D(idata[459]), .Q(\_zzLB[3][491] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][492] ( .G(n181), .D(idata[460]), .Q(\_zzLB[3][492] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][493] ( .G(n181), .D(idata[461]), .Q(\_zzLB[3][493] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][494] ( .G(n181), .D(idata[462]), .Q(\_zzLB[3][494] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][495] ( .G(n181), .D(idata[463]), .Q(\_zzLB[3][495] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][496] ( .G(n181), .D(idata[464]), .Q(\_zzLB[3][496] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][497] ( .G(n181), .D(idata[465]), .Q(\_zzLB[3][497] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][498] ( .G(n181), .D(idata[466]), .Q(\_zzLB[3][498] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][499] ( .G(n181), .D(idata[467]), .Q(\_zzLB[3][499] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][500] ( .G(n181), .D(idata[468]), .Q(\_zzLB[3][500] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][501] ( .G(n181), .D(idata[469]), .Q(\_zzLB[3][501] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][502] ( .G(n181), .D(idata[470]), .Q(\_zzLB[3][502] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][503] ( .G(n181), .D(idata[471]), .Q(\_zzLB[3][503] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][504] ( .G(n181), .D(idata[472]), .Q(\_zzLB[3][504] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][505] ( .G(n181), .D(idata[473]), .Q(\_zzLB[3][505] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][506] ( .G(n181), .D(idata[474]), .Q(\_zzLB[3][506] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][507] ( .G(n181), .D(idata[475]), .Q(\_zzLB[3][507] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][508] ( .G(n181), .D(idata[476]), .Q(\_zzLB[3][508] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][509] ( .G(n181), .D(idata[477]), .Q(\_zzLB[3][509] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][510] ( .G(n181), .D(idata[478]), .Q(\_zzLB[3][510] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][511] ( .G(n181), .D(idata[479]), .Q(\_zzLB[3][511] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][512] ( .G(n181), .D(idata[480]), .Q(\_zzLB[3][512] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][513] ( .G(n181), .D(idata[481]), .Q(\_zzLB[3][513] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][514] ( .G(n181), .D(idata[482]), .Q(\_zzLB[3][514] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][515] ( .G(n181), .D(idata[483]), .Q(\_zzLB[3][515] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][516] ( .G(n181), .D(idata[484]), .Q(\_zzLB[3][516] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][517] ( .G(n181), .D(idata[485]), .Q(\_zzLB[3][517] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][518] ( .G(n181), .D(idata[486]), .Q(\_zzLB[3][518] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][519] ( .G(n181), .D(idata[487]), .Q(\_zzLB[3][519] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][520] ( .G(n181), .D(idata[488]), .Q(\_zzLB[3][520] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][521] ( .G(n181), .D(idata[489]), .Q(\_zzLB[3][521] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][522] ( .G(n181), .D(idata[490]), .Q(\_zzLB[3][522] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][523] ( .G(n181), .D(idata[491]), .Q(\_zzLB[3][523] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][524] ( .G(n181), .D(idata[492]), .Q(\_zzLB[3][524] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][525] ( .G(n181), .D(idata[493]), .Q(\_zzLB[3][525] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][526] ( .G(n181), .D(idata[494]), .Q(\_zzLB[3][526] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][527] ( .G(n181), .D(idata[495]), .Q(\_zzLB[3][527] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][528] ( .G(n181), .D(idata[496]), .Q(\_zzLB[3][528] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][529] ( .G(n181), .D(idata[497]), .Q(\_zzLB[3][529] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][530] ( .G(n181), .D(idata[498]), .Q(\_zzLB[3][530] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][531] ( .G(n181), .D(idata[499]), .Q(\_zzLB[3][531] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][532] ( .G(n181), .D(idata[500]), .Q(\_zzLB[3][532] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][533] ( .G(n181), .D(idata[501]), .Q(\_zzLB[3][533] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][534] ( .G(n181), .D(idata[502]), .Q(\_zzLB[3][534] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][535] ( .G(n181), .D(idata[503]), .Q(\_zzLB[3][535] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][536] ( .G(n181), .D(idata[504]), .Q(\_zzLB[3][536] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][537] ( .G(n181), .D(idata[505]), .Q(\_zzLB[3][537] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][538] ( .G(n181), .D(idata[506]), .Q(\_zzLB[3][538] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][539] ( .G(n181), .D(idata[507]), .Q(\_zzLB[3][539] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][540] ( .G(n181), .D(idata[508]), .Q(\_zzLB[3][540] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][541] ( .G(n181), .D(idata[509]), .Q(\_zzLB[3][541] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][542] ( .G(n181), .D(idata[510]), .Q(\_zzLB[3][542] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][543] ( .G(n181), .D(idata[511]), .Q(\_zzLB[3][543] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][544] ( .G(n181), .D(idata[512]), .Q(\_zzLB[3][544] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][545] ( .G(n181), .D(idata[513]), .Q(\_zzLB[3][545] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][546] ( .G(n181), .D(idata[514]), .Q(\_zzLB[3][546] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][547] ( .G(n181), .D(idata[515]), .Q(\_zzLB[3][547] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][548] ( .G(n181), .D(idata[516]), .Q(\_zzLB[3][548] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][549] ( .G(n181), .D(idata[517]), .Q(\_zzLB[3][549] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][550] ( .G(n181), .D(idata[518]), .Q(\_zzLB[3][550] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][551] ( .G(n181), .D(idata[519]), .Q(\_zzLB[3][551] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][552] ( .G(n181), .D(idata[520]), .Q(\_zzLB[3][552] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][553] ( .G(n181), .D(idata[521]), .Q(\_zzLB[3][553] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][554] ( .G(n181), .D(idata[522]), .Q(\_zzLB[3][554] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][555] ( .G(n181), .D(idata[523]), .Q(\_zzLB[3][555] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][556] ( .G(n181), .D(idata[524]), .Q(\_zzLB[3][556] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][557] ( .G(n181), .D(idata[525]), .Q(\_zzLB[3][557] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][558] ( .G(n181), .D(idata[526]), .Q(\_zzLB[3][558] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][559] ( .G(n181), .D(idata[527]), .Q(\_zzLB[3][559] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][560] ( .G(n181), .D(idata[528]), .Q(\_zzLB[3][560] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][561] ( .G(n181), .D(idata[529]), .Q(\_zzLB[3][561] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][562] ( .G(n181), .D(idata[530]), .Q(\_zzLB[3][562] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][563] ( .G(n181), .D(idata[531]), .Q(\_zzLB[3][563] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][564] ( .G(n181), .D(idata[532]), .Q(\_zzLB[3][564] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][565] ( .G(n181), .D(idata[533]), .Q(\_zzLB[3][565] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][566] ( .G(n181), .D(idata[534]), .Q(\_zzLB[3][566] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][567] ( .G(n181), .D(idata[535]), .Q(\_zzLB[3][567] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][568] ( .G(n181), .D(idata[536]), .Q(\_zzLB[3][568] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][569] ( .G(n181), .D(idata[537]), .Q(\_zzLB[3][569] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][570] ( .G(n181), .D(idata[538]), .Q(\_zzLB[3][570] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][571] ( .G(n181), .D(idata[539]), .Q(\_zzLB[3][571] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][572] ( .G(n181), .D(idata[540]), .Q(\_zzLB[3][572] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][573] ( .G(n181), .D(idata[541]), .Q(\_zzLB[3][573] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][574] ( .G(n181), .D(idata[542]), .Q(\_zzLB[3][574] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][575] ( .G(n181), .D(idata[543]), .Q(\_zzLB[3][575] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][576] ( .G(n181), .D(idata[544]), .Q(\_zzLB[3][576] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][577] ( .G(n181), .D(idata[545]), .Q(\_zzLB[3][577] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][578] ( .G(n181), .D(idata[546]), .Q(\_zzLB[3][578] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][579] ( .G(n181), .D(idata[547]), .Q(\_zzLB[3][579] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][580] ( .G(n181), .D(idata[548]), .Q(\_zzLB[3][580] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][581] ( .G(n181), .D(idata[549]), .Q(\_zzLB[3][581] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][582] ( .G(n181), .D(idata[550]), .Q(\_zzLB[3][582] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][583] ( .G(n181), .D(idata[551]), .Q(\_zzLB[3][583] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][584] ( .G(n181), .D(idata[552]), .Q(\_zzLB[3][584] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][585] ( .G(n181), .D(idata[553]), .Q(\_zzLB[3][585] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][586] ( .G(n181), .D(idata[554]), .Q(\_zzLB[3][586] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][587] ( .G(n181), .D(idata[555]), .Q(\_zzLB[3][587] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][588] ( .G(n181), .D(idata[556]), .Q(\_zzLB[3][588] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][589] ( .G(n181), .D(idata[557]), .Q(\_zzLB[3][589] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][590] ( .G(n181), .D(idata[558]), .Q(\_zzLB[3][590] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][591] ( .G(n181), .D(idata[559]), .Q(\_zzLB[3][591] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][592] ( .G(n181), .D(ireq), .Q(\_zzLB[3][592] ), .QN( ));
Q_MX04 U3660 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][0] ), .A1(\_zzLB[1][0] ), .A2(\_zzLB[2][0] ), .A3(\_zzLB[3][0] ), .Z(olen[0]));
Q_MX04 U3661 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][1] ), .A1(\_zzLB[1][1] ), .A2(\_zzLB[2][1] ), .A3(\_zzLB[3][1] ), .Z(olen[1]));
Q_MX04 U3662 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][2] ), .A1(\_zzLB[1][2] ), .A2(\_zzLB[2][2] ), .A3(\_zzLB[3][2] ), .Z(olen[2]));
Q_MX04 U3663 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][3] ), .A1(\_zzLB[1][3] ), .A2(\_zzLB[2][3] ), .A3(\_zzLB[3][3] ), .Z(olen[3]));
Q_MX04 U3664 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][4] ), .A1(\_zzLB[1][4] ), .A2(\_zzLB[2][4] ), .A3(\_zzLB[3][4] ), .Z(olen[4]));
Q_MX04 U3665 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][5] ), .A1(\_zzLB[1][5] ), .A2(\_zzLB[2][5] ), .A3(\_zzLB[3][5] ), .Z(olen[5]));
Q_MX04 U3666 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][6] ), .A1(\_zzLB[1][6] ), .A2(\_zzLB[2][6] ), .A3(\_zzLB[3][6] ), .Z(olen[6]));
Q_MX04 U3667 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][7] ), .A1(\_zzLB[1][7] ), .A2(\_zzLB[2][7] ), .A3(\_zzLB[3][7] ), .Z(olen[7]));
Q_MX04 U3668 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][8] ), .A1(\_zzLB[1][8] ), .A2(\_zzLB[2][8] ), .A3(\_zzLB[3][8] ), .Z(olen[8]));
Q_MX04 U3669 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][9] ), .A1(\_zzLB[1][9] ), .A2(\_zzLB[2][9] ), .A3(\_zzLB[3][9] ), .Z(olen[9]));
Q_MX04 U3670 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][10] ), .A1(\_zzLB[1][10] ), .A2(\_zzLB[2][10] ), .A3(\_zzLB[3][10] ), .Z(olen[10]));
Q_MX04 U3671 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][11] ), .A1(\_zzLB[1][11] ), .A2(\_zzLB[2][11] ), .A3(\_zzLB[3][11] ), .Z(olen[11]));
Q_MX04 U3672 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][12] ), .A1(\_zzLB[1][12] ), .A2(\_zzLB[2][12] ), .A3(\_zzLB[3][12] ), .Z(ocbid[0]));
Q_MX04 U3673 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][13] ), .A1(\_zzLB[1][13] ), .A2(\_zzLB[2][13] ), .A3(\_zzLB[3][13] ), .Z(ocbid[1]));
Q_MX04 U3674 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][14] ), .A1(\_zzLB[1][14] ), .A2(\_zzLB[2][14] ), .A3(\_zzLB[3][14] ), .Z(ocbid[2]));
Q_MX04 U3675 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][15] ), .A1(\_zzLB[1][15] ), .A2(\_zzLB[2][15] ), .A3(\_zzLB[3][15] ), .Z(ocbid[3]));
Q_MX04 U3676 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][16] ), .A1(\_zzLB[1][16] ), .A2(\_zzLB[2][16] ), .A3(\_zzLB[3][16] ), .Z(ocbid[4]));
Q_MX04 U3677 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][17] ), .A1(\_zzLB[1][17] ), .A2(\_zzLB[2][17] ), .A3(\_zzLB[3][17] ), .Z(ocbid[5]));
Q_MX04 U3678 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][18] ), .A1(\_zzLB[1][18] ), .A2(\_zzLB[2][18] ), .A3(\_zzLB[3][18] ), .Z(ocbid[6]));
Q_MX04 U3679 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][19] ), .A1(\_zzLB[1][19] ), .A2(\_zzLB[2][19] ), .A3(\_zzLB[3][19] ), .Z(ocbid[7]));
Q_MX04 U3680 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][20] ), .A1(\_zzLB[1][20] ), .A2(\_zzLB[2][20] ), .A3(\_zzLB[3][20] ), .Z(ocbid[8]));
Q_MX04 U3681 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][21] ), .A1(\_zzLB[1][21] ), .A2(\_zzLB[2][21] ), .A3(\_zzLB[3][21] ), .Z(ocbid[9]));
Q_MX04 U3682 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][22] ), .A1(\_zzLB[1][22] ), .A2(\_zzLB[2][22] ), .A3(\_zzLB[3][22] ), .Z(ocbid[10]));
Q_MX04 U3683 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][23] ), .A1(\_zzLB[1][23] ), .A2(\_zzLB[2][23] ), .A3(\_zzLB[3][23] ), .Z(ocbid[11]));
Q_MX04 U3684 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][24] ), .A1(\_zzLB[1][24] ), .A2(\_zzLB[2][24] ), .A3(\_zzLB[3][24] ), .Z(ocbid[12]));
Q_MX04 U3685 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][25] ), .A1(\_zzLB[1][25] ), .A2(\_zzLB[2][25] ), .A3(\_zzLB[3][25] ), .Z(ocbid[13]));
Q_MX04 U3686 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][26] ), .A1(\_zzLB[1][26] ), .A2(\_zzLB[2][26] ), .A3(\_zzLB[3][26] ), .Z(ocbid[14]));
Q_MX04 U3687 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][27] ), .A1(\_zzLB[1][27] ), .A2(\_zzLB[2][27] ), .A3(\_zzLB[3][27] ), .Z(ocbid[15]));
Q_MX04 U3688 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][28] ), .A1(\_zzLB[1][28] ), .A2(\_zzLB[2][28] ), .A3(\_zzLB[3][28] ), .Z(ocbid[16]));
Q_MX04 U3689 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][29] ), .A1(\_zzLB[1][29] ), .A2(\_zzLB[2][29] ), .A3(\_zzLB[3][29] ), .Z(ocbid[17]));
Q_MX04 U3690 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][30] ), .A1(\_zzLB[1][30] ), .A2(\_zzLB[2][30] ), .A3(\_zzLB[3][30] ), .Z(ocbid[18]));
Q_MX04 U3691 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][31] ), .A1(\_zzLB[1][31] ), .A2(\_zzLB[2][31] ), .A3(\_zzLB[3][31] ), .Z(ocbid[19]));
Q_MX04 U3692 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][32] ), .A1(\_zzLB[1][32] ), .A2(\_zzLB[2][32] ), .A3(\_zzLB[3][32] ), .Z(odata[0]));
Q_MX04 U3693 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][33] ), .A1(\_zzLB[1][33] ), .A2(\_zzLB[2][33] ), .A3(\_zzLB[3][33] ), .Z(odata[1]));
Q_MX04 U3694 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][34] ), .A1(\_zzLB[1][34] ), .A2(\_zzLB[2][34] ), .A3(\_zzLB[3][34] ), .Z(odata[2]));
Q_MX04 U3695 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][35] ), .A1(\_zzLB[1][35] ), .A2(\_zzLB[2][35] ), .A3(\_zzLB[3][35] ), .Z(odata[3]));
Q_MX04 U3696 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][36] ), .A1(\_zzLB[1][36] ), .A2(\_zzLB[2][36] ), .A3(\_zzLB[3][36] ), .Z(odata[4]));
Q_MX04 U3697 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][37] ), .A1(\_zzLB[1][37] ), .A2(\_zzLB[2][37] ), .A3(\_zzLB[3][37] ), .Z(odata[5]));
Q_MX04 U3698 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][38] ), .A1(\_zzLB[1][38] ), .A2(\_zzLB[2][38] ), .A3(\_zzLB[3][38] ), .Z(odata[6]));
Q_MX04 U3699 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][39] ), .A1(\_zzLB[1][39] ), .A2(\_zzLB[2][39] ), .A3(\_zzLB[3][39] ), .Z(odata[7]));
Q_MX04 U3700 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][40] ), .A1(\_zzLB[1][40] ), .A2(\_zzLB[2][40] ), .A3(\_zzLB[3][40] ), .Z(odata[8]));
Q_MX04 U3701 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][41] ), .A1(\_zzLB[1][41] ), .A2(\_zzLB[2][41] ), .A3(\_zzLB[3][41] ), .Z(odata[9]));
Q_MX04 U3702 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][42] ), .A1(\_zzLB[1][42] ), .A2(\_zzLB[2][42] ), .A3(\_zzLB[3][42] ), .Z(odata[10]));
Q_MX04 U3703 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][43] ), .A1(\_zzLB[1][43] ), .A2(\_zzLB[2][43] ), .A3(\_zzLB[3][43] ), .Z(odata[11]));
Q_MX04 U3704 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][44] ), .A1(\_zzLB[1][44] ), .A2(\_zzLB[2][44] ), .A3(\_zzLB[3][44] ), .Z(odata[12]));
Q_MX04 U3705 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][45] ), .A1(\_zzLB[1][45] ), .A2(\_zzLB[2][45] ), .A3(\_zzLB[3][45] ), .Z(odata[13]));
Q_MX04 U3706 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][46] ), .A1(\_zzLB[1][46] ), .A2(\_zzLB[2][46] ), .A3(\_zzLB[3][46] ), .Z(odata[14]));
Q_MX04 U3707 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][47] ), .A1(\_zzLB[1][47] ), .A2(\_zzLB[2][47] ), .A3(\_zzLB[3][47] ), .Z(odata[15]));
Q_MX04 U3708 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][48] ), .A1(\_zzLB[1][48] ), .A2(\_zzLB[2][48] ), .A3(\_zzLB[3][48] ), .Z(odata[16]));
Q_MX04 U3709 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][49] ), .A1(\_zzLB[1][49] ), .A2(\_zzLB[2][49] ), .A3(\_zzLB[3][49] ), .Z(odata[17]));
Q_MX04 U3710 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][50] ), .A1(\_zzLB[1][50] ), .A2(\_zzLB[2][50] ), .A3(\_zzLB[3][50] ), .Z(odata[18]));
Q_MX04 U3711 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][51] ), .A1(\_zzLB[1][51] ), .A2(\_zzLB[2][51] ), .A3(\_zzLB[3][51] ), .Z(odata[19]));
Q_MX04 U3712 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][52] ), .A1(\_zzLB[1][52] ), .A2(\_zzLB[2][52] ), .A3(\_zzLB[3][52] ), .Z(odata[20]));
Q_MX04 U3713 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][53] ), .A1(\_zzLB[1][53] ), .A2(\_zzLB[2][53] ), .A3(\_zzLB[3][53] ), .Z(odata[21]));
Q_MX04 U3714 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][54] ), .A1(\_zzLB[1][54] ), .A2(\_zzLB[2][54] ), .A3(\_zzLB[3][54] ), .Z(odata[22]));
Q_MX04 U3715 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][55] ), .A1(\_zzLB[1][55] ), .A2(\_zzLB[2][55] ), .A3(\_zzLB[3][55] ), .Z(odata[23]));
Q_MX04 U3716 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][56] ), .A1(\_zzLB[1][56] ), .A2(\_zzLB[2][56] ), .A3(\_zzLB[3][56] ), .Z(odata[24]));
Q_MX04 U3717 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][57] ), .A1(\_zzLB[1][57] ), .A2(\_zzLB[2][57] ), .A3(\_zzLB[3][57] ), .Z(odata[25]));
Q_MX04 U3718 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][58] ), .A1(\_zzLB[1][58] ), .A2(\_zzLB[2][58] ), .A3(\_zzLB[3][58] ), .Z(odata[26]));
Q_MX04 U3719 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][59] ), .A1(\_zzLB[1][59] ), .A2(\_zzLB[2][59] ), .A3(\_zzLB[3][59] ), .Z(odata[27]));
Q_MX04 U3720 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][60] ), .A1(\_zzLB[1][60] ), .A2(\_zzLB[2][60] ), .A3(\_zzLB[3][60] ), .Z(odata[28]));
Q_MX04 U3721 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][61] ), .A1(\_zzLB[1][61] ), .A2(\_zzLB[2][61] ), .A3(\_zzLB[3][61] ), .Z(odata[29]));
Q_MX04 U3722 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][62] ), .A1(\_zzLB[1][62] ), .A2(\_zzLB[2][62] ), .A3(\_zzLB[3][62] ), .Z(odata[30]));
Q_MX04 U3723 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][63] ), .A1(\_zzLB[1][63] ), .A2(\_zzLB[2][63] ), .A3(\_zzLB[3][63] ), .Z(odata[31]));
Q_MX04 U3724 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][64] ), .A1(\_zzLB[1][64] ), .A2(\_zzLB[2][64] ), .A3(\_zzLB[3][64] ), .Z(odata[32]));
Q_MX04 U3725 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][65] ), .A1(\_zzLB[1][65] ), .A2(\_zzLB[2][65] ), .A3(\_zzLB[3][65] ), .Z(odata[33]));
Q_MX04 U3726 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][66] ), .A1(\_zzLB[1][66] ), .A2(\_zzLB[2][66] ), .A3(\_zzLB[3][66] ), .Z(odata[34]));
Q_MX04 U3727 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][67] ), .A1(\_zzLB[1][67] ), .A2(\_zzLB[2][67] ), .A3(\_zzLB[3][67] ), .Z(odata[35]));
Q_MX04 U3728 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][68] ), .A1(\_zzLB[1][68] ), .A2(\_zzLB[2][68] ), .A3(\_zzLB[3][68] ), .Z(odata[36]));
Q_MX04 U3729 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][69] ), .A1(\_zzLB[1][69] ), .A2(\_zzLB[2][69] ), .A3(\_zzLB[3][69] ), .Z(odata[37]));
Q_MX04 U3730 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][70] ), .A1(\_zzLB[1][70] ), .A2(\_zzLB[2][70] ), .A3(\_zzLB[3][70] ), .Z(odata[38]));
Q_MX04 U3731 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][71] ), .A1(\_zzLB[1][71] ), .A2(\_zzLB[2][71] ), .A3(\_zzLB[3][71] ), .Z(odata[39]));
Q_MX04 U3732 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][72] ), .A1(\_zzLB[1][72] ), .A2(\_zzLB[2][72] ), .A3(\_zzLB[3][72] ), .Z(odata[40]));
Q_MX04 U3733 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][73] ), .A1(\_zzLB[1][73] ), .A2(\_zzLB[2][73] ), .A3(\_zzLB[3][73] ), .Z(odata[41]));
Q_MX04 U3734 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][74] ), .A1(\_zzLB[1][74] ), .A2(\_zzLB[2][74] ), .A3(\_zzLB[3][74] ), .Z(odata[42]));
Q_MX04 U3735 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][75] ), .A1(\_zzLB[1][75] ), .A2(\_zzLB[2][75] ), .A3(\_zzLB[3][75] ), .Z(odata[43]));
Q_MX04 U3736 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][76] ), .A1(\_zzLB[1][76] ), .A2(\_zzLB[2][76] ), .A3(\_zzLB[3][76] ), .Z(odata[44]));
Q_MX04 U3737 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][77] ), .A1(\_zzLB[1][77] ), .A2(\_zzLB[2][77] ), .A3(\_zzLB[3][77] ), .Z(odata[45]));
Q_MX04 U3738 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][78] ), .A1(\_zzLB[1][78] ), .A2(\_zzLB[2][78] ), .A3(\_zzLB[3][78] ), .Z(odata[46]));
Q_MX04 U3739 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][79] ), .A1(\_zzLB[1][79] ), .A2(\_zzLB[2][79] ), .A3(\_zzLB[3][79] ), .Z(odata[47]));
Q_MX04 U3740 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][80] ), .A1(\_zzLB[1][80] ), .A2(\_zzLB[2][80] ), .A3(\_zzLB[3][80] ), .Z(odata[48]));
Q_MX04 U3741 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][81] ), .A1(\_zzLB[1][81] ), .A2(\_zzLB[2][81] ), .A3(\_zzLB[3][81] ), .Z(odata[49]));
Q_MX04 U3742 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][82] ), .A1(\_zzLB[1][82] ), .A2(\_zzLB[2][82] ), .A3(\_zzLB[3][82] ), .Z(odata[50]));
Q_MX04 U3743 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][83] ), .A1(\_zzLB[1][83] ), .A2(\_zzLB[2][83] ), .A3(\_zzLB[3][83] ), .Z(odata[51]));
Q_MX04 U3744 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][84] ), .A1(\_zzLB[1][84] ), .A2(\_zzLB[2][84] ), .A3(\_zzLB[3][84] ), .Z(odata[52]));
Q_MX04 U3745 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][85] ), .A1(\_zzLB[1][85] ), .A2(\_zzLB[2][85] ), .A3(\_zzLB[3][85] ), .Z(odata[53]));
Q_MX04 U3746 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][86] ), .A1(\_zzLB[1][86] ), .A2(\_zzLB[2][86] ), .A3(\_zzLB[3][86] ), .Z(odata[54]));
Q_MX04 U3747 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][87] ), .A1(\_zzLB[1][87] ), .A2(\_zzLB[2][87] ), .A3(\_zzLB[3][87] ), .Z(odata[55]));
Q_MX04 U3748 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][88] ), .A1(\_zzLB[1][88] ), .A2(\_zzLB[2][88] ), .A3(\_zzLB[3][88] ), .Z(odata[56]));
Q_MX04 U3749 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][89] ), .A1(\_zzLB[1][89] ), .A2(\_zzLB[2][89] ), .A3(\_zzLB[3][89] ), .Z(odata[57]));
Q_MX04 U3750 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][90] ), .A1(\_zzLB[1][90] ), .A2(\_zzLB[2][90] ), .A3(\_zzLB[3][90] ), .Z(odata[58]));
Q_MX04 U3751 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][91] ), .A1(\_zzLB[1][91] ), .A2(\_zzLB[2][91] ), .A3(\_zzLB[3][91] ), .Z(odata[59]));
Q_MX04 U3752 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][92] ), .A1(\_zzLB[1][92] ), .A2(\_zzLB[2][92] ), .A3(\_zzLB[3][92] ), .Z(odata[60]));
Q_MX04 U3753 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][93] ), .A1(\_zzLB[1][93] ), .A2(\_zzLB[2][93] ), .A3(\_zzLB[3][93] ), .Z(odata[61]));
Q_MX04 U3754 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][94] ), .A1(\_zzLB[1][94] ), .A2(\_zzLB[2][94] ), .A3(\_zzLB[3][94] ), .Z(odata[62]));
Q_MX04 U3755 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][95] ), .A1(\_zzLB[1][95] ), .A2(\_zzLB[2][95] ), .A3(\_zzLB[3][95] ), .Z(odata[63]));
Q_MX04 U3756 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][96] ), .A1(\_zzLB[1][96] ), .A2(\_zzLB[2][96] ), .A3(\_zzLB[3][96] ), .Z(odata[64]));
Q_MX04 U3757 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][97] ), .A1(\_zzLB[1][97] ), .A2(\_zzLB[2][97] ), .A3(\_zzLB[3][97] ), .Z(odata[65]));
Q_MX04 U3758 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][98] ), .A1(\_zzLB[1][98] ), .A2(\_zzLB[2][98] ), .A3(\_zzLB[3][98] ), .Z(odata[66]));
Q_MX04 U3759 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][99] ), .A1(\_zzLB[1][99] ), .A2(\_zzLB[2][99] ), .A3(\_zzLB[3][99] ), .Z(odata[67]));
Q_MX04 U3760 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][100] ), .A1(\_zzLB[1][100] ), .A2(\_zzLB[2][100] ), .A3(\_zzLB[3][100] ), .Z(odata[68]));
Q_MX04 U3761 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][101] ), .A1(\_zzLB[1][101] ), .A2(\_zzLB[2][101] ), .A3(\_zzLB[3][101] ), .Z(odata[69]));
Q_MX04 U3762 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][102] ), .A1(\_zzLB[1][102] ), .A2(\_zzLB[2][102] ), .A3(\_zzLB[3][102] ), .Z(odata[70]));
Q_MX04 U3763 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][103] ), .A1(\_zzLB[1][103] ), .A2(\_zzLB[2][103] ), .A3(\_zzLB[3][103] ), .Z(odata[71]));
Q_MX04 U3764 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][104] ), .A1(\_zzLB[1][104] ), .A2(\_zzLB[2][104] ), .A3(\_zzLB[3][104] ), .Z(odata[72]));
Q_MX04 U3765 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][105] ), .A1(\_zzLB[1][105] ), .A2(\_zzLB[2][105] ), .A3(\_zzLB[3][105] ), .Z(odata[73]));
Q_MX04 U3766 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][106] ), .A1(\_zzLB[1][106] ), .A2(\_zzLB[2][106] ), .A3(\_zzLB[3][106] ), .Z(odata[74]));
Q_MX04 U3767 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][107] ), .A1(\_zzLB[1][107] ), .A2(\_zzLB[2][107] ), .A3(\_zzLB[3][107] ), .Z(odata[75]));
Q_MX04 U3768 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][108] ), .A1(\_zzLB[1][108] ), .A2(\_zzLB[2][108] ), .A3(\_zzLB[3][108] ), .Z(odata[76]));
Q_MX04 U3769 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][109] ), .A1(\_zzLB[1][109] ), .A2(\_zzLB[2][109] ), .A3(\_zzLB[3][109] ), .Z(odata[77]));
Q_MX04 U3770 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][110] ), .A1(\_zzLB[1][110] ), .A2(\_zzLB[2][110] ), .A3(\_zzLB[3][110] ), .Z(odata[78]));
Q_MX04 U3771 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][111] ), .A1(\_zzLB[1][111] ), .A2(\_zzLB[2][111] ), .A3(\_zzLB[3][111] ), .Z(odata[79]));
Q_MX04 U3772 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][112] ), .A1(\_zzLB[1][112] ), .A2(\_zzLB[2][112] ), .A3(\_zzLB[3][112] ), .Z(odata[80]));
Q_MX04 U3773 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][113] ), .A1(\_zzLB[1][113] ), .A2(\_zzLB[2][113] ), .A3(\_zzLB[3][113] ), .Z(odata[81]));
Q_MX04 U3774 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][114] ), .A1(\_zzLB[1][114] ), .A2(\_zzLB[2][114] ), .A3(\_zzLB[3][114] ), .Z(odata[82]));
Q_MX04 U3775 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][115] ), .A1(\_zzLB[1][115] ), .A2(\_zzLB[2][115] ), .A3(\_zzLB[3][115] ), .Z(odata[83]));
Q_MX04 U3776 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][116] ), .A1(\_zzLB[1][116] ), .A2(\_zzLB[2][116] ), .A3(\_zzLB[3][116] ), .Z(odata[84]));
Q_MX04 U3777 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][117] ), .A1(\_zzLB[1][117] ), .A2(\_zzLB[2][117] ), .A3(\_zzLB[3][117] ), .Z(odata[85]));
Q_MX04 U3778 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][118] ), .A1(\_zzLB[1][118] ), .A2(\_zzLB[2][118] ), .A3(\_zzLB[3][118] ), .Z(odata[86]));
Q_MX04 U3779 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][119] ), .A1(\_zzLB[1][119] ), .A2(\_zzLB[2][119] ), .A3(\_zzLB[3][119] ), .Z(odata[87]));
Q_MX04 U3780 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][120] ), .A1(\_zzLB[1][120] ), .A2(\_zzLB[2][120] ), .A3(\_zzLB[3][120] ), .Z(odata[88]));
Q_MX04 U3781 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][121] ), .A1(\_zzLB[1][121] ), .A2(\_zzLB[2][121] ), .A3(\_zzLB[3][121] ), .Z(odata[89]));
Q_MX04 U3782 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][122] ), .A1(\_zzLB[1][122] ), .A2(\_zzLB[2][122] ), .A3(\_zzLB[3][122] ), .Z(odata[90]));
Q_MX04 U3783 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][123] ), .A1(\_zzLB[1][123] ), .A2(\_zzLB[2][123] ), .A3(\_zzLB[3][123] ), .Z(odata[91]));
Q_MX04 U3784 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][124] ), .A1(\_zzLB[1][124] ), .A2(\_zzLB[2][124] ), .A3(\_zzLB[3][124] ), .Z(odata[92]));
Q_MX04 U3785 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][125] ), .A1(\_zzLB[1][125] ), .A2(\_zzLB[2][125] ), .A3(\_zzLB[3][125] ), .Z(odata[93]));
Q_MX04 U3786 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][126] ), .A1(\_zzLB[1][126] ), .A2(\_zzLB[2][126] ), .A3(\_zzLB[3][126] ), .Z(odata[94]));
Q_MX04 U3787 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][127] ), .A1(\_zzLB[1][127] ), .A2(\_zzLB[2][127] ), .A3(\_zzLB[3][127] ), .Z(odata[95]));
Q_MX04 U3788 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][128] ), .A1(\_zzLB[1][128] ), .A2(\_zzLB[2][128] ), .A3(\_zzLB[3][128] ), .Z(odata[96]));
Q_MX04 U3789 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][129] ), .A1(\_zzLB[1][129] ), .A2(\_zzLB[2][129] ), .A3(\_zzLB[3][129] ), .Z(odata[97]));
Q_MX04 U3790 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][130] ), .A1(\_zzLB[1][130] ), .A2(\_zzLB[2][130] ), .A3(\_zzLB[3][130] ), .Z(odata[98]));
Q_MX04 U3791 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][131] ), .A1(\_zzLB[1][131] ), .A2(\_zzLB[2][131] ), .A3(\_zzLB[3][131] ), .Z(odata[99]));
Q_MX04 U3792 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][132] ), .A1(\_zzLB[1][132] ), .A2(\_zzLB[2][132] ), .A3(\_zzLB[3][132] ), .Z(odata[100]));
Q_MX04 U3793 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][133] ), .A1(\_zzLB[1][133] ), .A2(\_zzLB[2][133] ), .A3(\_zzLB[3][133] ), .Z(odata[101]));
Q_MX04 U3794 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][134] ), .A1(\_zzLB[1][134] ), .A2(\_zzLB[2][134] ), .A3(\_zzLB[3][134] ), .Z(odata[102]));
Q_MX04 U3795 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][135] ), .A1(\_zzLB[1][135] ), .A2(\_zzLB[2][135] ), .A3(\_zzLB[3][135] ), .Z(odata[103]));
Q_MX04 U3796 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][136] ), .A1(\_zzLB[1][136] ), .A2(\_zzLB[2][136] ), .A3(\_zzLB[3][136] ), .Z(odata[104]));
Q_MX04 U3797 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][137] ), .A1(\_zzLB[1][137] ), .A2(\_zzLB[2][137] ), .A3(\_zzLB[3][137] ), .Z(odata[105]));
Q_MX04 U3798 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][138] ), .A1(\_zzLB[1][138] ), .A2(\_zzLB[2][138] ), .A3(\_zzLB[3][138] ), .Z(odata[106]));
Q_MX04 U3799 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][139] ), .A1(\_zzLB[1][139] ), .A2(\_zzLB[2][139] ), .A3(\_zzLB[3][139] ), .Z(odata[107]));
Q_MX04 U3800 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][140] ), .A1(\_zzLB[1][140] ), .A2(\_zzLB[2][140] ), .A3(\_zzLB[3][140] ), .Z(odata[108]));
Q_MX04 U3801 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][141] ), .A1(\_zzLB[1][141] ), .A2(\_zzLB[2][141] ), .A3(\_zzLB[3][141] ), .Z(odata[109]));
Q_MX04 U3802 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][142] ), .A1(\_zzLB[1][142] ), .A2(\_zzLB[2][142] ), .A3(\_zzLB[3][142] ), .Z(odata[110]));
Q_MX04 U3803 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][143] ), .A1(\_zzLB[1][143] ), .A2(\_zzLB[2][143] ), .A3(\_zzLB[3][143] ), .Z(odata[111]));
Q_MX04 U3804 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][144] ), .A1(\_zzLB[1][144] ), .A2(\_zzLB[2][144] ), .A3(\_zzLB[3][144] ), .Z(odata[112]));
Q_MX04 U3805 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][145] ), .A1(\_zzLB[1][145] ), .A2(\_zzLB[2][145] ), .A3(\_zzLB[3][145] ), .Z(odata[113]));
Q_MX04 U3806 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][146] ), .A1(\_zzLB[1][146] ), .A2(\_zzLB[2][146] ), .A3(\_zzLB[3][146] ), .Z(odata[114]));
Q_MX04 U3807 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][147] ), .A1(\_zzLB[1][147] ), .A2(\_zzLB[2][147] ), .A3(\_zzLB[3][147] ), .Z(odata[115]));
Q_MX04 U3808 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][148] ), .A1(\_zzLB[1][148] ), .A2(\_zzLB[2][148] ), .A3(\_zzLB[3][148] ), .Z(odata[116]));
Q_MX04 U3809 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][149] ), .A1(\_zzLB[1][149] ), .A2(\_zzLB[2][149] ), .A3(\_zzLB[3][149] ), .Z(odata[117]));
Q_MX04 U3810 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][150] ), .A1(\_zzLB[1][150] ), .A2(\_zzLB[2][150] ), .A3(\_zzLB[3][150] ), .Z(odata[118]));
Q_MX04 U3811 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][151] ), .A1(\_zzLB[1][151] ), .A2(\_zzLB[2][151] ), .A3(\_zzLB[3][151] ), .Z(odata[119]));
Q_MX04 U3812 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][152] ), .A1(\_zzLB[1][152] ), .A2(\_zzLB[2][152] ), .A3(\_zzLB[3][152] ), .Z(odata[120]));
Q_MX04 U3813 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][153] ), .A1(\_zzLB[1][153] ), .A2(\_zzLB[2][153] ), .A3(\_zzLB[3][153] ), .Z(odata[121]));
Q_MX04 U3814 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][154] ), .A1(\_zzLB[1][154] ), .A2(\_zzLB[2][154] ), .A3(\_zzLB[3][154] ), .Z(odata[122]));
Q_MX04 U3815 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][155] ), .A1(\_zzLB[1][155] ), .A2(\_zzLB[2][155] ), .A3(\_zzLB[3][155] ), .Z(odata[123]));
Q_MX04 U3816 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][156] ), .A1(\_zzLB[1][156] ), .A2(\_zzLB[2][156] ), .A3(\_zzLB[3][156] ), .Z(odata[124]));
Q_MX04 U3817 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][157] ), .A1(\_zzLB[1][157] ), .A2(\_zzLB[2][157] ), .A3(\_zzLB[3][157] ), .Z(odata[125]));
Q_MX04 U3818 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][158] ), .A1(\_zzLB[1][158] ), .A2(\_zzLB[2][158] ), .A3(\_zzLB[3][158] ), .Z(odata[126]));
Q_MX04 U3819 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][159] ), .A1(\_zzLB[1][159] ), .A2(\_zzLB[2][159] ), .A3(\_zzLB[3][159] ), .Z(odata[127]));
Q_MX04 U3820 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][160] ), .A1(\_zzLB[1][160] ), .A2(\_zzLB[2][160] ), .A3(\_zzLB[3][160] ), .Z(odata[128]));
Q_MX04 U3821 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][161] ), .A1(\_zzLB[1][161] ), .A2(\_zzLB[2][161] ), .A3(\_zzLB[3][161] ), .Z(odata[129]));
Q_MX04 U3822 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][162] ), .A1(\_zzLB[1][162] ), .A2(\_zzLB[2][162] ), .A3(\_zzLB[3][162] ), .Z(odata[130]));
Q_MX04 U3823 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][163] ), .A1(\_zzLB[1][163] ), .A2(\_zzLB[2][163] ), .A3(\_zzLB[3][163] ), .Z(odata[131]));
Q_MX04 U3824 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][164] ), .A1(\_zzLB[1][164] ), .A2(\_zzLB[2][164] ), .A3(\_zzLB[3][164] ), .Z(odata[132]));
Q_MX04 U3825 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][165] ), .A1(\_zzLB[1][165] ), .A2(\_zzLB[2][165] ), .A3(\_zzLB[3][165] ), .Z(odata[133]));
Q_MX04 U3826 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][166] ), .A1(\_zzLB[1][166] ), .A2(\_zzLB[2][166] ), .A3(\_zzLB[3][166] ), .Z(odata[134]));
Q_MX04 U3827 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][167] ), .A1(\_zzLB[1][167] ), .A2(\_zzLB[2][167] ), .A3(\_zzLB[3][167] ), .Z(odata[135]));
Q_MX04 U3828 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][168] ), .A1(\_zzLB[1][168] ), .A2(\_zzLB[2][168] ), .A3(\_zzLB[3][168] ), .Z(odata[136]));
Q_MX04 U3829 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][169] ), .A1(\_zzLB[1][169] ), .A2(\_zzLB[2][169] ), .A3(\_zzLB[3][169] ), .Z(odata[137]));
Q_MX04 U3830 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][170] ), .A1(\_zzLB[1][170] ), .A2(\_zzLB[2][170] ), .A3(\_zzLB[3][170] ), .Z(odata[138]));
Q_MX04 U3831 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][171] ), .A1(\_zzLB[1][171] ), .A2(\_zzLB[2][171] ), .A3(\_zzLB[3][171] ), .Z(odata[139]));
Q_MX04 U3832 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][172] ), .A1(\_zzLB[1][172] ), .A2(\_zzLB[2][172] ), .A3(\_zzLB[3][172] ), .Z(odata[140]));
Q_MX04 U3833 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][173] ), .A1(\_zzLB[1][173] ), .A2(\_zzLB[2][173] ), .A3(\_zzLB[3][173] ), .Z(odata[141]));
Q_MX04 U3834 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][174] ), .A1(\_zzLB[1][174] ), .A2(\_zzLB[2][174] ), .A3(\_zzLB[3][174] ), .Z(odata[142]));
Q_MX04 U3835 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][175] ), .A1(\_zzLB[1][175] ), .A2(\_zzLB[2][175] ), .A3(\_zzLB[3][175] ), .Z(odata[143]));
Q_MX04 U3836 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][176] ), .A1(\_zzLB[1][176] ), .A2(\_zzLB[2][176] ), .A3(\_zzLB[3][176] ), .Z(odata[144]));
Q_MX04 U3837 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][177] ), .A1(\_zzLB[1][177] ), .A2(\_zzLB[2][177] ), .A3(\_zzLB[3][177] ), .Z(odata[145]));
Q_MX04 U3838 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][178] ), .A1(\_zzLB[1][178] ), .A2(\_zzLB[2][178] ), .A3(\_zzLB[3][178] ), .Z(odata[146]));
Q_MX04 U3839 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][179] ), .A1(\_zzLB[1][179] ), .A2(\_zzLB[2][179] ), .A3(\_zzLB[3][179] ), .Z(odata[147]));
Q_MX04 U3840 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][180] ), .A1(\_zzLB[1][180] ), .A2(\_zzLB[2][180] ), .A3(\_zzLB[3][180] ), .Z(odata[148]));
Q_MX04 U3841 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][181] ), .A1(\_zzLB[1][181] ), .A2(\_zzLB[2][181] ), .A3(\_zzLB[3][181] ), .Z(odata[149]));
Q_MX04 U3842 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][182] ), .A1(\_zzLB[1][182] ), .A2(\_zzLB[2][182] ), .A3(\_zzLB[3][182] ), .Z(odata[150]));
Q_MX04 U3843 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][183] ), .A1(\_zzLB[1][183] ), .A2(\_zzLB[2][183] ), .A3(\_zzLB[3][183] ), .Z(odata[151]));
Q_MX04 U3844 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][184] ), .A1(\_zzLB[1][184] ), .A2(\_zzLB[2][184] ), .A3(\_zzLB[3][184] ), .Z(odata[152]));
Q_MX04 U3845 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][185] ), .A1(\_zzLB[1][185] ), .A2(\_zzLB[2][185] ), .A3(\_zzLB[3][185] ), .Z(odata[153]));
Q_MX04 U3846 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][186] ), .A1(\_zzLB[1][186] ), .A2(\_zzLB[2][186] ), .A3(\_zzLB[3][186] ), .Z(odata[154]));
Q_MX04 U3847 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][187] ), .A1(\_zzLB[1][187] ), .A2(\_zzLB[2][187] ), .A3(\_zzLB[3][187] ), .Z(odata[155]));
Q_MX04 U3848 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][188] ), .A1(\_zzLB[1][188] ), .A2(\_zzLB[2][188] ), .A3(\_zzLB[3][188] ), .Z(odata[156]));
Q_MX04 U3849 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][189] ), .A1(\_zzLB[1][189] ), .A2(\_zzLB[2][189] ), .A3(\_zzLB[3][189] ), .Z(odata[157]));
Q_MX04 U3850 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][190] ), .A1(\_zzLB[1][190] ), .A2(\_zzLB[2][190] ), .A3(\_zzLB[3][190] ), .Z(odata[158]));
Q_MX04 U3851 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][191] ), .A1(\_zzLB[1][191] ), .A2(\_zzLB[2][191] ), .A3(\_zzLB[3][191] ), .Z(odata[159]));
Q_MX04 U3852 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][192] ), .A1(\_zzLB[1][192] ), .A2(\_zzLB[2][192] ), .A3(\_zzLB[3][192] ), .Z(odata[160]));
Q_MX04 U3853 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][193] ), .A1(\_zzLB[1][193] ), .A2(\_zzLB[2][193] ), .A3(\_zzLB[3][193] ), .Z(odata[161]));
Q_MX04 U3854 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][194] ), .A1(\_zzLB[1][194] ), .A2(\_zzLB[2][194] ), .A3(\_zzLB[3][194] ), .Z(odata[162]));
Q_MX04 U3855 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][195] ), .A1(\_zzLB[1][195] ), .A2(\_zzLB[2][195] ), .A3(\_zzLB[3][195] ), .Z(odata[163]));
Q_MX04 U3856 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][196] ), .A1(\_zzLB[1][196] ), .A2(\_zzLB[2][196] ), .A3(\_zzLB[3][196] ), .Z(odata[164]));
Q_MX04 U3857 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][197] ), .A1(\_zzLB[1][197] ), .A2(\_zzLB[2][197] ), .A3(\_zzLB[3][197] ), .Z(odata[165]));
Q_MX04 U3858 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][198] ), .A1(\_zzLB[1][198] ), .A2(\_zzLB[2][198] ), .A3(\_zzLB[3][198] ), .Z(odata[166]));
Q_MX04 U3859 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][199] ), .A1(\_zzLB[1][199] ), .A2(\_zzLB[2][199] ), .A3(\_zzLB[3][199] ), .Z(odata[167]));
Q_MX04 U3860 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][200] ), .A1(\_zzLB[1][200] ), .A2(\_zzLB[2][200] ), .A3(\_zzLB[3][200] ), .Z(odata[168]));
Q_MX04 U3861 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][201] ), .A1(\_zzLB[1][201] ), .A2(\_zzLB[2][201] ), .A3(\_zzLB[3][201] ), .Z(odata[169]));
Q_MX04 U3862 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][202] ), .A1(\_zzLB[1][202] ), .A2(\_zzLB[2][202] ), .A3(\_zzLB[3][202] ), .Z(odata[170]));
Q_MX04 U3863 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][203] ), .A1(\_zzLB[1][203] ), .A2(\_zzLB[2][203] ), .A3(\_zzLB[3][203] ), .Z(odata[171]));
Q_MX04 U3864 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][204] ), .A1(\_zzLB[1][204] ), .A2(\_zzLB[2][204] ), .A3(\_zzLB[3][204] ), .Z(odata[172]));
Q_MX04 U3865 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][205] ), .A1(\_zzLB[1][205] ), .A2(\_zzLB[2][205] ), .A3(\_zzLB[3][205] ), .Z(odata[173]));
Q_MX04 U3866 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][206] ), .A1(\_zzLB[1][206] ), .A2(\_zzLB[2][206] ), .A3(\_zzLB[3][206] ), .Z(odata[174]));
Q_MX04 U3867 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][207] ), .A1(\_zzLB[1][207] ), .A2(\_zzLB[2][207] ), .A3(\_zzLB[3][207] ), .Z(odata[175]));
Q_MX04 U3868 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][208] ), .A1(\_zzLB[1][208] ), .A2(\_zzLB[2][208] ), .A3(\_zzLB[3][208] ), .Z(odata[176]));
Q_MX04 U3869 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][209] ), .A1(\_zzLB[1][209] ), .A2(\_zzLB[2][209] ), .A3(\_zzLB[3][209] ), .Z(odata[177]));
Q_MX04 U3870 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][210] ), .A1(\_zzLB[1][210] ), .A2(\_zzLB[2][210] ), .A3(\_zzLB[3][210] ), .Z(odata[178]));
Q_MX04 U3871 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][211] ), .A1(\_zzLB[1][211] ), .A2(\_zzLB[2][211] ), .A3(\_zzLB[3][211] ), .Z(odata[179]));
Q_MX04 U3872 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][212] ), .A1(\_zzLB[1][212] ), .A2(\_zzLB[2][212] ), .A3(\_zzLB[3][212] ), .Z(odata[180]));
Q_MX04 U3873 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][213] ), .A1(\_zzLB[1][213] ), .A2(\_zzLB[2][213] ), .A3(\_zzLB[3][213] ), .Z(odata[181]));
Q_MX04 U3874 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][214] ), .A1(\_zzLB[1][214] ), .A2(\_zzLB[2][214] ), .A3(\_zzLB[3][214] ), .Z(odata[182]));
Q_MX04 U3875 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][215] ), .A1(\_zzLB[1][215] ), .A2(\_zzLB[2][215] ), .A3(\_zzLB[3][215] ), .Z(odata[183]));
Q_MX04 U3876 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][216] ), .A1(\_zzLB[1][216] ), .A2(\_zzLB[2][216] ), .A3(\_zzLB[3][216] ), .Z(odata[184]));
Q_MX04 U3877 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][217] ), .A1(\_zzLB[1][217] ), .A2(\_zzLB[2][217] ), .A3(\_zzLB[3][217] ), .Z(odata[185]));
Q_MX04 U3878 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][218] ), .A1(\_zzLB[1][218] ), .A2(\_zzLB[2][218] ), .A3(\_zzLB[3][218] ), .Z(odata[186]));
Q_MX04 U3879 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][219] ), .A1(\_zzLB[1][219] ), .A2(\_zzLB[2][219] ), .A3(\_zzLB[3][219] ), .Z(odata[187]));
Q_MX04 U3880 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][220] ), .A1(\_zzLB[1][220] ), .A2(\_zzLB[2][220] ), .A3(\_zzLB[3][220] ), .Z(odata[188]));
Q_MX04 U3881 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][221] ), .A1(\_zzLB[1][221] ), .A2(\_zzLB[2][221] ), .A3(\_zzLB[3][221] ), .Z(odata[189]));
Q_MX04 U3882 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][222] ), .A1(\_zzLB[1][222] ), .A2(\_zzLB[2][222] ), .A3(\_zzLB[3][222] ), .Z(odata[190]));
Q_MX04 U3883 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][223] ), .A1(\_zzLB[1][223] ), .A2(\_zzLB[2][223] ), .A3(\_zzLB[3][223] ), .Z(odata[191]));
Q_MX04 U3884 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][224] ), .A1(\_zzLB[1][224] ), .A2(\_zzLB[2][224] ), .A3(\_zzLB[3][224] ), .Z(odata[192]));
Q_MX04 U3885 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][225] ), .A1(\_zzLB[1][225] ), .A2(\_zzLB[2][225] ), .A3(\_zzLB[3][225] ), .Z(odata[193]));
Q_MX04 U3886 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][226] ), .A1(\_zzLB[1][226] ), .A2(\_zzLB[2][226] ), .A3(\_zzLB[3][226] ), .Z(odata[194]));
Q_MX04 U3887 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][227] ), .A1(\_zzLB[1][227] ), .A2(\_zzLB[2][227] ), .A3(\_zzLB[3][227] ), .Z(odata[195]));
Q_MX04 U3888 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][228] ), .A1(\_zzLB[1][228] ), .A2(\_zzLB[2][228] ), .A3(\_zzLB[3][228] ), .Z(odata[196]));
Q_MX04 U3889 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][229] ), .A1(\_zzLB[1][229] ), .A2(\_zzLB[2][229] ), .A3(\_zzLB[3][229] ), .Z(odata[197]));
Q_MX04 U3890 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][230] ), .A1(\_zzLB[1][230] ), .A2(\_zzLB[2][230] ), .A3(\_zzLB[3][230] ), .Z(odata[198]));
Q_MX04 U3891 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][231] ), .A1(\_zzLB[1][231] ), .A2(\_zzLB[2][231] ), .A3(\_zzLB[3][231] ), .Z(odata[199]));
Q_MX04 U3892 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][232] ), .A1(\_zzLB[1][232] ), .A2(\_zzLB[2][232] ), .A3(\_zzLB[3][232] ), .Z(odata[200]));
Q_MX04 U3893 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][233] ), .A1(\_zzLB[1][233] ), .A2(\_zzLB[2][233] ), .A3(\_zzLB[3][233] ), .Z(odata[201]));
Q_MX04 U3894 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][234] ), .A1(\_zzLB[1][234] ), .A2(\_zzLB[2][234] ), .A3(\_zzLB[3][234] ), .Z(odata[202]));
Q_MX04 U3895 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][235] ), .A1(\_zzLB[1][235] ), .A2(\_zzLB[2][235] ), .A3(\_zzLB[3][235] ), .Z(odata[203]));
Q_MX04 U3896 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][236] ), .A1(\_zzLB[1][236] ), .A2(\_zzLB[2][236] ), .A3(\_zzLB[3][236] ), .Z(odata[204]));
Q_MX04 U3897 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][237] ), .A1(\_zzLB[1][237] ), .A2(\_zzLB[2][237] ), .A3(\_zzLB[3][237] ), .Z(odata[205]));
Q_MX04 U3898 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][238] ), .A1(\_zzLB[1][238] ), .A2(\_zzLB[2][238] ), .A3(\_zzLB[3][238] ), .Z(odata[206]));
Q_MX04 U3899 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][239] ), .A1(\_zzLB[1][239] ), .A2(\_zzLB[2][239] ), .A3(\_zzLB[3][239] ), .Z(odata[207]));
Q_MX04 U3900 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][240] ), .A1(\_zzLB[1][240] ), .A2(\_zzLB[2][240] ), .A3(\_zzLB[3][240] ), .Z(odata[208]));
Q_MX04 U3901 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][241] ), .A1(\_zzLB[1][241] ), .A2(\_zzLB[2][241] ), .A3(\_zzLB[3][241] ), .Z(odata[209]));
Q_MX04 U3902 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][242] ), .A1(\_zzLB[1][242] ), .A2(\_zzLB[2][242] ), .A3(\_zzLB[3][242] ), .Z(odata[210]));
Q_MX04 U3903 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][243] ), .A1(\_zzLB[1][243] ), .A2(\_zzLB[2][243] ), .A3(\_zzLB[3][243] ), .Z(odata[211]));
Q_MX04 U3904 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][244] ), .A1(\_zzLB[1][244] ), .A2(\_zzLB[2][244] ), .A3(\_zzLB[3][244] ), .Z(odata[212]));
Q_MX04 U3905 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][245] ), .A1(\_zzLB[1][245] ), .A2(\_zzLB[2][245] ), .A3(\_zzLB[3][245] ), .Z(odata[213]));
Q_MX04 U3906 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][246] ), .A1(\_zzLB[1][246] ), .A2(\_zzLB[2][246] ), .A3(\_zzLB[3][246] ), .Z(odata[214]));
Q_MX04 U3907 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][247] ), .A1(\_zzLB[1][247] ), .A2(\_zzLB[2][247] ), .A3(\_zzLB[3][247] ), .Z(odata[215]));
Q_MX04 U3908 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][248] ), .A1(\_zzLB[1][248] ), .A2(\_zzLB[2][248] ), .A3(\_zzLB[3][248] ), .Z(odata[216]));
Q_MX04 U3909 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][249] ), .A1(\_zzLB[1][249] ), .A2(\_zzLB[2][249] ), .A3(\_zzLB[3][249] ), .Z(odata[217]));
Q_MX04 U3910 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][250] ), .A1(\_zzLB[1][250] ), .A2(\_zzLB[2][250] ), .A3(\_zzLB[3][250] ), .Z(odata[218]));
Q_MX04 U3911 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][251] ), .A1(\_zzLB[1][251] ), .A2(\_zzLB[2][251] ), .A3(\_zzLB[3][251] ), .Z(odata[219]));
Q_MX04 U3912 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][252] ), .A1(\_zzLB[1][252] ), .A2(\_zzLB[2][252] ), .A3(\_zzLB[3][252] ), .Z(odata[220]));
Q_MX04 U3913 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][253] ), .A1(\_zzLB[1][253] ), .A2(\_zzLB[2][253] ), .A3(\_zzLB[3][253] ), .Z(odata[221]));
Q_MX04 U3914 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][254] ), .A1(\_zzLB[1][254] ), .A2(\_zzLB[2][254] ), .A3(\_zzLB[3][254] ), .Z(odata[222]));
Q_MX04 U3915 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][255] ), .A1(\_zzLB[1][255] ), .A2(\_zzLB[2][255] ), .A3(\_zzLB[3][255] ), .Z(odata[223]));
Q_MX04 U3916 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][256] ), .A1(\_zzLB[1][256] ), .A2(\_zzLB[2][256] ), .A3(\_zzLB[3][256] ), .Z(odata[224]));
Q_MX04 U3917 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][257] ), .A1(\_zzLB[1][257] ), .A2(\_zzLB[2][257] ), .A3(\_zzLB[3][257] ), .Z(odata[225]));
Q_MX04 U3918 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][258] ), .A1(\_zzLB[1][258] ), .A2(\_zzLB[2][258] ), .A3(\_zzLB[3][258] ), .Z(odata[226]));
Q_MX04 U3919 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][259] ), .A1(\_zzLB[1][259] ), .A2(\_zzLB[2][259] ), .A3(\_zzLB[3][259] ), .Z(odata[227]));
Q_MX04 U3920 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][260] ), .A1(\_zzLB[1][260] ), .A2(\_zzLB[2][260] ), .A3(\_zzLB[3][260] ), .Z(odata[228]));
Q_MX04 U3921 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][261] ), .A1(\_zzLB[1][261] ), .A2(\_zzLB[2][261] ), .A3(\_zzLB[3][261] ), .Z(odata[229]));
Q_MX04 U3922 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][262] ), .A1(\_zzLB[1][262] ), .A2(\_zzLB[2][262] ), .A3(\_zzLB[3][262] ), .Z(odata[230]));
Q_MX04 U3923 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][263] ), .A1(\_zzLB[1][263] ), .A2(\_zzLB[2][263] ), .A3(\_zzLB[3][263] ), .Z(odata[231]));
Q_MX04 U3924 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][264] ), .A1(\_zzLB[1][264] ), .A2(\_zzLB[2][264] ), .A3(\_zzLB[3][264] ), .Z(odata[232]));
Q_MX04 U3925 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][265] ), .A1(\_zzLB[1][265] ), .A2(\_zzLB[2][265] ), .A3(\_zzLB[3][265] ), .Z(odata[233]));
Q_MX04 U3926 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][266] ), .A1(\_zzLB[1][266] ), .A2(\_zzLB[2][266] ), .A3(\_zzLB[3][266] ), .Z(odata[234]));
Q_MX04 U3927 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][267] ), .A1(\_zzLB[1][267] ), .A2(\_zzLB[2][267] ), .A3(\_zzLB[3][267] ), .Z(odata[235]));
Q_MX04 U3928 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][268] ), .A1(\_zzLB[1][268] ), .A2(\_zzLB[2][268] ), .A3(\_zzLB[3][268] ), .Z(odata[236]));
Q_MX04 U3929 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][269] ), .A1(\_zzLB[1][269] ), .A2(\_zzLB[2][269] ), .A3(\_zzLB[3][269] ), .Z(odata[237]));
Q_MX04 U3930 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][270] ), .A1(\_zzLB[1][270] ), .A2(\_zzLB[2][270] ), .A3(\_zzLB[3][270] ), .Z(odata[238]));
Q_MX04 U3931 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][271] ), .A1(\_zzLB[1][271] ), .A2(\_zzLB[2][271] ), .A3(\_zzLB[3][271] ), .Z(odata[239]));
Q_MX04 U3932 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][272] ), .A1(\_zzLB[1][272] ), .A2(\_zzLB[2][272] ), .A3(\_zzLB[3][272] ), .Z(odata[240]));
Q_MX04 U3933 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][273] ), .A1(\_zzLB[1][273] ), .A2(\_zzLB[2][273] ), .A3(\_zzLB[3][273] ), .Z(odata[241]));
Q_MX04 U3934 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][274] ), .A1(\_zzLB[1][274] ), .A2(\_zzLB[2][274] ), .A3(\_zzLB[3][274] ), .Z(odata[242]));
Q_MX04 U3935 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][275] ), .A1(\_zzLB[1][275] ), .A2(\_zzLB[2][275] ), .A3(\_zzLB[3][275] ), .Z(odata[243]));
Q_MX04 U3936 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][276] ), .A1(\_zzLB[1][276] ), .A2(\_zzLB[2][276] ), .A3(\_zzLB[3][276] ), .Z(odata[244]));
Q_MX04 U3937 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][277] ), .A1(\_zzLB[1][277] ), .A2(\_zzLB[2][277] ), .A3(\_zzLB[3][277] ), .Z(odata[245]));
Q_MX04 U3938 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][278] ), .A1(\_zzLB[1][278] ), .A2(\_zzLB[2][278] ), .A3(\_zzLB[3][278] ), .Z(odata[246]));
Q_MX04 U3939 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][279] ), .A1(\_zzLB[1][279] ), .A2(\_zzLB[2][279] ), .A3(\_zzLB[3][279] ), .Z(odata[247]));
Q_MX04 U3940 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][280] ), .A1(\_zzLB[1][280] ), .A2(\_zzLB[2][280] ), .A3(\_zzLB[3][280] ), .Z(odata[248]));
Q_MX04 U3941 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][281] ), .A1(\_zzLB[1][281] ), .A2(\_zzLB[2][281] ), .A3(\_zzLB[3][281] ), .Z(odata[249]));
Q_MX04 U3942 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][282] ), .A1(\_zzLB[1][282] ), .A2(\_zzLB[2][282] ), .A3(\_zzLB[3][282] ), .Z(odata[250]));
Q_MX04 U3943 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][283] ), .A1(\_zzLB[1][283] ), .A2(\_zzLB[2][283] ), .A3(\_zzLB[3][283] ), .Z(odata[251]));
Q_MX04 U3944 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][284] ), .A1(\_zzLB[1][284] ), .A2(\_zzLB[2][284] ), .A3(\_zzLB[3][284] ), .Z(odata[252]));
Q_MX04 U3945 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][285] ), .A1(\_zzLB[1][285] ), .A2(\_zzLB[2][285] ), .A3(\_zzLB[3][285] ), .Z(odata[253]));
Q_MX04 U3946 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][286] ), .A1(\_zzLB[1][286] ), .A2(\_zzLB[2][286] ), .A3(\_zzLB[3][286] ), .Z(odata[254]));
Q_MX04 U3947 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][287] ), .A1(\_zzLB[1][287] ), .A2(\_zzLB[2][287] ), .A3(\_zzLB[3][287] ), .Z(odata[255]));
Q_MX04 U3948 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][288] ), .A1(\_zzLB[1][288] ), .A2(\_zzLB[2][288] ), .A3(\_zzLB[3][288] ), .Z(odata[256]));
Q_MX04 U3949 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][289] ), .A1(\_zzLB[1][289] ), .A2(\_zzLB[2][289] ), .A3(\_zzLB[3][289] ), .Z(odata[257]));
Q_MX04 U3950 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][290] ), .A1(\_zzLB[1][290] ), .A2(\_zzLB[2][290] ), .A3(\_zzLB[3][290] ), .Z(odata[258]));
Q_MX04 U3951 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][291] ), .A1(\_zzLB[1][291] ), .A2(\_zzLB[2][291] ), .A3(\_zzLB[3][291] ), .Z(odata[259]));
Q_MX04 U3952 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][292] ), .A1(\_zzLB[1][292] ), .A2(\_zzLB[2][292] ), .A3(\_zzLB[3][292] ), .Z(odata[260]));
Q_MX04 U3953 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][293] ), .A1(\_zzLB[1][293] ), .A2(\_zzLB[2][293] ), .A3(\_zzLB[3][293] ), .Z(odata[261]));
Q_MX04 U3954 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][294] ), .A1(\_zzLB[1][294] ), .A2(\_zzLB[2][294] ), .A3(\_zzLB[3][294] ), .Z(odata[262]));
Q_MX04 U3955 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][295] ), .A1(\_zzLB[1][295] ), .A2(\_zzLB[2][295] ), .A3(\_zzLB[3][295] ), .Z(odata[263]));
Q_MX04 U3956 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][296] ), .A1(\_zzLB[1][296] ), .A2(\_zzLB[2][296] ), .A3(\_zzLB[3][296] ), .Z(odata[264]));
Q_MX04 U3957 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][297] ), .A1(\_zzLB[1][297] ), .A2(\_zzLB[2][297] ), .A3(\_zzLB[3][297] ), .Z(odata[265]));
Q_MX04 U3958 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][298] ), .A1(\_zzLB[1][298] ), .A2(\_zzLB[2][298] ), .A3(\_zzLB[3][298] ), .Z(odata[266]));
Q_MX04 U3959 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][299] ), .A1(\_zzLB[1][299] ), .A2(\_zzLB[2][299] ), .A3(\_zzLB[3][299] ), .Z(odata[267]));
Q_MX04 U3960 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][300] ), .A1(\_zzLB[1][300] ), .A2(\_zzLB[2][300] ), .A3(\_zzLB[3][300] ), .Z(odata[268]));
Q_MX04 U3961 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][301] ), .A1(\_zzLB[1][301] ), .A2(\_zzLB[2][301] ), .A3(\_zzLB[3][301] ), .Z(odata[269]));
Q_MX04 U3962 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][302] ), .A1(\_zzLB[1][302] ), .A2(\_zzLB[2][302] ), .A3(\_zzLB[3][302] ), .Z(odata[270]));
Q_MX04 U3963 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][303] ), .A1(\_zzLB[1][303] ), .A2(\_zzLB[2][303] ), .A3(\_zzLB[3][303] ), .Z(odata[271]));
Q_MX04 U3964 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][304] ), .A1(\_zzLB[1][304] ), .A2(\_zzLB[2][304] ), .A3(\_zzLB[3][304] ), .Z(odata[272]));
Q_MX04 U3965 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][305] ), .A1(\_zzLB[1][305] ), .A2(\_zzLB[2][305] ), .A3(\_zzLB[3][305] ), .Z(odata[273]));
Q_MX04 U3966 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][306] ), .A1(\_zzLB[1][306] ), .A2(\_zzLB[2][306] ), .A3(\_zzLB[3][306] ), .Z(odata[274]));
Q_MX04 U3967 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][307] ), .A1(\_zzLB[1][307] ), .A2(\_zzLB[2][307] ), .A3(\_zzLB[3][307] ), .Z(odata[275]));
Q_MX04 U3968 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][308] ), .A1(\_zzLB[1][308] ), .A2(\_zzLB[2][308] ), .A3(\_zzLB[3][308] ), .Z(odata[276]));
Q_MX04 U3969 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][309] ), .A1(\_zzLB[1][309] ), .A2(\_zzLB[2][309] ), .A3(\_zzLB[3][309] ), .Z(odata[277]));
Q_MX04 U3970 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][310] ), .A1(\_zzLB[1][310] ), .A2(\_zzLB[2][310] ), .A3(\_zzLB[3][310] ), .Z(odata[278]));
Q_MX04 U3971 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][311] ), .A1(\_zzLB[1][311] ), .A2(\_zzLB[2][311] ), .A3(\_zzLB[3][311] ), .Z(odata[279]));
Q_MX04 U3972 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][312] ), .A1(\_zzLB[1][312] ), .A2(\_zzLB[2][312] ), .A3(\_zzLB[3][312] ), .Z(odata[280]));
Q_MX04 U3973 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][313] ), .A1(\_zzLB[1][313] ), .A2(\_zzLB[2][313] ), .A3(\_zzLB[3][313] ), .Z(odata[281]));
Q_MX04 U3974 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][314] ), .A1(\_zzLB[1][314] ), .A2(\_zzLB[2][314] ), .A3(\_zzLB[3][314] ), .Z(odata[282]));
Q_MX04 U3975 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][315] ), .A1(\_zzLB[1][315] ), .A2(\_zzLB[2][315] ), .A3(\_zzLB[3][315] ), .Z(odata[283]));
Q_MX04 U3976 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][316] ), .A1(\_zzLB[1][316] ), .A2(\_zzLB[2][316] ), .A3(\_zzLB[3][316] ), .Z(odata[284]));
Q_MX04 U3977 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][317] ), .A1(\_zzLB[1][317] ), .A2(\_zzLB[2][317] ), .A3(\_zzLB[3][317] ), .Z(odata[285]));
Q_MX04 U3978 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][318] ), .A1(\_zzLB[1][318] ), .A2(\_zzLB[2][318] ), .A3(\_zzLB[3][318] ), .Z(odata[286]));
Q_MX04 U3979 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][319] ), .A1(\_zzLB[1][319] ), .A2(\_zzLB[2][319] ), .A3(\_zzLB[3][319] ), .Z(odata[287]));
Q_MX04 U3980 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][320] ), .A1(\_zzLB[1][320] ), .A2(\_zzLB[2][320] ), .A3(\_zzLB[3][320] ), .Z(odata[288]));
Q_MX04 U3981 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][321] ), .A1(\_zzLB[1][321] ), .A2(\_zzLB[2][321] ), .A3(\_zzLB[3][321] ), .Z(odata[289]));
Q_MX04 U3982 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][322] ), .A1(\_zzLB[1][322] ), .A2(\_zzLB[2][322] ), .A3(\_zzLB[3][322] ), .Z(odata[290]));
Q_MX04 U3983 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][323] ), .A1(\_zzLB[1][323] ), .A2(\_zzLB[2][323] ), .A3(\_zzLB[3][323] ), .Z(odata[291]));
Q_MX04 U3984 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][324] ), .A1(\_zzLB[1][324] ), .A2(\_zzLB[2][324] ), .A3(\_zzLB[3][324] ), .Z(odata[292]));
Q_MX04 U3985 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][325] ), .A1(\_zzLB[1][325] ), .A2(\_zzLB[2][325] ), .A3(\_zzLB[3][325] ), .Z(odata[293]));
Q_MX04 U3986 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][326] ), .A1(\_zzLB[1][326] ), .A2(\_zzLB[2][326] ), .A3(\_zzLB[3][326] ), .Z(odata[294]));
Q_MX04 U3987 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][327] ), .A1(\_zzLB[1][327] ), .A2(\_zzLB[2][327] ), .A3(\_zzLB[3][327] ), .Z(odata[295]));
Q_MX04 U3988 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][328] ), .A1(\_zzLB[1][328] ), .A2(\_zzLB[2][328] ), .A3(\_zzLB[3][328] ), .Z(odata[296]));
Q_MX04 U3989 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][329] ), .A1(\_zzLB[1][329] ), .A2(\_zzLB[2][329] ), .A3(\_zzLB[3][329] ), .Z(odata[297]));
Q_MX04 U3990 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][330] ), .A1(\_zzLB[1][330] ), .A2(\_zzLB[2][330] ), .A3(\_zzLB[3][330] ), .Z(odata[298]));
Q_MX04 U3991 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][331] ), .A1(\_zzLB[1][331] ), .A2(\_zzLB[2][331] ), .A3(\_zzLB[3][331] ), .Z(odata[299]));
Q_MX04 U3992 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][332] ), .A1(\_zzLB[1][332] ), .A2(\_zzLB[2][332] ), .A3(\_zzLB[3][332] ), .Z(odata[300]));
Q_MX04 U3993 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][333] ), .A1(\_zzLB[1][333] ), .A2(\_zzLB[2][333] ), .A3(\_zzLB[3][333] ), .Z(odata[301]));
Q_MX04 U3994 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][334] ), .A1(\_zzLB[1][334] ), .A2(\_zzLB[2][334] ), .A3(\_zzLB[3][334] ), .Z(odata[302]));
Q_MX04 U3995 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][335] ), .A1(\_zzLB[1][335] ), .A2(\_zzLB[2][335] ), .A3(\_zzLB[3][335] ), .Z(odata[303]));
Q_MX04 U3996 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][336] ), .A1(\_zzLB[1][336] ), .A2(\_zzLB[2][336] ), .A3(\_zzLB[3][336] ), .Z(odata[304]));
Q_MX04 U3997 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][337] ), .A1(\_zzLB[1][337] ), .A2(\_zzLB[2][337] ), .A3(\_zzLB[3][337] ), .Z(odata[305]));
Q_MX04 U3998 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][338] ), .A1(\_zzLB[1][338] ), .A2(\_zzLB[2][338] ), .A3(\_zzLB[3][338] ), .Z(odata[306]));
Q_MX04 U3999 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][339] ), .A1(\_zzLB[1][339] ), .A2(\_zzLB[2][339] ), .A3(\_zzLB[3][339] ), .Z(odata[307]));
Q_MX04 U4000 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][340] ), .A1(\_zzLB[1][340] ), .A2(\_zzLB[2][340] ), .A3(\_zzLB[3][340] ), .Z(odata[308]));
Q_MX04 U4001 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][341] ), .A1(\_zzLB[1][341] ), .A2(\_zzLB[2][341] ), .A3(\_zzLB[3][341] ), .Z(odata[309]));
Q_MX04 U4002 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][342] ), .A1(\_zzLB[1][342] ), .A2(\_zzLB[2][342] ), .A3(\_zzLB[3][342] ), .Z(odata[310]));
Q_MX04 U4003 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][343] ), .A1(\_zzLB[1][343] ), .A2(\_zzLB[2][343] ), .A3(\_zzLB[3][343] ), .Z(odata[311]));
Q_MX04 U4004 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][344] ), .A1(\_zzLB[1][344] ), .A2(\_zzLB[2][344] ), .A3(\_zzLB[3][344] ), .Z(odata[312]));
Q_MX04 U4005 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][345] ), .A1(\_zzLB[1][345] ), .A2(\_zzLB[2][345] ), .A3(\_zzLB[3][345] ), .Z(odata[313]));
Q_MX04 U4006 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][346] ), .A1(\_zzLB[1][346] ), .A2(\_zzLB[2][346] ), .A3(\_zzLB[3][346] ), .Z(odata[314]));
Q_MX04 U4007 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][347] ), .A1(\_zzLB[1][347] ), .A2(\_zzLB[2][347] ), .A3(\_zzLB[3][347] ), .Z(odata[315]));
Q_MX04 U4008 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][348] ), .A1(\_zzLB[1][348] ), .A2(\_zzLB[2][348] ), .A3(\_zzLB[3][348] ), .Z(odata[316]));
Q_MX04 U4009 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][349] ), .A1(\_zzLB[1][349] ), .A2(\_zzLB[2][349] ), .A3(\_zzLB[3][349] ), .Z(odata[317]));
Q_MX04 U4010 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][350] ), .A1(\_zzLB[1][350] ), .A2(\_zzLB[2][350] ), .A3(\_zzLB[3][350] ), .Z(odata[318]));
Q_MX04 U4011 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][351] ), .A1(\_zzLB[1][351] ), .A2(\_zzLB[2][351] ), .A3(\_zzLB[3][351] ), .Z(odata[319]));
Q_MX04 U4012 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][352] ), .A1(\_zzLB[1][352] ), .A2(\_zzLB[2][352] ), .A3(\_zzLB[3][352] ), .Z(odata[320]));
Q_MX04 U4013 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][353] ), .A1(\_zzLB[1][353] ), .A2(\_zzLB[2][353] ), .A3(\_zzLB[3][353] ), .Z(odata[321]));
Q_MX04 U4014 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][354] ), .A1(\_zzLB[1][354] ), .A2(\_zzLB[2][354] ), .A3(\_zzLB[3][354] ), .Z(odata[322]));
Q_MX04 U4015 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][355] ), .A1(\_zzLB[1][355] ), .A2(\_zzLB[2][355] ), .A3(\_zzLB[3][355] ), .Z(odata[323]));
Q_MX04 U4016 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][356] ), .A1(\_zzLB[1][356] ), .A2(\_zzLB[2][356] ), .A3(\_zzLB[3][356] ), .Z(odata[324]));
Q_MX04 U4017 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][357] ), .A1(\_zzLB[1][357] ), .A2(\_zzLB[2][357] ), .A3(\_zzLB[3][357] ), .Z(odata[325]));
Q_MX04 U4018 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][358] ), .A1(\_zzLB[1][358] ), .A2(\_zzLB[2][358] ), .A3(\_zzLB[3][358] ), .Z(odata[326]));
Q_MX04 U4019 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][359] ), .A1(\_zzLB[1][359] ), .A2(\_zzLB[2][359] ), .A3(\_zzLB[3][359] ), .Z(odata[327]));
Q_MX04 U4020 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][360] ), .A1(\_zzLB[1][360] ), .A2(\_zzLB[2][360] ), .A3(\_zzLB[3][360] ), .Z(odata[328]));
Q_MX04 U4021 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][361] ), .A1(\_zzLB[1][361] ), .A2(\_zzLB[2][361] ), .A3(\_zzLB[3][361] ), .Z(odata[329]));
Q_MX04 U4022 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][362] ), .A1(\_zzLB[1][362] ), .A2(\_zzLB[2][362] ), .A3(\_zzLB[3][362] ), .Z(odata[330]));
Q_MX04 U4023 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][363] ), .A1(\_zzLB[1][363] ), .A2(\_zzLB[2][363] ), .A3(\_zzLB[3][363] ), .Z(odata[331]));
Q_MX04 U4024 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][364] ), .A1(\_zzLB[1][364] ), .A2(\_zzLB[2][364] ), .A3(\_zzLB[3][364] ), .Z(odata[332]));
Q_MX04 U4025 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][365] ), .A1(\_zzLB[1][365] ), .A2(\_zzLB[2][365] ), .A3(\_zzLB[3][365] ), .Z(odata[333]));
Q_MX04 U4026 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][366] ), .A1(\_zzLB[1][366] ), .A2(\_zzLB[2][366] ), .A3(\_zzLB[3][366] ), .Z(odata[334]));
Q_MX04 U4027 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][367] ), .A1(\_zzLB[1][367] ), .A2(\_zzLB[2][367] ), .A3(\_zzLB[3][367] ), .Z(odata[335]));
Q_MX04 U4028 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][368] ), .A1(\_zzLB[1][368] ), .A2(\_zzLB[2][368] ), .A3(\_zzLB[3][368] ), .Z(odata[336]));
Q_MX04 U4029 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][369] ), .A1(\_zzLB[1][369] ), .A2(\_zzLB[2][369] ), .A3(\_zzLB[3][369] ), .Z(odata[337]));
Q_MX04 U4030 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][370] ), .A1(\_zzLB[1][370] ), .A2(\_zzLB[2][370] ), .A3(\_zzLB[3][370] ), .Z(odata[338]));
Q_MX04 U4031 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][371] ), .A1(\_zzLB[1][371] ), .A2(\_zzLB[2][371] ), .A3(\_zzLB[3][371] ), .Z(odata[339]));
Q_MX04 U4032 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][372] ), .A1(\_zzLB[1][372] ), .A2(\_zzLB[2][372] ), .A3(\_zzLB[3][372] ), .Z(odata[340]));
Q_MX04 U4033 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][373] ), .A1(\_zzLB[1][373] ), .A2(\_zzLB[2][373] ), .A3(\_zzLB[3][373] ), .Z(odata[341]));
Q_MX04 U4034 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][374] ), .A1(\_zzLB[1][374] ), .A2(\_zzLB[2][374] ), .A3(\_zzLB[3][374] ), .Z(odata[342]));
Q_MX04 U4035 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][375] ), .A1(\_zzLB[1][375] ), .A2(\_zzLB[2][375] ), .A3(\_zzLB[3][375] ), .Z(odata[343]));
Q_MX04 U4036 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][376] ), .A1(\_zzLB[1][376] ), .A2(\_zzLB[2][376] ), .A3(\_zzLB[3][376] ), .Z(odata[344]));
Q_MX04 U4037 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][377] ), .A1(\_zzLB[1][377] ), .A2(\_zzLB[2][377] ), .A3(\_zzLB[3][377] ), .Z(odata[345]));
Q_MX04 U4038 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][378] ), .A1(\_zzLB[1][378] ), .A2(\_zzLB[2][378] ), .A3(\_zzLB[3][378] ), .Z(odata[346]));
Q_MX04 U4039 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][379] ), .A1(\_zzLB[1][379] ), .A2(\_zzLB[2][379] ), .A3(\_zzLB[3][379] ), .Z(odata[347]));
Q_MX04 U4040 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][380] ), .A1(\_zzLB[1][380] ), .A2(\_zzLB[2][380] ), .A3(\_zzLB[3][380] ), .Z(odata[348]));
Q_MX04 U4041 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][381] ), .A1(\_zzLB[1][381] ), .A2(\_zzLB[2][381] ), .A3(\_zzLB[3][381] ), .Z(odata[349]));
Q_MX04 U4042 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][382] ), .A1(\_zzLB[1][382] ), .A2(\_zzLB[2][382] ), .A3(\_zzLB[3][382] ), .Z(odata[350]));
Q_MX04 U4043 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][383] ), .A1(\_zzLB[1][383] ), .A2(\_zzLB[2][383] ), .A3(\_zzLB[3][383] ), .Z(odata[351]));
Q_MX04 U4044 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][384] ), .A1(\_zzLB[1][384] ), .A2(\_zzLB[2][384] ), .A3(\_zzLB[3][384] ), .Z(odata[352]));
Q_MX04 U4045 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][385] ), .A1(\_zzLB[1][385] ), .A2(\_zzLB[2][385] ), .A3(\_zzLB[3][385] ), .Z(odata[353]));
Q_MX04 U4046 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][386] ), .A1(\_zzLB[1][386] ), .A2(\_zzLB[2][386] ), .A3(\_zzLB[3][386] ), .Z(odata[354]));
Q_MX04 U4047 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][387] ), .A1(\_zzLB[1][387] ), .A2(\_zzLB[2][387] ), .A3(\_zzLB[3][387] ), .Z(odata[355]));
Q_MX04 U4048 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][388] ), .A1(\_zzLB[1][388] ), .A2(\_zzLB[2][388] ), .A3(\_zzLB[3][388] ), .Z(odata[356]));
Q_MX04 U4049 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][389] ), .A1(\_zzLB[1][389] ), .A2(\_zzLB[2][389] ), .A3(\_zzLB[3][389] ), .Z(odata[357]));
Q_MX04 U4050 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][390] ), .A1(\_zzLB[1][390] ), .A2(\_zzLB[2][390] ), .A3(\_zzLB[3][390] ), .Z(odata[358]));
Q_MX04 U4051 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][391] ), .A1(\_zzLB[1][391] ), .A2(\_zzLB[2][391] ), .A3(\_zzLB[3][391] ), .Z(odata[359]));
Q_MX04 U4052 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][392] ), .A1(\_zzLB[1][392] ), .A2(\_zzLB[2][392] ), .A3(\_zzLB[3][392] ), .Z(odata[360]));
Q_MX04 U4053 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][393] ), .A1(\_zzLB[1][393] ), .A2(\_zzLB[2][393] ), .A3(\_zzLB[3][393] ), .Z(odata[361]));
Q_MX04 U4054 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][394] ), .A1(\_zzLB[1][394] ), .A2(\_zzLB[2][394] ), .A3(\_zzLB[3][394] ), .Z(odata[362]));
Q_MX04 U4055 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][395] ), .A1(\_zzLB[1][395] ), .A2(\_zzLB[2][395] ), .A3(\_zzLB[3][395] ), .Z(odata[363]));
Q_MX04 U4056 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][396] ), .A1(\_zzLB[1][396] ), .A2(\_zzLB[2][396] ), .A3(\_zzLB[3][396] ), .Z(odata[364]));
Q_MX04 U4057 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][397] ), .A1(\_zzLB[1][397] ), .A2(\_zzLB[2][397] ), .A3(\_zzLB[3][397] ), .Z(odata[365]));
Q_MX04 U4058 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][398] ), .A1(\_zzLB[1][398] ), .A2(\_zzLB[2][398] ), .A3(\_zzLB[3][398] ), .Z(odata[366]));
Q_MX04 U4059 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][399] ), .A1(\_zzLB[1][399] ), .A2(\_zzLB[2][399] ), .A3(\_zzLB[3][399] ), .Z(odata[367]));
Q_MX04 U4060 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][400] ), .A1(\_zzLB[1][400] ), .A2(\_zzLB[2][400] ), .A3(\_zzLB[3][400] ), .Z(odata[368]));
Q_MX04 U4061 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][401] ), .A1(\_zzLB[1][401] ), .A2(\_zzLB[2][401] ), .A3(\_zzLB[3][401] ), .Z(odata[369]));
Q_MX04 U4062 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][402] ), .A1(\_zzLB[1][402] ), .A2(\_zzLB[2][402] ), .A3(\_zzLB[3][402] ), .Z(odata[370]));
Q_MX04 U4063 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][403] ), .A1(\_zzLB[1][403] ), .A2(\_zzLB[2][403] ), .A3(\_zzLB[3][403] ), .Z(odata[371]));
Q_MX04 U4064 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][404] ), .A1(\_zzLB[1][404] ), .A2(\_zzLB[2][404] ), .A3(\_zzLB[3][404] ), .Z(odata[372]));
Q_MX04 U4065 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][405] ), .A1(\_zzLB[1][405] ), .A2(\_zzLB[2][405] ), .A3(\_zzLB[3][405] ), .Z(odata[373]));
Q_MX04 U4066 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][406] ), .A1(\_zzLB[1][406] ), .A2(\_zzLB[2][406] ), .A3(\_zzLB[3][406] ), .Z(odata[374]));
Q_MX04 U4067 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][407] ), .A1(\_zzLB[1][407] ), .A2(\_zzLB[2][407] ), .A3(\_zzLB[3][407] ), .Z(odata[375]));
Q_MX04 U4068 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][408] ), .A1(\_zzLB[1][408] ), .A2(\_zzLB[2][408] ), .A3(\_zzLB[3][408] ), .Z(odata[376]));
Q_MX04 U4069 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][409] ), .A1(\_zzLB[1][409] ), .A2(\_zzLB[2][409] ), .A3(\_zzLB[3][409] ), .Z(odata[377]));
Q_MX04 U4070 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][410] ), .A1(\_zzLB[1][410] ), .A2(\_zzLB[2][410] ), .A3(\_zzLB[3][410] ), .Z(odata[378]));
Q_MX04 U4071 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][411] ), .A1(\_zzLB[1][411] ), .A2(\_zzLB[2][411] ), .A3(\_zzLB[3][411] ), .Z(odata[379]));
Q_MX04 U4072 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][412] ), .A1(\_zzLB[1][412] ), .A2(\_zzLB[2][412] ), .A3(\_zzLB[3][412] ), .Z(odata[380]));
Q_MX04 U4073 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][413] ), .A1(\_zzLB[1][413] ), .A2(\_zzLB[2][413] ), .A3(\_zzLB[3][413] ), .Z(odata[381]));
Q_MX04 U4074 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][414] ), .A1(\_zzLB[1][414] ), .A2(\_zzLB[2][414] ), .A3(\_zzLB[3][414] ), .Z(odata[382]));
Q_MX04 U4075 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][415] ), .A1(\_zzLB[1][415] ), .A2(\_zzLB[2][415] ), .A3(\_zzLB[3][415] ), .Z(odata[383]));
Q_MX04 U4076 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][416] ), .A1(\_zzLB[1][416] ), .A2(\_zzLB[2][416] ), .A3(\_zzLB[3][416] ), .Z(odata[384]));
Q_MX04 U4077 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][417] ), .A1(\_zzLB[1][417] ), .A2(\_zzLB[2][417] ), .A3(\_zzLB[3][417] ), .Z(odata[385]));
Q_MX04 U4078 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][418] ), .A1(\_zzLB[1][418] ), .A2(\_zzLB[2][418] ), .A3(\_zzLB[3][418] ), .Z(odata[386]));
Q_MX04 U4079 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][419] ), .A1(\_zzLB[1][419] ), .A2(\_zzLB[2][419] ), .A3(\_zzLB[3][419] ), .Z(odata[387]));
Q_MX04 U4080 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][420] ), .A1(\_zzLB[1][420] ), .A2(\_zzLB[2][420] ), .A3(\_zzLB[3][420] ), .Z(odata[388]));
Q_MX04 U4081 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][421] ), .A1(\_zzLB[1][421] ), .A2(\_zzLB[2][421] ), .A3(\_zzLB[3][421] ), .Z(odata[389]));
Q_MX04 U4082 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][422] ), .A1(\_zzLB[1][422] ), .A2(\_zzLB[2][422] ), .A3(\_zzLB[3][422] ), .Z(odata[390]));
Q_MX04 U4083 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][423] ), .A1(\_zzLB[1][423] ), .A2(\_zzLB[2][423] ), .A3(\_zzLB[3][423] ), .Z(odata[391]));
Q_MX04 U4084 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][424] ), .A1(\_zzLB[1][424] ), .A2(\_zzLB[2][424] ), .A3(\_zzLB[3][424] ), .Z(odata[392]));
Q_MX04 U4085 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][425] ), .A1(\_zzLB[1][425] ), .A2(\_zzLB[2][425] ), .A3(\_zzLB[3][425] ), .Z(odata[393]));
Q_MX04 U4086 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][426] ), .A1(\_zzLB[1][426] ), .A2(\_zzLB[2][426] ), .A3(\_zzLB[3][426] ), .Z(odata[394]));
Q_MX04 U4087 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][427] ), .A1(\_zzLB[1][427] ), .A2(\_zzLB[2][427] ), .A3(\_zzLB[3][427] ), .Z(odata[395]));
Q_MX04 U4088 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][428] ), .A1(\_zzLB[1][428] ), .A2(\_zzLB[2][428] ), .A3(\_zzLB[3][428] ), .Z(odata[396]));
Q_MX04 U4089 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][429] ), .A1(\_zzLB[1][429] ), .A2(\_zzLB[2][429] ), .A3(\_zzLB[3][429] ), .Z(odata[397]));
Q_MX04 U4090 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][430] ), .A1(\_zzLB[1][430] ), .A2(\_zzLB[2][430] ), .A3(\_zzLB[3][430] ), .Z(odata[398]));
Q_MX04 U4091 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][431] ), .A1(\_zzLB[1][431] ), .A2(\_zzLB[2][431] ), .A3(\_zzLB[3][431] ), .Z(odata[399]));
Q_MX04 U4092 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][432] ), .A1(\_zzLB[1][432] ), .A2(\_zzLB[2][432] ), .A3(\_zzLB[3][432] ), .Z(odata[400]));
Q_MX04 U4093 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][433] ), .A1(\_zzLB[1][433] ), .A2(\_zzLB[2][433] ), .A3(\_zzLB[3][433] ), .Z(odata[401]));
Q_MX04 U4094 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][434] ), .A1(\_zzLB[1][434] ), .A2(\_zzLB[2][434] ), .A3(\_zzLB[3][434] ), .Z(odata[402]));
Q_MX04 U4095 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][435] ), .A1(\_zzLB[1][435] ), .A2(\_zzLB[2][435] ), .A3(\_zzLB[3][435] ), .Z(odata[403]));
Q_MX04 U4096 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][436] ), .A1(\_zzLB[1][436] ), .A2(\_zzLB[2][436] ), .A3(\_zzLB[3][436] ), .Z(odata[404]));
Q_MX04 U4097 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][437] ), .A1(\_zzLB[1][437] ), .A2(\_zzLB[2][437] ), .A3(\_zzLB[3][437] ), .Z(odata[405]));
Q_MX04 U4098 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][438] ), .A1(\_zzLB[1][438] ), .A2(\_zzLB[2][438] ), .A3(\_zzLB[3][438] ), .Z(odata[406]));
Q_MX04 U4099 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][439] ), .A1(\_zzLB[1][439] ), .A2(\_zzLB[2][439] ), .A3(\_zzLB[3][439] ), .Z(odata[407]));
Q_MX04 U4100 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][440] ), .A1(\_zzLB[1][440] ), .A2(\_zzLB[2][440] ), .A3(\_zzLB[3][440] ), .Z(odata[408]));
Q_MX04 U4101 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][441] ), .A1(\_zzLB[1][441] ), .A2(\_zzLB[2][441] ), .A3(\_zzLB[3][441] ), .Z(odata[409]));
Q_MX04 U4102 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][442] ), .A1(\_zzLB[1][442] ), .A2(\_zzLB[2][442] ), .A3(\_zzLB[3][442] ), .Z(odata[410]));
Q_MX04 U4103 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][443] ), .A1(\_zzLB[1][443] ), .A2(\_zzLB[2][443] ), .A3(\_zzLB[3][443] ), .Z(odata[411]));
Q_MX04 U4104 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][444] ), .A1(\_zzLB[1][444] ), .A2(\_zzLB[2][444] ), .A3(\_zzLB[3][444] ), .Z(odata[412]));
Q_MX04 U4105 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][445] ), .A1(\_zzLB[1][445] ), .A2(\_zzLB[2][445] ), .A3(\_zzLB[3][445] ), .Z(odata[413]));
Q_MX04 U4106 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][446] ), .A1(\_zzLB[1][446] ), .A2(\_zzLB[2][446] ), .A3(\_zzLB[3][446] ), .Z(odata[414]));
Q_MX04 U4107 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][447] ), .A1(\_zzLB[1][447] ), .A2(\_zzLB[2][447] ), .A3(\_zzLB[3][447] ), .Z(odata[415]));
Q_MX04 U4108 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][448] ), .A1(\_zzLB[1][448] ), .A2(\_zzLB[2][448] ), .A3(\_zzLB[3][448] ), .Z(odata[416]));
Q_MX04 U4109 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][449] ), .A1(\_zzLB[1][449] ), .A2(\_zzLB[2][449] ), .A3(\_zzLB[3][449] ), .Z(odata[417]));
Q_MX04 U4110 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][450] ), .A1(\_zzLB[1][450] ), .A2(\_zzLB[2][450] ), .A3(\_zzLB[3][450] ), .Z(odata[418]));
Q_MX04 U4111 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][451] ), .A1(\_zzLB[1][451] ), .A2(\_zzLB[2][451] ), .A3(\_zzLB[3][451] ), .Z(odata[419]));
Q_MX04 U4112 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][452] ), .A1(\_zzLB[1][452] ), .A2(\_zzLB[2][452] ), .A3(\_zzLB[3][452] ), .Z(odata[420]));
Q_MX04 U4113 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][453] ), .A1(\_zzLB[1][453] ), .A2(\_zzLB[2][453] ), .A3(\_zzLB[3][453] ), .Z(odata[421]));
Q_MX04 U4114 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][454] ), .A1(\_zzLB[1][454] ), .A2(\_zzLB[2][454] ), .A3(\_zzLB[3][454] ), .Z(odata[422]));
Q_MX04 U4115 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][455] ), .A1(\_zzLB[1][455] ), .A2(\_zzLB[2][455] ), .A3(\_zzLB[3][455] ), .Z(odata[423]));
Q_MX04 U4116 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][456] ), .A1(\_zzLB[1][456] ), .A2(\_zzLB[2][456] ), .A3(\_zzLB[3][456] ), .Z(odata[424]));
Q_MX04 U4117 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][457] ), .A1(\_zzLB[1][457] ), .A2(\_zzLB[2][457] ), .A3(\_zzLB[3][457] ), .Z(odata[425]));
Q_MX04 U4118 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][458] ), .A1(\_zzLB[1][458] ), .A2(\_zzLB[2][458] ), .A3(\_zzLB[3][458] ), .Z(odata[426]));
Q_MX04 U4119 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][459] ), .A1(\_zzLB[1][459] ), .A2(\_zzLB[2][459] ), .A3(\_zzLB[3][459] ), .Z(odata[427]));
Q_MX04 U4120 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][460] ), .A1(\_zzLB[1][460] ), .A2(\_zzLB[2][460] ), .A3(\_zzLB[3][460] ), .Z(odata[428]));
Q_MX04 U4121 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][461] ), .A1(\_zzLB[1][461] ), .A2(\_zzLB[2][461] ), .A3(\_zzLB[3][461] ), .Z(odata[429]));
Q_MX04 U4122 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][462] ), .A1(\_zzLB[1][462] ), .A2(\_zzLB[2][462] ), .A3(\_zzLB[3][462] ), .Z(odata[430]));
Q_MX04 U4123 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][463] ), .A1(\_zzLB[1][463] ), .A2(\_zzLB[2][463] ), .A3(\_zzLB[3][463] ), .Z(odata[431]));
Q_MX04 U4124 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][464] ), .A1(\_zzLB[1][464] ), .A2(\_zzLB[2][464] ), .A3(\_zzLB[3][464] ), .Z(odata[432]));
Q_MX04 U4125 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][465] ), .A1(\_zzLB[1][465] ), .A2(\_zzLB[2][465] ), .A3(\_zzLB[3][465] ), .Z(odata[433]));
Q_MX04 U4126 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][466] ), .A1(\_zzLB[1][466] ), .A2(\_zzLB[2][466] ), .A3(\_zzLB[3][466] ), .Z(odata[434]));
Q_MX04 U4127 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][467] ), .A1(\_zzLB[1][467] ), .A2(\_zzLB[2][467] ), .A3(\_zzLB[3][467] ), .Z(odata[435]));
Q_MX04 U4128 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][468] ), .A1(\_zzLB[1][468] ), .A2(\_zzLB[2][468] ), .A3(\_zzLB[3][468] ), .Z(odata[436]));
Q_MX04 U4129 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][469] ), .A1(\_zzLB[1][469] ), .A2(\_zzLB[2][469] ), .A3(\_zzLB[3][469] ), .Z(odata[437]));
Q_MX04 U4130 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][470] ), .A1(\_zzLB[1][470] ), .A2(\_zzLB[2][470] ), .A3(\_zzLB[3][470] ), .Z(odata[438]));
Q_MX04 U4131 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][471] ), .A1(\_zzLB[1][471] ), .A2(\_zzLB[2][471] ), .A3(\_zzLB[3][471] ), .Z(odata[439]));
Q_MX04 U4132 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][472] ), .A1(\_zzLB[1][472] ), .A2(\_zzLB[2][472] ), .A3(\_zzLB[3][472] ), .Z(odata[440]));
Q_MX04 U4133 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][473] ), .A1(\_zzLB[1][473] ), .A2(\_zzLB[2][473] ), .A3(\_zzLB[3][473] ), .Z(odata[441]));
Q_MX04 U4134 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][474] ), .A1(\_zzLB[1][474] ), .A2(\_zzLB[2][474] ), .A3(\_zzLB[3][474] ), .Z(odata[442]));
Q_MX04 U4135 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][475] ), .A1(\_zzLB[1][475] ), .A2(\_zzLB[2][475] ), .A3(\_zzLB[3][475] ), .Z(odata[443]));
Q_MX04 U4136 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][476] ), .A1(\_zzLB[1][476] ), .A2(\_zzLB[2][476] ), .A3(\_zzLB[3][476] ), .Z(odata[444]));
Q_MX04 U4137 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][477] ), .A1(\_zzLB[1][477] ), .A2(\_zzLB[2][477] ), .A3(\_zzLB[3][477] ), .Z(odata[445]));
Q_MX04 U4138 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][478] ), .A1(\_zzLB[1][478] ), .A2(\_zzLB[2][478] ), .A3(\_zzLB[3][478] ), .Z(odata[446]));
Q_MX04 U4139 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][479] ), .A1(\_zzLB[1][479] ), .A2(\_zzLB[2][479] ), .A3(\_zzLB[3][479] ), .Z(odata[447]));
Q_MX04 U4140 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][480] ), .A1(\_zzLB[1][480] ), .A2(\_zzLB[2][480] ), .A3(\_zzLB[3][480] ), .Z(odata[448]));
Q_MX04 U4141 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][481] ), .A1(\_zzLB[1][481] ), .A2(\_zzLB[2][481] ), .A3(\_zzLB[3][481] ), .Z(odata[449]));
Q_MX04 U4142 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][482] ), .A1(\_zzLB[1][482] ), .A2(\_zzLB[2][482] ), .A3(\_zzLB[3][482] ), .Z(odata[450]));
Q_MX04 U4143 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][483] ), .A1(\_zzLB[1][483] ), .A2(\_zzLB[2][483] ), .A3(\_zzLB[3][483] ), .Z(odata[451]));
Q_MX04 U4144 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][484] ), .A1(\_zzLB[1][484] ), .A2(\_zzLB[2][484] ), .A3(\_zzLB[3][484] ), .Z(odata[452]));
Q_MX04 U4145 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][485] ), .A1(\_zzLB[1][485] ), .A2(\_zzLB[2][485] ), .A3(\_zzLB[3][485] ), .Z(odata[453]));
Q_MX04 U4146 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][486] ), .A1(\_zzLB[1][486] ), .A2(\_zzLB[2][486] ), .A3(\_zzLB[3][486] ), .Z(odata[454]));
Q_MX04 U4147 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][487] ), .A1(\_zzLB[1][487] ), .A2(\_zzLB[2][487] ), .A3(\_zzLB[3][487] ), .Z(odata[455]));
Q_MX04 U4148 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][488] ), .A1(\_zzLB[1][488] ), .A2(\_zzLB[2][488] ), .A3(\_zzLB[3][488] ), .Z(odata[456]));
Q_MX04 U4149 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][489] ), .A1(\_zzLB[1][489] ), .A2(\_zzLB[2][489] ), .A3(\_zzLB[3][489] ), .Z(odata[457]));
Q_MX04 U4150 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][490] ), .A1(\_zzLB[1][490] ), .A2(\_zzLB[2][490] ), .A3(\_zzLB[3][490] ), .Z(odata[458]));
Q_MX04 U4151 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][491] ), .A1(\_zzLB[1][491] ), .A2(\_zzLB[2][491] ), .A3(\_zzLB[3][491] ), .Z(odata[459]));
Q_MX04 U4152 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][492] ), .A1(\_zzLB[1][492] ), .A2(\_zzLB[2][492] ), .A3(\_zzLB[3][492] ), .Z(odata[460]));
Q_MX04 U4153 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][493] ), .A1(\_zzLB[1][493] ), .A2(\_zzLB[2][493] ), .A3(\_zzLB[3][493] ), .Z(odata[461]));
Q_MX04 U4154 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][494] ), .A1(\_zzLB[1][494] ), .A2(\_zzLB[2][494] ), .A3(\_zzLB[3][494] ), .Z(odata[462]));
Q_MX04 U4155 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][495] ), .A1(\_zzLB[1][495] ), .A2(\_zzLB[2][495] ), .A3(\_zzLB[3][495] ), .Z(odata[463]));
Q_MX04 U4156 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][496] ), .A1(\_zzLB[1][496] ), .A2(\_zzLB[2][496] ), .A3(\_zzLB[3][496] ), .Z(odata[464]));
Q_MX04 U4157 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][497] ), .A1(\_zzLB[1][497] ), .A2(\_zzLB[2][497] ), .A3(\_zzLB[3][497] ), .Z(odata[465]));
Q_MX04 U4158 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][498] ), .A1(\_zzLB[1][498] ), .A2(\_zzLB[2][498] ), .A3(\_zzLB[3][498] ), .Z(odata[466]));
Q_MX04 U4159 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][499] ), .A1(\_zzLB[1][499] ), .A2(\_zzLB[2][499] ), .A3(\_zzLB[3][499] ), .Z(odata[467]));
Q_MX04 U4160 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][500] ), .A1(\_zzLB[1][500] ), .A2(\_zzLB[2][500] ), .A3(\_zzLB[3][500] ), .Z(odata[468]));
Q_MX04 U4161 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][501] ), .A1(\_zzLB[1][501] ), .A2(\_zzLB[2][501] ), .A3(\_zzLB[3][501] ), .Z(odata[469]));
Q_MX04 U4162 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][502] ), .A1(\_zzLB[1][502] ), .A2(\_zzLB[2][502] ), .A3(\_zzLB[3][502] ), .Z(odata[470]));
Q_MX04 U4163 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][503] ), .A1(\_zzLB[1][503] ), .A2(\_zzLB[2][503] ), .A3(\_zzLB[3][503] ), .Z(odata[471]));
Q_MX04 U4164 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][504] ), .A1(\_zzLB[1][504] ), .A2(\_zzLB[2][504] ), .A3(\_zzLB[3][504] ), .Z(odata[472]));
Q_MX04 U4165 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][505] ), .A1(\_zzLB[1][505] ), .A2(\_zzLB[2][505] ), .A3(\_zzLB[3][505] ), .Z(odata[473]));
Q_MX04 U4166 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][506] ), .A1(\_zzLB[1][506] ), .A2(\_zzLB[2][506] ), .A3(\_zzLB[3][506] ), .Z(odata[474]));
Q_MX04 U4167 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][507] ), .A1(\_zzLB[1][507] ), .A2(\_zzLB[2][507] ), .A3(\_zzLB[3][507] ), .Z(odata[475]));
Q_MX04 U4168 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][508] ), .A1(\_zzLB[1][508] ), .A2(\_zzLB[2][508] ), .A3(\_zzLB[3][508] ), .Z(odata[476]));
Q_MX04 U4169 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][509] ), .A1(\_zzLB[1][509] ), .A2(\_zzLB[2][509] ), .A3(\_zzLB[3][509] ), .Z(odata[477]));
Q_MX04 U4170 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][510] ), .A1(\_zzLB[1][510] ), .A2(\_zzLB[2][510] ), .A3(\_zzLB[3][510] ), .Z(odata[478]));
Q_MX04 U4171 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][511] ), .A1(\_zzLB[1][511] ), .A2(\_zzLB[2][511] ), .A3(\_zzLB[3][511] ), .Z(odata[479]));
Q_MX04 U4172 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][512] ), .A1(\_zzLB[1][512] ), .A2(\_zzLB[2][512] ), .A3(\_zzLB[3][512] ), .Z(odata[480]));
Q_MX04 U4173 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][513] ), .A1(\_zzLB[1][513] ), .A2(\_zzLB[2][513] ), .A3(\_zzLB[3][513] ), .Z(odata[481]));
Q_MX04 U4174 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][514] ), .A1(\_zzLB[1][514] ), .A2(\_zzLB[2][514] ), .A3(\_zzLB[3][514] ), .Z(odata[482]));
Q_MX04 U4175 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][515] ), .A1(\_zzLB[1][515] ), .A2(\_zzLB[2][515] ), .A3(\_zzLB[3][515] ), .Z(odata[483]));
Q_MX04 U4176 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][516] ), .A1(\_zzLB[1][516] ), .A2(\_zzLB[2][516] ), .A3(\_zzLB[3][516] ), .Z(odata[484]));
Q_MX04 U4177 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][517] ), .A1(\_zzLB[1][517] ), .A2(\_zzLB[2][517] ), .A3(\_zzLB[3][517] ), .Z(odata[485]));
Q_MX04 U4178 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][518] ), .A1(\_zzLB[1][518] ), .A2(\_zzLB[2][518] ), .A3(\_zzLB[3][518] ), .Z(odata[486]));
Q_MX04 U4179 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][519] ), .A1(\_zzLB[1][519] ), .A2(\_zzLB[2][519] ), .A3(\_zzLB[3][519] ), .Z(odata[487]));
Q_MX04 U4180 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][520] ), .A1(\_zzLB[1][520] ), .A2(\_zzLB[2][520] ), .A3(\_zzLB[3][520] ), .Z(odata[488]));
Q_MX04 U4181 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][521] ), .A1(\_zzLB[1][521] ), .A2(\_zzLB[2][521] ), .A3(\_zzLB[3][521] ), .Z(odata[489]));
Q_MX04 U4182 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][522] ), .A1(\_zzLB[1][522] ), .A2(\_zzLB[2][522] ), .A3(\_zzLB[3][522] ), .Z(odata[490]));
Q_MX04 U4183 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][523] ), .A1(\_zzLB[1][523] ), .A2(\_zzLB[2][523] ), .A3(\_zzLB[3][523] ), .Z(odata[491]));
Q_MX04 U4184 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][524] ), .A1(\_zzLB[1][524] ), .A2(\_zzLB[2][524] ), .A3(\_zzLB[3][524] ), .Z(odata[492]));
Q_MX04 U4185 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][525] ), .A1(\_zzLB[1][525] ), .A2(\_zzLB[2][525] ), .A3(\_zzLB[3][525] ), .Z(odata[493]));
Q_MX04 U4186 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][526] ), .A1(\_zzLB[1][526] ), .A2(\_zzLB[2][526] ), .A3(\_zzLB[3][526] ), .Z(odata[494]));
Q_MX04 U4187 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][527] ), .A1(\_zzLB[1][527] ), .A2(\_zzLB[2][527] ), .A3(\_zzLB[3][527] ), .Z(odata[495]));
Q_MX04 U4188 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][528] ), .A1(\_zzLB[1][528] ), .A2(\_zzLB[2][528] ), .A3(\_zzLB[3][528] ), .Z(odata[496]));
Q_MX04 U4189 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][529] ), .A1(\_zzLB[1][529] ), .A2(\_zzLB[2][529] ), .A3(\_zzLB[3][529] ), .Z(odata[497]));
Q_MX04 U4190 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][530] ), .A1(\_zzLB[1][530] ), .A2(\_zzLB[2][530] ), .A3(\_zzLB[3][530] ), .Z(odata[498]));
Q_MX04 U4191 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][531] ), .A1(\_zzLB[1][531] ), .A2(\_zzLB[2][531] ), .A3(\_zzLB[3][531] ), .Z(odata[499]));
Q_MX04 U4192 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][532] ), .A1(\_zzLB[1][532] ), .A2(\_zzLB[2][532] ), .A3(\_zzLB[3][532] ), .Z(odata[500]));
Q_MX04 U4193 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][533] ), .A1(\_zzLB[1][533] ), .A2(\_zzLB[2][533] ), .A3(\_zzLB[3][533] ), .Z(odata[501]));
Q_MX04 U4194 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][534] ), .A1(\_zzLB[1][534] ), .A2(\_zzLB[2][534] ), .A3(\_zzLB[3][534] ), .Z(odata[502]));
Q_MX04 U4195 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][535] ), .A1(\_zzLB[1][535] ), .A2(\_zzLB[2][535] ), .A3(\_zzLB[3][535] ), .Z(odata[503]));
Q_MX04 U4196 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][536] ), .A1(\_zzLB[1][536] ), .A2(\_zzLB[2][536] ), .A3(\_zzLB[3][536] ), .Z(odata[504]));
Q_MX04 U4197 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][537] ), .A1(\_zzLB[1][537] ), .A2(\_zzLB[2][537] ), .A3(\_zzLB[3][537] ), .Z(odata[505]));
Q_MX04 U4198 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][538] ), .A1(\_zzLB[1][538] ), .A2(\_zzLB[2][538] ), .A3(\_zzLB[3][538] ), .Z(odata[506]));
Q_MX04 U4199 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][539] ), .A1(\_zzLB[1][539] ), .A2(\_zzLB[2][539] ), .A3(\_zzLB[3][539] ), .Z(odata[507]));
Q_MX04 U4200 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][540] ), .A1(\_zzLB[1][540] ), .A2(\_zzLB[2][540] ), .A3(\_zzLB[3][540] ), .Z(odata[508]));
Q_MX04 U4201 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][541] ), .A1(\_zzLB[1][541] ), .A2(\_zzLB[2][541] ), .A3(\_zzLB[3][541] ), .Z(odata[509]));
Q_MX04 U4202 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][542] ), .A1(\_zzLB[1][542] ), .A2(\_zzLB[2][542] ), .A3(\_zzLB[3][542] ), .Z(odata[510]));
Q_MX04 U4203 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][543] ), .A1(\_zzLB[1][543] ), .A2(\_zzLB[2][543] ), .A3(\_zzLB[3][543] ), .Z(odata[511]));
Q_MX04 U4204 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][544] ), .A1(\_zzLB[1][544] ), .A2(\_zzLB[2][544] ), .A3(\_zzLB[3][544] ), .Z(odata[512]));
Q_MX04 U4205 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][545] ), .A1(\_zzLB[1][545] ), .A2(\_zzLB[2][545] ), .A3(\_zzLB[3][545] ), .Z(odata[513]));
Q_MX04 U4206 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][546] ), .A1(\_zzLB[1][546] ), .A2(\_zzLB[2][546] ), .A3(\_zzLB[3][546] ), .Z(odata[514]));
Q_MX04 U4207 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][547] ), .A1(\_zzLB[1][547] ), .A2(\_zzLB[2][547] ), .A3(\_zzLB[3][547] ), .Z(odata[515]));
Q_MX04 U4208 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][548] ), .A1(\_zzLB[1][548] ), .A2(\_zzLB[2][548] ), .A3(\_zzLB[3][548] ), .Z(odata[516]));
Q_MX04 U4209 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][549] ), .A1(\_zzLB[1][549] ), .A2(\_zzLB[2][549] ), .A3(\_zzLB[3][549] ), .Z(odata[517]));
Q_MX04 U4210 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][550] ), .A1(\_zzLB[1][550] ), .A2(\_zzLB[2][550] ), .A3(\_zzLB[3][550] ), .Z(odata[518]));
Q_MX04 U4211 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][551] ), .A1(\_zzLB[1][551] ), .A2(\_zzLB[2][551] ), .A3(\_zzLB[3][551] ), .Z(odata[519]));
Q_MX04 U4212 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][552] ), .A1(\_zzLB[1][552] ), .A2(\_zzLB[2][552] ), .A3(\_zzLB[3][552] ), .Z(odata[520]));
Q_MX04 U4213 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][553] ), .A1(\_zzLB[1][553] ), .A2(\_zzLB[2][553] ), .A3(\_zzLB[3][553] ), .Z(odata[521]));
Q_MX04 U4214 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][554] ), .A1(\_zzLB[1][554] ), .A2(\_zzLB[2][554] ), .A3(\_zzLB[3][554] ), .Z(odata[522]));
Q_MX04 U4215 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][555] ), .A1(\_zzLB[1][555] ), .A2(\_zzLB[2][555] ), .A3(\_zzLB[3][555] ), .Z(odata[523]));
Q_MX04 U4216 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][556] ), .A1(\_zzLB[1][556] ), .A2(\_zzLB[2][556] ), .A3(\_zzLB[3][556] ), .Z(odata[524]));
Q_MX04 U4217 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][557] ), .A1(\_zzLB[1][557] ), .A2(\_zzLB[2][557] ), .A3(\_zzLB[3][557] ), .Z(odata[525]));
Q_MX04 U4218 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][558] ), .A1(\_zzLB[1][558] ), .A2(\_zzLB[2][558] ), .A3(\_zzLB[3][558] ), .Z(odata[526]));
Q_MX04 U4219 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][559] ), .A1(\_zzLB[1][559] ), .A2(\_zzLB[2][559] ), .A3(\_zzLB[3][559] ), .Z(odata[527]));
Q_MX04 U4220 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][560] ), .A1(\_zzLB[1][560] ), .A2(\_zzLB[2][560] ), .A3(\_zzLB[3][560] ), .Z(odata[528]));
Q_MX04 U4221 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][561] ), .A1(\_zzLB[1][561] ), .A2(\_zzLB[2][561] ), .A3(\_zzLB[3][561] ), .Z(odata[529]));
Q_MX04 U4222 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][562] ), .A1(\_zzLB[1][562] ), .A2(\_zzLB[2][562] ), .A3(\_zzLB[3][562] ), .Z(odata[530]));
Q_MX04 U4223 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][563] ), .A1(\_zzLB[1][563] ), .A2(\_zzLB[2][563] ), .A3(\_zzLB[3][563] ), .Z(odata[531]));
Q_MX04 U4224 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][564] ), .A1(\_zzLB[1][564] ), .A2(\_zzLB[2][564] ), .A3(\_zzLB[3][564] ), .Z(odata[532]));
Q_MX04 U4225 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][565] ), .A1(\_zzLB[1][565] ), .A2(\_zzLB[2][565] ), .A3(\_zzLB[3][565] ), .Z(odata[533]));
Q_MX04 U4226 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][566] ), .A1(\_zzLB[1][566] ), .A2(\_zzLB[2][566] ), .A3(\_zzLB[3][566] ), .Z(odata[534]));
Q_MX04 U4227 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][567] ), .A1(\_zzLB[1][567] ), .A2(\_zzLB[2][567] ), .A3(\_zzLB[3][567] ), .Z(odata[535]));
Q_MX04 U4228 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][568] ), .A1(\_zzLB[1][568] ), .A2(\_zzLB[2][568] ), .A3(\_zzLB[3][568] ), .Z(odata[536]));
Q_MX04 U4229 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][569] ), .A1(\_zzLB[1][569] ), .A2(\_zzLB[2][569] ), .A3(\_zzLB[3][569] ), .Z(odata[537]));
Q_MX04 U4230 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][570] ), .A1(\_zzLB[1][570] ), .A2(\_zzLB[2][570] ), .A3(\_zzLB[3][570] ), .Z(odata[538]));
Q_MX04 U4231 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][571] ), .A1(\_zzLB[1][571] ), .A2(\_zzLB[2][571] ), .A3(\_zzLB[3][571] ), .Z(odata[539]));
Q_MX04 U4232 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][572] ), .A1(\_zzLB[1][572] ), .A2(\_zzLB[2][572] ), .A3(\_zzLB[3][572] ), .Z(odata[540]));
Q_MX04 U4233 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][573] ), .A1(\_zzLB[1][573] ), .A2(\_zzLB[2][573] ), .A3(\_zzLB[3][573] ), .Z(odata[541]));
Q_MX04 U4234 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][574] ), .A1(\_zzLB[1][574] ), .A2(\_zzLB[2][574] ), .A3(\_zzLB[3][574] ), .Z(odata[542]));
Q_MX04 U4235 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][575] ), .A1(\_zzLB[1][575] ), .A2(\_zzLB[2][575] ), .A3(\_zzLB[3][575] ), .Z(odata[543]));
Q_MX04 U4236 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][576] ), .A1(\_zzLB[1][576] ), .A2(\_zzLB[2][576] ), .A3(\_zzLB[3][576] ), .Z(odata[544]));
Q_MX04 U4237 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][577] ), .A1(\_zzLB[1][577] ), .A2(\_zzLB[2][577] ), .A3(\_zzLB[3][577] ), .Z(odata[545]));
Q_MX04 U4238 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][578] ), .A1(\_zzLB[1][578] ), .A2(\_zzLB[2][578] ), .A3(\_zzLB[3][578] ), .Z(odata[546]));
Q_MX04 U4239 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][579] ), .A1(\_zzLB[1][579] ), .A2(\_zzLB[2][579] ), .A3(\_zzLB[3][579] ), .Z(odata[547]));
Q_MX04 U4240 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][580] ), .A1(\_zzLB[1][580] ), .A2(\_zzLB[2][580] ), .A3(\_zzLB[3][580] ), .Z(odata[548]));
Q_MX04 U4241 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][581] ), .A1(\_zzLB[1][581] ), .A2(\_zzLB[2][581] ), .A3(\_zzLB[3][581] ), .Z(odata[549]));
Q_MX04 U4242 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][582] ), .A1(\_zzLB[1][582] ), .A2(\_zzLB[2][582] ), .A3(\_zzLB[3][582] ), .Z(odata[550]));
Q_MX04 U4243 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][583] ), .A1(\_zzLB[1][583] ), .A2(\_zzLB[2][583] ), .A3(\_zzLB[3][583] ), .Z(odata[551]));
Q_MX04 U4244 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][584] ), .A1(\_zzLB[1][584] ), .A2(\_zzLB[2][584] ), .A3(\_zzLB[3][584] ), .Z(odata[552]));
Q_MX04 U4245 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][585] ), .A1(\_zzLB[1][585] ), .A2(\_zzLB[2][585] ), .A3(\_zzLB[3][585] ), .Z(odata[553]));
Q_MX04 U4246 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][586] ), .A1(\_zzLB[1][586] ), .A2(\_zzLB[2][586] ), .A3(\_zzLB[3][586] ), .Z(odata[554]));
Q_MX04 U4247 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][587] ), .A1(\_zzLB[1][587] ), .A2(\_zzLB[2][587] ), .A3(\_zzLB[3][587] ), .Z(odata[555]));
Q_MX04 U4248 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][588] ), .A1(\_zzLB[1][588] ), .A2(\_zzLB[2][588] ), .A3(\_zzLB[3][588] ), .Z(odata[556]));
Q_MX04 U4249 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][589] ), .A1(\_zzLB[1][589] ), .A2(\_zzLB[2][589] ), .A3(\_zzLB[3][589] ), .Z(odata[557]));
Q_MX04 U4250 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][590] ), .A1(\_zzLB[1][590] ), .A2(\_zzLB[2][590] ), .A3(\_zzLB[3][590] ), .Z(odata[558]));
Q_MX04 U4251 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][591] ), .A1(\_zzLB[1][591] ), .A2(\_zzLB[2][591] ), .A3(\_zzLB[3][591] ), .Z(odata[559]));
Q_MX04 U4252 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][592] ), .A1(\_zzLB[1][592] ), .A2(\_zzLB[2][592] ), .A3(\_zzLB[3][592] ), .Z(oreq));
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m1 "_zzLB 1 592 0 0 3"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_NON_CMM "1"
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE "ixc_gfifo_port"
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE_LIB "IXCOM_TEMP_LIBRARY"
// pragma CVASTRPROP MODULE HDLICE PROP_IXCOM_MOD TRUE
endmodule
