architecture module of cr_kme_regs_flops is
  component ixc_assign
    generic (
      W : integer := 1
    ) ;
    port (
      L : out std_logic_vector((W - 1) downto 0) ;
    R : in std_logic_vector((W - 1) downto 0) := (others => 'X') ) ;
  end component ;

  signal DUMMY0 : std_logic_vector(0 to 31) ;
  signal DUMMY1 : std_logic_vector(0 to 31) ;
  signal DUMMY2 : std_logic_vector(0 to 31) ;
  signal DUMMY3 : std_logic_vector(0 to 31) ;
  signal DUMMY4 : std_logic_vector(0 to 12) ;
  signal DUMMY5 : std_logic_vector(0 to 11) ;
  signal DUMMY6 : std_logic_vector(0 to 1) ;
  signal DUMMY7 : std_logic_vector(0 to 31) ;
  signal DUMMY8 : std_logic_vector(0 to 31) ;
  signal DUMMY9 : std_logic_vector(0 to 31) ;
  signal DUMMY10 : std_logic_vector(0 to 12) ;
  signal DUMMY11 : std_logic_vector(0 to 11) ;
  signal DUMMY12 : std_logic_vector(0 to 1) ;
  signal DUMMY13 : std_logic_vector(0 to 31) ;
  signal DUMMY14 : std_logic_vector(0 to 31) ;
  signal DUMMY15 : std_logic_vector(0 to 31) ;
  signal DUMMY16 : std_logic_vector(0 to 12) ;
  signal DUMMY17 : std_logic_vector(0 to 11) ;
  signal DUMMY18 : std_logic_vector(0 to 1) ;
  signal DUMMY19 : std_logic_vector(0 to 31) ;
  signal DUMMY20 : std_logic_vector(0 to 31) ;
  signal DUMMY21 : std_logic_vector(0 to 31) ;
  signal DUMMY22 : std_logic_vector(0 to 12) ;
  signal DUMMY23 : std_logic_vector(0 to 11) ;
  signal DUMMY24 : std_logic_vector(0 to 1) ;
  signal DUMMY25 : std_logic_vector(0 to 31) ;
  signal DUMMY26 : std_logic_vector(0 to 31) ;
  signal DUMMY27 : std_logic_vector(0 to 31) ;
  signal DUMMY28 : std_logic_vector(0 to 12) ;
  signal DUMMY29 : std_logic_vector(0 to 11) ;
  signal DUMMY30 : std_logic_vector(0 to 1) ;
  signal DUMMY31 : std_logic_vector(0 to 31) ;
  signal DUMMY32 : std_logic_vector(0 to 31) ;
  signal DUMMY33 : std_logic_vector(0 to 31) ;
  signal DUMMY34 : std_logic_vector(0 to 12) ;
  signal DUMMY35 : std_logic_vector(0 to 11) ;
  signal DUMMY36 : std_logic_vector(0 to 1) ;
  signal DUMMY37 : std_logic_vector(0 to 31) ;
  signal DUMMY38 : std_logic_vector(0 to 31) ;
  signal DUMMY39 : std_logic_vector(0 to 31) ;
  signal DUMMY40 : std_logic_vector(0 to 12) ;
  signal DUMMY41 : std_logic_vector(0 to 11) ;
  signal DUMMY42 : std_logic_vector(0 to 1) ;
  signal DUMMY43 : std_logic_vector(0 to 31) ;
  signal DUMMY44 : std_logic_vector(0 to 31) ;
  signal DUMMY45 : std_logic_vector(0 to 31) ;
  signal DUMMY46 : std_logic_vector(0 to 12) ;
  signal DUMMY47 : std_logic_vector(0 to 11) ;
  signal DUMMY48 : std_logic_vector(0 to 1) ;
  signal DUMMY49 : std_logic_vector(0 to 31) ;
  signal DUMMY50 : std_logic_vector(0 to 31) ;
  signal DUMMY51 : std_logic_vector(0 to 18) ;
  signal DUMMY52 : std_logic_vector(0 to 20) ;
  signal DUMMY53 : std_logic_vector(0 to 16) ;
  signal DUMMY54 : std_logic_vector(0 to 17) ;
  signal DUMMY55 : std_logic_vector(0 to 15) ;
  signal DUMMY56 : std_logic_vector(0 to 31) ;
  signal DUMMY57 : std_logic_vector(0 to 31) ;
  signal DUMMY58 : std_logic_vector(0 to 31) ;
  signal DUMMY59 : std_logic_vector(0 to 31) ;
  signal DUMMY60 : std_logic_vector(0 to 31) ;
  signal DUMMY61 : std_logic_vector(0 to 31) ;
  signal DUMMY62 : std_logic_vector(0 to 31) ;
  signal DUMMY63 : std_logic_vector(0 to 31) ;
  signal DUMMY64 : std_logic_vector(0 to 15) ;
  signal DUMMY65 : std_logic_vector(0 to 31) ;
  signal DUMMY66 : std_logic_vector(0 to 31) ;
  signal DUMMY67 : std_logic_vector(0 to 31) ;
  signal DUMMY68 : std_logic_vector(0 to 31) ;
  signal DUMMY69 : std_logic_vector(0 to 31) ;
  signal DUMMY70 : std_logic_vector(0 to 31) ;
  signal DUMMY71 : std_logic_vector(0 to 31) ;
  signal DUMMY72 : std_logic_vector(0 to 31) ;
  signal DUMMY73 : std_logic_vector(0 to 15) ;
  signal DUMMY74 : std_logic_vector(0 to 31) ;
  signal DUMMY75 : std_logic_vector(0 to 31) ;
  signal DUMMY76 : std_logic_vector(0 to 31) ;
  signal DUMMY77 : std_logic_vector(0 to 31) ;
  signal DUMMY78 : std_logic_vector(0 to 31) ;
  signal DUMMY79 : std_logic_vector(0 to 31) ;
  signal DUMMY80 : std_logic_vector(0 to 31) ;
  signal DUMMY81 : std_logic_vector(0 to 31) ;
  signal DUMMY82 : std_logic_vector(0 to 15) ;
  signal DUMMY83 : std_logic_vector(0 to 31) ;
  signal DUMMY84 : std_logic_vector(0 to 31) ;
  signal DUMMY85 : std_logic_vector(0 to 31) ;
  signal DUMMY86 : std_logic_vector(0 to 31) ;
  signal DUMMY87 : std_logic_vector(0 to 31) ;
  signal DUMMY88 : std_logic_vector(0 to 31) ;
  signal DUMMY89 : std_logic_vector(0 to 31) ;
  signal DUMMY90 : std_logic_vector(0 to 31) ;
  signal DUMMY91 : std_logic_vector(0 to 15) ;
  signal DUMMY92 : std_logic_vector(0 to 31) ;
  signal DUMMY93 : std_logic_vector(0 to 31) ;
  signal DUMMY94 : std_logic_vector(0 to 31) ;
  signal DUMMY95 : std_logic_vector(0 to 31) ;
  signal DUMMY96 : std_logic_vector(0 to 31) ;
  signal DUMMY97 : std_logic_vector(0 to 31) ;
  signal DUMMY98 : std_logic_vector(0 to 31) ;
  signal DUMMY99 : std_logic_vector(0 to 31) ;
  signal DUMMY100 : std_logic_vector(0 to 15) ;
  signal DUMMY101 : std_logic_vector(0 to 31) ;
  signal DUMMY102 : std_logic_vector(0 to 31) ;
  signal DUMMY103 : std_logic_vector(0 to 31) ;
  signal DUMMY104 : std_logic_vector(0 to 31) ;
  signal DUMMY105 : std_logic_vector(0 to 31) ;
  signal DUMMY106 : std_logic_vector(0 to 31) ;
  signal DUMMY107 : std_logic_vector(0 to 31) ;
  signal DUMMY108 : std_logic_vector(0 to 31) ;
  signal DUMMY109 : std_logic_vector(0 to 15) ;
  signal DUMMY110 : std_logic_vector(0 to 31) ;
  signal DUMMY111 : std_logic_vector(0 to 31) ;
  signal DUMMY112 : std_logic_vector(0 to 31) ;
  signal DUMMY113 : std_logic_vector(0 to 31) ;
  signal DUMMY114 : std_logic_vector(0 to 31) ;
  signal DUMMY115 : std_logic_vector(0 to 31) ;
  signal DUMMY116 : std_logic_vector(0 to 31) ;
  signal DUMMY117 : std_logic_vector(0 to 31) ;
  signal DUMMY118 : std_logic_vector(0 to 15) ;
  signal DUMMY119 : std_logic_vector(0 to 31) ;
  signal DUMMY120 : std_logic_vector(0 to 31) ;
  signal DUMMY121 : std_logic_vector(0 to 31) ;
  signal DUMMY122 : std_logic_vector(0 to 31) ;
  signal DUMMY123 : std_logic_vector(0 to 31) ;
  signal DUMMY124 : std_logic_vector(0 to 31) ;
  signal DUMMY125 : std_logic_vector(0 to 31) ;
  signal DUMMY126 : std_logic_vector(0 to 31) ;
  signal DUMMY127 : std_logic_vector(0 to 1) ;
  signal DUMMY128 : std_logic_vector(0 to 31) ;
  signal DUMMY129 : std_logic_vector(0 to 31) ;
  signal DUMMY130 : std_logic_vector(0 to 31) ;
  signal DUMMY131 : std_logic_vector(0 to 31) ;
  signal DUMMY132 : std_logic_vector(0 to 31) ;
  signal DUMMY133 : std_logic_vector(0 to 31) ;
  signal DUMMY134 : std_logic_vector(0 to 31) ;
  signal DUMMY135 : std_logic_vector(0 to 31) ;
  signal DUMMY136 : std_logic_vector(0 to 31) ;
  signal DUMMY137 : std_logic_vector(0 to 31) ;
  signal DUMMY138 : std_logic_vector(0 to 31) ;
  signal DUMMY139 : std_logic_vector(0 to 31) ;
  signal DUMMY140 : std_logic_vector(0 to 31) ;
  signal DUMMY141 : std_logic_vector(0 to 15) ;
  signal DUMMY142 : std_logic_vector(0 to 31) ;
  signal DUMMY143 : std_logic_vector(0 to 31) ;
  signal DUMMY144 : std_logic_vector(0 to 31) ;
  signal DUMMY145 : std_logic_vector(0 to 31) ;
  signal DUMMY146 : std_logic_vector(0 to 31) ;
  signal DUMMY147 : std_logic_vector(0 to 31) ;
  signal DUMMY148 : std_logic_vector(0 to 31) ;
  signal DUMMY149 : std_logic_vector(0 to 31) ;
  signal DUMMY150 : std_logic_vector(0 to 31) ;
  signal DUMMY151 : std_logic_vector(0 to 31) ;
  signal DUMMY152 : std_logic_vector(0 to 31) ;
  signal DUMMY153 : std_logic_vector(0 to 31) ;
  signal DUMMY154 : std_logic_vector(0 to 31) ;
  signal DUMMY155 : std_logic_vector(0 to 15) ;
  signal DUMMY156 : std_logic_vector(0 to 4) ;
  signal DUMMY157 : std_logic_vector(0 to 4) ;
  signal DUMMY158 : std_logic_vector(0 to 7) ;
  signal DUMMY159 : std_logic_vector(0 to 6) ;
  signal DUMMY160 : std_logic_vector(0 to 31) ;
  signal DUMMY161 : std_logic_vector(0 to 31) ;
  signal DUMMY162 : std_logic_vector(0 to 31) ;
  signal DUMMY163 : std_logic_vector(0 to 31) ;
  signal DUMMY164 : std_logic_vector(0 to 28) ;
  signal DUMMY165 : std_logic_vector(0 to 10) ;
  signal DUMMY166 : std_logic_vector(0 to 31) ;
  signal DUMMY167 : std_logic_vector(0 to 31) ;
  signal DUMMY168 : std_logic_vector(0 to 9) ;
  signal DUMMY169 : std_logic_vector(0 to 9) ;
  signal DUMMY170 : std_logic_vector(0 to 9) ;
  signal DUMMY171 : std_logic_vector(0 to 9) ;
  signal DUMMY172 : std_logic_vector(0 to 15) ;
  signal DUMMY173 : std_logic_vector(0 to 8) ;
  signal DUMMY174 : std_logic_vector(0 to 31) ;
  signal DUMMY175 : std_logic_vector(0 to 31) ;
  signal DUMMY176 : std_logic_vector(0 to 31) ;
  signal DUMMY177 : std_logic_vector(0 to 8) ;
  signal DUMMY178 : std_logic_vector(0 to 31) ;
  signal DUMMY179 : std_logic_vector(0 to 31) ;
  signal DUMMY180 : std_logic_vector(0 to 8) ;
  signal DUMMY181 : std_logic_vector(0 to 6) ;
  signal DUMMY182 : std_logic_vector(0 to 6) ;
  signal DUMMY183 : std_logic_vector(0 to 6) ;
  signal DUMMY184 : std_logic_vector(0 to 31) ;
  signal DUMMY185 : std_logic_vector(0 to 31) ;
  signal DUMMY186 : std_logic_vector(0 to 8) ;
  signal DUMMY187 : std_logic_vector(0 to 31) ;

begin
  _zz_strnp_0 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY0
      ,o_spare_config
    ) ;
  _zz_strnp_1 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY1
      ,o_cceip0_out_ia_wdata_part0
    ) ;
  _zz_strnp_2 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY2
      ,o_cceip0_out_ia_wdata_part1
    ) ;
  _zz_strnp_3 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY3
      ,o_cceip0_out_ia_wdata_part2
    ) ;
  _zz_strnp_4 : ixc_assign
    generic map(W => 13)
    port map (
       DUMMY4
      ,o_cceip0_out_ia_config
    ) ;
  _zz_strnp_5 : ixc_assign
    generic map(W => 12)
    port map (
       DUMMY5
      ,o_cceip0_out_im_config
    ) ;
  _zz_strnp_6 : ixc_assign
    generic map(W => 2)
    port map (
       DUMMY6
      ,o_cceip0_out_im_read_done
    ) ;
  _zz_strnp_7 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY7
      ,o_cceip1_out_ia_wdata_part0
    ) ;
  _zz_strnp_8 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY8
      ,o_cceip1_out_ia_wdata_part1
    ) ;
  _zz_strnp_9 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY9
      ,o_cceip1_out_ia_wdata_part2
    ) ;
  _zz_strnp_10 : ixc_assign
    generic map(W => 13)
    port map (
       DUMMY10
      ,o_cceip1_out_ia_config
    ) ;
  _zz_strnp_11 : ixc_assign
    generic map(W => 12)
    port map (
       DUMMY11
      ,o_cceip1_out_im_config
    ) ;
  _zz_strnp_12 : ixc_assign
    generic map(W => 2)
    port map (
       DUMMY12
      ,o_cceip1_out_im_read_done
    ) ;
  _zz_strnp_13 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY13
      ,o_cceip2_out_ia_wdata_part0
    ) ;
  _zz_strnp_14 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY14
      ,o_cceip2_out_ia_wdata_part1
    ) ;
  _zz_strnp_15 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY15
      ,o_cceip2_out_ia_wdata_part2
    ) ;
  _zz_strnp_16 : ixc_assign
    generic map(W => 13)
    port map (
       DUMMY16
      ,o_cceip2_out_ia_config
    ) ;
  _zz_strnp_17 : ixc_assign
    generic map(W => 12)
    port map (
       DUMMY17
      ,o_cceip2_out_im_config
    ) ;
  _zz_strnp_18 : ixc_assign
    generic map(W => 2)
    port map (
       DUMMY18
      ,o_cceip2_out_im_read_done
    ) ;
  _zz_strnp_19 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY19
      ,o_cceip3_out_ia_wdata_part0
    ) ;
  _zz_strnp_20 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY20
      ,o_cceip3_out_ia_wdata_part1
    ) ;
  _zz_strnp_21 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY21
      ,o_cceip3_out_ia_wdata_part2
    ) ;
  _zz_strnp_22 : ixc_assign
    generic map(W => 13)
    port map (
       DUMMY22
      ,o_cceip3_out_ia_config
    ) ;
  _zz_strnp_23 : ixc_assign
    generic map(W => 12)
    port map (
       DUMMY23
      ,o_cceip3_out_im_config
    ) ;
  _zz_strnp_24 : ixc_assign
    generic map(W => 2)
    port map (
       DUMMY24
      ,o_cceip3_out_im_read_done
    ) ;
  _zz_strnp_25 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY25
      ,o_cddip0_out_ia_wdata_part0
    ) ;
  _zz_strnp_26 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY26
      ,o_cddip0_out_ia_wdata_part1
    ) ;
  _zz_strnp_27 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY27
      ,o_cddip0_out_ia_wdata_part2
    ) ;
  _zz_strnp_28 : ixc_assign
    generic map(W => 13)
    port map (
       DUMMY28
      ,o_cddip0_out_ia_config
    ) ;
  _zz_strnp_29 : ixc_assign
    generic map(W => 12)
    port map (
       DUMMY29
      ,o_cddip0_out_im_config
    ) ;
  _zz_strnp_30 : ixc_assign
    generic map(W => 2)
    port map (
       DUMMY30
      ,o_cddip0_out_im_read_done
    ) ;
  _zz_strnp_31 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY31
      ,o_cddip1_out_ia_wdata_part0
    ) ;
  _zz_strnp_32 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY32
      ,o_cddip1_out_ia_wdata_part1
    ) ;
  _zz_strnp_33 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY33
      ,o_cddip1_out_ia_wdata_part2
    ) ;
  _zz_strnp_34 : ixc_assign
    generic map(W => 13)
    port map (
       DUMMY34
      ,o_cddip1_out_ia_config
    ) ;
  _zz_strnp_35 : ixc_assign
    generic map(W => 12)
    port map (
       DUMMY35
      ,o_cddip1_out_im_config
    ) ;
  _zz_strnp_36 : ixc_assign
    generic map(W => 2)
    port map (
       DUMMY36
      ,o_cddip1_out_im_read_done
    ) ;
  _zz_strnp_37 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY37
      ,o_cddip2_out_ia_wdata_part0
    ) ;
  _zz_strnp_38 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY38
      ,o_cddip2_out_ia_wdata_part1
    ) ;
  _zz_strnp_39 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY39
      ,o_cddip2_out_ia_wdata_part2
    ) ;
  _zz_strnp_40 : ixc_assign
    generic map(W => 13)
    port map (
       DUMMY40
      ,o_cddip2_out_ia_config
    ) ;
  _zz_strnp_41 : ixc_assign
    generic map(W => 12)
    port map (
       DUMMY41
      ,o_cddip2_out_im_config
    ) ;
  _zz_strnp_42 : ixc_assign
    generic map(W => 2)
    port map (
       DUMMY42
      ,o_cddip2_out_im_read_done
    ) ;
  _zz_strnp_43 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY43
      ,o_cddip3_out_ia_wdata_part0
    ) ;
  _zz_strnp_44 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY44
      ,o_cddip3_out_ia_wdata_part1
    ) ;
  _zz_strnp_45 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY45
      ,o_cddip3_out_ia_wdata_part2
    ) ;
  _zz_strnp_46 : ixc_assign
    generic map(W => 13)
    port map (
       DUMMY46
      ,o_cddip3_out_ia_config
    ) ;
  _zz_strnp_47 : ixc_assign
    generic map(W => 12)
    port map (
       DUMMY47
      ,o_cddip3_out_im_config
    ) ;
  _zz_strnp_48 : ixc_assign
    generic map(W => 2)
    port map (
       DUMMY48
      ,o_cddip3_out_im_read_done
    ) ;
  _zz_strnp_49 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY49
      ,o_ckv_ia_wdata_part0
    ) ;
  _zz_strnp_50 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY50
      ,o_ckv_ia_wdata_part1
    ) ;
  _zz_strnp_51 : ixc_assign
    generic map(W => 19)
    port map (
       DUMMY51
      ,o_ckv_ia_config
    ) ;
  _zz_strnp_52 : ixc_assign
    generic map(W => 21)
    port map (
       DUMMY52
      ,o_kim_ia_wdata_part0
    ) ;
  _zz_strnp_53 : ixc_assign
    generic map(W => 17)
    port map (
       DUMMY53
      ,o_kim_ia_wdata_part1
    ) ;
  _zz_strnp_54 : ixc_assign
    generic map(W => 18)
    port map (
       DUMMY54
      ,o_kim_ia_config
    ) ;
  _zz_strnp_55 : ixc_assign
    generic map(W => 16)
    port map (
       DUMMY55
      ,o_label0_config
    ) ;
  _zz_strnp_56 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY56
      ,o_label0_data7
    ) ;
  _zz_strnp_57 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY57
      ,o_label0_data6
    ) ;
  _zz_strnp_58 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY58
      ,o_label0_data5
    ) ;
  _zz_strnp_59 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY59
      ,o_label0_data4
    ) ;
  _zz_strnp_60 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY60
      ,o_label0_data3
    ) ;
  _zz_strnp_61 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY61
      ,o_label0_data2
    ) ;
  _zz_strnp_62 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY62
      ,o_label0_data1
    ) ;
  _zz_strnp_63 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY63
      ,o_label0_data0
    ) ;
  _zz_strnp_64 : ixc_assign
    generic map(W => 16)
    port map (
       DUMMY64
      ,o_label1_config
    ) ;
  _zz_strnp_65 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY65
      ,o_label1_data7
    ) ;
  _zz_strnp_66 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY66
      ,o_label1_data6
    ) ;
  _zz_strnp_67 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY67
      ,o_label1_data5
    ) ;
  _zz_strnp_68 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY68
      ,o_label1_data4
    ) ;
  _zz_strnp_69 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY69
      ,o_label1_data3
    ) ;
  _zz_strnp_70 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY70
      ,o_label1_data2
    ) ;
  _zz_strnp_71 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY71
      ,o_label1_data1
    ) ;
  _zz_strnp_72 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY72
      ,o_label1_data0
    ) ;
  _zz_strnp_73 : ixc_assign
    generic map(W => 16)
    port map (
       DUMMY73
      ,o_label2_config
    ) ;
  _zz_strnp_74 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY74
      ,o_label2_data7
    ) ;
  _zz_strnp_75 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY75
      ,o_label2_data6
    ) ;
  _zz_strnp_76 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY76
      ,o_label2_data5
    ) ;
  _zz_strnp_77 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY77
      ,o_label2_data4
    ) ;
  _zz_strnp_78 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY78
      ,o_label2_data3
    ) ;
  _zz_strnp_79 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY79
      ,o_label2_data2
    ) ;
  _zz_strnp_80 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY80
      ,o_label2_data1
    ) ;
  _zz_strnp_81 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY81
      ,o_label2_data0
    ) ;
  _zz_strnp_82 : ixc_assign
    generic map(W => 16)
    port map (
       DUMMY82
      ,o_label3_config
    ) ;
  _zz_strnp_83 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY83
      ,o_label3_data7
    ) ;
  _zz_strnp_84 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY84
      ,o_label3_data6
    ) ;
  _zz_strnp_85 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY85
      ,o_label3_data5
    ) ;
  _zz_strnp_86 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY86
      ,o_label3_data4
    ) ;
  _zz_strnp_87 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY87
      ,o_label3_data3
    ) ;
  _zz_strnp_88 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY88
      ,o_label3_data2
    ) ;
  _zz_strnp_89 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY89
      ,o_label3_data1
    ) ;
  _zz_strnp_90 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY90
      ,o_label3_data0
    ) ;
  _zz_strnp_91 : ixc_assign
    generic map(W => 16)
    port map (
       DUMMY91
      ,o_label4_config
    ) ;
  _zz_strnp_92 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY92
      ,o_label4_data7
    ) ;
  _zz_strnp_93 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY93
      ,o_label4_data6
    ) ;
  _zz_strnp_94 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY94
      ,o_label4_data5
    ) ;
  _zz_strnp_95 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY95
      ,o_label4_data4
    ) ;
  _zz_strnp_96 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY96
      ,o_label4_data3
    ) ;
  _zz_strnp_97 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY97
      ,o_label4_data2
    ) ;
  _zz_strnp_98 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY98
      ,o_label4_data1
    ) ;
  _zz_strnp_99 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY99
      ,o_label4_data0
    ) ;
  _zz_strnp_100 : ixc_assign
    generic map(W => 16)
    port map (
       DUMMY100
      ,o_label5_config
    ) ;
  _zz_strnp_101 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY101
      ,o_label5_data7
    ) ;
  _zz_strnp_102 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY102
      ,o_label5_data6
    ) ;
  _zz_strnp_103 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY103
      ,o_label5_data5
    ) ;
  _zz_strnp_104 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY104
      ,o_label5_data4
    ) ;
  _zz_strnp_105 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY105
      ,o_label5_data3
    ) ;
  _zz_strnp_106 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY106
      ,o_label5_data2
    ) ;
  _zz_strnp_107 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY107
      ,o_label5_data1
    ) ;
  _zz_strnp_108 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY108
      ,o_label5_data0
    ) ;
  _zz_strnp_109 : ixc_assign
    generic map(W => 16)
    port map (
       DUMMY109
      ,o_label6_config
    ) ;
  _zz_strnp_110 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY110
      ,o_label6_data7
    ) ;
  _zz_strnp_111 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY111
      ,o_label6_data6
    ) ;
  _zz_strnp_112 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY112
      ,o_label6_data5
    ) ;
  _zz_strnp_113 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY113
      ,o_label6_data4
    ) ;
  _zz_strnp_114 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY114
      ,o_label6_data3
    ) ;
  _zz_strnp_115 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY115
      ,o_label6_data2
    ) ;
  _zz_strnp_116 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY116
      ,o_label6_data1
    ) ;
  _zz_strnp_117 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY117
      ,o_label6_data0
    ) ;
  _zz_strnp_118 : ixc_assign
    generic map(W => 16)
    port map (
       DUMMY118
      ,o_label7_config
    ) ;
  _zz_strnp_119 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY119
      ,o_label7_data7
    ) ;
  _zz_strnp_120 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY120
      ,o_label7_data6
    ) ;
  _zz_strnp_121 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY121
      ,o_label7_data5
    ) ;
  _zz_strnp_122 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY122
      ,o_label7_data4
    ) ;
  _zz_strnp_123 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY123
      ,o_label7_data3
    ) ;
  _zz_strnp_124 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY124
      ,o_label7_data2
    ) ;
  _zz_strnp_125 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY125
      ,o_label7_data1
    ) ;
  _zz_strnp_126 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY126
      ,o_label7_data0
    ) ;
  _zz_strnp_127 : ixc_assign
    generic map(W => 2)
    port map (
       DUMMY127
      ,o_kdf_drbg_ctrl
    ) ;
  _zz_strnp_128 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY128
      ,o_kdf_drbg_seed_0_state_key_31_0
    ) ;
  _zz_strnp_129 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY129
      ,o_kdf_drbg_seed_0_state_key_63_32
    ) ;
  _zz_strnp_130 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY130
      ,o_kdf_drbg_seed_0_state_key_95_64
    ) ;
  _zz_strnp_131 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY131
      ,o_kdf_drbg_seed_0_state_key_127_96
    ) ;
  _zz_strnp_132 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY132
      ,o_kdf_drbg_seed_0_state_key_159_128
    ) ;
  _zz_strnp_133 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY133
      ,o_kdf_drbg_seed_0_state_key_191_160
    ) ;
  _zz_strnp_134 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY134
      ,o_kdf_drbg_seed_0_state_key_223_192
    ) ;
  _zz_strnp_135 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY135
      ,o_kdf_drbg_seed_0_state_key_255_224
    ) ;
  _zz_strnp_136 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY136
      ,o_kdf_drbg_seed_0_state_value_31_0
    ) ;
  _zz_strnp_137 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY137
      ,o_kdf_drbg_seed_0_state_value_63_32
    ) ;
  _zz_strnp_138 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY138
      ,o_kdf_drbg_seed_0_state_value_95_64
    ) ;
  _zz_strnp_139 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY139
      ,o_kdf_drbg_seed_0_state_value_127_96
    ) ;
  _zz_strnp_140 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY140
      ,o_kdf_drbg_seed_0_reseed_interval_0
    ) ;
  _zz_strnp_141 : ixc_assign
    generic map(W => 16)
    port map (
       DUMMY141
      ,o_kdf_drbg_seed_0_reseed_interval_1
    ) ;
  _zz_strnp_142 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY142
      ,o_kdf_drbg_seed_1_state_key_31_0
    ) ;
  _zz_strnp_143 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY143
      ,o_kdf_drbg_seed_1_state_key_63_32
    ) ;
  _zz_strnp_144 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY144
      ,o_kdf_drbg_seed_1_state_key_95_64
    ) ;
  _zz_strnp_145 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY145
      ,o_kdf_drbg_seed_1_state_key_127_96
    ) ;
  _zz_strnp_146 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY146
      ,o_kdf_drbg_seed_1_state_key_159_128
    ) ;
  _zz_strnp_147 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY147
      ,o_kdf_drbg_seed_1_state_key_191_160
    ) ;
  _zz_strnp_148 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY148
      ,o_kdf_drbg_seed_1_state_key_223_192
    ) ;
  _zz_strnp_149 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY149
      ,o_kdf_drbg_seed_1_state_key_255_224
    ) ;
  _zz_strnp_150 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY150
      ,o_kdf_drbg_seed_1_state_value_31_0
    ) ;
  _zz_strnp_151 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY151
      ,o_kdf_drbg_seed_1_state_value_63_32
    ) ;
  _zz_strnp_152 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY152
      ,o_kdf_drbg_seed_1_state_value_95_64
    ) ;
  _zz_strnp_153 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY153
      ,o_kdf_drbg_seed_1_state_value_127_96
    ) ;
  _zz_strnp_154 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY154
      ,o_kdf_drbg_seed_1_reseed_interval_0
    ) ;
  _zz_strnp_155 : ixc_assign
    generic map(W => 16)
    port map (
       DUMMY155
      ,o_kdf_drbg_seed_1_reseed_interval_1
    ) ;
  _zz_strnp_156 : ixc_assign
    generic map(W => 5)
    port map (
       DUMMY156
      ,o_interrupt_status
    ) ;
  _zz_strnp_157 : ixc_assign
    generic map(W => 5)
    port map (
       DUMMY157
      ,o_interrupt_mask
    ) ;
  _zz_strnp_158 : ixc_assign
    generic map(W => 8)
    port map (
       DUMMY158
      ,o_engine_sticky_status
    ) ;
  _zz_strnp_159 : ixc_assign
    generic map(W => 7)
    port map (
       DUMMY159
      ,o_bimc_monitor_mask
    ) ;
  _zz_strnp_160 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY160
      ,o_bimc_ecc_uncorrectable_error_cnt
    ) ;
  _zz_strnp_161 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY161
      ,o_bimc_ecc_correctable_error_cnt
    ) ;
  _zz_strnp_162 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY162
      ,o_bimc_parity_error_cnt
    ) ;
  _zz_strnp_163 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY163
      ,o_bimc_global_config
    ) ;
  _zz_strnp_164 : ixc_assign
    generic map(W => 29)
    port map (
       DUMMY164
      ,o_bimc_eccpar_debug
    ) ;
  _zz_strnp_165 : ixc_assign
    generic map(W => 11)
    port map (
       DUMMY165
      ,o_bimc_cmd2
    ) ;
  _zz_strnp_166 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY166
      ,o_bimc_cmd1
    ) ;
  _zz_strnp_167 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY167
      ,o_bimc_cmd0
    ) ;
  _zz_strnp_168 : ixc_assign
    generic map(W => 10)
    port map (
       DUMMY168
      ,o_bimc_rxcmd2
    ) ;
  _zz_strnp_169 : ixc_assign
    generic map(W => 10)
    port map (
       DUMMY169
      ,o_bimc_rxrsp2
    ) ;
  _zz_strnp_170 : ixc_assign
    generic map(W => 10)
    port map (
       DUMMY170
      ,o_bimc_pollrsp2
    ) ;
  _zz_strnp_171 : ixc_assign
    generic map(W => 10)
    port map (
       DUMMY171
      ,o_bimc_dbgcmd2
    ) ;
  _zz_strnp_172 : ixc_assign
    generic map(W => 16)
    port map (
       DUMMY172
      ,o_im_consumed
    ) ;
  _zz_strnp_173 : ixc_assign
    generic map(W => 9)
    port map (
       DUMMY173
      ,o_tready_override
    ) ;
  _zz_strnp_174 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY174
      ,o_regs_sa_ctrl
    ) ;
  _zz_strnp_175 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY175
      ,o_sa_snapshot_ia_wdata_part0
    ) ;
  _zz_strnp_176 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY176
      ,o_sa_snapshot_ia_wdata_part1
    ) ;
  _zz_strnp_177 : ixc_assign
    generic map(W => 9)
    port map (
       DUMMY177
      ,o_sa_snapshot_ia_config
    ) ;
  _zz_strnp_178 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY178
      ,o_sa_count_ia_wdata_part0
    ) ;
  _zz_strnp_179 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY179
      ,o_sa_count_ia_wdata_part1
    ) ;
  _zz_strnp_180 : ixc_assign
    generic map(W => 9)
    port map (
       DUMMY180
      ,o_sa_count_ia_config
    ) ;
  _zz_strnp_181 : ixc_assign
    generic map(W => 7)
    port map (
       DUMMY181
      ,o_cceip_encrypt_kop_fifo_override
    ) ;
  _zz_strnp_182 : ixc_assign
    generic map(W => 7)
    port map (
       DUMMY182
      ,o_cceip_validate_kop_fifo_override
    ) ;
  _zz_strnp_183 : ixc_assign
    generic map(W => 7)
    port map (
       DUMMY183
      ,o_cddip_decrypt_kop_fifo_override
    ) ;
  _zz_strnp_184 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY184
      ,o_sa_global_ctrl
    ) ;
  _zz_strnp_185 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY185
      ,o_sa_ctrl_ia_wdata_part0
    ) ;
  _zz_strnp_186 : ixc_assign
    generic map(W => 9)
    port map (
       DUMMY186
      ,o_sa_ctrl_ia_config
    ) ;
  _zz_strnp_187 : ixc_assign
    generic map(W => 32)
    port map (
       DUMMY187
      ,o_kdf_test_key_size_config
    ) ;

  process --:o413
  (clk,i_reset_)
  begin
    if (i_reset_ = '0') then
      o_spare_config <= "00000000000000000000000000000000" ;
      o_cceip0_out_ia_wdata_part0(5 downto 0) <= "000000" ;
      o_cceip0_out_ia_wdata_part1 <= "00000000000000000000000000000000" ;
      o_cceip0_out_ia_wdata_part2 <= "00000000000000000000000000000000" ;
      o_cceip0_out_ia_config(8 downto 0) <= "000000000" ;
      o_cceip0_out_ia_config(12 downto 9) <= "0000" ;
      o_cceip0_out_im_config(9 downto 0) <= "1000000000" ;
      o_cceip0_out_im_config(11 downto 10) <= "11" ;
      o_cceip0_out_im_read_done(0 downto 0) <= "0" ;
      o_cceip0_out_im_read_done(1 downto 1) <= "0" ;
      o_cceip1_out_ia_wdata_part0(5 downto 0) <= "000000" ;
      o_cceip1_out_ia_wdata_part1 <= "00000000000000000000000000000000" ;
      o_cceip1_out_ia_wdata_part2 <= "00000000000000000000000000000000" ;
      o_cceip1_out_ia_config(8 downto 0) <= "000000000" ;
      o_cceip1_out_ia_config(12 downto 9) <= "0000" ;
      o_cceip1_out_im_config(9 downto 0) <= "1000000000" ;
      o_cceip1_out_im_config(11 downto 10) <= "11" ;
      o_cceip1_out_im_read_done(0 downto 0) <= "0" ;
      o_cceip1_out_im_read_done(1 downto 1) <= "0" ;
      o_cceip2_out_ia_wdata_part0(5 downto 0) <= "000000" ;
      o_cceip2_out_ia_wdata_part1 <= "00000000000000000000000000000000" ;
      o_cceip2_out_ia_wdata_part2 <= "00000000000000000000000000000000" ;
      o_cceip2_out_ia_config(8 downto 0) <= "000000000" ;
      o_cceip2_out_ia_config(12 downto 9) <= "0000" ;
      o_cceip2_out_im_config(9 downto 0) <= "1000000000" ;
      o_cceip2_out_im_config(11 downto 10) <= "11" ;
      o_cceip2_out_im_read_done(0 downto 0) <= "0" ;
      o_cceip2_out_im_read_done(1 downto 1) <= "0" ;
      o_cceip3_out_ia_wdata_part0(5 downto 0) <= "000000" ;
      o_cceip3_out_ia_wdata_part1 <= "00000000000000000000000000000000" ;
      o_cceip3_out_ia_wdata_part2 <= "00000000000000000000000000000000" ;
      o_cceip3_out_ia_config(8 downto 0) <= "000000000" ;
      o_cceip3_out_ia_config(12 downto 9) <= "0000" ;
      o_cceip3_out_im_config(9 downto 0) <= "1000000000" ;
      o_cceip3_out_im_config(11 downto 10) <= "11" ;
      o_cceip3_out_im_read_done(0 downto 0) <= "0" ;
      o_cceip3_out_im_read_done(1 downto 1) <= "0" ;
      o_cddip0_out_ia_wdata_part0(5 downto 0) <= "000000" ;
      o_cddip0_out_ia_wdata_part1 <= "00000000000000000000000000000000" ;
      o_cddip0_out_ia_wdata_part2 <= "00000000000000000000000000000000" ;
      o_cddip0_out_ia_config(8 downto 0) <= "000000000" ;
      o_cddip0_out_ia_config(12 downto 9) <= "0000" ;
      o_cddip0_out_im_config(9 downto 0) <= "1000000000" ;
      o_cddip0_out_im_config(11 downto 10) <= "11" ;
      o_cddip0_out_im_read_done(0 downto 0) <= "0" ;
      o_cddip0_out_im_read_done(1 downto 1) <= "0" ;
      o_cddip1_out_ia_wdata_part0(5 downto 0) <= "000000" ;
      o_cddip1_out_ia_wdata_part1 <= "00000000000000000000000000000000" ;
      o_cddip1_out_ia_wdata_part2 <= "00000000000000000000000000000000" ;
      o_cddip1_out_ia_config(8 downto 0) <= "000000000" ;
      o_cddip1_out_ia_config(12 downto 9) <= "0000" ;
      o_cddip1_out_im_config(9 downto 0) <= "1000000000" ;
      o_cddip1_out_im_config(11 downto 10) <= "11" ;
      o_cddip1_out_im_read_done(0 downto 0) <= "0" ;
      o_cddip1_out_im_read_done(1 downto 1) <= "0" ;
      o_cddip2_out_ia_wdata_part0(5 downto 0) <= "000000" ;
      o_cddip2_out_ia_wdata_part1 <= "00000000000000000000000000000000" ;
      o_cddip2_out_ia_wdata_part2 <= "00000000000000000000000000000000" ;
      o_cddip2_out_ia_config(8 downto 0) <= "000000000" ;
      o_cddip2_out_ia_config(12 downto 9) <= "0000" ;
      o_cddip2_out_im_config(9 downto 0) <= "1000000000" ;
      o_cddip2_out_im_config(11 downto 10) <= "11" ;
      o_cddip2_out_im_read_done(0 downto 0) <= "0" ;
      o_cddip2_out_im_read_done(1 downto 1) <= "0" ;
      o_cddip3_out_ia_wdata_part0(5 downto 0) <= "000000" ;
      o_cddip3_out_ia_wdata_part1 <= "00000000000000000000000000000000" ;
      o_cddip3_out_ia_wdata_part2 <= "00000000000000000000000000000000" ;
      o_cddip3_out_ia_config(8 downto 0) <= "000000000" ;
      o_cddip3_out_ia_config(12 downto 9) <= "0000" ;
      o_cddip3_out_im_config(9 downto 0) <= "1000000000" ;
      o_cddip3_out_im_config(11 downto 10) <= "11" ;
      o_cddip3_out_im_read_done(0 downto 0) <= "0" ;
      o_cddip3_out_im_read_done(1 downto 1) <= "0" ;
      o_ckv_ia_wdata_part0 <= "00000000000000000000000000000000" ;
      o_ckv_ia_wdata_part1 <= "00000000000000000000000000000000" ;
      o_ckv_ia_config(14 downto 0) <= "000000000000000" ;
      o_ckv_ia_config(18 downto 15) <= "0000" ;
      o_kim_ia_wdata_part0(14 downto 0) <= "000000000000000" ;
      o_kim_ia_wdata_part0(16 downto 15) <= "00" ;
      o_kim_ia_wdata_part0(19 downto 17) <= "000" ;
      o_kim_ia_wdata_part0(20 downto 20) <= "0" ;
      o_kim_ia_wdata_part1(0 downto 0) <= "0" ;
      o_kim_ia_wdata_part1(12 downto 1) <= "000000000000" ;
      o_kim_ia_wdata_part1(16 downto 13) <= "0000" ;
      o_kim_ia_config(13 downto 0) <= "00000000000000" ;
      o_kim_ia_config(17 downto 14) <= "0000" ;
      o_label0_config(7 downto 0) <= "00000000" ;
      o_label0_config(8 downto 8) <= "1" ;
      o_label0_config(14 downto 9) <= "000000" ;
      o_label0_config(15 downto 15) <= "0" ;
      o_label0_data7 <= "00000000000000000000000000000000" ;
      o_label0_data6 <= "00000000000000000000000000000000" ;
      o_label0_data5 <= "00000000000000000000000000000000" ;
      o_label0_data4 <= "00000000000000000000000000000000" ;
      o_label0_data3 <= "00000000000000000000000000000000" ;
      o_label0_data2 <= "00000000000000000000000000000000" ;
      o_label0_data1 <= "00000000000000000000000000000000" ;
      o_label0_data0 <= "00000000000000000000000000000000" ;
      o_label1_config(7 downto 0) <= "00000000" ;
      o_label1_config(8 downto 8) <= "1" ;
      o_label1_config(14 downto 9) <= "000000" ;
      o_label1_config(15 downto 15) <= "0" ;
      o_label1_data7 <= "00000000000000000000000000000000" ;
      o_label1_data6 <= "00000000000000000000000000000000" ;
      o_label1_data5 <= "00000000000000000000000000000000" ;
      o_label1_data4 <= "00000000000000000000000000000000" ;
      o_label1_data3 <= "00000000000000000000000000000000" ;
      o_label1_data2 <= "00000000000000000000000000000000" ;
      o_label1_data1 <= "00000000000000000000000000000000" ;
      o_label1_data0 <= "00000000000000000000000000000000" ;
      o_label2_config(7 downto 0) <= "00000000" ;
      o_label2_config(8 downto 8) <= "1" ;
      o_label2_config(14 downto 9) <= "000000" ;
      o_label2_config(15 downto 15) <= "0" ;
      o_label2_data7 <= "00000000000000000000000000000000" ;
      o_label2_data6 <= "00000000000000000000000000000000" ;
      o_label2_data5 <= "00000000000000000000000000000000" ;
      o_label2_data4 <= "00000000000000000000000000000000" ;
      o_label2_data3 <= "00000000000000000000000000000000" ;
      o_label2_data2 <= "00000000000000000000000000000000" ;
      o_label2_data1 <= "00000000000000000000000000000000" ;
      o_label2_data0 <= "00000000000000000000000000000000" ;
      o_label3_config(7 downto 0) <= "00000000" ;
      o_label3_config(8 downto 8) <= "1" ;
      o_label3_config(14 downto 9) <= "000000" ;
      o_label3_config(15 downto 15) <= "0" ;
      o_label3_data7 <= "00000000000000000000000000000000" ;
      o_label3_data6 <= "00000000000000000000000000000000" ;
      o_label3_data5 <= "00000000000000000000000000000000" ;
      o_label3_data4 <= "00000000000000000000000000000000" ;
      o_label3_data3 <= "00000000000000000000000000000000" ;
      o_label3_data2 <= "00000000000000000000000000000000" ;
      o_label3_data1 <= "00000000000000000000000000000000" ;
      o_label3_data0 <= "00000000000000000000000000000000" ;
      o_label4_config(7 downto 0) <= "00000000" ;
      o_label4_config(8 downto 8) <= "1" ;
      o_label4_config(14 downto 9) <= "000000" ;
      o_label4_config(15 downto 15) <= "0" ;
      o_label4_data7 <= "00000000000000000000000000000000" ;
      o_label4_data6 <= "00000000000000000000000000000000" ;
      o_label4_data5 <= "00000000000000000000000000000000" ;
      o_label4_data4 <= "00000000000000000000000000000000" ;
      o_label4_data3 <= "00000000000000000000000000000000" ;
      o_label4_data2 <= "00000000000000000000000000000000" ;
      o_label4_data1 <= "00000000000000000000000000000000" ;
      o_label4_data0 <= "00000000000000000000000000000000" ;
      o_label5_config(7 downto 0) <= "00000000" ;
      o_label5_config(8 downto 8) <= "1" ;
      o_label5_config(14 downto 9) <= "000000" ;
      o_label5_config(15 downto 15) <= "0" ;
      o_label5_data7 <= "00000000000000000000000000000000" ;
      o_label5_data6 <= "00000000000000000000000000000000" ;
      o_label5_data5 <= "00000000000000000000000000000000" ;
      o_label5_data4 <= "00000000000000000000000000000000" ;
      o_label5_data3 <= "00000000000000000000000000000000" ;
      o_label5_data2 <= "00000000000000000000000000000000" ;
      o_label5_data1 <= "00000000000000000000000000000000" ;
      o_label5_data0 <= "00000000000000000000000000000000" ;
      o_label6_config(7 downto 0) <= "00000000" ;
      o_label6_config(8 downto 8) <= "1" ;
      o_label6_config(14 downto 9) <= "000000" ;
      o_label6_config(15 downto 15) <= "0" ;
      o_label6_data7 <= "00000000000000000000000000000000" ;
      o_label6_data6 <= "00000000000000000000000000000000" ;
      o_label6_data5 <= "00000000000000000000000000000000" ;
      o_label6_data4 <= "00000000000000000000000000000000" ;
      o_label6_data3 <= "00000000000000000000000000000000" ;
      o_label6_data2 <= "00000000000000000000000000000000" ;
      o_label6_data1 <= "00000000000000000000000000000000" ;
      o_label6_data0 <= "00000000000000000000000000000000" ;
      o_label7_config(7 downto 0) <= "00000000" ;
      o_label7_config(8 downto 8) <= "1" ;
      o_label7_config(14 downto 9) <= "000000" ;
      o_label7_config(15 downto 15) <= "0" ;
      o_label7_data7 <= "00000000000000000000000000000000" ;
      o_label7_data6 <= "00000000000000000000000000000000" ;
      o_label7_data5 <= "00000000000000000000000000000000" ;
      o_label7_data4 <= "00000000000000000000000000000000" ;
      o_label7_data3 <= "00000000000000000000000000000000" ;
      o_label7_data2 <= "00000000000000000000000000000000" ;
      o_label7_data1 <= "00000000000000000000000000000000" ;
      o_label7_data0 <= "00000000000000000000000000000000" ;
      o_kdf_drbg_ctrl <= "00" ;
      o_kdf_drbg_seed_0_state_key_31_0 <= "00000000000000000000000000000000" ;
      o_kdf_drbg_seed_0_state_key_63_32 <= "00000000000000000000000000000000" ;
      o_kdf_drbg_seed_0_state_key_95_64 <= "00000000000000000000000000000000" ;
      o_kdf_drbg_seed_0_state_key_127_96 <= "00000000000000000000000000000000" ;
      o_kdf_drbg_seed_0_state_key_159_128 <= "00000000000000000000000000000000"
       ;
      o_kdf_drbg_seed_0_state_key_191_160 <= "00000000000000000000000000000000"
       ;
      o_kdf_drbg_seed_0_state_key_223_192 <= "00000000000000000000000000000000"
       ;
      o_kdf_drbg_seed_0_state_key_255_224 <= "00000000000000000000000000000000"
       ;
      o_kdf_drbg_seed_0_state_value_31_0 <= "00000000000000000000000000000000" ;
      o_kdf_drbg_seed_0_state_value_63_32 <= "00000000000000000000000000000000"
       ;
      o_kdf_drbg_seed_0_state_value_95_64 <= "00000000000000000000000000000000"
       ;
      o_kdf_drbg_seed_0_state_value_127_96 <= "00000000000000000000000000000000"
       ;
      o_kdf_drbg_seed_0_reseed_interval_0 <= "00000000000000000000000000000000"
       ;
      o_kdf_drbg_seed_0_reseed_interval_1 <= "0000000000000000" ;
      o_kdf_drbg_seed_1_state_key_31_0 <= "00000000000000000000000000000000" ;
      o_kdf_drbg_seed_1_state_key_63_32 <= "00000000000000000000000000000000" ;
      o_kdf_drbg_seed_1_state_key_95_64 <= "00000000000000000000000000000000" ;
      o_kdf_drbg_seed_1_state_key_127_96 <= "00000000000000000000000000000000" ;
      o_kdf_drbg_seed_1_state_key_159_128 <= "00000000000000000000000000000000"
       ;
      o_kdf_drbg_seed_1_state_key_191_160 <= "00000000000000000000000000000000"
       ;
      o_kdf_drbg_seed_1_state_key_223_192 <= "00000000000000000000000000000000"
       ;
      o_kdf_drbg_seed_1_state_key_255_224 <= "00000000000000000000000000000000"
       ;
      o_kdf_drbg_seed_1_state_value_31_0 <= "00000000000000000000000000000000" ;
      o_kdf_drbg_seed_1_state_value_63_32 <= "00000000000000000000000000000000"
       ;
      o_kdf_drbg_seed_1_state_value_95_64 <= "00000000000000000000000000000000"
       ;
      o_kdf_drbg_seed_1_state_value_127_96 <= "00000000000000000000000000000000"
       ;
      o_kdf_drbg_seed_1_reseed_interval_0 <= "00000000000000000000000000000000"
       ;
      o_kdf_drbg_seed_1_reseed_interval_1 <= "0000000000000000" ;
      o_interrupt_status(0 downto 0) <= "0" ;
      o_interrupt_status(1 downto 1) <= "0" ;
      o_interrupt_status(2 downto 2) <= "0" ;
      o_interrupt_status(3 downto 3) <= "0" ;
      o_interrupt_status(4 downto 4) <= "0" ;
      o_interrupt_mask(0 downto 0) <= "0" ;
      o_interrupt_mask(1 downto 1) <= "0" ;
      o_interrupt_mask(2 downto 2) <= "0" ;
      o_interrupt_mask(3 downto 3) <= "0" ;
      o_interrupt_mask(4 downto 4) <= "0" ;
      o_engine_sticky_status(0 downto 0) <= "0" ;
      o_engine_sticky_status(1 downto 1) <= "0" ;
      o_engine_sticky_status(2 downto 2) <= "0" ;
      o_engine_sticky_status(3 downto 3) <= "0" ;
      o_engine_sticky_status(4 downto 4) <= "0" ;
      o_engine_sticky_status(5 downto 5) <= "0" ;
      o_engine_sticky_status(6 downto 6) <= "0" ;
      o_engine_sticky_status(7 downto 7) <= "0" ;
      o_bimc_monitor_mask(0 downto 0) <= "0" ;
      o_bimc_monitor_mask(1 downto 1) <= "0" ;
      o_bimc_monitor_mask(2 downto 2) <= "0" ;
      o_bimc_monitor_mask(3 downto 3) <= "0" ;
      o_bimc_monitor_mask(4 downto 4) <= "0" ;
      o_bimc_monitor_mask(5 downto 5) <= "0" ;
      o_bimc_monitor_mask(6 downto 6) <= "0" ;
      o_bimc_ecc_uncorrectable_error_cnt <= "00000000000000000000000000000000" ;
      o_bimc_ecc_correctable_error_cnt <= "00000000000000000000000000000000" ;
      o_bimc_parity_error_cnt <= "00000000000000000000000000000000" ;
      o_bimc_global_config(0 downto 0) <= "1" ;
      o_bimc_global_config(1 downto 1) <= "0" ;
      o_bimc_global_config(2 downto 2) <= "0" ;
      o_bimc_global_config(3 downto 3) <= "0" ;
      o_bimc_global_config(4 downto 4) <= "0" ;
      o_bimc_global_config(5 downto 5) <= "0" ;
      o_bimc_global_config(31 downto 6) <= "00000000000000000000000000" ;
      o_bimc_eccpar_debug(11 downto 0) <= "000000000000" ;
      o_bimc_eccpar_debug(15 downto 12) <= "0000" ;
      o_bimc_eccpar_debug(17 downto 16) <= "00" ;
      o_bimc_eccpar_debug(19 downto 18) <= "00" ;
      o_bimc_eccpar_debug(21 downto 20) <= "00" ;
      o_bimc_eccpar_debug(22 downto 22) <= "0" ;
      o_bimc_eccpar_debug(23 downto 23) <= "0" ;
      o_bimc_eccpar_debug(27 downto 24) <= "0000" ;
      o_bimc_eccpar_debug(28 downto 28) <= "0" ;
      o_bimc_cmd2(7 downto 0) <= "00000000" ;
      o_bimc_cmd2(8 downto 8) <= "0" ;
      o_bimc_cmd2(9 downto 9) <= "0" ;
      o_bimc_cmd2(10 downto 10) <= "0" ;
      o_bimc_cmd1(15 downto 0) <= "0000000000000000" ;
      o_bimc_cmd1(27 downto 16) <= "000000000000" ;
      o_bimc_cmd1(31 downto 28) <= "0000" ;
      o_bimc_cmd0 <= "00000000000000000000000000000000" ;
      o_bimc_rxcmd2(7 downto 0) <= "00000000" ;
      o_bimc_rxcmd2(8 downto 8) <= "0" ;
      o_bimc_rxrsp2(7 downto 0) <= "00000000" ;
      o_bimc_rxrsp2(8 downto 8) <= "0" ;
      o_bimc_pollrsp2(7 downto 0) <= "00000000" ;
      o_bimc_pollrsp2(8 downto 8) <= "0" ;
      o_bimc_dbgcmd2(7 downto 0) <= "00000000" ;
      o_bimc_dbgcmd2(8 downto 8) <= "0" ;
      o_im_consumed(0 downto 0) <= "0" ;
      o_im_consumed(1 downto 1) <= "0" ;
      o_im_consumed(2 downto 2) <= "0" ;
      o_im_consumed(3 downto 3) <= "0" ;
      o_im_consumed(4 downto 4) <= "0" ;
      o_im_consumed(5 downto 5) <= "0" ;
      o_im_consumed(6 downto 6) <= "0" ;
      o_im_consumed(7 downto 7) <= "0" ;
      o_im_consumed(8 downto 8) <= "0" ;
      o_im_consumed(9 downto 9) <= "0" ;
      o_im_consumed(10 downto 10) <= "0" ;
      o_im_consumed(11 downto 11) <= "0" ;
      o_im_consumed(12 downto 12) <= "0" ;
      o_im_consumed(13 downto 13) <= "0" ;
      o_im_consumed(14 downto 14) <= "0" ;
      o_im_consumed(15 downto 15) <= "0" ;
      o_tready_override(0 downto 0) <= "0" ;
      o_tready_override(1 downto 1) <= "0" ;
      o_tready_override(2 downto 2) <= "0" ;
      o_tready_override(3 downto 3) <= "0" ;
      o_tready_override(4 downto 4) <= "0" ;
      o_tready_override(5 downto 5) <= "0" ;
      o_tready_override(6 downto 6) <= "0" ;
      o_tready_override(7 downto 7) <= "0" ;
      o_tready_override(8 downto 8) <= "0" ;
      o_regs_sa_ctrl(0 downto 0) <= "0" ;
      o_regs_sa_ctrl(1 downto 1) <= "0" ;
      o_regs_sa_ctrl(7 downto 2) <= "000000" ;
      o_regs_sa_ctrl(12 downto 8) <= "00000" ;
      o_regs_sa_ctrl(31 downto 13) <= "0000000000000000000" ;
      o_sa_snapshot_ia_wdata_part0(17 downto 0) <= "000000000000000000" ;
      o_sa_snapshot_ia_wdata_part0(31 downto 18) <= "00000000000000" ;
      o_sa_snapshot_ia_wdata_part1 <= "00000000000000000000000000000000" ;
      o_sa_snapshot_ia_config(4 downto 0) <= "00000" ;
      o_sa_snapshot_ia_config(8 downto 5) <= "0000" ;
      o_sa_count_ia_wdata_part0(17 downto 0) <= "000000000000000000" ;
      o_sa_count_ia_wdata_part0(31 downto 18) <= "00000000000000" ;
      o_sa_count_ia_wdata_part1 <= "00000000000000000000000000000000" ;
      o_sa_count_ia_config(4 downto 0) <= "00000" ;
      o_sa_count_ia_config(8 downto 5) <= "0000" ;
      o_cceip_encrypt_kop_fifo_override(0 downto 0) <= "0" ;
      o_cceip_encrypt_kop_fifo_override(1 downto 1) <= "0" ;
      o_cceip_encrypt_kop_fifo_override(2 downto 2) <= "0" ;
      o_cceip_encrypt_kop_fifo_override(3 downto 3) <= "0" ;
      o_cceip_encrypt_kop_fifo_override(4 downto 4) <= "0" ;
      o_cceip_encrypt_kop_fifo_override(5 downto 5) <= "0" ;
      o_cceip_encrypt_kop_fifo_override(6 downto 6) <= "0" ;
      o_cceip_validate_kop_fifo_override(0 downto 0) <= "0" ;
      o_cceip_validate_kop_fifo_override(1 downto 1) <= "0" ;
      o_cceip_validate_kop_fifo_override(2 downto 2) <= "0" ;
      o_cceip_validate_kop_fifo_override(3 downto 3) <= "0" ;
      o_cceip_validate_kop_fifo_override(4 downto 4) <= "0" ;
      o_cceip_validate_kop_fifo_override(5 downto 5) <= "0" ;
      o_cceip_validate_kop_fifo_override(6 downto 6) <= "0" ;
      o_cddip_decrypt_kop_fifo_override(0 downto 0) <= "0" ;
      o_cddip_decrypt_kop_fifo_override(1 downto 1) <= "0" ;
      o_cddip_decrypt_kop_fifo_override(2 downto 2) <= "0" ;
      o_cddip_decrypt_kop_fifo_override(3 downto 3) <= "0" ;
      o_cddip_decrypt_kop_fifo_override(4 downto 4) <= "0" ;
      o_cddip_decrypt_kop_fifo_override(5 downto 5) <= "0" ;
      o_cddip_decrypt_kop_fifo_override(6 downto 6) <= "0" ;
      o_sa_global_ctrl(0 downto 0) <= "0" ;
      o_sa_global_ctrl(1 downto 1) <= "0" ;
      o_sa_global_ctrl(31 downto 2) <= "000000000000000000000000000000" ;
      o_sa_ctrl_ia_wdata_part0(4 downto 0) <= "00000" ;
      o_sa_ctrl_ia_wdata_part0(31 downto 5) <= "000000000000000000000000000" ;
      o_sa_ctrl_ia_config(4 downto 0) <= "00000" ;
      o_sa_ctrl_ia_config(8 downto 5) <= "0000" ;
      o_kdf_test_key_size_config <= "00000000000000000000000000000000" ;
    elsif (clk'event and clk = '1') then
      if (i_sw_init = '1') then
        o_spare_config <= "00000000000000000000000000000000" ;
        o_cceip0_out_ia_wdata_part0(5 downto 0) <= "000000" ;
        o_cceip0_out_ia_wdata_part1 <= "00000000000000000000000000000000" ;
        o_cceip0_out_ia_wdata_part2 <= "00000000000000000000000000000000" ;
        o_cceip0_out_ia_config(8 downto 0) <= "000000000" ;
        o_cceip0_out_ia_config(12 downto 9) <= "0000" ;
        o_cceip0_out_im_config(9 downto 0) <= "1000000000" ;
        o_cceip0_out_im_config(11 downto 10) <= "11" ;
        o_cceip0_out_im_read_done(0 downto 0) <= "0" ;
        o_cceip0_out_im_read_done(1 downto 1) <= "0" ;
        o_cceip1_out_ia_wdata_part0(5 downto 0) <= "000000" ;
        o_cceip1_out_ia_wdata_part1 <= "00000000000000000000000000000000" ;
        o_cceip1_out_ia_wdata_part2 <= "00000000000000000000000000000000" ;
        o_cceip1_out_ia_config(8 downto 0) <= "000000000" ;
        o_cceip1_out_ia_config(12 downto 9) <= "0000" ;
        o_cceip1_out_im_config(9 downto 0) <= "1000000000" ;
        o_cceip1_out_im_config(11 downto 10) <= "11" ;
        o_cceip1_out_im_read_done(0 downto 0) <= "0" ;
        o_cceip1_out_im_read_done(1 downto 1) <= "0" ;
        o_cceip2_out_ia_wdata_part0(5 downto 0) <= "000000" ;
        o_cceip2_out_ia_wdata_part1 <= "00000000000000000000000000000000" ;
        o_cceip2_out_ia_wdata_part2 <= "00000000000000000000000000000000" ;
        o_cceip2_out_ia_config(8 downto 0) <= "000000000" ;
        o_cceip2_out_ia_config(12 downto 9) <= "0000" ;
        o_cceip2_out_im_config(9 downto 0) <= "1000000000" ;
        o_cceip2_out_im_config(11 downto 10) <= "11" ;
        o_cceip2_out_im_read_done(0 downto 0) <= "0" ;
        o_cceip2_out_im_read_done(1 downto 1) <= "0" ;
        o_cceip3_out_ia_wdata_part0(5 downto 0) <= "000000" ;
        o_cceip3_out_ia_wdata_part1 <= "00000000000000000000000000000000" ;
        o_cceip3_out_ia_wdata_part2 <= "00000000000000000000000000000000" ;
        o_cceip3_out_ia_config(8 downto 0) <= "000000000" ;
        o_cceip3_out_ia_config(12 downto 9) <= "0000" ;
        o_cceip3_out_im_config(9 downto 0) <= "1000000000" ;
        o_cceip3_out_im_config(11 downto 10) <= "11" ;
        o_cceip3_out_im_read_done(0 downto 0) <= "0" ;
        o_cceip3_out_im_read_done(1 downto 1) <= "0" ;
        o_cddip0_out_ia_wdata_part0(5 downto 0) <= "000000" ;
        o_cddip0_out_ia_wdata_part1 <= "00000000000000000000000000000000" ;
        o_cddip0_out_ia_wdata_part2 <= "00000000000000000000000000000000" ;
        o_cddip0_out_ia_config(8 downto 0) <= "000000000" ;
        o_cddip0_out_ia_config(12 downto 9) <= "0000" ;
        o_cddip0_out_im_config(9 downto 0) <= "1000000000" ;
        o_cddip0_out_im_config(11 downto 10) <= "11" ;
        o_cddip0_out_im_read_done(0 downto 0) <= "0" ;
        o_cddip0_out_im_read_done(1 downto 1) <= "0" ;
        o_cddip1_out_ia_wdata_part0(5 downto 0) <= "000000" ;
        o_cddip1_out_ia_wdata_part1 <= "00000000000000000000000000000000" ;
        o_cddip1_out_ia_wdata_part2 <= "00000000000000000000000000000000" ;
        o_cddip1_out_ia_config(8 downto 0) <= "000000000" ;
        o_cddip1_out_ia_config(12 downto 9) <= "0000" ;
        o_cddip1_out_im_config(9 downto 0) <= "1000000000" ;
        o_cddip1_out_im_config(11 downto 10) <= "11" ;
        o_cddip1_out_im_read_done(0 downto 0) <= "0" ;
        o_cddip1_out_im_read_done(1 downto 1) <= "0" ;
        o_cddip2_out_ia_wdata_part0(5 downto 0) <= "000000" ;
        o_cddip2_out_ia_wdata_part1 <= "00000000000000000000000000000000" ;
        o_cddip2_out_ia_wdata_part2 <= "00000000000000000000000000000000" ;
        o_cddip2_out_ia_config(8 downto 0) <= "000000000" ;
        o_cddip2_out_ia_config(12 downto 9) <= "0000" ;
        o_cddip2_out_im_config(9 downto 0) <= "1000000000" ;
        o_cddip2_out_im_config(11 downto 10) <= "11" ;
        o_cddip2_out_im_read_done(0 downto 0) <= "0" ;
        o_cddip2_out_im_read_done(1 downto 1) <= "0" ;
        o_cddip3_out_ia_wdata_part0(5 downto 0) <= "000000" ;
        o_cddip3_out_ia_wdata_part1 <= "00000000000000000000000000000000" ;
        o_cddip3_out_ia_wdata_part2 <= "00000000000000000000000000000000" ;
        o_cddip3_out_ia_config(8 downto 0) <= "000000000" ;
        o_cddip3_out_ia_config(12 downto 9) <= "0000" ;
        o_cddip3_out_im_config(9 downto 0) <= "1000000000" ;
        o_cddip3_out_im_config(11 downto 10) <= "11" ;
        o_cddip3_out_im_read_done(0 downto 0) <= "0" ;
        o_cddip3_out_im_read_done(1 downto 1) <= "0" ;
        o_ckv_ia_wdata_part0 <= "00000000000000000000000000000000" ;
        o_ckv_ia_wdata_part1 <= "00000000000000000000000000000000" ;
        o_ckv_ia_config(14 downto 0) <= "000000000000000" ;
        o_ckv_ia_config(18 downto 15) <= "0000" ;
        o_kim_ia_wdata_part0(14 downto 0) <= "000000000000000" ;
        o_kim_ia_wdata_part0(16 downto 15) <= "00" ;
        o_kim_ia_wdata_part0(19 downto 17) <= "000" ;
        o_kim_ia_wdata_part0(20 downto 20) <= "0" ;
        o_kim_ia_wdata_part1(0 downto 0) <= "0" ;
        o_kim_ia_wdata_part1(12 downto 1) <= "000000000000" ;
        o_kim_ia_wdata_part1(16 downto 13) <= "0000" ;
        o_kim_ia_config(13 downto 0) <= "00000000000000" ;
        o_kim_ia_config(17 downto 14) <= "0000" ;
        o_label0_config(7 downto 0) <= "00000000" ;
        o_label0_config(8 downto 8) <= "1" ;
        o_label0_config(14 downto 9) <= "000000" ;
        o_label0_config(15 downto 15) <= "0" ;
        o_label0_data7 <= "00000000000000000000000000000000" ;
        o_label0_data6 <= "00000000000000000000000000000000" ;
        o_label0_data5 <= "00000000000000000000000000000000" ;
        o_label0_data4 <= "00000000000000000000000000000000" ;
        o_label0_data3 <= "00000000000000000000000000000000" ;
        o_label0_data2 <= "00000000000000000000000000000000" ;
        o_label0_data1 <= "00000000000000000000000000000000" ;
        o_label0_data0 <= "00000000000000000000000000000000" ;
        o_label1_config(7 downto 0) <= "00000000" ;
        o_label1_config(8 downto 8) <= "1" ;
        o_label1_config(14 downto 9) <= "000000" ;
        o_label1_config(15 downto 15) <= "0" ;
        o_label1_data7 <= "00000000000000000000000000000000" ;
        o_label1_data6 <= "00000000000000000000000000000000" ;
        o_label1_data5 <= "00000000000000000000000000000000" ;
        o_label1_data4 <= "00000000000000000000000000000000" ;
        o_label1_data3 <= "00000000000000000000000000000000" ;
        o_label1_data2 <= "00000000000000000000000000000000" ;
        o_label1_data1 <= "00000000000000000000000000000000" ;
        o_label1_data0 <= "00000000000000000000000000000000" ;
        o_label2_config(7 downto 0) <= "00000000" ;
        o_label2_config(8 downto 8) <= "1" ;
        o_label2_config(14 downto 9) <= "000000" ;
        o_label2_config(15 downto 15) <= "0" ;
        o_label2_data7 <= "00000000000000000000000000000000" ;
        o_label2_data6 <= "00000000000000000000000000000000" ;
        o_label2_data5 <= "00000000000000000000000000000000" ;
        o_label2_data4 <= "00000000000000000000000000000000" ;
        o_label2_data3 <= "00000000000000000000000000000000" ;
        o_label2_data2 <= "00000000000000000000000000000000" ;
        o_label2_data1 <= "00000000000000000000000000000000" ;
        o_label2_data0 <= "00000000000000000000000000000000" ;
        o_label3_config(7 downto 0) <= "00000000" ;
        o_label3_config(8 downto 8) <= "1" ;
        o_label3_config(14 downto 9) <= "000000" ;
        o_label3_config(15 downto 15) <= "0" ;
        o_label3_data7 <= "00000000000000000000000000000000" ;
        o_label3_data6 <= "00000000000000000000000000000000" ;
        o_label3_data5 <= "00000000000000000000000000000000" ;
        o_label3_data4 <= "00000000000000000000000000000000" ;
        o_label3_data3 <= "00000000000000000000000000000000" ;
        o_label3_data2 <= "00000000000000000000000000000000" ;
        o_label3_data1 <= "00000000000000000000000000000000" ;
        o_label3_data0 <= "00000000000000000000000000000000" ;
        o_label4_config(7 downto 0) <= "00000000" ;
        o_label4_config(8 downto 8) <= "1" ;
        o_label4_config(14 downto 9) <= "000000" ;
        o_label4_config(15 downto 15) <= "0" ;
        o_label4_data7 <= "00000000000000000000000000000000" ;
        o_label4_data6 <= "00000000000000000000000000000000" ;
        o_label4_data5 <= "00000000000000000000000000000000" ;
        o_label4_data4 <= "00000000000000000000000000000000" ;
        o_label4_data3 <= "00000000000000000000000000000000" ;
        o_label4_data2 <= "00000000000000000000000000000000" ;
        o_label4_data1 <= "00000000000000000000000000000000" ;
        o_label4_data0 <= "00000000000000000000000000000000" ;
        o_label5_config(7 downto 0) <= "00000000" ;
        o_label5_config(8 downto 8) <= "1" ;
        o_label5_config(14 downto 9) <= "000000" ;
        o_label5_config(15 downto 15) <= "0" ;
        o_label5_data7 <= "00000000000000000000000000000000" ;
        o_label5_data6 <= "00000000000000000000000000000000" ;
        o_label5_data5 <= "00000000000000000000000000000000" ;
        o_label5_data4 <= "00000000000000000000000000000000" ;
        o_label5_data3 <= "00000000000000000000000000000000" ;
        o_label5_data2 <= "00000000000000000000000000000000" ;
        o_label5_data1 <= "00000000000000000000000000000000" ;
        o_label5_data0 <= "00000000000000000000000000000000" ;
        o_label6_config(7 downto 0) <= "00000000" ;
        o_label6_config(8 downto 8) <= "1" ;
        o_label6_config(14 downto 9) <= "000000" ;
        o_label6_config(15 downto 15) <= "0" ;
        o_label6_data7 <= "00000000000000000000000000000000" ;
        o_label6_data6 <= "00000000000000000000000000000000" ;
        o_label6_data5 <= "00000000000000000000000000000000" ;
        o_label6_data4 <= "00000000000000000000000000000000" ;
        o_label6_data3 <= "00000000000000000000000000000000" ;
        o_label6_data2 <= "00000000000000000000000000000000" ;
        o_label6_data1 <= "00000000000000000000000000000000" ;
        o_label6_data0 <= "00000000000000000000000000000000" ;
        o_label7_config(7 downto 0) <= "00000000" ;
        o_label7_config(8 downto 8) <= "1" ;
        o_label7_config(14 downto 9) <= "000000" ;
        o_label7_config(15 downto 15) <= "0" ;
        o_label7_data7 <= "00000000000000000000000000000000" ;
        o_label7_data6 <= "00000000000000000000000000000000" ;
        o_label7_data5 <= "00000000000000000000000000000000" ;
        o_label7_data4 <= "00000000000000000000000000000000" ;
        o_label7_data3 <= "00000000000000000000000000000000" ;
        o_label7_data2 <= "00000000000000000000000000000000" ;
        o_label7_data1 <= "00000000000000000000000000000000" ;
        o_label7_data0 <= "00000000000000000000000000000000" ;
        o_kdf_drbg_ctrl <= "00" ;
        o_kdf_drbg_seed_0_state_key_31_0 <= "00000000000000000000000000000000" ;
        o_kdf_drbg_seed_0_state_key_63_32 <= "00000000000000000000000000000000"
         ;
        o_kdf_drbg_seed_0_state_key_95_64 <= "00000000000000000000000000000000"
         ;
        o_kdf_drbg_seed_0_state_key_127_96 <= "00000000000000000000000000000000"
         ;
        o_kdf_drbg_seed_0_state_key_159_128 <=
         "00000000000000000000000000000000" ;
        o_kdf_drbg_seed_0_state_key_191_160 <=
         "00000000000000000000000000000000" ;
        o_kdf_drbg_seed_0_state_key_223_192 <=
         "00000000000000000000000000000000" ;
        o_kdf_drbg_seed_0_state_key_255_224 <=
         "00000000000000000000000000000000" ;
        o_kdf_drbg_seed_0_state_value_31_0 <= "00000000000000000000000000000000"
         ;
        o_kdf_drbg_seed_0_state_value_63_32 <=
         "00000000000000000000000000000000" ;
        o_kdf_drbg_seed_0_state_value_95_64 <=
         "00000000000000000000000000000000" ;
        o_kdf_drbg_seed_0_state_value_127_96 <=
         "00000000000000000000000000000000" ;
        o_kdf_drbg_seed_0_reseed_interval_0 <=
         "00000000000000000000000000000000" ;
        o_kdf_drbg_seed_0_reseed_interval_1 <= "0000000000000000" ;
        o_kdf_drbg_seed_1_state_key_31_0 <= "00000000000000000000000000000000" ;
        o_kdf_drbg_seed_1_state_key_63_32 <= "00000000000000000000000000000000"
         ;
        o_kdf_drbg_seed_1_state_key_95_64 <= "00000000000000000000000000000000"
         ;
        o_kdf_drbg_seed_1_state_key_127_96 <= "00000000000000000000000000000000"
         ;
        o_kdf_drbg_seed_1_state_key_159_128 <=
         "00000000000000000000000000000000" ;
        o_kdf_drbg_seed_1_state_key_191_160 <=
         "00000000000000000000000000000000" ;
        o_kdf_drbg_seed_1_state_key_223_192 <=
         "00000000000000000000000000000000" ;
        o_kdf_drbg_seed_1_state_key_255_224 <=
         "00000000000000000000000000000000" ;
        o_kdf_drbg_seed_1_state_value_31_0 <= "00000000000000000000000000000000"
         ;
        o_kdf_drbg_seed_1_state_value_63_32 <=
         "00000000000000000000000000000000" ;
        o_kdf_drbg_seed_1_state_value_95_64 <=
         "00000000000000000000000000000000" ;
        o_kdf_drbg_seed_1_state_value_127_96 <=
         "00000000000000000000000000000000" ;
        o_kdf_drbg_seed_1_reseed_interval_0 <=
         "00000000000000000000000000000000" ;
        o_kdf_drbg_seed_1_reseed_interval_1 <= "0000000000000000" ;
        o_interrupt_status(0 downto 0) <= "0" ;
        o_interrupt_status(1 downto 1) <= "0" ;
        o_interrupt_status(2 downto 2) <= "0" ;
        o_interrupt_status(3 downto 3) <= "0" ;
        o_interrupt_status(4 downto 4) <= "0" ;
        o_interrupt_mask(0 downto 0) <= "0" ;
        o_interrupt_mask(1 downto 1) <= "0" ;
        o_interrupt_mask(2 downto 2) <= "0" ;
        o_interrupt_mask(3 downto 3) <= "0" ;
        o_interrupt_mask(4 downto 4) <= "0" ;
        o_engine_sticky_status(0 downto 0) <= "0" ;
        o_engine_sticky_status(1 downto 1) <= "0" ;
        o_engine_sticky_status(2 downto 2) <= "0" ;
        o_engine_sticky_status(3 downto 3) <= "0" ;
        o_engine_sticky_status(4 downto 4) <= "0" ;
        o_engine_sticky_status(5 downto 5) <= "0" ;
        o_engine_sticky_status(6 downto 6) <= "0" ;
        o_engine_sticky_status(7 downto 7) <= "0" ;
        o_bimc_monitor_mask(0 downto 0) <= "0" ;
        o_bimc_monitor_mask(1 downto 1) <= "0" ;
        o_bimc_monitor_mask(2 downto 2) <= "0" ;
        o_bimc_monitor_mask(3 downto 3) <= "0" ;
        o_bimc_monitor_mask(4 downto 4) <= "0" ;
        o_bimc_monitor_mask(5 downto 5) <= "0" ;
        o_bimc_monitor_mask(6 downto 6) <= "0" ;
        o_bimc_ecc_uncorrectable_error_cnt <= "00000000000000000000000000000000"
         ;
        o_bimc_ecc_correctable_error_cnt <= "00000000000000000000000000000000" ;
        o_bimc_parity_error_cnt <= "00000000000000000000000000000000" ;
        o_bimc_global_config(0 downto 0) <= "1" ;
        o_bimc_global_config(1 downto 1) <= "0" ;
        o_bimc_global_config(2 downto 2) <= "0" ;
        o_bimc_global_config(3 downto 3) <= "0" ;
        o_bimc_global_config(4 downto 4) <= "0" ;
        o_bimc_global_config(5 downto 5) <= "0" ;
        o_bimc_global_config(31 downto 6) <= "00000000000000000000000000" ;
        o_bimc_eccpar_debug(11 downto 0) <= "000000000000" ;
        o_bimc_eccpar_debug(15 downto 12) <= "0000" ;
        o_bimc_eccpar_debug(17 downto 16) <= "00" ;
        o_bimc_eccpar_debug(19 downto 18) <= "00" ;
        o_bimc_eccpar_debug(21 downto 20) <= "00" ;
        o_bimc_eccpar_debug(22 downto 22) <= "0" ;
        o_bimc_eccpar_debug(23 downto 23) <= "0" ;
        o_bimc_eccpar_debug(27 downto 24) <= "0000" ;
        o_bimc_eccpar_debug(28 downto 28) <= "0" ;
        o_bimc_cmd2(7 downto 0) <= "00000000" ;
        o_bimc_cmd2(8 downto 8) <= "0" ;
        o_bimc_cmd2(9 downto 9) <= "0" ;
        o_bimc_cmd2(10 downto 10) <= "0" ;
        o_bimc_cmd1(15 downto 0) <= "0000000000000000" ;
        o_bimc_cmd1(27 downto 16) <= "000000000000" ;
        o_bimc_cmd1(31 downto 28) <= "0000" ;
        o_bimc_cmd0 <= "00000000000000000000000000000000" ;
        o_bimc_rxcmd2(7 downto 0) <= "00000000" ;
        o_bimc_rxcmd2(8 downto 8) <= "0" ;
        o_bimc_rxrsp2(7 downto 0) <= "00000000" ;
        o_bimc_rxrsp2(8 downto 8) <= "0" ;
        o_bimc_pollrsp2(7 downto 0) <= "00000000" ;
        o_bimc_pollrsp2(8 downto 8) <= "0" ;
        o_bimc_dbgcmd2(7 downto 0) <= "00000000" ;
        o_bimc_dbgcmd2(8 downto 8) <= "0" ;
        o_im_consumed(0 downto 0) <= "0" ;
        o_im_consumed(1 downto 1) <= "0" ;
        o_im_consumed(2 downto 2) <= "0" ;
        o_im_consumed(3 downto 3) <= "0" ;
        o_im_consumed(4 downto 4) <= "0" ;
        o_im_consumed(5 downto 5) <= "0" ;
        o_im_consumed(6 downto 6) <= "0" ;
        o_im_consumed(7 downto 7) <= "0" ;
        o_im_consumed(8 downto 8) <= "0" ;
        o_im_consumed(9 downto 9) <= "0" ;
        o_im_consumed(10 downto 10) <= "0" ;
        o_im_consumed(11 downto 11) <= "0" ;
        o_im_consumed(12 downto 12) <= "0" ;
        o_im_consumed(13 downto 13) <= "0" ;
        o_im_consumed(14 downto 14) <= "0" ;
        o_im_consumed(15 downto 15) <= "0" ;
        o_tready_override(0 downto 0) <= "0" ;
        o_tready_override(1 downto 1) <= "0" ;
        o_tready_override(2 downto 2) <= "0" ;
        o_tready_override(3 downto 3) <= "0" ;
        o_tready_override(4 downto 4) <= "0" ;
        o_tready_override(5 downto 5) <= "0" ;
        o_tready_override(6 downto 6) <= "0" ;
        o_tready_override(7 downto 7) <= "0" ;
        o_tready_override(8 downto 8) <= "0" ;
        o_regs_sa_ctrl(0 downto 0) <= "0" ;
        o_regs_sa_ctrl(1 downto 1) <= "0" ;
        o_regs_sa_ctrl(7 downto 2) <= "000000" ;
        o_regs_sa_ctrl(12 downto 8) <= "00000" ;
        o_regs_sa_ctrl(31 downto 13) <= "0000000000000000000" ;
        o_sa_snapshot_ia_wdata_part0(17 downto 0) <= "000000000000000000" ;
        o_sa_snapshot_ia_wdata_part0(31 downto 18) <= "00000000000000" ;
        o_sa_snapshot_ia_wdata_part1 <= "00000000000000000000000000000000" ;
        o_sa_snapshot_ia_config(4 downto 0) <= "00000" ;
        o_sa_snapshot_ia_config(8 downto 5) <= "0000" ;
        o_sa_count_ia_wdata_part0(17 downto 0) <= "000000000000000000" ;
        o_sa_count_ia_wdata_part0(31 downto 18) <= "00000000000000" ;
        o_sa_count_ia_wdata_part1 <= "00000000000000000000000000000000" ;
        o_sa_count_ia_config(4 downto 0) <= "00000" ;
        o_sa_count_ia_config(8 downto 5) <= "0000" ;
        o_cceip_encrypt_kop_fifo_override(0 downto 0) <= "0" ;
        o_cceip_encrypt_kop_fifo_override(1 downto 1) <= "0" ;
        o_cceip_encrypt_kop_fifo_override(2 downto 2) <= "0" ;
        o_cceip_encrypt_kop_fifo_override(3 downto 3) <= "0" ;
        o_cceip_encrypt_kop_fifo_override(4 downto 4) <= "0" ;
        o_cceip_encrypt_kop_fifo_override(5 downto 5) <= "0" ;
        o_cceip_encrypt_kop_fifo_override(6 downto 6) <= "0" ;
        o_cceip_validate_kop_fifo_override(0 downto 0) <= "0" ;
        o_cceip_validate_kop_fifo_override(1 downto 1) <= "0" ;
        o_cceip_validate_kop_fifo_override(2 downto 2) <= "0" ;
        o_cceip_validate_kop_fifo_override(3 downto 3) <= "0" ;
        o_cceip_validate_kop_fifo_override(4 downto 4) <= "0" ;
        o_cceip_validate_kop_fifo_override(5 downto 5) <= "0" ;
        o_cceip_validate_kop_fifo_override(6 downto 6) <= "0" ;
        o_cddip_decrypt_kop_fifo_override(0 downto 0) <= "0" ;
        o_cddip_decrypt_kop_fifo_override(1 downto 1) <= "0" ;
        o_cddip_decrypt_kop_fifo_override(2 downto 2) <= "0" ;
        o_cddip_decrypt_kop_fifo_override(3 downto 3) <= "0" ;
        o_cddip_decrypt_kop_fifo_override(4 downto 4) <= "0" ;
        o_cddip_decrypt_kop_fifo_override(5 downto 5) <= "0" ;
        o_cddip_decrypt_kop_fifo_override(6 downto 6) <= "0" ;
        o_sa_global_ctrl(0 downto 0) <= "0" ;
        o_sa_global_ctrl(1 downto 1) <= "0" ;
        o_sa_global_ctrl(31 downto 2) <= "000000000000000000000000000000" ;
        o_sa_ctrl_ia_wdata_part0(4 downto 0) <= "00000" ;
        o_sa_ctrl_ia_wdata_part0(31 downto 5) <= "000000000000000000000000000" ;
        o_sa_ctrl_ia_config(4 downto 0) <= "00000" ;
        o_sa_ctrl_ia_config(8 downto 5) <= "0000" ;
        o_kdf_test_key_size_config <= "00000000000000000000000000000000" ;
      else
        if (w_load_spare_config = '1') then
          o_spare_config <= f32_data ;
        end if;
        if (w_load_cceip0_out_ia_wdata_part0 = '1') then
          o_cceip0_out_ia_wdata_part0(5 downto 0) <= f32_data(5 downto 0) ;
        end if;
        if (w_load_cceip0_out_ia_wdata_part1 = '1') then
          o_cceip0_out_ia_wdata_part1 <= f32_data ;
        end if;
        if (w_load_cceip0_out_ia_wdata_part2 = '1') then
          o_cceip0_out_ia_wdata_part2 <= f32_data ;
        end if;
        if (w_load_cceip0_out_ia_config = '1') then
          o_cceip0_out_ia_config(8 downto 0) <= f32_data(8 downto 0) ;
        end if;
        if (w_load_cceip0_out_ia_config = '1') then
          o_cceip0_out_ia_config(12 downto 9) <= f32_data(31 downto 28) ;
        end if;
        if (w_load_cceip0_out_im_config = '1') then
          o_cceip0_out_im_config(9 downto 0) <= f32_data(9 downto 0) ;
        end if;
        if (w_load_cceip0_out_im_config = '1') then
          o_cceip0_out_im_config(11 downto 10) <= f32_data(31 downto 30) ;
        end if;
        if (w_load_cceip0_out_im_read_done = '1') then
          o_cceip0_out_im_read_done(0 downto 0) <= f32_data(30 downto 30) ;
        end if;
        if (w_load_cceip0_out_im_read_done = '1') then
          o_cceip0_out_im_read_done(1 downto 1) <= f32_data(31 downto 31) ;
        end if;
        if (w_load_cceip1_out_ia_wdata_part0 = '1') then
          o_cceip1_out_ia_wdata_part0(5 downto 0) <= f32_data(5 downto 0) ;
        end if;
        if (w_load_cceip1_out_ia_wdata_part1 = '1') then
          o_cceip1_out_ia_wdata_part1 <= f32_data ;
        end if;
        if (w_load_cceip1_out_ia_wdata_part2 = '1') then
          o_cceip1_out_ia_wdata_part2 <= f32_data ;
        end if;
        if (w_load_cceip1_out_ia_config = '1') then
          o_cceip1_out_ia_config(8 downto 0) <= f32_data(8 downto 0) ;
        end if;
        if (w_load_cceip1_out_ia_config = '1') then
          o_cceip1_out_ia_config(12 downto 9) <= f32_data(31 downto 28) ;
        end if;
        if (w_load_cceip1_out_im_config = '1') then
          o_cceip1_out_im_config(9 downto 0) <= f32_data(9 downto 0) ;
        end if;
        if (w_load_cceip1_out_im_config = '1') then
          o_cceip1_out_im_config(11 downto 10) <= f32_data(31 downto 30) ;
        end if;
        if (w_load_cceip1_out_im_read_done = '1') then
          o_cceip1_out_im_read_done(0 downto 0) <= f32_data(30 downto 30) ;
        end if;
        if (w_load_cceip1_out_im_read_done = '1') then
          o_cceip1_out_im_read_done(1 downto 1) <= f32_data(31 downto 31) ;
        end if;
        if (w_load_cceip2_out_ia_wdata_part0 = '1') then
          o_cceip2_out_ia_wdata_part0(5 downto 0) <= f32_data(5 downto 0) ;
        end if;
        if (w_load_cceip2_out_ia_wdata_part1 = '1') then
          o_cceip2_out_ia_wdata_part1 <= f32_data ;
        end if;
        if (w_load_cceip2_out_ia_wdata_part2 = '1') then
          o_cceip2_out_ia_wdata_part2 <= f32_data ;
        end if;
        if (w_load_cceip2_out_ia_config = '1') then
          o_cceip2_out_ia_config(8 downto 0) <= f32_data(8 downto 0) ;
        end if;
        if (w_load_cceip2_out_ia_config = '1') then
          o_cceip2_out_ia_config(12 downto 9) <= f32_data(31 downto 28) ;
        end if;
        if (w_load_cceip2_out_im_config = '1') then
          o_cceip2_out_im_config(9 downto 0) <= f32_data(9 downto 0) ;
        end if;
        if (w_load_cceip2_out_im_config = '1') then
          o_cceip2_out_im_config(11 downto 10) <= f32_data(31 downto 30) ;
        end if;
        if (w_load_cceip2_out_im_read_done = '1') then
          o_cceip2_out_im_read_done(0 downto 0) <= f32_data(30 downto 30) ;
        end if;
        if (w_load_cceip2_out_im_read_done = '1') then
          o_cceip2_out_im_read_done(1 downto 1) <= f32_data(31 downto 31) ;
        end if;
        if (w_load_cceip3_out_ia_wdata_part0 = '1') then
          o_cceip3_out_ia_wdata_part0(5 downto 0) <= f32_data(5 downto 0) ;
        end if;
        if (w_load_cceip3_out_ia_wdata_part1 = '1') then
          o_cceip3_out_ia_wdata_part1 <= f32_data ;
        end if;
        if (w_load_cceip3_out_ia_wdata_part2 = '1') then
          o_cceip3_out_ia_wdata_part2 <= f32_data ;
        end if;
        if (w_load_cceip3_out_ia_config = '1') then
          o_cceip3_out_ia_config(8 downto 0) <= f32_data(8 downto 0) ;
        end if;
        if (w_load_cceip3_out_ia_config = '1') then
          o_cceip3_out_ia_config(12 downto 9) <= f32_data(31 downto 28) ;
        end if;
        if (w_load_cceip3_out_im_config = '1') then
          o_cceip3_out_im_config(9 downto 0) <= f32_data(9 downto 0) ;
        end if;
        if (w_load_cceip3_out_im_config = '1') then
          o_cceip3_out_im_config(11 downto 10) <= f32_data(31 downto 30) ;
        end if;
        if (w_load_cceip3_out_im_read_done = '1') then
          o_cceip3_out_im_read_done(0 downto 0) <= f32_data(30 downto 30) ;
        end if;
        if (w_load_cceip3_out_im_read_done = '1') then
          o_cceip3_out_im_read_done(1 downto 1) <= f32_data(31 downto 31) ;
        end if;
        if (w_load_cddip0_out_ia_wdata_part0 = '1') then
          o_cddip0_out_ia_wdata_part0(5 downto 0) <= f32_data(5 downto 0) ;
        end if;
        if (w_load_cddip0_out_ia_wdata_part1 = '1') then
          o_cddip0_out_ia_wdata_part1 <= f32_data ;
        end if;
        if (w_load_cddip0_out_ia_wdata_part2 = '1') then
          o_cddip0_out_ia_wdata_part2 <= f32_data ;
        end if;
        if (w_load_cddip0_out_ia_config = '1') then
          o_cddip0_out_ia_config(8 downto 0) <= f32_data(8 downto 0) ;
        end if;
        if (w_load_cddip0_out_ia_config = '1') then
          o_cddip0_out_ia_config(12 downto 9) <= f32_data(31 downto 28) ;
        end if;
        if (w_load_cddip0_out_im_config = '1') then
          o_cddip0_out_im_config(9 downto 0) <= f32_data(9 downto 0) ;
        end if;
        if (w_load_cddip0_out_im_config = '1') then
          o_cddip0_out_im_config(11 downto 10) <= f32_data(31 downto 30) ;
        end if;
        if (w_load_cddip0_out_im_read_done = '1') then
          o_cddip0_out_im_read_done(0 downto 0) <= f32_data(30 downto 30) ;
        end if;
        if (w_load_cddip0_out_im_read_done = '1') then
          o_cddip0_out_im_read_done(1 downto 1) <= f32_data(31 downto 31) ;
        end if;
        if (w_load_cddip1_out_ia_wdata_part0 = '1') then
          o_cddip1_out_ia_wdata_part0(5 downto 0) <= f32_data(5 downto 0) ;
        end if;
        if (w_load_cddip1_out_ia_wdata_part1 = '1') then
          o_cddip1_out_ia_wdata_part1 <= f32_data ;
        end if;
        if (w_load_cddip1_out_ia_wdata_part2 = '1') then
          o_cddip1_out_ia_wdata_part2 <= f32_data ;
        end if;
        if (w_load_cddip1_out_ia_config = '1') then
          o_cddip1_out_ia_config(8 downto 0) <= f32_data(8 downto 0) ;
        end if;
        if (w_load_cddip1_out_ia_config = '1') then
          o_cddip1_out_ia_config(12 downto 9) <= f32_data(31 downto 28) ;
        end if;
        if (w_load_cddip1_out_im_config = '1') then
          o_cddip1_out_im_config(9 downto 0) <= f32_data(9 downto 0) ;
        end if;
        if (w_load_cddip1_out_im_config = '1') then
          o_cddip1_out_im_config(11 downto 10) <= f32_data(31 downto 30) ;
        end if;
        if (w_load_cddip1_out_im_read_done = '1') then
          o_cddip1_out_im_read_done(0 downto 0) <= f32_data(30 downto 30) ;
        end if;
        if (w_load_cddip1_out_im_read_done = '1') then
          o_cddip1_out_im_read_done(1 downto 1) <= f32_data(31 downto 31) ;
        end if;
        if (w_load_cddip2_out_ia_wdata_part0 = '1') then
          o_cddip2_out_ia_wdata_part0(5 downto 0) <= f32_data(5 downto 0) ;
        end if;
        if (w_load_cddip2_out_ia_wdata_part1 = '1') then
          o_cddip2_out_ia_wdata_part1 <= f32_data ;
        end if;
        if (w_load_cddip2_out_ia_wdata_part2 = '1') then
          o_cddip2_out_ia_wdata_part2 <= f32_data ;
        end if;
        if (w_load_cddip2_out_ia_config = '1') then
          o_cddip2_out_ia_config(8 downto 0) <= f32_data(8 downto 0) ;
        end if;
        if (w_load_cddip2_out_ia_config = '1') then
          o_cddip2_out_ia_config(12 downto 9) <= f32_data(31 downto 28) ;
        end if;
        if (w_load_cddip2_out_im_config = '1') then
          o_cddip2_out_im_config(9 downto 0) <= f32_data(9 downto 0) ;
        end if;
        if (w_load_cddip2_out_im_config = '1') then
          o_cddip2_out_im_config(11 downto 10) <= f32_data(31 downto 30) ;
        end if;
        if (w_load_cddip2_out_im_read_done = '1') then
          o_cddip2_out_im_read_done(0 downto 0) <= f32_data(30 downto 30) ;
        end if;
        if (w_load_cddip2_out_im_read_done = '1') then
          o_cddip2_out_im_read_done(1 downto 1) <= f32_data(31 downto 31) ;
        end if;
        if (w_load_cddip3_out_ia_wdata_part0 = '1') then
          o_cddip3_out_ia_wdata_part0(5 downto 0) <= f32_data(5 downto 0) ;
        end if;
        if (w_load_cddip3_out_ia_wdata_part1 = '1') then
          o_cddip3_out_ia_wdata_part1 <= f32_data ;
        end if;
        if (w_load_cddip3_out_ia_wdata_part2 = '1') then
          o_cddip3_out_ia_wdata_part2 <= f32_data ;
        end if;
        if (w_load_cddip3_out_ia_config = '1') then
          o_cddip3_out_ia_config(8 downto 0) <= f32_data(8 downto 0) ;
        end if;
        if (w_load_cddip3_out_ia_config = '1') then
          o_cddip3_out_ia_config(12 downto 9) <= f32_data(31 downto 28) ;
        end if;
        if (w_load_cddip3_out_im_config = '1') then
          o_cddip3_out_im_config(9 downto 0) <= f32_data(9 downto 0) ;
        end if;
        if (w_load_cddip3_out_im_config = '1') then
          o_cddip3_out_im_config(11 downto 10) <= f32_data(31 downto 30) ;
        end if;
        if (w_load_cddip3_out_im_read_done = '1') then
          o_cddip3_out_im_read_done(0 downto 0) <= f32_data(30 downto 30) ;
        end if;
        if (w_load_cddip3_out_im_read_done = '1') then
          o_cddip3_out_im_read_done(1 downto 1) <= f32_data(31 downto 31) ;
        end if;
        if (w_load_ckv_ia_wdata_part0 = '1') then
          o_ckv_ia_wdata_part0 <= f32_data ;
        end if;
        if (w_load_ckv_ia_wdata_part1 = '1') then
          o_ckv_ia_wdata_part1 <= f32_data ;
        end if;
        if (w_load_ckv_ia_config = '1') then
          o_ckv_ia_config(14 downto 0) <= f32_data(14 downto 0) ;
        end if;
        if (w_load_ckv_ia_config = '1') then
          o_ckv_ia_config(18 downto 15) <= f32_data(31 downto 28) ;
        end if;
        if (w_load_kim_ia_wdata_part0 = '1') then
          o_kim_ia_wdata_part0(14 downto 0) <= f32_data(14 downto 0) ;
        end if;
        if (w_load_kim_ia_wdata_part0 = '1') then
          o_kim_ia_wdata_part0(16 downto 15) <= f32_data(27 downto 26) ;
        end if;
        if (w_load_kim_ia_wdata_part0 = '1') then
          o_kim_ia_wdata_part0(19 downto 17) <= f32_data(30 downto 28) ;
        end if;
        if (w_load_kim_ia_wdata_part0 = '1') then
          o_kim_ia_wdata_part0(20 downto 20) <= f32_data(31 downto 31) ;
        end if;
        if (w_load_kim_ia_wdata_part1 = '1') then
          o_kim_ia_wdata_part1(0 downto 0) <= f32_data(0 downto 0) ;
        end if;
        if (w_load_kim_ia_wdata_part1 = '1') then
          o_kim_ia_wdata_part1(12 downto 1) <= f32_data(12 downto 1) ;
        end if;
        if (w_load_kim_ia_wdata_part1 = '1') then
          o_kim_ia_wdata_part1(16 downto 13) <= f32_data(31 downto 28) ;
        end if;
        if (w_load_kim_ia_config = '1') then
          o_kim_ia_config(13 downto 0) <= f32_data(13 downto 0) ;
        end if;
        if (w_load_kim_ia_config = '1') then
          o_kim_ia_config(17 downto 14) <= f32_data(31 downto 28) ;
        end if;
        if (w_load_label0_config = '1') then
          o_label0_config(7 downto 0) <= f32_data(7 downto 0) ;
        end if;
        if (w_load_label0_config = '1') then
          o_label0_config(8 downto 8) <= f32_data(8 downto 8) ;
        end if;
        if (w_load_label0_config = '1') then
          o_label0_config(14 downto 9) <= f32_data(30 downto 25) ;
        end if;
        if (w_load_label0_config = '1') then
          o_label0_config(15 downto 15) <= f32_data(31 downto 31) ;
        end if;
        if (w_load_label0_data7 = '1') then
          o_label0_data7 <= f32_data ;
        end if;
        if (w_load_label0_data6 = '1') then
          o_label0_data6 <= f32_data ;
        end if;
        if (w_load_label0_data5 = '1') then
          o_label0_data5 <= f32_data ;
        end if;
        if (w_load_label0_data4 = '1') then
          o_label0_data4 <= f32_data ;
        end if;
        if (w_load_label0_data3 = '1') then
          o_label0_data3 <= f32_data ;
        end if;
        if (w_load_label0_data2 = '1') then
          o_label0_data2 <= f32_data ;
        end if;
        if (w_load_label0_data1 = '1') then
          o_label0_data1 <= f32_data ;
        end if;
        if (w_load_label0_data0 = '1') then
          o_label0_data0 <= f32_data ;
        end if;
        if (w_load_label1_config = '1') then
          o_label1_config(7 downto 0) <= f32_data(7 downto 0) ;
        end if;
        if (w_load_label1_config = '1') then
          o_label1_config(8 downto 8) <= f32_data(8 downto 8) ;
        end if;
        if (w_load_label1_config = '1') then
          o_label1_config(14 downto 9) <= f32_data(30 downto 25) ;
        end if;
        if (w_load_label1_config = '1') then
          o_label1_config(15 downto 15) <= f32_data(31 downto 31) ;
        end if;
        if (w_load_label1_data7 = '1') then
          o_label1_data7 <= f32_data ;
        end if;
        if (w_load_label1_data6 = '1') then
          o_label1_data6 <= f32_data ;
        end if;
        if (w_load_label1_data5 = '1') then
          o_label1_data5 <= f32_data ;
        end if;
        if (w_load_label1_data4 = '1') then
          o_label1_data4 <= f32_data ;
        end if;
        if (w_load_label1_data3 = '1') then
          o_label1_data3 <= f32_data ;
        end if;
        if (w_load_label1_data2 = '1') then
          o_label1_data2 <= f32_data ;
        end if;
        if (w_load_label1_data1 = '1') then
          o_label1_data1 <= f32_data ;
        end if;
        if (w_load_label1_data0 = '1') then
          o_label1_data0 <= f32_data ;
        end if;
        if (w_load_label2_config = '1') then
          o_label2_config(7 downto 0) <= f32_data(7 downto 0) ;
        end if;
        if (w_load_label2_config = '1') then
          o_label2_config(8 downto 8) <= f32_data(8 downto 8) ;
        end if;
        if (w_load_label2_config = '1') then
          o_label2_config(14 downto 9) <= f32_data(30 downto 25) ;
        end if;
        if (w_load_label2_config = '1') then
          o_label2_config(15 downto 15) <= f32_data(31 downto 31) ;
        end if;
        if (w_load_label2_data7 = '1') then
          o_label2_data7 <= f32_data ;
        end if;
        if (w_load_label2_data6 = '1') then
          o_label2_data6 <= f32_data ;
        end if;
        if (w_load_label2_data5 = '1') then
          o_label2_data5 <= f32_data ;
        end if;
        if (w_load_label2_data4 = '1') then
          o_label2_data4 <= f32_data ;
        end if;
        if (w_load_label2_data3 = '1') then
          o_label2_data3 <= f32_data ;
        end if;
        if (w_load_label2_data2 = '1') then
          o_label2_data2 <= f32_data ;
        end if;
        if (w_load_label2_data1 = '1') then
          o_label2_data1 <= f32_data ;
        end if;
        if (w_load_label2_data0 = '1') then
          o_label2_data0 <= f32_data ;
        end if;
        if (w_load_label3_config = '1') then
          o_label3_config(7 downto 0) <= f32_data(7 downto 0) ;
        end if;
        if (w_load_label3_config = '1') then
          o_label3_config(8 downto 8) <= f32_data(8 downto 8) ;
        end if;
        if (w_load_label3_config = '1') then
          o_label3_config(14 downto 9) <= f32_data(30 downto 25) ;
        end if;
        if (w_load_label3_config = '1') then
          o_label3_config(15 downto 15) <= f32_data(31 downto 31) ;
        end if;
        if (w_load_label3_data7 = '1') then
          o_label3_data7 <= f32_data ;
        end if;
        if (w_load_label3_data6 = '1') then
          o_label3_data6 <= f32_data ;
        end if;
        if (w_load_label3_data5 = '1') then
          o_label3_data5 <= f32_data ;
        end if;
        if (w_load_label3_data4 = '1') then
          o_label3_data4 <= f32_data ;
        end if;
        if (w_load_label3_data3 = '1') then
          o_label3_data3 <= f32_data ;
        end if;
        if (w_load_label3_data2 = '1') then
          o_label3_data2 <= f32_data ;
        end if;
        if (w_load_label3_data1 = '1') then
          o_label3_data1 <= f32_data ;
        end if;
        if (w_load_label3_data0 = '1') then
          o_label3_data0 <= f32_data ;
        end if;
        if (w_load_label4_config = '1') then
          o_label4_config(7 downto 0) <= f32_data(7 downto 0) ;
        end if;
        if (w_load_label4_config = '1') then
          o_label4_config(8 downto 8) <= f32_data(8 downto 8) ;
        end if;
        if (w_load_label4_config = '1') then
          o_label4_config(14 downto 9) <= f32_data(30 downto 25) ;
        end if;
        if (w_load_label4_config = '1') then
          o_label4_config(15 downto 15) <= f32_data(31 downto 31) ;
        end if;
        if (w_load_label4_data7 = '1') then
          o_label4_data7 <= f32_data ;
        end if;
        if (w_load_label4_data6 = '1') then
          o_label4_data6 <= f32_data ;
        end if;
        if (w_load_label4_data5 = '1') then
          o_label4_data5 <= f32_data ;
        end if;
        if (w_load_label4_data4 = '1') then
          o_label4_data4 <= f32_data ;
        end if;
        if (w_load_label4_data3 = '1') then
          o_label4_data3 <= f32_data ;
        end if;
        if (w_load_label4_data2 = '1') then
          o_label4_data2 <= f32_data ;
        end if;
        if (w_load_label4_data1 = '1') then
          o_label4_data1 <= f32_data ;
        end if;
        if (w_load_label4_data0 = '1') then
          o_label4_data0 <= f32_data ;
        end if;
        if (w_load_label5_config = '1') then
          o_label5_config(7 downto 0) <= f32_data(7 downto 0) ;
        end if;
        if (w_load_label5_config = '1') then
          o_label5_config(8 downto 8) <= f32_data(8 downto 8) ;
        end if;
        if (w_load_label5_config = '1') then
          o_label5_config(14 downto 9) <= f32_data(30 downto 25) ;
        end if;
        if (w_load_label5_config = '1') then
          o_label5_config(15 downto 15) <= f32_data(31 downto 31) ;
        end if;
        if (w_load_label5_data7 = '1') then
          o_label5_data7 <= f32_data ;
        end if;
        if (w_load_label5_data6 = '1') then
          o_label5_data6 <= f32_data ;
        end if;
        if (w_load_label5_data5 = '1') then
          o_label5_data5 <= f32_data ;
        end if;
        if (w_load_label5_data4 = '1') then
          o_label5_data4 <= f32_data ;
        end if;
        if (w_load_label5_data3 = '1') then
          o_label5_data3 <= f32_data ;
        end if;
        if (w_load_label5_data2 = '1') then
          o_label5_data2 <= f32_data ;
        end if;
        if (w_load_label5_data1 = '1') then
          o_label5_data1 <= f32_data ;
        end if;
        if (w_load_label5_data0 = '1') then
          o_label5_data0 <= f32_data ;
        end if;
        if (w_load_label6_config = '1') then
          o_label6_config(7 downto 0) <= f32_data(7 downto 0) ;
        end if;
        if (w_load_label6_config = '1') then
          o_label6_config(8 downto 8) <= f32_data(8 downto 8) ;
        end if;
        if (w_load_label6_config = '1') then
          o_label6_config(14 downto 9) <= f32_data(30 downto 25) ;
        end if;
        if (w_load_label6_config = '1') then
          o_label6_config(15 downto 15) <= f32_data(31 downto 31) ;
        end if;
        if (w_load_label6_data7 = '1') then
          o_label6_data7 <= f32_data ;
        end if;
        if (w_load_label6_data6 = '1') then
          o_label6_data6 <= f32_data ;
        end if;
        if (w_load_label6_data5 = '1') then
          o_label6_data5 <= f32_data ;
        end if;
        if (w_load_label6_data4 = '1') then
          o_label6_data4 <= f32_data ;
        end if;
        if (w_load_label6_data3 = '1') then
          o_label6_data3 <= f32_data ;
        end if;
        if (w_load_label6_data2 = '1') then
          o_label6_data2 <= f32_data ;
        end if;
        if (w_load_label6_data1 = '1') then
          o_label6_data1 <= f32_data ;
        end if;
        if (w_load_label6_data0 = '1') then
          o_label6_data0 <= f32_data ;
        end if;
        if (w_load_label7_config = '1') then
          o_label7_config(7 downto 0) <= f32_data(7 downto 0) ;
        end if;
        if (w_load_label7_config = '1') then
          o_label7_config(8 downto 8) <= f32_data(8 downto 8) ;
        end if;
        if (w_load_label7_config = '1') then
          o_label7_config(14 downto 9) <= f32_data(30 downto 25) ;
        end if;
        if (w_load_label7_config = '1') then
          o_label7_config(15 downto 15) <= f32_data(31 downto 31) ;
        end if;
        if (w_load_label7_data7 = '1') then
          o_label7_data7 <= f32_data ;
        end if;
        if (w_load_label7_data6 = '1') then
          o_label7_data6 <= f32_data ;
        end if;
        if (w_load_label7_data5 = '1') then
          o_label7_data5 <= f32_data ;
        end if;
        if (w_load_label7_data4 = '1') then
          o_label7_data4 <= f32_data ;
        end if;
        if (w_load_label7_data3 = '1') then
          o_label7_data3 <= f32_data ;
        end if;
        if (w_load_label7_data2 = '1') then
          o_label7_data2 <= f32_data ;
        end if;
        if (w_load_label7_data1 = '1') then
          o_label7_data1 <= f32_data ;
        end if;
        if (w_load_label7_data0 = '1') then
          o_label7_data0 <= f32_data ;
        end if;
        if (w_load_kdf_drbg_ctrl = '1') then
          o_kdf_drbg_ctrl <= f32_data(1 downto 0) ;
        end if;
        if (w_load_kdf_drbg_seed_0_state_key_31_0 = '1') then
          o_kdf_drbg_seed_0_state_key_31_0 <= f32_data ;
        end if;
        if (w_load_kdf_drbg_seed_0_state_key_63_32 = '1') then
          o_kdf_drbg_seed_0_state_key_63_32 <= f32_data ;
        end if;
        if (w_load_kdf_drbg_seed_0_state_key_95_64 = '1') then
          o_kdf_drbg_seed_0_state_key_95_64 <= f32_data ;
        end if;
        if (w_load_kdf_drbg_seed_0_state_key_127_96 = '1') then
          o_kdf_drbg_seed_0_state_key_127_96 <= f32_data ;
        end if;
        if (w_load_kdf_drbg_seed_0_state_key_159_128 = '1') then
          o_kdf_drbg_seed_0_state_key_159_128 <= f32_data ;
        end if;
        if (w_load_kdf_drbg_seed_0_state_key_191_160 = '1') then
          o_kdf_drbg_seed_0_state_key_191_160 <= f32_data ;
        end if;
        if (w_load_kdf_drbg_seed_0_state_key_223_192 = '1') then
          o_kdf_drbg_seed_0_state_key_223_192 <= f32_data ;
        end if;
        if (w_load_kdf_drbg_seed_0_state_key_255_224 = '1') then
          o_kdf_drbg_seed_0_state_key_255_224 <= f32_data ;
        end if;
        if (w_load_kdf_drbg_seed_0_state_value_31_0 = '1') then
          o_kdf_drbg_seed_0_state_value_31_0 <= f32_data ;
        end if;
        if (w_load_kdf_drbg_seed_0_state_value_63_32 = '1') then
          o_kdf_drbg_seed_0_state_value_63_32 <= f32_data ;
        end if;
        if (w_load_kdf_drbg_seed_0_state_value_95_64 = '1') then
          o_kdf_drbg_seed_0_state_value_95_64 <= f32_data ;
        end if;
        if (w_load_kdf_drbg_seed_0_state_value_127_96 = '1') then
          o_kdf_drbg_seed_0_state_value_127_96 <= f32_data ;
        end if;
        if (w_load_kdf_drbg_seed_0_reseed_interval_0 = '1') then
          o_kdf_drbg_seed_0_reseed_interval_0 <= f32_data ;
        end if;
        if (w_load_kdf_drbg_seed_0_reseed_interval_1 = '1') then
          o_kdf_drbg_seed_0_reseed_interval_1 <= f32_data(15 downto 0) ;
        end if;
        if (w_load_kdf_drbg_seed_1_state_key_31_0 = '1') then
          o_kdf_drbg_seed_1_state_key_31_0 <= f32_data ;
        end if;
        if (w_load_kdf_drbg_seed_1_state_key_63_32 = '1') then
          o_kdf_drbg_seed_1_state_key_63_32 <= f32_data ;
        end if;
        if (w_load_kdf_drbg_seed_1_state_key_95_64 = '1') then
          o_kdf_drbg_seed_1_state_key_95_64 <= f32_data ;
        end if;
        if (w_load_kdf_drbg_seed_1_state_key_127_96 = '1') then
          o_kdf_drbg_seed_1_state_key_127_96 <= f32_data ;
        end if;
        if (w_load_kdf_drbg_seed_1_state_key_159_128 = '1') then
          o_kdf_drbg_seed_1_state_key_159_128 <= f32_data ;
        end if;
        if (w_load_kdf_drbg_seed_1_state_key_191_160 = '1') then
          o_kdf_drbg_seed_1_state_key_191_160 <= f32_data ;
        end if;
        if (w_load_kdf_drbg_seed_1_state_key_223_192 = '1') then
          o_kdf_drbg_seed_1_state_key_223_192 <= f32_data ;
        end if;
        if (w_load_kdf_drbg_seed_1_state_key_255_224 = '1') then
          o_kdf_drbg_seed_1_state_key_255_224 <= f32_data ;
        end if;
        if (w_load_kdf_drbg_seed_1_state_value_31_0 = '1') then
          o_kdf_drbg_seed_1_state_value_31_0 <= f32_data ;
        end if;
        if (w_load_kdf_drbg_seed_1_state_value_63_32 = '1') then
          o_kdf_drbg_seed_1_state_value_63_32 <= f32_data ;
        end if;
        if (w_load_kdf_drbg_seed_1_state_value_95_64 = '1') then
          o_kdf_drbg_seed_1_state_value_95_64 <= f32_data ;
        end if;
        if (w_load_kdf_drbg_seed_1_state_value_127_96 = '1') then
          o_kdf_drbg_seed_1_state_value_127_96 <= f32_data ;
        end if;
        if (w_load_kdf_drbg_seed_1_reseed_interval_0 = '1') then
          o_kdf_drbg_seed_1_reseed_interval_0 <= f32_data ;
        end if;
        if (w_load_kdf_drbg_seed_1_reseed_interval_1 = '1') then
          o_kdf_drbg_seed_1_reseed_interval_1 <= f32_data(15 downto 0) ;
        end if;
        if (w_load_interrupt_status = '1') then
          o_interrupt_status(0 downto 0) <= f32_data(0 downto 0) ;
        end if;
        if (w_load_interrupt_status = '1') then
          o_interrupt_status(1 downto 1) <= f32_data(1 downto 1) ;
        end if;
        if (w_load_interrupt_status = '1') then
          o_interrupt_status(2 downto 2) <= f32_data(2 downto 2) ;
        end if;
        if (w_load_interrupt_status = '1') then
          o_interrupt_status(3 downto 3) <= f32_data(3 downto 3) ;
        end if;
        if (w_load_interrupt_status = '1') then
          o_interrupt_status(4 downto 4) <= f32_data(4 downto 4) ;
        end if;
        if (w_load_interrupt_mask = '1') then
          o_interrupt_mask(0 downto 0) <= f32_data(0 downto 0) ;
        end if;
        if (w_load_interrupt_mask = '1') then
          o_interrupt_mask(1 downto 1) <= f32_data(1 downto 1) ;
        end if;
        if (w_load_interrupt_mask = '1') then
          o_interrupt_mask(2 downto 2) <= f32_data(2 downto 2) ;
        end if;
        if (w_load_interrupt_mask = '1') then
          o_interrupt_mask(3 downto 3) <= f32_data(3 downto 3) ;
        end if;
        if (w_load_interrupt_mask = '1') then
          o_interrupt_mask(4 downto 4) <= f32_data(4 downto 4) ;
        end if;
        if (w_load_engine_sticky_status = '1') then
          o_engine_sticky_status(0 downto 0) <= f32_data(0 downto 0) ;
        end if;
        if (w_load_engine_sticky_status = '1') then
          o_engine_sticky_status(1 downto 1) <= f32_data(1 downto 1) ;
        end if;
        if (w_load_engine_sticky_status = '1') then
          o_engine_sticky_status(2 downto 2) <= f32_data(2 downto 2) ;
        end if;
        if (w_load_engine_sticky_status = '1') then
          o_engine_sticky_status(3 downto 3) <= f32_data(3 downto 3) ;
        end if;
        if (w_load_engine_sticky_status = '1') then
          o_engine_sticky_status(4 downto 4) <= f32_data(4 downto 4) ;
        end if;
        if (w_load_engine_sticky_status = '1') then
          o_engine_sticky_status(5 downto 5) <= f32_data(5 downto 5) ;
        end if;
        if (w_load_engine_sticky_status = '1') then
          o_engine_sticky_status(6 downto 6) <= f32_data(6 downto 6) ;
        end if;
        if (w_load_engine_sticky_status = '1') then
          o_engine_sticky_status(7 downto 7) <= f32_data(7 downto 7) ;
        end if;
        if (w_load_bimc_monitor_mask = '1') then
          o_bimc_monitor_mask(0 downto 0) <= f32_data(0 downto 0) ;
        end if;
        if (w_load_bimc_monitor_mask = '1') then
          o_bimc_monitor_mask(1 downto 1) <= f32_data(1 downto 1) ;
        end if;
        if (w_load_bimc_monitor_mask = '1') then
          o_bimc_monitor_mask(2 downto 2) <= f32_data(2 downto 2) ;
        end if;
        if (w_load_bimc_monitor_mask = '1') then
          o_bimc_monitor_mask(3 downto 3) <= f32_data(3 downto 3) ;
        end if;
        if (w_load_bimc_monitor_mask = '1') then
          o_bimc_monitor_mask(4 downto 4) <= f32_data(4 downto 4) ;
        end if;
        if (w_load_bimc_monitor_mask = '1') then
          o_bimc_monitor_mask(5 downto 5) <= f32_data(5 downto 5) ;
        end if;
        if (w_load_bimc_monitor_mask = '1') then
          o_bimc_monitor_mask(6 downto 6) <= f32_data(6 downto 6) ;
        end if;
        if (w_load_bimc_ecc_uncorrectable_error_cnt = '1') then
          o_bimc_ecc_uncorrectable_error_cnt <= f32_data ;
        end if;
        if (w_load_bimc_ecc_correctable_error_cnt = '1') then
          o_bimc_ecc_correctable_error_cnt <= f32_data ;
        end if;
        if (w_load_bimc_parity_error_cnt = '1') then
          o_bimc_parity_error_cnt <= f32_data ;
        end if;
        if (w_load_bimc_global_config = '1') then
          o_bimc_global_config(0 downto 0) <= f32_data(0 downto 0) ;
        end if;
        if (w_load_bimc_global_config = '1') then
          o_bimc_global_config(1 downto 1) <= f32_data(1 downto 1) ;
        end if;
        if (w_load_bimc_global_config = '1') then
          o_bimc_global_config(2 downto 2) <= f32_data(2 downto 2) ;
        end if;
        if (w_load_bimc_global_config = '1') then
          o_bimc_global_config(3 downto 3) <= f32_data(3 downto 3) ;
        end if;
        if (w_load_bimc_global_config = '1') then
          o_bimc_global_config(4 downto 4) <= f32_data(4 downto 4) ;
        end if;
        if (w_load_bimc_global_config = '1') then
          o_bimc_global_config(5 downto 5) <= f32_data(5 downto 5) ;
        end if;
        if (w_load_bimc_global_config = '1') then
          o_bimc_global_config(31 downto 6) <= f32_data(31 downto 6) ;
        end if;
        if (w_load_bimc_eccpar_debug = '1') then
          o_bimc_eccpar_debug(11 downto 0) <= f32_data(11 downto 0) ;
        end if;
        if (w_load_bimc_eccpar_debug = '1') then
          o_bimc_eccpar_debug(15 downto 12) <= f32_data(15 downto 12) ;
        end if;
        if (w_load_bimc_eccpar_debug = '1') then
          o_bimc_eccpar_debug(17 downto 16) <= f32_data(17 downto 16) ;
        end if;
        if (w_load_bimc_eccpar_debug = '1') then
          o_bimc_eccpar_debug(19 downto 18) <= f32_data(19 downto 18) ;
        end if;
        if (w_load_bimc_eccpar_debug = '1') then
          o_bimc_eccpar_debug(21 downto 20) <= f32_data(21 downto 20) ;
        end if;
        if (w_load_bimc_eccpar_debug = '1') then
          o_bimc_eccpar_debug(22 downto 22) <= f32_data(22 downto 22) ;
        end if;
        if (w_load_bimc_eccpar_debug = '1') then
          o_bimc_eccpar_debug(23 downto 23) <= f32_data(23 downto 23) ;
        end if;
        if (w_load_bimc_eccpar_debug = '1') then
          o_bimc_eccpar_debug(27 downto 24) <= f32_data(27 downto 24) ;
        end if;
        if (w_load_bimc_eccpar_debug = '1') then
          o_bimc_eccpar_debug(28 downto 28) <= f32_data(28 downto 28) ;
        end if;
        if (w_load_bimc_cmd2 = '1') then
          o_bimc_cmd2(7 downto 0) <= f32_data(7 downto 0) ;
        end if;
        if (w_load_bimc_cmd2 = '1') then
          o_bimc_cmd2(8 downto 8) <= f32_data(8 downto 8) ;
        end if;
        if (w_load_bimc_cmd2 = '1') then
          o_bimc_cmd2(9 downto 9) <= f32_data(9 downto 9) ;
        end if;
        if (w_load_bimc_cmd2 = '1') then
          o_bimc_cmd2(10 downto 10) <= f32_data(10 downto 10) ;
        end if;
        if (w_load_bimc_cmd1 = '1') then
          o_bimc_cmd1(15 downto 0) <= f32_data(15 downto 0) ;
        end if;
        if (w_load_bimc_cmd1 = '1') then
          o_bimc_cmd1(27 downto 16) <= f32_data(27 downto 16) ;
        end if;
        if (w_load_bimc_cmd1 = '1') then
          o_bimc_cmd1(31 downto 28) <= f32_data(31 downto 28) ;
        end if;
        if (w_load_bimc_cmd0 = '1') then
          o_bimc_cmd0 <= f32_data ;
        end if;
        if (w_load_bimc_rxcmd2 = '1') then
          o_bimc_rxcmd2(7 downto 0) <= f32_data(7 downto 0) ;
        end if;
        if (w_load_bimc_rxcmd2 = '1') then
          o_bimc_rxcmd2(8 downto 8) <= f32_data(8 downto 8) ;
        end if;
        if (w_load_bimc_rxrsp2 = '1') then
          o_bimc_rxrsp2(7 downto 0) <= f32_data(7 downto 0) ;
        end if;
        if (w_load_bimc_rxrsp2 = '1') then
          o_bimc_rxrsp2(8 downto 8) <= f32_data(8 downto 8) ;
        end if;
        if (w_load_bimc_pollrsp2 = '1') then
          o_bimc_pollrsp2(7 downto 0) <= f32_data(7 downto 0) ;
        end if;
        if (w_load_bimc_pollrsp2 = '1') then
          o_bimc_pollrsp2(8 downto 8) <= f32_data(8 downto 8) ;
        end if;
        if (w_load_bimc_dbgcmd2 = '1') then
          o_bimc_dbgcmd2(7 downto 0) <= f32_data(7 downto 0) ;
        end if;
        if (w_load_bimc_dbgcmd2 = '1') then
          o_bimc_dbgcmd2(8 downto 8) <= f32_data(8 downto 8) ;
        end if;
        if (w_load_im_consumed = '1') then
          o_im_consumed(0 downto 0) <= f32_data(0 downto 0) ;
        end if;
        if (w_load_im_consumed = '1') then
          o_im_consumed(1 downto 1) <= f32_data(1 downto 1) ;
        end if;
        if (w_load_im_consumed = '1') then
          o_im_consumed(2 downto 2) <= f32_data(2 downto 2) ;
        end if;
        if (w_load_im_consumed = '1') then
          o_im_consumed(3 downto 3) <= f32_data(3 downto 3) ;
        end if;
        if (w_load_im_consumed = '1') then
          o_im_consumed(4 downto 4) <= f32_data(4 downto 4) ;
        end if;
        if (w_load_im_consumed = '1') then
          o_im_consumed(5 downto 5) <= f32_data(5 downto 5) ;
        end if;
        if (w_load_im_consumed = '1') then
          o_im_consumed(6 downto 6) <= f32_data(6 downto 6) ;
        end if;
        if (w_load_im_consumed = '1') then
          o_im_consumed(7 downto 7) <= f32_data(7 downto 7) ;
        end if;
        if (w_load_im_consumed = '1') then
          o_im_consumed(8 downto 8) <= f32_data(8 downto 8) ;
        end if;
        if (w_load_im_consumed = '1') then
          o_im_consumed(9 downto 9) <= f32_data(9 downto 9) ;
        end if;
        if (w_load_im_consumed = '1') then
          o_im_consumed(10 downto 10) <= f32_data(10 downto 10) ;
        end if;
        if (w_load_im_consumed = '1') then
          o_im_consumed(11 downto 11) <= f32_data(11 downto 11) ;
        end if;
        if (w_load_im_consumed = '1') then
          o_im_consumed(12 downto 12) <= f32_data(12 downto 12) ;
        end if;
        if (w_load_im_consumed = '1') then
          o_im_consumed(13 downto 13) <= f32_data(13 downto 13) ;
        end if;
        if (w_load_im_consumed = '1') then
          o_im_consumed(14 downto 14) <= f32_data(14 downto 14) ;
        end if;
        if (w_load_im_consumed = '1') then
          o_im_consumed(15 downto 15) <= f32_data(15 downto 15) ;
        end if;
        if (w_load_tready_override = '1') then
          o_tready_override(0 downto 0) <= f32_data(0 downto 0) ;
        end if;
        if (w_load_tready_override = '1') then
          o_tready_override(1 downto 1) <= f32_data(1 downto 1) ;
        end if;
        if (w_load_tready_override = '1') then
          o_tready_override(2 downto 2) <= f32_data(2 downto 2) ;
        end if;
        if (w_load_tready_override = '1') then
          o_tready_override(3 downto 3) <= f32_data(3 downto 3) ;
        end if;
        if (w_load_tready_override = '1') then
          o_tready_override(4 downto 4) <= f32_data(4 downto 4) ;
        end if;
        if (w_load_tready_override = '1') then
          o_tready_override(5 downto 5) <= f32_data(5 downto 5) ;
        end if;
        if (w_load_tready_override = '1') then
          o_tready_override(6 downto 6) <= f32_data(6 downto 6) ;
        end if;
        if (w_load_tready_override = '1') then
          o_tready_override(7 downto 7) <= f32_data(7 downto 7) ;
        end if;
        if (w_load_tready_override = '1') then
          o_tready_override(8 downto 8) <= f32_data(8 downto 8) ;
        end if;
        if (w_load_regs_sa_ctrl = '1') then
          o_regs_sa_ctrl(0 downto 0) <= f32_data(0 downto 0) ;
        end if;
        if (w_load_regs_sa_ctrl = '1') then
          o_regs_sa_ctrl(1 downto 1) <= f32_data(1 downto 1) ;
        end if;
        if (w_load_regs_sa_ctrl = '1') then
          o_regs_sa_ctrl(7 downto 2) <= f32_data(7 downto 2) ;
        end if;
        if (w_load_regs_sa_ctrl = '1') then
          o_regs_sa_ctrl(12 downto 8) <= f32_data(12 downto 8) ;
        end if;
        if (w_load_regs_sa_ctrl = '1') then
          o_regs_sa_ctrl(31 downto 13) <= f32_data(31 downto 13) ;
        end if;
        if (w_load_sa_snapshot_ia_wdata_part0 = '1') then
          o_sa_snapshot_ia_wdata_part0(17 downto 0) <= f32_data(17 downto 0) ;
        end if;
        if (w_load_sa_snapshot_ia_wdata_part0 = '1') then
          o_sa_snapshot_ia_wdata_part0(31 downto 18) <= f32_data(31 downto 18) ;
        end if;
        if (w_load_sa_snapshot_ia_wdata_part1 = '1') then
          o_sa_snapshot_ia_wdata_part1 <= f32_data ;
        end if;
        if (w_load_sa_snapshot_ia_config = '1') then
          o_sa_snapshot_ia_config(4 downto 0) <= f32_data(4 downto 0) ;
        end if;
        if (w_load_sa_snapshot_ia_config = '1') then
          o_sa_snapshot_ia_config(8 downto 5) <= f32_data(31 downto 28) ;
        end if;
        if (w_load_sa_count_ia_wdata_part0 = '1') then
          o_sa_count_ia_wdata_part0(17 downto 0) <= f32_data(17 downto 0) ;
        end if;
        if (w_load_sa_count_ia_wdata_part0 = '1') then
          o_sa_count_ia_wdata_part0(31 downto 18) <= f32_data(31 downto 18) ;
        end if;
        if (w_load_sa_count_ia_wdata_part1 = '1') then
          o_sa_count_ia_wdata_part1 <= f32_data ;
        end if;
        if (w_load_sa_count_ia_config = '1') then
          o_sa_count_ia_config(4 downto 0) <= f32_data(4 downto 0) ;
        end if;
        if (w_load_sa_count_ia_config = '1') then
          o_sa_count_ia_config(8 downto 5) <= f32_data(31 downto 28) ;
        end if;
        if (w_load_cceip_encrypt_kop_fifo_override = '1') then
          o_cceip_encrypt_kop_fifo_override(0 downto 0) <= f32_data(0 downto 0)
           ;
        end if;
        if (w_load_cceip_encrypt_kop_fifo_override = '1') then
          o_cceip_encrypt_kop_fifo_override(1 downto 1) <= f32_data(1 downto 1)
           ;
        end if;
        if (w_load_cceip_encrypt_kop_fifo_override = '1') then
          o_cceip_encrypt_kop_fifo_override(2 downto 2) <= f32_data(2 downto 2)
           ;
        end if;
        if (w_load_cceip_encrypt_kop_fifo_override = '1') then
          o_cceip_encrypt_kop_fifo_override(3 downto 3) <= f32_data(3 downto 3)
           ;
        end if;
        if (w_load_cceip_encrypt_kop_fifo_override = '1') then
          o_cceip_encrypt_kop_fifo_override(4 downto 4) <= f32_data(4 downto 4)
           ;
        end if;
        if (w_load_cceip_encrypt_kop_fifo_override = '1') then
          o_cceip_encrypt_kop_fifo_override(5 downto 5) <= f32_data(5 downto 5)
           ;
        end if;
        if (w_load_cceip_encrypt_kop_fifo_override = '1') then
          o_cceip_encrypt_kop_fifo_override(6 downto 6) <= f32_data(6 downto 6)
           ;
        end if;
        if (w_load_cceip_validate_kop_fifo_override = '1') then
          o_cceip_validate_kop_fifo_override(0 downto 0) <= f32_data(0 downto 0)
           ;
        end if;
        if (w_load_cceip_validate_kop_fifo_override = '1') then
          o_cceip_validate_kop_fifo_override(1 downto 1) <= f32_data(1 downto 1)
           ;
        end if;
        if (w_load_cceip_validate_kop_fifo_override = '1') then
          o_cceip_validate_kop_fifo_override(2 downto 2) <= f32_data(2 downto 2)
           ;
        end if;
        if (w_load_cceip_validate_kop_fifo_override = '1') then
          o_cceip_validate_kop_fifo_override(3 downto 3) <= f32_data(3 downto 3)
           ;
        end if;
        if (w_load_cceip_validate_kop_fifo_override = '1') then
          o_cceip_validate_kop_fifo_override(4 downto 4) <= f32_data(4 downto 4)
           ;
        end if;
        if (w_load_cceip_validate_kop_fifo_override = '1') then
          o_cceip_validate_kop_fifo_override(5 downto 5) <= f32_data(5 downto 5)
           ;
        end if;
        if (w_load_cceip_validate_kop_fifo_override = '1') then
          o_cceip_validate_kop_fifo_override(6 downto 6) <= f32_data(6 downto 6)
           ;
        end if;
        if (w_load_cddip_decrypt_kop_fifo_override = '1') then
          o_cddip_decrypt_kop_fifo_override(0 downto 0) <= f32_data(0 downto 0)
           ;
        end if;
        if (w_load_cddip_decrypt_kop_fifo_override = '1') then
          o_cddip_decrypt_kop_fifo_override(1 downto 1) <= f32_data(1 downto 1)
           ;
        end if;
        if (w_load_cddip_decrypt_kop_fifo_override = '1') then
          o_cddip_decrypt_kop_fifo_override(2 downto 2) <= f32_data(2 downto 2)
           ;
        end if;
        if (w_load_cddip_decrypt_kop_fifo_override = '1') then
          o_cddip_decrypt_kop_fifo_override(3 downto 3) <= f32_data(3 downto 3)
           ;
        end if;
        if (w_load_cddip_decrypt_kop_fifo_override = '1') then
          o_cddip_decrypt_kop_fifo_override(4 downto 4) <= f32_data(4 downto 4)
           ;
        end if;
        if (w_load_cddip_decrypt_kop_fifo_override = '1') then
          o_cddip_decrypt_kop_fifo_override(5 downto 5) <= f32_data(5 downto 5)
           ;
        end if;
        if (w_load_cddip_decrypt_kop_fifo_override = '1') then
          o_cddip_decrypt_kop_fifo_override(6 downto 6) <= f32_data(6 downto 6)
           ;
        end if;
        if (w_load_sa_global_ctrl = '1') then
          o_sa_global_ctrl(0 downto 0) <= f32_data(0 downto 0) ;
        end if;
        if (w_load_sa_global_ctrl = '1') then
          o_sa_global_ctrl(1 downto 1) <= f32_data(1 downto 1) ;
        end if;
        if (w_load_sa_global_ctrl = '1') then
          o_sa_global_ctrl(31 downto 2) <= f32_data(31 downto 2) ;
        end if;
        if (w_load_sa_ctrl_ia_wdata_part0 = '1') then
          o_sa_ctrl_ia_wdata_part0(4 downto 0) <= f32_data(4 downto 0) ;
        end if;
        if (w_load_sa_ctrl_ia_wdata_part0 = '1') then
          o_sa_ctrl_ia_wdata_part0(31 downto 5) <= f32_data(31 downto 5) ;
        end if;
        if (w_load_sa_ctrl_ia_config = '1') then
          o_sa_ctrl_ia_config(4 downto 0) <= f32_data(4 downto 0) ;
        end if;
        if (w_load_sa_ctrl_ia_config = '1') then
          o_sa_ctrl_ia_config(8 downto 5) <= f32_data(31 downto 28) ;
        end if;
        if (w_load_kdf_test_key_size_config = '1') then
          o_kdf_test_key_size_config <= f32_data ;
        end if;
      end if;
    end if ;
  end process ;

  process --:o1787
  (clk)
  begin
    if (clk'event and clk = '1') then
      if (w_load_cceip0_out_ia_wdata_part0 = '1') then
        o_cceip0_out_ia_wdata_part0(13 downto 6) <= f32_data(13 downto 6) ;
      end if;
      if (w_load_cceip0_out_ia_wdata_part0 = '1') then
        o_cceip0_out_ia_wdata_part0(14 downto 14) <= f32_data(14 downto 14) ;
      end if;
      if (w_load_cceip0_out_ia_wdata_part0 = '1') then
        o_cceip0_out_ia_wdata_part0(22 downto 15) <= f32_data(22 downto 15) ;
      end if;
      if (w_load_cceip0_out_ia_wdata_part0 = '1') then
        o_cceip0_out_ia_wdata_part0(30 downto 23) <= f32_data(30 downto 23) ;
      end if;
      if (w_load_cceip0_out_ia_wdata_part0 = '1') then
        o_cceip0_out_ia_wdata_part0(31 downto 31) <= f32_data(31 downto 31) ;
      end if;
      if (w_load_cceip1_out_ia_wdata_part0 = '1') then
        o_cceip1_out_ia_wdata_part0(13 downto 6) <= f32_data(13 downto 6) ;
      end if;
      if (w_load_cceip1_out_ia_wdata_part0 = '1') then
        o_cceip1_out_ia_wdata_part0(14 downto 14) <= f32_data(14 downto 14) ;
      end if;
      if (w_load_cceip1_out_ia_wdata_part0 = '1') then
        o_cceip1_out_ia_wdata_part0(22 downto 15) <= f32_data(22 downto 15) ;
      end if;
      if (w_load_cceip1_out_ia_wdata_part0 = '1') then
        o_cceip1_out_ia_wdata_part0(30 downto 23) <= f32_data(30 downto 23) ;
      end if;
      if (w_load_cceip1_out_ia_wdata_part0 = '1') then
        o_cceip1_out_ia_wdata_part0(31 downto 31) <= f32_data(31 downto 31) ;
      end if;
      if (w_load_cceip2_out_ia_wdata_part0 = '1') then
        o_cceip2_out_ia_wdata_part0(13 downto 6) <= f32_data(13 downto 6) ;
      end if;
      if (w_load_cceip2_out_ia_wdata_part0 = '1') then
        o_cceip2_out_ia_wdata_part0(14 downto 14) <= f32_data(14 downto 14) ;
      end if;
      if (w_load_cceip2_out_ia_wdata_part0 = '1') then
        o_cceip2_out_ia_wdata_part0(22 downto 15) <= f32_data(22 downto 15) ;
      end if;
      if (w_load_cceip2_out_ia_wdata_part0 = '1') then
        o_cceip2_out_ia_wdata_part0(30 downto 23) <= f32_data(30 downto 23) ;
      end if;
      if (w_load_cceip2_out_ia_wdata_part0 = '1') then
        o_cceip2_out_ia_wdata_part0(31 downto 31) <= f32_data(31 downto 31) ;
      end if;
      if (w_load_cceip3_out_ia_wdata_part0 = '1') then
        o_cceip3_out_ia_wdata_part0(13 downto 6) <= f32_data(13 downto 6) ;
      end if;
      if (w_load_cceip3_out_ia_wdata_part0 = '1') then
        o_cceip3_out_ia_wdata_part0(14 downto 14) <= f32_data(14 downto 14) ;
      end if;
      if (w_load_cceip3_out_ia_wdata_part0 = '1') then
        o_cceip3_out_ia_wdata_part0(22 downto 15) <= f32_data(22 downto 15) ;
      end if;
      if (w_load_cceip3_out_ia_wdata_part0 = '1') then
        o_cceip3_out_ia_wdata_part0(30 downto 23) <= f32_data(30 downto 23) ;
      end if;
      if (w_load_cceip3_out_ia_wdata_part0 = '1') then
        o_cceip3_out_ia_wdata_part0(31 downto 31) <= f32_data(31 downto 31) ;
      end if;
      if (w_load_cddip0_out_ia_wdata_part0 = '1') then
        o_cddip0_out_ia_wdata_part0(13 downto 6) <= f32_data(13 downto 6) ;
      end if;
      if (w_load_cddip0_out_ia_wdata_part0 = '1') then
        o_cddip0_out_ia_wdata_part0(14 downto 14) <= f32_data(14 downto 14) ;
      end if;
      if (w_load_cddip0_out_ia_wdata_part0 = '1') then
        o_cddip0_out_ia_wdata_part0(22 downto 15) <= f32_data(22 downto 15) ;
      end if;
      if (w_load_cddip0_out_ia_wdata_part0 = '1') then
        o_cddip0_out_ia_wdata_part0(30 downto 23) <= f32_data(30 downto 23) ;
      end if;
      if (w_load_cddip0_out_ia_wdata_part0 = '1') then
        o_cddip0_out_ia_wdata_part0(31 downto 31) <= f32_data(31 downto 31) ;
      end if;
      if (w_load_cddip1_out_ia_wdata_part0 = '1') then
        o_cddip1_out_ia_wdata_part0(13 downto 6) <= f32_data(13 downto 6) ;
      end if;
      if (w_load_cddip1_out_ia_wdata_part0 = '1') then
        o_cddip1_out_ia_wdata_part0(14 downto 14) <= f32_data(14 downto 14) ;
      end if;
      if (w_load_cddip1_out_ia_wdata_part0 = '1') then
        o_cddip1_out_ia_wdata_part0(22 downto 15) <= f32_data(22 downto 15) ;
      end if;
      if (w_load_cddip1_out_ia_wdata_part0 = '1') then
        o_cddip1_out_ia_wdata_part0(30 downto 23) <= f32_data(30 downto 23) ;
      end if;
      if (w_load_cddip1_out_ia_wdata_part0 = '1') then
        o_cddip1_out_ia_wdata_part0(31 downto 31) <= f32_data(31 downto 31) ;
      end if;
      if (w_load_cddip2_out_ia_wdata_part0 = '1') then
        o_cddip2_out_ia_wdata_part0(13 downto 6) <= f32_data(13 downto 6) ;
      end if;
      if (w_load_cddip2_out_ia_wdata_part0 = '1') then
        o_cddip2_out_ia_wdata_part0(14 downto 14) <= f32_data(14 downto 14) ;
      end if;
      if (w_load_cddip2_out_ia_wdata_part0 = '1') then
        o_cddip2_out_ia_wdata_part0(22 downto 15) <= f32_data(22 downto 15) ;
      end if;
      if (w_load_cddip2_out_ia_wdata_part0 = '1') then
        o_cddip2_out_ia_wdata_part0(30 downto 23) <= f32_data(30 downto 23) ;
      end if;
      if (w_load_cddip2_out_ia_wdata_part0 = '1') then
        o_cddip2_out_ia_wdata_part0(31 downto 31) <= f32_data(31 downto 31) ;
      end if;
      if (w_load_cddip3_out_ia_wdata_part0 = '1') then
        o_cddip3_out_ia_wdata_part0(13 downto 6) <= f32_data(13 downto 6) ;
      end if;
      if (w_load_cddip3_out_ia_wdata_part0 = '1') then
        o_cddip3_out_ia_wdata_part0(14 downto 14) <= f32_data(14 downto 14) ;
      end if;
      if (w_load_cddip3_out_ia_wdata_part0 = '1') then
        o_cddip3_out_ia_wdata_part0(22 downto 15) <= f32_data(22 downto 15) ;
      end if;
      if (w_load_cddip3_out_ia_wdata_part0 = '1') then
        o_cddip3_out_ia_wdata_part0(30 downto 23) <= f32_data(30 downto 23) ;
      end if;
      if (w_load_cddip3_out_ia_wdata_part0 = '1') then
        o_cddip3_out_ia_wdata_part0(31 downto 31) <= f32_data(31 downto 31) ;
      end if;
      if (w_load_bimc_rxcmd2 = '1') then
        o_bimc_rxcmd2(9 downto 9) <= f32_data(9 downto 9) ;
      end if;
      if (w_load_bimc_rxrsp2 = '1') then
        o_bimc_rxrsp2(9 downto 9) <= f32_data(9 downto 9) ;
      end if;
      if (w_load_bimc_pollrsp2 = '1') then
        o_bimc_pollrsp2(9 downto 9) <= f32_data(9 downto 9) ;
      end if;
      if (w_load_bimc_dbgcmd2 = '1') then
        o_bimc_dbgcmd2(9 downto 9) <= f32_data(9 downto 9) ;
      end if;
    end if ;
  end process ;
end module;
