// xc_work/v/144.sv
// /lan/cva_rel/ixcom23h1/23.03.131.s001/tools.lnx86/etc/ixcom/GFIFO.sv:89
// NOTE: This file corresponds to a module in the Hardware/DUT partition.
`timescale 1ps/1ps
module IXC_SV_GFIFO(input  [63:0] rdCnt );
IXC_SV_GFIFO_VXE_256 O(rdCnt); 
// pragma CVASTRPROP MODULE IXC_SV_GFIFO PROP_IXCOM_MOD TRUE
endmodule

